VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_08_sws
  CLASS BLOCK ;
  FOREIGN tt_um_08_sws ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    ANTENNAGATEAREA 200.000000 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    ANTENNAGATEAREA 550.000000 ;
    ANTENNADIFFAREA 2.900000 ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    ANTENNAGATEAREA 550.000000 ;
    ANTENNADIFFAREA 2.900000 ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    ANTENNADIFFAREA 29.000000 ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    ANTENNADIFFAREA 29.000000 ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    ANTENNAGATEAREA 918.296448 ;
    ANTENNADIFFAREA 1107.646118 ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 14.805 211.185 14.975 211.375 ;
        RECT 18.485 211.185 18.655 211.375 ;
        RECT 24.005 211.185 24.175 211.375 ;
        RECT 25.845 211.185 26.015 211.375 ;
        RECT 31.365 211.185 31.535 211.375 ;
        RECT 36.885 211.185 37.055 211.375 ;
        RECT 38.725 211.185 38.895 211.375 ;
        RECT 44.245 211.185 44.415 211.375 ;
        RECT 49.765 211.185 49.935 211.375 ;
        RECT 51.605 211.185 51.775 211.375 ;
        RECT 57.125 211.185 57.295 211.375 ;
        RECT 62.645 211.185 62.815 211.375 ;
        RECT 64.485 211.185 64.655 211.375 ;
        RECT 70.005 211.185 70.175 211.375 ;
        RECT 75.525 211.185 75.695 211.375 ;
        RECT 77.365 211.185 77.535 211.375 ;
        RECT 82.885 211.185 83.055 211.375 ;
        RECT 88.405 211.185 88.575 211.375 ;
        RECT 90.245 211.185 90.415 211.375 ;
        RECT 95.765 211.185 95.935 211.375 ;
        RECT 101.285 211.185 101.455 211.375 ;
        RECT 103.125 211.185 103.295 211.375 ;
        RECT 108.645 211.185 108.815 211.375 ;
        RECT 114.165 211.185 114.335 211.375 ;
        RECT 115.140 211.235 115.260 211.345 ;
        RECT 120.605 211.185 120.775 211.375 ;
        RECT 126.125 211.185 126.295 211.375 ;
        RECT 127.505 211.185 127.675 211.375 ;
        RECT 14.665 210.375 16.035 211.185 ;
        RECT 16.045 210.375 18.795 211.185 ;
        RECT 18.805 210.375 24.315 211.185 ;
        RECT 24.335 210.315 24.765 211.100 ;
        RECT 24.785 210.375 26.155 211.185 ;
        RECT 26.165 210.375 31.675 211.185 ;
        RECT 31.685 210.375 37.195 211.185 ;
        RECT 37.215 210.315 37.645 211.100 ;
        RECT 37.665 210.375 39.035 211.185 ;
        RECT 39.045 210.375 44.555 211.185 ;
        RECT 44.565 210.375 50.075 211.185 ;
        RECT 50.095 210.315 50.525 211.100 ;
        RECT 50.545 210.375 51.915 211.185 ;
        RECT 51.925 210.375 57.435 211.185 ;
        RECT 57.445 210.375 62.955 211.185 ;
        RECT 62.975 210.315 63.405 211.100 ;
        RECT 63.425 210.375 64.795 211.185 ;
        RECT 64.805 210.375 70.315 211.185 ;
        RECT 70.325 210.375 75.835 211.185 ;
        RECT 75.855 210.315 76.285 211.100 ;
        RECT 76.305 210.375 77.675 211.185 ;
        RECT 77.685 210.375 83.195 211.185 ;
        RECT 83.205 210.375 88.715 211.185 ;
        RECT 88.735 210.315 89.165 211.100 ;
        RECT 89.185 210.375 90.555 211.185 ;
        RECT 90.565 210.375 96.075 211.185 ;
        RECT 96.085 210.375 101.595 211.185 ;
        RECT 101.615 210.315 102.045 211.100 ;
        RECT 102.065 210.375 103.435 211.185 ;
        RECT 103.445 210.375 108.955 211.185 ;
        RECT 108.965 210.375 114.475 211.185 ;
        RECT 114.495 210.315 114.925 211.100 ;
        RECT 115.405 210.375 120.915 211.185 ;
        RECT 120.925 210.375 126.435 211.185 ;
        RECT 126.445 210.375 127.815 211.185 ;
      LAYER nwell ;
        RECT 14.470 207.155 128.010 209.985 ;
      LAYER pwell ;
        RECT 14.665 205.955 16.035 206.765 ;
        RECT 16.045 205.955 18.795 206.765 ;
        RECT 18.805 205.955 24.315 206.765 ;
        RECT 24.335 206.040 24.765 206.825 ;
        RECT 25.245 205.955 27.995 206.765 ;
        RECT 28.005 205.955 33.515 206.765 ;
        RECT 33.525 205.955 39.035 206.765 ;
        RECT 39.045 205.955 44.555 206.765 ;
        RECT 44.565 205.955 50.075 206.765 ;
        RECT 50.095 206.040 50.525 206.825 ;
        RECT 51.005 205.955 53.755 206.765 ;
        RECT 53.765 205.955 59.275 206.765 ;
        RECT 59.285 205.955 64.795 206.765 ;
        RECT 64.805 205.955 70.315 206.765 ;
        RECT 70.325 205.955 75.835 206.765 ;
        RECT 75.855 206.040 76.285 206.825 ;
        RECT 76.765 205.955 79.515 206.765 ;
        RECT 79.525 205.955 85.035 206.765 ;
        RECT 85.045 205.955 90.555 206.765 ;
        RECT 90.565 205.955 96.075 206.765 ;
        RECT 96.085 205.955 101.595 206.765 ;
        RECT 101.615 206.040 102.045 206.825 ;
        RECT 102.525 205.955 104.355 206.765 ;
        RECT 104.365 205.955 109.875 206.765 ;
        RECT 109.885 205.955 115.395 206.765 ;
        RECT 115.405 205.955 120.915 206.765 ;
        RECT 120.925 205.955 126.435 206.765 ;
        RECT 126.445 205.955 127.815 206.765 ;
        RECT 14.805 205.745 14.975 205.955 ;
        RECT 16.645 205.790 16.805 205.900 ;
        RECT 18.485 205.765 18.655 205.955 ;
        RECT 20.325 205.745 20.495 205.935 ;
        RECT 24.005 205.765 24.175 205.955 ;
        RECT 24.980 205.795 25.100 205.905 ;
        RECT 25.845 205.745 26.015 205.935 ;
        RECT 27.685 205.765 27.855 205.955 ;
        RECT 31.365 205.745 31.535 205.935 ;
        RECT 33.205 205.765 33.375 205.955 ;
        RECT 36.885 205.745 37.055 205.935 ;
        RECT 38.725 205.765 38.895 205.955 ;
        RECT 39.185 205.745 39.355 205.935 ;
        RECT 44.245 205.765 44.415 205.955 ;
        RECT 44.705 205.745 44.875 205.935 ;
        RECT 49.765 205.765 49.935 205.955 ;
        RECT 50.225 205.745 50.395 205.935 ;
        RECT 50.740 205.795 50.860 205.905 ;
        RECT 53.445 205.765 53.615 205.955 ;
        RECT 55.745 205.745 55.915 205.935 ;
        RECT 58.965 205.765 59.135 205.955 ;
        RECT 61.265 205.745 61.435 205.935 ;
        RECT 62.645 205.745 62.815 205.935 ;
        RECT 64.025 205.790 64.185 205.900 ;
        RECT 64.485 205.745 64.655 205.955 ;
        RECT 70.005 205.765 70.175 205.955 ;
        RECT 74.605 205.745 74.775 205.935 ;
        RECT 75.525 205.765 75.695 205.955 ;
        RECT 76.500 205.795 76.620 205.905 ;
        RECT 77.365 205.745 77.535 205.935 ;
        RECT 79.205 205.765 79.375 205.955 ;
        RECT 82.885 205.745 83.055 205.935 ;
        RECT 84.725 205.765 84.895 205.955 ;
        RECT 88.405 205.745 88.575 205.935 ;
        RECT 89.380 205.795 89.500 205.905 ;
        RECT 90.245 205.765 90.415 205.955 ;
        RECT 92.085 205.745 92.255 205.935 ;
        RECT 95.765 205.765 95.935 205.955 ;
        RECT 97.605 205.745 97.775 205.935 ;
        RECT 101.285 205.765 101.455 205.955 ;
        RECT 102.260 205.795 102.380 205.905 ;
        RECT 103.125 205.745 103.295 205.935 ;
        RECT 104.045 205.765 104.215 205.955 ;
        RECT 108.645 205.745 108.815 205.935 ;
        RECT 109.565 205.765 109.735 205.955 ;
        RECT 114.165 205.745 114.335 205.935 ;
        RECT 115.085 205.905 115.255 205.955 ;
        RECT 115.085 205.795 115.260 205.905 ;
        RECT 115.085 205.765 115.255 205.795 ;
        RECT 120.605 205.745 120.775 205.955 ;
        RECT 126.125 205.745 126.295 205.955 ;
        RECT 127.505 205.745 127.675 205.955 ;
        RECT 14.665 204.935 16.035 205.745 ;
        RECT 16.965 204.935 20.635 205.745 ;
        RECT 20.645 204.935 26.155 205.745 ;
        RECT 26.165 204.935 31.675 205.745 ;
        RECT 31.685 204.935 37.195 205.745 ;
        RECT 37.215 204.875 37.645 205.660 ;
        RECT 37.665 204.935 39.495 205.745 ;
        RECT 39.505 204.935 45.015 205.745 ;
        RECT 45.025 204.935 50.535 205.745 ;
        RECT 50.545 204.935 56.055 205.745 ;
        RECT 56.065 204.935 61.575 205.745 ;
        RECT 61.595 204.835 62.945 205.745 ;
        RECT 62.975 204.875 63.405 205.660 ;
        RECT 64.355 204.835 65.705 205.745 ;
        RECT 65.725 205.065 74.915 205.745 ;
        RECT 65.725 204.835 66.645 205.065 ;
        RECT 69.475 204.845 70.405 205.065 ;
        RECT 74.925 204.935 77.675 205.745 ;
        RECT 77.685 204.935 83.195 205.745 ;
        RECT 83.205 204.935 88.715 205.745 ;
        RECT 88.735 204.875 89.165 205.660 ;
        RECT 89.645 204.935 92.395 205.745 ;
        RECT 92.405 204.935 97.915 205.745 ;
        RECT 97.925 204.935 103.435 205.745 ;
        RECT 103.445 204.935 108.955 205.745 ;
        RECT 108.965 204.935 114.475 205.745 ;
        RECT 114.495 204.875 114.925 205.660 ;
        RECT 115.405 204.935 120.915 205.745 ;
        RECT 120.925 204.935 126.435 205.745 ;
        RECT 126.445 204.935 127.815 205.745 ;
      LAYER nwell ;
        RECT 14.470 201.715 128.010 204.545 ;
      LAYER pwell ;
        RECT 14.665 200.515 16.035 201.325 ;
        RECT 16.045 200.515 18.795 201.325 ;
        RECT 18.805 200.515 24.315 201.325 ;
        RECT 24.335 200.600 24.765 201.385 ;
        RECT 25.245 200.515 27.995 201.325 ;
        RECT 28.005 200.515 33.515 201.325 ;
        RECT 33.525 200.515 39.035 201.325 ;
        RECT 39.045 200.515 44.555 201.325 ;
        RECT 44.565 200.515 50.075 201.325 ;
        RECT 50.095 200.600 50.525 201.385 ;
        RECT 51.005 200.515 52.835 201.325 ;
        RECT 52.845 200.515 58.355 201.325 ;
        RECT 58.565 201.195 60.775 201.425 ;
        RECT 63.495 201.195 64.425 201.415 ;
        RECT 58.565 200.515 68.935 201.195 ;
        RECT 69.405 200.515 72.155 201.325 ;
        RECT 72.165 200.515 73.535 201.295 ;
        RECT 74.475 200.515 75.825 201.425 ;
        RECT 75.855 200.600 76.285 201.385 ;
        RECT 76.305 200.515 78.135 201.325 ;
        RECT 78.145 200.515 83.655 201.325 ;
        RECT 83.665 200.515 89.175 201.325 ;
        RECT 89.185 200.515 94.695 201.325 ;
        RECT 94.705 200.515 100.215 201.325 ;
        RECT 100.235 200.515 101.585 201.425 ;
        RECT 101.615 200.600 102.045 201.385 ;
        RECT 102.065 200.515 103.895 201.325 ;
        RECT 103.905 201.195 104.825 201.425 ;
        RECT 107.655 201.195 108.585 201.415 ;
        RECT 103.905 200.515 113.095 201.195 ;
        RECT 113.565 200.515 115.395 201.325 ;
        RECT 115.405 200.515 120.915 201.325 ;
        RECT 120.925 200.515 126.435 201.325 ;
        RECT 126.445 200.515 127.815 201.325 ;
        RECT 14.805 200.305 14.975 200.515 ;
        RECT 16.645 200.350 16.805 200.460 ;
        RECT 18.485 200.325 18.655 200.515 ;
        RECT 20.325 200.305 20.495 200.495 ;
        RECT 24.005 200.325 24.175 200.515 ;
        RECT 24.980 200.355 25.100 200.465 ;
        RECT 25.845 200.305 26.015 200.495 ;
        RECT 27.685 200.325 27.855 200.515 ;
        RECT 31.365 200.305 31.535 200.495 ;
        RECT 33.205 200.325 33.375 200.515 ;
        RECT 36.885 200.305 37.055 200.495 ;
        RECT 37.860 200.355 37.980 200.465 ;
        RECT 38.725 200.325 38.895 200.515 ;
        RECT 40.565 200.305 40.735 200.495 ;
        RECT 44.245 200.325 44.415 200.515 ;
        RECT 46.085 200.305 46.255 200.495 ;
        RECT 49.765 200.325 49.935 200.515 ;
        RECT 50.740 200.355 50.860 200.465 ;
        RECT 51.605 200.305 51.775 200.495 ;
        RECT 52.525 200.325 52.695 200.515 ;
        RECT 57.125 200.305 57.295 200.495 ;
        RECT 58.045 200.325 58.215 200.515 ;
        RECT 62.645 200.305 62.815 200.495 ;
        RECT 63.620 200.355 63.740 200.465 ;
        RECT 66.325 200.305 66.495 200.495 ;
        RECT 66.785 200.305 66.955 200.495 ;
        RECT 68.625 200.325 68.795 200.515 ;
        RECT 69.140 200.355 69.260 200.465 ;
        RECT 69.545 200.305 69.715 200.495 ;
        RECT 71.845 200.305 72.015 200.515 ;
        RECT 72.305 200.325 72.475 200.515 ;
        RECT 74.145 200.360 74.305 200.470 ;
        RECT 74.605 200.325 74.775 200.515 ;
        RECT 77.825 200.325 77.995 200.515 ;
        RECT 81.045 200.305 81.215 200.495 ;
        RECT 81.560 200.355 81.680 200.465 ;
        RECT 83.345 200.325 83.515 200.515 ;
        RECT 87.025 200.305 87.195 200.495 ;
        RECT 87.485 200.305 87.655 200.495 ;
        RECT 88.865 200.325 89.035 200.515 ;
        RECT 94.385 200.325 94.555 200.515 ;
        RECT 98.065 200.305 98.235 200.495 ;
        RECT 99.905 200.325 100.075 200.515 ;
        RECT 100.365 200.325 100.535 200.515 ;
        RECT 103.585 200.325 103.755 200.515 ;
        RECT 107.265 200.305 107.435 200.495 ;
        RECT 108.645 200.305 108.815 200.495 ;
        RECT 109.105 200.305 109.275 200.495 ;
        RECT 110.540 200.355 110.660 200.465 ;
        RECT 112.785 200.325 112.955 200.515 ;
        RECT 113.300 200.355 113.420 200.465 ;
        RECT 114.165 200.305 114.335 200.495 ;
        RECT 115.085 200.465 115.255 200.515 ;
        RECT 115.085 200.355 115.260 200.465 ;
        RECT 115.085 200.325 115.255 200.355 ;
        RECT 120.605 200.305 120.775 200.515 ;
        RECT 126.125 200.305 126.295 200.515 ;
        RECT 127.505 200.305 127.675 200.515 ;
        RECT 14.665 199.495 16.035 200.305 ;
        RECT 16.965 199.495 20.635 200.305 ;
        RECT 20.645 199.495 26.155 200.305 ;
        RECT 26.165 199.495 31.675 200.305 ;
        RECT 31.685 199.495 37.195 200.305 ;
        RECT 37.215 199.435 37.645 200.220 ;
        RECT 38.125 199.495 40.875 200.305 ;
        RECT 40.885 199.495 46.395 200.305 ;
        RECT 46.405 199.495 51.915 200.305 ;
        RECT 51.925 199.495 57.435 200.305 ;
        RECT 57.445 199.495 62.955 200.305 ;
        RECT 62.975 199.435 63.405 200.220 ;
        RECT 63.885 199.495 66.635 200.305 ;
        RECT 66.645 199.525 68.015 200.305 ;
        RECT 68.025 199.495 69.855 200.305 ;
        RECT 69.865 199.625 72.155 200.305 ;
        RECT 72.165 199.625 81.355 200.305 ;
        RECT 69.865 199.395 70.785 199.625 ;
        RECT 72.165 199.395 73.085 199.625 ;
        RECT 75.915 199.405 76.845 199.625 ;
        RECT 81.825 199.495 87.335 200.305 ;
        RECT 87.355 199.395 88.705 200.305 ;
        RECT 88.735 199.435 89.165 200.220 ;
        RECT 89.185 199.625 98.375 200.305 ;
        RECT 98.385 199.625 107.575 200.305 ;
        RECT 89.185 199.395 90.105 199.625 ;
        RECT 92.935 199.405 93.865 199.625 ;
        RECT 98.385 199.395 99.305 199.625 ;
        RECT 102.135 199.405 103.065 199.625 ;
        RECT 107.585 199.525 108.955 200.305 ;
        RECT 108.975 199.395 110.325 200.305 ;
        RECT 110.805 199.495 114.475 200.305 ;
        RECT 114.495 199.435 114.925 200.220 ;
        RECT 115.405 199.495 120.915 200.305 ;
        RECT 120.925 199.495 126.435 200.305 ;
        RECT 126.445 199.495 127.815 200.305 ;
      LAYER nwell ;
        RECT 14.470 196.275 128.010 199.105 ;
      LAYER pwell ;
        RECT 14.665 195.075 16.035 195.885 ;
        RECT 16.045 195.075 18.795 195.885 ;
        RECT 18.805 195.075 24.315 195.885 ;
        RECT 24.335 195.160 24.765 195.945 ;
        RECT 25.245 195.075 27.995 195.885 ;
        RECT 28.005 195.075 33.515 195.885 ;
        RECT 33.525 195.075 39.035 195.885 ;
        RECT 39.045 195.075 44.555 195.885 ;
        RECT 44.565 195.075 50.075 195.885 ;
        RECT 50.095 195.160 50.525 195.945 ;
        RECT 50.545 195.075 56.055 195.885 ;
        RECT 56.065 195.075 61.575 195.885 ;
        RECT 61.595 195.075 62.945 195.985 ;
        RECT 62.965 195.075 64.795 195.885 ;
        RECT 66.175 195.755 67.095 195.985 ;
        RECT 64.805 195.075 67.095 195.755 ;
        RECT 67.105 195.075 70.025 195.985 ;
        RECT 70.325 195.785 71.270 195.985 ;
        RECT 72.605 195.785 73.535 195.985 ;
        RECT 70.325 195.305 73.535 195.785 ;
        RECT 73.855 195.755 74.785 195.985 ;
        RECT 70.325 195.105 73.395 195.305 ;
        RECT 70.325 195.075 71.270 195.105 ;
        RECT 14.805 194.865 14.975 195.075 ;
        RECT 16.645 194.910 16.805 195.020 ;
        RECT 18.485 194.885 18.655 195.075 ;
        RECT 20.325 194.865 20.495 195.055 ;
        RECT 24.005 194.885 24.175 195.075 ;
        RECT 24.980 194.915 25.100 195.025 ;
        RECT 25.845 194.865 26.015 195.055 ;
        RECT 27.685 194.885 27.855 195.075 ;
        RECT 31.365 194.865 31.535 195.055 ;
        RECT 33.205 194.885 33.375 195.075 ;
        RECT 36.885 194.865 37.055 195.055 ;
        RECT 38.725 194.885 38.895 195.075 ;
        RECT 42.865 194.865 43.035 195.055 ;
        RECT 44.245 194.885 44.415 195.075 ;
        RECT 48.385 194.865 48.555 195.055 ;
        RECT 49.765 194.865 49.935 195.075 ;
        RECT 51.605 194.865 51.775 195.055 ;
        RECT 52.065 194.865 52.235 195.055 ;
        RECT 53.445 194.865 53.615 195.055 ;
        RECT 55.745 194.885 55.915 195.075 ;
        RECT 61.265 194.885 61.435 195.075 ;
        RECT 62.645 194.885 62.815 195.075 ;
        RECT 63.620 194.915 63.740 195.025 ;
        RECT 64.485 194.885 64.655 195.075 ;
        RECT 64.945 194.885 65.115 195.075 ;
        RECT 65.405 194.865 65.575 195.055 ;
        RECT 67.250 194.885 67.420 195.075 ;
        RECT 68.625 194.865 68.795 195.055 ;
        RECT 14.665 194.055 16.035 194.865 ;
        RECT 16.965 194.055 20.635 194.865 ;
        RECT 20.645 194.055 26.155 194.865 ;
        RECT 26.165 194.055 31.675 194.865 ;
        RECT 31.685 194.055 37.195 194.865 ;
        RECT 37.215 193.995 37.645 194.780 ;
        RECT 37.665 194.055 43.175 194.865 ;
        RECT 43.185 194.055 48.695 194.865 ;
        RECT 48.715 193.955 50.065 194.865 ;
        RECT 50.085 194.055 51.915 194.865 ;
        RECT 51.935 193.955 53.285 194.865 ;
        RECT 53.305 194.185 62.915 194.865 ;
        RECT 57.815 193.965 58.745 194.185 ;
        RECT 61.575 193.955 62.915 194.185 ;
        RECT 62.975 193.995 63.405 194.780 ;
        RECT 63.885 194.055 65.715 194.865 ;
        RECT 65.725 193.955 68.835 194.865 ;
        RECT 69.085 194.835 69.255 195.055 ;
        RECT 72.360 194.915 72.480 195.025 ;
        RECT 73.225 194.885 73.395 195.105 ;
        RECT 73.855 195.075 75.690 195.755 ;
        RECT 75.855 195.160 76.285 195.945 ;
        RECT 76.865 195.075 79.975 195.985 ;
        RECT 80.905 195.075 84.575 195.885 ;
        RECT 84.585 195.075 90.095 195.885 ;
        RECT 93.305 195.755 94.235 195.985 ;
        RECT 90.335 195.075 94.235 195.755 ;
        RECT 94.245 195.075 95.615 195.855 ;
        RECT 95.625 195.075 97.455 195.885 ;
        RECT 100.665 195.755 101.595 195.985 ;
        RECT 97.695 195.075 101.595 195.755 ;
        RECT 101.615 195.160 102.045 195.945 ;
        RECT 102.525 195.075 104.355 195.885 ;
        RECT 107.565 195.755 108.495 195.985 ;
        RECT 104.595 195.075 108.495 195.755 ;
        RECT 109.425 195.075 110.795 195.855 ;
        RECT 111.725 195.075 115.395 195.885 ;
        RECT 115.405 195.075 120.915 195.885 ;
        RECT 120.925 195.075 126.435 195.885 ;
        RECT 126.445 195.075 127.815 195.885 ;
        RECT 75.525 195.055 75.690 195.075 ;
        RECT 74.145 194.865 74.315 195.055 ;
        RECT 74.600 194.865 74.770 195.055 ;
        RECT 75.525 194.885 75.695 195.055 ;
        RECT 76.040 194.915 76.160 195.025 ;
        RECT 76.500 194.915 76.620 195.025 ;
        RECT 76.905 194.885 77.075 195.075 ;
        RECT 78.745 194.865 78.915 195.055 ;
        RECT 80.585 194.920 80.745 195.030 ;
        RECT 84.265 194.865 84.435 195.075 ;
        RECT 88.130 194.865 88.300 195.055 ;
        RECT 89.380 194.915 89.500 195.025 ;
        RECT 89.785 194.865 89.955 195.075 ;
        RECT 92.085 194.865 92.255 195.055 ;
        RECT 93.650 194.885 93.820 195.075 ;
        RECT 94.385 194.885 94.555 195.075 ;
        RECT 97.145 194.885 97.315 195.075 ;
        RECT 97.605 194.865 97.775 195.055 ;
        RECT 101.010 194.885 101.180 195.075 ;
        RECT 102.260 194.915 102.380 195.025 ;
        RECT 103.125 194.865 103.295 195.055 ;
        RECT 103.585 194.865 103.755 195.055 ;
        RECT 104.045 194.885 104.215 195.075 ;
        RECT 107.910 194.885 108.080 195.075 ;
        RECT 108.370 194.865 108.540 195.055 ;
        RECT 109.105 194.865 109.275 195.055 ;
        RECT 109.565 194.885 109.735 195.075 ;
        RECT 110.540 194.915 110.660 195.025 ;
        RECT 111.405 194.920 111.565 195.030 ;
        RECT 114.165 194.865 114.335 195.055 ;
        RECT 115.085 195.025 115.255 195.075 ;
        RECT 115.085 194.915 115.260 195.025 ;
        RECT 115.085 194.885 115.255 194.915 ;
        RECT 120.605 194.865 120.775 195.075 ;
        RECT 126.125 194.865 126.295 195.075 ;
        RECT 127.505 194.865 127.675 195.075 ;
        RECT 71.210 194.835 72.155 194.865 ;
        RECT 69.085 194.635 72.155 194.835 ;
        RECT 68.945 194.155 72.155 194.635 ;
        RECT 68.945 193.955 69.875 194.155 ;
        RECT 71.210 193.955 72.155 194.155 ;
        RECT 72.625 194.055 74.455 194.865 ;
        RECT 74.485 193.955 75.835 194.865 ;
        RECT 76.305 194.055 79.055 194.865 ;
        RECT 79.065 194.055 84.575 194.865 ;
        RECT 84.815 194.185 88.715 194.865 ;
        RECT 87.785 193.955 88.715 194.185 ;
        RECT 88.735 193.995 89.165 194.780 ;
        RECT 89.645 194.085 91.015 194.865 ;
        RECT 91.025 194.055 92.395 194.865 ;
        RECT 92.405 194.055 97.915 194.865 ;
        RECT 97.925 194.055 103.435 194.865 ;
        RECT 103.455 193.955 104.805 194.865 ;
        RECT 105.055 194.185 108.955 194.865 ;
        RECT 108.025 193.955 108.955 194.185 ;
        RECT 108.965 194.085 110.335 194.865 ;
        RECT 110.805 194.055 114.475 194.865 ;
        RECT 114.495 193.995 114.925 194.780 ;
        RECT 115.405 194.055 120.915 194.865 ;
        RECT 120.925 194.055 126.435 194.865 ;
        RECT 126.445 194.055 127.815 194.865 ;
      LAYER nwell ;
        RECT 14.470 190.835 128.010 193.665 ;
      LAYER pwell ;
        RECT 14.665 189.635 16.035 190.445 ;
        RECT 16.045 189.635 18.795 190.445 ;
        RECT 18.805 189.635 24.315 190.445 ;
        RECT 24.335 189.720 24.765 190.505 ;
        RECT 25.705 189.635 29.375 190.445 ;
        RECT 29.385 189.635 34.895 190.445 ;
        RECT 34.905 189.635 40.415 190.445 ;
        RECT 40.795 190.435 41.715 190.545 ;
        RECT 40.795 190.315 43.130 190.435 ;
        RECT 47.795 190.315 48.715 190.535 ;
        RECT 40.795 189.635 50.075 190.315 ;
        RECT 50.095 189.720 50.525 190.505 ;
        RECT 50.915 190.435 51.835 190.545 ;
        RECT 50.915 190.315 53.250 190.435 ;
        RECT 57.915 190.315 58.835 190.535 ;
        RECT 50.915 189.635 60.195 190.315 ;
        RECT 60.665 189.635 63.415 190.445 ;
        RECT 63.425 189.635 68.935 190.445 ;
        RECT 68.945 189.635 71.235 190.545 ;
        RECT 72.165 189.635 75.835 190.445 ;
        RECT 75.855 189.720 76.285 190.505 ;
        RECT 76.305 189.635 77.675 190.445 ;
        RECT 77.685 189.635 81.355 190.445 ;
        RECT 81.375 189.635 82.725 190.545 ;
        RECT 82.755 189.635 84.105 190.545 ;
        RECT 84.495 190.435 85.415 190.545 ;
        RECT 84.495 190.315 86.830 190.435 ;
        RECT 91.495 190.315 92.415 190.535 ;
        RECT 84.495 189.635 93.775 190.315 ;
        RECT 94.245 189.635 96.075 190.445 ;
        RECT 96.085 189.635 101.595 190.445 ;
        RECT 101.615 189.720 102.045 190.505 ;
        RECT 102.065 189.635 103.435 190.445 ;
        RECT 103.445 190.315 104.365 190.545 ;
        RECT 107.195 190.315 108.125 190.535 ;
        RECT 103.445 189.635 112.635 190.315 ;
        RECT 112.645 189.635 114.015 190.445 ;
        RECT 114.025 189.635 117.695 190.445 ;
        RECT 117.715 189.635 119.065 190.545 ;
        RECT 119.085 189.635 120.915 190.445 ;
        RECT 120.925 189.635 126.435 190.445 ;
        RECT 126.445 189.635 127.815 190.445 ;
        RECT 14.805 189.425 14.975 189.635 ;
        RECT 16.645 189.470 16.805 189.580 ;
        RECT 18.485 189.445 18.655 189.635 ;
        RECT 20.325 189.425 20.495 189.615 ;
        RECT 24.005 189.445 24.175 189.635 ;
        RECT 25.385 189.480 25.545 189.590 ;
        RECT 25.845 189.425 26.015 189.615 ;
        RECT 29.065 189.445 29.235 189.635 ;
        RECT 31.365 189.425 31.535 189.615 ;
        RECT 34.585 189.445 34.755 189.635 ;
        RECT 36.885 189.425 37.055 189.615 ;
        RECT 40.105 189.445 40.275 189.635 ;
        RECT 41.025 189.425 41.195 189.615 ;
        RECT 46.545 189.425 46.715 189.615 ;
        RECT 49.765 189.445 49.935 189.635 ;
        RECT 50.410 189.425 50.580 189.615 ;
        RECT 54.550 189.425 54.720 189.615 ;
        RECT 55.340 189.475 55.460 189.585 ;
        RECT 55.745 189.425 55.915 189.615 ;
        RECT 57.125 189.425 57.295 189.615 ;
        RECT 58.965 189.470 59.125 189.580 ;
        RECT 59.885 189.445 60.055 189.635 ;
        RECT 60.400 189.475 60.520 189.585 ;
        RECT 62.645 189.425 62.815 189.615 ;
        RECT 63.105 189.445 63.275 189.635 ;
        RECT 64.945 189.425 65.115 189.615 ;
        RECT 65.405 189.425 65.575 189.615 ;
        RECT 66.785 189.425 66.955 189.615 ;
        RECT 68.625 189.445 68.795 189.635 ;
        RECT 70.920 189.615 71.090 189.635 ;
        RECT 69.085 189.470 69.245 189.580 ;
        RECT 70.920 189.445 71.095 189.615 ;
        RECT 71.845 189.480 72.005 189.590 ;
        RECT 70.925 189.425 71.095 189.445 ;
        RECT 72.765 189.425 72.935 189.615 ;
        RECT 73.225 189.425 73.395 189.615 ;
        RECT 75.065 189.470 75.225 189.580 ;
        RECT 75.525 189.445 75.695 189.635 ;
        RECT 77.365 189.445 77.535 189.635 ;
        RECT 78.745 189.425 78.915 189.615 ;
        RECT 81.045 189.445 81.215 189.635 ;
        RECT 81.505 189.445 81.675 189.635 ;
        RECT 83.805 189.445 83.975 189.635 ;
        RECT 88.405 189.425 88.575 189.615 ;
        RECT 90.245 189.425 90.415 189.615 ;
        RECT 90.760 189.475 90.880 189.585 ;
        RECT 93.465 189.425 93.635 189.635 ;
        RECT 93.980 189.475 94.100 189.585 ;
        RECT 95.765 189.445 95.935 189.635 ;
        RECT 98.985 189.425 99.155 189.615 ;
        RECT 101.285 189.445 101.455 189.635 ;
        RECT 103.125 189.445 103.295 189.635 ;
        RECT 108.185 189.425 108.355 189.615 ;
        RECT 108.700 189.475 108.820 189.585 ;
        RECT 112.325 189.445 112.495 189.635 ;
        RECT 113.705 189.445 113.875 189.635 ;
        RECT 114.165 189.425 114.335 189.615 ;
        RECT 117.385 189.445 117.555 189.635 ;
        RECT 118.765 189.445 118.935 189.635 ;
        RECT 120.605 189.445 120.775 189.635 ;
        RECT 123.825 189.425 123.995 189.615 ;
        RECT 124.340 189.475 124.460 189.585 ;
        RECT 126.125 189.425 126.295 189.635 ;
        RECT 127.505 189.425 127.675 189.635 ;
        RECT 14.665 188.615 16.035 189.425 ;
        RECT 16.965 188.615 20.635 189.425 ;
        RECT 20.645 188.615 26.155 189.425 ;
        RECT 26.165 188.615 31.675 189.425 ;
        RECT 31.685 188.615 37.195 189.425 ;
        RECT 37.215 188.555 37.645 189.340 ;
        RECT 37.665 188.615 41.335 189.425 ;
        RECT 41.345 188.615 46.855 189.425 ;
        RECT 47.095 188.745 50.995 189.425 ;
        RECT 51.235 188.745 55.135 189.425 ;
        RECT 50.065 188.515 50.995 188.745 ;
        RECT 54.205 188.515 55.135 188.745 ;
        RECT 55.615 188.515 56.965 189.425 ;
        RECT 56.985 188.645 58.355 189.425 ;
        RECT 59.285 188.615 62.955 189.425 ;
        RECT 62.975 188.555 63.405 189.340 ;
        RECT 63.425 188.615 65.255 189.425 ;
        RECT 65.275 188.515 66.625 189.425 ;
        RECT 66.645 188.745 68.475 189.425 ;
        RECT 69.405 188.745 71.235 189.425 ;
        RECT 69.405 188.515 70.750 188.745 ;
        RECT 71.245 188.615 73.075 189.425 ;
        RECT 73.095 188.515 74.445 189.425 ;
        RECT 75.385 188.615 79.055 189.425 ;
        RECT 79.435 188.745 88.715 189.425 ;
        RECT 79.435 188.625 81.770 188.745 ;
        RECT 79.435 188.515 80.355 188.625 ;
        RECT 86.435 188.525 87.355 188.745 ;
        RECT 88.735 188.555 89.165 189.340 ;
        RECT 89.185 188.645 90.555 189.425 ;
        RECT 91.025 188.615 93.775 189.425 ;
        RECT 93.785 188.615 99.295 189.425 ;
        RECT 99.305 188.745 108.495 189.425 ;
        RECT 99.305 188.515 100.225 188.745 ;
        RECT 103.055 188.525 103.985 188.745 ;
        RECT 108.965 188.615 114.475 189.425 ;
        RECT 114.495 188.555 114.925 189.340 ;
        RECT 114.945 188.745 124.135 189.425 ;
        RECT 114.945 188.515 115.865 188.745 ;
        RECT 118.695 188.525 119.625 188.745 ;
        RECT 124.605 188.615 126.435 189.425 ;
        RECT 126.445 188.615 127.815 189.425 ;
      LAYER nwell ;
        RECT 14.470 185.395 128.010 188.225 ;
      LAYER pwell ;
        RECT 14.665 184.195 16.035 185.005 ;
        RECT 16.045 184.195 18.795 185.005 ;
        RECT 18.805 184.195 24.315 185.005 ;
        RECT 24.335 184.280 24.765 185.065 ;
        RECT 24.785 184.195 26.615 185.005 ;
        RECT 26.625 184.195 32.135 185.005 ;
        RECT 32.155 184.195 33.505 185.105 ;
        RECT 33.525 184.195 35.355 185.005 ;
        RECT 35.365 184.875 36.295 185.105 ;
        RECT 35.365 184.195 39.265 184.875 ;
        RECT 39.505 184.195 41.335 185.005 ;
        RECT 44.545 184.875 45.475 185.105 ;
        RECT 41.575 184.195 45.475 184.875 ;
        RECT 46.405 184.195 50.075 185.005 ;
        RECT 50.095 184.280 50.525 185.065 ;
        RECT 52.755 184.995 53.675 185.105 ;
        RECT 50.545 184.195 51.915 184.975 ;
        RECT 52.755 184.875 55.090 184.995 ;
        RECT 59.755 184.875 60.675 185.095 ;
        RECT 65.705 184.875 66.635 185.105 ;
        RECT 52.755 184.195 62.035 184.875 ;
        RECT 62.965 184.195 66.635 184.875 ;
        RECT 66.645 184.875 67.565 185.105 ;
        RECT 70.395 184.875 71.325 185.095 ;
        RECT 66.645 184.195 75.835 184.875 ;
        RECT 75.855 184.280 76.285 185.065 ;
        RECT 76.305 184.195 77.675 185.005 ;
        RECT 77.685 184.195 81.355 185.005 ;
        RECT 81.375 184.195 82.725 185.105 ;
        RECT 85.945 184.875 86.875 185.105 ;
        RECT 82.975 184.195 86.875 184.875 ;
        RECT 86.885 184.195 88.255 185.005 ;
        RECT 88.265 184.195 91.935 185.005 ;
        RECT 91.945 184.195 97.455 185.005 ;
        RECT 100.665 184.875 101.595 185.105 ;
        RECT 97.695 184.195 101.595 184.875 ;
        RECT 101.615 184.280 102.045 185.065 ;
        RECT 105.725 184.875 106.655 185.105 ;
        RECT 102.755 184.195 106.655 184.875 ;
        RECT 106.675 184.195 108.025 185.105 ;
        RECT 108.045 184.195 109.415 184.975 ;
        RECT 109.885 184.195 113.555 185.005 ;
        RECT 113.575 184.195 114.925 185.105 ;
        RECT 114.945 184.875 115.865 185.105 ;
        RECT 118.695 184.875 119.625 185.095 ;
        RECT 114.945 184.195 124.135 184.875 ;
        RECT 124.145 184.195 125.515 184.975 ;
        RECT 126.445 184.195 127.815 185.005 ;
        RECT 14.805 183.985 14.975 184.195 ;
        RECT 16.645 184.030 16.805 184.140 ;
        RECT 18.485 184.005 18.655 184.195 ;
        RECT 22.165 183.985 22.335 184.175 ;
        RECT 24.005 184.005 24.175 184.195 ;
        RECT 26.305 184.005 26.475 184.195 ;
        RECT 27.685 183.985 27.855 184.175 ;
        RECT 31.825 184.005 31.995 184.195 ;
        RECT 33.205 184.005 33.375 184.195 ;
        RECT 35.045 184.005 35.215 184.195 ;
        RECT 35.780 184.005 35.950 184.195 ;
        RECT 36.885 183.985 37.055 184.175 ;
        RECT 41.025 184.005 41.195 184.195 ;
        RECT 44.890 184.005 45.060 184.195 ;
        RECT 46.085 184.040 46.245 184.150 ;
        RECT 46.545 183.985 46.715 184.175 ;
        RECT 49.765 184.005 49.935 184.195 ;
        RECT 51.605 184.005 51.775 184.195 ;
        RECT 52.065 184.145 52.235 184.175 ;
        RECT 52.065 184.035 52.240 184.145 ;
        RECT 52.065 183.985 52.235 184.035 ;
        RECT 57.585 183.985 57.755 184.175 ;
        RECT 58.045 183.985 58.215 184.175 ;
        RECT 61.725 184.005 61.895 184.195 ;
        RECT 62.645 183.985 62.815 184.175 ;
        RECT 63.105 184.005 63.275 184.195 ;
        RECT 64.945 183.985 65.115 184.175 ;
        RECT 65.405 183.985 65.575 184.175 ;
        RECT 71.385 183.985 71.555 184.175 ;
        RECT 71.900 184.035 72.020 184.145 ;
        RECT 74.605 183.985 74.775 184.175 ;
        RECT 75.070 183.985 75.240 184.175 ;
        RECT 75.525 184.005 75.695 184.195 ;
        RECT 77.365 184.005 77.535 184.195 ;
        RECT 78.285 184.030 78.445 184.140 ;
        RECT 81.045 184.005 81.215 184.195 ;
        RECT 82.425 184.005 82.595 184.195 ;
        RECT 86.290 184.005 86.460 184.195 ;
        RECT 87.485 183.985 87.655 184.175 ;
        RECT 87.945 184.005 88.115 184.195 ;
        RECT 88.405 184.030 88.565 184.140 ;
        RECT 90.245 183.985 90.415 184.175 ;
        RECT 90.705 183.985 90.875 184.175 ;
        RECT 91.625 184.005 91.795 184.195 ;
        RECT 92.085 183.985 92.255 184.175 ;
        RECT 97.145 184.005 97.315 184.195 ;
        RECT 101.010 184.005 101.180 184.195 ;
        RECT 102.205 184.145 102.375 184.175 ;
        RECT 102.205 184.035 102.380 184.145 ;
        RECT 102.205 183.985 102.375 184.035 ;
        RECT 103.585 183.985 103.755 184.175 ;
        RECT 106.070 184.005 106.240 184.195 ;
        RECT 107.265 183.985 107.435 184.175 ;
        RECT 107.725 183.985 107.895 184.195 ;
        RECT 109.105 184.005 109.275 184.195 ;
        RECT 109.620 184.035 109.740 184.145 ;
        RECT 112.510 183.985 112.680 184.175 ;
        RECT 113.245 184.005 113.415 184.195 ;
        RECT 113.705 184.005 113.875 184.195 ;
        RECT 114.165 183.985 114.335 184.175 ;
        RECT 118.490 183.985 118.660 184.175 ;
        RECT 119.280 184.035 119.400 184.145 ;
        RECT 119.685 183.985 119.855 184.175 ;
        RECT 123.825 184.005 123.995 184.195 ;
        RECT 125.205 184.005 125.375 184.195 ;
        RECT 126.125 183.985 126.295 184.175 ;
        RECT 127.505 183.985 127.675 184.195 ;
        RECT 14.665 183.175 16.035 183.985 ;
        RECT 16.965 183.175 22.475 183.985 ;
        RECT 22.485 183.175 27.995 183.985 ;
        RECT 28.005 183.305 37.195 183.985 ;
        RECT 28.005 183.075 28.925 183.305 ;
        RECT 31.755 183.085 32.685 183.305 ;
        RECT 37.215 183.115 37.645 183.900 ;
        RECT 37.665 183.305 46.855 183.985 ;
        RECT 37.665 183.075 38.585 183.305 ;
        RECT 41.415 183.085 42.345 183.305 ;
        RECT 46.865 183.175 52.375 183.985 ;
        RECT 52.385 183.175 57.895 183.985 ;
        RECT 57.905 183.205 59.275 183.985 ;
        RECT 59.285 183.175 62.955 183.985 ;
        RECT 62.975 183.115 63.405 183.900 ;
        RECT 63.425 183.175 65.255 183.985 ;
        RECT 65.265 183.305 67.095 183.985 ;
        RECT 67.115 183.945 68.035 183.985 ;
        RECT 67.105 183.755 68.035 183.945 ;
        RECT 70.125 183.755 71.695 183.985 ;
        RECT 67.105 183.395 71.695 183.755 ;
        RECT 65.750 183.075 67.095 183.305 ;
        RECT 67.115 183.305 71.695 183.395 ;
        RECT 67.115 183.075 70.115 183.305 ;
        RECT 72.165 183.175 74.915 183.985 ;
        RECT 74.925 183.075 77.535 183.985 ;
        RECT 78.605 183.305 87.795 183.985 ;
        RECT 78.605 183.075 79.525 183.305 ;
        RECT 82.355 183.085 83.285 183.305 ;
        RECT 88.735 183.115 89.165 183.900 ;
        RECT 89.185 183.175 90.555 183.985 ;
        RECT 90.565 183.205 91.935 183.985 ;
        RECT 91.955 183.075 93.305 183.985 ;
        RECT 93.325 183.305 102.515 183.985 ;
        RECT 93.325 183.075 94.245 183.305 ;
        RECT 97.075 183.085 98.005 183.305 ;
        RECT 102.525 183.205 103.895 183.985 ;
        RECT 103.905 183.175 107.575 183.985 ;
        RECT 107.595 183.075 108.945 183.985 ;
        RECT 109.195 183.305 113.095 183.985 ;
        RECT 112.165 183.075 113.095 183.305 ;
        RECT 113.105 183.175 114.475 183.985 ;
        RECT 114.495 183.115 114.925 183.900 ;
        RECT 115.175 183.305 119.075 183.985 ;
        RECT 118.145 183.075 119.075 183.305 ;
        RECT 119.545 183.205 120.915 183.985 ;
        RECT 120.925 183.175 126.435 183.985 ;
        RECT 126.445 183.175 127.815 183.985 ;
      LAYER nwell ;
        RECT 14.470 179.955 128.010 182.785 ;
      LAYER pwell ;
        RECT 14.665 178.755 16.035 179.565 ;
        RECT 16.045 178.755 17.415 179.565 ;
        RECT 17.425 178.755 22.935 179.565 ;
        RECT 22.955 178.755 24.305 179.665 ;
        RECT 24.335 178.840 24.765 179.625 ;
        RECT 29.295 179.435 30.225 179.655 ;
        RECT 33.055 179.435 33.975 179.665 ;
        RECT 24.785 178.755 33.975 179.435 ;
        RECT 33.985 178.755 35.815 179.565 ;
        RECT 35.835 178.755 37.185 179.665 ;
        RECT 37.205 178.755 38.575 179.535 ;
        RECT 39.505 178.755 43.175 179.565 ;
        RECT 43.185 178.755 44.555 179.535 ;
        RECT 45.025 178.755 48.695 179.565 ;
        RECT 48.715 178.755 50.065 179.665 ;
        RECT 50.095 178.840 50.525 179.625 ;
        RECT 50.545 178.755 52.375 179.565 ;
        RECT 52.395 178.755 53.745 179.665 ;
        RECT 56.965 179.435 57.895 179.665 ;
        RECT 53.995 178.755 57.895 179.435 ;
        RECT 57.905 178.755 59.275 179.535 ;
        RECT 59.285 178.755 64.795 179.565 ;
        RECT 64.805 178.755 70.315 179.565 ;
        RECT 70.325 178.755 75.835 179.565 ;
        RECT 75.855 178.840 76.285 179.625 ;
        RECT 77.225 178.755 79.835 179.665 ;
        RECT 83.185 179.435 84.115 179.665 ;
        RECT 80.215 178.755 84.115 179.435 ;
        RECT 84.125 179.435 85.045 179.665 ;
        RECT 87.875 179.435 88.805 179.655 ;
        RECT 84.125 178.755 93.315 179.435 ;
        RECT 93.325 178.755 96.075 179.565 ;
        RECT 96.085 178.755 101.595 179.565 ;
        RECT 101.615 178.840 102.045 179.625 ;
        RECT 102.985 178.755 108.495 179.565 ;
        RECT 108.505 179.435 109.425 179.665 ;
        RECT 112.255 179.435 113.185 179.655 ;
        RECT 120.905 179.435 121.835 179.665 ;
        RECT 108.505 178.755 117.695 179.435 ;
        RECT 117.935 178.755 121.835 179.435 ;
        RECT 122.765 178.755 126.435 179.565 ;
        RECT 126.445 178.755 127.815 179.565 ;
        RECT 14.805 178.545 14.975 178.755 ;
        RECT 16.645 178.590 16.805 178.700 ;
        RECT 17.105 178.565 17.275 178.755 ;
        RECT 22.165 178.545 22.335 178.735 ;
        RECT 22.625 178.565 22.795 178.755 ;
        RECT 23.085 178.565 23.255 178.755 ;
        RECT 24.925 178.565 25.095 178.755 ;
        RECT 27.685 178.545 27.855 178.735 ;
        RECT 29.065 178.545 29.235 178.735 ;
        RECT 29.800 178.545 29.970 178.735 ;
        RECT 35.505 178.565 35.675 178.755 ;
        RECT 35.965 178.565 36.135 178.755 ;
        RECT 36.885 178.545 37.055 178.735 ;
        RECT 38.265 178.565 38.435 178.755 ;
        RECT 39.185 178.600 39.345 178.710 ;
        RECT 42.865 178.545 43.035 178.755 ;
        RECT 43.325 178.565 43.495 178.755 ;
        RECT 44.760 178.595 44.880 178.705 ;
        RECT 48.385 178.565 48.555 178.755 ;
        RECT 49.765 178.565 49.935 178.755 ;
        RECT 52.065 178.565 52.235 178.755 ;
        RECT 52.525 178.545 52.695 178.755 ;
        RECT 57.310 178.565 57.480 178.755 ;
        RECT 58.045 178.565 58.215 178.755 ;
        RECT 62.185 178.545 62.355 178.735 ;
        RECT 62.700 178.595 62.820 178.705 ;
        RECT 64.485 178.565 64.655 178.755 ;
        RECT 64.945 178.545 65.115 178.735 ;
        RECT 70.005 178.565 70.175 178.755 ;
        RECT 70.465 178.545 70.635 178.735 ;
        RECT 70.925 178.565 71.095 178.735 ;
        RECT 75.525 178.565 75.695 178.755 ;
        RECT 76.905 178.600 77.065 178.710 ;
        RECT 77.370 178.565 77.540 178.755 ;
        RECT 71.025 178.545 71.095 178.565 ;
        RECT 79.205 178.545 79.375 178.735 ;
        RECT 79.665 178.545 79.835 178.735 ;
        RECT 83.530 178.565 83.700 178.755 ;
        RECT 89.600 178.545 89.770 178.735 ;
        RECT 93.005 178.565 93.175 178.755 ;
        RECT 93.520 178.595 93.640 178.705 ;
        RECT 95.765 178.565 95.935 178.755 ;
        RECT 98.985 178.545 99.155 178.735 ;
        RECT 100.365 178.545 100.535 178.735 ;
        RECT 101.285 178.565 101.455 178.755 ;
        RECT 101.745 178.545 101.915 178.735 ;
        RECT 102.665 178.600 102.825 178.710 ;
        RECT 108.185 178.565 108.355 178.755 ;
        RECT 111.000 178.595 111.120 178.705 ;
        RECT 112.785 178.545 112.955 178.735 ;
        RECT 113.245 178.545 113.415 178.735 ;
        RECT 115.140 178.595 115.260 178.705 ;
        RECT 117.385 178.565 117.555 178.755 ;
        RECT 120.605 178.545 120.775 178.735 ;
        RECT 121.250 178.565 121.420 178.755 ;
        RECT 122.445 178.600 122.605 178.710 ;
        RECT 126.125 178.545 126.295 178.755 ;
        RECT 127.505 178.545 127.675 178.755 ;
        RECT 14.665 177.735 16.035 178.545 ;
        RECT 16.965 177.735 22.475 178.545 ;
        RECT 22.485 177.735 27.995 178.545 ;
        RECT 28.005 177.765 29.375 178.545 ;
        RECT 29.385 177.865 33.285 178.545 ;
        RECT 29.385 177.635 30.315 177.865 ;
        RECT 33.525 177.735 37.195 178.545 ;
        RECT 37.215 177.675 37.645 178.460 ;
        RECT 37.665 177.735 43.175 178.545 ;
        RECT 43.555 177.865 52.835 178.545 ;
        RECT 53.215 177.865 62.495 178.545 ;
        RECT 43.555 177.745 45.890 177.865 ;
        RECT 43.555 177.635 44.475 177.745 ;
        RECT 50.555 177.645 51.475 177.865 ;
        RECT 53.215 177.745 55.550 177.865 ;
        RECT 53.215 177.635 54.135 177.745 ;
        RECT 60.215 177.645 61.135 177.865 ;
        RECT 62.975 177.675 63.405 178.460 ;
        RECT 63.425 177.735 65.255 178.545 ;
        RECT 65.265 177.735 70.775 178.545 ;
        RECT 71.025 178.315 73.295 178.545 ;
        RECT 71.025 177.635 73.780 178.315 ;
        RECT 74.005 177.735 79.515 178.545 ;
        RECT 79.525 177.865 88.630 178.545 ;
        RECT 88.735 177.675 89.165 178.460 ;
        RECT 89.185 177.865 93.085 178.545 ;
        RECT 89.185 177.635 90.115 177.865 ;
        RECT 93.785 177.735 99.295 178.545 ;
        RECT 99.315 177.635 100.665 178.545 ;
        RECT 101.605 177.865 110.710 178.545 ;
        RECT 111.265 177.735 113.095 178.545 ;
        RECT 113.105 177.765 114.475 178.545 ;
        RECT 114.495 177.675 114.925 178.460 ;
        RECT 115.405 177.735 120.915 178.545 ;
        RECT 120.925 177.735 126.435 178.545 ;
        RECT 126.445 177.735 127.815 178.545 ;
      LAYER nwell ;
        RECT 14.470 174.515 128.010 177.345 ;
      LAYER pwell ;
        RECT 14.665 173.315 16.035 174.125 ;
        RECT 16.045 173.315 18.795 174.125 ;
        RECT 18.805 173.315 24.315 174.125 ;
        RECT 24.335 173.400 24.765 174.185 ;
        RECT 24.785 173.315 28.455 174.125 ;
        RECT 31.665 173.995 32.595 174.225 ;
        RECT 28.695 173.315 32.595 173.995 ;
        RECT 32.605 173.315 33.975 174.125 ;
        RECT 33.995 173.315 35.345 174.225 ;
        RECT 35.365 173.995 36.285 174.225 ;
        RECT 39.115 173.995 40.045 174.215 ;
        RECT 48.685 173.995 49.615 174.225 ;
        RECT 35.365 173.315 44.555 173.995 ;
        RECT 45.715 173.315 49.615 173.995 ;
        RECT 50.095 173.400 50.525 174.185 ;
        RECT 50.545 173.315 51.915 174.095 ;
        RECT 51.925 173.315 53.295 174.125 ;
        RECT 56.505 173.995 57.435 174.225 ;
        RECT 53.535 173.315 57.435 173.995 ;
        RECT 57.905 173.315 61.575 174.125 ;
        RECT 61.585 173.315 67.095 174.125 ;
        RECT 67.345 173.545 70.100 174.225 ;
        RECT 71.905 173.995 74.905 174.225 ;
        RECT 70.325 173.905 74.905 173.995 ;
        RECT 70.325 173.545 74.915 173.905 ;
        RECT 67.345 173.315 69.615 173.545 ;
        RECT 70.325 173.315 71.895 173.545 ;
        RECT 73.985 173.355 74.915 173.545 ;
        RECT 75.855 173.400 76.285 174.185 ;
        RECT 76.520 173.545 79.275 174.225 ;
        RECT 73.985 173.315 74.905 173.355 ;
        RECT 77.005 173.315 79.275 173.545 ;
        RECT 79.525 173.315 82.265 173.995 ;
        RECT 82.745 173.315 85.495 174.125 ;
        RECT 85.505 173.315 86.875 174.095 ;
        RECT 86.895 173.315 88.245 174.225 ;
        RECT 96.915 173.995 97.845 174.215 ;
        RECT 100.675 173.995 101.595 174.225 ;
        RECT 89.195 173.315 91.935 173.995 ;
        RECT 92.405 173.315 101.595 173.995 ;
        RECT 101.615 173.400 102.045 174.185 ;
        RECT 102.085 173.315 113.095 174.225 ;
        RECT 113.565 173.315 115.395 174.125 ;
        RECT 118.605 173.995 119.535 174.225 ;
        RECT 115.635 173.315 119.535 173.995 ;
        RECT 119.555 173.315 120.905 174.225 ;
        RECT 121.845 173.315 123.215 174.095 ;
        RECT 123.685 173.315 126.435 174.125 ;
        RECT 126.445 173.315 127.815 174.125 ;
        RECT 14.805 173.105 14.975 173.315 ;
        RECT 16.240 173.155 16.360 173.265 ;
        RECT 18.485 173.125 18.655 173.315 ;
        RECT 21.705 173.105 21.875 173.295 ;
        RECT 22.165 173.105 22.335 173.295 ;
        RECT 24.005 173.125 24.175 173.315 ;
        RECT 28.145 173.125 28.315 173.315 ;
        RECT 32.010 173.125 32.180 173.315 ;
        RECT 32.285 173.105 32.455 173.295 ;
        RECT 33.665 173.105 33.835 173.315 ;
        RECT 34.125 173.125 34.295 173.315 ;
        RECT 35.505 173.105 35.675 173.295 ;
        RECT 35.965 173.105 36.135 173.295 ;
        RECT 38.080 173.105 38.250 173.295 ;
        RECT 44.245 173.125 44.415 173.315 ;
        RECT 45.165 173.160 45.325 173.270 ;
        RECT 49.030 173.125 49.200 173.315 ;
        RECT 49.820 173.155 49.940 173.265 ;
        RECT 50.685 173.105 50.855 173.315 ;
        RECT 52.985 173.125 53.155 173.315 ;
        RECT 53.445 173.105 53.615 173.295 ;
        RECT 53.960 173.155 54.080 173.265 ;
        RECT 56.665 173.105 56.835 173.295 ;
        RECT 56.850 173.125 57.020 173.315 ;
        RECT 57.640 173.155 57.760 173.265 ;
        RECT 59.425 173.105 59.595 173.295 ;
        RECT 59.940 173.155 60.060 173.265 ;
        RECT 61.265 173.125 61.435 173.315 ;
        RECT 62.645 173.105 62.815 173.295 ;
        RECT 64.025 173.150 64.185 173.260 ;
        RECT 65.865 173.105 66.035 173.295 ;
        RECT 66.325 173.105 66.495 173.295 ;
        RECT 66.785 173.125 66.955 173.315 ;
        RECT 67.345 173.295 67.415 173.315 ;
        RECT 67.245 173.125 67.415 173.295 ;
        RECT 68.220 173.155 68.340 173.265 ;
        RECT 70.005 173.105 70.175 173.295 ;
        RECT 70.465 173.105 70.635 173.315 ;
        RECT 79.205 173.295 79.275 173.315 ;
        RECT 71.845 173.125 72.015 173.295 ;
        RECT 75.525 173.160 75.685 173.270 ;
        RECT 71.945 173.105 72.015 173.125 ;
        RECT 75.985 173.105 76.155 173.295 ;
        RECT 76.445 173.105 76.615 173.295 ;
        RECT 79.205 173.125 79.375 173.295 ;
        RECT 79.665 173.125 79.835 173.315 ;
        RECT 82.480 173.155 82.600 173.265 ;
        RECT 85.185 173.125 85.355 173.315 ;
        RECT 85.645 173.125 85.815 173.315 ;
        RECT 87.945 173.125 88.115 173.315 ;
        RECT 88.405 173.105 88.575 173.295 ;
        RECT 88.865 173.160 89.025 173.270 ;
        RECT 89.380 173.155 89.500 173.265 ;
        RECT 91.165 173.105 91.335 173.295 ;
        RECT 91.625 173.125 91.795 173.315 ;
        RECT 92.140 173.155 92.260 173.265 ;
        RECT 92.545 173.125 92.715 173.315 ;
        RECT 96.685 173.105 96.855 173.295 ;
        RECT 100.550 173.105 100.720 173.295 ;
        RECT 101.745 173.150 101.905 173.260 ;
        RECT 103.125 173.105 103.295 173.295 ;
        RECT 108.645 173.105 108.815 173.295 ;
        RECT 109.110 173.105 109.280 173.295 ;
        RECT 112.780 173.125 112.950 173.315 ;
        RECT 113.300 173.155 113.420 173.265 ;
        RECT 114.165 173.105 114.335 173.295 ;
        RECT 115.085 173.265 115.255 173.315 ;
        RECT 115.085 173.155 115.260 173.265 ;
        RECT 115.085 173.125 115.255 173.155 ;
        RECT 115.545 173.105 115.715 173.295 ;
        RECT 118.950 173.125 119.120 173.315 ;
        RECT 119.685 173.125 119.855 173.315 ;
        RECT 121.525 173.160 121.685 173.270 ;
        RECT 121.985 173.125 122.155 173.315 ;
        RECT 123.420 173.155 123.540 173.265 ;
        RECT 125.665 173.105 125.835 173.295 ;
        RECT 126.125 173.265 126.295 173.315 ;
        RECT 126.125 173.155 126.300 173.265 ;
        RECT 126.125 173.125 126.295 173.155 ;
        RECT 127.505 173.105 127.675 173.315 ;
        RECT 14.665 172.295 16.035 173.105 ;
        RECT 16.505 172.295 22.015 173.105 ;
        RECT 22.035 172.195 23.385 173.105 ;
        RECT 23.405 172.425 32.595 173.105 ;
        RECT 23.405 172.195 24.325 172.425 ;
        RECT 27.155 172.205 28.085 172.425 ;
        RECT 32.605 172.325 33.975 173.105 ;
        RECT 33.985 172.295 35.815 173.105 ;
        RECT 35.825 172.325 37.195 173.105 ;
        RECT 37.215 172.235 37.645 173.020 ;
        RECT 37.665 172.425 41.565 173.105 ;
        RECT 41.890 172.425 50.995 173.105 ;
        RECT 37.665 172.195 38.595 172.425 ;
        RECT 51.665 172.295 53.755 173.105 ;
        RECT 54.225 172.295 56.975 173.105 ;
        RECT 56.995 172.425 59.735 173.105 ;
        RECT 60.205 172.295 62.955 173.105 ;
        RECT 62.975 172.235 63.405 173.020 ;
        RECT 64.345 172.425 66.175 173.105 ;
        RECT 66.185 172.425 68.015 173.105 ;
        RECT 64.345 172.195 65.690 172.425 ;
        RECT 66.670 172.195 68.015 172.425 ;
        RECT 68.485 172.295 70.315 173.105 ;
        RECT 70.335 172.195 71.685 173.105 ;
        RECT 71.945 172.875 74.215 173.105 ;
        RECT 71.945 172.195 74.700 172.875 ;
        RECT 74.925 172.295 76.295 173.105 ;
        RECT 76.305 172.425 79.045 173.105 ;
        RECT 79.435 172.425 88.715 173.105 ;
        RECT 79.435 172.305 81.770 172.425 ;
        RECT 79.435 172.195 80.355 172.305 ;
        RECT 86.435 172.205 87.355 172.425 ;
        RECT 88.735 172.235 89.165 173.020 ;
        RECT 89.645 172.295 91.475 173.105 ;
        RECT 91.485 172.295 96.995 173.105 ;
        RECT 97.235 172.425 101.135 173.105 ;
        RECT 100.205 172.195 101.135 172.425 ;
        RECT 102.065 172.325 103.435 173.105 ;
        RECT 103.445 172.295 108.955 173.105 ;
        RECT 108.965 172.195 112.440 173.105 ;
        RECT 112.645 172.295 114.475 173.105 ;
        RECT 114.495 172.235 114.925 173.020 ;
        RECT 115.405 172.325 116.775 173.105 ;
        RECT 116.785 172.425 125.975 173.105 ;
        RECT 116.785 172.195 117.705 172.425 ;
        RECT 120.535 172.205 121.465 172.425 ;
        RECT 126.445 172.295 127.815 173.105 ;
      LAYER nwell ;
        RECT 14.470 169.075 128.010 171.905 ;
      LAYER pwell ;
        RECT 14.665 167.875 16.035 168.685 ;
        RECT 16.045 167.875 21.555 168.685 ;
        RECT 21.575 167.875 22.925 168.785 ;
        RECT 22.945 167.875 24.315 168.685 ;
        RECT 24.335 167.960 24.765 168.745 ;
        RECT 25.245 167.875 27.995 168.685 ;
        RECT 28.005 167.875 33.515 168.685 ;
        RECT 33.525 167.875 39.035 168.685 ;
        RECT 39.185 167.875 41.795 168.785 ;
        RECT 42.920 167.875 46.395 168.785 ;
        RECT 46.405 167.875 49.880 168.785 ;
        RECT 50.095 167.960 50.525 168.745 ;
        RECT 50.545 167.875 51.915 168.685 ;
        RECT 51.925 167.875 55.400 168.785 ;
        RECT 56.065 167.875 61.575 168.685 ;
        RECT 61.595 167.875 64.335 168.555 ;
        RECT 64.345 167.875 65.715 168.685 ;
        RECT 66.210 168.555 67.555 168.785 ;
        RECT 65.725 167.875 67.555 168.555 ;
        RECT 68.485 167.875 71.205 168.785 ;
        RECT 71.285 167.875 75.835 168.785 ;
        RECT 75.855 167.960 76.285 168.745 ;
        RECT 76.305 167.875 78.135 168.685 ;
        RECT 78.145 167.875 83.655 168.685 ;
        RECT 86.865 168.555 87.795 168.785 ;
        RECT 83.895 167.875 87.795 168.555 ;
        RECT 87.815 167.875 89.165 168.785 ;
        RECT 89.185 167.875 90.555 168.655 ;
        RECT 90.565 167.875 91.935 168.685 ;
        RECT 91.945 167.875 97.455 168.685 ;
        RECT 100.665 168.555 101.595 168.785 ;
        RECT 97.695 167.875 101.595 168.555 ;
        RECT 101.615 167.960 102.045 168.745 ;
        RECT 102.985 167.875 104.355 168.655 ;
        RECT 104.825 167.875 108.300 168.785 ;
        RECT 108.505 167.875 110.335 168.685 ;
        RECT 113.545 168.555 114.475 168.785 ;
        RECT 110.575 167.875 114.475 168.555 ;
        RECT 114.855 168.675 115.775 168.785 ;
        RECT 114.855 168.555 117.190 168.675 ;
        RECT 121.855 168.555 122.775 168.775 ;
        RECT 114.855 167.875 124.135 168.555 ;
        RECT 124.145 167.875 125.975 168.555 ;
        RECT 126.445 167.875 127.815 168.685 ;
        RECT 14.805 167.665 14.975 167.875 ;
        RECT 17.565 167.665 17.735 167.855 ;
        RECT 21.245 167.685 21.415 167.875 ;
        RECT 22.625 167.685 22.795 167.875 ;
        RECT 24.005 167.685 24.175 167.875 ;
        RECT 24.980 167.715 25.100 167.825 ;
        RECT 26.765 167.665 26.935 167.855 ;
        RECT 27.685 167.685 27.855 167.875 ;
        RECT 28.605 167.665 28.775 167.855 ;
        RECT 33.205 167.685 33.375 167.875 ;
        RECT 34.125 167.665 34.295 167.855 ;
        RECT 36.885 167.665 37.055 167.855 ;
        RECT 37.805 167.665 37.975 167.855 ;
        RECT 38.725 167.685 38.895 167.875 ;
        RECT 39.645 167.710 39.805 167.820 ;
        RECT 41.480 167.685 41.650 167.875 ;
        RECT 42.405 167.720 42.565 167.830 ;
        RECT 43.320 167.665 43.490 167.855 ;
        RECT 46.080 167.685 46.250 167.875 ;
        RECT 46.550 167.685 46.720 167.875 ;
        RECT 47.000 167.665 47.170 167.855 ;
        RECT 50.680 167.665 50.850 167.855 ;
        RECT 51.150 167.665 51.320 167.855 ;
        RECT 51.605 167.685 51.775 167.875 ;
        RECT 52.070 167.685 52.240 167.875 ;
        RECT 55.800 167.715 55.920 167.825 ;
        RECT 57.120 167.665 57.290 167.855 ;
        RECT 57.640 167.715 57.760 167.825 ;
        RECT 61.265 167.665 61.435 167.875 ;
        RECT 61.725 167.665 61.895 167.855 ;
        RECT 63.620 167.715 63.740 167.825 ;
        RECT 64.025 167.685 64.195 167.875 ;
        RECT 65.405 167.665 65.575 167.875 ;
        RECT 65.865 167.665 66.035 167.875 ;
        RECT 68.165 167.710 68.325 167.830 ;
        RECT 68.625 167.685 68.795 167.875 ;
        RECT 73.685 167.665 73.855 167.855 ;
        RECT 75.525 167.665 75.695 167.875 ;
        RECT 76.040 167.715 76.160 167.825 ;
        RECT 77.825 167.685 77.995 167.875 ;
        RECT 83.345 167.855 83.515 167.875 ;
        RECT 79.660 167.665 79.830 167.855 ;
        RECT 83.340 167.685 83.515 167.855 ;
        RECT 83.860 167.715 83.980 167.825 ;
        RECT 83.340 167.665 83.510 167.685 ;
        RECT 84.540 167.665 84.710 167.855 ;
        RECT 87.210 167.685 87.380 167.875 ;
        RECT 88.460 167.715 88.580 167.825 ;
        RECT 88.865 167.685 89.035 167.875 ;
        RECT 90.245 167.685 90.415 167.875 ;
        RECT 91.625 167.685 91.795 167.875 ;
        RECT 92.545 167.665 92.715 167.855 ;
        RECT 93.005 167.665 93.175 167.855 ;
        RECT 94.845 167.710 95.005 167.820 ;
        RECT 95.305 167.665 95.475 167.855 ;
        RECT 97.145 167.685 97.315 167.875 ;
        RECT 101.010 167.685 101.180 167.875 ;
        RECT 102.665 167.720 102.825 167.830 ;
        RECT 103.125 167.685 103.295 167.875 ;
        RECT 104.560 167.715 104.680 167.825 ;
        RECT 104.970 167.685 105.140 167.875 ;
        RECT 105.885 167.665 106.055 167.855 ;
        RECT 107.725 167.665 107.895 167.855 ;
        RECT 108.190 167.665 108.360 167.855 ;
        RECT 110.025 167.685 110.195 167.875 ;
        RECT 113.890 167.685 114.060 167.875 ;
        RECT 114.165 167.665 114.335 167.855 ;
        RECT 115.545 167.710 115.705 167.820 ;
        RECT 116.005 167.665 116.175 167.855 ;
        RECT 119.680 167.665 119.850 167.855 ;
        RECT 120.605 167.710 120.765 167.820 ;
        RECT 123.825 167.685 123.995 167.875 ;
        RECT 125.665 167.685 125.835 167.875 ;
        RECT 126.125 167.825 126.295 167.855 ;
        RECT 126.125 167.715 126.300 167.825 ;
        RECT 126.125 167.665 126.295 167.715 ;
        RECT 127.505 167.665 127.675 167.875 ;
        RECT 14.665 166.855 16.035 167.665 ;
        RECT 16.045 166.855 17.875 167.665 ;
        RECT 17.885 166.985 27.075 167.665 ;
        RECT 17.885 166.755 18.805 166.985 ;
        RECT 21.635 166.765 22.565 166.985 ;
        RECT 27.085 166.855 28.915 167.665 ;
        RECT 28.925 166.855 34.435 167.665 ;
        RECT 34.455 166.985 37.195 167.665 ;
        RECT 37.215 166.795 37.645 167.580 ;
        RECT 37.665 166.885 39.035 167.665 ;
        RECT 40.160 166.755 43.635 167.665 ;
        RECT 43.840 166.755 47.315 167.665 ;
        RECT 47.520 166.755 50.995 167.665 ;
        RECT 51.005 166.755 54.480 167.665 ;
        RECT 54.825 166.755 57.435 167.665 ;
        RECT 57.905 166.855 61.575 167.665 ;
        RECT 61.595 166.755 62.945 167.665 ;
        RECT 62.975 166.795 63.405 167.580 ;
        RECT 63.885 166.855 65.715 167.665 ;
        RECT 65.725 166.985 67.555 167.665 ;
        RECT 66.210 166.755 67.555 166.985 ;
        RECT 68.485 166.855 73.995 167.665 ;
        RECT 74.005 166.985 75.835 167.665 ;
        RECT 74.005 166.755 75.350 166.985 ;
        RECT 76.500 166.755 79.975 167.665 ;
        RECT 80.180 166.755 83.655 167.665 ;
        RECT 84.125 166.985 88.025 167.665 ;
        RECT 84.125 166.755 85.055 166.985 ;
        RECT 88.735 166.795 89.165 167.580 ;
        RECT 89.185 166.855 92.855 167.665 ;
        RECT 92.865 166.885 94.235 167.665 ;
        RECT 95.175 166.755 96.525 167.665 ;
        RECT 96.915 166.985 106.195 167.665 ;
        RECT 96.915 166.865 99.250 166.985 ;
        RECT 96.915 166.755 97.835 166.865 ;
        RECT 103.915 166.765 104.835 166.985 ;
        RECT 106.205 166.855 108.035 167.665 ;
        RECT 108.045 166.755 111.520 167.665 ;
        RECT 111.725 166.855 114.475 167.665 ;
        RECT 114.495 166.795 114.925 167.580 ;
        RECT 115.875 166.755 117.225 167.665 ;
        RECT 117.385 166.755 119.995 167.665 ;
        RECT 120.925 166.855 126.435 167.665 ;
        RECT 126.445 166.855 127.815 167.665 ;
      LAYER nwell ;
        RECT 14.470 163.635 128.010 166.465 ;
      LAYER pwell ;
        RECT 14.665 162.435 16.035 163.245 ;
        RECT 16.505 162.435 20.175 163.245 ;
        RECT 23.385 163.115 24.315 163.345 ;
        RECT 20.415 162.435 24.315 163.115 ;
        RECT 24.335 162.520 24.765 163.305 ;
        RECT 24.785 162.435 26.155 163.215 ;
        RECT 26.625 162.435 28.455 163.245 ;
        RECT 28.475 162.435 29.825 163.345 ;
        RECT 29.855 162.435 31.205 163.345 ;
        RECT 31.225 163.115 32.145 163.345 ;
        RECT 34.975 163.115 35.905 163.335 ;
        RECT 31.225 162.435 40.415 163.115 ;
        RECT 41.080 162.435 44.555 163.345 ;
        RECT 44.760 162.435 48.235 163.345 ;
        RECT 48.245 162.435 50.075 163.245 ;
        RECT 50.095 162.520 50.525 163.305 ;
        RECT 50.545 162.435 54.215 163.245 ;
        RECT 54.225 162.435 59.735 163.245 ;
        RECT 60.115 163.235 61.035 163.345 ;
        RECT 60.115 163.115 62.450 163.235 ;
        RECT 67.115 163.115 68.035 163.335 ;
        RECT 60.115 162.435 69.395 163.115 ;
        RECT 70.325 162.435 73.995 163.245 ;
        RECT 74.005 163.115 75.350 163.345 ;
        RECT 74.005 162.435 75.835 163.115 ;
        RECT 75.855 162.520 76.285 163.305 ;
        RECT 76.305 162.435 79.055 163.245 ;
        RECT 79.065 162.435 82.540 163.345 ;
        RECT 83.575 163.235 84.495 163.345 ;
        RECT 83.575 163.115 85.910 163.235 ;
        RECT 90.575 163.115 91.495 163.335 ;
        RECT 92.865 163.115 93.795 163.345 ;
        RECT 83.575 162.435 92.855 163.115 ;
        RECT 92.865 162.435 96.765 163.115 ;
        RECT 97.925 162.435 101.400 163.345 ;
        RECT 101.615 162.520 102.045 163.305 ;
        RECT 102.525 162.435 108.035 163.245 ;
        RECT 108.045 162.435 111.520 163.345 ;
        RECT 111.725 162.435 115.200 163.345 ;
        RECT 115.405 162.435 120.915 163.245 ;
        RECT 120.925 162.435 126.435 163.245 ;
        RECT 126.445 162.435 127.815 163.245 ;
        RECT 14.805 162.225 14.975 162.435 ;
        RECT 16.240 162.275 16.360 162.385 ;
        RECT 16.645 162.270 16.805 162.380 ;
        RECT 19.865 162.245 20.035 162.435 ;
        RECT 23.730 162.245 23.900 162.435 ;
        RECT 24.925 162.245 25.095 162.435 ;
        RECT 25.845 162.225 26.015 162.415 ;
        RECT 26.360 162.275 26.480 162.385 ;
        RECT 28.145 162.245 28.315 162.435 ;
        RECT 28.605 162.245 28.775 162.435 ;
        RECT 29.985 162.245 30.155 162.435 ;
        RECT 35.045 162.225 35.215 162.415 ;
        RECT 36.885 162.245 37.055 162.415 ;
        RECT 38.080 162.225 38.250 162.415 ;
        RECT 40.105 162.245 40.275 162.435 ;
        RECT 40.620 162.275 40.740 162.385 ;
        RECT 42.405 162.270 42.565 162.380 ;
        RECT 44.240 162.245 44.410 162.435 ;
        RECT 47.920 162.415 48.090 162.435 ;
        RECT 47.920 162.245 48.095 162.415 ;
        RECT 47.925 162.225 48.095 162.245 ;
        RECT 48.390 162.225 48.560 162.415 ;
        RECT 49.765 162.245 49.935 162.435 ;
        RECT 53.905 162.245 54.075 162.435 ;
        RECT 57.125 162.225 57.295 162.415 ;
        RECT 58.505 162.225 58.675 162.415 ;
        RECT 59.425 162.245 59.595 162.435 ;
        RECT 62.370 162.225 62.540 162.415 ;
        RECT 63.620 162.275 63.740 162.385 ;
        RECT 64.025 162.225 64.195 162.415 ;
        RECT 68.165 162.225 68.335 162.415 ;
        RECT 69.085 162.245 69.255 162.435 ;
        RECT 70.005 162.280 70.165 162.390 ;
        RECT 72.765 162.225 72.935 162.415 ;
        RECT 73.685 162.245 73.855 162.435 ;
        RECT 74.605 162.225 74.775 162.415 ;
        RECT 75.525 162.245 75.695 162.435 ;
        RECT 75.985 162.225 76.155 162.415 ;
        RECT 78.745 162.245 78.915 162.435 ;
        RECT 79.210 162.245 79.380 162.435 ;
        RECT 79.665 162.225 79.835 162.415 ;
        RECT 82.940 162.275 83.060 162.385 ;
        RECT 83.340 162.225 83.510 162.415 ;
        RECT 84.265 162.270 84.425 162.380 ;
        RECT 84.725 162.225 84.895 162.415 ;
        RECT 87.025 162.225 87.195 162.415 ;
        RECT 87.485 162.225 87.655 162.415 ;
        RECT 92.545 162.245 92.715 162.435 ;
        RECT 93.280 162.245 93.450 162.435 ;
        RECT 97.605 162.280 97.765 162.390 ;
        RECT 98.070 162.245 98.240 162.435 ;
        RECT 98.525 162.225 98.695 162.415 ;
        RECT 102.205 162.385 102.375 162.415 ;
        RECT 102.205 162.275 102.380 162.385 ;
        RECT 102.205 162.225 102.375 162.275 ;
        RECT 105.880 162.225 106.050 162.415 ;
        RECT 107.725 162.245 107.895 162.435 ;
        RECT 108.190 162.245 108.360 162.435 ;
        RECT 108.645 162.225 108.815 162.415 ;
        RECT 111.870 162.245 112.040 162.435 ;
        RECT 114.165 162.225 114.335 162.415 ;
        RECT 118.305 162.225 118.475 162.415 ;
        RECT 118.765 162.225 118.935 162.415 ;
        RECT 120.605 162.245 120.775 162.435 ;
        RECT 126.125 162.225 126.295 162.435 ;
        RECT 127.505 162.225 127.675 162.435 ;
        RECT 14.665 161.415 16.035 162.225 ;
        RECT 16.965 161.545 26.155 162.225 ;
        RECT 26.250 161.545 35.355 162.225 ;
        RECT 35.365 161.545 36.730 162.225 ;
        RECT 16.965 161.315 17.885 161.545 ;
        RECT 20.715 161.325 21.645 161.545 ;
        RECT 37.215 161.355 37.645 162.140 ;
        RECT 37.665 161.545 41.565 162.225 ;
        RECT 37.665 161.315 38.595 161.545 ;
        RECT 42.725 161.415 48.235 162.225 ;
        RECT 48.245 161.315 51.720 162.225 ;
        RECT 51.925 161.415 57.435 162.225 ;
        RECT 57.455 161.315 58.805 162.225 ;
        RECT 59.055 161.545 62.955 162.225 ;
        RECT 62.025 161.315 62.955 161.545 ;
        RECT 62.975 161.355 63.405 162.140 ;
        RECT 63.885 161.445 65.255 162.225 ;
        RECT 65.265 161.315 68.475 162.225 ;
        RECT 69.405 161.415 73.075 162.225 ;
        RECT 73.085 161.545 74.915 162.225 ;
        RECT 73.085 161.315 74.430 161.545 ;
        RECT 74.925 161.415 76.295 162.225 ;
        RECT 76.305 161.415 79.975 162.225 ;
        RECT 80.180 161.315 83.655 162.225 ;
        RECT 84.585 161.445 85.955 162.225 ;
        RECT 85.975 161.315 87.325 162.225 ;
        RECT 87.355 161.315 88.705 162.225 ;
        RECT 88.735 161.355 89.165 162.140 ;
        RECT 89.555 161.545 98.835 162.225 ;
        RECT 89.555 161.425 91.890 161.545 ;
        RECT 89.555 161.315 90.475 161.425 ;
        RECT 96.555 161.325 97.475 161.545 ;
        RECT 98.845 161.415 102.515 162.225 ;
        RECT 102.720 161.315 106.195 162.225 ;
        RECT 106.205 161.415 108.955 162.225 ;
        RECT 108.965 161.415 114.475 162.225 ;
        RECT 114.495 161.355 114.925 162.140 ;
        RECT 114.945 161.415 118.615 162.225 ;
        RECT 118.635 161.315 119.985 162.225 ;
        RECT 120.925 161.415 126.435 162.225 ;
        RECT 126.445 161.415 127.815 162.225 ;
      LAYER nwell ;
        RECT 14.470 158.195 128.010 161.025 ;
      LAYER pwell ;
        RECT 14.665 156.995 16.035 157.805 ;
        RECT 16.045 156.995 17.415 157.805 ;
        RECT 17.435 156.995 18.785 157.905 ;
        RECT 18.815 156.995 20.165 157.905 ;
        RECT 23.385 157.675 24.315 157.905 ;
        RECT 20.415 156.995 24.315 157.675 ;
        RECT 24.335 157.080 24.765 157.865 ;
        RECT 24.785 156.995 26.155 157.775 ;
        RECT 26.625 156.995 30.295 157.805 ;
        RECT 30.675 157.795 31.595 157.905 ;
        RECT 30.675 157.675 33.010 157.795 ;
        RECT 37.675 157.675 38.595 157.895 ;
        RECT 30.675 156.995 39.955 157.675 ;
        RECT 39.965 156.995 41.335 157.775 ;
        RECT 41.345 156.995 42.715 157.805 ;
        RECT 42.725 156.995 46.395 157.805 ;
        RECT 46.405 156.995 49.880 157.905 ;
        RECT 50.095 157.080 50.525 157.865 ;
        RECT 51.005 156.995 52.835 157.805 ;
        RECT 52.845 156.995 58.355 157.805 ;
        RECT 58.735 157.795 59.655 157.905 ;
        RECT 58.735 157.675 61.070 157.795 ;
        RECT 65.735 157.675 66.655 157.895 ;
        RECT 68.945 157.675 70.290 157.905 ;
        RECT 70.785 157.675 72.130 157.905 ;
        RECT 73.110 157.675 74.455 157.905 ;
        RECT 58.735 156.995 68.015 157.675 ;
        RECT 68.945 156.995 70.775 157.675 ;
        RECT 70.785 156.995 72.615 157.675 ;
        RECT 72.625 156.995 74.455 157.675 ;
        RECT 74.465 156.995 75.835 157.805 ;
        RECT 75.855 157.080 76.285 157.865 ;
        RECT 76.790 157.675 78.135 157.905 ;
        RECT 76.305 156.995 78.135 157.675 ;
        RECT 78.145 156.995 79.515 157.805 ;
        RECT 79.525 156.995 85.035 157.805 ;
        RECT 85.045 156.995 90.555 157.805 ;
        RECT 90.565 156.995 96.075 157.805 ;
        RECT 96.085 156.995 101.595 157.805 ;
        RECT 101.615 157.080 102.045 157.865 ;
        RECT 103.180 156.995 106.655 157.905 ;
        RECT 107.585 157.705 108.530 157.905 ;
        RECT 107.585 157.025 110.335 157.705 ;
        RECT 107.585 156.995 108.530 157.025 ;
        RECT 14.805 156.785 14.975 156.995 ;
        RECT 17.105 156.805 17.275 156.995 ;
        RECT 17.565 156.785 17.735 156.975 ;
        RECT 18.485 156.805 18.655 156.995 ;
        RECT 18.945 156.805 19.115 156.995 ;
        RECT 23.730 156.805 23.900 156.995 ;
        RECT 25.845 156.805 26.015 156.995 ;
        RECT 26.360 156.835 26.480 156.945 ;
        RECT 26.765 156.785 26.935 156.975 ;
        RECT 28.145 156.785 28.315 156.975 ;
        RECT 29.065 156.830 29.225 156.940 ;
        RECT 29.985 156.805 30.155 156.995 ;
        RECT 32.745 156.785 32.915 156.975 ;
        RECT 36.610 156.785 36.780 156.975 ;
        RECT 38.725 156.785 38.895 156.975 ;
        RECT 39.645 156.805 39.815 156.995 ;
        RECT 41.025 156.805 41.195 156.995 ;
        RECT 42.405 156.785 42.575 156.995 ;
        RECT 14.665 155.975 16.035 156.785 ;
        RECT 16.045 155.975 17.875 156.785 ;
        RECT 17.885 156.105 27.075 156.785 ;
        RECT 17.885 155.875 18.805 156.105 ;
        RECT 21.635 155.885 22.565 156.105 ;
        RECT 27.085 156.005 28.455 156.785 ;
        RECT 29.385 155.975 33.055 156.785 ;
        RECT 33.295 156.105 37.195 156.785 ;
        RECT 36.265 155.875 37.195 156.105 ;
        RECT 37.215 155.915 37.645 156.700 ;
        RECT 37.665 155.975 39.035 156.785 ;
        RECT 39.045 155.975 42.715 156.785 ;
        RECT 42.725 156.755 43.670 156.785 ;
        RECT 45.160 156.755 45.330 156.975 ;
        RECT 45.630 156.785 45.800 156.975 ;
        RECT 46.085 156.805 46.255 156.995 ;
        RECT 46.550 156.805 46.720 156.995 ;
        RECT 52.525 156.975 52.695 156.995 ;
        RECT 50.740 156.835 50.860 156.945 ;
        RECT 52.520 156.805 52.695 156.975 ;
        RECT 53.445 156.830 53.605 156.940 ;
        RECT 58.045 156.805 58.215 156.995 ;
        RECT 52.520 156.785 52.690 156.805 ;
        RECT 58.965 156.785 59.135 156.975 ;
        RECT 62.640 156.785 62.810 156.975 ;
        RECT 64.485 156.785 64.655 156.975 ;
        RECT 64.945 156.785 65.115 156.975 ;
        RECT 67.705 156.805 67.875 156.995 ;
        RECT 68.625 156.840 68.785 156.950 ;
        RECT 70.465 156.805 70.635 156.995 ;
        RECT 72.305 156.805 72.475 156.995 ;
        RECT 72.765 156.805 72.935 156.995 ;
        RECT 75.525 156.785 75.695 156.995 ;
        RECT 76.445 156.805 76.615 156.995 ;
        RECT 77.365 156.785 77.535 156.975 ;
        RECT 79.205 156.805 79.375 156.995 ;
        RECT 82.885 156.785 83.055 156.975 ;
        RECT 84.725 156.805 84.895 156.995 ;
        RECT 88.405 156.785 88.575 156.975 ;
        RECT 89.785 156.830 89.945 156.940 ;
        RECT 90.245 156.805 90.415 156.995 ;
        RECT 93.465 156.785 93.635 156.975 ;
        RECT 93.925 156.785 94.095 156.975 ;
        RECT 95.360 156.835 95.480 156.945 ;
        RECT 95.765 156.805 95.935 156.995 ;
        RECT 97.145 156.785 97.315 156.975 ;
        RECT 97.610 156.785 97.780 156.975 ;
        RECT 101.285 156.945 101.455 156.995 ;
        RECT 101.285 156.835 101.460 156.945 ;
        RECT 102.665 156.840 102.825 156.950 ;
        RECT 101.285 156.805 101.455 156.835 ;
        RECT 104.960 156.785 105.130 156.975 ;
        RECT 106.340 156.805 106.510 156.995 ;
        RECT 110.020 156.975 110.190 157.025 ;
        RECT 110.345 156.995 113.820 157.905 ;
        RECT 114.025 156.995 115.395 157.805 ;
        RECT 115.405 157.675 116.325 157.905 ;
        RECT 119.155 157.675 120.085 157.895 ;
        RECT 115.405 156.995 124.595 157.675 ;
        RECT 124.605 156.995 126.435 157.805 ;
        RECT 126.445 156.995 127.815 157.805 ;
        RECT 107.265 156.840 107.425 156.950 ;
        RECT 108.640 156.785 108.810 156.975 ;
        RECT 110.020 156.805 110.195 156.975 ;
        RECT 110.490 156.805 110.660 156.995 ;
        RECT 110.025 156.785 110.195 156.805 ;
        RECT 113.890 156.785 114.060 156.975 ;
        RECT 115.085 156.945 115.255 156.995 ;
        RECT 115.085 156.835 115.260 156.945 ;
        RECT 115.085 156.805 115.255 156.835 ;
        RECT 115.545 156.785 115.715 156.975 ;
        RECT 124.285 156.805 124.455 156.995 ;
        RECT 126.125 156.785 126.295 156.995 ;
        RECT 127.505 156.785 127.675 156.995 ;
        RECT 42.725 156.075 45.475 156.755 ;
        RECT 42.725 155.875 43.670 156.075 ;
        RECT 45.485 155.875 48.960 156.785 ;
        RECT 49.360 155.875 52.835 156.785 ;
        RECT 53.765 155.975 59.275 156.785 ;
        RECT 59.480 155.875 62.955 156.785 ;
        RECT 62.975 155.915 63.405 156.700 ;
        RECT 63.425 155.975 64.795 156.785 ;
        RECT 64.815 155.875 66.165 156.785 ;
        RECT 66.555 156.105 75.835 156.785 ;
        RECT 75.845 156.105 77.675 156.785 ;
        RECT 66.555 155.985 68.890 156.105 ;
        RECT 66.555 155.875 67.475 155.985 ;
        RECT 73.555 155.885 74.475 156.105 ;
        RECT 75.845 155.875 77.190 156.105 ;
        RECT 77.685 155.975 83.195 156.785 ;
        RECT 83.205 155.975 88.715 156.785 ;
        RECT 88.735 155.915 89.165 156.700 ;
        RECT 90.105 155.975 93.775 156.785 ;
        RECT 93.785 156.005 95.155 156.785 ;
        RECT 95.625 155.975 97.455 156.785 ;
        RECT 97.465 155.875 100.940 156.785 ;
        RECT 101.800 155.875 105.275 156.785 ;
        RECT 105.480 155.875 108.955 156.785 ;
        RECT 108.965 155.975 110.335 156.785 ;
        RECT 110.575 156.105 114.475 156.785 ;
        RECT 113.545 155.875 114.475 156.105 ;
        RECT 114.495 155.915 114.925 156.700 ;
        RECT 115.415 155.875 116.765 156.785 ;
        RECT 117.155 156.105 126.435 156.785 ;
        RECT 117.155 155.985 119.490 156.105 ;
        RECT 117.155 155.875 118.075 155.985 ;
        RECT 124.155 155.885 125.075 156.105 ;
        RECT 126.445 155.975 127.815 156.785 ;
      LAYER nwell ;
        RECT 14.470 152.755 128.010 155.585 ;
      LAYER pwell ;
        RECT 14.665 151.555 16.035 152.365 ;
        RECT 16.505 151.555 20.175 152.365 ;
        RECT 23.385 152.235 24.315 152.465 ;
        RECT 20.415 151.555 24.315 152.235 ;
        RECT 24.335 151.640 24.765 152.425 ;
        RECT 24.785 151.555 26.155 152.365 ;
        RECT 26.165 151.555 29.835 152.365 ;
        RECT 29.845 151.555 35.355 152.365 ;
        RECT 38.565 152.235 39.495 152.465 ;
        RECT 35.595 151.555 39.495 152.235 ;
        RECT 39.965 151.555 43.635 152.365 ;
        RECT 43.645 152.265 44.590 152.465 ;
        RECT 43.645 151.585 46.395 152.265 ;
        RECT 43.645 151.555 44.590 151.585 ;
        RECT 14.805 151.345 14.975 151.555 ;
        RECT 16.240 151.395 16.360 151.505 ;
        RECT 19.865 151.365 20.035 151.555 ;
        RECT 23.730 151.365 23.900 151.555 ;
        RECT 25.385 151.345 25.555 151.535 ;
        RECT 25.845 151.505 26.015 151.555 ;
        RECT 25.845 151.395 26.020 151.505 ;
        RECT 25.845 151.365 26.015 151.395 ;
        RECT 27.685 151.345 27.855 151.535 ;
        RECT 28.145 151.345 28.315 151.535 ;
        RECT 29.525 151.365 29.695 151.555 ;
        RECT 35.045 151.365 35.215 151.555 ;
        RECT 38.265 151.390 38.425 151.500 ;
        RECT 38.910 151.365 39.080 151.555 ;
        RECT 39.645 151.505 39.815 151.535 ;
        RECT 39.645 151.395 39.820 151.505 ;
        RECT 39.645 151.345 39.815 151.395 ;
        RECT 40.565 151.390 40.725 151.500 ;
        RECT 43.325 151.365 43.495 151.555 ;
        RECT 46.080 151.535 46.250 151.585 ;
        RECT 46.600 151.555 50.075 152.465 ;
        RECT 50.095 151.640 50.525 152.425 ;
        RECT 50.545 151.555 54.020 152.465 ;
        RECT 54.685 151.555 58.355 152.365 ;
        RECT 58.365 151.555 61.840 152.465 ;
        RECT 62.505 151.555 65.255 152.365 ;
        RECT 68.465 152.235 69.395 152.465 ;
        RECT 65.495 151.555 69.395 152.235 ;
        RECT 69.405 151.555 70.775 152.335 ;
        RECT 74.490 152.235 75.835 152.465 ;
        RECT 70.795 151.555 73.535 152.235 ;
        RECT 74.005 151.555 75.835 152.235 ;
        RECT 75.855 151.640 76.285 152.425 ;
        RECT 76.305 151.555 79.025 152.465 ;
        RECT 79.065 151.555 81.815 152.365 ;
        RECT 81.825 151.555 84.565 152.235 ;
        RECT 85.045 151.555 86.875 152.365 ;
        RECT 86.895 151.555 88.245 152.465 ;
        RECT 88.265 152.235 89.185 152.465 ;
        RECT 92.015 152.235 92.945 152.455 ;
        RECT 88.265 151.555 97.455 152.235 ;
        RECT 97.925 151.555 101.595 152.365 ;
        RECT 101.615 151.640 102.045 152.425 ;
        RECT 102.720 151.555 106.195 152.465 ;
        RECT 106.205 151.555 109.680 152.465 ;
        RECT 111.000 151.555 114.475 152.465 ;
        RECT 114.485 151.555 116.315 152.365 ;
        RECT 119.525 152.235 120.455 152.465 ;
        RECT 116.555 151.555 120.455 152.235 ;
        RECT 120.465 151.555 121.835 152.335 ;
        RECT 121.845 151.555 123.215 152.335 ;
        RECT 123.685 151.555 126.435 152.365 ;
        RECT 126.445 151.555 127.815 152.365 ;
        RECT 46.080 151.365 46.255 151.535 ;
        RECT 46.085 151.345 46.255 151.365 ;
        RECT 14.665 150.535 16.035 151.345 ;
        RECT 16.505 150.665 25.695 151.345 ;
        RECT 16.505 150.435 17.425 150.665 ;
        RECT 20.255 150.445 21.185 150.665 ;
        RECT 26.165 150.535 27.995 151.345 ;
        RECT 28.005 150.665 37.195 151.345 ;
        RECT 32.515 150.445 33.445 150.665 ;
        RECT 36.275 150.435 37.195 150.665 ;
        RECT 37.215 150.475 37.645 151.260 ;
        RECT 38.585 150.565 39.955 151.345 ;
        RECT 40.885 150.535 46.395 151.345 ;
        RECT 46.405 151.315 47.350 151.345 ;
        RECT 48.840 151.315 49.010 151.535 ;
        RECT 49.760 151.365 49.930 151.555 ;
        RECT 50.690 151.365 50.860 151.555 ;
        RECT 49.165 151.315 50.110 151.345 ;
        RECT 51.600 151.315 51.770 151.535 ;
        RECT 54.365 151.505 54.535 151.535 ;
        RECT 54.365 151.395 54.540 151.505 ;
        RECT 54.365 151.345 54.535 151.395 ;
        RECT 54.830 151.345 55.000 151.535 ;
        RECT 58.045 151.365 58.215 151.555 ;
        RECT 58.510 151.345 58.680 151.555 ;
        RECT 62.240 151.395 62.360 151.505 ;
        RECT 62.645 151.390 62.805 151.500 ;
        RECT 64.945 151.365 65.115 151.555 ;
        RECT 68.810 151.365 68.980 151.555 ;
        RECT 69.545 151.365 69.715 151.555 ;
        RECT 72.305 151.345 72.475 151.535 ;
        RECT 73.225 151.365 73.395 151.555 ;
        RECT 73.740 151.395 73.860 151.505 ;
        RECT 74.145 151.345 74.315 151.555 ;
        RECT 75.985 151.345 76.155 151.535 ;
        RECT 76.445 151.505 76.615 151.555 ;
        RECT 76.445 151.395 76.620 151.505 ;
        RECT 76.445 151.365 76.615 151.395 ;
        RECT 80.120 151.345 80.290 151.535 ;
        RECT 80.590 151.345 80.760 151.535 ;
        RECT 81.505 151.365 81.675 151.555 ;
        RECT 81.965 151.365 82.135 151.555 ;
        RECT 84.780 151.500 84.900 151.505 ;
        RECT 84.725 151.395 84.900 151.500 ;
        RECT 84.725 151.390 84.885 151.395 ;
        RECT 86.565 151.365 86.735 151.555 ;
        RECT 87.025 151.365 87.195 151.555 ;
        RECT 88.405 151.345 88.575 151.535 ;
        RECT 92.730 151.345 92.900 151.535 ;
        RECT 94.385 151.345 94.555 151.535 ;
        RECT 97.145 151.365 97.315 151.555 ;
        RECT 97.660 151.395 97.780 151.505 ;
        RECT 98.065 151.345 98.235 151.535 ;
        RECT 101.285 151.365 101.455 151.555 ;
        RECT 102.260 151.395 102.380 151.505 ;
        RECT 103.585 151.345 103.755 151.535 ;
        RECT 46.405 150.635 49.155 151.315 ;
        RECT 49.165 150.635 51.915 151.315 ;
        RECT 46.405 150.435 47.350 150.635 ;
        RECT 49.165 150.435 50.110 150.635 ;
        RECT 51.925 150.535 54.675 151.345 ;
        RECT 54.685 150.435 58.160 151.345 ;
        RECT 58.365 150.435 61.840 151.345 ;
        RECT 62.975 150.475 63.405 151.260 ;
        RECT 63.510 150.665 72.615 151.345 ;
        RECT 72.625 150.665 74.455 151.345 ;
        RECT 74.465 150.665 76.295 151.345 ;
        RECT 72.625 150.435 73.970 150.665 ;
        RECT 74.465 150.435 75.810 150.665 ;
        RECT 76.960 150.435 80.435 151.345 ;
        RECT 80.445 150.435 83.920 151.345 ;
        RECT 85.045 150.535 88.715 151.345 ;
        RECT 88.735 150.475 89.165 151.260 ;
        RECT 89.415 150.665 93.315 151.345 ;
        RECT 92.385 150.435 93.315 150.665 ;
        RECT 93.325 150.535 94.695 151.345 ;
        RECT 94.705 150.535 98.375 151.345 ;
        RECT 98.385 150.535 103.895 151.345 ;
        RECT 104.050 151.315 104.220 151.535 ;
        RECT 105.880 151.365 106.050 151.555 ;
        RECT 106.350 151.365 106.520 151.555 ;
        RECT 114.160 151.535 114.330 151.555 ;
        RECT 109.105 151.345 109.275 151.535 ;
        RECT 105.710 151.315 106.655 151.345 ;
        RECT 103.905 150.635 106.655 151.315 ;
        RECT 105.710 150.435 106.655 150.635 ;
        RECT 106.665 150.535 109.415 151.345 ;
        RECT 109.570 151.315 109.740 151.535 ;
        RECT 110.485 151.400 110.645 151.510 ;
        RECT 112.380 151.395 112.500 151.505 ;
        RECT 114.160 151.365 114.335 151.535 ;
        RECT 115.140 151.395 115.260 151.505 ;
        RECT 116.005 151.365 116.175 151.555 ;
        RECT 119.870 151.365 120.040 151.555 ;
        RECT 114.165 151.345 114.335 151.365 ;
        RECT 120.605 151.345 120.775 151.555 ;
        RECT 121.985 151.365 122.155 151.555 ;
        RECT 123.420 151.395 123.540 151.505 ;
        RECT 126.125 151.345 126.295 151.555 ;
        RECT 127.505 151.345 127.675 151.555 ;
        RECT 111.230 151.315 112.175 151.345 ;
        RECT 109.425 150.635 112.175 151.315 ;
        RECT 111.230 150.435 112.175 150.635 ;
        RECT 112.645 150.535 114.475 151.345 ;
        RECT 114.495 150.475 114.925 151.260 ;
        RECT 115.405 150.535 120.915 151.345 ;
        RECT 120.925 150.535 126.435 151.345 ;
        RECT 126.445 150.535 127.815 151.345 ;
      LAYER nwell ;
        RECT 14.470 147.315 128.010 150.145 ;
      LAYER pwell ;
        RECT 14.665 146.115 16.035 146.925 ;
        RECT 16.045 146.115 18.795 146.925 ;
        RECT 18.815 146.115 20.165 147.025 ;
        RECT 23.385 146.795 24.315 147.025 ;
        RECT 20.415 146.115 24.315 146.795 ;
        RECT 24.335 146.200 24.765 146.985 ;
        RECT 25.245 146.115 27.075 146.925 ;
        RECT 27.085 146.115 32.595 146.925 ;
        RECT 32.615 146.115 33.965 147.025 ;
        RECT 33.985 146.115 35.355 146.895 ;
        RECT 36.285 146.115 41.795 146.925 ;
        RECT 41.805 146.115 44.415 147.025 ;
        RECT 44.565 146.115 50.075 146.925 ;
        RECT 50.095 146.200 50.525 146.985 ;
        RECT 51.005 146.115 54.675 146.925 ;
        RECT 54.685 146.115 60.195 146.925 ;
        RECT 60.215 146.115 61.565 147.025 ;
        RECT 62.045 146.115 64.795 146.925 ;
        RECT 64.805 146.115 66.175 146.895 ;
        RECT 66.185 146.115 67.555 146.925 ;
        RECT 67.565 146.115 71.235 146.925 ;
        RECT 71.730 146.795 73.075 147.025 ;
        RECT 74.030 146.795 75.375 147.025 ;
        RECT 71.245 146.115 73.075 146.795 ;
        RECT 73.545 146.115 75.375 146.795 ;
        RECT 75.855 146.200 76.285 146.985 ;
        RECT 76.790 146.795 78.135 147.025 ;
        RECT 76.305 146.115 78.135 146.795 ;
        RECT 78.800 146.115 82.275 147.025 ;
        RECT 82.285 146.115 85.760 147.025 ;
        RECT 86.885 146.115 92.395 146.925 ;
        RECT 92.415 146.115 93.765 147.025 ;
        RECT 93.785 146.115 95.155 146.925 ;
        RECT 95.165 146.825 96.110 147.025 ;
        RECT 95.165 146.145 97.915 146.825 ;
        RECT 95.165 146.115 96.110 146.145 ;
        RECT 14.805 145.905 14.975 146.115 ;
        RECT 16.645 145.950 16.805 146.060 ;
        RECT 17.105 145.905 17.275 146.095 ;
        RECT 18.485 145.925 18.655 146.115 ;
        RECT 19.865 145.925 20.035 146.115 ;
        RECT 23.730 145.925 23.900 146.115 ;
        RECT 24.980 145.955 25.100 146.065 ;
        RECT 26.765 145.925 26.935 146.115 ;
        RECT 27.225 145.905 27.395 146.095 ;
        RECT 32.285 145.925 32.455 146.115 ;
        RECT 32.745 145.925 32.915 146.115 ;
        RECT 34.125 145.925 34.295 146.115 ;
        RECT 35.965 145.960 36.125 146.070 ;
        RECT 36.425 145.905 36.595 146.095 ;
        RECT 36.940 145.955 37.060 146.065 ;
        RECT 41.210 145.905 41.380 146.095 ;
        RECT 41.485 145.925 41.655 146.115 ;
        RECT 41.950 145.925 42.120 146.115 ;
        RECT 45.620 145.905 45.790 146.095 ;
        RECT 46.090 145.905 46.260 146.095 ;
        RECT 49.765 146.065 49.935 146.115 ;
        RECT 49.765 145.955 49.940 146.065 ;
        RECT 50.740 145.955 50.860 146.065 ;
        RECT 49.765 145.925 49.935 145.955 ;
        RECT 53.445 145.905 53.615 146.095 ;
        RECT 54.365 145.925 54.535 146.115 ;
        RECT 59.885 145.925 60.055 146.115 ;
        RECT 61.265 145.925 61.435 146.115 ;
        RECT 61.780 145.955 61.900 146.065 ;
        RECT 62.645 145.905 62.815 146.095 ;
        RECT 63.840 145.905 64.010 146.095 ;
        RECT 64.485 145.925 64.655 146.115 ;
        RECT 65.865 145.925 66.035 146.115 ;
        RECT 67.245 145.925 67.415 146.115 ;
        RECT 67.705 145.905 67.875 146.095 ;
        RECT 69.140 145.955 69.260 146.065 ;
        RECT 69.545 145.905 69.715 146.095 ;
        RECT 70.925 145.925 71.095 146.115 ;
        RECT 71.385 145.925 71.555 146.115 ;
        RECT 73.280 145.955 73.400 146.065 ;
        RECT 73.685 145.925 73.855 146.115 ;
        RECT 74.145 145.905 74.315 146.095 ;
        RECT 75.580 145.955 75.700 146.065 ;
        RECT 76.445 145.925 76.615 146.115 ;
        RECT 78.340 145.955 78.460 146.065 ;
        RECT 79.665 145.905 79.835 146.095 ;
        RECT 80.130 145.905 80.300 146.095 ;
        RECT 81.960 145.925 82.130 146.115 ;
        RECT 82.430 145.925 82.600 146.115 ;
        RECT 84.265 145.950 84.425 146.060 ;
        RECT 86.565 145.960 86.725 146.070 ;
        RECT 88.130 145.905 88.300 146.095 ;
        RECT 92.085 145.925 92.255 146.115 ;
        RECT 93.465 145.925 93.635 146.115 ;
        RECT 94.845 145.925 95.015 146.115 ;
        RECT 97.600 145.925 97.770 146.145 ;
        RECT 97.925 146.115 101.400 147.025 ;
        RECT 101.615 146.200 102.045 146.985 ;
        RECT 102.065 146.115 107.575 146.925 ;
        RECT 109.390 146.825 110.335 147.025 ;
        RECT 107.585 146.145 110.335 146.825 ;
        RECT 98.070 145.925 98.240 146.115 ;
        RECT 98.525 145.905 98.695 146.095 ;
        RECT 99.040 145.955 99.160 146.065 ;
        RECT 104.505 145.905 104.675 146.095 ;
        RECT 14.665 145.095 16.035 145.905 ;
        RECT 16.965 145.125 18.335 145.905 ;
        RECT 18.345 145.225 27.535 145.905 ;
        RECT 27.545 145.225 36.735 145.905 ;
        RECT 18.345 144.995 19.265 145.225 ;
        RECT 22.095 145.005 23.025 145.225 ;
        RECT 27.545 144.995 28.465 145.225 ;
        RECT 31.295 145.005 32.225 145.225 ;
        RECT 37.215 145.035 37.645 145.820 ;
        RECT 37.895 145.225 41.795 145.905 ;
        RECT 40.865 144.995 41.795 145.225 ;
        RECT 42.460 144.995 45.935 145.905 ;
        RECT 45.945 144.995 49.420 145.905 ;
        RECT 50.085 145.095 53.755 145.905 ;
        RECT 53.765 145.225 62.955 145.905 ;
        RECT 53.765 144.995 54.685 145.225 ;
        RECT 57.515 145.005 58.445 145.225 ;
        RECT 62.975 145.035 63.405 145.820 ;
        RECT 63.425 145.225 67.325 145.905 ;
        RECT 63.425 144.995 64.355 145.225 ;
        RECT 67.575 144.995 68.925 145.905 ;
        RECT 69.405 145.125 70.775 145.905 ;
        RECT 70.785 145.095 74.455 145.905 ;
        RECT 74.465 145.095 79.975 145.905 ;
        RECT 79.985 144.995 83.460 145.905 ;
        RECT 84.815 145.225 88.715 145.905 ;
        RECT 87.785 144.995 88.715 145.225 ;
        RECT 88.735 145.035 89.165 145.820 ;
        RECT 89.555 145.225 98.835 145.905 ;
        RECT 89.555 145.105 91.890 145.225 ;
        RECT 89.555 144.995 90.475 145.105 ;
        RECT 96.555 145.005 97.475 145.225 ;
        RECT 99.305 145.095 104.815 145.905 ;
        RECT 104.970 145.875 105.140 146.095 ;
        RECT 107.265 145.925 107.435 146.115 ;
        RECT 107.730 145.905 107.900 146.145 ;
        RECT 109.390 146.115 110.335 146.145 ;
        RECT 110.345 146.115 113.820 147.025 ;
        RECT 114.485 146.115 116.315 146.925 ;
        RECT 119.525 146.795 120.455 147.025 ;
        RECT 116.555 146.115 120.455 146.795 ;
        RECT 120.465 146.115 121.835 146.925 ;
        RECT 121.845 146.115 123.215 146.895 ;
        RECT 123.685 146.115 126.435 146.925 ;
        RECT 126.445 146.115 127.815 146.925 ;
        RECT 110.490 145.925 110.660 146.115 ;
        RECT 111.460 145.955 111.580 146.065 ;
        RECT 111.870 145.905 112.040 146.095 ;
        RECT 114.220 145.955 114.340 146.065 ;
        RECT 115.140 145.955 115.260 146.065 ;
        RECT 115.545 145.905 115.715 146.095 ;
        RECT 116.005 145.925 116.175 146.115 ;
        RECT 119.870 145.925 120.040 146.115 ;
        RECT 121.525 145.925 121.695 146.115 ;
        RECT 121.985 145.925 122.155 146.115 ;
        RECT 123.420 145.955 123.540 146.065 ;
        RECT 126.125 145.905 126.295 146.115 ;
        RECT 127.505 145.905 127.675 146.115 ;
        RECT 106.630 145.875 107.575 145.905 ;
        RECT 104.825 145.195 107.575 145.875 ;
        RECT 106.630 144.995 107.575 145.195 ;
        RECT 107.585 144.995 111.060 145.905 ;
        RECT 111.725 144.995 114.335 145.905 ;
        RECT 114.495 145.035 114.925 145.820 ;
        RECT 115.415 144.995 116.765 145.905 ;
        RECT 117.155 145.225 126.435 145.905 ;
        RECT 117.155 145.105 119.490 145.225 ;
        RECT 117.155 144.995 118.075 145.105 ;
        RECT 124.155 145.005 125.075 145.225 ;
        RECT 126.445 145.095 127.815 145.905 ;
      LAYER nwell ;
        RECT 14.470 141.875 128.010 144.705 ;
      LAYER pwell ;
        RECT 14.665 140.675 16.035 141.485 ;
        RECT 16.045 140.675 18.795 141.485 ;
        RECT 18.815 140.675 20.165 141.585 ;
        RECT 20.185 141.355 21.115 141.585 ;
        RECT 20.185 140.675 24.085 141.355 ;
        RECT 24.335 140.760 24.765 141.545 ;
        RECT 25.245 140.675 26.615 141.455 ;
        RECT 26.625 140.675 29.375 141.485 ;
        RECT 29.395 140.675 30.745 141.585 ;
        RECT 30.775 140.675 32.125 141.585 ;
        RECT 32.145 141.355 33.065 141.585 ;
        RECT 35.895 141.355 36.825 141.575 ;
        RECT 32.145 140.675 41.335 141.355 ;
        RECT 41.345 140.675 42.715 141.455 ;
        RECT 42.920 140.675 46.395 141.585 ;
        RECT 46.600 140.675 50.075 141.585 ;
        RECT 50.095 140.760 50.525 141.545 ;
        RECT 52.350 141.385 53.295 141.585 ;
        RECT 50.545 140.705 53.295 141.385 ;
        RECT 14.805 140.465 14.975 140.675 ;
        RECT 16.240 140.515 16.360 140.625 ;
        RECT 18.485 140.485 18.655 140.675 ;
        RECT 19.865 140.485 20.035 140.675 ;
        RECT 20.600 140.485 20.770 140.675 ;
        RECT 21.705 140.465 21.875 140.655 ;
        RECT 24.980 140.515 25.100 140.625 ;
        RECT 25.385 140.485 25.555 140.675 ;
        RECT 27.225 140.465 27.395 140.655 ;
        RECT 29.065 140.485 29.235 140.675 ;
        RECT 29.525 140.485 29.695 140.675 ;
        RECT 30.905 140.485 31.075 140.675 ;
        RECT 32.745 140.465 32.915 140.655 ;
        RECT 33.480 140.465 33.650 140.655 ;
        RECT 41.025 140.485 41.195 140.675 ;
        RECT 42.405 140.485 42.575 140.675 ;
        RECT 46.080 140.655 46.250 140.675 ;
        RECT 42.865 140.465 43.035 140.655 ;
        RECT 14.665 139.655 16.035 140.465 ;
        RECT 16.505 139.655 22.015 140.465 ;
        RECT 22.025 139.655 27.535 140.465 ;
        RECT 27.545 139.655 33.055 140.465 ;
        RECT 33.065 139.785 36.965 140.465 ;
        RECT 33.065 139.555 33.995 139.785 ;
        RECT 37.215 139.595 37.645 140.380 ;
        RECT 37.665 139.655 43.175 140.465 ;
        RECT 43.185 140.435 44.130 140.465 ;
        RECT 45.620 140.435 45.790 140.655 ;
        RECT 46.080 140.485 46.260 140.655 ;
        RECT 49.760 140.625 49.930 140.675 ;
        RECT 49.760 140.515 49.940 140.625 ;
        RECT 49.760 140.485 49.930 140.515 ;
        RECT 50.690 140.485 50.860 140.705 ;
        RECT 52.350 140.675 53.295 140.705 ;
        RECT 53.305 140.675 56.055 141.485 ;
        RECT 56.065 140.675 59.540 141.585 ;
        RECT 63.865 141.355 64.795 141.585 ;
        RECT 60.895 140.675 64.795 141.355 ;
        RECT 65.175 141.475 66.095 141.585 ;
        RECT 65.175 141.355 67.510 141.475 ;
        RECT 72.175 141.355 73.095 141.575 ;
        RECT 65.175 140.675 74.455 141.355 ;
        RECT 74.465 140.675 75.835 141.485 ;
        RECT 75.855 140.760 76.285 141.545 ;
        RECT 76.305 141.385 77.250 141.585 ;
        RECT 79.065 141.385 80.010 141.585 ;
        RECT 76.305 140.705 79.055 141.385 ;
        RECT 79.065 140.705 81.815 141.385 ;
        RECT 76.305 140.675 77.250 140.705 ;
        RECT 46.090 140.465 46.260 140.485 ;
        RECT 51.605 140.465 51.775 140.655 ;
        RECT 55.745 140.485 55.915 140.675 ;
        RECT 56.210 140.485 56.380 140.675 ;
        RECT 57.125 140.465 57.295 140.655 ;
        RECT 57.590 140.465 57.760 140.655 ;
        RECT 60.345 140.520 60.505 140.630 ;
        RECT 62.645 140.465 62.815 140.655 ;
        RECT 64.210 140.485 64.380 140.675 ;
        RECT 64.485 140.465 64.655 140.655 ;
        RECT 68.165 140.465 68.335 140.655 ;
        RECT 68.625 140.465 68.795 140.655 ;
        RECT 70.925 140.465 71.095 140.655 ;
        RECT 71.385 140.465 71.555 140.655 ;
        RECT 73.685 140.465 73.855 140.655 ;
        RECT 74.145 140.485 74.315 140.675 ;
        RECT 75.525 140.485 75.695 140.675 ;
        RECT 77.365 140.465 77.535 140.655 ;
        RECT 78.740 140.485 78.910 140.705 ;
        RECT 79.065 140.675 80.010 140.705 ;
        RECT 81.500 140.485 81.670 140.705 ;
        RECT 81.825 140.675 85.300 141.585 ;
        RECT 85.965 140.675 91.475 141.485 ;
        RECT 91.485 140.675 92.855 141.455 ;
        RECT 92.865 140.675 94.235 141.455 ;
        RECT 94.245 140.675 96.075 141.485 ;
        RECT 96.085 140.675 101.595 141.485 ;
        RECT 101.615 140.760 102.045 141.545 ;
        RECT 102.065 140.675 103.435 141.485 ;
        RECT 103.445 140.675 107.115 141.485 ;
        RECT 110.325 141.355 111.255 141.585 ;
        RECT 107.355 140.675 111.255 141.355 ;
        RECT 111.725 140.675 113.555 141.485 ;
        RECT 113.575 140.675 114.925 141.585 ;
        RECT 115.315 141.475 116.235 141.585 ;
        RECT 115.315 141.355 117.650 141.475 ;
        RECT 122.315 141.355 123.235 141.575 ;
        RECT 115.315 140.675 124.595 141.355 ;
        RECT 124.605 140.675 126.435 141.485 ;
        RECT 126.445 140.675 127.815 141.485 ;
        RECT 81.970 140.485 82.140 140.675 ;
        RECT 82.885 140.465 83.055 140.655 ;
        RECT 85.700 140.515 85.820 140.625 ;
        RECT 88.405 140.465 88.575 140.655 ;
        RECT 91.165 140.485 91.335 140.675 ;
        RECT 91.625 140.485 91.795 140.675 ;
        RECT 93.005 140.485 93.175 140.675 ;
        RECT 95.765 140.485 95.935 140.675 ;
        RECT 98.525 140.465 98.695 140.655 ;
        RECT 99.445 140.510 99.605 140.620 ;
        RECT 101.285 140.485 101.455 140.675 ;
        RECT 103.125 140.465 103.295 140.675 ;
        RECT 106.805 140.485 106.975 140.675 ;
        RECT 110.670 140.485 110.840 140.675 ;
        RECT 111.460 140.515 111.580 140.625 ;
        RECT 112.785 140.465 112.955 140.655 ;
        RECT 113.245 140.485 113.415 140.675 ;
        RECT 113.705 140.485 113.875 140.675 ;
        RECT 114.165 140.465 114.335 140.655 ;
        RECT 115.140 140.515 115.260 140.625 ;
        RECT 118.950 140.465 119.120 140.655 ;
        RECT 119.740 140.515 119.860 140.625 ;
        RECT 120.145 140.465 120.315 140.655 ;
        RECT 122.445 140.465 122.615 140.655 ;
        RECT 124.285 140.485 124.455 140.675 ;
        RECT 126.125 140.465 126.295 140.675 ;
        RECT 127.505 140.465 127.675 140.675 ;
        RECT 43.185 139.755 45.935 140.435 ;
        RECT 43.185 139.555 44.130 139.755 ;
        RECT 45.945 139.555 49.420 140.465 ;
        RECT 50.085 139.655 51.915 140.465 ;
        RECT 51.925 139.655 57.435 140.465 ;
        RECT 57.445 139.555 60.920 140.465 ;
        RECT 61.125 139.655 62.955 140.465 ;
        RECT 62.975 139.595 63.405 140.380 ;
        RECT 63.425 139.655 64.795 140.465 ;
        RECT 64.805 139.655 68.475 140.465 ;
        RECT 68.495 139.555 69.845 140.465 ;
        RECT 69.865 139.655 71.235 140.465 ;
        RECT 71.245 139.685 72.615 140.465 ;
        RECT 72.625 139.655 73.995 140.465 ;
        RECT 74.005 139.655 77.675 140.465 ;
        RECT 77.685 139.655 83.195 140.465 ;
        RECT 83.205 139.655 88.715 140.465 ;
        RECT 88.735 139.595 89.165 140.380 ;
        RECT 89.555 139.785 98.835 140.465 ;
        RECT 89.555 139.665 91.890 139.785 ;
        RECT 89.555 139.555 90.475 139.665 ;
        RECT 96.555 139.565 97.475 139.785 ;
        RECT 99.765 139.655 103.435 140.465 ;
        RECT 103.815 139.785 113.095 140.465 ;
        RECT 103.815 139.665 106.150 139.785 ;
        RECT 103.815 139.555 104.735 139.665 ;
        RECT 110.815 139.565 111.735 139.785 ;
        RECT 113.105 139.655 114.475 140.465 ;
        RECT 114.495 139.595 114.925 140.380 ;
        RECT 115.635 139.785 119.535 140.465 ;
        RECT 118.605 139.555 119.535 139.785 ;
        RECT 120.005 139.685 121.375 140.465 ;
        RECT 121.385 139.655 122.755 140.465 ;
        RECT 122.765 139.655 126.435 140.465 ;
        RECT 126.445 139.655 127.815 140.465 ;
      LAYER nwell ;
        RECT 14.470 136.435 128.010 139.265 ;
      LAYER pwell ;
        RECT 14.665 135.235 16.035 136.045 ;
        RECT 16.045 135.235 18.795 136.045 ;
        RECT 18.805 135.235 24.315 136.045 ;
        RECT 24.335 135.320 24.765 136.105 ;
        RECT 48.465 136.055 49.415 136.145 ;
        RECT 25.245 135.235 30.755 136.045 ;
        RECT 30.765 135.235 36.275 136.045 ;
        RECT 36.285 135.235 41.795 136.045 ;
        RECT 41.805 135.235 47.315 136.045 ;
        RECT 47.485 135.235 49.415 136.055 ;
        RECT 50.095 135.320 50.525 136.105 ;
        RECT 51.005 135.235 56.515 136.045 ;
        RECT 56.525 135.235 62.035 136.045 ;
        RECT 65.245 135.915 66.175 136.145 ;
        RECT 62.275 135.235 66.175 135.915 ;
        RECT 66.555 136.035 67.475 136.145 ;
        RECT 66.555 135.915 68.890 136.035 ;
        RECT 73.555 135.915 74.475 136.135 ;
        RECT 66.555 135.235 75.835 135.915 ;
        RECT 75.855 135.320 76.285 136.105 ;
        RECT 77.225 135.235 80.895 136.045 ;
        RECT 82.710 135.945 83.655 136.145 ;
        RECT 80.905 135.265 83.655 135.945 ;
        RECT 14.805 135.025 14.975 135.235 ;
        RECT 16.240 135.075 16.360 135.185 ;
        RECT 18.025 135.025 18.195 135.215 ;
        RECT 18.485 135.045 18.655 135.235 ;
        RECT 23.545 135.025 23.715 135.215 ;
        RECT 24.005 135.045 24.175 135.235 ;
        RECT 24.980 135.075 25.100 135.185 ;
        RECT 30.445 135.045 30.615 135.235 ;
        RECT 33.205 135.025 33.375 135.215 ;
        RECT 34.585 135.025 34.755 135.215 ;
        RECT 35.045 135.025 35.215 135.215 ;
        RECT 35.965 135.045 36.135 135.235 ;
        RECT 36.885 135.070 37.045 135.180 ;
        RECT 40.105 135.025 40.275 135.215 ;
        RECT 40.565 135.045 40.735 135.215 ;
        RECT 41.485 135.045 41.655 135.235 ;
        RECT 42.865 135.045 43.035 135.215 ;
        RECT 40.585 135.025 40.735 135.045 ;
        RECT 42.885 135.025 43.035 135.045 ;
        RECT 47.005 135.045 47.175 135.235 ;
        RECT 47.485 135.215 47.635 135.235 ;
        RECT 47.465 135.045 47.640 135.215 ;
        RECT 49.820 135.075 49.940 135.185 ;
        RECT 50.740 135.075 50.860 135.185 ;
        RECT 47.005 135.025 47.155 135.045 ;
        RECT 14.665 134.215 16.035 135.025 ;
        RECT 16.505 134.215 18.335 135.025 ;
        RECT 18.345 134.215 23.855 135.025 ;
        RECT 24.235 134.345 33.515 135.025 ;
        RECT 24.235 134.225 26.570 134.345 ;
        RECT 24.235 134.115 25.155 134.225 ;
        RECT 31.235 134.125 32.155 134.345 ;
        RECT 33.525 134.215 34.895 135.025 ;
        RECT 34.915 134.115 36.265 135.025 ;
        RECT 37.215 134.155 37.645 134.940 ;
        RECT 37.665 134.215 40.415 135.025 ;
        RECT 40.585 134.205 42.515 135.025 ;
        RECT 42.885 134.205 44.815 135.025 ;
        RECT 41.565 134.115 42.515 134.205 ;
        RECT 43.865 134.115 44.815 134.205 ;
        RECT 45.225 134.205 47.155 135.025 ;
        RECT 47.470 134.995 47.640 135.045 ;
        RECT 51.605 135.025 51.775 135.215 ;
        RECT 56.205 135.045 56.375 135.235 ;
        RECT 57.125 135.025 57.295 135.215 ;
        RECT 57.590 135.025 57.760 135.215 ;
        RECT 61.725 135.045 61.895 135.235 ;
        RECT 62.645 135.025 62.815 135.215 ;
        RECT 64.025 135.070 64.185 135.180 ;
        RECT 65.590 135.045 65.760 135.235 ;
        RECT 67.705 135.025 67.875 135.215 ;
        RECT 73.225 135.025 73.395 135.215 ;
        RECT 75.525 135.045 75.695 135.235 ;
        RECT 76.905 135.080 77.065 135.190 ;
        RECT 78.745 135.025 78.915 135.215 ;
        RECT 80.585 135.045 80.755 135.235 ;
        RECT 81.050 135.045 81.220 135.265 ;
        RECT 82.710 135.235 83.655 135.265 ;
        RECT 84.585 135.235 88.255 136.045 ;
        RECT 91.465 135.915 92.395 136.145 ;
        RECT 88.495 135.235 92.395 135.915 ;
        RECT 92.415 135.235 93.765 136.145 ;
        RECT 93.785 135.235 97.455 136.045 ;
        RECT 100.665 135.915 101.595 136.145 ;
        RECT 97.695 135.235 101.595 135.915 ;
        RECT 101.615 135.320 102.045 136.105 ;
        RECT 102.065 135.235 103.895 136.045 ;
        RECT 103.905 135.235 105.275 136.015 ;
        RECT 105.285 135.235 106.655 136.045 ;
        RECT 106.675 135.235 108.025 136.145 ;
        RECT 108.045 135.235 109.875 136.045 ;
        RECT 109.885 135.235 111.255 136.015 ;
        RECT 111.725 135.235 115.395 136.045 ;
        RECT 115.405 135.235 120.915 136.045 ;
        RECT 120.925 135.235 126.435 136.045 ;
        RECT 126.445 135.235 127.815 136.045 ;
        RECT 82.420 135.025 82.590 135.215 ;
        RECT 82.890 135.025 83.060 135.215 ;
        RECT 84.265 135.080 84.425 135.190 ;
        RECT 86.620 135.075 86.740 135.185 ;
        RECT 87.945 135.045 88.115 135.235 ;
        RECT 88.405 135.025 88.575 135.215 ;
        RECT 91.810 135.045 91.980 135.235 ;
        RECT 92.730 135.025 92.900 135.215 ;
        RECT 93.465 135.025 93.635 135.235 ;
        RECT 94.900 135.075 95.020 135.185 ;
        RECT 96.685 135.025 96.855 135.215 ;
        RECT 97.145 135.045 97.315 135.235 ;
        RECT 101.010 135.045 101.180 135.235 ;
        RECT 103.585 135.045 103.755 135.235 ;
        RECT 104.045 135.045 104.215 135.235 ;
        RECT 106.345 135.025 106.515 135.235 ;
        RECT 106.805 135.045 106.975 135.235 ;
        RECT 109.105 135.025 109.275 135.215 ;
        RECT 109.565 135.045 109.735 135.235 ;
        RECT 110.025 135.045 110.195 135.235 ;
        RECT 111.405 135.185 111.575 135.215 ;
        RECT 111.405 135.075 111.580 135.185 ;
        RECT 111.405 135.045 111.575 135.075 ;
        RECT 113.705 135.045 113.875 135.215 ;
        RECT 115.085 135.185 115.255 135.235 ;
        RECT 114.220 135.075 114.340 135.185 ;
        RECT 115.085 135.075 115.260 135.185 ;
        RECT 115.085 135.045 115.255 135.075 ;
        RECT 111.405 135.025 111.555 135.045 ;
        RECT 113.705 135.025 113.855 135.045 ;
        RECT 120.605 135.025 120.775 135.235 ;
        RECT 126.125 135.025 126.295 135.235 ;
        RECT 127.505 135.025 127.675 135.235 ;
        RECT 49.130 134.995 50.075 135.025 ;
        RECT 47.325 134.315 50.075 134.995 ;
        RECT 45.225 134.115 46.175 134.205 ;
        RECT 49.130 134.115 50.075 134.315 ;
        RECT 50.085 134.215 51.915 135.025 ;
        RECT 51.925 134.215 57.435 135.025 ;
        RECT 57.445 134.115 60.920 135.025 ;
        RECT 61.125 134.215 62.955 135.025 ;
        RECT 62.975 134.155 63.405 134.940 ;
        RECT 64.345 134.215 68.015 135.025 ;
        RECT 68.025 134.215 73.535 135.025 ;
        RECT 73.545 134.215 79.055 135.025 ;
        RECT 79.260 134.115 82.735 135.025 ;
        RECT 82.745 134.115 86.220 135.025 ;
        RECT 86.885 134.215 88.715 135.025 ;
        RECT 88.735 134.155 89.165 134.940 ;
        RECT 89.415 134.345 93.315 135.025 ;
        RECT 92.385 134.115 93.315 134.345 ;
        RECT 93.325 134.245 94.695 135.025 ;
        RECT 95.165 134.215 96.995 135.025 ;
        RECT 97.375 134.345 106.655 135.025 ;
        RECT 97.375 134.225 99.710 134.345 ;
        RECT 97.375 134.115 98.295 134.225 ;
        RECT 104.375 134.125 105.295 134.345 ;
        RECT 106.665 134.215 109.415 135.025 ;
        RECT 109.625 134.205 111.555 135.025 ;
        RECT 111.925 134.205 113.855 135.025 ;
        RECT 109.625 134.115 110.575 134.205 ;
        RECT 111.925 134.115 112.875 134.205 ;
        RECT 114.495 134.155 114.925 134.940 ;
        RECT 115.405 134.215 120.915 135.025 ;
        RECT 120.925 134.215 126.435 135.025 ;
        RECT 126.445 134.215 127.815 135.025 ;
      LAYER nwell ;
        RECT 14.470 130.995 128.010 133.825 ;
      LAYER pwell ;
        RECT 14.665 129.795 16.035 130.605 ;
        RECT 16.045 129.795 18.795 130.605 ;
        RECT 18.815 129.795 20.165 130.705 ;
        RECT 23.385 130.475 24.315 130.705 ;
        RECT 20.415 129.795 24.315 130.475 ;
        RECT 24.335 129.880 24.765 130.665 ;
        RECT 24.785 129.795 26.155 130.575 ;
        RECT 26.175 129.795 27.525 130.705 ;
        RECT 30.745 130.475 31.675 130.705 ;
        RECT 27.775 129.795 31.675 130.475 ;
        RECT 32.055 130.595 32.975 130.705 ;
        RECT 32.055 130.475 34.390 130.595 ;
        RECT 39.055 130.475 39.975 130.695 ;
        RECT 42.265 130.475 43.195 130.705 ;
        RECT 46.865 130.505 47.810 130.705 ;
        RECT 32.055 129.795 41.335 130.475 ;
        RECT 42.265 129.795 46.165 130.475 ;
        RECT 46.865 129.825 49.615 130.505 ;
        RECT 50.095 129.880 50.525 130.665 ;
        RECT 50.745 130.615 51.695 130.705 ;
        RECT 46.865 129.795 47.810 129.825 ;
        RECT 14.805 129.585 14.975 129.795 ;
        RECT 16.240 129.635 16.360 129.745 ;
        RECT 18.485 129.605 18.655 129.795 ;
        RECT 19.865 129.605 20.035 129.795 ;
        RECT 23.730 129.605 23.900 129.795 ;
        RECT 25.845 129.585 26.015 129.795 ;
        RECT 26.305 129.745 26.475 129.795 ;
        RECT 26.305 129.635 26.480 129.745 ;
        RECT 26.305 129.605 26.475 129.635 ;
        RECT 31.090 129.605 31.260 129.795 ;
        RECT 31.825 129.585 31.995 129.775 ;
        RECT 33.205 129.585 33.375 129.775 ;
        RECT 36.885 129.585 37.055 129.775 ;
        RECT 41.025 129.585 41.195 129.795 ;
        RECT 41.945 129.640 42.105 129.750 ;
        RECT 42.405 129.585 42.575 129.775 ;
        RECT 42.680 129.605 42.850 129.795 ;
        RECT 49.300 129.775 49.470 129.825 ;
        RECT 50.745 129.795 52.675 130.615 ;
        RECT 53.765 129.795 57.240 130.705 ;
        RECT 57.445 129.795 60.920 130.705 ;
        RECT 61.585 129.795 65.255 130.605 ;
        RECT 68.465 130.475 69.395 130.705 ;
        RECT 65.495 129.795 69.395 130.475 ;
        RECT 69.405 129.795 70.775 130.575 ;
        RECT 70.785 129.795 72.615 130.475 ;
        RECT 72.625 129.795 74.455 130.475 ;
        RECT 74.465 129.795 75.835 130.605 ;
        RECT 75.855 129.880 76.285 130.665 ;
        RECT 76.305 129.795 79.975 130.605 ;
        RECT 79.985 130.505 80.930 130.705 ;
        RECT 79.985 129.825 82.735 130.505 ;
        RECT 79.985 129.795 80.930 129.825 ;
        RECT 52.525 129.775 52.675 129.795 ;
        RECT 42.865 129.605 43.035 129.775 ;
        RECT 46.600 129.635 46.720 129.745 ;
        RECT 42.885 129.585 43.035 129.605 ;
        RECT 14.665 128.775 16.035 129.585 ;
        RECT 16.875 128.905 26.155 129.585 ;
        RECT 16.875 128.785 19.210 128.905 ;
        RECT 16.875 128.675 17.795 128.785 ;
        RECT 23.875 128.685 24.795 128.905 ;
        RECT 26.625 128.775 32.135 129.585 ;
        RECT 32.145 128.805 33.515 129.585 ;
        RECT 33.525 128.775 37.195 129.585 ;
        RECT 37.215 128.715 37.645 129.500 ;
        RECT 37.665 128.775 41.335 129.585 ;
        RECT 41.345 128.805 42.715 129.585 ;
        RECT 42.885 128.765 44.815 129.585 ;
        RECT 43.865 128.675 44.815 128.765 ;
        RECT 45.025 129.555 45.970 129.585 ;
        RECT 47.460 129.555 47.630 129.775 ;
        RECT 49.300 129.605 49.475 129.775 ;
        RECT 49.820 129.635 49.940 129.745 ;
        RECT 49.305 129.585 49.475 129.605 ;
        RECT 45.025 128.875 47.775 129.555 ;
        RECT 45.025 128.675 45.970 128.875 ;
        RECT 47.785 128.775 49.615 129.585 ;
        RECT 49.625 129.555 50.570 129.585 ;
        RECT 52.060 129.555 52.230 129.775 ;
        RECT 52.525 129.605 52.695 129.775 ;
        RECT 53.445 129.585 53.615 129.775 ;
        RECT 53.910 129.605 54.080 129.795 ;
        RECT 56.205 129.585 56.375 129.775 ;
        RECT 56.720 129.635 56.840 129.745 ;
        RECT 57.130 129.585 57.300 129.775 ;
        RECT 57.590 129.605 57.760 129.795 ;
        RECT 61.320 129.740 61.440 129.745 ;
        RECT 61.265 129.635 61.440 129.740 ;
        RECT 61.265 129.630 61.425 129.635 ;
        RECT 61.725 129.585 61.895 129.775 ;
        RECT 63.565 129.585 63.735 129.775 ;
        RECT 64.945 129.605 65.115 129.795 ;
        RECT 68.810 129.605 68.980 129.795 ;
        RECT 69.545 129.605 69.715 129.795 ;
        RECT 72.305 129.605 72.475 129.795 ;
        RECT 74.145 129.585 74.315 129.795 ;
        RECT 75.525 129.605 75.695 129.795 ;
        RECT 76.445 129.605 76.615 129.775 ;
        RECT 79.665 129.605 79.835 129.795 ;
        RECT 76.445 129.585 76.595 129.605 ;
        RECT 81.965 129.585 82.135 129.775 ;
        RECT 82.420 129.605 82.590 129.825 ;
        RECT 82.745 129.795 84.115 130.605 ;
        RECT 84.125 129.795 87.795 130.605 ;
        RECT 88.175 130.595 89.095 130.705 ;
        RECT 88.175 130.475 90.510 130.595 ;
        RECT 95.175 130.475 96.095 130.695 ;
        RECT 88.175 129.795 97.455 130.475 ;
        RECT 97.465 129.795 100.215 130.605 ;
        RECT 100.235 129.795 101.585 130.705 ;
        RECT 101.615 129.880 102.045 130.665 ;
        RECT 104.105 130.615 105.055 130.705 ;
        RECT 106.405 130.615 107.355 130.705 ;
        RECT 102.065 129.795 103.895 130.605 ;
        RECT 104.105 129.795 106.035 130.615 ;
        RECT 106.405 129.795 108.335 130.615 ;
        RECT 111.705 130.475 112.635 130.705 ;
        RECT 108.735 129.795 112.635 130.475 ;
        RECT 112.845 130.615 113.795 130.705 ;
        RECT 112.845 129.795 114.775 130.615 ;
        RECT 118.605 130.475 119.535 130.705 ;
        RECT 115.635 129.795 119.535 130.475 ;
        RECT 119.545 129.795 120.915 130.605 ;
        RECT 120.925 129.795 126.435 130.605 ;
        RECT 126.445 129.795 127.815 130.605 ;
        RECT 83.805 129.605 83.975 129.795 ;
        RECT 84.265 129.605 84.435 129.775 ;
        RECT 84.780 129.635 84.900 129.745 ;
        RECT 87.485 129.605 87.655 129.795 ;
        RECT 84.265 129.585 84.415 129.605 ;
        RECT 88.405 129.585 88.575 129.775 ;
        RECT 89.380 129.635 89.500 129.745 ;
        RECT 92.085 129.585 92.255 129.775 ;
        RECT 93.465 129.585 93.635 129.775 ;
        RECT 97.145 129.605 97.315 129.795 ;
        RECT 98.985 129.585 99.155 129.775 ;
        RECT 99.905 129.605 100.075 129.795 ;
        RECT 100.365 129.605 100.535 129.795 ;
        RECT 101.285 129.605 101.455 129.775 ;
        RECT 101.285 129.585 101.435 129.605 ;
        RECT 103.125 129.585 103.295 129.775 ;
        RECT 103.585 129.585 103.755 129.795 ;
        RECT 105.885 129.775 106.035 129.795 ;
        RECT 108.185 129.775 108.335 129.795 ;
        RECT 105.885 129.605 106.055 129.775 ;
        RECT 108.185 129.605 108.355 129.775 ;
        RECT 112.050 129.605 112.220 129.795 ;
        RECT 114.625 129.775 114.775 129.795 ;
        RECT 112.840 129.635 112.960 129.745 ;
        RECT 113.245 129.585 113.415 129.775 ;
        RECT 114.625 129.605 114.795 129.775 ;
        RECT 115.085 129.745 115.255 129.775 ;
        RECT 115.085 129.635 115.260 129.745 ;
        RECT 115.085 129.585 115.255 129.635 ;
        RECT 118.950 129.605 119.120 129.795 ;
        RECT 120.605 129.605 120.775 129.795 ;
        RECT 125.665 129.585 125.835 129.775 ;
        RECT 126.125 129.745 126.295 129.795 ;
        RECT 126.125 129.635 126.300 129.745 ;
        RECT 126.125 129.605 126.295 129.635 ;
        RECT 127.505 129.585 127.675 129.795 ;
        RECT 49.625 128.875 52.375 129.555 ;
        RECT 49.625 128.675 50.570 128.875 ;
        RECT 52.385 128.775 53.755 129.585 ;
        RECT 53.775 128.905 56.515 129.585 ;
        RECT 56.985 128.675 60.460 129.585 ;
        RECT 61.595 128.675 62.945 129.585 ;
        RECT 62.975 128.715 63.405 129.500 ;
        RECT 63.435 128.675 64.785 129.585 ;
        RECT 65.175 128.905 74.455 129.585 ;
        RECT 65.175 128.785 67.510 128.905 ;
        RECT 65.175 128.675 66.095 128.785 ;
        RECT 72.175 128.685 73.095 128.905 ;
        RECT 74.665 128.765 76.595 129.585 ;
        RECT 76.765 128.775 82.275 129.585 ;
        RECT 82.485 128.765 84.415 129.585 ;
        RECT 85.045 128.775 88.715 129.585 ;
        RECT 74.665 128.675 75.615 128.765 ;
        RECT 82.485 128.675 83.435 128.765 ;
        RECT 88.735 128.715 89.165 129.500 ;
        RECT 89.645 128.775 92.395 129.585 ;
        RECT 92.415 128.675 93.765 129.585 ;
        RECT 93.785 128.775 99.295 129.585 ;
        RECT 99.505 128.765 101.435 129.585 ;
        RECT 101.605 128.775 103.435 129.585 ;
        RECT 103.445 128.905 112.550 129.585 ;
        RECT 99.505 128.675 100.455 128.765 ;
        RECT 113.115 128.675 114.465 129.585 ;
        RECT 114.495 128.715 114.925 129.500 ;
        RECT 114.955 128.675 116.305 129.585 ;
        RECT 116.695 128.905 125.975 129.585 ;
        RECT 116.695 128.785 119.030 128.905 ;
        RECT 116.695 128.675 117.615 128.785 ;
        RECT 123.695 128.685 124.615 128.905 ;
        RECT 126.445 128.775 127.815 129.585 ;
      LAYER nwell ;
        RECT 14.470 125.555 128.010 128.385 ;
      LAYER pwell ;
        RECT 14.665 124.355 16.035 125.165 ;
        RECT 16.045 124.355 18.795 125.165 ;
        RECT 18.805 124.355 20.175 125.135 ;
        RECT 20.185 125.035 21.115 125.265 ;
        RECT 20.185 124.355 24.085 125.035 ;
        RECT 24.335 124.440 24.765 125.225 ;
        RECT 25.705 125.035 26.635 125.265 ;
        RECT 25.705 124.355 29.605 125.035 ;
        RECT 30.305 124.355 33.055 125.165 ;
        RECT 36.265 125.035 37.195 125.265 ;
        RECT 40.645 125.175 41.595 125.265 ;
        RECT 42.945 125.175 43.895 125.265 ;
        RECT 45.245 125.175 46.195 125.265 ;
        RECT 48.925 125.175 49.875 125.265 ;
        RECT 33.295 124.355 37.195 125.035 ;
        RECT 37.665 124.355 39.495 125.165 ;
        RECT 39.665 124.355 41.595 125.175 ;
        RECT 41.965 124.355 43.895 125.175 ;
        RECT 44.265 124.355 46.195 125.175 ;
        RECT 46.405 124.355 47.775 125.165 ;
        RECT 47.945 124.355 49.875 125.175 ;
        RECT 50.095 124.440 50.525 125.225 ;
        RECT 50.545 124.355 51.915 125.165 ;
        RECT 51.925 124.355 55.595 125.165 ;
        RECT 55.605 124.355 61.115 125.165 ;
        RECT 61.495 125.155 62.415 125.265 ;
        RECT 61.495 125.035 63.830 125.155 ;
        RECT 68.495 125.035 69.415 125.255 ;
        RECT 61.495 124.355 70.775 125.035 ;
        RECT 70.785 124.355 72.155 125.135 ;
        RECT 73.085 124.355 75.825 125.035 ;
        RECT 75.855 124.440 76.285 125.225 ;
        RECT 78.345 125.175 79.295 125.265 ;
        RECT 81.585 125.175 82.535 125.265 ;
        RECT 76.305 124.355 78.135 125.165 ;
        RECT 78.345 124.355 80.275 125.175 ;
        RECT 14.805 124.145 14.975 124.355 ;
        RECT 18.485 124.165 18.655 124.355 ;
        RECT 18.945 124.165 19.115 124.355 ;
        RECT 20.600 124.165 20.770 124.355 ;
        RECT 25.385 124.145 25.555 124.335 ;
        RECT 25.900 124.195 26.020 124.305 ;
        RECT 26.120 124.165 26.290 124.355 ;
        RECT 27.685 124.145 27.855 124.335 ;
        RECT 30.040 124.195 30.160 124.305 ;
        RECT 32.745 124.165 32.915 124.355 ;
        RECT 36.610 124.165 36.780 124.355 ;
        RECT 36.885 124.145 37.055 124.335 ;
        RECT 37.400 124.195 37.520 124.305 ;
        RECT 37.860 124.195 37.980 124.305 ;
        RECT 39.185 124.165 39.355 124.355 ;
        RECT 39.665 124.335 39.815 124.355 ;
        RECT 41.965 124.335 42.115 124.355 ;
        RECT 44.265 124.335 44.415 124.355 ;
        RECT 39.645 124.145 39.815 124.335 ;
        RECT 41.945 124.165 42.115 124.335 ;
        RECT 44.245 124.165 44.415 124.335 ;
        RECT 45.165 124.145 45.335 124.335 ;
        RECT 47.465 124.165 47.635 124.355 ;
        RECT 47.945 124.335 48.095 124.355 ;
        RECT 47.925 124.165 48.095 124.335 ;
        RECT 50.685 124.145 50.855 124.335 ;
        RECT 51.605 124.165 51.775 124.355 ;
        RECT 54.550 124.145 54.720 124.335 ;
        RECT 55.285 124.165 55.455 124.355 ;
        RECT 55.745 124.190 55.905 124.300 ;
        RECT 58.500 124.145 58.670 124.335 ;
        RECT 59.020 124.195 59.140 124.305 ;
        RECT 60.805 124.165 60.975 124.355 ;
        RECT 61.725 124.145 61.895 124.335 ;
        RECT 62.645 124.190 62.805 124.300 ;
        RECT 66.970 124.145 67.140 124.335 ;
        RECT 68.625 124.145 68.795 124.335 ;
        RECT 70.465 124.165 70.635 124.355 ;
        RECT 71.845 124.165 72.015 124.355 ;
        RECT 72.305 124.145 72.475 124.335 ;
        RECT 72.765 124.200 72.925 124.310 ;
        RECT 73.225 124.165 73.395 124.355 ;
        RECT 77.825 124.145 77.995 124.355 ;
        RECT 80.125 124.335 80.275 124.355 ;
        RECT 80.605 124.355 82.535 125.175 ;
        RECT 82.945 125.175 83.895 125.265 ;
        RECT 82.945 124.355 84.875 125.175 ;
        RECT 85.505 124.355 91.015 125.165 ;
        RECT 91.025 124.355 96.535 125.165 ;
        RECT 96.545 124.355 97.915 125.135 ;
        RECT 97.925 124.355 101.595 125.165 ;
        RECT 101.615 124.440 102.045 125.225 ;
        RECT 102.535 124.355 103.885 125.265 ;
        RECT 104.275 125.155 105.195 125.265 ;
        RECT 104.275 125.035 106.610 125.155 ;
        RECT 111.275 125.035 112.195 125.255 ;
        RECT 115.775 125.155 116.695 125.265 ;
        RECT 104.275 124.355 113.555 125.035 ;
        RECT 113.565 124.355 114.935 125.135 ;
        RECT 115.775 125.035 118.110 125.155 ;
        RECT 122.775 125.035 123.695 125.255 ;
        RECT 115.775 124.355 125.055 125.035 ;
        RECT 125.065 124.355 126.435 125.135 ;
        RECT 126.445 124.355 127.815 125.165 ;
        RECT 80.605 124.335 80.755 124.355 ;
        RECT 84.725 124.335 84.875 124.355 ;
        RECT 80.125 124.165 80.295 124.335 ;
        RECT 80.585 124.165 80.755 124.335 ;
        RECT 81.690 124.145 81.860 124.335 ;
        RECT 84.725 124.165 84.895 124.335 ;
        RECT 85.240 124.195 85.360 124.305 ;
        RECT 85.830 124.145 86.000 124.335 ;
        RECT 86.620 124.195 86.740 124.305 ;
        RECT 88.405 124.145 88.575 124.335 ;
        RECT 90.245 124.145 90.415 124.335 ;
        RECT 90.705 124.145 90.875 124.355 ;
        RECT 95.490 124.145 95.660 124.335 ;
        RECT 96.225 124.165 96.395 124.355 ;
        RECT 96.685 124.165 96.855 124.355 ;
        RECT 101.285 124.165 101.455 124.355 ;
        RECT 102.260 124.195 102.380 124.305 ;
        RECT 102.665 124.165 102.835 124.355 ;
        RECT 105.425 124.145 105.595 124.335 ;
        RECT 106.160 124.145 106.330 124.335 ;
        RECT 110.485 124.190 110.645 124.300 ;
        RECT 112.325 124.165 112.495 124.335 ;
        RECT 113.245 124.165 113.415 124.355 ;
        RECT 114.165 124.145 114.335 124.335 ;
        RECT 114.625 124.165 114.795 124.355 ;
        RECT 115.140 124.195 115.260 124.305 ;
        RECT 118.950 124.145 119.120 124.335 ;
        RECT 120.605 124.145 120.775 124.335 ;
        RECT 121.065 124.145 121.235 124.335 ;
        RECT 122.500 124.195 122.620 124.305 ;
        RECT 124.745 124.165 124.915 124.355 ;
        RECT 126.125 124.145 126.295 124.355 ;
        RECT 127.505 124.145 127.675 124.355 ;
        RECT 14.665 123.335 16.035 124.145 ;
        RECT 16.415 123.465 25.695 124.145 ;
        RECT 16.415 123.345 18.750 123.465 ;
        RECT 16.415 123.235 17.335 123.345 ;
        RECT 23.415 123.245 24.335 123.465 ;
        RECT 26.165 123.335 27.995 124.145 ;
        RECT 28.090 123.465 37.195 124.145 ;
        RECT 37.215 123.275 37.645 124.060 ;
        RECT 38.125 123.335 39.955 124.145 ;
        RECT 39.965 123.335 45.475 124.145 ;
        RECT 45.485 123.335 50.995 124.145 ;
        RECT 51.235 123.465 55.135 124.145 ;
        RECT 54.205 123.235 55.135 123.465 ;
        RECT 56.205 123.235 58.815 124.145 ;
        RECT 59.945 123.335 62.035 124.145 ;
        RECT 62.975 123.275 63.405 124.060 ;
        RECT 63.655 123.465 67.555 124.145 ;
        RECT 66.625 123.235 67.555 123.465 ;
        RECT 67.565 123.335 68.935 124.145 ;
        RECT 68.945 123.335 72.615 124.145 ;
        RECT 72.625 123.335 78.135 124.145 ;
        RECT 78.375 123.465 82.275 124.145 ;
        RECT 82.515 123.465 86.415 124.145 ;
        RECT 81.345 123.235 82.275 123.465 ;
        RECT 85.485 123.235 86.415 123.465 ;
        RECT 86.885 123.335 88.715 124.145 ;
        RECT 88.735 123.275 89.165 124.060 ;
        RECT 89.185 123.335 90.555 124.145 ;
        RECT 90.575 123.235 91.925 124.145 ;
        RECT 92.175 123.465 96.075 124.145 ;
        RECT 95.145 123.235 96.075 123.465 ;
        RECT 96.455 123.465 105.735 124.145 ;
        RECT 105.745 123.465 109.645 124.145 ;
        RECT 110.805 123.465 112.170 124.145 ;
        RECT 96.455 123.345 98.790 123.465 ;
        RECT 96.455 123.235 97.375 123.345 ;
        RECT 103.455 123.245 104.375 123.465 ;
        RECT 105.745 123.235 106.675 123.465 ;
        RECT 112.645 123.335 114.475 124.145 ;
        RECT 114.495 123.275 114.925 124.060 ;
        RECT 115.635 123.465 119.535 124.145 ;
        RECT 118.605 123.235 119.535 123.465 ;
        RECT 119.545 123.335 120.915 124.145 ;
        RECT 120.925 123.365 122.295 124.145 ;
        RECT 122.765 123.335 126.435 124.145 ;
        RECT 126.445 123.335 127.815 124.145 ;
      LAYER nwell ;
        RECT 14.470 120.115 128.010 122.945 ;
      LAYER pwell ;
        RECT 14.665 118.915 16.035 119.725 ;
        RECT 16.505 118.915 19.255 119.725 ;
        RECT 19.275 118.915 20.625 119.825 ;
        RECT 21.105 118.915 22.935 119.725 ;
        RECT 22.945 118.915 24.315 119.695 ;
        RECT 24.335 119.000 24.765 119.785 ;
        RECT 26.145 119.595 27.065 119.815 ;
        RECT 33.145 119.715 34.065 119.825 ;
        RECT 31.730 119.595 34.065 119.715 ;
        RECT 24.785 118.915 34.065 119.595 ;
        RECT 34.455 118.915 35.805 119.825 ;
        RECT 36.195 119.715 37.115 119.825 ;
        RECT 36.195 119.595 38.530 119.715 ;
        RECT 43.195 119.595 44.115 119.815 ;
        RECT 49.145 119.595 50.075 119.825 ;
        RECT 36.195 118.915 45.475 119.595 ;
        RECT 46.175 118.915 50.075 119.595 ;
        RECT 50.095 119.000 50.525 119.785 ;
        RECT 51.005 118.915 52.835 119.725 ;
        RECT 52.845 118.915 61.950 119.595 ;
        RECT 62.045 118.915 63.415 119.725 ;
        RECT 66.625 119.595 67.555 119.825 ;
        RECT 63.655 118.915 67.555 119.595 ;
        RECT 68.025 118.915 69.395 119.695 ;
        RECT 70.325 118.915 75.835 119.725 ;
        RECT 75.855 119.000 76.285 119.785 ;
        RECT 76.775 118.915 78.125 119.825 ;
        RECT 78.515 119.715 79.435 119.825 ;
        RECT 78.515 119.595 80.850 119.715 ;
        RECT 85.515 119.595 86.435 119.815 ;
        RECT 90.015 119.715 90.935 119.825 ;
        RECT 78.515 118.915 87.795 119.595 ;
        RECT 87.805 118.915 89.175 119.695 ;
        RECT 90.015 119.595 92.350 119.715 ;
        RECT 97.015 119.595 97.935 119.815 ;
        RECT 90.015 118.915 99.295 119.595 ;
        RECT 99.305 118.915 100.260 119.595 ;
        RECT 101.615 119.000 102.045 119.785 ;
        RECT 102.065 118.915 103.895 119.725 ;
        RECT 103.905 118.915 105.275 119.695 ;
        RECT 105.285 118.915 107.115 119.725 ;
        RECT 107.125 118.915 112.635 119.725 ;
        RECT 112.645 118.915 118.155 119.725 ;
        RECT 118.175 118.915 119.525 119.825 ;
        RECT 119.545 118.915 120.915 119.695 ;
        RECT 120.925 118.915 126.435 119.725 ;
        RECT 126.445 118.915 127.815 119.725 ;
        RECT 14.805 118.705 14.975 118.915 ;
        RECT 16.240 118.755 16.360 118.865 ;
        RECT 17.565 118.705 17.735 118.895 ;
        RECT 18.945 118.725 19.115 118.915 ;
        RECT 20.325 118.725 20.495 118.915 ;
        RECT 20.840 118.755 20.960 118.865 ;
        RECT 21.430 118.705 21.600 118.895 ;
        RECT 22.165 118.705 22.335 118.895 ;
        RECT 22.625 118.725 22.795 118.915 ;
        RECT 23.085 118.725 23.255 118.915 ;
        RECT 24.925 118.725 25.095 118.915 ;
        RECT 31.825 118.705 31.995 118.895 ;
        RECT 34.585 118.725 34.755 118.915 ;
        RECT 36.610 118.705 36.780 118.895 ;
        RECT 37.805 118.705 37.975 118.895 ;
        RECT 39.185 118.705 39.355 118.895 ;
        RECT 45.165 118.725 45.335 118.915 ;
        RECT 45.680 118.755 45.800 118.865 ;
        RECT 49.490 118.725 49.660 118.915 ;
        RECT 49.765 118.705 49.935 118.895 ;
        RECT 50.740 118.755 50.860 118.865 ;
        RECT 52.525 118.725 52.695 118.915 ;
        RECT 52.985 118.725 53.155 118.915 ;
        RECT 59.425 118.705 59.595 118.895 ;
        RECT 59.940 118.755 60.060 118.865 ;
        RECT 62.645 118.705 62.815 118.895 ;
        RECT 63.105 118.725 63.275 118.915 ;
        RECT 64.025 118.750 64.185 118.860 ;
        RECT 66.970 118.725 67.140 118.915 ;
        RECT 67.760 118.755 67.880 118.865 ;
        RECT 68.165 118.725 68.335 118.915 ;
        RECT 70.005 118.760 70.165 118.870 ;
        RECT 73.685 118.705 73.855 118.895 ;
        RECT 74.200 118.755 74.320 118.865 ;
        RECT 75.525 118.725 75.695 118.915 ;
        RECT 75.985 118.705 76.155 118.895 ;
        RECT 76.500 118.755 76.620 118.865 ;
        RECT 76.905 118.725 77.075 118.915 ;
        RECT 85.645 118.705 85.815 118.895 ;
        RECT 87.025 118.705 87.195 118.895 ;
        RECT 87.485 118.705 87.655 118.915 ;
        RECT 88.865 118.725 89.035 118.915 ;
        RECT 89.325 118.865 89.495 118.895 ;
        RECT 89.325 118.755 89.500 118.865 ;
        RECT 89.325 118.705 89.495 118.755 ;
        RECT 98.525 118.705 98.695 118.895 ;
        RECT 98.985 118.725 99.155 118.915 ;
        RECT 100.365 118.725 100.535 118.895 ;
        RECT 101.285 118.760 101.445 118.870 ;
        RECT 103.125 118.705 103.295 118.895 ;
        RECT 103.585 118.705 103.755 118.915 ;
        RECT 104.965 118.725 105.135 118.915 ;
        RECT 106.805 118.725 106.975 118.915 ;
        RECT 108.370 118.705 108.540 118.895 ;
        RECT 110.025 118.705 110.195 118.895 ;
        RECT 112.325 118.725 112.495 118.915 ;
        RECT 113.890 118.705 114.060 118.895 ;
        RECT 117.845 118.725 118.015 118.915 ;
        RECT 118.305 118.725 118.475 118.915 ;
        RECT 119.685 118.725 119.855 118.915 ;
        RECT 124.285 118.705 124.455 118.895 ;
        RECT 126.125 118.705 126.295 118.915 ;
        RECT 127.505 118.705 127.675 118.915 ;
        RECT 14.665 117.895 16.035 118.705 ;
        RECT 16.045 117.895 17.875 118.705 ;
        RECT 18.115 118.025 22.015 118.705 ;
        RECT 22.025 118.025 31.305 118.705 ;
        RECT 21.085 117.795 22.015 118.025 ;
        RECT 23.385 117.805 24.305 118.025 ;
        RECT 28.970 117.905 31.305 118.025 ;
        RECT 30.385 117.795 31.305 117.905 ;
        RECT 31.695 117.795 33.045 118.705 ;
        RECT 33.295 118.025 37.195 118.705 ;
        RECT 36.265 117.795 37.195 118.025 ;
        RECT 37.215 117.835 37.645 118.620 ;
        RECT 37.665 117.925 39.035 118.705 ;
        RECT 39.045 117.925 40.415 118.705 ;
        RECT 40.795 118.025 50.075 118.705 ;
        RECT 50.455 118.025 59.735 118.705 ;
        RECT 40.795 117.905 43.130 118.025 ;
        RECT 40.795 117.795 41.715 117.905 ;
        RECT 47.795 117.805 48.715 118.025 ;
        RECT 50.455 117.905 52.790 118.025 ;
        RECT 50.455 117.795 51.375 117.905 ;
        RECT 57.455 117.805 58.375 118.025 ;
        RECT 60.205 117.895 62.955 118.705 ;
        RECT 62.975 117.835 63.405 118.620 ;
        RECT 64.715 118.025 73.995 118.705 ;
        RECT 64.715 117.905 67.050 118.025 ;
        RECT 64.715 117.795 65.635 117.905 ;
        RECT 71.715 117.805 72.635 118.025 ;
        RECT 74.465 117.895 76.295 118.705 ;
        RECT 76.675 118.025 85.955 118.705 ;
        RECT 76.675 117.905 79.010 118.025 ;
        RECT 76.675 117.795 77.595 117.905 ;
        RECT 83.675 117.805 84.595 118.025 ;
        RECT 85.965 117.895 87.335 118.705 ;
        RECT 87.355 117.795 88.705 118.705 ;
        RECT 88.735 117.835 89.165 118.620 ;
        RECT 89.185 118.025 98.290 118.705 ;
        RECT 98.395 117.795 99.745 118.705 ;
        RECT 99.765 117.895 103.435 118.705 ;
        RECT 103.455 117.795 104.805 118.705 ;
        RECT 105.055 118.025 108.955 118.705 ;
        RECT 108.025 117.795 108.955 118.025 ;
        RECT 108.965 117.895 110.335 118.705 ;
        RECT 110.575 118.025 114.475 118.705 ;
        RECT 113.545 117.795 114.475 118.025 ;
        RECT 114.495 117.835 114.925 118.620 ;
        RECT 115.315 118.025 124.595 118.705 ;
        RECT 115.315 117.905 117.650 118.025 ;
        RECT 115.315 117.795 116.235 117.905 ;
        RECT 122.315 117.805 123.235 118.025 ;
        RECT 124.605 117.895 126.435 118.705 ;
        RECT 126.445 117.895 127.815 118.705 ;
      LAYER nwell ;
        RECT 14.470 114.675 128.010 117.505 ;
      LAYER pwell ;
        RECT 14.665 113.475 16.035 114.285 ;
        RECT 16.965 113.475 22.475 114.285 ;
        RECT 22.495 113.475 23.845 114.385 ;
        RECT 24.335 113.560 24.765 114.345 ;
        RECT 24.795 113.475 26.145 114.385 ;
        RECT 26.625 113.475 27.995 114.255 ;
        RECT 28.465 113.475 32.135 114.285 ;
        RECT 32.515 114.275 33.435 114.385 ;
        RECT 32.515 114.155 34.850 114.275 ;
        RECT 39.515 114.155 40.435 114.375 ;
        RECT 32.515 113.475 41.795 114.155 ;
        RECT 41.805 113.475 44.555 114.285 ;
        RECT 44.565 113.475 50.075 114.285 ;
        RECT 50.095 113.560 50.525 114.345 ;
        RECT 51.015 113.475 52.365 114.385 ;
        RECT 52.395 113.475 53.745 114.385 ;
        RECT 53.765 113.475 55.135 114.255 ;
        RECT 55.605 113.475 56.975 114.255 ;
        RECT 57.445 113.475 61.115 114.285 ;
        RECT 61.135 113.475 62.485 114.385 ;
        RECT 62.875 114.275 63.795 114.385 ;
        RECT 62.875 114.155 65.210 114.275 ;
        RECT 69.875 114.155 70.795 114.375 ;
        RECT 62.875 113.475 72.155 114.155 ;
        RECT 72.175 113.475 73.525 114.385 ;
        RECT 74.005 113.475 75.835 114.285 ;
        RECT 75.855 113.560 76.285 114.345 ;
        RECT 76.765 113.475 79.515 114.285 ;
        RECT 79.535 113.475 80.885 114.385 ;
        RECT 80.905 113.475 82.735 114.285 ;
        RECT 82.745 113.475 84.115 114.255 ;
        RECT 84.125 113.475 87.795 114.285 ;
        RECT 88.175 114.275 89.095 114.385 ;
        RECT 88.175 114.155 90.510 114.275 ;
        RECT 95.175 114.155 96.095 114.375 ;
        RECT 88.175 113.475 97.455 114.155 ;
        RECT 97.925 113.475 101.595 114.285 ;
        RECT 101.615 113.560 102.045 114.345 ;
        RECT 102.525 113.475 104.355 114.285 ;
        RECT 104.735 114.275 105.655 114.385 ;
        RECT 104.735 114.155 107.070 114.275 ;
        RECT 111.735 114.155 112.655 114.375 ;
        RECT 104.735 113.475 114.015 114.155 ;
        RECT 114.025 113.475 115.395 114.285 ;
        RECT 115.405 113.475 120.915 114.285 ;
        RECT 120.925 113.475 126.435 114.285 ;
        RECT 126.445 113.475 127.815 114.285 ;
        RECT 14.805 113.265 14.975 113.475 ;
        RECT 16.240 113.315 16.360 113.425 ;
        RECT 16.645 113.320 16.805 113.430 ;
        RECT 18.025 113.265 18.195 113.455 ;
        RECT 22.165 113.285 22.335 113.475 ;
        RECT 22.625 113.285 22.795 113.475 ;
        RECT 24.060 113.315 24.180 113.425 ;
        RECT 24.925 113.285 25.095 113.475 ;
        RECT 26.360 113.315 26.480 113.425 ;
        RECT 27.685 113.285 27.855 113.475 ;
        RECT 28.200 113.315 28.320 113.425 ;
        RECT 28.605 113.265 28.775 113.455 ;
        RECT 29.985 113.265 30.155 113.455 ;
        RECT 31.825 113.285 31.995 113.475 ;
        RECT 33.665 113.265 33.835 113.455 ;
        RECT 35.045 113.265 35.215 113.455 ;
        RECT 35.560 113.315 35.680 113.425 ;
        RECT 36.885 113.265 37.055 113.455 ;
        RECT 41.485 113.285 41.655 113.475 ;
        RECT 42.865 113.265 43.035 113.455 ;
        RECT 44.245 113.265 44.415 113.475 ;
        RECT 45.165 113.310 45.325 113.420 ;
        RECT 45.625 113.265 45.795 113.455 ;
        RECT 47.925 113.265 48.095 113.455 ;
        RECT 49.765 113.285 49.935 113.475 ;
        RECT 50.740 113.315 50.860 113.425 ;
        RECT 51.605 113.265 51.775 113.455 ;
        RECT 52.065 113.285 52.235 113.475 ;
        RECT 52.525 113.285 52.695 113.475 ;
        RECT 54.825 113.285 54.995 113.475 ;
        RECT 55.340 113.315 55.460 113.425 ;
        RECT 55.745 113.285 55.915 113.475 ;
        RECT 57.125 113.425 57.295 113.455 ;
        RECT 57.125 113.315 57.300 113.425 ;
        RECT 57.125 113.265 57.295 113.315 ;
        RECT 60.805 113.285 60.975 113.475 ;
        RECT 61.265 113.285 61.435 113.475 ;
        RECT 62.645 113.265 62.815 113.455 ;
        RECT 64.485 113.265 64.655 113.455 ;
        RECT 68.350 113.265 68.520 113.455 ;
        RECT 69.140 113.315 69.260 113.425 ;
        RECT 69.545 113.265 69.715 113.455 ;
        RECT 70.980 113.315 71.100 113.425 ;
        RECT 71.845 113.285 72.015 113.475 ;
        RECT 73.225 113.285 73.395 113.475 ;
        RECT 73.685 113.425 73.855 113.455 ;
        RECT 73.685 113.315 73.860 113.425 ;
        RECT 73.685 113.265 73.855 113.315 ;
        RECT 75.525 113.285 75.695 113.475 ;
        RECT 76.500 113.315 76.620 113.425 ;
        RECT 79.205 113.265 79.375 113.475 ;
        RECT 79.665 113.285 79.835 113.475 ;
        RECT 80.585 113.265 80.755 113.455 ;
        RECT 81.100 113.315 81.220 113.425 ;
        RECT 82.425 113.285 82.595 113.475 ;
        RECT 82.885 113.265 83.055 113.475 ;
        RECT 87.485 113.285 87.655 113.475 ;
        RECT 88.405 113.265 88.575 113.455 ;
        RECT 92.730 113.265 92.900 113.455 ;
        RECT 93.465 113.265 93.635 113.455 ;
        RECT 97.145 113.285 97.315 113.475 ;
        RECT 97.660 113.315 97.780 113.425 ;
        RECT 98.065 113.265 98.235 113.455 ;
        RECT 101.285 113.285 101.455 113.475 ;
        RECT 102.260 113.315 102.380 113.425 ;
        RECT 103.585 113.265 103.755 113.455 ;
        RECT 104.045 113.285 104.215 113.475 ;
        RECT 109.105 113.265 109.275 113.455 ;
        RECT 109.565 113.265 109.735 113.455 ;
        RECT 113.705 113.285 113.875 113.475 ;
        RECT 114.165 113.265 114.335 113.455 ;
        RECT 115.085 113.425 115.255 113.475 ;
        RECT 115.085 113.315 115.260 113.425 ;
        RECT 115.085 113.285 115.255 113.315 ;
        RECT 118.765 113.265 118.935 113.455 ;
        RECT 119.225 113.265 119.395 113.455 ;
        RECT 120.605 113.265 120.775 113.475 ;
        RECT 122.905 113.265 123.075 113.455 ;
        RECT 123.420 113.315 123.540 113.425 ;
        RECT 126.125 113.265 126.295 113.475 ;
        RECT 127.505 113.265 127.675 113.475 ;
        RECT 14.665 112.455 16.035 113.265 ;
        RECT 16.505 112.455 18.335 113.265 ;
        RECT 18.545 112.585 28.915 113.265 ;
        RECT 18.545 112.355 20.755 112.585 ;
        RECT 23.475 112.365 24.405 112.585 ;
        RECT 28.925 112.455 30.295 113.265 ;
        RECT 30.305 112.455 33.975 113.265 ;
        RECT 33.995 112.355 35.345 113.265 ;
        RECT 35.825 112.485 37.195 113.265 ;
        RECT 37.215 112.395 37.645 113.180 ;
        RECT 37.665 112.455 43.175 113.265 ;
        RECT 43.185 112.485 44.555 113.265 ;
        RECT 45.485 112.485 46.855 113.265 ;
        RECT 46.865 112.455 48.235 113.265 ;
        RECT 48.245 112.455 51.915 113.265 ;
        RECT 51.925 112.455 57.435 113.265 ;
        RECT 57.445 112.455 62.955 113.265 ;
        RECT 62.975 112.395 63.405 113.180 ;
        RECT 63.425 112.455 64.795 113.265 ;
        RECT 65.035 112.585 68.935 113.265 ;
        RECT 68.005 112.355 68.935 112.585 ;
        RECT 69.405 112.485 70.775 113.265 ;
        RECT 71.245 112.455 73.995 113.265 ;
        RECT 74.005 112.455 79.515 113.265 ;
        RECT 79.535 112.355 80.885 113.265 ;
        RECT 81.365 112.455 83.195 113.265 ;
        RECT 83.205 112.455 88.715 113.265 ;
        RECT 88.735 112.395 89.165 113.180 ;
        RECT 89.415 112.585 93.315 113.265 ;
        RECT 92.385 112.355 93.315 112.585 ;
        RECT 93.325 112.485 94.695 113.265 ;
        RECT 94.705 112.455 98.375 113.265 ;
        RECT 98.385 112.455 103.895 113.265 ;
        RECT 103.905 112.455 109.415 113.265 ;
        RECT 109.425 112.485 110.795 113.265 ;
        RECT 110.805 112.455 114.475 113.265 ;
        RECT 114.495 112.395 114.925 113.180 ;
        RECT 115.405 112.455 119.075 113.265 ;
        RECT 119.095 112.355 120.445 113.265 ;
        RECT 120.465 112.485 121.835 113.265 ;
        RECT 121.845 112.485 123.215 113.265 ;
        RECT 123.685 112.455 126.435 113.265 ;
        RECT 126.445 112.455 127.815 113.265 ;
      LAYER nwell ;
        RECT 14.470 109.235 128.010 112.065 ;
      LAYER pwell ;
        RECT 14.665 108.035 16.035 108.845 ;
        RECT 16.045 108.035 17.415 108.845 ;
        RECT 17.425 108.035 22.935 108.845 ;
        RECT 22.945 108.035 24.315 108.815 ;
        RECT 24.335 108.120 24.765 108.905 ;
        RECT 24.985 108.715 27.195 108.945 ;
        RECT 29.915 108.715 30.845 108.935 ;
        RECT 36.485 108.715 38.695 108.945 ;
        RECT 41.415 108.715 42.345 108.935 ;
        RECT 24.985 108.035 35.355 108.715 ;
        RECT 36.485 108.035 46.855 108.715 ;
        RECT 46.865 108.035 48.235 108.815 ;
        RECT 48.245 108.035 50.075 108.845 ;
        RECT 50.095 108.120 50.525 108.905 ;
        RECT 51.465 108.035 55.135 108.845 ;
        RECT 55.145 108.035 56.515 108.815 ;
        RECT 56.525 108.035 60.195 108.845 ;
        RECT 60.205 108.035 62.815 108.945 ;
        RECT 63.425 108.035 64.795 108.815 ;
        RECT 65.265 108.035 68.015 108.845 ;
        RECT 68.025 108.035 69.395 108.815 ;
        RECT 69.405 108.035 70.775 108.845 ;
        RECT 70.785 108.035 74.455 108.845 ;
        RECT 74.475 108.035 75.825 108.945 ;
        RECT 75.855 108.120 76.285 108.905 ;
        RECT 76.775 108.035 78.125 108.945 ;
        RECT 78.145 108.035 80.755 108.945 ;
        RECT 80.905 108.035 82.275 108.815 ;
        RECT 82.285 108.035 83.655 108.815 ;
        RECT 84.585 108.035 88.255 108.845 ;
        RECT 88.275 108.035 89.625 108.945 ;
        RECT 89.645 108.035 91.015 108.815 ;
        RECT 91.225 108.715 93.435 108.945 ;
        RECT 96.155 108.715 97.085 108.935 ;
        RECT 91.225 108.035 101.595 108.715 ;
        RECT 101.615 108.120 102.045 108.905 ;
        RECT 102.065 108.035 103.435 108.815 ;
        RECT 104.375 108.035 105.725 108.945 ;
        RECT 106.665 108.035 108.035 108.815 ;
        RECT 108.045 108.035 109.415 108.845 ;
        RECT 109.425 108.035 110.795 108.815 ;
        RECT 110.805 108.035 114.475 108.845 ;
        RECT 114.485 108.035 115.855 108.815 ;
        RECT 120.375 108.715 121.305 108.935 ;
        RECT 124.025 108.715 126.235 108.945 ;
        RECT 115.865 108.035 126.235 108.715 ;
        RECT 126.445 108.035 127.815 108.845 ;
        RECT 14.805 107.825 14.975 108.035 ;
        RECT 16.240 107.875 16.360 107.985 ;
        RECT 17.105 107.845 17.275 108.035 ;
        RECT 19.865 107.825 20.035 108.015 ;
        RECT 21.245 107.825 21.415 108.015 ;
        RECT 22.165 107.870 22.325 107.980 ;
        RECT 22.625 107.845 22.795 108.035 ;
        RECT 23.085 107.845 23.255 108.035 ;
        RECT 23.545 107.825 23.715 108.015 ;
        RECT 34.125 107.825 34.295 108.015 ;
        RECT 34.585 107.825 34.755 108.015 ;
        RECT 35.045 107.845 35.215 108.035 ;
        RECT 35.965 107.825 36.135 108.015 ;
        RECT 37.860 107.875 37.980 107.985 ;
        RECT 46.545 107.845 46.715 108.035 ;
        RECT 47.925 107.845 48.095 108.035 ;
        RECT 48.385 107.825 48.555 108.015 ;
        RECT 49.765 107.825 49.935 108.035 ;
        RECT 51.145 107.825 51.315 108.015 ;
        RECT 54.825 107.845 54.995 108.035 ;
        RECT 55.285 107.845 55.455 108.035 ;
        RECT 59.885 107.845 60.055 108.035 ;
        RECT 60.350 107.845 60.520 108.035 ;
        RECT 61.725 107.825 61.895 108.015 ;
        RECT 62.645 107.870 62.805 107.980 ;
        RECT 63.160 107.875 63.280 107.985 ;
        RECT 63.565 107.845 63.735 108.035 ;
        RECT 65.000 107.875 65.120 107.985 ;
        RECT 67.705 107.845 67.875 108.035 ;
        RECT 68.165 107.845 68.335 108.035 ;
        RECT 70.465 107.845 70.635 108.035 ;
        RECT 73.685 107.825 73.855 108.015 ;
        RECT 74.145 107.845 74.315 108.035 ;
        RECT 74.605 107.870 74.765 107.980 ;
        RECT 75.525 107.845 75.695 108.035 ;
        RECT 76.500 107.875 76.620 107.985 ;
        RECT 77.825 107.845 77.995 108.035 ;
        RECT 78.290 107.845 78.460 108.035 ;
        RECT 81.045 107.845 81.215 108.035 ;
        RECT 82.425 107.845 82.595 108.035 ;
        RECT 84.265 107.880 84.425 107.990 ;
        RECT 85.185 107.825 85.355 108.015 ;
        RECT 85.645 107.825 85.815 108.015 ;
        RECT 87.025 107.825 87.195 108.015 ;
        RECT 87.945 107.845 88.115 108.035 ;
        RECT 88.405 107.985 88.575 108.035 ;
        RECT 88.405 107.875 88.580 107.985 ;
        RECT 88.405 107.845 88.575 107.875 ;
        RECT 89.325 107.825 89.495 108.015 ;
        RECT 89.785 107.845 89.955 108.035 ;
        RECT 99.960 107.875 100.080 107.985 ;
        RECT 101.285 107.845 101.455 108.035 ;
        RECT 103.125 107.845 103.295 108.035 ;
        RECT 104.045 107.880 104.205 107.990 ;
        RECT 105.425 107.845 105.595 108.035 ;
        RECT 106.345 107.880 106.505 107.990 ;
        RECT 106.805 107.845 106.975 108.035 ;
        RECT 109.105 107.845 109.275 108.035 ;
        RECT 110.485 107.825 110.655 108.035 ;
        RECT 111.865 107.825 112.035 108.015 ;
        RECT 112.785 107.870 112.945 107.980 ;
        RECT 113.245 107.825 113.415 108.015 ;
        RECT 114.165 107.845 114.335 108.035 ;
        RECT 114.625 107.845 114.795 108.035 ;
        RECT 115.545 107.870 115.705 107.980 ;
        RECT 116.005 107.845 116.175 108.035 ;
        RECT 126.125 107.825 126.295 108.015 ;
        RECT 127.505 107.825 127.675 108.035 ;
        RECT 14.665 107.015 16.035 107.825 ;
        RECT 16.505 107.015 20.175 107.825 ;
        RECT 20.195 106.915 21.545 107.825 ;
        RECT 22.495 106.915 23.845 107.825 ;
        RECT 24.065 107.145 34.435 107.825 ;
        RECT 24.065 106.915 26.275 107.145 ;
        RECT 28.995 106.925 29.925 107.145 ;
        RECT 34.455 106.915 35.805 107.825 ;
        RECT 35.835 106.915 37.185 107.825 ;
        RECT 37.215 106.955 37.645 107.740 ;
        RECT 38.325 107.145 48.695 107.825 ;
        RECT 38.325 106.915 40.535 107.145 ;
        RECT 43.255 106.925 44.185 107.145 ;
        RECT 48.715 106.915 50.065 107.825 ;
        RECT 50.085 107.045 51.455 107.825 ;
        RECT 51.665 107.145 62.035 107.825 ;
        RECT 51.665 106.915 53.875 107.145 ;
        RECT 56.595 106.925 57.525 107.145 ;
        RECT 62.975 106.955 63.405 107.740 ;
        RECT 63.625 107.145 73.995 107.825 ;
        RECT 75.125 107.145 85.495 107.825 ;
        RECT 63.625 106.915 65.835 107.145 ;
        RECT 68.555 106.925 69.485 107.145 ;
        RECT 75.125 106.915 77.335 107.145 ;
        RECT 80.055 106.925 80.985 107.145 ;
        RECT 85.515 106.915 86.865 107.825 ;
        RECT 86.885 107.045 88.255 107.825 ;
        RECT 88.735 106.955 89.165 107.740 ;
        RECT 89.185 107.145 99.555 107.825 ;
        RECT 93.695 106.925 94.625 107.145 ;
        RECT 97.345 106.915 99.555 107.145 ;
        RECT 100.425 107.145 110.795 107.825 ;
        RECT 100.425 106.915 102.635 107.145 ;
        RECT 105.355 106.925 106.285 107.145 ;
        RECT 110.815 106.915 112.165 107.825 ;
        RECT 113.115 106.915 114.465 107.825 ;
        RECT 114.495 106.955 114.925 107.740 ;
        RECT 116.065 107.145 126.435 107.825 ;
        RECT 116.065 106.915 118.275 107.145 ;
        RECT 120.995 106.925 121.925 107.145 ;
        RECT 126.445 107.015 127.815 107.825 ;
      LAYER nwell ;
        RECT 14.470 103.795 128.010 106.625 ;
      LAYER pwell ;
        RECT 14.665 102.595 16.035 103.405 ;
        RECT 16.045 102.595 18.795 103.405 ;
        RECT 18.805 102.595 24.315 103.405 ;
        RECT 24.335 102.680 24.765 103.465 ;
        RECT 24.785 102.595 26.155 103.405 ;
        RECT 26.175 102.595 27.525 103.505 ;
        RECT 27.545 102.595 28.915 103.375 ;
        RECT 29.125 103.275 31.335 103.505 ;
        RECT 34.055 103.275 34.985 103.495 ;
        RECT 44.015 103.275 44.945 103.495 ;
        RECT 47.665 103.275 49.875 103.505 ;
        RECT 29.125 102.595 39.495 103.275 ;
        RECT 39.505 102.595 49.875 103.275 ;
        RECT 50.095 102.680 50.525 103.465 ;
        RECT 50.545 102.595 51.915 103.405 ;
        RECT 51.925 102.595 55.595 103.405 ;
        RECT 55.615 102.595 56.965 103.505 ;
        RECT 56.985 102.595 58.355 103.405 ;
        RECT 58.565 103.275 60.775 103.505 ;
        RECT 63.495 103.275 64.425 103.495 ;
        RECT 58.565 102.595 68.935 103.275 ;
        RECT 68.945 102.595 70.315 103.405 ;
        RECT 70.325 102.595 75.835 103.405 ;
        RECT 75.855 102.680 76.285 103.465 ;
        RECT 76.505 103.275 78.715 103.505 ;
        RECT 81.435 103.275 82.365 103.495 ;
        RECT 87.085 103.275 89.295 103.505 ;
        RECT 92.015 103.275 92.945 103.495 ;
        RECT 76.505 102.595 86.875 103.275 ;
        RECT 87.085 102.595 97.455 103.275 ;
        RECT 98.395 102.595 99.745 103.505 ;
        RECT 99.765 102.595 101.595 103.405 ;
        RECT 101.615 102.680 102.045 103.465 ;
        RECT 102.065 102.595 103.435 103.405 ;
        RECT 107.955 103.275 108.885 103.495 ;
        RECT 111.605 103.275 113.815 103.505 ;
        RECT 103.445 102.595 113.815 103.275 ;
        RECT 114.225 103.275 116.435 103.505 ;
        RECT 119.155 103.275 120.085 103.495 ;
        RECT 114.225 102.595 124.595 103.275 ;
        RECT 125.065 102.595 126.435 103.375 ;
        RECT 126.445 102.595 127.815 103.405 ;
        RECT 14.805 102.385 14.975 102.595 ;
        RECT 18.485 102.385 18.655 102.595 ;
        RECT 24.005 102.385 24.175 102.595 ;
        RECT 25.845 102.385 26.015 102.595 ;
        RECT 26.305 102.405 26.475 102.595 ;
        RECT 28.605 102.405 28.775 102.595 ;
        RECT 31.365 102.385 31.535 102.575 ;
        RECT 36.885 102.385 37.055 102.575 ;
        RECT 38.725 102.385 38.895 102.575 ;
        RECT 39.185 102.405 39.355 102.595 ;
        RECT 39.645 102.405 39.815 102.595 ;
        RECT 44.245 102.385 44.415 102.575 ;
        RECT 49.765 102.385 49.935 102.575 ;
        RECT 51.605 102.405 51.775 102.595 ;
        RECT 55.285 102.405 55.455 102.595 ;
        RECT 55.745 102.385 55.915 102.575 ;
        RECT 56.665 102.405 56.835 102.595 ;
        RECT 58.045 102.405 58.215 102.595 ;
        RECT 61.265 102.385 61.435 102.575 ;
        RECT 61.725 102.385 61.895 102.575 ;
        RECT 64.025 102.430 64.185 102.540 ;
        RECT 64.485 102.385 64.655 102.575 ;
        RECT 66.325 102.430 66.485 102.540 ;
        RECT 68.625 102.405 68.795 102.595 ;
        RECT 70.005 102.385 70.175 102.595 ;
        RECT 75.525 102.385 75.695 102.595 ;
        RECT 77.365 102.385 77.535 102.575 ;
        RECT 82.885 102.385 83.055 102.575 ;
        RECT 86.565 102.405 86.735 102.595 ;
        RECT 88.405 102.385 88.575 102.575 ;
        RECT 90.245 102.385 90.415 102.575 ;
        RECT 95.765 102.385 95.935 102.575 ;
        RECT 97.145 102.405 97.315 102.595 ;
        RECT 98.065 102.440 98.225 102.550 ;
        RECT 99.445 102.405 99.615 102.595 ;
        RECT 101.285 102.385 101.455 102.595 ;
        RECT 103.125 102.385 103.295 102.595 ;
        RECT 103.585 102.405 103.755 102.595 ;
        RECT 108.645 102.385 108.815 102.575 ;
        RECT 114.165 102.385 114.335 102.575 ;
        RECT 115.140 102.435 115.260 102.545 ;
        RECT 118.765 102.385 118.935 102.575 ;
        RECT 119.225 102.385 119.395 102.575 ;
        RECT 120.660 102.435 120.780 102.545 ;
        RECT 124.285 102.405 124.455 102.595 ;
        RECT 126.115 102.575 126.285 102.595 ;
        RECT 124.800 102.435 124.920 102.545 ;
        RECT 126.115 102.405 126.295 102.575 ;
        RECT 126.125 102.385 126.295 102.405 ;
        RECT 127.505 102.385 127.675 102.595 ;
        RECT 14.665 101.575 16.035 102.385 ;
        RECT 16.045 101.575 18.795 102.385 ;
        RECT 18.805 101.575 24.315 102.385 ;
        RECT 24.335 101.515 24.765 102.300 ;
        RECT 24.785 101.575 26.155 102.385 ;
        RECT 26.165 101.575 31.675 102.385 ;
        RECT 31.685 101.575 37.195 102.385 ;
        RECT 37.215 101.515 37.645 102.300 ;
        RECT 37.665 101.575 39.035 102.385 ;
        RECT 39.045 101.575 44.555 102.385 ;
        RECT 44.565 101.575 50.075 102.385 ;
        RECT 50.095 101.515 50.525 102.300 ;
        RECT 50.545 101.575 56.055 102.385 ;
        RECT 56.065 101.575 61.575 102.385 ;
        RECT 61.595 101.475 62.945 102.385 ;
        RECT 62.975 101.515 63.405 102.300 ;
        RECT 64.355 101.475 65.705 102.385 ;
        RECT 66.645 101.575 70.315 102.385 ;
        RECT 70.325 101.575 75.835 102.385 ;
        RECT 75.855 101.515 76.285 102.300 ;
        RECT 76.305 101.575 77.675 102.385 ;
        RECT 77.685 101.575 83.195 102.385 ;
        RECT 83.205 101.575 88.715 102.385 ;
        RECT 88.735 101.515 89.165 102.300 ;
        RECT 89.185 101.575 90.555 102.385 ;
        RECT 90.565 101.575 96.075 102.385 ;
        RECT 96.085 101.575 101.595 102.385 ;
        RECT 101.615 101.515 102.045 102.300 ;
        RECT 102.065 101.575 103.435 102.385 ;
        RECT 103.445 101.575 108.955 102.385 ;
        RECT 108.965 101.575 114.475 102.385 ;
        RECT 114.495 101.515 114.925 102.300 ;
        RECT 115.405 101.575 119.075 102.385 ;
        RECT 119.095 101.475 120.445 102.385 ;
        RECT 120.925 101.575 126.435 102.385 ;
        RECT 126.445 101.575 127.815 102.385 ;
      LAYER nwell ;
        RECT 14.470 99.580 128.010 101.185 ;
        RECT 20.485 54.580 29.875 66.420 ;
        RECT 31.685 54.590 41.075 66.430 ;
        RECT 42.905 54.560 52.295 66.400 ;
        RECT 54.155 54.540 63.545 66.380 ;
        RECT 65.375 54.530 74.765 66.370 ;
        RECT 76.615 54.520 86.005 66.360 ;
        RECT 87.865 54.530 97.255 66.370 ;
        RECT 99.145 54.520 108.535 66.360 ;
        RECT 110.415 54.520 119.805 66.360 ;
        RECT 121.665 54.520 131.055 66.360 ;
        RECT 132.415 54.490 139.375 66.330 ;
        RECT 20.655 49.020 23.115 53.210 ;
      LAYER pwell ;
        RECT 20.555 45.340 22.915 48.340 ;
      LAYER nwell ;
        RECT 24.735 45.940 29.125 53.130 ;
        RECT 31.855 49.030 34.315 53.220 ;
      LAYER pwell ;
        RECT 31.755 45.350 34.115 48.350 ;
      LAYER nwell ;
        RECT 35.935 45.950 40.325 53.140 ;
        RECT 43.075 49.000 45.535 53.190 ;
      LAYER pwell ;
        RECT 42.975 45.320 45.335 48.320 ;
      LAYER nwell ;
        RECT 47.155 45.920 51.545 53.110 ;
        RECT 54.325 48.980 56.785 53.170 ;
      LAYER pwell ;
        RECT 54.225 45.300 56.585 48.300 ;
      LAYER nwell ;
        RECT 58.405 45.900 62.795 53.090 ;
        RECT 65.545 48.970 68.005 53.160 ;
      LAYER pwell ;
        RECT 65.445 45.290 67.805 48.290 ;
      LAYER nwell ;
        RECT 69.625 45.890 74.015 53.080 ;
        RECT 76.785 48.960 79.245 53.150 ;
      LAYER pwell ;
        RECT 76.685 45.280 79.045 48.280 ;
      LAYER nwell ;
        RECT 80.865 45.880 85.255 53.070 ;
        RECT 88.035 48.970 90.495 53.160 ;
      LAYER pwell ;
        RECT 87.935 45.290 90.295 48.290 ;
      LAYER nwell ;
        RECT 92.115 45.890 96.505 53.080 ;
        RECT 99.315 48.960 101.775 53.150 ;
      LAYER pwell ;
        RECT 99.215 45.280 101.575 48.280 ;
      LAYER nwell ;
        RECT 103.395 45.880 107.785 53.070 ;
        RECT 110.585 48.960 113.045 53.150 ;
      LAYER pwell ;
        RECT 110.485 45.280 112.845 48.280 ;
      LAYER nwell ;
        RECT 114.665 45.880 119.055 53.070 ;
        RECT 121.835 48.960 124.295 53.150 ;
      LAYER pwell ;
        RECT 121.735 45.280 124.095 48.280 ;
      LAYER nwell ;
        RECT 125.915 45.880 130.305 53.070 ;
        RECT 19.615 32.280 24.005 39.470 ;
      LAYER pwell ;
        RECT 25.825 37.070 28.185 40.070 ;
      LAYER nwell ;
        RECT 25.625 32.200 28.085 36.390 ;
        RECT 30.895 32.280 35.285 39.470 ;
      LAYER pwell ;
        RECT 37.105 37.070 39.465 40.070 ;
      LAYER nwell ;
        RECT 36.905 32.200 39.365 36.390 ;
        RECT 42.185 32.260 46.575 39.450 ;
      LAYER pwell ;
        RECT 48.395 37.050 50.755 40.050 ;
      LAYER nwell ;
        RECT 48.195 32.180 50.655 36.370 ;
        RECT 53.405 32.260 57.795 39.450 ;
      LAYER pwell ;
        RECT 59.615 37.050 61.975 40.050 ;
      LAYER nwell ;
        RECT 59.415 32.180 61.875 36.370 ;
        RECT 64.605 32.260 68.995 39.450 ;
      LAYER pwell ;
        RECT 70.815 37.050 73.175 40.050 ;
      LAYER nwell ;
        RECT 70.615 32.180 73.075 36.370 ;
        RECT 75.895 32.250 80.285 39.440 ;
      LAYER pwell ;
        RECT 82.105 37.040 84.465 40.040 ;
      LAYER nwell ;
        RECT 81.905 32.170 84.365 36.360 ;
        RECT 87.135 32.270 91.525 39.460 ;
      LAYER pwell ;
        RECT 93.345 37.060 95.705 40.060 ;
      LAYER nwell ;
        RECT 93.145 32.190 95.605 36.380 ;
        RECT 98.345 32.290 102.735 39.480 ;
      LAYER pwell ;
        RECT 104.555 37.080 106.915 40.080 ;
      LAYER nwell ;
        RECT 104.355 32.210 106.815 36.400 ;
        RECT 109.545 32.330 113.935 39.520 ;
      LAYER pwell ;
        RECT 115.755 37.120 118.115 40.120 ;
      LAYER nwell ;
        RECT 115.555 32.250 118.015 36.440 ;
        RECT 120.755 32.350 125.145 39.540 ;
      LAYER pwell ;
        RECT 126.965 37.140 129.325 40.140 ;
      LAYER nwell ;
        RECT 126.765 32.270 129.225 36.460 ;
        RECT 18.865 18.990 28.255 30.830 ;
        RECT 30.145 18.990 39.535 30.830 ;
        RECT 41.435 18.970 50.825 30.810 ;
        RECT 52.655 18.970 62.045 30.810 ;
        RECT 63.855 18.970 73.245 30.810 ;
        RECT 75.145 18.960 84.535 30.800 ;
        RECT 86.385 18.980 95.775 30.820 ;
        RECT 97.595 19.000 106.985 30.840 ;
        RECT 108.795 19.040 118.185 30.880 ;
        RECT 120.005 19.060 129.395 30.900 ;
        RECT 131.725 19.030 138.685 30.870 ;
      LAYER li1 ;
        RECT 14.660 211.205 127.820 211.375 ;
        RECT 14.745 210.455 15.955 211.205 ;
        RECT 14.745 209.915 15.265 210.455 ;
        RECT 16.125 210.435 18.715 211.205 ;
        RECT 18.890 210.660 24.235 211.205 ;
        RECT 15.435 209.745 15.955 210.285 ;
        RECT 14.745 208.655 15.955 209.745 ;
        RECT 16.125 209.745 17.335 210.265 ;
        RECT 17.505 209.915 18.715 210.435 ;
        RECT 16.125 208.655 18.715 209.745 ;
        RECT 20.480 209.090 20.830 210.340 ;
        RECT 22.310 209.830 22.650 210.660 ;
        RECT 24.405 210.480 24.695 211.205 ;
        RECT 24.865 210.455 26.075 211.205 ;
        RECT 26.250 210.660 31.595 211.205 ;
        RECT 31.770 210.660 37.115 211.205 ;
        RECT 18.890 208.655 24.235 209.090 ;
        RECT 24.405 208.655 24.695 209.820 ;
        RECT 24.865 209.745 25.385 210.285 ;
        RECT 25.555 209.915 26.075 210.455 ;
        RECT 24.865 208.655 26.075 209.745 ;
        RECT 27.840 209.090 28.190 210.340 ;
        RECT 29.670 209.830 30.010 210.660 ;
        RECT 33.360 209.090 33.710 210.340 ;
        RECT 35.190 209.830 35.530 210.660 ;
        RECT 37.285 210.480 37.575 211.205 ;
        RECT 37.745 210.455 38.955 211.205 ;
        RECT 39.130 210.660 44.475 211.205 ;
        RECT 44.650 210.660 49.995 211.205 ;
        RECT 26.250 208.655 31.595 209.090 ;
        RECT 31.770 208.655 37.115 209.090 ;
        RECT 37.285 208.655 37.575 209.820 ;
        RECT 37.745 209.745 38.265 210.285 ;
        RECT 38.435 209.915 38.955 210.455 ;
        RECT 37.745 208.655 38.955 209.745 ;
        RECT 40.720 209.090 41.070 210.340 ;
        RECT 42.550 209.830 42.890 210.660 ;
        RECT 46.240 209.090 46.590 210.340 ;
        RECT 48.070 209.830 48.410 210.660 ;
        RECT 50.165 210.480 50.455 211.205 ;
        RECT 50.625 210.455 51.835 211.205 ;
        RECT 52.010 210.660 57.355 211.205 ;
        RECT 57.530 210.660 62.875 211.205 ;
        RECT 39.130 208.655 44.475 209.090 ;
        RECT 44.650 208.655 49.995 209.090 ;
        RECT 50.165 208.655 50.455 209.820 ;
        RECT 50.625 209.745 51.145 210.285 ;
        RECT 51.315 209.915 51.835 210.455 ;
        RECT 50.625 208.655 51.835 209.745 ;
        RECT 53.600 209.090 53.950 210.340 ;
        RECT 55.430 209.830 55.770 210.660 ;
        RECT 59.120 209.090 59.470 210.340 ;
        RECT 60.950 209.830 61.290 210.660 ;
        RECT 63.045 210.480 63.335 211.205 ;
        RECT 63.505 210.455 64.715 211.205 ;
        RECT 64.890 210.660 70.235 211.205 ;
        RECT 70.410 210.660 75.755 211.205 ;
        RECT 52.010 208.655 57.355 209.090 ;
        RECT 57.530 208.655 62.875 209.090 ;
        RECT 63.045 208.655 63.335 209.820 ;
        RECT 63.505 209.745 64.025 210.285 ;
        RECT 64.195 209.915 64.715 210.455 ;
        RECT 63.505 208.655 64.715 209.745 ;
        RECT 66.480 209.090 66.830 210.340 ;
        RECT 68.310 209.830 68.650 210.660 ;
        RECT 72.000 209.090 72.350 210.340 ;
        RECT 73.830 209.830 74.170 210.660 ;
        RECT 75.925 210.480 76.215 211.205 ;
        RECT 76.385 210.455 77.595 211.205 ;
        RECT 77.770 210.660 83.115 211.205 ;
        RECT 83.290 210.660 88.635 211.205 ;
        RECT 64.890 208.655 70.235 209.090 ;
        RECT 70.410 208.655 75.755 209.090 ;
        RECT 75.925 208.655 76.215 209.820 ;
        RECT 76.385 209.745 76.905 210.285 ;
        RECT 77.075 209.915 77.595 210.455 ;
        RECT 76.385 208.655 77.595 209.745 ;
        RECT 79.360 209.090 79.710 210.340 ;
        RECT 81.190 209.830 81.530 210.660 ;
        RECT 84.880 209.090 85.230 210.340 ;
        RECT 86.710 209.830 87.050 210.660 ;
        RECT 88.805 210.480 89.095 211.205 ;
        RECT 89.265 210.455 90.475 211.205 ;
        RECT 90.650 210.660 95.995 211.205 ;
        RECT 96.170 210.660 101.515 211.205 ;
        RECT 77.770 208.655 83.115 209.090 ;
        RECT 83.290 208.655 88.635 209.090 ;
        RECT 88.805 208.655 89.095 209.820 ;
        RECT 89.265 209.745 89.785 210.285 ;
        RECT 89.955 209.915 90.475 210.455 ;
        RECT 89.265 208.655 90.475 209.745 ;
        RECT 92.240 209.090 92.590 210.340 ;
        RECT 94.070 209.830 94.410 210.660 ;
        RECT 97.760 209.090 98.110 210.340 ;
        RECT 99.590 209.830 99.930 210.660 ;
        RECT 101.685 210.480 101.975 211.205 ;
        RECT 102.145 210.455 103.355 211.205 ;
        RECT 103.530 210.660 108.875 211.205 ;
        RECT 109.050 210.660 114.395 211.205 ;
        RECT 90.650 208.655 95.995 209.090 ;
        RECT 96.170 208.655 101.515 209.090 ;
        RECT 101.685 208.655 101.975 209.820 ;
        RECT 102.145 209.745 102.665 210.285 ;
        RECT 102.835 209.915 103.355 210.455 ;
        RECT 102.145 208.655 103.355 209.745 ;
        RECT 105.120 209.090 105.470 210.340 ;
        RECT 106.950 209.830 107.290 210.660 ;
        RECT 110.640 209.090 110.990 210.340 ;
        RECT 112.470 209.830 112.810 210.660 ;
        RECT 114.565 210.480 114.855 211.205 ;
        RECT 115.490 210.660 120.835 211.205 ;
        RECT 121.010 210.660 126.355 211.205 ;
        RECT 103.530 208.655 108.875 209.090 ;
        RECT 109.050 208.655 114.395 209.090 ;
        RECT 114.565 208.655 114.855 209.820 ;
        RECT 117.080 209.090 117.430 210.340 ;
        RECT 118.910 209.830 119.250 210.660 ;
        RECT 122.600 209.090 122.950 210.340 ;
        RECT 124.430 209.830 124.770 210.660 ;
        RECT 126.525 210.455 127.735 211.205 ;
        RECT 126.525 209.745 127.045 210.285 ;
        RECT 127.215 209.915 127.735 210.455 ;
        RECT 115.490 208.655 120.835 209.090 ;
        RECT 121.010 208.655 126.355 209.090 ;
        RECT 126.525 208.655 127.735 209.745 ;
        RECT 14.660 208.485 127.820 208.655 ;
        RECT 14.745 207.395 15.955 208.485 ;
        RECT 14.745 206.685 15.265 207.225 ;
        RECT 15.435 206.855 15.955 207.395 ;
        RECT 16.125 207.395 18.715 208.485 ;
        RECT 18.890 208.050 24.235 208.485 ;
        RECT 16.125 206.875 17.335 207.395 ;
        RECT 17.505 206.705 18.715 207.225 ;
        RECT 20.480 206.800 20.830 208.050 ;
        RECT 24.405 207.320 24.695 208.485 ;
        RECT 25.325 207.395 27.915 208.485 ;
        RECT 28.090 208.050 33.435 208.485 ;
        RECT 33.610 208.050 38.955 208.485 ;
        RECT 39.130 208.050 44.475 208.485 ;
        RECT 44.650 208.050 49.995 208.485 ;
        RECT 14.745 205.935 15.955 206.685 ;
        RECT 16.125 205.935 18.715 206.705 ;
        RECT 22.310 206.480 22.650 207.310 ;
        RECT 25.325 206.875 26.535 207.395 ;
        RECT 26.705 206.705 27.915 207.225 ;
        RECT 29.680 206.800 30.030 208.050 ;
        RECT 18.890 205.935 24.235 206.480 ;
        RECT 24.405 205.935 24.695 206.660 ;
        RECT 25.325 205.935 27.915 206.705 ;
        RECT 31.510 206.480 31.850 207.310 ;
        RECT 35.200 206.800 35.550 208.050 ;
        RECT 37.030 206.480 37.370 207.310 ;
        RECT 40.720 206.800 41.070 208.050 ;
        RECT 42.550 206.480 42.890 207.310 ;
        RECT 46.240 206.800 46.590 208.050 ;
        RECT 50.165 207.320 50.455 208.485 ;
        RECT 51.085 207.395 53.675 208.485 ;
        RECT 53.850 208.050 59.195 208.485 ;
        RECT 59.370 208.050 64.715 208.485 ;
        RECT 64.890 208.050 70.235 208.485 ;
        RECT 70.410 208.050 75.755 208.485 ;
        RECT 48.070 206.480 48.410 207.310 ;
        RECT 51.085 206.875 52.295 207.395 ;
        RECT 52.465 206.705 53.675 207.225 ;
        RECT 55.440 206.800 55.790 208.050 ;
        RECT 28.090 205.935 33.435 206.480 ;
        RECT 33.610 205.935 38.955 206.480 ;
        RECT 39.130 205.935 44.475 206.480 ;
        RECT 44.650 205.935 49.995 206.480 ;
        RECT 50.165 205.935 50.455 206.660 ;
        RECT 51.085 205.935 53.675 206.705 ;
        RECT 57.270 206.480 57.610 207.310 ;
        RECT 60.960 206.800 61.310 208.050 ;
        RECT 62.790 206.480 63.130 207.310 ;
        RECT 66.480 206.800 66.830 208.050 ;
        RECT 68.310 206.480 68.650 207.310 ;
        RECT 72.000 206.800 72.350 208.050 ;
        RECT 75.925 207.320 76.215 208.485 ;
        RECT 76.845 207.395 79.435 208.485 ;
        RECT 79.610 208.050 84.955 208.485 ;
        RECT 85.130 208.050 90.475 208.485 ;
        RECT 90.650 208.050 95.995 208.485 ;
        RECT 96.170 208.050 101.515 208.485 ;
        RECT 73.830 206.480 74.170 207.310 ;
        RECT 76.845 206.875 78.055 207.395 ;
        RECT 78.225 206.705 79.435 207.225 ;
        RECT 81.200 206.800 81.550 208.050 ;
        RECT 53.850 205.935 59.195 206.480 ;
        RECT 59.370 205.935 64.715 206.480 ;
        RECT 64.890 205.935 70.235 206.480 ;
        RECT 70.410 205.935 75.755 206.480 ;
        RECT 75.925 205.935 76.215 206.660 ;
        RECT 76.845 205.935 79.435 206.705 ;
        RECT 83.030 206.480 83.370 207.310 ;
        RECT 86.720 206.800 87.070 208.050 ;
        RECT 88.550 206.480 88.890 207.310 ;
        RECT 92.240 206.800 92.590 208.050 ;
        RECT 94.070 206.480 94.410 207.310 ;
        RECT 97.760 206.800 98.110 208.050 ;
        RECT 101.685 207.320 101.975 208.485 ;
        RECT 102.605 207.395 104.275 208.485 ;
        RECT 104.450 208.050 109.795 208.485 ;
        RECT 109.970 208.050 115.315 208.485 ;
        RECT 115.490 208.050 120.835 208.485 ;
        RECT 121.010 208.050 126.355 208.485 ;
        RECT 99.590 206.480 99.930 207.310 ;
        RECT 102.605 206.875 103.355 207.395 ;
        RECT 103.525 206.705 104.275 207.225 ;
        RECT 106.040 206.800 106.390 208.050 ;
        RECT 79.610 205.935 84.955 206.480 ;
        RECT 85.130 205.935 90.475 206.480 ;
        RECT 90.650 205.935 95.995 206.480 ;
        RECT 96.170 205.935 101.515 206.480 ;
        RECT 101.685 205.935 101.975 206.660 ;
        RECT 102.605 205.935 104.275 206.705 ;
        RECT 107.870 206.480 108.210 207.310 ;
        RECT 111.560 206.800 111.910 208.050 ;
        RECT 113.390 206.480 113.730 207.310 ;
        RECT 117.080 206.800 117.430 208.050 ;
        RECT 118.910 206.480 119.250 207.310 ;
        RECT 122.600 206.800 122.950 208.050 ;
        RECT 126.525 207.395 127.735 208.485 ;
        RECT 124.430 206.480 124.770 207.310 ;
        RECT 126.525 206.855 127.045 207.395 ;
        RECT 127.215 206.685 127.735 207.225 ;
        RECT 104.450 205.935 109.795 206.480 ;
        RECT 109.970 205.935 115.315 206.480 ;
        RECT 115.490 205.935 120.835 206.480 ;
        RECT 121.010 205.935 126.355 206.480 ;
        RECT 126.525 205.935 127.735 206.685 ;
        RECT 14.660 205.765 127.820 205.935 ;
        RECT 14.745 205.015 15.955 205.765 ;
        RECT 14.745 204.475 15.265 205.015 ;
        RECT 17.045 204.995 20.555 205.765 ;
        RECT 20.730 205.220 26.075 205.765 ;
        RECT 26.250 205.220 31.595 205.765 ;
        RECT 31.770 205.220 37.115 205.765 ;
        RECT 15.435 204.305 15.955 204.845 ;
        RECT 14.745 203.215 15.955 204.305 ;
        RECT 17.045 204.305 18.735 204.825 ;
        RECT 18.905 204.475 20.555 204.995 ;
        RECT 17.045 203.215 20.555 204.305 ;
        RECT 22.320 203.650 22.670 204.900 ;
        RECT 24.150 204.390 24.490 205.220 ;
        RECT 27.840 203.650 28.190 204.900 ;
        RECT 29.670 204.390 30.010 205.220 ;
        RECT 33.360 203.650 33.710 204.900 ;
        RECT 35.190 204.390 35.530 205.220 ;
        RECT 37.285 205.040 37.575 205.765 ;
        RECT 37.745 204.995 39.415 205.765 ;
        RECT 39.590 205.220 44.935 205.765 ;
        RECT 45.110 205.220 50.455 205.765 ;
        RECT 50.630 205.220 55.975 205.765 ;
        RECT 56.150 205.220 61.495 205.765 ;
        RECT 20.730 203.215 26.075 203.650 ;
        RECT 26.250 203.215 31.595 203.650 ;
        RECT 31.770 203.215 37.115 203.650 ;
        RECT 37.285 203.215 37.575 204.380 ;
        RECT 37.745 204.305 38.495 204.825 ;
        RECT 38.665 204.475 39.415 204.995 ;
        RECT 37.745 203.215 39.415 204.305 ;
        RECT 41.180 203.650 41.530 204.900 ;
        RECT 43.010 204.390 43.350 205.220 ;
        RECT 46.700 203.650 47.050 204.900 ;
        RECT 48.530 204.390 48.870 205.220 ;
        RECT 52.220 203.650 52.570 204.900 ;
        RECT 54.050 204.390 54.390 205.220 ;
        RECT 57.740 203.650 58.090 204.900 ;
        RECT 59.570 204.390 59.910 205.220 ;
        RECT 61.725 204.945 61.935 205.765 ;
        RECT 62.105 204.965 62.435 205.595 ;
        RECT 62.105 204.365 62.355 204.965 ;
        RECT 62.605 204.945 62.835 205.765 ;
        RECT 63.045 205.040 63.335 205.765 ;
        RECT 64.465 204.945 64.695 205.765 ;
        RECT 64.865 204.965 65.195 205.595 ;
        RECT 62.525 204.525 62.855 204.775 ;
        RECT 64.445 204.525 64.775 204.775 ;
        RECT 39.590 203.215 44.935 203.650 ;
        RECT 45.110 203.215 50.455 203.650 ;
        RECT 50.630 203.215 55.975 203.650 ;
        RECT 56.150 203.215 61.495 203.650 ;
        RECT 61.725 203.215 61.935 204.355 ;
        RECT 62.105 203.385 62.435 204.365 ;
        RECT 62.605 203.215 62.835 204.355 ;
        RECT 63.045 203.215 63.335 204.380 ;
        RECT 64.945 204.365 65.195 204.965 ;
        RECT 65.365 204.945 65.575 205.765 ;
        RECT 65.810 205.055 66.065 205.585 ;
        RECT 66.235 205.305 66.540 205.765 ;
        RECT 66.785 205.385 67.855 205.555 ;
        RECT 64.465 203.215 64.695 204.355 ;
        RECT 64.865 203.385 65.195 204.365 ;
        RECT 65.810 204.405 66.020 205.055 ;
        RECT 66.785 205.030 67.105 205.385 ;
        RECT 66.780 204.855 67.105 205.030 ;
        RECT 66.190 204.555 67.105 204.855 ;
        RECT 67.275 204.815 67.515 205.215 ;
        RECT 67.685 205.155 67.855 205.385 ;
        RECT 68.025 205.325 68.215 205.765 ;
        RECT 68.385 205.315 69.335 205.595 ;
        RECT 69.555 205.405 69.905 205.575 ;
        RECT 67.685 204.985 68.215 205.155 ;
        RECT 66.190 204.525 66.930 204.555 ;
        RECT 65.365 203.215 65.575 204.355 ;
        RECT 65.810 203.525 66.065 204.405 ;
        RECT 66.235 203.215 66.540 204.355 ;
        RECT 66.760 203.935 66.930 204.525 ;
        RECT 67.275 204.445 67.815 204.815 ;
        RECT 67.995 204.705 68.215 204.985 ;
        RECT 68.385 204.535 68.555 205.315 ;
        RECT 68.150 204.365 68.555 204.535 ;
        RECT 68.725 204.525 69.075 205.145 ;
        RECT 68.150 204.275 68.320 204.365 ;
        RECT 69.245 204.355 69.455 205.145 ;
        RECT 67.100 204.105 68.320 204.275 ;
        RECT 68.780 204.195 69.455 204.355 ;
        RECT 66.760 203.765 67.560 203.935 ;
        RECT 66.880 203.215 67.210 203.595 ;
        RECT 67.390 203.475 67.560 203.765 ;
        RECT 68.150 203.725 68.320 204.105 ;
        RECT 68.490 204.185 69.455 204.195 ;
        RECT 69.645 205.015 69.905 205.405 ;
        RECT 70.115 205.305 70.445 205.765 ;
        RECT 71.320 205.375 72.175 205.545 ;
        RECT 72.380 205.375 72.875 205.545 ;
        RECT 73.045 205.405 73.375 205.765 ;
        RECT 69.645 204.325 69.815 205.015 ;
        RECT 69.985 204.665 70.155 204.845 ;
        RECT 70.325 204.835 71.115 205.085 ;
        RECT 71.320 204.665 71.490 205.375 ;
        RECT 71.660 204.865 72.015 205.085 ;
        RECT 69.985 204.495 71.675 204.665 ;
        RECT 68.490 203.895 68.950 204.185 ;
        RECT 69.645 204.155 71.145 204.325 ;
        RECT 69.645 204.015 69.815 204.155 ;
        RECT 69.255 203.845 69.815 204.015 ;
        RECT 67.730 203.215 67.980 203.675 ;
        RECT 68.150 203.385 69.020 203.725 ;
        RECT 69.255 203.385 69.425 203.845 ;
        RECT 70.260 203.815 71.335 203.985 ;
        RECT 69.595 203.215 69.965 203.675 ;
        RECT 70.260 203.475 70.430 203.815 ;
        RECT 70.600 203.215 70.930 203.645 ;
        RECT 71.165 203.475 71.335 203.815 ;
        RECT 71.505 203.715 71.675 204.495 ;
        RECT 71.845 204.275 72.015 204.865 ;
        RECT 72.185 204.465 72.535 205.085 ;
        RECT 71.845 203.885 72.310 204.275 ;
        RECT 72.705 204.015 72.875 205.375 ;
        RECT 73.045 204.185 73.505 205.235 ;
        RECT 72.480 203.845 72.875 204.015 ;
        RECT 72.480 203.715 72.650 203.845 ;
        RECT 71.505 203.385 72.185 203.715 ;
        RECT 72.400 203.385 72.650 203.715 ;
        RECT 72.820 203.215 73.070 203.675 ;
        RECT 73.240 203.400 73.565 204.185 ;
        RECT 73.735 203.385 73.905 205.505 ;
        RECT 74.075 205.385 74.405 205.765 ;
        RECT 74.575 205.215 74.830 205.505 ;
        RECT 74.080 205.045 74.830 205.215 ;
        RECT 74.080 204.055 74.310 205.045 ;
        RECT 75.005 204.995 77.595 205.765 ;
        RECT 77.770 205.220 83.115 205.765 ;
        RECT 83.290 205.220 88.635 205.765 ;
        RECT 74.480 204.225 74.830 204.875 ;
        RECT 75.005 204.305 76.215 204.825 ;
        RECT 76.385 204.475 77.595 204.995 ;
        RECT 74.080 203.885 74.830 204.055 ;
        RECT 74.075 203.215 74.405 203.715 ;
        RECT 74.575 203.385 74.830 203.885 ;
        RECT 75.005 203.215 77.595 204.305 ;
        RECT 79.360 203.650 79.710 204.900 ;
        RECT 81.190 204.390 81.530 205.220 ;
        RECT 84.880 203.650 85.230 204.900 ;
        RECT 86.710 204.390 87.050 205.220 ;
        RECT 88.805 205.040 89.095 205.765 ;
        RECT 89.725 204.995 92.315 205.765 ;
        RECT 92.490 205.220 97.835 205.765 ;
        RECT 98.010 205.220 103.355 205.765 ;
        RECT 103.530 205.220 108.875 205.765 ;
        RECT 109.050 205.220 114.395 205.765 ;
        RECT 77.770 203.215 83.115 203.650 ;
        RECT 83.290 203.215 88.635 203.650 ;
        RECT 88.805 203.215 89.095 204.380 ;
        RECT 89.725 204.305 90.935 204.825 ;
        RECT 91.105 204.475 92.315 204.995 ;
        RECT 89.725 203.215 92.315 204.305 ;
        RECT 94.080 203.650 94.430 204.900 ;
        RECT 95.910 204.390 96.250 205.220 ;
        RECT 99.600 203.650 99.950 204.900 ;
        RECT 101.430 204.390 101.770 205.220 ;
        RECT 105.120 203.650 105.470 204.900 ;
        RECT 106.950 204.390 107.290 205.220 ;
        RECT 110.640 203.650 110.990 204.900 ;
        RECT 112.470 204.390 112.810 205.220 ;
        RECT 114.565 205.040 114.855 205.765 ;
        RECT 115.490 205.220 120.835 205.765 ;
        RECT 121.010 205.220 126.355 205.765 ;
        RECT 92.490 203.215 97.835 203.650 ;
        RECT 98.010 203.215 103.355 203.650 ;
        RECT 103.530 203.215 108.875 203.650 ;
        RECT 109.050 203.215 114.395 203.650 ;
        RECT 114.565 203.215 114.855 204.380 ;
        RECT 117.080 203.650 117.430 204.900 ;
        RECT 118.910 204.390 119.250 205.220 ;
        RECT 122.600 203.650 122.950 204.900 ;
        RECT 124.430 204.390 124.770 205.220 ;
        RECT 126.525 205.015 127.735 205.765 ;
        RECT 126.525 204.305 127.045 204.845 ;
        RECT 127.215 204.475 127.735 205.015 ;
        RECT 115.490 203.215 120.835 203.650 ;
        RECT 121.010 203.215 126.355 203.650 ;
        RECT 126.525 203.215 127.735 204.305 ;
        RECT 14.660 203.045 127.820 203.215 ;
        RECT 14.745 201.955 15.955 203.045 ;
        RECT 14.745 201.245 15.265 201.785 ;
        RECT 15.435 201.415 15.955 201.955 ;
        RECT 16.125 201.955 18.715 203.045 ;
        RECT 18.890 202.610 24.235 203.045 ;
        RECT 16.125 201.435 17.335 201.955 ;
        RECT 17.505 201.265 18.715 201.785 ;
        RECT 20.480 201.360 20.830 202.610 ;
        RECT 24.405 201.880 24.695 203.045 ;
        RECT 25.325 201.955 27.915 203.045 ;
        RECT 28.090 202.610 33.435 203.045 ;
        RECT 33.610 202.610 38.955 203.045 ;
        RECT 39.130 202.610 44.475 203.045 ;
        RECT 44.650 202.610 49.995 203.045 ;
        RECT 14.745 200.495 15.955 201.245 ;
        RECT 16.125 200.495 18.715 201.265 ;
        RECT 22.310 201.040 22.650 201.870 ;
        RECT 25.325 201.435 26.535 201.955 ;
        RECT 26.705 201.265 27.915 201.785 ;
        RECT 29.680 201.360 30.030 202.610 ;
        RECT 18.890 200.495 24.235 201.040 ;
        RECT 24.405 200.495 24.695 201.220 ;
        RECT 25.325 200.495 27.915 201.265 ;
        RECT 31.510 201.040 31.850 201.870 ;
        RECT 35.200 201.360 35.550 202.610 ;
        RECT 37.030 201.040 37.370 201.870 ;
        RECT 40.720 201.360 41.070 202.610 ;
        RECT 42.550 201.040 42.890 201.870 ;
        RECT 46.240 201.360 46.590 202.610 ;
        RECT 50.165 201.880 50.455 203.045 ;
        RECT 51.085 201.955 52.755 203.045 ;
        RECT 52.930 202.610 58.275 203.045 ;
        RECT 48.070 201.040 48.410 201.870 ;
        RECT 51.085 201.435 51.835 201.955 ;
        RECT 52.005 201.265 52.755 201.785 ;
        RECT 54.520 201.360 54.870 202.610 ;
        RECT 58.755 202.205 58.925 203.045 ;
        RECT 59.135 202.035 59.385 202.875 ;
        RECT 59.595 202.205 59.765 203.045 ;
        RECT 59.935 202.035 60.225 202.875 ;
        RECT 28.090 200.495 33.435 201.040 ;
        RECT 33.610 200.495 38.955 201.040 ;
        RECT 39.130 200.495 44.475 201.040 ;
        RECT 44.650 200.495 49.995 201.040 ;
        RECT 50.165 200.495 50.455 201.220 ;
        RECT 51.085 200.495 52.755 201.265 ;
        RECT 56.350 201.040 56.690 201.870 ;
        RECT 58.500 201.865 60.225 202.035 ;
        RECT 60.435 201.985 60.605 203.045 ;
        RECT 60.900 202.665 61.230 203.045 ;
        RECT 61.410 202.495 61.580 202.785 ;
        RECT 61.750 202.585 62.000 203.045 ;
        RECT 60.780 202.325 61.580 202.495 ;
        RECT 62.170 202.535 63.040 202.875 ;
        RECT 58.500 201.315 58.910 201.865 ;
        RECT 60.780 201.705 60.950 202.325 ;
        RECT 62.170 202.155 62.340 202.535 ;
        RECT 63.275 202.415 63.445 202.875 ;
        RECT 63.615 202.585 63.985 203.045 ;
        RECT 64.280 202.445 64.450 202.785 ;
        RECT 64.620 202.615 64.950 203.045 ;
        RECT 65.185 202.445 65.355 202.785 ;
        RECT 61.120 201.985 62.340 202.155 ;
        RECT 62.510 202.075 62.970 202.365 ;
        RECT 63.275 202.245 63.835 202.415 ;
        RECT 64.280 202.275 65.355 202.445 ;
        RECT 65.525 202.545 66.205 202.875 ;
        RECT 66.420 202.545 66.670 202.875 ;
        RECT 66.840 202.585 67.090 203.045 ;
        RECT 63.665 202.105 63.835 202.245 ;
        RECT 62.510 202.065 63.475 202.075 ;
        RECT 62.170 201.895 62.340 201.985 ;
        RECT 62.800 201.905 63.475 202.065 ;
        RECT 60.780 201.695 61.125 201.705 ;
        RECT 59.095 201.485 61.125 201.695 ;
        RECT 58.500 201.145 60.265 201.315 ;
        RECT 52.930 200.495 58.275 201.040 ;
        RECT 58.755 200.495 58.925 200.965 ;
        RECT 59.095 200.665 59.425 201.145 ;
        RECT 59.595 200.495 59.765 200.965 ;
        RECT 59.935 200.665 60.265 201.145 ;
        RECT 60.435 200.495 60.605 201.305 ;
        RECT 60.800 201.230 61.125 201.485 ;
        RECT 60.805 200.875 61.125 201.230 ;
        RECT 61.295 201.445 61.835 201.815 ;
        RECT 62.170 201.725 62.575 201.895 ;
        RECT 61.295 201.045 61.535 201.445 ;
        RECT 62.015 201.275 62.235 201.555 ;
        RECT 61.705 201.105 62.235 201.275 ;
        RECT 61.705 200.875 61.875 201.105 ;
        RECT 62.405 200.945 62.575 201.725 ;
        RECT 62.745 201.115 63.095 201.735 ;
        RECT 63.265 201.115 63.475 201.905 ;
        RECT 63.665 201.935 65.165 202.105 ;
        RECT 63.665 201.245 63.835 201.935 ;
        RECT 65.525 201.765 65.695 202.545 ;
        RECT 66.500 202.415 66.670 202.545 ;
        RECT 64.005 201.595 65.695 201.765 ;
        RECT 65.865 201.985 66.330 202.375 ;
        RECT 66.500 202.245 66.895 202.415 ;
        RECT 64.005 201.415 64.175 201.595 ;
        RECT 60.805 200.705 61.875 200.875 ;
        RECT 62.045 200.495 62.235 200.935 ;
        RECT 62.405 200.665 63.355 200.945 ;
        RECT 63.665 200.855 63.925 201.245 ;
        RECT 64.345 201.175 65.135 201.425 ;
        RECT 63.575 200.685 63.925 200.855 ;
        RECT 64.135 200.495 64.465 200.955 ;
        RECT 65.340 200.885 65.510 201.595 ;
        RECT 65.865 201.395 66.035 201.985 ;
        RECT 65.680 201.175 66.035 201.395 ;
        RECT 66.205 201.175 66.555 201.795 ;
        RECT 66.725 200.885 66.895 202.245 ;
        RECT 67.260 202.075 67.585 202.860 ;
        RECT 67.065 201.025 67.525 202.075 ;
        RECT 65.340 200.715 66.195 200.885 ;
        RECT 66.400 200.715 66.895 200.885 ;
        RECT 67.065 200.495 67.395 200.855 ;
        RECT 67.755 200.755 67.925 202.875 ;
        RECT 68.095 202.545 68.425 203.045 ;
        RECT 68.595 202.375 68.850 202.875 ;
        RECT 68.100 202.205 68.850 202.375 ;
        RECT 68.100 201.215 68.330 202.205 ;
        RECT 68.500 201.385 68.850 202.035 ;
        RECT 69.485 201.955 72.075 203.045 ;
        RECT 72.335 202.115 72.505 202.875 ;
        RECT 72.685 202.285 73.015 203.045 ;
        RECT 69.485 201.435 70.695 201.955 ;
        RECT 72.335 201.945 73.000 202.115 ;
        RECT 73.185 201.970 73.455 202.875 ;
        RECT 72.830 201.800 73.000 201.945 ;
        RECT 70.865 201.265 72.075 201.785 ;
        RECT 72.265 201.395 72.595 201.765 ;
        RECT 72.830 201.470 73.115 201.800 ;
        RECT 68.100 201.045 68.850 201.215 ;
        RECT 68.095 200.495 68.425 200.875 ;
        RECT 68.595 200.755 68.850 201.045 ;
        RECT 69.485 200.495 72.075 201.265 ;
        RECT 72.830 201.215 73.000 201.470 ;
        RECT 72.335 201.045 73.000 201.215 ;
        RECT 73.285 201.170 73.455 201.970 ;
        RECT 74.585 201.905 74.815 203.045 ;
        RECT 74.985 201.895 75.315 202.875 ;
        RECT 75.485 201.905 75.695 203.045 ;
        RECT 74.565 201.485 74.895 201.735 ;
        RECT 72.335 200.665 72.505 201.045 ;
        RECT 72.685 200.495 73.015 200.875 ;
        RECT 73.195 200.665 73.455 201.170 ;
        RECT 74.585 200.495 74.815 201.315 ;
        RECT 75.065 201.295 75.315 201.895 ;
        RECT 75.925 201.880 76.215 203.045 ;
        RECT 76.385 201.955 78.055 203.045 ;
        RECT 78.230 202.610 83.575 203.045 ;
        RECT 83.750 202.610 89.095 203.045 ;
        RECT 89.270 202.610 94.615 203.045 ;
        RECT 94.790 202.610 100.135 203.045 ;
        RECT 76.385 201.435 77.135 201.955 ;
        RECT 74.985 200.665 75.315 201.295 ;
        RECT 75.485 200.495 75.695 201.315 ;
        RECT 77.305 201.265 78.055 201.785 ;
        RECT 79.820 201.360 80.170 202.610 ;
        RECT 75.925 200.495 76.215 201.220 ;
        RECT 76.385 200.495 78.055 201.265 ;
        RECT 81.650 201.040 81.990 201.870 ;
        RECT 85.340 201.360 85.690 202.610 ;
        RECT 87.170 201.040 87.510 201.870 ;
        RECT 90.860 201.360 91.210 202.610 ;
        RECT 92.690 201.040 93.030 201.870 ;
        RECT 96.380 201.360 96.730 202.610 ;
        RECT 100.345 201.905 100.575 203.045 ;
        RECT 100.745 201.895 101.075 202.875 ;
        RECT 101.245 201.905 101.455 203.045 ;
        RECT 98.210 201.040 98.550 201.870 ;
        RECT 100.325 201.485 100.655 201.735 ;
        RECT 78.230 200.495 83.575 201.040 ;
        RECT 83.750 200.495 89.095 201.040 ;
        RECT 89.270 200.495 94.615 201.040 ;
        RECT 94.790 200.495 100.135 201.040 ;
        RECT 100.345 200.495 100.575 201.315 ;
        RECT 100.825 201.295 101.075 201.895 ;
        RECT 101.685 201.880 101.975 203.045 ;
        RECT 102.145 201.955 103.815 203.045 ;
        RECT 102.145 201.435 102.895 201.955 ;
        RECT 103.990 201.855 104.245 202.735 ;
        RECT 104.415 201.905 104.720 203.045 ;
        RECT 105.060 202.665 105.390 203.045 ;
        RECT 105.570 202.495 105.740 202.785 ;
        RECT 105.910 202.585 106.160 203.045 ;
        RECT 104.940 202.325 105.740 202.495 ;
        RECT 106.330 202.535 107.200 202.875 ;
        RECT 100.745 200.665 101.075 201.295 ;
        RECT 101.245 200.495 101.455 201.315 ;
        RECT 103.065 201.265 103.815 201.785 ;
        RECT 101.685 200.495 101.975 201.220 ;
        RECT 102.145 200.495 103.815 201.265 ;
        RECT 103.990 201.205 104.200 201.855 ;
        RECT 104.940 201.735 105.110 202.325 ;
        RECT 106.330 202.155 106.500 202.535 ;
        RECT 107.435 202.415 107.605 202.875 ;
        RECT 107.775 202.585 108.145 203.045 ;
        RECT 108.440 202.445 108.610 202.785 ;
        RECT 108.780 202.615 109.110 203.045 ;
        RECT 109.345 202.445 109.515 202.785 ;
        RECT 105.280 201.985 106.500 202.155 ;
        RECT 106.670 202.075 107.130 202.365 ;
        RECT 107.435 202.245 107.995 202.415 ;
        RECT 108.440 202.275 109.515 202.445 ;
        RECT 109.685 202.545 110.365 202.875 ;
        RECT 110.580 202.545 110.830 202.875 ;
        RECT 111.000 202.585 111.250 203.045 ;
        RECT 107.825 202.105 107.995 202.245 ;
        RECT 106.670 202.065 107.635 202.075 ;
        RECT 106.330 201.895 106.500 201.985 ;
        RECT 106.960 201.905 107.635 202.065 ;
        RECT 104.370 201.705 105.110 201.735 ;
        RECT 104.370 201.405 105.285 201.705 ;
        RECT 104.960 201.230 105.285 201.405 ;
        RECT 103.990 200.675 104.245 201.205 ;
        RECT 104.415 200.495 104.720 200.955 ;
        RECT 104.965 200.875 105.285 201.230 ;
        RECT 105.455 201.445 105.995 201.815 ;
        RECT 106.330 201.725 106.735 201.895 ;
        RECT 105.455 201.045 105.695 201.445 ;
        RECT 106.175 201.275 106.395 201.555 ;
        RECT 105.865 201.105 106.395 201.275 ;
        RECT 105.865 200.875 106.035 201.105 ;
        RECT 106.565 200.945 106.735 201.725 ;
        RECT 106.905 201.115 107.255 201.735 ;
        RECT 107.425 201.115 107.635 201.905 ;
        RECT 107.825 201.935 109.325 202.105 ;
        RECT 107.825 201.245 107.995 201.935 ;
        RECT 109.685 201.765 109.855 202.545 ;
        RECT 110.660 202.415 110.830 202.545 ;
        RECT 108.165 201.595 109.855 201.765 ;
        RECT 110.025 201.985 110.490 202.375 ;
        RECT 110.660 202.245 111.055 202.415 ;
        RECT 108.165 201.415 108.335 201.595 ;
        RECT 104.965 200.705 106.035 200.875 ;
        RECT 106.205 200.495 106.395 200.935 ;
        RECT 106.565 200.665 107.515 200.945 ;
        RECT 107.825 200.855 108.085 201.245 ;
        RECT 108.505 201.175 109.295 201.425 ;
        RECT 107.735 200.685 108.085 200.855 ;
        RECT 108.295 200.495 108.625 200.955 ;
        RECT 109.500 200.885 109.670 201.595 ;
        RECT 110.025 201.395 110.195 201.985 ;
        RECT 109.840 201.175 110.195 201.395 ;
        RECT 110.365 201.175 110.715 201.795 ;
        RECT 110.885 200.885 111.055 202.245 ;
        RECT 111.420 202.075 111.745 202.860 ;
        RECT 111.225 201.025 111.685 202.075 ;
        RECT 109.500 200.715 110.355 200.885 ;
        RECT 110.560 200.715 111.055 200.885 ;
        RECT 111.225 200.495 111.555 200.855 ;
        RECT 111.915 200.755 112.085 202.875 ;
        RECT 112.255 202.545 112.585 203.045 ;
        RECT 112.755 202.375 113.010 202.875 ;
        RECT 112.260 202.205 113.010 202.375 ;
        RECT 112.260 201.215 112.490 202.205 ;
        RECT 112.660 201.385 113.010 202.035 ;
        RECT 113.645 201.955 115.315 203.045 ;
        RECT 115.490 202.610 120.835 203.045 ;
        RECT 121.010 202.610 126.355 203.045 ;
        RECT 113.645 201.435 114.395 201.955 ;
        RECT 114.565 201.265 115.315 201.785 ;
        RECT 117.080 201.360 117.430 202.610 ;
        RECT 112.260 201.045 113.010 201.215 ;
        RECT 112.255 200.495 112.585 200.875 ;
        RECT 112.755 200.755 113.010 201.045 ;
        RECT 113.645 200.495 115.315 201.265 ;
        RECT 118.910 201.040 119.250 201.870 ;
        RECT 122.600 201.360 122.950 202.610 ;
        RECT 126.525 201.955 127.735 203.045 ;
        RECT 124.430 201.040 124.770 201.870 ;
        RECT 126.525 201.415 127.045 201.955 ;
        RECT 127.215 201.245 127.735 201.785 ;
        RECT 115.490 200.495 120.835 201.040 ;
        RECT 121.010 200.495 126.355 201.040 ;
        RECT 126.525 200.495 127.735 201.245 ;
        RECT 14.660 200.325 127.820 200.495 ;
        RECT 14.745 199.575 15.955 200.325 ;
        RECT 14.745 199.035 15.265 199.575 ;
        RECT 17.045 199.555 20.555 200.325 ;
        RECT 20.730 199.780 26.075 200.325 ;
        RECT 26.250 199.780 31.595 200.325 ;
        RECT 31.770 199.780 37.115 200.325 ;
        RECT 15.435 198.865 15.955 199.405 ;
        RECT 14.745 197.775 15.955 198.865 ;
        RECT 17.045 198.865 18.735 199.385 ;
        RECT 18.905 199.035 20.555 199.555 ;
        RECT 17.045 197.775 20.555 198.865 ;
        RECT 22.320 198.210 22.670 199.460 ;
        RECT 24.150 198.950 24.490 199.780 ;
        RECT 27.840 198.210 28.190 199.460 ;
        RECT 29.670 198.950 30.010 199.780 ;
        RECT 33.360 198.210 33.710 199.460 ;
        RECT 35.190 198.950 35.530 199.780 ;
        RECT 37.285 199.600 37.575 200.325 ;
        RECT 38.205 199.555 40.795 200.325 ;
        RECT 40.970 199.780 46.315 200.325 ;
        RECT 46.490 199.780 51.835 200.325 ;
        RECT 52.010 199.780 57.355 200.325 ;
        RECT 57.530 199.780 62.875 200.325 ;
        RECT 20.730 197.775 26.075 198.210 ;
        RECT 26.250 197.775 31.595 198.210 ;
        RECT 31.770 197.775 37.115 198.210 ;
        RECT 37.285 197.775 37.575 198.940 ;
        RECT 38.205 198.865 39.415 199.385 ;
        RECT 39.585 199.035 40.795 199.555 ;
        RECT 38.205 197.775 40.795 198.865 ;
        RECT 42.560 198.210 42.910 199.460 ;
        RECT 44.390 198.950 44.730 199.780 ;
        RECT 48.080 198.210 48.430 199.460 ;
        RECT 49.910 198.950 50.250 199.780 ;
        RECT 53.600 198.210 53.950 199.460 ;
        RECT 55.430 198.950 55.770 199.780 ;
        RECT 59.120 198.210 59.470 199.460 ;
        RECT 60.950 198.950 61.290 199.780 ;
        RECT 63.045 199.600 63.335 200.325 ;
        RECT 63.965 199.555 66.555 200.325 ;
        RECT 66.815 199.775 66.985 200.155 ;
        RECT 67.165 199.945 67.495 200.325 ;
        RECT 66.815 199.605 67.480 199.775 ;
        RECT 67.675 199.650 67.935 200.155 ;
        RECT 40.970 197.775 46.315 198.210 ;
        RECT 46.490 197.775 51.835 198.210 ;
        RECT 52.010 197.775 57.355 198.210 ;
        RECT 57.530 197.775 62.875 198.210 ;
        RECT 63.045 197.775 63.335 198.940 ;
        RECT 63.965 198.865 65.175 199.385 ;
        RECT 65.345 199.035 66.555 199.555 ;
        RECT 66.745 199.055 67.075 199.425 ;
        RECT 67.310 199.350 67.480 199.605 ;
        RECT 67.310 199.020 67.595 199.350 ;
        RECT 67.310 198.875 67.480 199.020 ;
        RECT 63.965 197.775 66.555 198.865 ;
        RECT 66.815 198.705 67.480 198.875 ;
        RECT 67.765 198.850 67.935 199.650 ;
        RECT 68.105 199.555 69.775 200.325 ;
        RECT 66.815 197.945 66.985 198.705 ;
        RECT 67.165 197.775 67.495 198.535 ;
        RECT 67.665 197.945 67.935 198.850 ;
        RECT 68.105 198.865 68.855 199.385 ;
        RECT 69.025 199.035 69.775 199.555 ;
        RECT 69.945 199.675 70.205 200.155 ;
        RECT 70.375 199.785 70.625 200.325 ;
        RECT 68.105 197.775 69.775 198.865 ;
        RECT 69.945 198.645 70.115 199.675 ;
        RECT 70.795 199.645 71.015 200.105 ;
        RECT 70.765 199.620 71.015 199.645 ;
        RECT 70.285 199.025 70.515 199.420 ;
        RECT 70.685 199.195 71.015 199.620 ;
        RECT 71.185 199.945 72.075 200.115 ;
        RECT 71.185 199.220 71.355 199.945 ;
        RECT 71.525 199.390 72.075 199.775 ;
        RECT 72.250 199.615 72.505 200.145 ;
        RECT 72.675 199.865 72.980 200.325 ;
        RECT 73.225 199.945 74.295 200.115 ;
        RECT 71.185 199.150 72.075 199.220 ;
        RECT 71.180 199.125 72.075 199.150 ;
        RECT 71.170 199.110 72.075 199.125 ;
        RECT 71.165 199.095 72.075 199.110 ;
        RECT 71.155 199.090 72.075 199.095 ;
        RECT 71.150 199.080 72.075 199.090 ;
        RECT 71.145 199.070 72.075 199.080 ;
        RECT 71.135 199.065 72.075 199.070 ;
        RECT 71.125 199.055 72.075 199.065 ;
        RECT 71.115 199.050 72.075 199.055 ;
        RECT 71.115 199.045 71.450 199.050 ;
        RECT 71.100 199.040 71.450 199.045 ;
        RECT 71.085 199.030 71.450 199.040 ;
        RECT 71.060 199.025 71.450 199.030 ;
        RECT 70.285 199.020 71.450 199.025 ;
        RECT 70.285 198.985 71.420 199.020 ;
        RECT 70.285 198.960 71.385 198.985 ;
        RECT 70.285 198.930 71.355 198.960 ;
        RECT 70.285 198.900 71.335 198.930 ;
        RECT 70.285 198.870 71.315 198.900 ;
        RECT 70.285 198.860 71.245 198.870 ;
        RECT 70.285 198.850 71.220 198.860 ;
        RECT 70.285 198.835 71.200 198.850 ;
        RECT 70.285 198.820 71.180 198.835 ;
        RECT 70.390 198.810 71.175 198.820 ;
        RECT 70.390 198.775 71.160 198.810 ;
        RECT 69.945 197.945 70.220 198.645 ;
        RECT 70.390 198.525 71.145 198.775 ;
        RECT 71.315 198.455 71.645 198.700 ;
        RECT 71.815 198.600 72.075 199.050 ;
        RECT 72.250 198.965 72.460 199.615 ;
        RECT 73.225 199.590 73.545 199.945 ;
        RECT 73.220 199.415 73.545 199.590 ;
        RECT 72.630 199.115 73.545 199.415 ;
        RECT 73.715 199.375 73.955 199.775 ;
        RECT 74.125 199.715 74.295 199.945 ;
        RECT 74.465 199.885 74.655 200.325 ;
        RECT 74.825 199.875 75.775 200.155 ;
        RECT 75.995 199.965 76.345 200.135 ;
        RECT 74.125 199.545 74.655 199.715 ;
        RECT 72.630 199.085 73.370 199.115 ;
        RECT 71.460 198.430 71.645 198.455 ;
        RECT 71.460 198.330 72.075 198.430 ;
        RECT 70.390 197.775 70.645 198.320 ;
        RECT 70.815 197.945 71.295 198.285 ;
        RECT 71.470 197.775 72.075 198.330 ;
        RECT 72.250 198.085 72.505 198.965 ;
        RECT 72.675 197.775 72.980 198.915 ;
        RECT 73.200 198.495 73.370 199.085 ;
        RECT 73.715 199.005 74.255 199.375 ;
        RECT 74.435 199.265 74.655 199.545 ;
        RECT 74.825 199.095 74.995 199.875 ;
        RECT 74.590 198.925 74.995 199.095 ;
        RECT 75.165 199.085 75.515 199.705 ;
        RECT 74.590 198.835 74.760 198.925 ;
        RECT 75.685 198.915 75.895 199.705 ;
        RECT 73.540 198.665 74.760 198.835 ;
        RECT 75.220 198.755 75.895 198.915 ;
        RECT 73.200 198.325 74.000 198.495 ;
        RECT 73.320 197.775 73.650 198.155 ;
        RECT 73.830 198.035 74.000 198.325 ;
        RECT 74.590 198.285 74.760 198.665 ;
        RECT 74.930 198.745 75.895 198.755 ;
        RECT 76.085 199.575 76.345 199.965 ;
        RECT 76.555 199.865 76.885 200.325 ;
        RECT 77.760 199.935 78.615 200.105 ;
        RECT 78.820 199.935 79.315 200.105 ;
        RECT 79.485 199.965 79.815 200.325 ;
        RECT 76.085 198.885 76.255 199.575 ;
        RECT 76.425 199.225 76.595 199.405 ;
        RECT 76.765 199.395 77.555 199.645 ;
        RECT 77.760 199.225 77.930 199.935 ;
        RECT 78.100 199.425 78.455 199.645 ;
        RECT 76.425 199.055 78.115 199.225 ;
        RECT 74.930 198.455 75.390 198.745 ;
        RECT 76.085 198.715 77.585 198.885 ;
        RECT 76.085 198.575 76.255 198.715 ;
        RECT 75.695 198.405 76.255 198.575 ;
        RECT 74.170 197.775 74.420 198.235 ;
        RECT 74.590 197.945 75.460 198.285 ;
        RECT 75.695 197.945 75.865 198.405 ;
        RECT 76.700 198.375 77.775 198.545 ;
        RECT 76.035 197.775 76.405 198.235 ;
        RECT 76.700 198.035 76.870 198.375 ;
        RECT 77.040 197.775 77.370 198.205 ;
        RECT 77.605 198.035 77.775 198.375 ;
        RECT 77.945 198.275 78.115 199.055 ;
        RECT 78.285 198.835 78.455 199.425 ;
        RECT 78.625 199.025 78.975 199.645 ;
        RECT 78.285 198.445 78.750 198.835 ;
        RECT 79.145 198.575 79.315 199.935 ;
        RECT 79.485 198.745 79.945 199.795 ;
        RECT 78.920 198.405 79.315 198.575 ;
        RECT 78.920 198.275 79.090 198.405 ;
        RECT 77.945 197.945 78.625 198.275 ;
        RECT 78.840 197.945 79.090 198.275 ;
        RECT 79.260 197.775 79.510 198.235 ;
        RECT 79.680 197.960 80.005 198.745 ;
        RECT 80.175 197.945 80.345 200.065 ;
        RECT 80.515 199.945 80.845 200.325 ;
        RECT 81.015 199.775 81.270 200.065 ;
        RECT 81.910 199.780 87.255 200.325 ;
        RECT 80.520 199.605 81.270 199.775 ;
        RECT 80.520 198.615 80.750 199.605 ;
        RECT 80.920 198.785 81.270 199.435 ;
        RECT 80.520 198.445 81.270 198.615 ;
        RECT 80.515 197.775 80.845 198.275 ;
        RECT 81.015 197.945 81.270 198.445 ;
        RECT 83.500 198.210 83.850 199.460 ;
        RECT 85.330 198.950 85.670 199.780 ;
        RECT 87.465 199.505 87.695 200.325 ;
        RECT 87.865 199.525 88.195 200.155 ;
        RECT 87.445 199.085 87.775 199.335 ;
        RECT 87.945 198.925 88.195 199.525 ;
        RECT 88.365 199.505 88.575 200.325 ;
        RECT 88.805 199.600 89.095 200.325 ;
        RECT 89.270 199.615 89.525 200.145 ;
        RECT 89.695 199.865 90.000 200.325 ;
        RECT 90.245 199.945 91.315 200.115 ;
        RECT 89.270 198.965 89.480 199.615 ;
        RECT 90.245 199.590 90.565 199.945 ;
        RECT 90.240 199.415 90.565 199.590 ;
        RECT 89.650 199.115 90.565 199.415 ;
        RECT 90.735 199.375 90.975 199.775 ;
        RECT 91.145 199.715 91.315 199.945 ;
        RECT 91.485 199.885 91.675 200.325 ;
        RECT 91.845 199.875 92.795 200.155 ;
        RECT 93.015 199.965 93.365 200.135 ;
        RECT 91.145 199.545 91.675 199.715 ;
        RECT 89.650 199.085 90.390 199.115 ;
        RECT 81.910 197.775 87.255 198.210 ;
        RECT 87.465 197.775 87.695 198.915 ;
        RECT 87.865 197.945 88.195 198.925 ;
        RECT 88.365 197.775 88.575 198.915 ;
        RECT 88.805 197.775 89.095 198.940 ;
        RECT 89.270 198.085 89.525 198.965 ;
        RECT 89.695 197.775 90.000 198.915 ;
        RECT 90.220 198.495 90.390 199.085 ;
        RECT 90.735 199.005 91.275 199.375 ;
        RECT 91.455 199.265 91.675 199.545 ;
        RECT 91.845 199.095 92.015 199.875 ;
        RECT 91.610 198.925 92.015 199.095 ;
        RECT 92.185 199.085 92.535 199.705 ;
        RECT 91.610 198.835 91.780 198.925 ;
        RECT 92.705 198.915 92.915 199.705 ;
        RECT 90.560 198.665 91.780 198.835 ;
        RECT 92.240 198.755 92.915 198.915 ;
        RECT 90.220 198.325 91.020 198.495 ;
        RECT 90.340 197.775 90.670 198.155 ;
        RECT 90.850 198.035 91.020 198.325 ;
        RECT 91.610 198.285 91.780 198.665 ;
        RECT 91.950 198.745 92.915 198.755 ;
        RECT 93.105 199.575 93.365 199.965 ;
        RECT 93.575 199.865 93.905 200.325 ;
        RECT 94.780 199.935 95.635 200.105 ;
        RECT 95.840 199.935 96.335 200.105 ;
        RECT 96.505 199.965 96.835 200.325 ;
        RECT 93.105 198.885 93.275 199.575 ;
        RECT 93.445 199.225 93.615 199.405 ;
        RECT 93.785 199.395 94.575 199.645 ;
        RECT 94.780 199.225 94.950 199.935 ;
        RECT 95.120 199.425 95.475 199.645 ;
        RECT 93.445 199.055 95.135 199.225 ;
        RECT 91.950 198.455 92.410 198.745 ;
        RECT 93.105 198.715 94.605 198.885 ;
        RECT 93.105 198.575 93.275 198.715 ;
        RECT 92.715 198.405 93.275 198.575 ;
        RECT 91.190 197.775 91.440 198.235 ;
        RECT 91.610 197.945 92.480 198.285 ;
        RECT 92.715 197.945 92.885 198.405 ;
        RECT 93.720 198.375 94.795 198.545 ;
        RECT 93.055 197.775 93.425 198.235 ;
        RECT 93.720 198.035 93.890 198.375 ;
        RECT 94.060 197.775 94.390 198.205 ;
        RECT 94.625 198.035 94.795 198.375 ;
        RECT 94.965 198.275 95.135 199.055 ;
        RECT 95.305 198.835 95.475 199.425 ;
        RECT 95.645 199.025 95.995 199.645 ;
        RECT 95.305 198.445 95.770 198.835 ;
        RECT 96.165 198.575 96.335 199.935 ;
        RECT 96.505 198.745 96.965 199.795 ;
        RECT 95.940 198.405 96.335 198.575 ;
        RECT 95.940 198.275 96.110 198.405 ;
        RECT 94.965 197.945 95.645 198.275 ;
        RECT 95.860 197.945 96.110 198.275 ;
        RECT 96.280 197.775 96.530 198.235 ;
        RECT 96.700 197.960 97.025 198.745 ;
        RECT 97.195 197.945 97.365 200.065 ;
        RECT 97.535 199.945 97.865 200.325 ;
        RECT 98.035 199.775 98.290 200.065 ;
        RECT 97.540 199.605 98.290 199.775 ;
        RECT 98.470 199.615 98.725 200.145 ;
        RECT 98.895 199.865 99.200 200.325 ;
        RECT 99.445 199.945 100.515 200.115 ;
        RECT 97.540 198.615 97.770 199.605 ;
        RECT 97.940 198.785 98.290 199.435 ;
        RECT 98.470 198.965 98.680 199.615 ;
        RECT 99.445 199.590 99.765 199.945 ;
        RECT 99.440 199.415 99.765 199.590 ;
        RECT 98.850 199.115 99.765 199.415 ;
        RECT 99.935 199.375 100.175 199.775 ;
        RECT 100.345 199.715 100.515 199.945 ;
        RECT 100.685 199.885 100.875 200.325 ;
        RECT 101.045 199.875 101.995 200.155 ;
        RECT 102.215 199.965 102.565 200.135 ;
        RECT 100.345 199.545 100.875 199.715 ;
        RECT 98.850 199.085 99.590 199.115 ;
        RECT 97.540 198.445 98.290 198.615 ;
        RECT 97.535 197.775 97.865 198.275 ;
        RECT 98.035 197.945 98.290 198.445 ;
        RECT 98.470 198.085 98.725 198.965 ;
        RECT 98.895 197.775 99.200 198.915 ;
        RECT 99.420 198.495 99.590 199.085 ;
        RECT 99.935 199.005 100.475 199.375 ;
        RECT 100.655 199.265 100.875 199.545 ;
        RECT 101.045 199.095 101.215 199.875 ;
        RECT 100.810 198.925 101.215 199.095 ;
        RECT 101.385 199.085 101.735 199.705 ;
        RECT 100.810 198.835 100.980 198.925 ;
        RECT 101.905 198.915 102.115 199.705 ;
        RECT 99.760 198.665 100.980 198.835 ;
        RECT 101.440 198.755 102.115 198.915 ;
        RECT 99.420 198.325 100.220 198.495 ;
        RECT 99.540 197.775 99.870 198.155 ;
        RECT 100.050 198.035 100.220 198.325 ;
        RECT 100.810 198.285 100.980 198.665 ;
        RECT 101.150 198.745 102.115 198.755 ;
        RECT 102.305 199.575 102.565 199.965 ;
        RECT 102.775 199.865 103.105 200.325 ;
        RECT 103.980 199.935 104.835 200.105 ;
        RECT 105.040 199.935 105.535 200.105 ;
        RECT 105.705 199.965 106.035 200.325 ;
        RECT 102.305 198.885 102.475 199.575 ;
        RECT 102.645 199.225 102.815 199.405 ;
        RECT 102.985 199.395 103.775 199.645 ;
        RECT 103.980 199.225 104.150 199.935 ;
        RECT 104.320 199.425 104.675 199.645 ;
        RECT 102.645 199.055 104.335 199.225 ;
        RECT 101.150 198.455 101.610 198.745 ;
        RECT 102.305 198.715 103.805 198.885 ;
        RECT 102.305 198.575 102.475 198.715 ;
        RECT 101.915 198.405 102.475 198.575 ;
        RECT 100.390 197.775 100.640 198.235 ;
        RECT 100.810 197.945 101.680 198.285 ;
        RECT 101.915 197.945 102.085 198.405 ;
        RECT 102.920 198.375 103.995 198.545 ;
        RECT 102.255 197.775 102.625 198.235 ;
        RECT 102.920 198.035 103.090 198.375 ;
        RECT 103.260 197.775 103.590 198.205 ;
        RECT 103.825 198.035 103.995 198.375 ;
        RECT 104.165 198.275 104.335 199.055 ;
        RECT 104.505 198.835 104.675 199.425 ;
        RECT 104.845 199.025 105.195 199.645 ;
        RECT 104.505 198.445 104.970 198.835 ;
        RECT 105.365 198.575 105.535 199.935 ;
        RECT 105.705 198.745 106.165 199.795 ;
        RECT 105.140 198.405 105.535 198.575 ;
        RECT 105.140 198.275 105.310 198.405 ;
        RECT 104.165 197.945 104.845 198.275 ;
        RECT 105.060 197.945 105.310 198.275 ;
        RECT 105.480 197.775 105.730 198.235 ;
        RECT 105.900 197.960 106.225 198.745 ;
        RECT 106.395 197.945 106.565 200.065 ;
        RECT 106.735 199.945 107.065 200.325 ;
        RECT 107.235 199.775 107.490 200.065 ;
        RECT 106.740 199.605 107.490 199.775 ;
        RECT 107.665 199.650 107.925 200.155 ;
        RECT 108.105 199.945 108.435 200.325 ;
        RECT 108.615 199.775 108.785 200.155 ;
        RECT 106.740 198.615 106.970 199.605 ;
        RECT 107.140 198.785 107.490 199.435 ;
        RECT 107.665 198.850 107.835 199.650 ;
        RECT 108.120 199.605 108.785 199.775 ;
        RECT 108.120 199.350 108.290 199.605 ;
        RECT 109.085 199.505 109.315 200.325 ;
        RECT 109.485 199.525 109.815 200.155 ;
        RECT 108.005 199.020 108.290 199.350 ;
        RECT 108.525 199.055 108.855 199.425 ;
        RECT 109.065 199.085 109.395 199.335 ;
        RECT 108.120 198.875 108.290 199.020 ;
        RECT 109.565 198.925 109.815 199.525 ;
        RECT 109.985 199.505 110.195 200.325 ;
        RECT 110.885 199.555 114.395 200.325 ;
        RECT 114.565 199.600 114.855 200.325 ;
        RECT 115.490 199.780 120.835 200.325 ;
        RECT 121.010 199.780 126.355 200.325 ;
        RECT 106.740 198.445 107.490 198.615 ;
        RECT 106.735 197.775 107.065 198.275 ;
        RECT 107.235 197.945 107.490 198.445 ;
        RECT 107.665 197.945 107.935 198.850 ;
        RECT 108.120 198.705 108.785 198.875 ;
        RECT 108.105 197.775 108.435 198.535 ;
        RECT 108.615 197.945 108.785 198.705 ;
        RECT 109.085 197.775 109.315 198.915 ;
        RECT 109.485 197.945 109.815 198.925 ;
        RECT 109.985 197.775 110.195 198.915 ;
        RECT 110.885 198.865 112.575 199.385 ;
        RECT 112.745 199.035 114.395 199.555 ;
        RECT 110.885 197.775 114.395 198.865 ;
        RECT 114.565 197.775 114.855 198.940 ;
        RECT 117.080 198.210 117.430 199.460 ;
        RECT 118.910 198.950 119.250 199.780 ;
        RECT 122.600 198.210 122.950 199.460 ;
        RECT 124.430 198.950 124.770 199.780 ;
        RECT 126.525 199.575 127.735 200.325 ;
        RECT 126.525 198.865 127.045 199.405 ;
        RECT 127.215 199.035 127.735 199.575 ;
        RECT 115.490 197.775 120.835 198.210 ;
        RECT 121.010 197.775 126.355 198.210 ;
        RECT 126.525 197.775 127.735 198.865 ;
        RECT 14.660 197.605 127.820 197.775 ;
        RECT 14.745 196.515 15.955 197.605 ;
        RECT 14.745 195.805 15.265 196.345 ;
        RECT 15.435 195.975 15.955 196.515 ;
        RECT 16.125 196.515 18.715 197.605 ;
        RECT 18.890 197.170 24.235 197.605 ;
        RECT 16.125 195.995 17.335 196.515 ;
        RECT 17.505 195.825 18.715 196.345 ;
        RECT 20.480 195.920 20.830 197.170 ;
        RECT 24.405 196.440 24.695 197.605 ;
        RECT 25.325 196.515 27.915 197.605 ;
        RECT 28.090 197.170 33.435 197.605 ;
        RECT 33.610 197.170 38.955 197.605 ;
        RECT 39.130 197.170 44.475 197.605 ;
        RECT 44.650 197.170 49.995 197.605 ;
        RECT 14.745 195.055 15.955 195.805 ;
        RECT 16.125 195.055 18.715 195.825 ;
        RECT 22.310 195.600 22.650 196.430 ;
        RECT 25.325 195.995 26.535 196.515 ;
        RECT 26.705 195.825 27.915 196.345 ;
        RECT 29.680 195.920 30.030 197.170 ;
        RECT 18.890 195.055 24.235 195.600 ;
        RECT 24.405 195.055 24.695 195.780 ;
        RECT 25.325 195.055 27.915 195.825 ;
        RECT 31.510 195.600 31.850 196.430 ;
        RECT 35.200 195.920 35.550 197.170 ;
        RECT 37.030 195.600 37.370 196.430 ;
        RECT 40.720 195.920 41.070 197.170 ;
        RECT 42.550 195.600 42.890 196.430 ;
        RECT 46.240 195.920 46.590 197.170 ;
        RECT 50.165 196.440 50.455 197.605 ;
        RECT 50.630 197.170 55.975 197.605 ;
        RECT 56.150 197.170 61.495 197.605 ;
        RECT 48.070 195.600 48.410 196.430 ;
        RECT 52.220 195.920 52.570 197.170 ;
        RECT 28.090 195.055 33.435 195.600 ;
        RECT 33.610 195.055 38.955 195.600 ;
        RECT 39.130 195.055 44.475 195.600 ;
        RECT 44.650 195.055 49.995 195.600 ;
        RECT 50.165 195.055 50.455 195.780 ;
        RECT 54.050 195.600 54.390 196.430 ;
        RECT 57.740 195.920 58.090 197.170 ;
        RECT 61.725 196.465 61.935 197.605 ;
        RECT 62.105 196.455 62.435 197.435 ;
        RECT 62.605 196.465 62.835 197.605 ;
        RECT 63.045 196.515 64.715 197.605 ;
        RECT 64.885 197.050 65.490 197.605 ;
        RECT 65.665 197.095 66.145 197.435 ;
        RECT 66.315 197.060 66.570 197.605 ;
        RECT 64.885 196.950 65.500 197.050 ;
        RECT 65.315 196.925 65.500 196.950 ;
        RECT 59.570 195.600 59.910 196.430 ;
        RECT 50.630 195.055 55.975 195.600 ;
        RECT 56.150 195.055 61.495 195.600 ;
        RECT 61.725 195.055 61.935 195.875 ;
        RECT 62.105 195.855 62.355 196.455 ;
        RECT 62.525 196.045 62.855 196.295 ;
        RECT 63.045 195.995 63.795 196.515 ;
        RECT 62.105 195.225 62.435 195.855 ;
        RECT 62.605 195.055 62.835 195.875 ;
        RECT 63.965 195.825 64.715 196.345 ;
        RECT 64.885 196.330 65.145 196.780 ;
        RECT 65.315 196.680 65.645 196.925 ;
        RECT 65.815 196.605 66.570 196.855 ;
        RECT 66.740 196.735 67.015 197.435 ;
        RECT 65.800 196.570 66.570 196.605 ;
        RECT 65.785 196.560 66.570 196.570 ;
        RECT 65.780 196.545 66.675 196.560 ;
        RECT 65.760 196.530 66.675 196.545 ;
        RECT 65.740 196.520 66.675 196.530 ;
        RECT 65.715 196.510 66.675 196.520 ;
        RECT 65.645 196.480 66.675 196.510 ;
        RECT 65.625 196.450 66.675 196.480 ;
        RECT 65.605 196.420 66.675 196.450 ;
        RECT 65.575 196.395 66.675 196.420 ;
        RECT 65.540 196.360 66.675 196.395 ;
        RECT 65.510 196.355 66.675 196.360 ;
        RECT 65.510 196.350 65.900 196.355 ;
        RECT 65.510 196.340 65.875 196.350 ;
        RECT 65.510 196.335 65.860 196.340 ;
        RECT 65.510 196.330 65.845 196.335 ;
        RECT 64.885 196.325 65.845 196.330 ;
        RECT 64.885 196.315 65.835 196.325 ;
        RECT 64.885 196.310 65.825 196.315 ;
        RECT 64.885 196.300 65.815 196.310 ;
        RECT 64.885 196.290 65.810 196.300 ;
        RECT 64.885 196.285 65.805 196.290 ;
        RECT 64.885 196.270 65.795 196.285 ;
        RECT 64.885 196.255 65.790 196.270 ;
        RECT 64.885 196.230 65.780 196.255 ;
        RECT 64.885 196.160 65.775 196.230 ;
        RECT 63.045 195.055 64.715 195.825 ;
        RECT 64.885 195.605 65.435 195.990 ;
        RECT 65.605 195.435 65.775 196.160 ;
        RECT 64.885 195.265 65.775 195.435 ;
        RECT 65.945 195.760 66.275 196.185 ;
        RECT 66.445 195.960 66.675 196.355 ;
        RECT 65.945 195.275 66.165 195.760 ;
        RECT 66.845 195.705 67.015 196.735 ;
        RECT 66.335 195.055 66.585 195.595 ;
        RECT 66.755 195.225 67.015 195.705 ;
        RECT 67.195 196.545 67.525 197.395 ;
        RECT 67.195 195.780 67.385 196.545 ;
        RECT 67.695 196.465 67.945 197.605 ;
        RECT 68.135 196.965 68.385 197.385 ;
        RECT 68.615 197.135 68.945 197.605 ;
        RECT 69.175 196.965 69.425 197.385 ;
        RECT 68.135 196.795 69.425 196.965 ;
        RECT 69.605 196.965 69.935 197.395 ;
        RECT 69.605 196.795 70.060 196.965 ;
        RECT 68.125 196.295 68.340 196.625 ;
        RECT 67.555 195.965 67.865 196.295 ;
        RECT 68.035 195.965 68.340 196.295 ;
        RECT 68.515 195.965 68.800 196.625 ;
        RECT 68.995 195.965 69.260 196.625 ;
        RECT 69.475 195.965 69.720 196.625 ;
        RECT 67.695 195.795 67.865 195.965 ;
        RECT 69.890 195.795 70.060 196.795 ;
        RECT 67.195 195.270 67.525 195.780 ;
        RECT 67.695 195.625 70.060 195.795 ;
        RECT 70.405 196.465 70.680 197.435 ;
        RECT 70.890 196.805 71.170 197.605 ;
        RECT 71.340 197.095 72.955 197.425 ;
        RECT 71.340 196.755 72.515 196.925 ;
        RECT 71.340 196.635 71.510 196.755 ;
        RECT 70.850 196.465 71.510 196.635 ;
        RECT 70.405 195.730 70.575 196.465 ;
        RECT 70.850 196.295 71.020 196.465 ;
        RECT 71.770 196.295 72.015 196.585 ;
        RECT 72.185 196.465 72.515 196.755 ;
        RECT 72.775 196.295 72.945 196.855 ;
        RECT 73.195 196.465 73.455 197.605 ;
        RECT 73.660 196.815 74.195 197.435 ;
        RECT 70.745 195.965 71.020 196.295 ;
        RECT 71.190 195.965 72.015 196.295 ;
        RECT 72.230 195.965 72.945 196.295 ;
        RECT 73.115 196.045 73.450 196.295 ;
        RECT 70.850 195.795 71.020 195.965 ;
        RECT 72.695 195.875 72.945 195.965 ;
        RECT 67.695 195.055 68.025 195.455 ;
        RECT 69.075 195.285 69.405 195.625 ;
        RECT 69.575 195.055 69.905 195.455 ;
        RECT 70.405 195.385 70.680 195.730 ;
        RECT 70.850 195.625 72.515 195.795 ;
        RECT 70.870 195.055 71.245 195.455 ;
        RECT 71.415 195.275 71.585 195.625 ;
        RECT 71.755 195.055 72.085 195.455 ;
        RECT 72.255 195.225 72.515 195.625 ;
        RECT 72.695 195.455 73.025 195.875 ;
        RECT 73.195 195.055 73.455 195.875 ;
        RECT 73.660 195.795 73.975 196.815 ;
        RECT 74.365 196.805 74.695 197.605 ;
        RECT 75.180 196.635 75.570 196.810 ;
        RECT 74.145 196.465 75.570 196.635 ;
        RECT 74.145 195.965 74.315 196.465 ;
        RECT 73.660 195.225 74.275 195.795 ;
        RECT 74.565 195.735 74.830 196.295 ;
        RECT 75.000 195.565 75.170 196.465 ;
        RECT 75.925 196.440 76.215 197.605 ;
        RECT 76.845 197.095 77.145 197.605 ;
        RECT 77.315 196.925 77.645 197.435 ;
        RECT 77.815 197.095 78.445 197.605 ;
        RECT 79.025 197.095 79.405 197.265 ;
        RECT 79.575 197.095 79.875 197.605 ;
        RECT 79.235 196.925 79.405 197.095 ;
        RECT 76.845 196.755 79.065 196.925 ;
        RECT 75.340 195.735 75.695 196.295 ;
        RECT 76.845 195.795 77.015 196.755 ;
        RECT 77.185 196.415 78.725 196.585 ;
        RECT 77.185 195.965 77.430 196.415 ;
        RECT 77.690 196.045 78.385 196.245 ;
        RECT 78.555 196.215 78.725 196.415 ;
        RECT 78.895 196.555 79.065 196.755 ;
        RECT 79.235 196.725 79.895 196.925 ;
        RECT 78.895 196.385 79.555 196.555 ;
        RECT 78.555 196.045 79.155 196.215 ;
        RECT 79.385 195.965 79.555 196.385 ;
        RECT 74.445 195.055 74.660 195.565 ;
        RECT 74.890 195.235 75.170 195.565 ;
        RECT 75.350 195.055 75.590 195.565 ;
        RECT 75.925 195.055 76.215 195.780 ;
        RECT 76.845 195.250 77.310 195.795 ;
        RECT 77.815 195.055 77.985 195.875 ;
        RECT 78.155 195.795 79.065 195.875 ;
        RECT 79.725 195.795 79.895 196.725 ;
        RECT 80.985 196.515 84.495 197.605 ;
        RECT 84.670 197.170 90.015 197.605 ;
        RECT 80.985 195.995 82.675 196.515 ;
        RECT 82.845 195.825 84.495 196.345 ;
        RECT 86.260 195.920 86.610 197.170 ;
        RECT 90.185 196.845 90.700 197.255 ;
        RECT 90.935 196.845 91.105 197.605 ;
        RECT 91.275 197.265 93.305 197.435 ;
        RECT 78.155 195.705 79.405 195.795 ;
        RECT 78.155 195.225 78.485 195.705 ;
        RECT 78.895 195.625 79.405 195.705 ;
        RECT 78.655 195.055 79.005 195.445 ;
        RECT 79.175 195.225 79.405 195.625 ;
        RECT 79.575 195.315 79.895 195.795 ;
        RECT 80.985 195.055 84.495 195.825 ;
        RECT 88.090 195.600 88.430 196.430 ;
        RECT 90.185 196.035 90.525 196.845 ;
        RECT 91.275 196.600 91.445 197.265 ;
        RECT 91.840 196.925 92.965 197.095 ;
        RECT 90.695 196.410 91.445 196.600 ;
        RECT 91.615 196.585 92.625 196.755 ;
        RECT 90.185 195.865 91.415 196.035 ;
        RECT 84.670 195.055 90.015 195.600 ;
        RECT 90.460 195.260 90.705 195.865 ;
        RECT 90.925 195.055 91.435 195.590 ;
        RECT 91.615 195.225 91.805 196.585 ;
        RECT 91.975 195.565 92.250 196.385 ;
        RECT 92.455 195.785 92.625 196.585 ;
        RECT 92.795 195.795 92.965 196.925 ;
        RECT 93.135 196.295 93.305 197.265 ;
        RECT 93.475 196.465 93.645 197.605 ;
        RECT 93.815 196.465 94.150 197.435 ;
        RECT 94.415 196.675 94.585 197.435 ;
        RECT 94.765 196.845 95.095 197.605 ;
        RECT 94.415 196.505 95.080 196.675 ;
        RECT 95.265 196.530 95.535 197.435 ;
        RECT 93.135 195.965 93.330 196.295 ;
        RECT 93.555 195.965 93.810 196.295 ;
        RECT 93.555 195.795 93.725 195.965 ;
        RECT 93.980 195.795 94.150 196.465 ;
        RECT 94.910 196.360 95.080 196.505 ;
        RECT 94.345 195.955 94.675 196.325 ;
        RECT 94.910 196.030 95.195 196.360 ;
        RECT 92.795 195.625 93.725 195.795 ;
        RECT 92.795 195.590 92.970 195.625 ;
        RECT 91.975 195.395 92.255 195.565 ;
        RECT 91.975 195.225 92.250 195.395 ;
        RECT 92.440 195.225 92.970 195.590 ;
        RECT 93.395 195.055 93.725 195.455 ;
        RECT 93.895 195.225 94.150 195.795 ;
        RECT 94.910 195.775 95.080 196.030 ;
        RECT 94.415 195.605 95.080 195.775 ;
        RECT 95.365 195.730 95.535 196.530 ;
        RECT 95.705 196.515 97.375 197.605 ;
        RECT 97.545 196.845 98.060 197.255 ;
        RECT 98.295 196.845 98.465 197.605 ;
        RECT 98.635 197.265 100.665 197.435 ;
        RECT 95.705 195.995 96.455 196.515 ;
        RECT 96.625 195.825 97.375 196.345 ;
        RECT 97.545 196.035 97.885 196.845 ;
        RECT 98.635 196.600 98.805 197.265 ;
        RECT 99.200 196.925 100.325 197.095 ;
        RECT 98.055 196.410 98.805 196.600 ;
        RECT 98.975 196.585 99.985 196.755 ;
        RECT 97.545 195.865 98.775 196.035 ;
        RECT 94.415 195.225 94.585 195.605 ;
        RECT 94.765 195.055 95.095 195.435 ;
        RECT 95.275 195.225 95.535 195.730 ;
        RECT 95.705 195.055 97.375 195.825 ;
        RECT 97.820 195.260 98.065 195.865 ;
        RECT 98.285 195.055 98.795 195.590 ;
        RECT 98.975 195.225 99.165 196.585 ;
        RECT 99.335 196.245 99.610 196.385 ;
        RECT 99.335 196.075 99.615 196.245 ;
        RECT 99.335 195.225 99.610 196.075 ;
        RECT 99.815 195.785 99.985 196.585 ;
        RECT 100.155 195.795 100.325 196.925 ;
        RECT 100.495 196.295 100.665 197.265 ;
        RECT 100.835 196.465 101.005 197.605 ;
        RECT 101.175 196.465 101.510 197.435 ;
        RECT 100.495 195.965 100.690 196.295 ;
        RECT 100.915 195.965 101.170 196.295 ;
        RECT 100.915 195.795 101.085 195.965 ;
        RECT 101.340 195.795 101.510 196.465 ;
        RECT 101.685 196.440 101.975 197.605 ;
        RECT 102.605 196.515 104.275 197.605 ;
        RECT 104.445 196.845 104.960 197.255 ;
        RECT 105.195 196.845 105.365 197.605 ;
        RECT 105.535 197.265 107.565 197.435 ;
        RECT 102.605 195.995 103.355 196.515 ;
        RECT 103.525 195.825 104.275 196.345 ;
        RECT 104.445 196.035 104.785 196.845 ;
        RECT 105.535 196.600 105.705 197.265 ;
        RECT 106.100 196.925 107.225 197.095 ;
        RECT 104.955 196.410 105.705 196.600 ;
        RECT 105.875 196.585 106.885 196.755 ;
        RECT 104.445 195.865 105.675 196.035 ;
        RECT 100.155 195.625 101.085 195.795 ;
        RECT 100.155 195.590 100.330 195.625 ;
        RECT 99.800 195.225 100.330 195.590 ;
        RECT 100.755 195.055 101.085 195.455 ;
        RECT 101.255 195.225 101.510 195.795 ;
        RECT 101.685 195.055 101.975 195.780 ;
        RECT 102.605 195.055 104.275 195.825 ;
        RECT 104.720 195.260 104.965 195.865 ;
        RECT 105.185 195.055 105.695 195.590 ;
        RECT 105.875 195.225 106.065 196.585 ;
        RECT 106.235 195.905 106.510 196.385 ;
        RECT 106.235 195.735 106.515 195.905 ;
        RECT 106.715 195.785 106.885 196.585 ;
        RECT 107.055 195.795 107.225 196.925 ;
        RECT 107.395 196.295 107.565 197.265 ;
        RECT 107.735 196.465 107.905 197.605 ;
        RECT 108.075 196.465 108.410 197.435 ;
        RECT 109.595 196.675 109.765 197.435 ;
        RECT 109.945 196.845 110.275 197.605 ;
        RECT 109.595 196.505 110.260 196.675 ;
        RECT 110.445 196.530 110.715 197.435 ;
        RECT 107.395 195.965 107.590 196.295 ;
        RECT 107.815 195.965 108.070 196.295 ;
        RECT 107.815 195.795 107.985 195.965 ;
        RECT 108.240 195.795 108.410 196.465 ;
        RECT 110.090 196.360 110.260 196.505 ;
        RECT 109.525 195.955 109.855 196.325 ;
        RECT 110.090 196.030 110.375 196.360 ;
        RECT 106.235 195.225 106.510 195.735 ;
        RECT 107.055 195.625 107.985 195.795 ;
        RECT 107.055 195.590 107.230 195.625 ;
        RECT 106.700 195.225 107.230 195.590 ;
        RECT 107.655 195.055 107.985 195.455 ;
        RECT 108.155 195.225 108.410 195.795 ;
        RECT 110.090 195.775 110.260 196.030 ;
        RECT 109.595 195.605 110.260 195.775 ;
        RECT 110.545 195.730 110.715 196.530 ;
        RECT 111.805 196.515 115.315 197.605 ;
        RECT 115.490 197.170 120.835 197.605 ;
        RECT 121.010 197.170 126.355 197.605 ;
        RECT 111.805 195.995 113.495 196.515 ;
        RECT 113.665 195.825 115.315 196.345 ;
        RECT 117.080 195.920 117.430 197.170 ;
        RECT 109.595 195.225 109.765 195.605 ;
        RECT 109.945 195.055 110.275 195.435 ;
        RECT 110.455 195.225 110.715 195.730 ;
        RECT 111.805 195.055 115.315 195.825 ;
        RECT 118.910 195.600 119.250 196.430 ;
        RECT 122.600 195.920 122.950 197.170 ;
        RECT 126.525 196.515 127.735 197.605 ;
        RECT 124.430 195.600 124.770 196.430 ;
        RECT 126.525 195.975 127.045 196.515 ;
        RECT 127.215 195.805 127.735 196.345 ;
        RECT 115.490 195.055 120.835 195.600 ;
        RECT 121.010 195.055 126.355 195.600 ;
        RECT 126.525 195.055 127.735 195.805 ;
        RECT 14.660 194.885 127.820 195.055 ;
        RECT 14.745 194.135 15.955 194.885 ;
        RECT 14.745 193.595 15.265 194.135 ;
        RECT 17.045 194.115 20.555 194.885 ;
        RECT 20.730 194.340 26.075 194.885 ;
        RECT 26.250 194.340 31.595 194.885 ;
        RECT 31.770 194.340 37.115 194.885 ;
        RECT 15.435 193.425 15.955 193.965 ;
        RECT 14.745 192.335 15.955 193.425 ;
        RECT 17.045 193.425 18.735 193.945 ;
        RECT 18.905 193.595 20.555 194.115 ;
        RECT 17.045 192.335 20.555 193.425 ;
        RECT 22.320 192.770 22.670 194.020 ;
        RECT 24.150 193.510 24.490 194.340 ;
        RECT 27.840 192.770 28.190 194.020 ;
        RECT 29.670 193.510 30.010 194.340 ;
        RECT 33.360 192.770 33.710 194.020 ;
        RECT 35.190 193.510 35.530 194.340 ;
        RECT 37.285 194.160 37.575 194.885 ;
        RECT 37.750 194.340 43.095 194.885 ;
        RECT 43.270 194.340 48.615 194.885 ;
        RECT 20.730 192.335 26.075 192.770 ;
        RECT 26.250 192.335 31.595 192.770 ;
        RECT 31.770 192.335 37.115 192.770 ;
        RECT 37.285 192.335 37.575 193.500 ;
        RECT 39.340 192.770 39.690 194.020 ;
        RECT 41.170 193.510 41.510 194.340 ;
        RECT 44.860 192.770 45.210 194.020 ;
        RECT 46.690 193.510 47.030 194.340 ;
        RECT 48.845 194.065 49.055 194.885 ;
        RECT 49.225 194.085 49.555 194.715 ;
        RECT 49.225 193.485 49.475 194.085 ;
        RECT 49.725 194.065 49.955 194.885 ;
        RECT 50.165 194.115 51.835 194.885 ;
        RECT 49.645 193.645 49.975 193.895 ;
        RECT 37.750 192.335 43.095 192.770 ;
        RECT 43.270 192.335 48.615 192.770 ;
        RECT 48.845 192.335 49.055 193.475 ;
        RECT 49.225 192.505 49.555 193.485 ;
        RECT 49.725 192.335 49.955 193.475 ;
        RECT 50.165 193.425 50.915 193.945 ;
        RECT 51.085 193.595 51.835 194.115 ;
        RECT 52.045 194.065 52.275 194.885 ;
        RECT 52.445 194.085 52.775 194.715 ;
        RECT 52.025 193.645 52.355 193.895 ;
        RECT 52.525 193.485 52.775 194.085 ;
        RECT 52.945 194.065 53.155 194.885 ;
        RECT 53.390 194.335 53.645 194.625 ;
        RECT 53.815 194.505 54.145 194.885 ;
        RECT 53.390 194.165 54.140 194.335 ;
        RECT 50.165 192.335 51.835 193.425 ;
        RECT 52.045 192.335 52.275 193.475 ;
        RECT 52.445 192.505 52.775 193.485 ;
        RECT 52.945 192.335 53.155 193.475 ;
        RECT 53.390 193.345 53.740 193.995 ;
        RECT 53.910 193.175 54.140 194.165 ;
        RECT 53.390 193.005 54.140 193.175 ;
        RECT 53.390 192.505 53.645 193.005 ;
        RECT 53.815 192.335 54.145 192.835 ;
        RECT 54.315 192.505 54.485 194.625 ;
        RECT 54.845 194.525 55.175 194.885 ;
        RECT 55.345 194.495 55.840 194.665 ;
        RECT 56.045 194.495 56.900 194.665 ;
        RECT 54.715 193.305 55.175 194.355 ;
        RECT 54.655 192.520 54.980 193.305 ;
        RECT 55.345 193.135 55.515 194.495 ;
        RECT 55.685 193.585 56.035 194.205 ;
        RECT 56.205 193.985 56.560 194.205 ;
        RECT 56.205 193.395 56.375 193.985 ;
        RECT 56.730 193.785 56.900 194.495 ;
        RECT 57.775 194.425 58.105 194.885 ;
        RECT 58.315 194.525 58.665 194.695 ;
        RECT 57.105 193.955 57.895 194.205 ;
        RECT 58.315 194.135 58.575 194.525 ;
        RECT 58.885 194.435 59.835 194.715 ;
        RECT 60.005 194.445 60.195 194.885 ;
        RECT 60.365 194.505 61.435 194.675 ;
        RECT 58.065 193.785 58.235 193.965 ;
        RECT 55.345 192.965 55.740 193.135 ;
        RECT 55.910 193.005 56.375 193.395 ;
        RECT 56.545 193.615 58.235 193.785 ;
        RECT 55.570 192.835 55.740 192.965 ;
        RECT 56.545 192.835 56.715 193.615 ;
        RECT 58.405 193.445 58.575 194.135 ;
        RECT 57.075 193.275 58.575 193.445 ;
        RECT 58.765 193.475 58.975 194.265 ;
        RECT 59.145 193.645 59.495 194.265 ;
        RECT 59.665 193.655 59.835 194.435 ;
        RECT 60.365 194.275 60.535 194.505 ;
        RECT 60.005 194.105 60.535 194.275 ;
        RECT 60.005 193.825 60.225 194.105 ;
        RECT 60.705 193.935 60.945 194.335 ;
        RECT 59.665 193.485 60.070 193.655 ;
        RECT 60.405 193.565 60.945 193.935 ;
        RECT 61.115 194.150 61.435 194.505 ;
        RECT 61.680 194.425 61.985 194.885 ;
        RECT 62.155 194.175 62.405 194.705 ;
        RECT 61.115 193.975 61.440 194.150 ;
        RECT 61.115 193.675 62.030 193.975 ;
        RECT 61.290 193.645 62.030 193.675 ;
        RECT 58.765 193.315 59.440 193.475 ;
        RECT 59.900 193.395 60.070 193.485 ;
        RECT 58.765 193.305 59.730 193.315 ;
        RECT 58.405 193.135 58.575 193.275 ;
        RECT 55.150 192.335 55.400 192.795 ;
        RECT 55.570 192.505 55.820 192.835 ;
        RECT 56.035 192.505 56.715 192.835 ;
        RECT 56.885 192.935 57.960 193.105 ;
        RECT 58.405 192.965 58.965 193.135 ;
        RECT 59.270 193.015 59.730 193.305 ;
        RECT 59.900 193.225 61.120 193.395 ;
        RECT 56.885 192.595 57.055 192.935 ;
        RECT 57.290 192.335 57.620 192.765 ;
        RECT 57.790 192.595 57.960 192.935 ;
        RECT 58.255 192.335 58.625 192.795 ;
        RECT 58.795 192.505 58.965 192.965 ;
        RECT 59.900 192.845 60.070 193.225 ;
        RECT 61.290 193.055 61.460 193.645 ;
        RECT 62.200 193.525 62.405 194.175 ;
        RECT 62.575 194.130 62.825 194.885 ;
        RECT 63.045 194.160 63.335 194.885 ;
        RECT 63.965 194.115 65.635 194.885 ;
        RECT 59.200 192.505 60.070 192.845 ;
        RECT 60.660 192.885 61.460 193.055 ;
        RECT 60.240 192.335 60.490 192.795 ;
        RECT 60.660 192.595 60.830 192.885 ;
        RECT 61.010 192.335 61.340 192.715 ;
        RECT 61.680 192.335 61.985 193.475 ;
        RECT 62.155 192.645 62.405 193.525 ;
        RECT 62.575 192.335 62.825 193.475 ;
        RECT 63.045 192.335 63.335 193.500 ;
        RECT 63.965 193.425 64.715 193.945 ;
        RECT 64.885 193.595 65.635 194.115 ;
        RECT 65.805 194.145 66.125 194.625 ;
        RECT 66.295 194.315 66.525 194.715 ;
        RECT 66.695 194.495 67.045 194.885 ;
        RECT 66.295 194.235 66.805 194.315 ;
        RECT 67.215 194.235 67.545 194.715 ;
        RECT 66.295 194.145 67.545 194.235 ;
        RECT 63.965 192.335 65.635 193.425 ;
        RECT 65.805 193.215 65.975 194.145 ;
        RECT 66.635 194.065 67.545 194.145 ;
        RECT 67.715 194.065 67.885 194.885 ;
        RECT 68.390 194.145 68.855 194.690 ;
        RECT 66.145 193.555 66.315 193.975 ;
        RECT 66.545 193.725 67.145 193.895 ;
        RECT 66.145 193.385 66.805 193.555 ;
        RECT 65.805 193.015 66.465 193.215 ;
        RECT 66.635 193.185 66.805 193.385 ;
        RECT 66.975 193.525 67.145 193.725 ;
        RECT 67.315 193.695 68.010 193.895 ;
        RECT 68.270 193.525 68.515 193.975 ;
        RECT 66.975 193.355 68.515 193.525 ;
        RECT 68.685 193.185 68.855 194.145 ;
        RECT 69.025 194.065 69.285 194.885 ;
        RECT 69.455 194.065 69.785 194.485 ;
        RECT 69.965 194.315 70.225 194.715 ;
        RECT 70.395 194.485 70.725 194.885 ;
        RECT 70.895 194.315 71.065 194.665 ;
        RECT 71.235 194.485 71.610 194.885 ;
        RECT 69.965 194.145 71.630 194.315 ;
        RECT 71.800 194.210 72.075 194.555 ;
        RECT 69.535 193.975 69.785 194.065 ;
        RECT 71.460 193.975 71.630 194.145 ;
        RECT 69.030 193.645 69.365 193.895 ;
        RECT 69.535 193.645 70.250 193.975 ;
        RECT 70.465 193.645 71.290 193.975 ;
        RECT 71.460 193.645 71.735 193.975 ;
        RECT 66.635 193.015 68.855 193.185 ;
        RECT 66.295 192.845 66.465 193.015 ;
        RECT 65.825 192.335 66.125 192.845 ;
        RECT 66.295 192.675 66.675 192.845 ;
        RECT 67.255 192.335 67.885 192.845 ;
        RECT 68.055 192.505 68.385 193.015 ;
        RECT 68.555 192.335 68.855 192.845 ;
        RECT 69.025 192.335 69.285 193.475 ;
        RECT 69.535 193.085 69.705 193.645 ;
        RECT 69.965 193.185 70.295 193.475 ;
        RECT 70.465 193.355 70.710 193.645 ;
        RECT 71.460 193.475 71.630 193.645 ;
        RECT 71.905 193.475 72.075 194.210 ;
        RECT 72.705 194.115 74.375 194.885 ;
        RECT 70.970 193.305 71.630 193.475 ;
        RECT 70.970 193.185 71.140 193.305 ;
        RECT 69.965 193.015 71.140 193.185 ;
        RECT 69.525 192.515 71.140 192.845 ;
        RECT 71.310 192.335 71.590 193.135 ;
        RECT 71.800 192.505 72.075 193.475 ;
        RECT 72.705 193.425 73.455 193.945 ;
        RECT 73.625 193.595 74.375 194.115 ;
        RECT 74.545 194.085 74.855 194.885 ;
        RECT 75.060 194.085 75.755 194.715 ;
        RECT 76.385 194.115 78.975 194.885 ;
        RECT 79.150 194.340 84.495 194.885 ;
        RECT 74.555 193.645 74.890 193.915 ;
        RECT 75.060 193.485 75.230 194.085 ;
        RECT 75.400 193.645 75.735 193.895 ;
        RECT 72.705 192.335 74.375 193.425 ;
        RECT 74.545 192.335 74.825 193.475 ;
        RECT 74.995 192.505 75.325 193.485 ;
        RECT 75.495 192.335 75.755 193.475 ;
        RECT 76.385 193.425 77.595 193.945 ;
        RECT 77.765 193.595 78.975 194.115 ;
        RECT 76.385 192.335 78.975 193.425 ;
        RECT 80.740 192.770 81.090 194.020 ;
        RECT 82.570 193.510 82.910 194.340 ;
        RECT 84.940 194.075 85.185 194.680 ;
        RECT 85.405 194.350 85.915 194.885 ;
        RECT 84.665 193.905 85.895 194.075 ;
        RECT 84.665 193.095 85.005 193.905 ;
        RECT 85.175 193.340 85.925 193.530 ;
        RECT 79.150 192.335 84.495 192.770 ;
        RECT 84.665 192.685 85.180 193.095 ;
        RECT 85.415 192.335 85.585 193.095 ;
        RECT 85.755 192.675 85.925 193.340 ;
        RECT 86.095 193.355 86.285 194.715 ;
        RECT 86.455 193.865 86.730 194.715 ;
        RECT 86.920 194.350 87.450 194.715 ;
        RECT 87.875 194.485 88.205 194.885 ;
        RECT 87.275 194.315 87.450 194.350 ;
        RECT 86.455 193.695 86.735 193.865 ;
        RECT 86.455 193.555 86.730 193.695 ;
        RECT 86.935 193.355 87.105 194.155 ;
        RECT 86.095 193.185 87.105 193.355 ;
        RECT 87.275 194.145 88.205 194.315 ;
        RECT 88.375 194.145 88.630 194.715 ;
        RECT 88.805 194.160 89.095 194.885 ;
        RECT 89.815 194.335 89.985 194.715 ;
        RECT 90.165 194.505 90.495 194.885 ;
        RECT 89.815 194.165 90.480 194.335 ;
        RECT 90.675 194.210 90.935 194.715 ;
        RECT 87.275 193.015 87.445 194.145 ;
        RECT 88.035 193.975 88.205 194.145 ;
        RECT 86.320 192.845 87.445 193.015 ;
        RECT 87.615 193.645 87.810 193.975 ;
        RECT 88.035 193.645 88.290 193.975 ;
        RECT 87.615 192.675 87.785 193.645 ;
        RECT 88.460 193.475 88.630 194.145 ;
        RECT 89.745 193.615 90.075 193.985 ;
        RECT 90.310 193.910 90.480 194.165 ;
        RECT 90.310 193.580 90.595 193.910 ;
        RECT 85.755 192.505 87.785 192.675 ;
        RECT 87.955 192.335 88.125 193.475 ;
        RECT 88.295 192.505 88.630 193.475 ;
        RECT 88.805 192.335 89.095 193.500 ;
        RECT 90.310 193.435 90.480 193.580 ;
        RECT 89.815 193.265 90.480 193.435 ;
        RECT 90.765 193.410 90.935 194.210 ;
        RECT 91.105 194.135 92.315 194.885 ;
        RECT 92.490 194.340 97.835 194.885 ;
        RECT 98.010 194.340 103.355 194.885 ;
        RECT 89.815 192.505 89.985 193.265 ;
        RECT 90.165 192.335 90.495 193.095 ;
        RECT 90.665 192.505 90.935 193.410 ;
        RECT 91.105 193.425 91.625 193.965 ;
        RECT 91.795 193.595 92.315 194.135 ;
        RECT 91.105 192.335 92.315 193.425 ;
        RECT 94.080 192.770 94.430 194.020 ;
        RECT 95.910 193.510 96.250 194.340 ;
        RECT 99.600 192.770 99.950 194.020 ;
        RECT 101.430 193.510 101.770 194.340 ;
        RECT 103.565 194.065 103.795 194.885 ;
        RECT 103.965 194.085 104.295 194.715 ;
        RECT 103.545 193.645 103.875 193.895 ;
        RECT 104.045 193.485 104.295 194.085 ;
        RECT 104.465 194.065 104.675 194.885 ;
        RECT 105.180 194.075 105.425 194.680 ;
        RECT 105.645 194.350 106.155 194.885 ;
        RECT 92.490 192.335 97.835 192.770 ;
        RECT 98.010 192.335 103.355 192.770 ;
        RECT 103.565 192.335 103.795 193.475 ;
        RECT 103.965 192.505 104.295 193.485 ;
        RECT 104.905 193.905 106.135 194.075 ;
        RECT 104.465 192.335 104.675 193.475 ;
        RECT 104.905 193.095 105.245 193.905 ;
        RECT 105.415 193.340 106.165 193.530 ;
        RECT 104.905 192.685 105.420 193.095 ;
        RECT 105.655 192.335 105.825 193.095 ;
        RECT 105.995 192.675 106.165 193.340 ;
        RECT 106.335 193.355 106.525 194.715 ;
        RECT 106.695 194.205 106.970 194.715 ;
        RECT 107.160 194.350 107.690 194.715 ;
        RECT 108.115 194.485 108.445 194.885 ;
        RECT 107.515 194.315 107.690 194.350 ;
        RECT 106.695 194.035 106.975 194.205 ;
        RECT 106.695 193.555 106.970 194.035 ;
        RECT 107.175 193.355 107.345 194.155 ;
        RECT 106.335 193.185 107.345 193.355 ;
        RECT 107.515 194.145 108.445 194.315 ;
        RECT 108.615 194.145 108.870 194.715 ;
        RECT 109.135 194.335 109.305 194.715 ;
        RECT 109.485 194.505 109.815 194.885 ;
        RECT 109.135 194.165 109.800 194.335 ;
        RECT 109.995 194.210 110.255 194.715 ;
        RECT 107.515 193.015 107.685 194.145 ;
        RECT 108.275 193.975 108.445 194.145 ;
        RECT 106.560 192.845 107.685 193.015 ;
        RECT 107.855 193.645 108.050 193.975 ;
        RECT 108.275 193.645 108.530 193.975 ;
        RECT 107.855 192.675 108.025 193.645 ;
        RECT 108.700 193.475 108.870 194.145 ;
        RECT 109.065 193.615 109.395 193.985 ;
        RECT 109.630 193.910 109.800 194.165 ;
        RECT 105.995 192.505 108.025 192.675 ;
        RECT 108.195 192.335 108.365 193.475 ;
        RECT 108.535 192.505 108.870 193.475 ;
        RECT 109.630 193.580 109.915 193.910 ;
        RECT 109.630 193.435 109.800 193.580 ;
        RECT 109.135 193.265 109.800 193.435 ;
        RECT 110.085 193.410 110.255 194.210 ;
        RECT 110.885 194.115 114.395 194.885 ;
        RECT 114.565 194.160 114.855 194.885 ;
        RECT 115.490 194.340 120.835 194.885 ;
        RECT 121.010 194.340 126.355 194.885 ;
        RECT 109.135 192.505 109.305 193.265 ;
        RECT 109.485 192.335 109.815 193.095 ;
        RECT 109.985 192.505 110.255 193.410 ;
        RECT 110.885 193.425 112.575 193.945 ;
        RECT 112.745 193.595 114.395 194.115 ;
        RECT 110.885 192.335 114.395 193.425 ;
        RECT 114.565 192.335 114.855 193.500 ;
        RECT 117.080 192.770 117.430 194.020 ;
        RECT 118.910 193.510 119.250 194.340 ;
        RECT 122.600 192.770 122.950 194.020 ;
        RECT 124.430 193.510 124.770 194.340 ;
        RECT 126.525 194.135 127.735 194.885 ;
        RECT 126.525 193.425 127.045 193.965 ;
        RECT 127.215 193.595 127.735 194.135 ;
        RECT 115.490 192.335 120.835 192.770 ;
        RECT 121.010 192.335 126.355 192.770 ;
        RECT 126.525 192.335 127.735 193.425 ;
        RECT 14.660 192.165 127.820 192.335 ;
        RECT 14.745 191.075 15.955 192.165 ;
        RECT 14.745 190.365 15.265 190.905 ;
        RECT 15.435 190.535 15.955 191.075 ;
        RECT 16.125 191.075 18.715 192.165 ;
        RECT 18.890 191.730 24.235 192.165 ;
        RECT 16.125 190.555 17.335 191.075 ;
        RECT 17.505 190.385 18.715 190.905 ;
        RECT 20.480 190.480 20.830 191.730 ;
        RECT 24.405 191.000 24.695 192.165 ;
        RECT 25.785 191.075 29.295 192.165 ;
        RECT 29.470 191.730 34.815 192.165 ;
        RECT 34.990 191.730 40.335 192.165 ;
        RECT 14.745 189.615 15.955 190.365 ;
        RECT 16.125 189.615 18.715 190.385 ;
        RECT 22.310 190.160 22.650 190.990 ;
        RECT 25.785 190.555 27.475 191.075 ;
        RECT 27.645 190.385 29.295 190.905 ;
        RECT 31.060 190.480 31.410 191.730 ;
        RECT 18.890 189.615 24.235 190.160 ;
        RECT 24.405 189.615 24.695 190.340 ;
        RECT 25.785 189.615 29.295 190.385 ;
        RECT 32.890 190.160 33.230 190.990 ;
        RECT 36.580 190.480 36.930 191.730 ;
        RECT 40.880 191.185 41.135 191.855 ;
        RECT 41.315 191.365 41.600 192.165 ;
        RECT 41.780 191.445 42.110 191.955 ;
        RECT 40.880 191.145 41.060 191.185 ;
        RECT 38.410 190.160 38.750 190.990 ;
        RECT 40.795 190.975 41.060 191.145 ;
        RECT 40.880 190.325 41.060 190.975 ;
        RECT 41.780 190.855 42.030 191.445 ;
        RECT 42.380 191.295 42.550 191.905 ;
        RECT 42.720 191.475 43.050 192.165 ;
        RECT 43.280 191.615 43.520 191.905 ;
        RECT 43.720 191.785 44.140 192.165 ;
        RECT 44.320 191.695 44.950 191.945 ;
        RECT 45.420 191.785 45.750 192.165 ;
        RECT 44.320 191.615 44.490 191.695 ;
        RECT 45.920 191.615 46.090 191.905 ;
        RECT 46.270 191.785 46.650 192.165 ;
        RECT 46.890 191.780 47.720 191.950 ;
        RECT 43.280 191.445 44.490 191.615 ;
        RECT 41.230 190.525 42.030 190.855 ;
        RECT 29.470 189.615 34.815 190.160 ;
        RECT 34.990 189.615 40.335 190.160 ;
        RECT 40.880 189.795 41.135 190.325 ;
        RECT 41.315 189.615 41.600 190.075 ;
        RECT 41.780 189.875 42.030 190.525 ;
        RECT 42.230 191.275 42.550 191.295 ;
        RECT 42.230 191.105 44.150 191.275 ;
        RECT 42.230 190.210 42.420 191.105 ;
        RECT 44.320 190.935 44.490 191.445 ;
        RECT 44.660 191.185 45.180 191.495 ;
        RECT 42.590 190.765 44.490 190.935 ;
        RECT 42.590 190.705 42.920 190.765 ;
        RECT 43.070 190.535 43.400 190.595 ;
        RECT 42.740 190.265 43.400 190.535 ;
        RECT 42.230 189.880 42.550 190.210 ;
        RECT 42.730 189.615 43.390 190.095 ;
        RECT 43.590 190.005 43.760 190.765 ;
        RECT 44.660 190.595 44.840 191.005 ;
        RECT 43.930 190.425 44.260 190.545 ;
        RECT 45.010 190.425 45.180 191.185 ;
        RECT 43.930 190.255 45.180 190.425 ;
        RECT 45.350 191.365 46.720 191.615 ;
        RECT 45.350 190.595 45.540 191.365 ;
        RECT 46.470 191.105 46.720 191.365 ;
        RECT 45.710 190.935 45.960 191.095 ;
        RECT 46.890 190.935 47.060 191.780 ;
        RECT 47.955 191.495 48.125 191.995 ;
        RECT 48.295 191.665 48.625 192.165 ;
        RECT 47.230 191.105 47.730 191.485 ;
        RECT 47.955 191.325 48.650 191.495 ;
        RECT 45.710 190.765 47.060 190.935 ;
        RECT 46.640 190.725 47.060 190.765 ;
        RECT 45.350 190.255 45.770 190.595 ;
        RECT 46.060 190.265 46.470 190.595 ;
        RECT 43.590 189.835 44.440 190.005 ;
        RECT 45.000 189.615 45.320 190.075 ;
        RECT 45.520 189.825 45.770 190.255 ;
        RECT 46.060 189.615 46.470 190.055 ;
        RECT 46.640 189.995 46.810 190.725 ;
        RECT 46.980 190.175 47.330 190.545 ;
        RECT 47.510 190.235 47.730 191.105 ;
        RECT 47.900 190.535 48.310 191.155 ;
        RECT 48.480 190.355 48.650 191.325 ;
        RECT 47.955 190.165 48.650 190.355 ;
        RECT 46.640 189.795 47.655 189.995 ;
        RECT 47.955 189.835 48.125 190.165 ;
        RECT 48.295 189.615 48.625 189.995 ;
        RECT 48.840 189.875 49.065 191.995 ;
        RECT 49.235 191.665 49.565 192.165 ;
        RECT 49.735 191.495 49.905 191.995 ;
        RECT 49.240 191.325 49.905 191.495 ;
        RECT 49.240 190.335 49.470 191.325 ;
        RECT 49.640 190.505 49.990 191.155 ;
        RECT 50.165 191.000 50.455 192.165 ;
        RECT 51.000 191.185 51.255 191.855 ;
        RECT 51.435 191.365 51.720 192.165 ;
        RECT 51.900 191.445 52.230 191.955 ;
        RECT 49.240 190.165 49.905 190.335 ;
        RECT 49.235 189.615 49.565 189.995 ;
        RECT 49.735 189.875 49.905 190.165 ;
        RECT 50.165 189.615 50.455 190.340 ;
        RECT 51.000 190.325 51.180 191.185 ;
        RECT 51.900 190.855 52.150 191.445 ;
        RECT 52.500 191.295 52.670 191.905 ;
        RECT 52.840 191.475 53.170 192.165 ;
        RECT 53.400 191.615 53.640 191.905 ;
        RECT 53.840 191.785 54.260 192.165 ;
        RECT 54.440 191.695 55.070 191.945 ;
        RECT 55.540 191.785 55.870 192.165 ;
        RECT 54.440 191.615 54.610 191.695 ;
        RECT 56.040 191.615 56.210 191.905 ;
        RECT 56.390 191.785 56.770 192.165 ;
        RECT 57.010 191.780 57.840 191.950 ;
        RECT 53.400 191.445 54.610 191.615 ;
        RECT 51.350 190.525 52.150 190.855 ;
        RECT 51.000 190.125 51.255 190.325 ;
        RECT 50.915 189.955 51.255 190.125 ;
        RECT 51.000 189.795 51.255 189.955 ;
        RECT 51.435 189.615 51.720 190.075 ;
        RECT 51.900 189.875 52.150 190.525 ;
        RECT 52.350 191.275 52.670 191.295 ;
        RECT 52.350 191.105 54.270 191.275 ;
        RECT 52.350 190.210 52.540 191.105 ;
        RECT 54.440 190.935 54.610 191.445 ;
        RECT 54.780 191.185 55.300 191.495 ;
        RECT 52.710 190.765 54.610 190.935 ;
        RECT 52.710 190.705 53.040 190.765 ;
        RECT 53.190 190.535 53.520 190.595 ;
        RECT 52.860 190.265 53.520 190.535 ;
        RECT 52.350 189.880 52.670 190.210 ;
        RECT 52.850 189.615 53.510 190.095 ;
        RECT 53.710 190.005 53.880 190.765 ;
        RECT 54.780 190.595 54.960 191.005 ;
        RECT 54.050 190.425 54.380 190.545 ;
        RECT 55.130 190.425 55.300 191.185 ;
        RECT 54.050 190.255 55.300 190.425 ;
        RECT 55.470 191.365 56.840 191.615 ;
        RECT 55.470 190.595 55.660 191.365 ;
        RECT 56.590 191.105 56.840 191.365 ;
        RECT 55.830 190.935 56.080 191.095 ;
        RECT 57.010 190.935 57.180 191.780 ;
        RECT 58.075 191.495 58.245 191.995 ;
        RECT 58.415 191.665 58.745 192.165 ;
        RECT 57.350 191.105 57.850 191.485 ;
        RECT 58.075 191.325 58.770 191.495 ;
        RECT 55.830 190.765 57.180 190.935 ;
        RECT 56.760 190.725 57.180 190.765 ;
        RECT 55.470 190.255 55.890 190.595 ;
        RECT 56.180 190.265 56.590 190.595 ;
        RECT 53.710 189.835 54.560 190.005 ;
        RECT 55.120 189.615 55.440 190.075 ;
        RECT 55.640 189.825 55.890 190.255 ;
        RECT 56.180 189.615 56.590 190.055 ;
        RECT 56.760 189.995 56.930 190.725 ;
        RECT 57.100 190.175 57.450 190.545 ;
        RECT 57.630 190.235 57.850 191.105 ;
        RECT 58.020 190.535 58.430 191.155 ;
        RECT 58.600 190.355 58.770 191.325 ;
        RECT 58.075 190.165 58.770 190.355 ;
        RECT 56.760 189.795 57.775 189.995 ;
        RECT 58.075 189.835 58.245 190.165 ;
        RECT 58.415 189.615 58.745 189.995 ;
        RECT 58.960 189.875 59.185 191.995 ;
        RECT 59.355 191.665 59.685 192.165 ;
        RECT 59.855 191.495 60.025 191.995 ;
        RECT 59.360 191.325 60.025 191.495 ;
        RECT 59.360 190.335 59.590 191.325 ;
        RECT 59.760 190.505 60.110 191.155 ;
        RECT 60.745 191.075 63.335 192.165 ;
        RECT 63.510 191.730 68.855 192.165 ;
        RECT 60.745 190.555 61.955 191.075 ;
        RECT 62.125 190.385 63.335 190.905 ;
        RECT 65.100 190.480 65.450 191.730 ;
        RECT 69.045 191.365 69.325 192.165 ;
        RECT 69.525 191.195 69.855 191.995 ;
        RECT 70.055 191.365 70.225 192.165 ;
        RECT 70.395 191.195 70.725 191.995 ;
        RECT 59.360 190.165 60.025 190.335 ;
        RECT 59.355 189.615 59.685 189.995 ;
        RECT 59.855 189.875 60.025 190.165 ;
        RECT 60.745 189.615 63.335 190.385 ;
        RECT 66.930 190.160 67.270 190.990 ;
        RECT 69.025 190.525 69.265 191.195 ;
        RECT 69.445 191.025 70.725 191.195 ;
        RECT 70.895 191.025 71.155 192.165 ;
        RECT 72.245 191.075 75.755 192.165 ;
        RECT 69.445 190.355 69.615 191.025 ;
        RECT 69.785 190.525 70.095 190.855 ;
        RECT 70.265 190.525 70.645 190.855 ;
        RECT 70.845 190.525 71.130 190.855 ;
        RECT 72.245 190.555 73.935 191.075 ;
        RECT 75.925 191.000 76.215 192.165 ;
        RECT 76.385 191.075 77.595 192.165 ;
        RECT 77.765 191.075 81.275 192.165 ;
        RECT 69.890 190.355 70.095 190.525 ;
        RECT 63.510 189.615 68.855 190.160 ;
        RECT 69.025 189.785 69.720 190.355 ;
        RECT 69.890 189.830 70.240 190.355 ;
        RECT 70.430 189.830 70.645 190.525 ;
        RECT 74.105 190.385 75.755 190.905 ;
        RECT 76.385 190.535 76.905 191.075 ;
        RECT 70.815 189.615 71.150 190.355 ;
        RECT 72.245 189.615 75.755 190.385 ;
        RECT 77.075 190.365 77.595 190.905 ;
        RECT 77.765 190.555 79.455 191.075 ;
        RECT 81.485 191.025 81.715 192.165 ;
        RECT 81.885 191.015 82.215 191.995 ;
        RECT 82.385 191.025 82.595 192.165 ;
        RECT 82.885 191.025 83.095 192.165 ;
        RECT 79.625 190.385 81.275 190.905 ;
        RECT 81.465 190.605 81.795 190.855 ;
        RECT 75.925 189.615 76.215 190.340 ;
        RECT 76.385 189.615 77.595 190.365 ;
        RECT 77.765 189.615 81.275 190.385 ;
        RECT 81.485 189.615 81.715 190.435 ;
        RECT 81.965 190.415 82.215 191.015 ;
        RECT 83.265 191.015 83.595 191.995 ;
        RECT 83.765 191.025 83.995 192.165 ;
        RECT 84.580 191.185 84.835 191.855 ;
        RECT 85.015 191.365 85.300 192.165 ;
        RECT 85.480 191.445 85.810 191.955 ;
        RECT 84.580 191.145 84.760 191.185 ;
        RECT 81.885 189.785 82.215 190.415 ;
        RECT 82.385 189.615 82.595 190.435 ;
        RECT 82.885 189.615 83.095 190.435 ;
        RECT 83.265 190.415 83.515 191.015 ;
        RECT 84.495 190.975 84.760 191.145 ;
        RECT 83.685 190.605 84.015 190.855 ;
        RECT 83.265 189.785 83.595 190.415 ;
        RECT 83.765 189.615 83.995 190.435 ;
        RECT 84.580 190.325 84.760 190.975 ;
        RECT 85.480 190.855 85.730 191.445 ;
        RECT 86.080 191.295 86.250 191.905 ;
        RECT 86.420 191.475 86.750 192.165 ;
        RECT 86.980 191.615 87.220 191.905 ;
        RECT 87.420 191.785 87.840 192.165 ;
        RECT 88.020 191.695 88.650 191.945 ;
        RECT 89.120 191.785 89.450 192.165 ;
        RECT 88.020 191.615 88.190 191.695 ;
        RECT 89.620 191.615 89.790 191.905 ;
        RECT 89.970 191.785 90.350 192.165 ;
        RECT 90.590 191.780 91.420 191.950 ;
        RECT 86.980 191.445 88.190 191.615 ;
        RECT 84.930 190.525 85.730 190.855 ;
        RECT 84.580 189.795 84.835 190.325 ;
        RECT 85.015 189.615 85.300 190.075 ;
        RECT 85.480 189.875 85.730 190.525 ;
        RECT 85.930 191.275 86.250 191.295 ;
        RECT 85.930 191.105 87.850 191.275 ;
        RECT 85.930 190.210 86.120 191.105 ;
        RECT 88.020 190.935 88.190 191.445 ;
        RECT 88.360 191.185 88.880 191.495 ;
        RECT 86.290 190.765 88.190 190.935 ;
        RECT 86.290 190.705 86.620 190.765 ;
        RECT 86.770 190.535 87.100 190.595 ;
        RECT 86.440 190.265 87.100 190.535 ;
        RECT 85.930 189.880 86.250 190.210 ;
        RECT 86.430 189.615 87.090 190.095 ;
        RECT 87.290 190.005 87.460 190.765 ;
        RECT 88.360 190.595 88.540 191.005 ;
        RECT 87.630 190.425 87.960 190.545 ;
        RECT 88.710 190.425 88.880 191.185 ;
        RECT 87.630 190.255 88.880 190.425 ;
        RECT 89.050 191.365 90.420 191.615 ;
        RECT 89.050 190.595 89.240 191.365 ;
        RECT 90.170 191.105 90.420 191.365 ;
        RECT 89.410 190.935 89.660 191.095 ;
        RECT 90.590 190.935 90.760 191.780 ;
        RECT 91.655 191.495 91.825 191.995 ;
        RECT 91.995 191.665 92.325 192.165 ;
        RECT 90.930 191.105 91.430 191.485 ;
        RECT 91.655 191.325 92.350 191.495 ;
        RECT 89.410 190.765 90.760 190.935 ;
        RECT 90.340 190.725 90.760 190.765 ;
        RECT 89.050 190.255 89.470 190.595 ;
        RECT 89.760 190.265 90.170 190.595 ;
        RECT 87.290 189.835 88.140 190.005 ;
        RECT 88.700 189.615 89.020 190.075 ;
        RECT 89.220 189.825 89.470 190.255 ;
        RECT 89.760 189.615 90.170 190.055 ;
        RECT 90.340 189.995 90.510 190.725 ;
        RECT 90.680 190.175 91.030 190.545 ;
        RECT 91.210 190.235 91.430 191.105 ;
        RECT 91.600 190.535 92.010 191.155 ;
        RECT 92.180 190.355 92.350 191.325 ;
        RECT 91.655 190.165 92.350 190.355 ;
        RECT 90.340 189.795 91.355 189.995 ;
        RECT 91.655 189.835 91.825 190.165 ;
        RECT 91.995 189.615 92.325 189.995 ;
        RECT 92.540 189.875 92.765 191.995 ;
        RECT 92.935 191.665 93.265 192.165 ;
        RECT 93.435 191.495 93.605 191.995 ;
        RECT 92.940 191.325 93.605 191.495 ;
        RECT 92.940 190.335 93.170 191.325 ;
        RECT 93.340 190.505 93.690 191.155 ;
        RECT 94.325 191.075 95.995 192.165 ;
        RECT 96.170 191.730 101.515 192.165 ;
        RECT 94.325 190.555 95.075 191.075 ;
        RECT 95.245 190.385 95.995 190.905 ;
        RECT 97.760 190.480 98.110 191.730 ;
        RECT 101.685 191.000 101.975 192.165 ;
        RECT 102.145 191.075 103.355 192.165 ;
        RECT 92.940 190.165 93.605 190.335 ;
        RECT 92.935 189.615 93.265 189.995 ;
        RECT 93.435 189.875 93.605 190.165 ;
        RECT 94.325 189.615 95.995 190.385 ;
        RECT 99.590 190.160 99.930 190.990 ;
        RECT 102.145 190.535 102.665 191.075 ;
        RECT 103.530 190.975 103.785 191.855 ;
        RECT 103.955 191.025 104.260 192.165 ;
        RECT 104.600 191.785 104.930 192.165 ;
        RECT 105.110 191.615 105.280 191.905 ;
        RECT 105.450 191.705 105.700 192.165 ;
        RECT 104.480 191.445 105.280 191.615 ;
        RECT 105.870 191.655 106.740 191.995 ;
        RECT 102.835 190.365 103.355 190.905 ;
        RECT 96.170 189.615 101.515 190.160 ;
        RECT 101.685 189.615 101.975 190.340 ;
        RECT 102.145 189.615 103.355 190.365 ;
        RECT 103.530 190.325 103.740 190.975 ;
        RECT 104.480 190.855 104.650 191.445 ;
        RECT 105.870 191.275 106.040 191.655 ;
        RECT 106.975 191.535 107.145 191.995 ;
        RECT 107.315 191.705 107.685 192.165 ;
        RECT 107.980 191.565 108.150 191.905 ;
        RECT 108.320 191.735 108.650 192.165 ;
        RECT 108.885 191.565 109.055 191.905 ;
        RECT 104.820 191.105 106.040 191.275 ;
        RECT 106.210 191.195 106.670 191.485 ;
        RECT 106.975 191.365 107.535 191.535 ;
        RECT 107.980 191.395 109.055 191.565 ;
        RECT 109.225 191.665 109.905 191.995 ;
        RECT 110.120 191.665 110.370 191.995 ;
        RECT 110.540 191.705 110.790 192.165 ;
        RECT 107.365 191.225 107.535 191.365 ;
        RECT 106.210 191.185 107.175 191.195 ;
        RECT 105.870 191.015 106.040 191.105 ;
        RECT 106.500 191.025 107.175 191.185 ;
        RECT 103.910 190.825 104.650 190.855 ;
        RECT 103.910 190.525 104.825 190.825 ;
        RECT 104.500 190.350 104.825 190.525 ;
        RECT 103.530 189.795 103.785 190.325 ;
        RECT 103.955 189.615 104.260 190.075 ;
        RECT 104.505 189.995 104.825 190.350 ;
        RECT 104.995 190.565 105.535 190.935 ;
        RECT 105.870 190.845 106.275 191.015 ;
        RECT 104.995 190.165 105.235 190.565 ;
        RECT 105.715 190.395 105.935 190.675 ;
        RECT 105.405 190.225 105.935 190.395 ;
        RECT 105.405 189.995 105.575 190.225 ;
        RECT 106.105 190.065 106.275 190.845 ;
        RECT 106.445 190.235 106.795 190.855 ;
        RECT 106.965 190.235 107.175 191.025 ;
        RECT 107.365 191.055 108.865 191.225 ;
        RECT 107.365 190.365 107.535 191.055 ;
        RECT 109.225 190.885 109.395 191.665 ;
        RECT 110.200 191.535 110.370 191.665 ;
        RECT 107.705 190.715 109.395 190.885 ;
        RECT 109.565 191.105 110.030 191.495 ;
        RECT 110.200 191.365 110.595 191.535 ;
        RECT 107.705 190.535 107.875 190.715 ;
        RECT 104.505 189.825 105.575 189.995 ;
        RECT 105.745 189.615 105.935 190.055 ;
        RECT 106.105 189.785 107.055 190.065 ;
        RECT 107.365 189.975 107.625 190.365 ;
        RECT 108.045 190.295 108.835 190.545 ;
        RECT 107.275 189.805 107.625 189.975 ;
        RECT 107.835 189.615 108.165 190.075 ;
        RECT 109.040 190.005 109.210 190.715 ;
        RECT 109.565 190.515 109.735 191.105 ;
        RECT 109.380 190.295 109.735 190.515 ;
        RECT 109.905 190.295 110.255 190.915 ;
        RECT 110.425 190.005 110.595 191.365 ;
        RECT 110.960 191.195 111.285 191.980 ;
        RECT 110.765 190.145 111.225 191.195 ;
        RECT 109.040 189.835 109.895 190.005 ;
        RECT 110.100 189.835 110.595 190.005 ;
        RECT 110.765 189.615 111.095 189.975 ;
        RECT 111.455 189.875 111.625 191.995 ;
        RECT 111.795 191.665 112.125 192.165 ;
        RECT 112.295 191.495 112.550 191.995 ;
        RECT 111.800 191.325 112.550 191.495 ;
        RECT 111.800 190.335 112.030 191.325 ;
        RECT 112.200 190.505 112.550 191.155 ;
        RECT 112.725 191.075 113.935 192.165 ;
        RECT 114.105 191.075 117.615 192.165 ;
        RECT 112.725 190.535 113.245 191.075 ;
        RECT 113.415 190.365 113.935 190.905 ;
        RECT 114.105 190.555 115.795 191.075 ;
        RECT 117.845 191.025 118.055 192.165 ;
        RECT 118.225 191.015 118.555 191.995 ;
        RECT 118.725 191.025 118.955 192.165 ;
        RECT 119.165 191.075 120.835 192.165 ;
        RECT 121.010 191.730 126.355 192.165 ;
        RECT 115.965 190.385 117.615 190.905 ;
        RECT 111.800 190.165 112.550 190.335 ;
        RECT 111.795 189.615 112.125 189.995 ;
        RECT 112.295 189.875 112.550 190.165 ;
        RECT 112.725 189.615 113.935 190.365 ;
        RECT 114.105 189.615 117.615 190.385 ;
        RECT 117.845 189.615 118.055 190.435 ;
        RECT 118.225 190.415 118.475 191.015 ;
        RECT 118.645 190.605 118.975 190.855 ;
        RECT 119.165 190.555 119.915 191.075 ;
        RECT 118.225 189.785 118.555 190.415 ;
        RECT 118.725 189.615 118.955 190.435 ;
        RECT 120.085 190.385 120.835 190.905 ;
        RECT 122.600 190.480 122.950 191.730 ;
        RECT 126.525 191.075 127.735 192.165 ;
        RECT 119.165 189.615 120.835 190.385 ;
        RECT 124.430 190.160 124.770 190.990 ;
        RECT 126.525 190.535 127.045 191.075 ;
        RECT 127.215 190.365 127.735 190.905 ;
        RECT 121.010 189.615 126.355 190.160 ;
        RECT 126.525 189.615 127.735 190.365 ;
        RECT 14.660 189.445 127.820 189.615 ;
        RECT 14.745 188.695 15.955 189.445 ;
        RECT 14.745 188.155 15.265 188.695 ;
        RECT 17.045 188.675 20.555 189.445 ;
        RECT 20.730 188.900 26.075 189.445 ;
        RECT 26.250 188.900 31.595 189.445 ;
        RECT 31.770 188.900 37.115 189.445 ;
        RECT 15.435 187.985 15.955 188.525 ;
        RECT 14.745 186.895 15.955 187.985 ;
        RECT 17.045 187.985 18.735 188.505 ;
        RECT 18.905 188.155 20.555 188.675 ;
        RECT 17.045 186.895 20.555 187.985 ;
        RECT 22.320 187.330 22.670 188.580 ;
        RECT 24.150 188.070 24.490 188.900 ;
        RECT 27.840 187.330 28.190 188.580 ;
        RECT 29.670 188.070 30.010 188.900 ;
        RECT 33.360 187.330 33.710 188.580 ;
        RECT 35.190 188.070 35.530 188.900 ;
        RECT 37.285 188.720 37.575 189.445 ;
        RECT 37.745 188.675 41.255 189.445 ;
        RECT 41.430 188.900 46.775 189.445 ;
        RECT 20.730 186.895 26.075 187.330 ;
        RECT 26.250 186.895 31.595 187.330 ;
        RECT 31.770 186.895 37.115 187.330 ;
        RECT 37.285 186.895 37.575 188.060 ;
        RECT 37.745 187.985 39.435 188.505 ;
        RECT 39.605 188.155 41.255 188.675 ;
        RECT 37.745 186.895 41.255 187.985 ;
        RECT 43.020 187.330 43.370 188.580 ;
        RECT 44.850 188.070 45.190 188.900 ;
        RECT 47.220 188.635 47.465 189.240 ;
        RECT 47.685 188.910 48.195 189.445 ;
        RECT 46.945 188.465 48.175 188.635 ;
        RECT 46.945 187.655 47.285 188.465 ;
        RECT 47.455 187.900 48.205 188.090 ;
        RECT 41.430 186.895 46.775 187.330 ;
        RECT 46.945 187.245 47.460 187.655 ;
        RECT 47.695 186.895 47.865 187.655 ;
        RECT 48.035 187.235 48.205 187.900 ;
        RECT 48.375 187.915 48.565 189.275 ;
        RECT 48.735 188.425 49.010 189.275 ;
        RECT 49.200 188.910 49.730 189.275 ;
        RECT 50.155 189.045 50.485 189.445 ;
        RECT 49.555 188.875 49.730 188.910 ;
        RECT 48.735 188.255 49.015 188.425 ;
        RECT 48.735 188.115 49.010 188.255 ;
        RECT 49.215 187.915 49.385 188.715 ;
        RECT 48.375 187.745 49.385 187.915 ;
        RECT 49.555 188.705 50.485 188.875 ;
        RECT 50.655 188.705 50.910 189.275 ;
        RECT 49.555 187.575 49.725 188.705 ;
        RECT 50.315 188.535 50.485 188.705 ;
        RECT 48.600 187.405 49.725 187.575 ;
        RECT 49.895 188.205 50.090 188.535 ;
        RECT 50.315 188.205 50.570 188.535 ;
        RECT 49.895 187.235 50.065 188.205 ;
        RECT 50.740 188.035 50.910 188.705 ;
        RECT 51.360 188.635 51.605 189.240 ;
        RECT 51.825 188.910 52.335 189.445 ;
        RECT 48.035 187.065 50.065 187.235 ;
        RECT 50.235 186.895 50.405 188.035 ;
        RECT 50.575 187.065 50.910 188.035 ;
        RECT 51.085 188.465 52.315 188.635 ;
        RECT 51.085 187.655 51.425 188.465 ;
        RECT 51.595 187.900 52.345 188.090 ;
        RECT 51.085 187.245 51.600 187.655 ;
        RECT 51.835 186.895 52.005 187.655 ;
        RECT 52.175 187.235 52.345 187.900 ;
        RECT 52.515 187.915 52.705 189.275 ;
        RECT 52.875 188.425 53.150 189.275 ;
        RECT 53.340 188.910 53.870 189.275 ;
        RECT 54.295 189.045 54.625 189.445 ;
        RECT 53.695 188.875 53.870 188.910 ;
        RECT 52.875 188.255 53.155 188.425 ;
        RECT 52.875 188.115 53.150 188.255 ;
        RECT 53.355 187.915 53.525 188.715 ;
        RECT 52.515 187.745 53.525 187.915 ;
        RECT 53.695 188.705 54.625 188.875 ;
        RECT 54.795 188.705 55.050 189.275 ;
        RECT 53.695 187.575 53.865 188.705 ;
        RECT 54.455 188.535 54.625 188.705 ;
        RECT 52.740 187.405 53.865 187.575 ;
        RECT 54.035 188.205 54.230 188.535 ;
        RECT 54.455 188.205 54.710 188.535 ;
        RECT 54.035 187.235 54.205 188.205 ;
        RECT 54.880 188.035 55.050 188.705 ;
        RECT 55.725 188.625 55.955 189.445 ;
        RECT 56.125 188.645 56.455 189.275 ;
        RECT 55.705 188.205 56.035 188.455 ;
        RECT 56.205 188.045 56.455 188.645 ;
        RECT 56.625 188.625 56.835 189.445 ;
        RECT 57.155 188.895 57.325 189.275 ;
        RECT 57.505 189.065 57.835 189.445 ;
        RECT 57.155 188.725 57.820 188.895 ;
        RECT 58.015 188.770 58.275 189.275 ;
        RECT 57.085 188.175 57.415 188.545 ;
        RECT 57.650 188.470 57.820 188.725 ;
        RECT 52.175 187.065 54.205 187.235 ;
        RECT 54.375 186.895 54.545 188.035 ;
        RECT 54.715 187.065 55.050 188.035 ;
        RECT 55.725 186.895 55.955 188.035 ;
        RECT 56.125 187.065 56.455 188.045 ;
        RECT 57.650 188.140 57.935 188.470 ;
        RECT 56.625 186.895 56.835 188.035 ;
        RECT 57.650 187.995 57.820 188.140 ;
        RECT 57.155 187.825 57.820 187.995 ;
        RECT 58.105 187.970 58.275 188.770 ;
        RECT 59.365 188.675 62.875 189.445 ;
        RECT 63.045 188.720 63.335 189.445 ;
        RECT 63.505 188.675 65.175 189.445 ;
        RECT 57.155 187.065 57.325 187.825 ;
        RECT 57.505 186.895 57.835 187.655 ;
        RECT 58.005 187.065 58.275 187.970 ;
        RECT 59.365 187.985 61.055 188.505 ;
        RECT 61.225 188.155 62.875 188.675 ;
        RECT 59.365 186.895 62.875 187.985 ;
        RECT 63.045 186.895 63.335 188.060 ;
        RECT 63.505 187.985 64.255 188.505 ;
        RECT 64.425 188.155 65.175 188.675 ;
        RECT 65.385 188.625 65.615 189.445 ;
        RECT 65.785 188.645 66.115 189.275 ;
        RECT 65.365 188.205 65.695 188.455 ;
        RECT 65.865 188.045 66.115 188.645 ;
        RECT 66.285 188.625 66.495 189.445 ;
        RECT 66.725 188.945 66.985 189.275 ;
        RECT 67.195 188.965 67.470 189.445 ;
        RECT 63.505 186.895 65.175 187.985 ;
        RECT 65.385 186.895 65.615 188.035 ;
        RECT 65.785 187.065 66.115 188.045 ;
        RECT 66.725 188.035 66.895 188.945 ;
        RECT 67.680 188.875 67.885 189.275 ;
        RECT 68.055 189.045 68.390 189.445 ;
        RECT 67.065 188.205 67.425 188.785 ;
        RECT 67.680 188.705 68.365 188.875 ;
        RECT 67.605 188.035 67.855 188.535 ;
        RECT 66.285 186.895 66.495 188.035 ;
        RECT 66.725 187.865 67.855 188.035 ;
        RECT 66.725 187.095 66.995 187.865 ;
        RECT 68.025 187.675 68.365 188.705 ;
        RECT 69.490 188.605 69.750 189.445 ;
        RECT 69.925 188.700 70.180 189.275 ;
        RECT 70.350 189.065 70.680 189.445 ;
        RECT 70.895 188.895 71.065 189.275 ;
        RECT 70.350 188.725 71.065 188.895 ;
        RECT 67.165 186.895 67.495 187.675 ;
        RECT 67.700 187.500 68.365 187.675 ;
        RECT 67.700 187.095 67.885 187.500 ;
        RECT 68.055 186.895 68.390 187.320 ;
        RECT 69.490 186.895 69.750 188.045 ;
        RECT 69.925 187.970 70.095 188.700 ;
        RECT 70.350 188.535 70.520 188.725 ;
        RECT 71.325 188.675 72.995 189.445 ;
        RECT 70.265 188.205 70.520 188.535 ;
        RECT 70.350 187.995 70.520 188.205 ;
        RECT 70.800 188.175 71.155 188.545 ;
        RECT 69.925 187.065 70.180 187.970 ;
        RECT 70.350 187.825 71.065 187.995 ;
        RECT 70.350 186.895 70.680 187.655 ;
        RECT 70.895 187.065 71.065 187.825 ;
        RECT 71.325 187.985 72.075 188.505 ;
        RECT 72.245 188.155 72.995 188.675 ;
        RECT 73.205 188.625 73.435 189.445 ;
        RECT 73.605 188.645 73.935 189.275 ;
        RECT 73.185 188.205 73.515 188.455 ;
        RECT 73.685 188.045 73.935 188.645 ;
        RECT 74.105 188.625 74.315 189.445 ;
        RECT 75.465 188.675 78.975 189.445 ;
        RECT 71.325 186.895 72.995 187.985 ;
        RECT 73.205 186.895 73.435 188.035 ;
        RECT 73.605 187.065 73.935 188.045 ;
        RECT 74.105 186.895 74.315 188.035 ;
        RECT 75.465 187.985 77.155 188.505 ;
        RECT 77.325 188.155 78.975 188.675 ;
        RECT 79.520 188.735 79.775 189.265 ;
        RECT 79.955 188.985 80.240 189.445 ;
        RECT 79.520 188.085 79.700 188.735 ;
        RECT 80.420 188.535 80.670 189.185 ;
        RECT 79.870 188.205 80.670 188.535 ;
        RECT 75.465 186.895 78.975 187.985 ;
        RECT 79.435 187.915 79.700 188.085 ;
        RECT 79.520 187.875 79.700 187.915 ;
        RECT 79.520 187.205 79.775 187.875 ;
        RECT 79.955 186.895 80.240 187.695 ;
        RECT 80.420 187.615 80.670 188.205 ;
        RECT 80.870 188.850 81.190 189.180 ;
        RECT 81.370 188.965 82.030 189.445 ;
        RECT 82.230 189.055 83.080 189.225 ;
        RECT 80.870 187.955 81.060 188.850 ;
        RECT 81.380 188.525 82.040 188.795 ;
        RECT 81.710 188.465 82.040 188.525 ;
        RECT 81.230 188.295 81.560 188.355 ;
        RECT 82.230 188.295 82.400 189.055 ;
        RECT 83.640 188.985 83.960 189.445 ;
        RECT 84.160 188.805 84.410 189.235 ;
        RECT 84.700 189.005 85.110 189.445 ;
        RECT 85.280 189.065 86.295 189.265 ;
        RECT 82.570 188.635 83.820 188.805 ;
        RECT 82.570 188.515 82.900 188.635 ;
        RECT 81.230 188.125 83.130 188.295 ;
        RECT 80.870 187.785 82.790 187.955 ;
        RECT 80.870 187.765 81.190 187.785 ;
        RECT 80.420 187.105 80.750 187.615 ;
        RECT 81.020 187.155 81.190 187.765 ;
        RECT 82.960 187.615 83.130 188.125 ;
        RECT 83.300 188.055 83.480 188.465 ;
        RECT 83.650 187.875 83.820 188.635 ;
        RECT 81.360 186.895 81.690 187.585 ;
        RECT 81.920 187.445 83.130 187.615 ;
        RECT 83.300 187.565 83.820 187.875 ;
        RECT 83.990 188.465 84.410 188.805 ;
        RECT 84.700 188.465 85.110 188.795 ;
        RECT 83.990 187.695 84.180 188.465 ;
        RECT 85.280 188.335 85.450 189.065 ;
        RECT 86.595 188.895 86.765 189.225 ;
        RECT 86.935 189.065 87.265 189.445 ;
        RECT 85.620 188.515 85.970 188.885 ;
        RECT 85.280 188.295 85.700 188.335 ;
        RECT 84.350 188.125 85.700 188.295 ;
        RECT 84.350 187.965 84.600 188.125 ;
        RECT 85.110 187.695 85.360 187.955 ;
        RECT 83.990 187.445 85.360 187.695 ;
        RECT 81.920 187.155 82.160 187.445 ;
        RECT 82.960 187.365 83.130 187.445 ;
        RECT 82.360 186.895 82.780 187.275 ;
        RECT 82.960 187.115 83.590 187.365 ;
        RECT 84.060 186.895 84.390 187.275 ;
        RECT 84.560 187.155 84.730 187.445 ;
        RECT 85.530 187.280 85.700 188.125 ;
        RECT 86.150 187.955 86.370 188.825 ;
        RECT 86.595 188.705 87.290 188.895 ;
        RECT 85.870 187.575 86.370 187.955 ;
        RECT 86.540 187.905 86.950 188.525 ;
        RECT 87.120 187.735 87.290 188.705 ;
        RECT 86.595 187.565 87.290 187.735 ;
        RECT 84.910 186.895 85.290 187.275 ;
        RECT 85.530 187.110 86.360 187.280 ;
        RECT 86.595 187.065 86.765 187.565 ;
        RECT 86.935 186.895 87.265 187.395 ;
        RECT 87.480 187.065 87.705 189.185 ;
        RECT 87.875 189.065 88.205 189.445 ;
        RECT 88.375 188.895 88.545 189.185 ;
        RECT 87.880 188.725 88.545 188.895 ;
        RECT 87.880 187.735 88.110 188.725 ;
        RECT 88.805 188.720 89.095 189.445 ;
        RECT 89.265 188.770 89.525 189.275 ;
        RECT 89.705 189.065 90.035 189.445 ;
        RECT 90.215 188.895 90.385 189.275 ;
        RECT 88.280 187.905 88.630 188.555 ;
        RECT 87.880 187.565 88.545 187.735 ;
        RECT 87.875 186.895 88.205 187.395 ;
        RECT 88.375 187.065 88.545 187.565 ;
        RECT 88.805 186.895 89.095 188.060 ;
        RECT 89.265 187.970 89.435 188.770 ;
        RECT 89.720 188.725 90.385 188.895 ;
        RECT 89.720 188.470 89.890 188.725 ;
        RECT 91.105 188.675 93.695 189.445 ;
        RECT 93.870 188.900 99.215 189.445 ;
        RECT 89.605 188.140 89.890 188.470 ;
        RECT 90.125 188.175 90.455 188.545 ;
        RECT 89.720 187.995 89.890 188.140 ;
        RECT 89.265 187.065 89.535 187.970 ;
        RECT 89.720 187.825 90.385 187.995 ;
        RECT 89.705 186.895 90.035 187.655 ;
        RECT 90.215 187.065 90.385 187.825 ;
        RECT 91.105 187.985 92.315 188.505 ;
        RECT 92.485 188.155 93.695 188.675 ;
        RECT 91.105 186.895 93.695 187.985 ;
        RECT 95.460 187.330 95.810 188.580 ;
        RECT 97.290 188.070 97.630 188.900 ;
        RECT 99.390 188.735 99.645 189.265 ;
        RECT 99.815 188.985 100.120 189.445 ;
        RECT 100.365 189.065 101.435 189.235 ;
        RECT 99.390 188.085 99.600 188.735 ;
        RECT 100.365 188.710 100.685 189.065 ;
        RECT 100.360 188.535 100.685 188.710 ;
        RECT 99.770 188.235 100.685 188.535 ;
        RECT 100.855 188.495 101.095 188.895 ;
        RECT 101.265 188.835 101.435 189.065 ;
        RECT 101.605 189.005 101.795 189.445 ;
        RECT 101.965 188.995 102.915 189.275 ;
        RECT 103.135 189.085 103.485 189.255 ;
        RECT 101.265 188.665 101.795 188.835 ;
        RECT 99.770 188.205 100.510 188.235 ;
        RECT 93.870 186.895 99.215 187.330 ;
        RECT 99.390 187.205 99.645 188.085 ;
        RECT 99.815 186.895 100.120 188.035 ;
        RECT 100.340 187.615 100.510 188.205 ;
        RECT 100.855 188.125 101.395 188.495 ;
        RECT 101.575 188.385 101.795 188.665 ;
        RECT 101.965 188.215 102.135 188.995 ;
        RECT 101.730 188.045 102.135 188.215 ;
        RECT 102.305 188.205 102.655 188.825 ;
        RECT 101.730 187.955 101.900 188.045 ;
        RECT 102.825 188.035 103.035 188.825 ;
        RECT 100.680 187.785 101.900 187.955 ;
        RECT 102.360 187.875 103.035 188.035 ;
        RECT 100.340 187.445 101.140 187.615 ;
        RECT 100.460 186.895 100.790 187.275 ;
        RECT 100.970 187.155 101.140 187.445 ;
        RECT 101.730 187.405 101.900 187.785 ;
        RECT 102.070 187.865 103.035 187.875 ;
        RECT 103.225 188.695 103.485 189.085 ;
        RECT 103.695 188.985 104.025 189.445 ;
        RECT 104.900 189.055 105.755 189.225 ;
        RECT 105.960 189.055 106.455 189.225 ;
        RECT 106.625 189.085 106.955 189.445 ;
        RECT 103.225 188.005 103.395 188.695 ;
        RECT 103.565 188.345 103.735 188.525 ;
        RECT 103.905 188.515 104.695 188.765 ;
        RECT 104.900 188.345 105.070 189.055 ;
        RECT 105.240 188.545 105.595 188.765 ;
        RECT 103.565 188.175 105.255 188.345 ;
        RECT 102.070 187.575 102.530 187.865 ;
        RECT 103.225 187.835 104.725 188.005 ;
        RECT 103.225 187.695 103.395 187.835 ;
        RECT 102.835 187.525 103.395 187.695 ;
        RECT 101.310 186.895 101.560 187.355 ;
        RECT 101.730 187.065 102.600 187.405 ;
        RECT 102.835 187.065 103.005 187.525 ;
        RECT 103.840 187.495 104.915 187.665 ;
        RECT 103.175 186.895 103.545 187.355 ;
        RECT 103.840 187.155 104.010 187.495 ;
        RECT 104.180 186.895 104.510 187.325 ;
        RECT 104.745 187.155 104.915 187.495 ;
        RECT 105.085 187.395 105.255 188.175 ;
        RECT 105.425 187.955 105.595 188.545 ;
        RECT 105.765 188.145 106.115 188.765 ;
        RECT 105.425 187.565 105.890 187.955 ;
        RECT 106.285 187.695 106.455 189.055 ;
        RECT 106.625 187.865 107.085 188.915 ;
        RECT 106.060 187.525 106.455 187.695 ;
        RECT 106.060 187.395 106.230 187.525 ;
        RECT 105.085 187.065 105.765 187.395 ;
        RECT 105.980 187.065 106.230 187.395 ;
        RECT 106.400 186.895 106.650 187.355 ;
        RECT 106.820 187.080 107.145 187.865 ;
        RECT 107.315 187.065 107.485 189.185 ;
        RECT 107.655 189.065 107.985 189.445 ;
        RECT 108.155 188.895 108.410 189.185 ;
        RECT 109.050 188.900 114.395 189.445 ;
        RECT 107.660 188.725 108.410 188.895 ;
        RECT 107.660 187.735 107.890 188.725 ;
        RECT 108.060 187.905 108.410 188.555 ;
        RECT 107.660 187.565 108.410 187.735 ;
        RECT 107.655 186.895 107.985 187.395 ;
        RECT 108.155 187.065 108.410 187.565 ;
        RECT 110.640 187.330 110.990 188.580 ;
        RECT 112.470 188.070 112.810 188.900 ;
        RECT 114.565 188.720 114.855 189.445 ;
        RECT 115.030 188.735 115.285 189.265 ;
        RECT 115.455 188.985 115.760 189.445 ;
        RECT 116.005 189.065 117.075 189.235 ;
        RECT 115.030 188.085 115.240 188.735 ;
        RECT 116.005 188.710 116.325 189.065 ;
        RECT 116.000 188.535 116.325 188.710 ;
        RECT 115.410 188.235 116.325 188.535 ;
        RECT 116.495 188.495 116.735 188.895 ;
        RECT 116.905 188.835 117.075 189.065 ;
        RECT 117.245 189.005 117.435 189.445 ;
        RECT 117.605 188.995 118.555 189.275 ;
        RECT 118.775 189.085 119.125 189.255 ;
        RECT 116.905 188.665 117.435 188.835 ;
        RECT 115.410 188.205 116.150 188.235 ;
        RECT 109.050 186.895 114.395 187.330 ;
        RECT 114.565 186.895 114.855 188.060 ;
        RECT 115.030 187.205 115.285 188.085 ;
        RECT 115.455 186.895 115.760 188.035 ;
        RECT 115.980 187.615 116.150 188.205 ;
        RECT 116.495 188.125 117.035 188.495 ;
        RECT 117.215 188.385 117.435 188.665 ;
        RECT 117.605 188.215 117.775 188.995 ;
        RECT 117.370 188.045 117.775 188.215 ;
        RECT 117.945 188.205 118.295 188.825 ;
        RECT 117.370 187.955 117.540 188.045 ;
        RECT 118.465 188.035 118.675 188.825 ;
        RECT 116.320 187.785 117.540 187.955 ;
        RECT 118.000 187.875 118.675 188.035 ;
        RECT 115.980 187.445 116.780 187.615 ;
        RECT 116.100 186.895 116.430 187.275 ;
        RECT 116.610 187.155 116.780 187.445 ;
        RECT 117.370 187.405 117.540 187.785 ;
        RECT 117.710 187.865 118.675 187.875 ;
        RECT 118.865 188.695 119.125 189.085 ;
        RECT 119.335 188.985 119.665 189.445 ;
        RECT 120.540 189.055 121.395 189.225 ;
        RECT 121.600 189.055 122.095 189.225 ;
        RECT 122.265 189.085 122.595 189.445 ;
        RECT 118.865 188.005 119.035 188.695 ;
        RECT 119.205 188.345 119.375 188.525 ;
        RECT 119.545 188.515 120.335 188.765 ;
        RECT 120.540 188.345 120.710 189.055 ;
        RECT 120.880 188.545 121.235 188.765 ;
        RECT 119.205 188.175 120.895 188.345 ;
        RECT 117.710 187.575 118.170 187.865 ;
        RECT 118.865 187.835 120.365 188.005 ;
        RECT 118.865 187.695 119.035 187.835 ;
        RECT 118.475 187.525 119.035 187.695 ;
        RECT 116.950 186.895 117.200 187.355 ;
        RECT 117.370 187.065 118.240 187.405 ;
        RECT 118.475 187.065 118.645 187.525 ;
        RECT 119.480 187.495 120.555 187.665 ;
        RECT 118.815 186.895 119.185 187.355 ;
        RECT 119.480 187.155 119.650 187.495 ;
        RECT 119.820 186.895 120.150 187.325 ;
        RECT 120.385 187.155 120.555 187.495 ;
        RECT 120.725 187.395 120.895 188.175 ;
        RECT 121.065 187.955 121.235 188.545 ;
        RECT 121.405 188.145 121.755 188.765 ;
        RECT 121.065 187.565 121.530 187.955 ;
        RECT 121.925 187.695 122.095 189.055 ;
        RECT 122.265 187.865 122.725 188.915 ;
        RECT 121.700 187.525 122.095 187.695 ;
        RECT 121.700 187.395 121.870 187.525 ;
        RECT 120.725 187.065 121.405 187.395 ;
        RECT 121.620 187.065 121.870 187.395 ;
        RECT 122.040 186.895 122.290 187.355 ;
        RECT 122.460 187.080 122.785 187.865 ;
        RECT 122.955 187.065 123.125 189.185 ;
        RECT 123.295 189.065 123.625 189.445 ;
        RECT 123.795 188.895 124.050 189.185 ;
        RECT 123.300 188.725 124.050 188.895 ;
        RECT 123.300 187.735 123.530 188.725 ;
        RECT 124.685 188.675 126.355 189.445 ;
        RECT 126.525 188.695 127.735 189.445 ;
        RECT 123.700 187.905 124.050 188.555 ;
        RECT 124.685 187.985 125.435 188.505 ;
        RECT 125.605 188.155 126.355 188.675 ;
        RECT 126.525 187.985 127.045 188.525 ;
        RECT 127.215 188.155 127.735 188.695 ;
        RECT 123.300 187.565 124.050 187.735 ;
        RECT 123.295 186.895 123.625 187.395 ;
        RECT 123.795 187.065 124.050 187.565 ;
        RECT 124.685 186.895 126.355 187.985 ;
        RECT 126.525 186.895 127.735 187.985 ;
        RECT 14.660 186.725 127.820 186.895 ;
        RECT 14.745 185.635 15.955 186.725 ;
        RECT 14.745 184.925 15.265 185.465 ;
        RECT 15.435 185.095 15.955 185.635 ;
        RECT 16.125 185.635 18.715 186.725 ;
        RECT 18.890 186.290 24.235 186.725 ;
        RECT 16.125 185.115 17.335 185.635 ;
        RECT 17.505 184.945 18.715 185.465 ;
        RECT 20.480 185.040 20.830 186.290 ;
        RECT 24.405 185.560 24.695 186.725 ;
        RECT 24.865 185.635 26.535 186.725 ;
        RECT 26.710 186.290 32.055 186.725 ;
        RECT 14.745 184.175 15.955 184.925 ;
        RECT 16.125 184.175 18.715 184.945 ;
        RECT 22.310 184.720 22.650 185.550 ;
        RECT 24.865 185.115 25.615 185.635 ;
        RECT 25.785 184.945 26.535 185.465 ;
        RECT 28.300 185.040 28.650 186.290 ;
        RECT 32.285 185.585 32.495 186.725 ;
        RECT 32.665 185.575 32.995 186.555 ;
        RECT 33.165 185.585 33.395 186.725 ;
        RECT 33.605 185.635 35.275 186.725 ;
        RECT 18.890 184.175 24.235 184.720 ;
        RECT 24.405 184.175 24.695 184.900 ;
        RECT 24.865 184.175 26.535 184.945 ;
        RECT 30.130 184.720 30.470 185.550 ;
        RECT 26.710 184.175 32.055 184.720 ;
        RECT 32.285 184.175 32.495 184.995 ;
        RECT 32.665 184.975 32.915 185.575 ;
        RECT 33.085 185.165 33.415 185.415 ;
        RECT 33.605 185.115 34.355 185.635 ;
        RECT 35.450 185.585 35.785 186.555 ;
        RECT 35.955 185.585 36.125 186.725 ;
        RECT 36.295 186.385 38.325 186.555 ;
        RECT 32.665 184.345 32.995 184.975 ;
        RECT 33.165 184.175 33.395 184.995 ;
        RECT 34.525 184.945 35.275 185.465 ;
        RECT 33.605 184.175 35.275 184.945 ;
        RECT 35.450 184.915 35.620 185.585 ;
        RECT 36.295 185.415 36.465 186.385 ;
        RECT 35.790 185.085 36.045 185.415 ;
        RECT 36.270 185.085 36.465 185.415 ;
        RECT 36.635 186.045 37.760 186.215 ;
        RECT 35.875 184.915 36.045 185.085 ;
        RECT 36.635 184.915 36.805 186.045 ;
        RECT 35.450 184.345 35.705 184.915 ;
        RECT 35.875 184.745 36.805 184.915 ;
        RECT 36.975 185.705 37.985 185.875 ;
        RECT 36.975 184.905 37.145 185.705 ;
        RECT 37.350 185.025 37.625 185.505 ;
        RECT 37.345 184.855 37.625 185.025 ;
        RECT 36.630 184.710 36.805 184.745 ;
        RECT 35.875 184.175 36.205 184.575 ;
        RECT 36.630 184.345 37.160 184.710 ;
        RECT 37.350 184.345 37.625 184.855 ;
        RECT 37.795 184.345 37.985 185.705 ;
        RECT 38.155 185.720 38.325 186.385 ;
        RECT 38.495 185.965 38.665 186.725 ;
        RECT 38.900 185.965 39.415 186.375 ;
        RECT 38.155 185.530 38.905 185.720 ;
        RECT 39.075 185.155 39.415 185.965 ;
        RECT 38.185 184.985 39.415 185.155 ;
        RECT 39.585 185.635 41.255 186.725 ;
        RECT 41.425 185.965 41.940 186.375 ;
        RECT 42.175 185.965 42.345 186.725 ;
        RECT 42.515 186.385 44.545 186.555 ;
        RECT 39.585 185.115 40.335 185.635 ;
        RECT 38.165 184.175 38.675 184.710 ;
        RECT 38.895 184.380 39.140 184.985 ;
        RECT 40.505 184.945 41.255 185.465 ;
        RECT 41.425 185.155 41.765 185.965 ;
        RECT 42.515 185.720 42.685 186.385 ;
        RECT 43.080 186.045 44.205 186.215 ;
        RECT 41.935 185.530 42.685 185.720 ;
        RECT 42.855 185.705 43.865 185.875 ;
        RECT 41.425 184.985 42.655 185.155 ;
        RECT 39.585 184.175 41.255 184.945 ;
        RECT 41.700 184.380 41.945 184.985 ;
        RECT 42.165 184.175 42.675 184.710 ;
        RECT 42.855 184.345 43.045 185.705 ;
        RECT 43.215 185.365 43.490 185.505 ;
        RECT 43.215 185.195 43.495 185.365 ;
        RECT 43.215 184.345 43.490 185.195 ;
        RECT 43.695 184.905 43.865 185.705 ;
        RECT 44.035 184.915 44.205 186.045 ;
        RECT 44.375 185.415 44.545 186.385 ;
        RECT 44.715 185.585 44.885 186.725 ;
        RECT 45.055 185.585 45.390 186.555 ;
        RECT 44.375 185.085 44.570 185.415 ;
        RECT 44.795 185.085 45.050 185.415 ;
        RECT 44.795 184.915 44.965 185.085 ;
        RECT 45.220 184.915 45.390 185.585 ;
        RECT 46.485 185.635 49.995 186.725 ;
        RECT 46.485 185.115 48.175 185.635 ;
        RECT 50.165 185.560 50.455 186.725 ;
        RECT 50.625 185.650 50.895 186.555 ;
        RECT 51.065 185.965 51.395 186.725 ;
        RECT 51.575 185.795 51.745 186.555 ;
        RECT 48.345 184.945 49.995 185.465 ;
        RECT 44.035 184.745 44.965 184.915 ;
        RECT 44.035 184.710 44.210 184.745 ;
        RECT 43.680 184.345 44.210 184.710 ;
        RECT 44.635 184.175 44.965 184.575 ;
        RECT 45.135 184.345 45.390 184.915 ;
        RECT 46.485 184.175 49.995 184.945 ;
        RECT 50.165 184.175 50.455 184.900 ;
        RECT 50.625 184.850 50.795 185.650 ;
        RECT 51.080 185.625 51.745 185.795 ;
        RECT 52.840 185.745 53.095 186.415 ;
        RECT 53.275 185.925 53.560 186.725 ;
        RECT 53.740 186.005 54.070 186.515 ;
        RECT 51.080 185.480 51.250 185.625 ;
        RECT 50.965 185.150 51.250 185.480 ;
        RECT 51.080 184.895 51.250 185.150 ;
        RECT 51.485 185.075 51.815 185.445 ;
        RECT 50.625 184.345 50.885 184.850 ;
        RECT 51.080 184.725 51.745 184.895 ;
        RECT 51.065 184.175 51.395 184.555 ;
        RECT 51.575 184.345 51.745 184.725 ;
        RECT 52.840 184.885 53.020 185.745 ;
        RECT 53.740 185.415 53.990 186.005 ;
        RECT 54.340 185.855 54.510 186.465 ;
        RECT 54.680 186.035 55.010 186.725 ;
        RECT 55.240 186.175 55.480 186.465 ;
        RECT 55.680 186.345 56.100 186.725 ;
        RECT 56.280 186.255 56.910 186.505 ;
        RECT 57.380 186.345 57.710 186.725 ;
        RECT 56.280 186.175 56.450 186.255 ;
        RECT 57.880 186.175 58.050 186.465 ;
        RECT 58.230 186.345 58.610 186.725 ;
        RECT 58.850 186.340 59.680 186.510 ;
        RECT 55.240 186.005 56.450 186.175 ;
        RECT 53.190 185.085 53.990 185.415 ;
        RECT 52.840 184.685 53.095 184.885 ;
        RECT 52.755 184.515 53.095 184.685 ;
        RECT 52.840 184.355 53.095 184.515 ;
        RECT 53.275 184.175 53.560 184.635 ;
        RECT 53.740 184.435 53.990 185.085 ;
        RECT 54.190 185.835 54.510 185.855 ;
        RECT 54.190 185.665 56.110 185.835 ;
        RECT 54.190 184.770 54.380 185.665 ;
        RECT 56.280 185.495 56.450 186.005 ;
        RECT 56.620 185.745 57.140 186.055 ;
        RECT 54.550 185.325 56.450 185.495 ;
        RECT 54.550 185.265 54.880 185.325 ;
        RECT 55.030 185.095 55.360 185.155 ;
        RECT 54.700 184.825 55.360 185.095 ;
        RECT 54.190 184.440 54.510 184.770 ;
        RECT 54.690 184.175 55.350 184.655 ;
        RECT 55.550 184.565 55.720 185.325 ;
        RECT 56.620 185.155 56.800 185.565 ;
        RECT 55.890 184.985 56.220 185.105 ;
        RECT 56.970 184.985 57.140 185.745 ;
        RECT 55.890 184.815 57.140 184.985 ;
        RECT 57.310 185.925 58.680 186.175 ;
        RECT 57.310 185.155 57.500 185.925 ;
        RECT 58.430 185.665 58.680 185.925 ;
        RECT 57.670 185.495 57.920 185.655 ;
        RECT 58.850 185.495 59.020 186.340 ;
        RECT 59.915 186.055 60.085 186.555 ;
        RECT 60.255 186.225 60.585 186.725 ;
        RECT 59.190 185.665 59.690 186.045 ;
        RECT 59.915 185.885 60.610 186.055 ;
        RECT 57.670 185.325 59.020 185.495 ;
        RECT 58.600 185.285 59.020 185.325 ;
        RECT 57.310 184.815 57.730 185.155 ;
        RECT 58.020 184.825 58.430 185.155 ;
        RECT 55.550 184.395 56.400 184.565 ;
        RECT 56.960 184.175 57.280 184.635 ;
        RECT 57.480 184.385 57.730 184.815 ;
        RECT 58.020 184.175 58.430 184.615 ;
        RECT 58.600 184.555 58.770 185.285 ;
        RECT 58.940 184.735 59.290 185.105 ;
        RECT 59.470 184.795 59.690 185.665 ;
        RECT 59.860 185.095 60.270 185.715 ;
        RECT 60.440 184.915 60.610 185.885 ;
        RECT 59.915 184.725 60.610 184.915 ;
        RECT 58.600 184.355 59.615 184.555 ;
        RECT 59.915 184.395 60.085 184.725 ;
        RECT 60.255 184.175 60.585 184.555 ;
        RECT 60.800 184.435 61.025 186.555 ;
        RECT 61.195 186.225 61.525 186.725 ;
        RECT 61.695 186.055 61.865 186.555 ;
        RECT 61.200 185.885 61.865 186.055 ;
        RECT 63.130 186.105 63.305 186.555 ;
        RECT 63.475 186.285 63.805 186.725 ;
        RECT 64.110 186.135 64.280 186.555 ;
        RECT 64.515 186.315 65.185 186.725 ;
        RECT 65.400 186.135 65.570 186.555 ;
        RECT 65.770 186.315 66.100 186.725 ;
        RECT 63.130 185.935 63.760 186.105 ;
        RECT 61.200 184.895 61.430 185.885 ;
        RECT 61.600 185.065 61.950 185.715 ;
        RECT 63.045 185.085 63.410 185.765 ;
        RECT 63.590 185.415 63.760 185.935 ;
        RECT 64.110 185.965 66.125 186.135 ;
        RECT 63.590 185.085 63.940 185.415 ;
        RECT 63.590 184.915 63.760 185.085 ;
        RECT 61.200 184.725 61.865 184.895 ;
        RECT 61.195 184.175 61.525 184.555 ;
        RECT 61.695 184.435 61.865 184.725 ;
        RECT 63.130 184.745 63.760 184.915 ;
        RECT 63.130 184.345 63.305 184.745 ;
        RECT 64.110 184.675 64.280 185.965 ;
        RECT 63.475 184.175 63.805 184.555 ;
        RECT 64.050 184.345 64.280 184.675 ;
        RECT 64.480 184.510 64.760 185.785 ;
        RECT 64.985 184.685 65.255 185.785 ;
        RECT 65.445 184.755 65.785 185.785 ;
        RECT 65.955 185.415 66.125 185.965 ;
        RECT 66.295 185.585 66.555 186.555 ;
        RECT 65.955 185.085 66.215 185.415 ;
        RECT 66.385 184.895 66.555 185.585 ;
        RECT 64.945 184.515 65.255 184.685 ;
        RECT 64.985 184.510 65.255 184.515 ;
        RECT 65.715 184.175 66.045 184.555 ;
        RECT 66.215 184.430 66.555 184.895 ;
        RECT 66.730 185.535 66.985 186.415 ;
        RECT 67.155 185.585 67.460 186.725 ;
        RECT 67.800 186.345 68.130 186.725 ;
        RECT 68.310 186.175 68.480 186.465 ;
        RECT 68.650 186.265 68.900 186.725 ;
        RECT 67.680 186.005 68.480 186.175 ;
        RECT 69.070 186.215 69.940 186.555 ;
        RECT 66.730 184.885 66.940 185.535 ;
        RECT 67.680 185.415 67.850 186.005 ;
        RECT 69.070 185.835 69.240 186.215 ;
        RECT 70.175 186.095 70.345 186.555 ;
        RECT 70.515 186.265 70.885 186.725 ;
        RECT 71.180 186.125 71.350 186.465 ;
        RECT 71.520 186.295 71.850 186.725 ;
        RECT 72.085 186.125 72.255 186.465 ;
        RECT 68.020 185.665 69.240 185.835 ;
        RECT 69.410 185.755 69.870 186.045 ;
        RECT 70.175 185.925 70.735 186.095 ;
        RECT 71.180 185.955 72.255 186.125 ;
        RECT 72.425 186.225 73.105 186.555 ;
        RECT 73.320 186.225 73.570 186.555 ;
        RECT 73.740 186.265 73.990 186.725 ;
        RECT 70.565 185.785 70.735 185.925 ;
        RECT 69.410 185.745 70.375 185.755 ;
        RECT 69.070 185.575 69.240 185.665 ;
        RECT 69.700 185.585 70.375 185.745 ;
        RECT 67.110 185.385 67.850 185.415 ;
        RECT 67.110 185.085 68.025 185.385 ;
        RECT 67.700 184.910 68.025 185.085 ;
        RECT 66.215 184.385 66.550 184.430 ;
        RECT 66.730 184.355 66.985 184.885 ;
        RECT 67.155 184.175 67.460 184.635 ;
        RECT 67.705 184.555 68.025 184.910 ;
        RECT 68.195 185.125 68.735 185.495 ;
        RECT 69.070 185.405 69.475 185.575 ;
        RECT 68.195 184.725 68.435 185.125 ;
        RECT 68.915 184.955 69.135 185.235 ;
        RECT 68.605 184.785 69.135 184.955 ;
        RECT 68.605 184.555 68.775 184.785 ;
        RECT 69.305 184.625 69.475 185.405 ;
        RECT 69.645 184.795 69.995 185.415 ;
        RECT 70.165 184.795 70.375 185.585 ;
        RECT 70.565 185.615 72.065 185.785 ;
        RECT 70.565 184.925 70.735 185.615 ;
        RECT 72.425 185.445 72.595 186.225 ;
        RECT 73.400 186.095 73.570 186.225 ;
        RECT 70.905 185.275 72.595 185.445 ;
        RECT 72.765 185.665 73.230 186.055 ;
        RECT 73.400 185.925 73.795 186.095 ;
        RECT 70.905 185.095 71.075 185.275 ;
        RECT 67.705 184.385 68.775 184.555 ;
        RECT 68.945 184.175 69.135 184.615 ;
        RECT 69.305 184.345 70.255 184.625 ;
        RECT 70.565 184.535 70.825 184.925 ;
        RECT 71.245 184.855 72.035 185.105 ;
        RECT 70.475 184.365 70.825 184.535 ;
        RECT 71.035 184.175 71.365 184.635 ;
        RECT 72.240 184.565 72.410 185.275 ;
        RECT 72.765 185.075 72.935 185.665 ;
        RECT 72.580 184.855 72.935 185.075 ;
        RECT 73.105 184.855 73.455 185.475 ;
        RECT 73.625 184.565 73.795 185.925 ;
        RECT 74.160 185.755 74.485 186.540 ;
        RECT 73.965 184.705 74.425 185.755 ;
        RECT 72.240 184.395 73.095 184.565 ;
        RECT 73.300 184.395 73.795 184.565 ;
        RECT 73.965 184.175 74.295 184.535 ;
        RECT 74.655 184.435 74.825 186.555 ;
        RECT 74.995 186.225 75.325 186.725 ;
        RECT 75.495 186.055 75.750 186.555 ;
        RECT 75.000 185.885 75.750 186.055 ;
        RECT 75.000 184.895 75.230 185.885 ;
        RECT 75.400 185.065 75.750 185.715 ;
        RECT 75.925 185.560 76.215 186.725 ;
        RECT 76.385 185.635 77.595 186.725 ;
        RECT 77.765 185.635 81.275 186.725 ;
        RECT 76.385 185.095 76.905 185.635 ;
        RECT 77.075 184.925 77.595 185.465 ;
        RECT 77.765 185.115 79.455 185.635 ;
        RECT 81.505 185.585 81.715 186.725 ;
        RECT 81.885 185.575 82.215 186.555 ;
        RECT 82.385 185.585 82.615 186.725 ;
        RECT 82.825 185.965 83.340 186.375 ;
        RECT 83.575 185.965 83.745 186.725 ;
        RECT 83.915 186.385 85.945 186.555 ;
        RECT 79.625 184.945 81.275 185.465 ;
        RECT 75.000 184.725 75.750 184.895 ;
        RECT 74.995 184.175 75.325 184.555 ;
        RECT 75.495 184.435 75.750 184.725 ;
        RECT 75.925 184.175 76.215 184.900 ;
        RECT 76.385 184.175 77.595 184.925 ;
        RECT 77.765 184.175 81.275 184.945 ;
        RECT 81.505 184.175 81.715 184.995 ;
        RECT 81.885 184.975 82.135 185.575 ;
        RECT 82.305 185.165 82.635 185.415 ;
        RECT 82.825 185.155 83.165 185.965 ;
        RECT 83.915 185.720 84.085 186.385 ;
        RECT 84.480 186.045 85.605 186.215 ;
        RECT 83.335 185.530 84.085 185.720 ;
        RECT 84.255 185.705 85.265 185.875 ;
        RECT 81.885 184.345 82.215 184.975 ;
        RECT 82.385 184.175 82.615 184.995 ;
        RECT 82.825 184.985 84.055 185.155 ;
        RECT 83.100 184.380 83.345 184.985 ;
        RECT 83.565 184.175 84.075 184.710 ;
        RECT 84.255 184.345 84.445 185.705 ;
        RECT 84.615 185.025 84.890 185.505 ;
        RECT 84.615 184.855 84.895 185.025 ;
        RECT 85.095 184.905 85.265 185.705 ;
        RECT 85.435 184.915 85.605 186.045 ;
        RECT 85.775 185.415 85.945 186.385 ;
        RECT 86.115 185.585 86.285 186.725 ;
        RECT 86.455 185.585 86.790 186.555 ;
        RECT 85.775 185.085 85.970 185.415 ;
        RECT 86.195 185.085 86.450 185.415 ;
        RECT 86.195 184.915 86.365 185.085 ;
        RECT 86.620 184.915 86.790 185.585 ;
        RECT 86.965 185.635 88.175 186.725 ;
        RECT 88.345 185.635 91.855 186.725 ;
        RECT 92.030 186.290 97.375 186.725 ;
        RECT 86.965 185.095 87.485 185.635 ;
        RECT 87.655 184.925 88.175 185.465 ;
        RECT 88.345 185.115 90.035 185.635 ;
        RECT 90.205 184.945 91.855 185.465 ;
        RECT 93.620 185.040 93.970 186.290 ;
        RECT 97.545 185.965 98.060 186.375 ;
        RECT 98.295 185.965 98.465 186.725 ;
        RECT 98.635 186.385 100.665 186.555 ;
        RECT 84.615 184.345 84.890 184.855 ;
        RECT 85.435 184.745 86.365 184.915 ;
        RECT 85.435 184.710 85.610 184.745 ;
        RECT 85.080 184.345 85.610 184.710 ;
        RECT 86.035 184.175 86.365 184.575 ;
        RECT 86.535 184.345 86.790 184.915 ;
        RECT 86.965 184.175 88.175 184.925 ;
        RECT 88.345 184.175 91.855 184.945 ;
        RECT 95.450 184.720 95.790 185.550 ;
        RECT 97.545 185.155 97.885 185.965 ;
        RECT 98.635 185.720 98.805 186.385 ;
        RECT 99.200 186.045 100.325 186.215 ;
        RECT 98.055 185.530 98.805 185.720 ;
        RECT 98.975 185.705 99.985 185.875 ;
        RECT 97.545 184.985 98.775 185.155 ;
        RECT 92.030 184.175 97.375 184.720 ;
        RECT 97.820 184.380 98.065 184.985 ;
        RECT 98.285 184.175 98.795 184.710 ;
        RECT 98.975 184.345 99.165 185.705 ;
        RECT 99.335 185.365 99.610 185.505 ;
        RECT 99.335 185.195 99.615 185.365 ;
        RECT 99.335 184.345 99.610 185.195 ;
        RECT 99.815 184.905 99.985 185.705 ;
        RECT 100.155 184.915 100.325 186.045 ;
        RECT 100.495 185.415 100.665 186.385 ;
        RECT 100.835 185.585 101.005 186.725 ;
        RECT 101.175 185.585 101.510 186.555 ;
        RECT 100.495 185.085 100.690 185.415 ;
        RECT 100.915 185.085 101.170 185.415 ;
        RECT 100.915 184.915 101.085 185.085 ;
        RECT 101.340 184.915 101.510 185.585 ;
        RECT 101.685 185.560 101.975 186.725 ;
        RECT 102.605 185.965 103.120 186.375 ;
        RECT 103.355 185.965 103.525 186.725 ;
        RECT 103.695 186.385 105.725 186.555 ;
        RECT 102.605 185.155 102.945 185.965 ;
        RECT 103.695 185.720 103.865 186.385 ;
        RECT 104.260 186.045 105.385 186.215 ;
        RECT 103.115 185.530 103.865 185.720 ;
        RECT 104.035 185.705 105.045 185.875 ;
        RECT 102.605 184.985 103.835 185.155 ;
        RECT 100.155 184.745 101.085 184.915 ;
        RECT 100.155 184.710 100.330 184.745 ;
        RECT 99.800 184.345 100.330 184.710 ;
        RECT 100.755 184.175 101.085 184.575 ;
        RECT 101.255 184.345 101.510 184.915 ;
        RECT 101.685 184.175 101.975 184.900 ;
        RECT 102.880 184.380 103.125 184.985 ;
        RECT 103.345 184.175 103.855 184.710 ;
        RECT 104.035 184.345 104.225 185.705 ;
        RECT 104.395 184.685 104.670 185.505 ;
        RECT 104.875 184.905 105.045 185.705 ;
        RECT 105.215 184.915 105.385 186.045 ;
        RECT 105.555 185.415 105.725 186.385 ;
        RECT 105.895 185.585 106.065 186.725 ;
        RECT 106.235 185.585 106.570 186.555 ;
        RECT 106.805 185.585 107.015 186.725 ;
        RECT 105.555 185.085 105.750 185.415 ;
        RECT 105.975 185.085 106.230 185.415 ;
        RECT 105.975 184.915 106.145 185.085 ;
        RECT 106.400 184.915 106.570 185.585 ;
        RECT 107.185 185.575 107.515 186.555 ;
        RECT 107.685 185.585 107.915 186.725 ;
        RECT 108.125 185.650 108.395 186.555 ;
        RECT 108.565 185.965 108.895 186.725 ;
        RECT 109.075 185.795 109.245 186.555 ;
        RECT 105.215 184.745 106.145 184.915 ;
        RECT 105.215 184.710 105.390 184.745 ;
        RECT 104.395 184.515 104.675 184.685 ;
        RECT 104.395 184.345 104.670 184.515 ;
        RECT 104.860 184.345 105.390 184.710 ;
        RECT 105.815 184.175 106.145 184.575 ;
        RECT 106.315 184.345 106.570 184.915 ;
        RECT 106.805 184.175 107.015 184.995 ;
        RECT 107.185 184.975 107.435 185.575 ;
        RECT 107.605 185.165 107.935 185.415 ;
        RECT 107.185 184.345 107.515 184.975 ;
        RECT 107.685 184.175 107.915 184.995 ;
        RECT 108.125 184.850 108.295 185.650 ;
        RECT 108.580 185.625 109.245 185.795 ;
        RECT 109.965 185.635 113.475 186.725 ;
        RECT 108.580 185.480 108.750 185.625 ;
        RECT 108.465 185.150 108.750 185.480 ;
        RECT 108.580 184.895 108.750 185.150 ;
        RECT 108.985 185.075 109.315 185.445 ;
        RECT 109.965 185.115 111.655 185.635 ;
        RECT 113.685 185.585 113.915 186.725 ;
        RECT 114.085 185.575 114.415 186.555 ;
        RECT 114.585 185.585 114.795 186.725 ;
        RECT 111.825 184.945 113.475 185.465 ;
        RECT 113.665 185.165 113.995 185.415 ;
        RECT 108.125 184.345 108.385 184.850 ;
        RECT 108.580 184.725 109.245 184.895 ;
        RECT 108.565 184.175 108.895 184.555 ;
        RECT 109.075 184.345 109.245 184.725 ;
        RECT 109.965 184.175 113.475 184.945 ;
        RECT 113.685 184.175 113.915 184.995 ;
        RECT 114.165 184.975 114.415 185.575 ;
        RECT 115.030 185.535 115.285 186.415 ;
        RECT 115.455 185.585 115.760 186.725 ;
        RECT 116.100 186.345 116.430 186.725 ;
        RECT 116.610 186.175 116.780 186.465 ;
        RECT 116.950 186.265 117.200 186.725 ;
        RECT 115.980 186.005 116.780 186.175 ;
        RECT 117.370 186.215 118.240 186.555 ;
        RECT 114.085 184.345 114.415 184.975 ;
        RECT 114.585 184.175 114.795 184.995 ;
        RECT 115.030 184.885 115.240 185.535 ;
        RECT 115.980 185.415 116.150 186.005 ;
        RECT 117.370 185.835 117.540 186.215 ;
        RECT 118.475 186.095 118.645 186.555 ;
        RECT 118.815 186.265 119.185 186.725 ;
        RECT 119.480 186.125 119.650 186.465 ;
        RECT 119.820 186.295 120.150 186.725 ;
        RECT 120.385 186.125 120.555 186.465 ;
        RECT 116.320 185.665 117.540 185.835 ;
        RECT 117.710 185.755 118.170 186.045 ;
        RECT 118.475 185.925 119.035 186.095 ;
        RECT 119.480 185.955 120.555 186.125 ;
        RECT 120.725 186.225 121.405 186.555 ;
        RECT 121.620 186.225 121.870 186.555 ;
        RECT 122.040 186.265 122.290 186.725 ;
        RECT 118.865 185.785 119.035 185.925 ;
        RECT 117.710 185.745 118.675 185.755 ;
        RECT 117.370 185.575 117.540 185.665 ;
        RECT 118.000 185.585 118.675 185.745 ;
        RECT 115.410 185.385 116.150 185.415 ;
        RECT 115.410 185.085 116.325 185.385 ;
        RECT 116.000 184.910 116.325 185.085 ;
        RECT 115.030 184.355 115.285 184.885 ;
        RECT 115.455 184.175 115.760 184.635 ;
        RECT 116.005 184.555 116.325 184.910 ;
        RECT 116.495 185.125 117.035 185.495 ;
        RECT 117.370 185.405 117.775 185.575 ;
        RECT 116.495 184.725 116.735 185.125 ;
        RECT 117.215 184.955 117.435 185.235 ;
        RECT 116.905 184.785 117.435 184.955 ;
        RECT 116.905 184.555 117.075 184.785 ;
        RECT 117.605 184.625 117.775 185.405 ;
        RECT 117.945 184.795 118.295 185.415 ;
        RECT 118.465 184.795 118.675 185.585 ;
        RECT 118.865 185.615 120.365 185.785 ;
        RECT 118.865 184.925 119.035 185.615 ;
        RECT 120.725 185.445 120.895 186.225 ;
        RECT 121.700 186.095 121.870 186.225 ;
        RECT 119.205 185.275 120.895 185.445 ;
        RECT 121.065 185.665 121.530 186.055 ;
        RECT 121.700 185.925 122.095 186.095 ;
        RECT 119.205 185.095 119.375 185.275 ;
        RECT 116.005 184.385 117.075 184.555 ;
        RECT 117.245 184.175 117.435 184.615 ;
        RECT 117.605 184.345 118.555 184.625 ;
        RECT 118.865 184.535 119.125 184.925 ;
        RECT 119.545 184.855 120.335 185.105 ;
        RECT 118.775 184.365 119.125 184.535 ;
        RECT 119.335 184.175 119.665 184.635 ;
        RECT 120.540 184.565 120.710 185.275 ;
        RECT 121.065 185.075 121.235 185.665 ;
        RECT 120.880 184.855 121.235 185.075 ;
        RECT 121.405 184.855 121.755 185.475 ;
        RECT 121.925 184.565 122.095 185.925 ;
        RECT 122.460 185.755 122.785 186.540 ;
        RECT 122.265 184.705 122.725 185.755 ;
        RECT 120.540 184.395 121.395 184.565 ;
        RECT 121.600 184.395 122.095 184.565 ;
        RECT 122.265 184.175 122.595 184.535 ;
        RECT 122.955 184.435 123.125 186.555 ;
        RECT 123.295 186.225 123.625 186.725 ;
        RECT 123.795 186.055 124.050 186.555 ;
        RECT 123.300 185.885 124.050 186.055 ;
        RECT 123.300 184.895 123.530 185.885 ;
        RECT 123.700 185.065 124.050 185.715 ;
        RECT 124.225 185.650 124.495 186.555 ;
        RECT 124.665 185.965 124.995 186.725 ;
        RECT 125.175 185.795 125.345 186.555 ;
        RECT 123.300 184.725 124.050 184.895 ;
        RECT 123.295 184.175 123.625 184.555 ;
        RECT 123.795 184.435 124.050 184.725 ;
        RECT 124.225 184.850 124.395 185.650 ;
        RECT 124.680 185.625 125.345 185.795 ;
        RECT 126.525 185.635 127.735 186.725 ;
        RECT 124.680 185.480 124.850 185.625 ;
        RECT 124.565 185.150 124.850 185.480 ;
        RECT 124.680 184.895 124.850 185.150 ;
        RECT 125.085 185.075 125.415 185.445 ;
        RECT 126.525 185.095 127.045 185.635 ;
        RECT 127.215 184.925 127.735 185.465 ;
        RECT 124.225 184.345 124.485 184.850 ;
        RECT 124.680 184.725 125.345 184.895 ;
        RECT 124.665 184.175 124.995 184.555 ;
        RECT 125.175 184.345 125.345 184.725 ;
        RECT 126.525 184.175 127.735 184.925 ;
        RECT 14.660 184.005 127.820 184.175 ;
        RECT 14.745 183.255 15.955 184.005 ;
        RECT 17.050 183.460 22.395 184.005 ;
        RECT 22.570 183.460 27.915 184.005 ;
        RECT 14.745 182.715 15.265 183.255 ;
        RECT 15.435 182.545 15.955 183.085 ;
        RECT 14.745 181.455 15.955 182.545 ;
        RECT 18.640 181.890 18.990 183.140 ;
        RECT 20.470 182.630 20.810 183.460 ;
        RECT 24.160 181.890 24.510 183.140 ;
        RECT 25.990 182.630 26.330 183.460 ;
        RECT 28.090 183.295 28.345 183.825 ;
        RECT 28.515 183.545 28.820 184.005 ;
        RECT 29.065 183.625 30.135 183.795 ;
        RECT 28.090 182.645 28.300 183.295 ;
        RECT 29.065 183.270 29.385 183.625 ;
        RECT 29.060 183.095 29.385 183.270 ;
        RECT 28.470 182.795 29.385 183.095 ;
        RECT 29.555 183.055 29.795 183.455 ;
        RECT 29.965 183.395 30.135 183.625 ;
        RECT 30.305 183.565 30.495 184.005 ;
        RECT 30.665 183.555 31.615 183.835 ;
        RECT 31.835 183.645 32.185 183.815 ;
        RECT 29.965 183.225 30.495 183.395 ;
        RECT 28.470 182.765 29.210 182.795 ;
        RECT 17.050 181.455 22.395 181.890 ;
        RECT 22.570 181.455 27.915 181.890 ;
        RECT 28.090 181.765 28.345 182.645 ;
        RECT 28.515 181.455 28.820 182.595 ;
        RECT 29.040 182.175 29.210 182.765 ;
        RECT 29.555 182.685 30.095 183.055 ;
        RECT 30.275 182.945 30.495 183.225 ;
        RECT 30.665 182.775 30.835 183.555 ;
        RECT 30.430 182.605 30.835 182.775 ;
        RECT 31.005 182.765 31.355 183.385 ;
        RECT 30.430 182.515 30.600 182.605 ;
        RECT 31.525 182.595 31.735 183.385 ;
        RECT 29.380 182.345 30.600 182.515 ;
        RECT 31.060 182.435 31.735 182.595 ;
        RECT 29.040 182.005 29.840 182.175 ;
        RECT 29.160 181.455 29.490 181.835 ;
        RECT 29.670 181.715 29.840 182.005 ;
        RECT 30.430 181.965 30.600 182.345 ;
        RECT 30.770 182.425 31.735 182.435 ;
        RECT 31.925 183.255 32.185 183.645 ;
        RECT 32.395 183.545 32.725 184.005 ;
        RECT 33.600 183.615 34.455 183.785 ;
        RECT 34.660 183.615 35.155 183.785 ;
        RECT 35.325 183.645 35.655 184.005 ;
        RECT 31.925 182.565 32.095 183.255 ;
        RECT 32.265 182.905 32.435 183.085 ;
        RECT 32.605 183.075 33.395 183.325 ;
        RECT 33.600 182.905 33.770 183.615 ;
        RECT 33.940 183.105 34.295 183.325 ;
        RECT 32.265 182.735 33.955 182.905 ;
        RECT 30.770 182.135 31.230 182.425 ;
        RECT 31.925 182.395 33.425 182.565 ;
        RECT 31.925 182.255 32.095 182.395 ;
        RECT 31.535 182.085 32.095 182.255 ;
        RECT 30.010 181.455 30.260 181.915 ;
        RECT 30.430 181.625 31.300 181.965 ;
        RECT 31.535 181.625 31.705 182.085 ;
        RECT 32.540 182.055 33.615 182.225 ;
        RECT 31.875 181.455 32.245 181.915 ;
        RECT 32.540 181.715 32.710 182.055 ;
        RECT 32.880 181.455 33.210 181.885 ;
        RECT 33.445 181.715 33.615 182.055 ;
        RECT 33.785 181.955 33.955 182.735 ;
        RECT 34.125 182.515 34.295 183.105 ;
        RECT 34.465 182.705 34.815 183.325 ;
        RECT 34.125 182.125 34.590 182.515 ;
        RECT 34.985 182.255 35.155 183.615 ;
        RECT 35.325 182.425 35.785 183.475 ;
        RECT 34.760 182.085 35.155 182.255 ;
        RECT 34.760 181.955 34.930 182.085 ;
        RECT 33.785 181.625 34.465 181.955 ;
        RECT 34.680 181.625 34.930 181.955 ;
        RECT 35.100 181.455 35.350 181.915 ;
        RECT 35.520 181.640 35.845 182.425 ;
        RECT 36.015 181.625 36.185 183.745 ;
        RECT 36.355 183.625 36.685 184.005 ;
        RECT 36.855 183.455 37.110 183.745 ;
        RECT 36.360 183.285 37.110 183.455 ;
        RECT 36.360 182.295 36.590 183.285 ;
        RECT 37.285 183.280 37.575 184.005 ;
        RECT 37.750 183.295 38.005 183.825 ;
        RECT 38.175 183.545 38.480 184.005 ;
        RECT 38.725 183.625 39.795 183.795 ;
        RECT 36.760 182.465 37.110 183.115 ;
        RECT 37.750 182.645 37.960 183.295 ;
        RECT 38.725 183.270 39.045 183.625 ;
        RECT 38.720 183.095 39.045 183.270 ;
        RECT 38.130 182.795 39.045 183.095 ;
        RECT 39.215 183.055 39.455 183.455 ;
        RECT 39.625 183.395 39.795 183.625 ;
        RECT 39.965 183.565 40.155 184.005 ;
        RECT 40.325 183.555 41.275 183.835 ;
        RECT 41.495 183.645 41.845 183.815 ;
        RECT 39.625 183.225 40.155 183.395 ;
        RECT 38.130 182.765 38.870 182.795 ;
        RECT 36.360 182.125 37.110 182.295 ;
        RECT 36.355 181.455 36.685 181.955 ;
        RECT 36.855 181.625 37.110 182.125 ;
        RECT 37.285 181.455 37.575 182.620 ;
        RECT 37.750 181.765 38.005 182.645 ;
        RECT 38.175 181.455 38.480 182.595 ;
        RECT 38.700 182.175 38.870 182.765 ;
        RECT 39.215 182.685 39.755 183.055 ;
        RECT 39.935 182.945 40.155 183.225 ;
        RECT 40.325 182.775 40.495 183.555 ;
        RECT 40.090 182.605 40.495 182.775 ;
        RECT 40.665 182.765 41.015 183.385 ;
        RECT 40.090 182.515 40.260 182.605 ;
        RECT 41.185 182.595 41.395 183.385 ;
        RECT 39.040 182.345 40.260 182.515 ;
        RECT 40.720 182.435 41.395 182.595 ;
        RECT 38.700 182.005 39.500 182.175 ;
        RECT 38.820 181.455 39.150 181.835 ;
        RECT 39.330 181.715 39.500 182.005 ;
        RECT 40.090 181.965 40.260 182.345 ;
        RECT 40.430 182.425 41.395 182.435 ;
        RECT 41.585 183.255 41.845 183.645 ;
        RECT 42.055 183.545 42.385 184.005 ;
        RECT 43.260 183.615 44.115 183.785 ;
        RECT 44.320 183.615 44.815 183.785 ;
        RECT 44.985 183.645 45.315 184.005 ;
        RECT 41.585 182.565 41.755 183.255 ;
        RECT 41.925 182.905 42.095 183.085 ;
        RECT 42.265 183.075 43.055 183.325 ;
        RECT 43.260 182.905 43.430 183.615 ;
        RECT 43.600 183.105 43.955 183.325 ;
        RECT 41.925 182.735 43.615 182.905 ;
        RECT 40.430 182.135 40.890 182.425 ;
        RECT 41.585 182.395 43.085 182.565 ;
        RECT 41.585 182.255 41.755 182.395 ;
        RECT 41.195 182.085 41.755 182.255 ;
        RECT 39.670 181.455 39.920 181.915 ;
        RECT 40.090 181.625 40.960 181.965 ;
        RECT 41.195 181.625 41.365 182.085 ;
        RECT 42.200 182.055 43.275 182.225 ;
        RECT 41.535 181.455 41.905 181.915 ;
        RECT 42.200 181.715 42.370 182.055 ;
        RECT 42.540 181.455 42.870 181.885 ;
        RECT 43.105 181.715 43.275 182.055 ;
        RECT 43.445 181.955 43.615 182.735 ;
        RECT 43.785 182.515 43.955 183.105 ;
        RECT 44.125 182.705 44.475 183.325 ;
        RECT 43.785 182.125 44.250 182.515 ;
        RECT 44.645 182.255 44.815 183.615 ;
        RECT 44.985 182.425 45.445 183.475 ;
        RECT 44.420 182.085 44.815 182.255 ;
        RECT 44.420 181.955 44.590 182.085 ;
        RECT 43.445 181.625 44.125 181.955 ;
        RECT 44.340 181.625 44.590 181.955 ;
        RECT 44.760 181.455 45.010 181.915 ;
        RECT 45.180 181.640 45.505 182.425 ;
        RECT 45.675 181.625 45.845 183.745 ;
        RECT 46.015 183.625 46.345 184.005 ;
        RECT 46.515 183.455 46.770 183.745 ;
        RECT 46.950 183.460 52.295 184.005 ;
        RECT 52.470 183.460 57.815 184.005 ;
        RECT 46.020 183.285 46.770 183.455 ;
        RECT 46.020 182.295 46.250 183.285 ;
        RECT 46.420 182.465 46.770 183.115 ;
        RECT 46.020 182.125 46.770 182.295 ;
        RECT 46.015 181.455 46.345 181.955 ;
        RECT 46.515 181.625 46.770 182.125 ;
        RECT 48.540 181.890 48.890 183.140 ;
        RECT 50.370 182.630 50.710 183.460 ;
        RECT 54.060 181.890 54.410 183.140 ;
        RECT 55.890 182.630 56.230 183.460 ;
        RECT 58.075 183.455 58.245 183.835 ;
        RECT 58.425 183.625 58.755 184.005 ;
        RECT 58.075 183.285 58.740 183.455 ;
        RECT 58.935 183.330 59.195 183.835 ;
        RECT 58.005 182.735 58.335 183.105 ;
        RECT 58.570 183.030 58.740 183.285 ;
        RECT 58.570 182.700 58.855 183.030 ;
        RECT 58.570 182.555 58.740 182.700 ;
        RECT 58.075 182.385 58.740 182.555 ;
        RECT 59.025 182.530 59.195 183.330 ;
        RECT 59.365 183.235 62.875 184.005 ;
        RECT 63.045 183.280 63.335 184.005 ;
        RECT 63.505 183.235 65.175 184.005 ;
        RECT 65.435 183.455 65.605 183.835 ;
        RECT 65.820 183.625 66.150 184.005 ;
        RECT 65.435 183.285 66.150 183.455 ;
        RECT 46.950 181.455 52.295 181.890 ;
        RECT 52.470 181.455 57.815 181.890 ;
        RECT 58.075 181.625 58.245 182.385 ;
        RECT 58.425 181.455 58.755 182.215 ;
        RECT 58.925 181.625 59.195 182.530 ;
        RECT 59.365 182.545 61.055 183.065 ;
        RECT 61.225 182.715 62.875 183.235 ;
        RECT 59.365 181.455 62.875 182.545 ;
        RECT 63.045 181.455 63.335 182.620 ;
        RECT 63.505 182.545 64.255 183.065 ;
        RECT 64.425 182.715 65.175 183.235 ;
        RECT 65.345 182.735 65.700 183.105 ;
        RECT 65.980 183.095 66.150 183.285 ;
        RECT 66.320 183.260 66.575 183.835 ;
        RECT 65.980 182.765 66.235 183.095 ;
        RECT 65.980 182.555 66.150 182.765 ;
        RECT 63.505 181.455 65.175 182.545 ;
        RECT 65.435 182.385 66.150 182.555 ;
        RECT 66.405 182.530 66.575 183.260 ;
        RECT 66.750 183.165 67.010 184.005 ;
        RECT 65.435 181.625 65.605 182.385 ;
        RECT 65.820 181.455 66.150 182.215 ;
        RECT 66.320 181.625 66.575 182.530 ;
        RECT 66.750 181.455 67.010 182.605 ;
        RECT 67.185 181.625 67.445 183.835 ;
        RECT 67.615 183.625 67.945 184.005 ;
        RECT 68.155 183.095 68.350 183.670 ;
        RECT 68.620 183.095 68.805 183.675 ;
        RECT 67.615 182.175 67.785 183.095 ;
        RECT 68.095 182.765 68.350 183.095 ;
        RECT 68.575 182.765 68.805 183.095 ;
        RECT 69.055 183.665 70.535 183.835 ;
        RECT 69.055 182.765 69.225 183.665 ;
        RECT 69.395 183.165 69.945 183.495 ;
        RECT 70.135 183.335 70.535 183.665 ;
        RECT 70.715 183.625 71.045 184.005 ;
        RECT 71.355 183.505 71.615 183.835 ;
        RECT 68.155 182.455 68.350 182.765 ;
        RECT 68.620 182.455 68.805 182.765 ;
        RECT 69.395 182.175 69.565 183.165 ;
        RECT 70.135 182.855 70.305 183.335 ;
        RECT 70.885 183.145 71.095 183.325 ;
        RECT 70.475 182.975 71.095 183.145 ;
        RECT 67.615 182.005 69.565 182.175 ;
        RECT 69.735 182.685 70.305 182.855 ;
        RECT 71.445 182.805 71.615 183.505 ;
        RECT 72.245 183.235 74.835 184.005 ;
        RECT 69.735 182.175 69.905 182.685 ;
        RECT 70.485 182.635 71.615 182.805 ;
        RECT 70.485 182.515 70.655 182.635 ;
        RECT 70.075 182.345 70.655 182.515 ;
        RECT 69.735 182.005 70.475 182.175 ;
        RECT 70.925 182.135 71.275 182.465 ;
        RECT 67.615 181.455 67.945 181.835 ;
        RECT 68.370 181.625 68.540 182.005 ;
        RECT 68.800 181.455 69.130 181.835 ;
        RECT 69.325 181.625 69.495 182.005 ;
        RECT 69.705 181.455 70.035 181.835 ;
        RECT 70.285 181.625 70.475 182.005 ;
        RECT 71.445 181.955 71.615 182.635 ;
        RECT 70.715 181.455 71.045 181.835 ;
        RECT 71.355 181.625 71.615 181.955 ;
        RECT 72.245 182.545 73.455 183.065 ;
        RECT 73.625 182.715 74.835 183.235 ;
        RECT 75.095 183.355 75.265 183.835 ;
        RECT 75.445 183.525 75.685 184.005 ;
        RECT 75.935 183.355 76.105 183.835 ;
        RECT 76.275 183.525 76.605 184.005 ;
        RECT 76.775 183.355 76.945 183.835 ;
        RECT 75.095 183.185 75.730 183.355 ;
        RECT 75.935 183.185 76.945 183.355 ;
        RECT 77.115 183.205 77.445 184.005 ;
        RECT 78.690 183.295 78.945 183.825 ;
        RECT 79.115 183.545 79.420 184.005 ;
        RECT 79.665 183.625 80.735 183.795 ;
        RECT 75.560 183.015 75.730 183.185 ;
        RECT 76.445 183.155 76.945 183.185 ;
        RECT 75.010 182.775 75.390 183.015 ;
        RECT 75.560 182.845 76.060 183.015 ;
        RECT 75.560 182.605 75.730 182.845 ;
        RECT 76.450 182.645 76.945 183.155 ;
        RECT 72.245 181.455 74.835 182.545 ;
        RECT 75.015 182.435 75.730 182.605 ;
        RECT 75.935 182.475 76.945 182.645 ;
        RECT 78.690 182.645 78.900 183.295 ;
        RECT 79.665 183.270 79.985 183.625 ;
        RECT 79.660 183.095 79.985 183.270 ;
        RECT 79.070 182.795 79.985 183.095 ;
        RECT 80.155 183.055 80.395 183.455 ;
        RECT 80.565 183.395 80.735 183.625 ;
        RECT 80.905 183.565 81.095 184.005 ;
        RECT 81.265 183.555 82.215 183.835 ;
        RECT 82.435 183.645 82.785 183.815 ;
        RECT 80.565 183.225 81.095 183.395 ;
        RECT 79.070 182.765 79.810 182.795 ;
        RECT 75.015 181.625 75.345 182.435 ;
        RECT 75.515 181.455 75.755 182.255 ;
        RECT 75.935 181.625 76.105 182.475 ;
        RECT 76.275 181.455 76.605 182.255 ;
        RECT 76.775 181.625 76.945 182.475 ;
        RECT 77.115 181.455 77.445 182.605 ;
        RECT 78.690 181.765 78.945 182.645 ;
        RECT 79.115 181.455 79.420 182.595 ;
        RECT 79.640 182.175 79.810 182.765 ;
        RECT 80.155 182.685 80.695 183.055 ;
        RECT 80.875 182.945 81.095 183.225 ;
        RECT 81.265 182.775 81.435 183.555 ;
        RECT 81.030 182.605 81.435 182.775 ;
        RECT 81.605 182.765 81.955 183.385 ;
        RECT 81.030 182.515 81.200 182.605 ;
        RECT 82.125 182.595 82.335 183.385 ;
        RECT 79.980 182.345 81.200 182.515 ;
        RECT 81.660 182.435 82.335 182.595 ;
        RECT 79.640 182.005 80.440 182.175 ;
        RECT 79.760 181.455 80.090 181.835 ;
        RECT 80.270 181.715 80.440 182.005 ;
        RECT 81.030 181.965 81.200 182.345 ;
        RECT 81.370 182.425 82.335 182.435 ;
        RECT 82.525 183.255 82.785 183.645 ;
        RECT 82.995 183.545 83.325 184.005 ;
        RECT 84.200 183.615 85.055 183.785 ;
        RECT 85.260 183.615 85.755 183.785 ;
        RECT 85.925 183.645 86.255 184.005 ;
        RECT 82.525 182.565 82.695 183.255 ;
        RECT 82.865 182.905 83.035 183.085 ;
        RECT 83.205 183.075 83.995 183.325 ;
        RECT 84.200 182.905 84.370 183.615 ;
        RECT 84.540 183.105 84.895 183.325 ;
        RECT 82.865 182.735 84.555 182.905 ;
        RECT 81.370 182.135 81.830 182.425 ;
        RECT 82.525 182.395 84.025 182.565 ;
        RECT 82.525 182.255 82.695 182.395 ;
        RECT 82.135 182.085 82.695 182.255 ;
        RECT 80.610 181.455 80.860 181.915 ;
        RECT 81.030 181.625 81.900 181.965 ;
        RECT 82.135 181.625 82.305 182.085 ;
        RECT 83.140 182.055 84.215 182.225 ;
        RECT 82.475 181.455 82.845 181.915 ;
        RECT 83.140 181.715 83.310 182.055 ;
        RECT 83.480 181.455 83.810 181.885 ;
        RECT 84.045 181.715 84.215 182.055 ;
        RECT 84.385 181.955 84.555 182.735 ;
        RECT 84.725 182.515 84.895 183.105 ;
        RECT 85.065 182.705 85.415 183.325 ;
        RECT 84.725 182.125 85.190 182.515 ;
        RECT 85.585 182.255 85.755 183.615 ;
        RECT 85.925 182.425 86.385 183.475 ;
        RECT 85.360 182.085 85.755 182.255 ;
        RECT 85.360 181.955 85.530 182.085 ;
        RECT 84.385 181.625 85.065 181.955 ;
        RECT 85.280 181.625 85.530 181.955 ;
        RECT 85.700 181.455 85.950 181.915 ;
        RECT 86.120 181.640 86.445 182.425 ;
        RECT 86.615 181.625 86.785 183.745 ;
        RECT 86.955 183.625 87.285 184.005 ;
        RECT 87.455 183.455 87.710 183.745 ;
        RECT 86.960 183.285 87.710 183.455 ;
        RECT 86.960 182.295 87.190 183.285 ;
        RECT 88.805 183.280 89.095 184.005 ;
        RECT 89.265 183.255 90.475 184.005 ;
        RECT 90.735 183.455 90.905 183.835 ;
        RECT 91.085 183.625 91.415 184.005 ;
        RECT 90.735 183.285 91.400 183.455 ;
        RECT 91.595 183.330 91.855 183.835 ;
        RECT 87.360 182.465 87.710 183.115 ;
        RECT 86.960 182.125 87.710 182.295 ;
        RECT 86.955 181.455 87.285 181.955 ;
        RECT 87.455 181.625 87.710 182.125 ;
        RECT 88.805 181.455 89.095 182.620 ;
        RECT 89.265 182.545 89.785 183.085 ;
        RECT 89.955 182.715 90.475 183.255 ;
        RECT 90.665 182.735 90.995 183.105 ;
        RECT 91.230 183.030 91.400 183.285 ;
        RECT 91.230 182.700 91.515 183.030 ;
        RECT 91.230 182.555 91.400 182.700 ;
        RECT 89.265 181.455 90.475 182.545 ;
        RECT 90.735 182.385 91.400 182.555 ;
        RECT 91.685 182.530 91.855 183.330 ;
        RECT 92.065 183.185 92.295 184.005 ;
        RECT 92.465 183.205 92.795 183.835 ;
        RECT 92.045 182.765 92.375 183.015 ;
        RECT 92.545 182.605 92.795 183.205 ;
        RECT 92.965 183.185 93.175 184.005 ;
        RECT 93.410 183.295 93.665 183.825 ;
        RECT 93.835 183.545 94.140 184.005 ;
        RECT 94.385 183.625 95.455 183.795 ;
        RECT 90.735 181.625 90.905 182.385 ;
        RECT 91.085 181.455 91.415 182.215 ;
        RECT 91.585 181.625 91.855 182.530 ;
        RECT 92.065 181.455 92.295 182.595 ;
        RECT 92.465 181.625 92.795 182.605 ;
        RECT 93.410 182.645 93.620 183.295 ;
        RECT 94.385 183.270 94.705 183.625 ;
        RECT 94.380 183.095 94.705 183.270 ;
        RECT 93.790 182.795 94.705 183.095 ;
        RECT 94.875 183.055 95.115 183.455 ;
        RECT 95.285 183.395 95.455 183.625 ;
        RECT 95.625 183.565 95.815 184.005 ;
        RECT 95.985 183.555 96.935 183.835 ;
        RECT 97.155 183.645 97.505 183.815 ;
        RECT 95.285 183.225 95.815 183.395 ;
        RECT 93.790 182.765 94.530 182.795 ;
        RECT 92.965 181.455 93.175 182.595 ;
        RECT 93.410 181.765 93.665 182.645 ;
        RECT 93.835 181.455 94.140 182.595 ;
        RECT 94.360 182.175 94.530 182.765 ;
        RECT 94.875 182.685 95.415 183.055 ;
        RECT 95.595 182.945 95.815 183.225 ;
        RECT 95.985 182.775 96.155 183.555 ;
        RECT 95.750 182.605 96.155 182.775 ;
        RECT 96.325 182.765 96.675 183.385 ;
        RECT 95.750 182.515 95.920 182.605 ;
        RECT 96.845 182.595 97.055 183.385 ;
        RECT 94.700 182.345 95.920 182.515 ;
        RECT 96.380 182.435 97.055 182.595 ;
        RECT 94.360 182.005 95.160 182.175 ;
        RECT 94.480 181.455 94.810 181.835 ;
        RECT 94.990 181.715 95.160 182.005 ;
        RECT 95.750 181.965 95.920 182.345 ;
        RECT 96.090 182.425 97.055 182.435 ;
        RECT 97.245 183.255 97.505 183.645 ;
        RECT 97.715 183.545 98.045 184.005 ;
        RECT 98.920 183.615 99.775 183.785 ;
        RECT 99.980 183.615 100.475 183.785 ;
        RECT 100.645 183.645 100.975 184.005 ;
        RECT 97.245 182.565 97.415 183.255 ;
        RECT 97.585 182.905 97.755 183.085 ;
        RECT 97.925 183.075 98.715 183.325 ;
        RECT 98.920 182.905 99.090 183.615 ;
        RECT 99.260 183.105 99.615 183.325 ;
        RECT 97.585 182.735 99.275 182.905 ;
        RECT 96.090 182.135 96.550 182.425 ;
        RECT 97.245 182.395 98.745 182.565 ;
        RECT 97.245 182.255 97.415 182.395 ;
        RECT 96.855 182.085 97.415 182.255 ;
        RECT 95.330 181.455 95.580 181.915 ;
        RECT 95.750 181.625 96.620 181.965 ;
        RECT 96.855 181.625 97.025 182.085 ;
        RECT 97.860 182.055 98.935 182.225 ;
        RECT 97.195 181.455 97.565 181.915 ;
        RECT 97.860 181.715 98.030 182.055 ;
        RECT 98.200 181.455 98.530 181.885 ;
        RECT 98.765 181.715 98.935 182.055 ;
        RECT 99.105 181.955 99.275 182.735 ;
        RECT 99.445 182.515 99.615 183.105 ;
        RECT 99.785 182.705 100.135 183.325 ;
        RECT 99.445 182.125 99.910 182.515 ;
        RECT 100.305 182.255 100.475 183.615 ;
        RECT 100.645 182.425 101.105 183.475 ;
        RECT 100.080 182.085 100.475 182.255 ;
        RECT 100.080 181.955 100.250 182.085 ;
        RECT 99.105 181.625 99.785 181.955 ;
        RECT 100.000 181.625 100.250 181.955 ;
        RECT 100.420 181.455 100.670 181.915 ;
        RECT 100.840 181.640 101.165 182.425 ;
        RECT 101.335 181.625 101.505 183.745 ;
        RECT 101.675 183.625 102.005 184.005 ;
        RECT 102.175 183.455 102.430 183.745 ;
        RECT 101.680 183.285 102.430 183.455 ;
        RECT 102.605 183.330 102.865 183.835 ;
        RECT 103.045 183.625 103.375 184.005 ;
        RECT 103.555 183.455 103.725 183.835 ;
        RECT 101.680 182.295 101.910 183.285 ;
        RECT 102.080 182.465 102.430 183.115 ;
        RECT 102.605 182.530 102.775 183.330 ;
        RECT 103.060 183.285 103.725 183.455 ;
        RECT 103.060 183.030 103.230 183.285 ;
        RECT 103.985 183.235 107.495 184.005 ;
        RECT 102.945 182.700 103.230 183.030 ;
        RECT 103.465 182.735 103.795 183.105 ;
        RECT 103.060 182.555 103.230 182.700 ;
        RECT 101.680 182.125 102.430 182.295 ;
        RECT 101.675 181.455 102.005 181.955 ;
        RECT 102.175 181.625 102.430 182.125 ;
        RECT 102.605 181.625 102.875 182.530 ;
        RECT 103.060 182.385 103.725 182.555 ;
        RECT 103.045 181.455 103.375 182.215 ;
        RECT 103.555 181.625 103.725 182.385 ;
        RECT 103.985 182.545 105.675 183.065 ;
        RECT 105.845 182.715 107.495 183.235 ;
        RECT 107.705 183.185 107.935 184.005 ;
        RECT 108.105 183.205 108.435 183.835 ;
        RECT 107.685 182.765 108.015 183.015 ;
        RECT 108.185 182.605 108.435 183.205 ;
        RECT 108.605 183.185 108.815 184.005 ;
        RECT 109.320 183.195 109.565 183.800 ;
        RECT 109.785 183.470 110.295 184.005 ;
        RECT 103.985 181.455 107.495 182.545 ;
        RECT 107.705 181.455 107.935 182.595 ;
        RECT 108.105 181.625 108.435 182.605 ;
        RECT 109.045 183.025 110.275 183.195 ;
        RECT 108.605 181.455 108.815 182.595 ;
        RECT 109.045 182.215 109.385 183.025 ;
        RECT 109.555 182.460 110.305 182.650 ;
        RECT 109.045 181.805 109.560 182.215 ;
        RECT 109.795 181.455 109.965 182.215 ;
        RECT 110.135 181.795 110.305 182.460 ;
        RECT 110.475 182.475 110.665 183.835 ;
        RECT 110.835 183.325 111.110 183.835 ;
        RECT 111.300 183.470 111.830 183.835 ;
        RECT 112.255 183.605 112.585 184.005 ;
        RECT 111.655 183.435 111.830 183.470 ;
        RECT 110.835 183.155 111.115 183.325 ;
        RECT 110.835 182.675 111.110 183.155 ;
        RECT 111.315 182.475 111.485 183.275 ;
        RECT 110.475 182.305 111.485 182.475 ;
        RECT 111.655 183.265 112.585 183.435 ;
        RECT 112.755 183.265 113.010 183.835 ;
        RECT 111.655 182.135 111.825 183.265 ;
        RECT 112.415 183.095 112.585 183.265 ;
        RECT 110.700 181.965 111.825 182.135 ;
        RECT 111.995 182.765 112.190 183.095 ;
        RECT 112.415 182.765 112.670 183.095 ;
        RECT 111.995 181.795 112.165 182.765 ;
        RECT 112.840 182.595 113.010 183.265 ;
        RECT 113.185 183.255 114.395 184.005 ;
        RECT 114.565 183.280 114.855 184.005 ;
        RECT 110.135 181.625 112.165 181.795 ;
        RECT 112.335 181.455 112.505 182.595 ;
        RECT 112.675 181.625 113.010 182.595 ;
        RECT 113.185 182.545 113.705 183.085 ;
        RECT 113.875 182.715 114.395 183.255 ;
        RECT 115.300 183.195 115.545 183.800 ;
        RECT 115.765 183.470 116.275 184.005 ;
        RECT 115.025 183.025 116.255 183.195 ;
        RECT 113.185 181.455 114.395 182.545 ;
        RECT 114.565 181.455 114.855 182.620 ;
        RECT 115.025 182.215 115.365 183.025 ;
        RECT 115.535 182.460 116.285 182.650 ;
        RECT 115.025 181.805 115.540 182.215 ;
        RECT 115.775 181.455 115.945 182.215 ;
        RECT 116.115 181.795 116.285 182.460 ;
        RECT 116.455 182.475 116.645 183.835 ;
        RECT 116.815 182.985 117.090 183.835 ;
        RECT 117.280 183.470 117.810 183.835 ;
        RECT 118.235 183.605 118.565 184.005 ;
        RECT 117.635 183.435 117.810 183.470 ;
        RECT 116.815 182.815 117.095 182.985 ;
        RECT 116.815 182.675 117.090 182.815 ;
        RECT 117.295 182.475 117.465 183.275 ;
        RECT 116.455 182.305 117.465 182.475 ;
        RECT 117.635 183.265 118.565 183.435 ;
        RECT 118.735 183.265 118.990 183.835 ;
        RECT 119.715 183.455 119.885 183.835 ;
        RECT 120.065 183.625 120.395 184.005 ;
        RECT 119.715 183.285 120.380 183.455 ;
        RECT 120.575 183.330 120.835 183.835 ;
        RECT 121.010 183.460 126.355 184.005 ;
        RECT 117.635 182.135 117.805 183.265 ;
        RECT 118.395 183.095 118.565 183.265 ;
        RECT 116.680 181.965 117.805 182.135 ;
        RECT 117.975 182.765 118.170 183.095 ;
        RECT 118.395 182.765 118.650 183.095 ;
        RECT 117.975 181.795 118.145 182.765 ;
        RECT 118.820 182.595 118.990 183.265 ;
        RECT 119.645 182.735 119.975 183.105 ;
        RECT 120.210 183.030 120.380 183.285 ;
        RECT 116.115 181.625 118.145 181.795 ;
        RECT 118.315 181.455 118.485 182.595 ;
        RECT 118.655 181.625 118.990 182.595 ;
        RECT 120.210 182.700 120.495 183.030 ;
        RECT 120.210 182.555 120.380 182.700 ;
        RECT 119.715 182.385 120.380 182.555 ;
        RECT 120.665 182.530 120.835 183.330 ;
        RECT 119.715 181.625 119.885 182.385 ;
        RECT 120.065 181.455 120.395 182.215 ;
        RECT 120.565 181.625 120.835 182.530 ;
        RECT 122.600 181.890 122.950 183.140 ;
        RECT 124.430 182.630 124.770 183.460 ;
        RECT 126.525 183.255 127.735 184.005 ;
        RECT 126.525 182.545 127.045 183.085 ;
        RECT 127.215 182.715 127.735 183.255 ;
        RECT 121.010 181.455 126.355 181.890 ;
        RECT 126.525 181.455 127.735 182.545 ;
        RECT 14.660 181.285 127.820 181.455 ;
        RECT 14.745 180.195 15.955 181.285 ;
        RECT 14.745 179.485 15.265 180.025 ;
        RECT 15.435 179.655 15.955 180.195 ;
        RECT 16.125 180.195 17.335 181.285 ;
        RECT 17.510 180.850 22.855 181.285 ;
        RECT 16.125 179.655 16.645 180.195 ;
        RECT 16.815 179.485 17.335 180.025 ;
        RECT 19.100 179.600 19.450 180.850 ;
        RECT 23.065 180.145 23.295 181.285 ;
        RECT 23.465 180.135 23.795 181.115 ;
        RECT 23.965 180.145 24.175 181.285 ;
        RECT 14.745 178.735 15.955 179.485 ;
        RECT 16.125 178.735 17.335 179.485 ;
        RECT 20.930 179.280 21.270 180.110 ;
        RECT 23.045 179.725 23.375 179.975 ;
        RECT 17.510 178.735 22.855 179.280 ;
        RECT 23.065 178.735 23.295 179.555 ;
        RECT 23.545 179.535 23.795 180.135 ;
        RECT 24.405 180.120 24.695 181.285 ;
        RECT 24.870 180.615 25.125 181.115 ;
        RECT 25.295 180.785 25.625 181.285 ;
        RECT 24.870 180.445 25.620 180.615 ;
        RECT 24.870 179.625 25.220 180.275 ;
        RECT 23.465 178.905 23.795 179.535 ;
        RECT 23.965 178.735 24.175 179.555 ;
        RECT 24.405 178.735 24.695 179.460 ;
        RECT 25.390 179.455 25.620 180.445 ;
        RECT 24.870 179.285 25.620 179.455 ;
        RECT 24.870 178.995 25.125 179.285 ;
        RECT 25.295 178.735 25.625 179.115 ;
        RECT 25.795 178.995 25.965 181.115 ;
        RECT 26.135 180.315 26.460 181.100 ;
        RECT 26.630 180.825 26.880 181.285 ;
        RECT 27.050 180.785 27.300 181.115 ;
        RECT 27.515 180.785 28.195 181.115 ;
        RECT 27.050 180.655 27.220 180.785 ;
        RECT 26.825 180.485 27.220 180.655 ;
        RECT 26.195 179.265 26.655 180.315 ;
        RECT 26.825 179.125 26.995 180.485 ;
        RECT 27.390 180.225 27.855 180.615 ;
        RECT 27.165 179.415 27.515 180.035 ;
        RECT 27.685 179.635 27.855 180.225 ;
        RECT 28.025 180.005 28.195 180.785 ;
        RECT 28.365 180.685 28.535 181.025 ;
        RECT 28.770 180.855 29.100 181.285 ;
        RECT 29.270 180.685 29.440 181.025 ;
        RECT 29.735 180.825 30.105 181.285 ;
        RECT 28.365 180.515 29.440 180.685 ;
        RECT 30.275 180.655 30.445 181.115 ;
        RECT 30.680 180.775 31.550 181.115 ;
        RECT 31.720 180.825 31.970 181.285 ;
        RECT 29.885 180.485 30.445 180.655 ;
        RECT 29.885 180.345 30.055 180.485 ;
        RECT 28.555 180.175 30.055 180.345 ;
        RECT 30.750 180.315 31.210 180.605 ;
        RECT 28.025 179.835 29.715 180.005 ;
        RECT 27.685 179.415 28.040 179.635 ;
        RECT 28.210 179.125 28.380 179.835 ;
        RECT 28.585 179.415 29.375 179.665 ;
        RECT 29.545 179.655 29.715 179.835 ;
        RECT 29.885 179.485 30.055 180.175 ;
        RECT 26.325 178.735 26.655 179.095 ;
        RECT 26.825 178.955 27.320 179.125 ;
        RECT 27.525 178.955 28.380 179.125 ;
        RECT 29.255 178.735 29.585 179.195 ;
        RECT 29.795 179.095 30.055 179.485 ;
        RECT 30.245 180.305 31.210 180.315 ;
        RECT 31.380 180.395 31.550 180.775 ;
        RECT 32.140 180.735 32.310 181.025 ;
        RECT 32.490 180.905 32.820 181.285 ;
        RECT 32.140 180.565 32.940 180.735 ;
        RECT 30.245 180.145 30.920 180.305 ;
        RECT 31.380 180.225 32.600 180.395 ;
        RECT 30.245 179.355 30.455 180.145 ;
        RECT 31.380 180.135 31.550 180.225 ;
        RECT 30.625 179.355 30.975 179.975 ;
        RECT 31.145 179.965 31.550 180.135 ;
        RECT 31.145 179.185 31.315 179.965 ;
        RECT 31.485 179.515 31.705 179.795 ;
        RECT 31.885 179.685 32.425 180.055 ;
        RECT 32.770 179.975 32.940 180.565 ;
        RECT 33.160 180.145 33.465 181.285 ;
        RECT 33.635 180.095 33.890 180.975 ;
        RECT 32.770 179.945 33.510 179.975 ;
        RECT 31.485 179.345 32.015 179.515 ;
        RECT 29.795 178.925 30.145 179.095 ;
        RECT 30.365 178.905 31.315 179.185 ;
        RECT 31.485 178.735 31.675 179.175 ;
        RECT 31.845 179.115 32.015 179.345 ;
        RECT 32.185 179.285 32.425 179.685 ;
        RECT 32.595 179.645 33.510 179.945 ;
        RECT 32.595 179.470 32.920 179.645 ;
        RECT 32.595 179.115 32.915 179.470 ;
        RECT 33.680 179.445 33.890 180.095 ;
        RECT 34.065 180.195 35.735 181.285 ;
        RECT 34.065 179.675 34.815 180.195 ;
        RECT 35.945 180.145 36.175 181.285 ;
        RECT 36.345 180.135 36.675 181.115 ;
        RECT 36.845 180.145 37.055 181.285 ;
        RECT 37.285 180.210 37.555 181.115 ;
        RECT 37.725 180.525 38.055 181.285 ;
        RECT 38.235 180.355 38.405 181.115 ;
        RECT 34.985 179.505 35.735 180.025 ;
        RECT 35.925 179.725 36.255 179.975 ;
        RECT 31.845 178.945 32.915 179.115 ;
        RECT 33.160 178.735 33.465 179.195 ;
        RECT 33.635 178.915 33.890 179.445 ;
        RECT 34.065 178.735 35.735 179.505 ;
        RECT 35.945 178.735 36.175 179.555 ;
        RECT 36.425 179.535 36.675 180.135 ;
        RECT 36.345 178.905 36.675 179.535 ;
        RECT 36.845 178.735 37.055 179.555 ;
        RECT 37.285 179.410 37.455 180.210 ;
        RECT 37.740 180.185 38.405 180.355 ;
        RECT 39.585 180.195 43.095 181.285 ;
        RECT 43.355 180.355 43.525 181.115 ;
        RECT 43.705 180.525 44.035 181.285 ;
        RECT 37.740 180.040 37.910 180.185 ;
        RECT 37.625 179.710 37.910 180.040 ;
        RECT 37.740 179.455 37.910 179.710 ;
        RECT 38.145 179.635 38.475 180.005 ;
        RECT 39.585 179.675 41.275 180.195 ;
        RECT 43.355 180.185 44.020 180.355 ;
        RECT 44.205 180.210 44.475 181.115 ;
        RECT 43.850 180.040 44.020 180.185 ;
        RECT 41.445 179.505 43.095 180.025 ;
        RECT 43.285 179.635 43.615 180.005 ;
        RECT 43.850 179.710 44.135 180.040 ;
        RECT 37.285 178.905 37.545 179.410 ;
        RECT 37.740 179.285 38.405 179.455 ;
        RECT 37.725 178.735 38.055 179.115 ;
        RECT 38.235 178.905 38.405 179.285 ;
        RECT 39.585 178.735 43.095 179.505 ;
        RECT 43.850 179.455 44.020 179.710 ;
        RECT 43.355 179.285 44.020 179.455 ;
        RECT 44.305 179.410 44.475 180.210 ;
        RECT 45.105 180.195 48.615 181.285 ;
        RECT 45.105 179.675 46.795 180.195 ;
        RECT 48.845 180.145 49.055 181.285 ;
        RECT 49.225 180.135 49.555 181.115 ;
        RECT 49.725 180.145 49.955 181.285 ;
        RECT 46.965 179.505 48.615 180.025 ;
        RECT 43.355 178.905 43.525 179.285 ;
        RECT 43.705 178.735 44.035 179.115 ;
        RECT 44.215 178.905 44.475 179.410 ;
        RECT 45.105 178.735 48.615 179.505 ;
        RECT 48.845 178.735 49.055 179.555 ;
        RECT 49.225 179.535 49.475 180.135 ;
        RECT 50.165 180.120 50.455 181.285 ;
        RECT 50.625 180.195 52.295 181.285 ;
        RECT 49.645 179.725 49.975 179.975 ;
        RECT 50.625 179.675 51.375 180.195 ;
        RECT 52.505 180.145 52.735 181.285 ;
        RECT 52.905 180.135 53.235 181.115 ;
        RECT 53.405 180.145 53.615 181.285 ;
        RECT 53.845 180.525 54.360 180.935 ;
        RECT 54.595 180.525 54.765 181.285 ;
        RECT 54.935 180.945 56.965 181.115 ;
        RECT 49.225 178.905 49.555 179.535 ;
        RECT 49.725 178.735 49.955 179.555 ;
        RECT 51.545 179.505 52.295 180.025 ;
        RECT 52.485 179.725 52.815 179.975 ;
        RECT 50.165 178.735 50.455 179.460 ;
        RECT 50.625 178.735 52.295 179.505 ;
        RECT 52.505 178.735 52.735 179.555 ;
        RECT 52.985 179.535 53.235 180.135 ;
        RECT 53.845 179.715 54.185 180.525 ;
        RECT 54.935 180.280 55.105 180.945 ;
        RECT 55.500 180.605 56.625 180.775 ;
        RECT 54.355 180.090 55.105 180.280 ;
        RECT 55.275 180.265 56.285 180.435 ;
        RECT 52.905 178.905 53.235 179.535 ;
        RECT 53.405 178.735 53.615 179.555 ;
        RECT 53.845 179.545 55.075 179.715 ;
        RECT 54.120 178.940 54.365 179.545 ;
        RECT 54.585 178.735 55.095 179.270 ;
        RECT 55.275 178.905 55.465 180.265 ;
        RECT 55.635 179.585 55.910 180.065 ;
        RECT 55.635 179.415 55.915 179.585 ;
        RECT 56.115 179.465 56.285 180.265 ;
        RECT 56.455 179.475 56.625 180.605 ;
        RECT 56.795 179.975 56.965 180.945 ;
        RECT 57.135 180.145 57.305 181.285 ;
        RECT 57.475 180.145 57.810 181.115 ;
        RECT 58.075 180.355 58.245 181.115 ;
        RECT 58.425 180.525 58.755 181.285 ;
        RECT 58.075 180.185 58.740 180.355 ;
        RECT 58.925 180.210 59.195 181.115 ;
        RECT 59.370 180.850 64.715 181.285 ;
        RECT 64.890 180.850 70.235 181.285 ;
        RECT 70.410 180.850 75.755 181.285 ;
        RECT 56.795 179.645 56.990 179.975 ;
        RECT 57.215 179.645 57.470 179.975 ;
        RECT 57.215 179.475 57.385 179.645 ;
        RECT 57.640 179.475 57.810 180.145 ;
        RECT 58.570 180.040 58.740 180.185 ;
        RECT 58.005 179.635 58.335 180.005 ;
        RECT 58.570 179.710 58.855 180.040 ;
        RECT 55.635 178.905 55.910 179.415 ;
        RECT 56.455 179.305 57.385 179.475 ;
        RECT 56.455 179.270 56.630 179.305 ;
        RECT 56.100 178.905 56.630 179.270 ;
        RECT 57.055 178.735 57.385 179.135 ;
        RECT 57.555 178.905 57.810 179.475 ;
        RECT 58.570 179.455 58.740 179.710 ;
        RECT 58.075 179.285 58.740 179.455 ;
        RECT 59.025 179.410 59.195 180.210 ;
        RECT 60.960 179.600 61.310 180.850 ;
        RECT 58.075 178.905 58.245 179.285 ;
        RECT 58.425 178.735 58.755 179.115 ;
        RECT 58.935 178.905 59.195 179.410 ;
        RECT 62.790 179.280 63.130 180.110 ;
        RECT 66.480 179.600 66.830 180.850 ;
        RECT 68.310 179.280 68.650 180.110 ;
        RECT 72.000 179.600 72.350 180.850 ;
        RECT 75.925 180.120 76.215 181.285 ;
        RECT 77.315 180.305 77.645 181.115 ;
        RECT 77.815 180.485 78.055 181.285 ;
        RECT 77.315 180.135 78.030 180.305 ;
        RECT 73.830 179.280 74.170 180.110 ;
        RECT 77.310 179.725 77.690 179.965 ;
        RECT 77.860 179.895 78.030 180.135 ;
        RECT 78.235 180.265 78.405 181.115 ;
        RECT 78.575 180.485 78.905 181.285 ;
        RECT 79.075 180.265 79.245 181.115 ;
        RECT 78.235 180.095 79.245 180.265 ;
        RECT 79.415 180.135 79.745 181.285 ;
        RECT 80.065 180.525 80.580 180.935 ;
        RECT 80.815 180.525 80.985 181.285 ;
        RECT 81.155 180.945 83.185 181.115 ;
        RECT 78.750 179.925 79.245 180.095 ;
        RECT 77.860 179.725 78.360 179.895 ;
        RECT 78.745 179.755 79.245 179.925 ;
        RECT 77.860 179.555 78.030 179.725 ;
        RECT 78.750 179.555 79.245 179.755 ;
        RECT 59.370 178.735 64.715 179.280 ;
        RECT 64.890 178.735 70.235 179.280 ;
        RECT 70.410 178.735 75.755 179.280 ;
        RECT 75.925 178.735 76.215 179.460 ;
        RECT 77.395 179.385 78.030 179.555 ;
        RECT 78.235 179.385 79.245 179.555 ;
        RECT 80.065 179.715 80.405 180.525 ;
        RECT 81.155 180.280 81.325 180.945 ;
        RECT 81.720 180.605 82.845 180.775 ;
        RECT 80.575 180.090 81.325 180.280 ;
        RECT 81.495 180.265 82.505 180.435 ;
        RECT 80.065 179.545 81.295 179.715 ;
        RECT 77.395 178.905 77.565 179.385 ;
        RECT 77.745 178.735 77.985 179.215 ;
        RECT 78.235 178.905 78.405 179.385 ;
        RECT 78.575 178.735 78.905 179.215 ;
        RECT 79.075 178.905 79.245 179.385 ;
        RECT 79.415 178.735 79.745 179.535 ;
        RECT 80.340 178.940 80.585 179.545 ;
        RECT 80.805 178.735 81.315 179.270 ;
        RECT 81.495 178.905 81.685 180.265 ;
        RECT 81.855 179.585 82.130 180.065 ;
        RECT 81.855 179.415 82.135 179.585 ;
        RECT 82.335 179.465 82.505 180.265 ;
        RECT 82.675 179.475 82.845 180.605 ;
        RECT 83.015 179.975 83.185 180.945 ;
        RECT 83.355 180.145 83.525 181.285 ;
        RECT 83.695 180.145 84.030 181.115 ;
        RECT 83.015 179.645 83.210 179.975 ;
        RECT 83.435 179.645 83.690 179.975 ;
        RECT 83.435 179.475 83.605 179.645 ;
        RECT 83.860 179.475 84.030 180.145 ;
        RECT 81.855 178.905 82.130 179.415 ;
        RECT 82.675 179.305 83.605 179.475 ;
        RECT 82.675 179.270 82.850 179.305 ;
        RECT 82.320 178.905 82.850 179.270 ;
        RECT 83.275 178.735 83.605 179.135 ;
        RECT 83.775 178.905 84.030 179.475 ;
        RECT 84.210 180.095 84.465 180.975 ;
        RECT 84.635 180.145 84.940 181.285 ;
        RECT 85.280 180.905 85.610 181.285 ;
        RECT 85.790 180.735 85.960 181.025 ;
        RECT 86.130 180.825 86.380 181.285 ;
        RECT 85.160 180.565 85.960 180.735 ;
        RECT 86.550 180.775 87.420 181.115 ;
        RECT 84.210 179.445 84.420 180.095 ;
        RECT 85.160 179.975 85.330 180.565 ;
        RECT 86.550 180.395 86.720 180.775 ;
        RECT 87.655 180.655 87.825 181.115 ;
        RECT 87.995 180.825 88.365 181.285 ;
        RECT 88.660 180.685 88.830 181.025 ;
        RECT 89.000 180.855 89.330 181.285 ;
        RECT 89.565 180.685 89.735 181.025 ;
        RECT 85.500 180.225 86.720 180.395 ;
        RECT 86.890 180.315 87.350 180.605 ;
        RECT 87.655 180.485 88.215 180.655 ;
        RECT 88.660 180.515 89.735 180.685 ;
        RECT 89.905 180.785 90.585 181.115 ;
        RECT 90.800 180.785 91.050 181.115 ;
        RECT 91.220 180.825 91.470 181.285 ;
        RECT 88.045 180.345 88.215 180.485 ;
        RECT 86.890 180.305 87.855 180.315 ;
        RECT 86.550 180.135 86.720 180.225 ;
        RECT 87.180 180.145 87.855 180.305 ;
        RECT 84.590 179.945 85.330 179.975 ;
        RECT 84.590 179.645 85.505 179.945 ;
        RECT 85.180 179.470 85.505 179.645 ;
        RECT 84.210 178.915 84.465 179.445 ;
        RECT 84.635 178.735 84.940 179.195 ;
        RECT 85.185 179.115 85.505 179.470 ;
        RECT 85.675 179.685 86.215 180.055 ;
        RECT 86.550 179.965 86.955 180.135 ;
        RECT 85.675 179.285 85.915 179.685 ;
        RECT 86.395 179.515 86.615 179.795 ;
        RECT 86.085 179.345 86.615 179.515 ;
        RECT 86.085 179.115 86.255 179.345 ;
        RECT 86.785 179.185 86.955 179.965 ;
        RECT 87.125 179.355 87.475 179.975 ;
        RECT 87.645 179.355 87.855 180.145 ;
        RECT 88.045 180.175 89.545 180.345 ;
        RECT 88.045 179.485 88.215 180.175 ;
        RECT 89.905 180.005 90.075 180.785 ;
        RECT 90.880 180.655 91.050 180.785 ;
        RECT 88.385 179.835 90.075 180.005 ;
        RECT 90.245 180.225 90.710 180.615 ;
        RECT 90.880 180.485 91.275 180.655 ;
        RECT 88.385 179.655 88.555 179.835 ;
        RECT 85.185 178.945 86.255 179.115 ;
        RECT 86.425 178.735 86.615 179.175 ;
        RECT 86.785 178.905 87.735 179.185 ;
        RECT 88.045 179.095 88.305 179.485 ;
        RECT 88.725 179.415 89.515 179.665 ;
        RECT 87.955 178.925 88.305 179.095 ;
        RECT 88.515 178.735 88.845 179.195 ;
        RECT 89.720 179.125 89.890 179.835 ;
        RECT 90.245 179.635 90.415 180.225 ;
        RECT 90.060 179.415 90.415 179.635 ;
        RECT 90.585 179.415 90.935 180.035 ;
        RECT 91.105 179.125 91.275 180.485 ;
        RECT 91.640 180.315 91.965 181.100 ;
        RECT 91.445 179.265 91.905 180.315 ;
        RECT 89.720 178.955 90.575 179.125 ;
        RECT 90.780 178.955 91.275 179.125 ;
        RECT 91.445 178.735 91.775 179.095 ;
        RECT 92.135 178.995 92.305 181.115 ;
        RECT 92.475 180.785 92.805 181.285 ;
        RECT 92.975 180.615 93.230 181.115 ;
        RECT 92.480 180.445 93.230 180.615 ;
        RECT 92.480 179.455 92.710 180.445 ;
        RECT 92.880 179.625 93.230 180.275 ;
        RECT 93.405 180.195 95.995 181.285 ;
        RECT 96.170 180.850 101.515 181.285 ;
        RECT 93.405 179.675 94.615 180.195 ;
        RECT 94.785 179.505 95.995 180.025 ;
        RECT 97.760 179.600 98.110 180.850 ;
        RECT 101.685 180.120 101.975 181.285 ;
        RECT 103.070 180.850 108.415 181.285 ;
        RECT 92.480 179.285 93.230 179.455 ;
        RECT 92.475 178.735 92.805 179.115 ;
        RECT 92.975 178.995 93.230 179.285 ;
        RECT 93.405 178.735 95.995 179.505 ;
        RECT 99.590 179.280 99.930 180.110 ;
        RECT 104.660 179.600 105.010 180.850 ;
        RECT 96.170 178.735 101.515 179.280 ;
        RECT 101.685 178.735 101.975 179.460 ;
        RECT 106.490 179.280 106.830 180.110 ;
        RECT 108.590 180.095 108.845 180.975 ;
        RECT 109.015 180.145 109.320 181.285 ;
        RECT 109.660 180.905 109.990 181.285 ;
        RECT 110.170 180.735 110.340 181.025 ;
        RECT 110.510 180.825 110.760 181.285 ;
        RECT 109.540 180.565 110.340 180.735 ;
        RECT 110.930 180.775 111.800 181.115 ;
        RECT 108.590 179.445 108.800 180.095 ;
        RECT 109.540 179.975 109.710 180.565 ;
        RECT 110.930 180.395 111.100 180.775 ;
        RECT 112.035 180.655 112.205 181.115 ;
        RECT 112.375 180.825 112.745 181.285 ;
        RECT 113.040 180.685 113.210 181.025 ;
        RECT 113.380 180.855 113.710 181.285 ;
        RECT 113.945 180.685 114.115 181.025 ;
        RECT 109.880 180.225 111.100 180.395 ;
        RECT 111.270 180.315 111.730 180.605 ;
        RECT 112.035 180.485 112.595 180.655 ;
        RECT 113.040 180.515 114.115 180.685 ;
        RECT 114.285 180.785 114.965 181.115 ;
        RECT 115.180 180.785 115.430 181.115 ;
        RECT 115.600 180.825 115.850 181.285 ;
        RECT 112.425 180.345 112.595 180.485 ;
        RECT 111.270 180.305 112.235 180.315 ;
        RECT 110.930 180.135 111.100 180.225 ;
        RECT 111.560 180.145 112.235 180.305 ;
        RECT 108.970 179.945 109.710 179.975 ;
        RECT 108.970 179.645 109.885 179.945 ;
        RECT 109.560 179.470 109.885 179.645 ;
        RECT 103.070 178.735 108.415 179.280 ;
        RECT 108.590 178.915 108.845 179.445 ;
        RECT 109.015 178.735 109.320 179.195 ;
        RECT 109.565 179.115 109.885 179.470 ;
        RECT 110.055 179.685 110.595 180.055 ;
        RECT 110.930 179.965 111.335 180.135 ;
        RECT 110.055 179.285 110.295 179.685 ;
        RECT 110.775 179.515 110.995 179.795 ;
        RECT 110.465 179.345 110.995 179.515 ;
        RECT 110.465 179.115 110.635 179.345 ;
        RECT 111.165 179.185 111.335 179.965 ;
        RECT 111.505 179.355 111.855 179.975 ;
        RECT 112.025 179.355 112.235 180.145 ;
        RECT 112.425 180.175 113.925 180.345 ;
        RECT 112.425 179.485 112.595 180.175 ;
        RECT 114.285 180.005 114.455 180.785 ;
        RECT 115.260 180.655 115.430 180.785 ;
        RECT 112.765 179.835 114.455 180.005 ;
        RECT 114.625 180.225 115.090 180.615 ;
        RECT 115.260 180.485 115.655 180.655 ;
        RECT 112.765 179.655 112.935 179.835 ;
        RECT 109.565 178.945 110.635 179.115 ;
        RECT 110.805 178.735 110.995 179.175 ;
        RECT 111.165 178.905 112.115 179.185 ;
        RECT 112.425 179.095 112.685 179.485 ;
        RECT 113.105 179.415 113.895 179.665 ;
        RECT 112.335 178.925 112.685 179.095 ;
        RECT 112.895 178.735 113.225 179.195 ;
        RECT 114.100 179.125 114.270 179.835 ;
        RECT 114.625 179.635 114.795 180.225 ;
        RECT 114.440 179.415 114.795 179.635 ;
        RECT 114.965 179.415 115.315 180.035 ;
        RECT 115.485 179.125 115.655 180.485 ;
        RECT 116.020 180.315 116.345 181.100 ;
        RECT 115.825 179.265 116.285 180.315 ;
        RECT 114.100 178.955 114.955 179.125 ;
        RECT 115.160 178.955 115.655 179.125 ;
        RECT 115.825 178.735 116.155 179.095 ;
        RECT 116.515 178.995 116.685 181.115 ;
        RECT 116.855 180.785 117.185 181.285 ;
        RECT 117.355 180.615 117.610 181.115 ;
        RECT 116.860 180.445 117.610 180.615 ;
        RECT 117.785 180.525 118.300 180.935 ;
        RECT 118.535 180.525 118.705 181.285 ;
        RECT 118.875 180.945 120.905 181.115 ;
        RECT 116.860 179.455 117.090 180.445 ;
        RECT 117.260 179.625 117.610 180.275 ;
        RECT 117.785 179.715 118.125 180.525 ;
        RECT 118.875 180.280 119.045 180.945 ;
        RECT 119.440 180.605 120.565 180.775 ;
        RECT 118.295 180.090 119.045 180.280 ;
        RECT 119.215 180.265 120.225 180.435 ;
        RECT 117.785 179.545 119.015 179.715 ;
        RECT 116.860 179.285 117.610 179.455 ;
        RECT 116.855 178.735 117.185 179.115 ;
        RECT 117.355 178.995 117.610 179.285 ;
        RECT 118.060 178.940 118.305 179.545 ;
        RECT 118.525 178.735 119.035 179.270 ;
        RECT 119.215 178.905 119.405 180.265 ;
        RECT 119.575 179.925 119.850 180.065 ;
        RECT 119.575 179.755 119.855 179.925 ;
        RECT 119.575 178.905 119.850 179.755 ;
        RECT 120.055 179.465 120.225 180.265 ;
        RECT 120.395 179.475 120.565 180.605 ;
        RECT 120.735 179.975 120.905 180.945 ;
        RECT 121.075 180.145 121.245 181.285 ;
        RECT 121.415 180.145 121.750 181.115 ;
        RECT 120.735 179.645 120.930 179.975 ;
        RECT 121.155 179.645 121.410 179.975 ;
        RECT 121.155 179.475 121.325 179.645 ;
        RECT 121.580 179.475 121.750 180.145 ;
        RECT 122.845 180.195 126.355 181.285 ;
        RECT 126.525 180.195 127.735 181.285 ;
        RECT 122.845 179.675 124.535 180.195 ;
        RECT 124.705 179.505 126.355 180.025 ;
        RECT 126.525 179.655 127.045 180.195 ;
        RECT 120.395 179.305 121.325 179.475 ;
        RECT 120.395 179.270 120.570 179.305 ;
        RECT 120.040 178.905 120.570 179.270 ;
        RECT 120.995 178.735 121.325 179.135 ;
        RECT 121.495 178.905 121.750 179.475 ;
        RECT 122.845 178.735 126.355 179.505 ;
        RECT 127.215 179.485 127.735 180.025 ;
        RECT 126.525 178.735 127.735 179.485 ;
        RECT 14.660 178.565 127.820 178.735 ;
        RECT 14.745 177.815 15.955 178.565 ;
        RECT 17.050 178.020 22.395 178.565 ;
        RECT 22.570 178.020 27.915 178.565 ;
        RECT 14.745 177.275 15.265 177.815 ;
        RECT 15.435 177.105 15.955 177.645 ;
        RECT 14.745 176.015 15.955 177.105 ;
        RECT 18.640 176.450 18.990 177.700 ;
        RECT 20.470 177.190 20.810 178.020 ;
        RECT 24.160 176.450 24.510 177.700 ;
        RECT 25.990 177.190 26.330 178.020 ;
        RECT 28.085 177.890 28.345 178.395 ;
        RECT 28.525 178.185 28.855 178.565 ;
        RECT 29.035 178.015 29.205 178.395 ;
        RECT 28.085 177.090 28.255 177.890 ;
        RECT 28.540 177.845 29.205 178.015 ;
        RECT 28.540 177.590 28.710 177.845 ;
        RECT 29.470 177.825 29.725 178.395 ;
        RECT 29.895 178.165 30.225 178.565 ;
        RECT 30.650 178.030 31.180 178.395 ;
        RECT 30.650 177.995 30.825 178.030 ;
        RECT 29.895 177.825 30.825 177.995 ;
        RECT 28.425 177.260 28.710 177.590 ;
        RECT 28.945 177.295 29.275 177.665 ;
        RECT 28.540 177.115 28.710 177.260 ;
        RECT 29.470 177.155 29.640 177.825 ;
        RECT 29.895 177.655 30.065 177.825 ;
        RECT 29.810 177.325 30.065 177.655 ;
        RECT 30.290 177.325 30.485 177.655 ;
        RECT 17.050 176.015 22.395 176.450 ;
        RECT 22.570 176.015 27.915 176.450 ;
        RECT 28.085 176.185 28.355 177.090 ;
        RECT 28.540 176.945 29.205 177.115 ;
        RECT 28.525 176.015 28.855 176.775 ;
        RECT 29.035 176.185 29.205 176.945 ;
        RECT 29.470 176.185 29.805 177.155 ;
        RECT 29.975 176.015 30.145 177.155 ;
        RECT 30.315 176.355 30.485 177.325 ;
        RECT 30.655 176.695 30.825 177.825 ;
        RECT 30.995 177.035 31.165 177.835 ;
        RECT 31.370 177.545 31.645 178.395 ;
        RECT 31.365 177.375 31.645 177.545 ;
        RECT 31.370 177.235 31.645 177.375 ;
        RECT 31.815 177.035 32.005 178.395 ;
        RECT 32.185 178.030 32.695 178.565 ;
        RECT 32.915 177.755 33.160 178.360 ;
        RECT 33.605 177.795 37.115 178.565 ;
        RECT 37.285 177.840 37.575 178.565 ;
        RECT 37.750 178.020 43.095 178.565 ;
        RECT 32.205 177.585 33.435 177.755 ;
        RECT 30.995 176.865 32.005 177.035 ;
        RECT 32.175 177.020 32.925 177.210 ;
        RECT 30.655 176.525 31.780 176.695 ;
        RECT 32.175 176.355 32.345 177.020 ;
        RECT 33.095 176.775 33.435 177.585 ;
        RECT 30.315 176.185 32.345 176.355 ;
        RECT 32.515 176.015 32.685 176.775 ;
        RECT 32.920 176.365 33.435 176.775 ;
        RECT 33.605 177.105 35.295 177.625 ;
        RECT 35.465 177.275 37.115 177.795 ;
        RECT 33.605 176.015 37.115 177.105 ;
        RECT 37.285 176.015 37.575 177.180 ;
        RECT 39.340 176.450 39.690 177.700 ;
        RECT 41.170 177.190 41.510 178.020 ;
        RECT 43.640 177.855 43.895 178.385 ;
        RECT 44.075 178.105 44.360 178.565 ;
        RECT 43.640 176.995 43.820 177.855 ;
        RECT 44.540 177.655 44.790 178.305 ;
        RECT 43.990 177.325 44.790 177.655 ;
        RECT 43.640 176.525 43.895 176.995 ;
        RECT 37.750 176.015 43.095 176.450 ;
        RECT 43.555 176.355 43.895 176.525 ;
        RECT 43.640 176.325 43.895 176.355 ;
        RECT 44.075 176.015 44.360 176.815 ;
        RECT 44.540 176.735 44.790 177.325 ;
        RECT 44.990 177.970 45.310 178.300 ;
        RECT 45.490 178.085 46.150 178.565 ;
        RECT 46.350 178.175 47.200 178.345 ;
        RECT 44.990 177.075 45.180 177.970 ;
        RECT 45.500 177.645 46.160 177.915 ;
        RECT 45.830 177.585 46.160 177.645 ;
        RECT 45.350 177.415 45.680 177.475 ;
        RECT 46.350 177.415 46.520 178.175 ;
        RECT 47.760 178.105 48.080 178.565 ;
        RECT 48.280 177.925 48.530 178.355 ;
        RECT 48.820 178.125 49.230 178.565 ;
        RECT 49.400 178.185 50.415 178.385 ;
        RECT 46.690 177.755 47.940 177.925 ;
        RECT 46.690 177.635 47.020 177.755 ;
        RECT 45.350 177.245 47.250 177.415 ;
        RECT 44.990 176.905 46.910 177.075 ;
        RECT 44.990 176.885 45.310 176.905 ;
        RECT 44.540 176.225 44.870 176.735 ;
        RECT 45.140 176.275 45.310 176.885 ;
        RECT 47.080 176.735 47.250 177.245 ;
        RECT 47.420 177.175 47.600 177.585 ;
        RECT 47.770 176.995 47.940 177.755 ;
        RECT 45.480 176.015 45.810 176.705 ;
        RECT 46.040 176.565 47.250 176.735 ;
        RECT 47.420 176.685 47.940 176.995 ;
        RECT 48.110 177.585 48.530 177.925 ;
        RECT 48.820 177.585 49.230 177.915 ;
        RECT 48.110 176.815 48.300 177.585 ;
        RECT 49.400 177.455 49.570 178.185 ;
        RECT 50.715 178.015 50.885 178.345 ;
        RECT 51.055 178.185 51.385 178.565 ;
        RECT 49.740 177.635 50.090 178.005 ;
        RECT 49.400 177.415 49.820 177.455 ;
        RECT 48.470 177.245 49.820 177.415 ;
        RECT 48.470 177.085 48.720 177.245 ;
        RECT 49.230 176.815 49.480 177.075 ;
        RECT 48.110 176.565 49.480 176.815 ;
        RECT 46.040 176.275 46.280 176.565 ;
        RECT 47.080 176.485 47.250 176.565 ;
        RECT 46.480 176.015 46.900 176.395 ;
        RECT 47.080 176.235 47.710 176.485 ;
        RECT 48.180 176.015 48.510 176.395 ;
        RECT 48.680 176.275 48.850 176.565 ;
        RECT 49.650 176.400 49.820 177.245 ;
        RECT 50.270 177.075 50.490 177.945 ;
        RECT 50.715 177.825 51.410 178.015 ;
        RECT 49.990 176.695 50.490 177.075 ;
        RECT 50.660 177.025 51.070 177.645 ;
        RECT 51.240 176.855 51.410 177.825 ;
        RECT 50.715 176.685 51.410 176.855 ;
        RECT 49.030 176.015 49.410 176.395 ;
        RECT 49.650 176.230 50.480 176.400 ;
        RECT 50.715 176.185 50.885 176.685 ;
        RECT 51.055 176.015 51.385 176.515 ;
        RECT 51.600 176.185 51.825 178.305 ;
        RECT 51.995 178.185 52.325 178.565 ;
        RECT 52.495 178.015 52.665 178.305 ;
        RECT 52.000 177.845 52.665 178.015 ;
        RECT 53.300 177.855 53.555 178.385 ;
        RECT 53.735 178.105 54.020 178.565 ;
        RECT 52.000 176.855 52.230 177.845 ;
        RECT 52.400 177.025 52.750 177.675 ;
        RECT 53.300 176.995 53.480 177.855 ;
        RECT 54.200 177.655 54.450 178.305 ;
        RECT 53.650 177.325 54.450 177.655 ;
        RECT 52.000 176.685 52.665 176.855 ;
        RECT 51.995 176.015 52.325 176.515 ;
        RECT 52.495 176.185 52.665 176.685 ;
        RECT 53.300 176.525 53.555 176.995 ;
        RECT 53.215 176.355 53.555 176.525 ;
        RECT 53.300 176.325 53.555 176.355 ;
        RECT 53.735 176.015 54.020 176.815 ;
        RECT 54.200 176.735 54.450 177.325 ;
        RECT 54.650 177.970 54.970 178.300 ;
        RECT 55.150 178.085 55.810 178.565 ;
        RECT 56.010 178.175 56.860 178.345 ;
        RECT 54.650 177.075 54.840 177.970 ;
        RECT 55.160 177.645 55.820 177.915 ;
        RECT 55.490 177.585 55.820 177.645 ;
        RECT 55.010 177.415 55.340 177.475 ;
        RECT 56.010 177.415 56.180 178.175 ;
        RECT 57.420 178.105 57.740 178.565 ;
        RECT 57.940 177.925 58.190 178.355 ;
        RECT 58.480 178.125 58.890 178.565 ;
        RECT 59.060 178.185 60.075 178.385 ;
        RECT 56.350 177.755 57.600 177.925 ;
        RECT 56.350 177.635 56.680 177.755 ;
        RECT 55.010 177.245 56.910 177.415 ;
        RECT 54.650 176.905 56.570 177.075 ;
        RECT 54.650 176.885 54.970 176.905 ;
        RECT 54.200 176.225 54.530 176.735 ;
        RECT 54.800 176.275 54.970 176.885 ;
        RECT 56.740 176.735 56.910 177.245 ;
        RECT 57.080 177.175 57.260 177.585 ;
        RECT 57.430 176.995 57.600 177.755 ;
        RECT 55.140 176.015 55.470 176.705 ;
        RECT 55.700 176.565 56.910 176.735 ;
        RECT 57.080 176.685 57.600 176.995 ;
        RECT 57.770 177.585 58.190 177.925 ;
        RECT 58.480 177.585 58.890 177.915 ;
        RECT 57.770 176.815 57.960 177.585 ;
        RECT 59.060 177.455 59.230 178.185 ;
        RECT 60.375 178.015 60.545 178.345 ;
        RECT 60.715 178.185 61.045 178.565 ;
        RECT 59.400 177.635 59.750 178.005 ;
        RECT 59.060 177.415 59.480 177.455 ;
        RECT 58.130 177.245 59.480 177.415 ;
        RECT 58.130 177.085 58.380 177.245 ;
        RECT 58.890 176.815 59.140 177.075 ;
        RECT 57.770 176.565 59.140 176.815 ;
        RECT 55.700 176.275 55.940 176.565 ;
        RECT 56.740 176.485 56.910 176.565 ;
        RECT 56.140 176.015 56.560 176.395 ;
        RECT 56.740 176.235 57.370 176.485 ;
        RECT 57.840 176.015 58.170 176.395 ;
        RECT 58.340 176.275 58.510 176.565 ;
        RECT 59.310 176.400 59.480 177.245 ;
        RECT 59.930 177.075 60.150 177.945 ;
        RECT 60.375 177.825 61.070 178.015 ;
        RECT 59.650 176.695 60.150 177.075 ;
        RECT 60.320 177.025 60.730 177.645 ;
        RECT 60.900 176.855 61.070 177.825 ;
        RECT 60.375 176.685 61.070 176.855 ;
        RECT 58.690 176.015 59.070 176.395 ;
        RECT 59.310 176.230 60.140 176.400 ;
        RECT 60.375 176.185 60.545 176.685 ;
        RECT 60.715 176.015 61.045 176.515 ;
        RECT 61.260 176.185 61.485 178.305 ;
        RECT 61.655 178.185 61.985 178.565 ;
        RECT 62.155 178.015 62.325 178.305 ;
        RECT 61.660 177.845 62.325 178.015 ;
        RECT 61.660 176.855 61.890 177.845 ;
        RECT 63.045 177.840 63.335 178.565 ;
        RECT 63.505 177.795 65.175 178.565 ;
        RECT 65.350 178.020 70.695 178.565 ;
        RECT 71.135 178.170 71.465 178.565 ;
        RECT 62.060 177.025 62.410 177.675 ;
        RECT 61.660 176.685 62.325 176.855 ;
        RECT 61.655 176.015 61.985 176.515 ;
        RECT 62.155 176.185 62.325 176.685 ;
        RECT 63.045 176.015 63.335 177.180 ;
        RECT 63.505 177.105 64.255 177.625 ;
        RECT 64.425 177.275 65.175 177.795 ;
        RECT 63.505 176.015 65.175 177.105 ;
        RECT 66.940 176.450 67.290 177.700 ;
        RECT 68.770 177.190 69.110 178.020 ;
        RECT 71.635 177.995 71.835 178.350 ;
        RECT 72.005 178.165 72.335 178.565 ;
        RECT 72.505 177.995 72.705 178.340 ;
        RECT 70.865 177.825 72.705 177.995 ;
        RECT 72.875 177.825 73.205 178.565 ;
        RECT 73.440 177.995 73.610 178.245 ;
        RECT 74.090 178.020 79.435 178.565 ;
        RECT 79.605 178.055 79.910 178.565 ;
        RECT 73.440 177.825 73.915 177.995 ;
        RECT 65.350 176.015 70.695 176.450 ;
        RECT 70.865 176.200 71.125 177.825 ;
        RECT 71.305 176.855 71.525 177.655 ;
        RECT 71.765 177.035 72.065 177.655 ;
        RECT 72.235 177.035 72.565 177.655 ;
        RECT 72.735 177.035 73.055 177.655 ;
        RECT 73.225 177.035 73.575 177.655 ;
        RECT 73.745 176.855 73.915 177.825 ;
        RECT 71.305 176.645 73.915 176.855 ;
        RECT 72.875 176.015 73.205 176.465 ;
        RECT 75.680 176.450 76.030 177.700 ;
        RECT 77.510 177.190 77.850 178.020 ;
        RECT 79.605 177.325 79.920 177.885 ;
        RECT 80.090 177.575 80.340 178.385 ;
        RECT 80.510 178.040 80.770 178.565 ;
        RECT 80.950 177.575 81.200 178.385 ;
        RECT 81.370 178.005 81.630 178.565 ;
        RECT 81.800 177.915 82.060 178.370 ;
        RECT 82.230 178.085 82.490 178.565 ;
        RECT 82.660 177.915 82.920 178.370 ;
        RECT 83.090 178.085 83.350 178.565 ;
        RECT 83.520 177.915 83.780 178.370 ;
        RECT 83.950 178.085 84.195 178.565 ;
        RECT 84.365 177.915 84.640 178.370 ;
        RECT 84.810 178.085 85.055 178.565 ;
        RECT 85.225 177.915 85.485 178.370 ;
        RECT 85.665 178.085 85.915 178.565 ;
        RECT 86.085 177.915 86.345 178.370 ;
        RECT 86.525 178.085 86.775 178.565 ;
        RECT 86.945 177.915 87.205 178.370 ;
        RECT 87.385 178.085 87.645 178.565 ;
        RECT 87.815 177.915 88.075 178.370 ;
        RECT 88.245 178.085 88.545 178.565 ;
        RECT 81.800 177.745 88.545 177.915 ;
        RECT 88.805 177.840 89.095 178.565 ;
        RECT 80.090 177.325 87.210 177.575 ;
        RECT 74.090 176.015 79.435 176.450 ;
        RECT 79.615 176.015 79.910 176.825 ;
        RECT 80.090 176.185 80.335 177.325 ;
        RECT 80.510 176.015 80.770 176.825 ;
        RECT 80.950 176.190 81.200 177.325 ;
        RECT 87.380 177.155 88.545 177.745 ;
        RECT 89.270 177.825 89.525 178.395 ;
        RECT 89.695 178.165 90.025 178.565 ;
        RECT 90.450 178.030 90.980 178.395 ;
        RECT 90.450 177.995 90.625 178.030 ;
        RECT 89.695 177.825 90.625 177.995 ;
        RECT 81.800 176.930 88.545 177.155 ;
        RECT 81.800 176.915 87.205 176.930 ;
        RECT 81.370 176.020 81.630 176.815 ;
        RECT 81.800 176.190 82.060 176.915 ;
        RECT 82.230 176.020 82.490 176.745 ;
        RECT 82.660 176.190 82.920 176.915 ;
        RECT 83.090 176.020 83.350 176.745 ;
        RECT 83.520 176.190 83.780 176.915 ;
        RECT 83.950 176.020 84.210 176.745 ;
        RECT 84.380 176.190 84.640 176.915 ;
        RECT 84.810 176.020 85.055 176.745 ;
        RECT 85.225 176.190 85.485 176.915 ;
        RECT 85.670 176.020 85.915 176.745 ;
        RECT 86.085 176.190 86.345 176.915 ;
        RECT 86.530 176.020 86.775 176.745 ;
        RECT 86.945 176.190 87.205 176.915 ;
        RECT 87.390 176.020 87.645 176.745 ;
        RECT 87.815 176.190 88.105 176.930 ;
        RECT 81.370 176.015 87.645 176.020 ;
        RECT 88.275 176.015 88.545 176.760 ;
        RECT 88.805 176.015 89.095 177.180 ;
        RECT 89.270 177.155 89.440 177.825 ;
        RECT 89.695 177.655 89.865 177.825 ;
        RECT 89.610 177.325 89.865 177.655 ;
        RECT 90.090 177.325 90.285 177.655 ;
        RECT 89.270 176.185 89.605 177.155 ;
        RECT 89.775 176.015 89.945 177.155 ;
        RECT 90.115 176.355 90.285 177.325 ;
        RECT 90.455 176.695 90.625 177.825 ;
        RECT 90.795 177.035 90.965 177.835 ;
        RECT 91.170 177.545 91.445 178.395 ;
        RECT 91.165 177.375 91.445 177.545 ;
        RECT 91.170 177.235 91.445 177.375 ;
        RECT 91.615 177.035 91.805 178.395 ;
        RECT 91.985 178.030 92.495 178.565 ;
        RECT 92.715 177.755 92.960 178.360 ;
        RECT 93.870 178.020 99.215 178.565 ;
        RECT 92.005 177.585 93.235 177.755 ;
        RECT 90.795 176.865 91.805 177.035 ;
        RECT 91.975 177.020 92.725 177.210 ;
        RECT 90.455 176.525 91.580 176.695 ;
        RECT 91.975 176.355 92.145 177.020 ;
        RECT 92.895 176.775 93.235 177.585 ;
        RECT 90.115 176.185 92.145 176.355 ;
        RECT 92.315 176.015 92.485 176.775 ;
        RECT 92.720 176.365 93.235 176.775 ;
        RECT 95.460 176.450 95.810 177.700 ;
        RECT 97.290 177.190 97.630 178.020 ;
        RECT 99.445 177.745 99.655 178.565 ;
        RECT 99.825 177.765 100.155 178.395 ;
        RECT 99.825 177.165 100.075 177.765 ;
        RECT 100.325 177.745 100.555 178.565 ;
        RECT 101.685 178.055 101.990 178.565 ;
        RECT 100.245 177.325 100.575 177.575 ;
        RECT 101.685 177.325 102.000 177.885 ;
        RECT 102.170 177.575 102.420 178.385 ;
        RECT 102.590 178.040 102.850 178.565 ;
        RECT 103.030 177.575 103.280 178.385 ;
        RECT 103.450 178.005 103.710 178.565 ;
        RECT 103.880 177.915 104.140 178.370 ;
        RECT 104.310 178.085 104.570 178.565 ;
        RECT 104.740 177.915 105.000 178.370 ;
        RECT 105.170 178.085 105.430 178.565 ;
        RECT 105.600 177.915 105.860 178.370 ;
        RECT 106.030 178.085 106.275 178.565 ;
        RECT 106.445 177.915 106.720 178.370 ;
        RECT 106.890 178.085 107.135 178.565 ;
        RECT 107.305 177.915 107.565 178.370 ;
        RECT 107.745 178.085 107.995 178.565 ;
        RECT 108.165 177.915 108.425 178.370 ;
        RECT 108.605 178.085 108.855 178.565 ;
        RECT 109.025 177.915 109.285 178.370 ;
        RECT 109.465 178.085 109.725 178.565 ;
        RECT 109.895 177.915 110.155 178.370 ;
        RECT 110.325 178.085 110.625 178.565 ;
        RECT 103.880 177.745 110.625 177.915 ;
        RECT 111.345 177.795 113.015 178.565 ;
        RECT 113.275 178.015 113.445 178.395 ;
        RECT 113.625 178.185 113.955 178.565 ;
        RECT 113.275 177.845 113.940 178.015 ;
        RECT 114.135 177.890 114.395 178.395 ;
        RECT 102.170 177.325 109.290 177.575 ;
        RECT 93.870 176.015 99.215 176.450 ;
        RECT 99.445 176.015 99.655 177.155 ;
        RECT 99.825 176.185 100.155 177.165 ;
        RECT 100.325 176.015 100.555 177.155 ;
        RECT 101.695 176.015 101.990 176.825 ;
        RECT 102.170 176.185 102.415 177.325 ;
        RECT 102.590 176.015 102.850 176.825 ;
        RECT 103.030 176.190 103.280 177.325 ;
        RECT 109.460 177.205 110.625 177.745 ;
        RECT 109.460 177.155 110.655 177.205 ;
        RECT 103.880 177.035 110.655 177.155 ;
        RECT 111.345 177.105 112.095 177.625 ;
        RECT 112.265 177.275 113.015 177.795 ;
        RECT 113.205 177.295 113.535 177.665 ;
        RECT 113.770 177.590 113.940 177.845 ;
        RECT 113.770 177.260 114.055 177.590 ;
        RECT 113.770 177.115 113.940 177.260 ;
        RECT 103.880 176.930 110.625 177.035 ;
        RECT 103.880 176.915 109.285 176.930 ;
        RECT 103.450 176.020 103.710 176.815 ;
        RECT 103.880 176.190 104.140 176.915 ;
        RECT 104.310 176.020 104.570 176.745 ;
        RECT 104.740 176.190 105.000 176.915 ;
        RECT 105.170 176.020 105.430 176.745 ;
        RECT 105.600 176.190 105.860 176.915 ;
        RECT 106.030 176.020 106.290 176.745 ;
        RECT 106.460 176.190 106.720 176.915 ;
        RECT 106.890 176.020 107.135 176.745 ;
        RECT 107.305 176.190 107.565 176.915 ;
        RECT 107.750 176.020 107.995 176.745 ;
        RECT 108.165 176.190 108.425 176.915 ;
        RECT 108.610 176.020 108.855 176.745 ;
        RECT 109.025 176.190 109.285 176.915 ;
        RECT 109.470 176.020 109.725 176.745 ;
        RECT 109.895 176.190 110.185 176.930 ;
        RECT 103.450 176.015 109.725 176.020 ;
        RECT 110.355 176.015 110.625 176.760 ;
        RECT 111.345 176.015 113.015 177.105 ;
        RECT 113.275 176.945 113.940 177.115 ;
        RECT 114.225 177.090 114.395 177.890 ;
        RECT 114.565 177.840 114.855 178.565 ;
        RECT 115.490 178.020 120.835 178.565 ;
        RECT 121.010 178.020 126.355 178.565 ;
        RECT 113.275 176.185 113.445 176.945 ;
        RECT 113.625 176.015 113.955 176.775 ;
        RECT 114.125 176.185 114.395 177.090 ;
        RECT 114.565 176.015 114.855 177.180 ;
        RECT 117.080 176.450 117.430 177.700 ;
        RECT 118.910 177.190 119.250 178.020 ;
        RECT 122.600 176.450 122.950 177.700 ;
        RECT 124.430 177.190 124.770 178.020 ;
        RECT 126.525 177.815 127.735 178.565 ;
        RECT 126.525 177.105 127.045 177.645 ;
        RECT 127.215 177.275 127.735 177.815 ;
        RECT 115.490 176.015 120.835 176.450 ;
        RECT 121.010 176.015 126.355 176.450 ;
        RECT 126.525 176.015 127.735 177.105 ;
        RECT 14.660 175.845 127.820 176.015 ;
        RECT 14.745 174.755 15.955 175.845 ;
        RECT 14.745 174.045 15.265 174.585 ;
        RECT 15.435 174.215 15.955 174.755 ;
        RECT 16.125 174.755 18.715 175.845 ;
        RECT 18.890 175.410 24.235 175.845 ;
        RECT 16.125 174.235 17.335 174.755 ;
        RECT 17.505 174.065 18.715 174.585 ;
        RECT 20.480 174.160 20.830 175.410 ;
        RECT 24.405 174.680 24.695 175.845 ;
        RECT 24.865 174.755 28.375 175.845 ;
        RECT 28.545 175.085 29.060 175.495 ;
        RECT 29.295 175.085 29.465 175.845 ;
        RECT 29.635 175.505 31.665 175.675 ;
        RECT 14.745 173.295 15.955 174.045 ;
        RECT 16.125 173.295 18.715 174.065 ;
        RECT 22.310 173.840 22.650 174.670 ;
        RECT 24.865 174.235 26.555 174.755 ;
        RECT 26.725 174.065 28.375 174.585 ;
        RECT 28.545 174.275 28.885 175.085 ;
        RECT 29.635 174.840 29.805 175.505 ;
        RECT 30.200 175.165 31.325 175.335 ;
        RECT 29.055 174.650 29.805 174.840 ;
        RECT 29.975 174.825 30.985 174.995 ;
        RECT 28.545 174.105 29.775 174.275 ;
        RECT 18.890 173.295 24.235 173.840 ;
        RECT 24.405 173.295 24.695 174.020 ;
        RECT 24.865 173.295 28.375 174.065 ;
        RECT 28.820 173.500 29.065 174.105 ;
        RECT 29.285 173.295 29.795 173.830 ;
        RECT 29.975 173.465 30.165 174.825 ;
        RECT 30.335 174.485 30.610 174.625 ;
        RECT 30.335 174.315 30.615 174.485 ;
        RECT 30.335 173.465 30.610 174.315 ;
        RECT 30.815 174.025 30.985 174.825 ;
        RECT 31.155 174.035 31.325 175.165 ;
        RECT 31.495 174.535 31.665 175.505 ;
        RECT 31.835 174.705 32.005 175.845 ;
        RECT 32.175 174.705 32.510 175.675 ;
        RECT 31.495 174.205 31.690 174.535 ;
        RECT 31.915 174.205 32.170 174.535 ;
        RECT 31.915 174.035 32.085 174.205 ;
        RECT 32.340 174.035 32.510 174.705 ;
        RECT 32.685 174.755 33.895 175.845 ;
        RECT 32.685 174.215 33.205 174.755 ;
        RECT 34.105 174.705 34.335 175.845 ;
        RECT 34.505 174.695 34.835 175.675 ;
        RECT 35.005 174.705 35.215 175.845 ;
        RECT 33.375 174.045 33.895 174.585 ;
        RECT 34.085 174.285 34.415 174.535 ;
        RECT 31.155 173.865 32.085 174.035 ;
        RECT 31.155 173.830 31.330 173.865 ;
        RECT 30.800 173.465 31.330 173.830 ;
        RECT 31.755 173.295 32.085 173.695 ;
        RECT 32.255 173.465 32.510 174.035 ;
        RECT 32.685 173.295 33.895 174.045 ;
        RECT 34.105 173.295 34.335 174.115 ;
        RECT 34.585 174.095 34.835 174.695 ;
        RECT 35.450 174.655 35.705 175.535 ;
        RECT 35.875 174.705 36.180 175.845 ;
        RECT 36.520 175.465 36.850 175.845 ;
        RECT 37.030 175.295 37.200 175.585 ;
        RECT 37.370 175.385 37.620 175.845 ;
        RECT 36.400 175.125 37.200 175.295 ;
        RECT 37.790 175.335 38.660 175.675 ;
        RECT 34.505 173.465 34.835 174.095 ;
        RECT 35.005 173.295 35.215 174.115 ;
        RECT 35.450 174.005 35.660 174.655 ;
        RECT 36.400 174.535 36.570 175.125 ;
        RECT 37.790 174.955 37.960 175.335 ;
        RECT 38.895 175.215 39.065 175.675 ;
        RECT 39.235 175.385 39.605 175.845 ;
        RECT 39.900 175.245 40.070 175.585 ;
        RECT 40.240 175.415 40.570 175.845 ;
        RECT 40.805 175.245 40.975 175.585 ;
        RECT 36.740 174.785 37.960 174.955 ;
        RECT 38.130 174.875 38.590 175.165 ;
        RECT 38.895 175.045 39.455 175.215 ;
        RECT 39.900 175.075 40.975 175.245 ;
        RECT 41.145 175.345 41.825 175.675 ;
        RECT 42.040 175.345 42.290 175.675 ;
        RECT 42.460 175.385 42.710 175.845 ;
        RECT 39.285 174.905 39.455 175.045 ;
        RECT 38.130 174.865 39.095 174.875 ;
        RECT 37.790 174.695 37.960 174.785 ;
        RECT 38.420 174.705 39.095 174.865 ;
        RECT 35.830 174.505 36.570 174.535 ;
        RECT 35.830 174.205 36.745 174.505 ;
        RECT 36.420 174.030 36.745 174.205 ;
        RECT 35.450 173.475 35.705 174.005 ;
        RECT 35.875 173.295 36.180 173.755 ;
        RECT 36.425 173.675 36.745 174.030 ;
        RECT 36.915 174.245 37.455 174.615 ;
        RECT 37.790 174.525 38.195 174.695 ;
        RECT 36.915 173.845 37.155 174.245 ;
        RECT 37.635 174.075 37.855 174.355 ;
        RECT 37.325 173.905 37.855 174.075 ;
        RECT 37.325 173.675 37.495 173.905 ;
        RECT 38.025 173.745 38.195 174.525 ;
        RECT 38.365 173.915 38.715 174.535 ;
        RECT 38.885 173.915 39.095 174.705 ;
        RECT 39.285 174.735 40.785 174.905 ;
        RECT 39.285 174.045 39.455 174.735 ;
        RECT 41.145 174.565 41.315 175.345 ;
        RECT 42.120 175.215 42.290 175.345 ;
        RECT 39.625 174.395 41.315 174.565 ;
        RECT 41.485 174.785 41.950 175.175 ;
        RECT 42.120 175.045 42.515 175.215 ;
        RECT 39.625 174.215 39.795 174.395 ;
        RECT 36.425 173.505 37.495 173.675 ;
        RECT 37.665 173.295 37.855 173.735 ;
        RECT 38.025 173.465 38.975 173.745 ;
        RECT 39.285 173.655 39.545 174.045 ;
        RECT 39.965 173.975 40.755 174.225 ;
        RECT 39.195 173.485 39.545 173.655 ;
        RECT 39.755 173.295 40.085 173.755 ;
        RECT 40.960 173.685 41.130 174.395 ;
        RECT 41.485 174.195 41.655 174.785 ;
        RECT 41.300 173.975 41.655 174.195 ;
        RECT 41.825 173.975 42.175 174.595 ;
        RECT 42.345 173.685 42.515 175.045 ;
        RECT 42.880 174.875 43.205 175.660 ;
        RECT 42.685 173.825 43.145 174.875 ;
        RECT 40.960 173.515 41.815 173.685 ;
        RECT 42.020 173.515 42.515 173.685 ;
        RECT 42.685 173.295 43.015 173.655 ;
        RECT 43.375 173.555 43.545 175.675 ;
        RECT 43.715 175.345 44.045 175.845 ;
        RECT 44.215 175.175 44.470 175.675 ;
        RECT 43.720 175.005 44.470 175.175 ;
        RECT 45.565 175.085 46.080 175.495 ;
        RECT 46.315 175.085 46.485 175.845 ;
        RECT 46.655 175.505 48.685 175.675 ;
        RECT 43.720 174.015 43.950 175.005 ;
        RECT 44.120 174.185 44.470 174.835 ;
        RECT 45.565 174.275 45.905 175.085 ;
        RECT 46.655 174.840 46.825 175.505 ;
        RECT 47.220 175.165 48.345 175.335 ;
        RECT 46.075 174.650 46.825 174.840 ;
        RECT 46.995 174.825 48.005 174.995 ;
        RECT 45.565 174.105 46.795 174.275 ;
        RECT 43.720 173.845 44.470 174.015 ;
        RECT 43.715 173.295 44.045 173.675 ;
        RECT 44.215 173.555 44.470 173.845 ;
        RECT 45.840 173.500 46.085 174.105 ;
        RECT 46.305 173.295 46.815 173.830 ;
        RECT 46.995 173.465 47.185 174.825 ;
        RECT 47.355 174.485 47.630 174.625 ;
        RECT 47.355 174.315 47.635 174.485 ;
        RECT 47.355 173.465 47.630 174.315 ;
        RECT 47.835 174.025 48.005 174.825 ;
        RECT 48.175 174.035 48.345 175.165 ;
        RECT 48.515 174.535 48.685 175.505 ;
        RECT 48.855 174.705 49.025 175.845 ;
        RECT 49.195 174.705 49.530 175.675 ;
        RECT 48.515 174.205 48.710 174.535 ;
        RECT 48.935 174.205 49.190 174.535 ;
        RECT 48.935 174.035 49.105 174.205 ;
        RECT 49.360 174.035 49.530 174.705 ;
        RECT 50.165 174.680 50.455 175.845 ;
        RECT 50.715 174.915 50.885 175.675 ;
        RECT 51.065 175.085 51.395 175.845 ;
        RECT 50.715 174.745 51.380 174.915 ;
        RECT 51.565 174.770 51.835 175.675 ;
        RECT 51.210 174.600 51.380 174.745 ;
        RECT 50.645 174.195 50.975 174.565 ;
        RECT 51.210 174.270 51.495 174.600 ;
        RECT 48.175 173.865 49.105 174.035 ;
        RECT 48.175 173.830 48.350 173.865 ;
        RECT 47.820 173.465 48.350 173.830 ;
        RECT 48.775 173.295 49.105 173.695 ;
        RECT 49.275 173.465 49.530 174.035 ;
        RECT 50.165 173.295 50.455 174.020 ;
        RECT 51.210 174.015 51.380 174.270 ;
        RECT 50.715 173.845 51.380 174.015 ;
        RECT 51.665 173.970 51.835 174.770 ;
        RECT 52.005 174.755 53.215 175.845 ;
        RECT 53.385 175.085 53.900 175.495 ;
        RECT 54.135 175.085 54.305 175.845 ;
        RECT 54.475 175.505 56.505 175.675 ;
        RECT 52.005 174.215 52.525 174.755 ;
        RECT 52.695 174.045 53.215 174.585 ;
        RECT 53.385 174.275 53.725 175.085 ;
        RECT 54.475 174.840 54.645 175.505 ;
        RECT 55.040 175.165 56.165 175.335 ;
        RECT 53.895 174.650 54.645 174.840 ;
        RECT 54.815 174.825 55.825 174.995 ;
        RECT 53.385 174.105 54.615 174.275 ;
        RECT 50.715 173.465 50.885 173.845 ;
        RECT 51.065 173.295 51.395 173.675 ;
        RECT 51.575 173.465 51.835 173.970 ;
        RECT 52.005 173.295 53.215 174.045 ;
        RECT 53.660 173.500 53.905 174.105 ;
        RECT 54.125 173.295 54.635 173.830 ;
        RECT 54.815 173.465 55.005 174.825 ;
        RECT 55.175 174.145 55.450 174.625 ;
        RECT 55.175 173.975 55.455 174.145 ;
        RECT 55.655 174.025 55.825 174.825 ;
        RECT 55.995 174.035 56.165 175.165 ;
        RECT 56.335 174.535 56.505 175.505 ;
        RECT 56.675 174.705 56.845 175.845 ;
        RECT 57.015 174.705 57.350 175.675 ;
        RECT 56.335 174.205 56.530 174.535 ;
        RECT 56.755 174.205 57.010 174.535 ;
        RECT 56.755 174.035 56.925 174.205 ;
        RECT 57.180 174.035 57.350 174.705 ;
        RECT 57.985 174.755 61.495 175.845 ;
        RECT 61.670 175.410 67.015 175.845 ;
        RECT 57.985 174.235 59.675 174.755 ;
        RECT 59.845 174.065 61.495 174.585 ;
        RECT 63.260 174.160 63.610 175.410 ;
        RECT 55.175 173.465 55.450 173.975 ;
        RECT 55.995 173.865 56.925 174.035 ;
        RECT 55.995 173.830 56.170 173.865 ;
        RECT 55.640 173.465 56.170 173.830 ;
        RECT 56.595 173.295 56.925 173.695 ;
        RECT 57.095 173.465 57.350 174.035 ;
        RECT 57.985 173.295 61.495 174.065 ;
        RECT 65.090 173.840 65.430 174.670 ;
        RECT 67.185 174.035 67.445 175.660 ;
        RECT 69.195 175.395 69.525 175.845 ;
        RECT 70.405 175.345 70.665 175.675 ;
        RECT 70.975 175.465 71.305 175.845 ;
        RECT 67.625 175.005 70.235 175.215 ;
        RECT 67.625 174.205 67.845 175.005 ;
        RECT 68.085 174.205 68.385 174.825 ;
        RECT 68.555 174.205 68.885 174.825 ;
        RECT 69.055 174.205 69.375 174.825 ;
        RECT 69.545 174.205 69.895 174.825 ;
        RECT 70.065 174.035 70.235 175.005 ;
        RECT 67.185 173.865 69.025 174.035 ;
        RECT 61.670 173.295 67.015 173.840 ;
        RECT 67.455 173.295 67.785 173.690 ;
        RECT 67.955 173.510 68.155 173.865 ;
        RECT 68.325 173.295 68.655 173.695 ;
        RECT 68.825 173.520 69.025 173.865 ;
        RECT 69.195 173.295 69.525 174.035 ;
        RECT 69.760 173.865 70.235 174.035 ;
        RECT 70.405 174.665 70.575 175.345 ;
        RECT 71.545 175.295 71.735 175.675 ;
        RECT 71.985 175.465 72.315 175.845 ;
        RECT 72.525 175.295 72.695 175.675 ;
        RECT 72.890 175.465 73.220 175.845 ;
        RECT 73.480 175.295 73.650 175.675 ;
        RECT 74.075 175.465 74.405 175.845 ;
        RECT 70.745 174.835 71.095 175.165 ;
        RECT 71.545 175.125 72.285 175.295 ;
        RECT 71.365 174.785 71.945 174.955 ;
        RECT 71.365 174.665 71.535 174.785 ;
        RECT 70.405 174.495 71.535 174.665 ;
        RECT 72.115 174.615 72.285 175.125 ;
        RECT 69.760 173.615 69.930 173.865 ;
        RECT 70.405 173.795 70.575 174.495 ;
        RECT 71.715 174.445 72.285 174.615 ;
        RECT 72.455 175.125 74.405 175.295 ;
        RECT 70.925 174.155 71.545 174.325 ;
        RECT 70.925 173.975 71.135 174.155 ;
        RECT 71.715 173.965 71.885 174.445 ;
        RECT 72.455 174.135 72.625 175.125 ;
        RECT 73.215 174.535 73.400 174.845 ;
        RECT 73.670 174.535 73.865 174.845 ;
        RECT 70.405 173.465 70.665 173.795 ;
        RECT 70.975 173.295 71.305 173.675 ;
        RECT 71.485 173.635 71.885 173.965 ;
        RECT 72.075 173.805 72.625 174.135 ;
        RECT 72.795 173.635 72.965 174.535 ;
        RECT 71.485 173.465 72.965 173.635 ;
        RECT 73.215 174.205 73.445 174.535 ;
        RECT 73.670 174.205 73.925 174.535 ;
        RECT 74.235 174.205 74.405 175.125 ;
        RECT 73.215 173.625 73.400 174.205 ;
        RECT 73.670 173.630 73.865 174.205 ;
        RECT 74.075 173.295 74.405 173.675 ;
        RECT 74.575 173.465 74.835 175.675 ;
        RECT 75.925 174.680 76.215 175.845 ;
        RECT 77.095 175.395 77.425 175.845 ;
        RECT 76.385 175.005 78.995 175.215 ;
        RECT 76.385 174.035 76.555 175.005 ;
        RECT 76.725 174.205 77.075 174.825 ;
        RECT 77.245 174.205 77.565 174.825 ;
        RECT 77.735 174.205 78.065 174.825 ;
        RECT 78.235 174.205 78.535 174.825 ;
        RECT 78.775 174.205 78.995 175.005 ;
        RECT 79.175 174.035 79.435 175.660 ;
        RECT 75.925 173.295 76.215 174.020 ;
        RECT 76.385 173.865 76.860 174.035 ;
        RECT 76.690 173.615 76.860 173.865 ;
        RECT 77.095 173.295 77.425 174.035 ;
        RECT 77.595 173.865 79.435 174.035 ;
        RECT 79.605 174.875 79.915 175.675 ;
        RECT 80.085 175.045 80.395 175.845 ;
        RECT 80.565 175.215 80.825 175.675 ;
        RECT 80.995 175.385 81.250 175.845 ;
        RECT 81.425 175.215 81.685 175.675 ;
        RECT 80.565 175.045 81.685 175.215 ;
        RECT 79.605 174.705 80.635 174.875 ;
        RECT 77.595 173.520 77.795 173.865 ;
        RECT 77.965 173.295 78.295 173.695 ;
        RECT 78.465 173.510 78.665 173.865 ;
        RECT 79.605 173.795 79.775 174.705 ;
        RECT 79.945 173.965 80.295 174.535 ;
        RECT 80.465 174.455 80.635 174.705 ;
        RECT 81.425 174.795 81.685 175.045 ;
        RECT 81.855 174.975 82.140 175.845 ;
        RECT 81.425 174.625 82.180 174.795 ;
        RECT 80.465 174.285 81.605 174.455 ;
        RECT 81.775 174.115 82.180 174.625 ;
        RECT 82.825 174.755 85.415 175.845 ;
        RECT 85.675 174.915 85.845 175.675 ;
        RECT 86.025 175.085 86.355 175.845 ;
        RECT 82.825 174.235 84.035 174.755 ;
        RECT 85.675 174.745 86.340 174.915 ;
        RECT 86.525 174.770 86.795 175.675 ;
        RECT 86.170 174.600 86.340 174.745 ;
        RECT 80.530 173.945 82.180 174.115 ;
        RECT 84.205 174.065 85.415 174.585 ;
        RECT 85.605 174.195 85.935 174.565 ;
        RECT 86.170 174.270 86.455 174.600 ;
        RECT 78.835 173.295 79.165 173.690 ;
        RECT 79.605 173.465 79.905 173.795 ;
        RECT 80.075 173.295 80.350 173.775 ;
        RECT 80.530 173.555 80.825 173.945 ;
        RECT 80.995 173.295 81.250 173.775 ;
        RECT 81.425 173.555 81.685 173.945 ;
        RECT 81.855 173.295 82.135 173.775 ;
        RECT 82.825 173.295 85.415 174.065 ;
        RECT 86.170 174.015 86.340 174.270 ;
        RECT 85.675 173.845 86.340 174.015 ;
        RECT 86.625 173.970 86.795 174.770 ;
        RECT 87.025 174.705 87.235 175.845 ;
        RECT 87.405 174.695 87.735 175.675 ;
        RECT 87.905 174.705 88.135 175.845 ;
        RECT 89.320 174.975 89.605 175.845 ;
        RECT 89.775 175.215 90.035 175.675 ;
        RECT 90.210 175.385 90.465 175.845 ;
        RECT 90.635 175.215 90.895 175.675 ;
        RECT 89.775 175.045 90.895 175.215 ;
        RECT 91.065 175.045 91.375 175.845 ;
        RECT 89.775 174.795 90.035 175.045 ;
        RECT 91.545 174.875 91.855 175.675 ;
        RECT 92.490 175.175 92.745 175.675 ;
        RECT 92.915 175.345 93.245 175.845 ;
        RECT 92.490 175.005 93.240 175.175 ;
        RECT 85.675 173.465 85.845 173.845 ;
        RECT 86.025 173.295 86.355 173.675 ;
        RECT 86.535 173.465 86.795 173.970 ;
        RECT 87.025 173.295 87.235 174.115 ;
        RECT 87.405 174.095 87.655 174.695 ;
        RECT 89.280 174.625 90.035 174.795 ;
        RECT 90.825 174.705 91.855 174.875 ;
        RECT 87.825 174.285 88.155 174.535 ;
        RECT 89.280 174.115 89.685 174.625 ;
        RECT 90.825 174.455 90.995 174.705 ;
        RECT 89.855 174.285 90.995 174.455 ;
        RECT 87.405 173.465 87.735 174.095 ;
        RECT 87.905 173.295 88.135 174.115 ;
        RECT 89.280 173.945 90.930 174.115 ;
        RECT 91.165 173.965 91.515 174.535 ;
        RECT 89.325 173.295 89.605 173.775 ;
        RECT 89.775 173.555 90.035 173.945 ;
        RECT 90.210 173.295 90.465 173.775 ;
        RECT 90.635 173.555 90.930 173.945 ;
        RECT 91.685 173.795 91.855 174.705 ;
        RECT 92.490 174.185 92.840 174.835 ;
        RECT 93.010 174.015 93.240 175.005 ;
        RECT 91.110 173.295 91.385 173.775 ;
        RECT 91.555 173.465 91.855 173.795 ;
        RECT 92.490 173.845 93.240 174.015 ;
        RECT 92.490 173.555 92.745 173.845 ;
        RECT 92.915 173.295 93.245 173.675 ;
        RECT 93.415 173.555 93.585 175.675 ;
        RECT 93.755 174.875 94.080 175.660 ;
        RECT 94.250 175.385 94.500 175.845 ;
        RECT 94.670 175.345 94.920 175.675 ;
        RECT 95.135 175.345 95.815 175.675 ;
        RECT 94.670 175.215 94.840 175.345 ;
        RECT 94.445 175.045 94.840 175.215 ;
        RECT 93.815 173.825 94.275 174.875 ;
        RECT 94.445 173.685 94.615 175.045 ;
        RECT 95.010 174.785 95.475 175.175 ;
        RECT 94.785 173.975 95.135 174.595 ;
        RECT 95.305 174.195 95.475 174.785 ;
        RECT 95.645 174.565 95.815 175.345 ;
        RECT 95.985 175.245 96.155 175.585 ;
        RECT 96.390 175.415 96.720 175.845 ;
        RECT 96.890 175.245 97.060 175.585 ;
        RECT 97.355 175.385 97.725 175.845 ;
        RECT 95.985 175.075 97.060 175.245 ;
        RECT 97.895 175.215 98.065 175.675 ;
        RECT 98.300 175.335 99.170 175.675 ;
        RECT 99.340 175.385 99.590 175.845 ;
        RECT 97.505 175.045 98.065 175.215 ;
        RECT 97.505 174.905 97.675 175.045 ;
        RECT 96.175 174.735 97.675 174.905 ;
        RECT 98.370 174.875 98.830 175.165 ;
        RECT 95.645 174.395 97.335 174.565 ;
        RECT 95.305 173.975 95.660 174.195 ;
        RECT 95.830 173.685 96.000 174.395 ;
        RECT 96.205 173.975 96.995 174.225 ;
        RECT 97.165 174.215 97.335 174.395 ;
        RECT 97.505 174.045 97.675 174.735 ;
        RECT 93.945 173.295 94.275 173.655 ;
        RECT 94.445 173.515 94.940 173.685 ;
        RECT 95.145 173.515 96.000 173.685 ;
        RECT 96.875 173.295 97.205 173.755 ;
        RECT 97.415 173.655 97.675 174.045 ;
        RECT 97.865 174.865 98.830 174.875 ;
        RECT 99.000 174.955 99.170 175.335 ;
        RECT 99.760 175.295 99.930 175.585 ;
        RECT 100.110 175.465 100.440 175.845 ;
        RECT 99.760 175.125 100.560 175.295 ;
        RECT 97.865 174.705 98.540 174.865 ;
        RECT 99.000 174.785 100.220 174.955 ;
        RECT 97.865 173.915 98.075 174.705 ;
        RECT 99.000 174.695 99.170 174.785 ;
        RECT 98.245 173.915 98.595 174.535 ;
        RECT 98.765 174.525 99.170 174.695 ;
        RECT 98.765 173.745 98.935 174.525 ;
        RECT 99.105 174.075 99.325 174.355 ;
        RECT 99.505 174.245 100.045 174.615 ;
        RECT 100.390 174.535 100.560 175.125 ;
        RECT 100.780 174.705 101.085 175.845 ;
        RECT 101.255 174.655 101.510 175.535 ;
        RECT 101.685 174.680 101.975 175.845 ;
        RECT 102.255 175.045 102.425 175.845 ;
        RECT 102.595 174.825 102.925 175.675 ;
        RECT 103.095 175.045 103.265 175.845 ;
        RECT 103.435 174.825 103.765 175.675 ;
        RECT 103.935 175.045 104.105 175.845 ;
        RECT 104.275 174.825 104.605 175.675 ;
        RECT 104.775 175.045 104.945 175.845 ;
        RECT 105.115 174.825 105.445 175.675 ;
        RECT 105.615 175.045 105.785 175.845 ;
        RECT 105.955 174.825 106.285 175.675 ;
        RECT 106.455 175.045 106.625 175.845 ;
        RECT 106.795 174.825 107.125 175.675 ;
        RECT 107.295 175.045 107.465 175.845 ;
        RECT 107.635 174.825 107.965 175.675 ;
        RECT 108.135 175.045 108.305 175.845 ;
        RECT 108.475 174.825 108.805 175.675 ;
        RECT 108.975 175.045 109.145 175.845 ;
        RECT 109.315 174.825 109.645 175.675 ;
        RECT 109.815 175.045 109.985 175.845 ;
        RECT 110.155 174.825 110.485 175.675 ;
        RECT 110.655 175.045 110.825 175.845 ;
        RECT 110.995 174.825 111.325 175.675 ;
        RECT 111.495 174.995 111.665 175.845 ;
        RECT 111.835 174.825 112.165 175.675 ;
        RECT 112.335 174.995 112.505 175.845 ;
        RECT 112.675 174.825 113.005 175.675 ;
        RECT 100.390 174.505 101.130 174.535 ;
        RECT 99.105 173.905 99.635 174.075 ;
        RECT 97.415 173.485 97.765 173.655 ;
        RECT 97.985 173.465 98.935 173.745 ;
        RECT 99.105 173.295 99.295 173.735 ;
        RECT 99.465 173.675 99.635 173.905 ;
        RECT 99.805 173.845 100.045 174.245 ;
        RECT 100.215 174.205 101.130 174.505 ;
        RECT 100.215 174.030 100.540 174.205 ;
        RECT 100.215 173.675 100.535 174.030 ;
        RECT 101.300 174.005 101.510 174.655 ;
        RECT 102.145 174.655 108.805 174.825 ;
        RECT 108.975 174.655 111.325 174.825 ;
        RECT 111.495 174.655 113.005 174.825 ;
        RECT 113.645 174.755 115.315 175.845 ;
        RECT 115.485 175.085 116.000 175.495 ;
        RECT 116.235 175.085 116.405 175.845 ;
        RECT 116.575 175.505 118.605 175.675 ;
        RECT 102.145 174.115 102.420 174.655 ;
        RECT 108.975 174.485 109.150 174.655 ;
        RECT 111.495 174.485 111.665 174.655 ;
        RECT 102.590 174.285 109.150 174.485 ;
        RECT 109.355 174.285 111.665 174.485 ;
        RECT 111.835 174.285 113.010 174.485 ;
        RECT 108.975 174.115 109.150 174.285 ;
        RECT 111.495 174.115 111.665 174.285 ;
        RECT 113.645 174.235 114.395 174.755 ;
        RECT 99.465 173.505 100.535 173.675 ;
        RECT 100.780 173.295 101.085 173.755 ;
        RECT 101.255 173.475 101.510 174.005 ;
        RECT 101.685 173.295 101.975 174.020 ;
        RECT 102.145 173.945 108.805 174.115 ;
        RECT 108.975 173.945 111.325 174.115 ;
        RECT 111.495 173.945 113.005 174.115 ;
        RECT 114.565 174.065 115.315 174.585 ;
        RECT 115.485 174.275 115.825 175.085 ;
        RECT 116.575 174.840 116.745 175.505 ;
        RECT 117.140 175.165 118.265 175.335 ;
        RECT 115.995 174.650 116.745 174.840 ;
        RECT 116.915 174.825 117.925 174.995 ;
        RECT 115.485 174.105 116.715 174.275 ;
        RECT 102.255 173.295 102.425 173.775 ;
        RECT 102.595 173.470 102.925 173.945 ;
        RECT 103.095 173.295 103.265 173.775 ;
        RECT 103.435 173.470 103.765 173.945 ;
        RECT 103.935 173.295 104.105 173.775 ;
        RECT 104.275 173.470 104.605 173.945 ;
        RECT 104.775 173.295 104.945 173.775 ;
        RECT 105.115 173.470 105.445 173.945 ;
        RECT 105.615 173.295 105.785 173.775 ;
        RECT 105.955 173.470 106.285 173.945 ;
        RECT 106.455 173.295 106.625 173.775 ;
        RECT 106.795 173.470 107.125 173.945 ;
        RECT 106.875 173.465 107.045 173.470 ;
        RECT 107.295 173.295 107.465 173.775 ;
        RECT 107.635 173.470 107.965 173.945 ;
        RECT 107.715 173.465 107.885 173.470 ;
        RECT 108.135 173.295 108.305 173.775 ;
        RECT 108.475 173.470 108.805 173.945 ;
        RECT 108.555 173.465 108.805 173.470 ;
        RECT 108.975 173.295 109.145 173.775 ;
        RECT 109.315 173.470 109.645 173.945 ;
        RECT 109.815 173.295 109.985 173.775 ;
        RECT 110.155 173.470 110.485 173.945 ;
        RECT 110.655 173.295 110.825 173.775 ;
        RECT 110.995 173.470 111.325 173.945 ;
        RECT 111.495 173.295 111.665 173.775 ;
        RECT 111.835 173.470 112.165 173.945 ;
        RECT 112.335 173.295 112.505 173.775 ;
        RECT 112.675 173.470 113.005 173.945 ;
        RECT 113.645 173.295 115.315 174.065 ;
        RECT 115.760 173.500 116.005 174.105 ;
        RECT 116.225 173.295 116.735 173.830 ;
        RECT 116.915 173.465 117.105 174.825 ;
        RECT 117.275 174.485 117.550 174.625 ;
        RECT 117.275 174.315 117.555 174.485 ;
        RECT 117.275 173.465 117.550 174.315 ;
        RECT 117.755 174.025 117.925 174.825 ;
        RECT 118.095 174.035 118.265 175.165 ;
        RECT 118.435 174.535 118.605 175.505 ;
        RECT 118.775 174.705 118.945 175.845 ;
        RECT 119.115 174.705 119.450 175.675 ;
        RECT 119.665 174.705 119.895 175.845 ;
        RECT 118.435 174.205 118.630 174.535 ;
        RECT 118.855 174.205 119.110 174.535 ;
        RECT 118.855 174.035 119.025 174.205 ;
        RECT 119.280 174.035 119.450 174.705 ;
        RECT 120.065 174.695 120.395 175.675 ;
        RECT 120.565 174.705 120.775 175.845 ;
        RECT 122.015 174.915 122.185 175.675 ;
        RECT 122.365 175.085 122.695 175.845 ;
        RECT 122.015 174.745 122.680 174.915 ;
        RECT 122.865 174.770 123.135 175.675 ;
        RECT 119.645 174.285 119.975 174.535 ;
        RECT 118.095 173.865 119.025 174.035 ;
        RECT 118.095 173.830 118.270 173.865 ;
        RECT 117.740 173.465 118.270 173.830 ;
        RECT 118.695 173.295 119.025 173.695 ;
        RECT 119.195 173.465 119.450 174.035 ;
        RECT 119.665 173.295 119.895 174.115 ;
        RECT 120.145 174.095 120.395 174.695 ;
        RECT 122.510 174.600 122.680 174.745 ;
        RECT 121.945 174.195 122.275 174.565 ;
        RECT 122.510 174.270 122.795 174.600 ;
        RECT 120.065 173.465 120.395 174.095 ;
        RECT 120.565 173.295 120.775 174.115 ;
        RECT 122.510 174.015 122.680 174.270 ;
        RECT 122.015 173.845 122.680 174.015 ;
        RECT 122.965 173.970 123.135 174.770 ;
        RECT 123.765 174.755 126.355 175.845 ;
        RECT 126.525 174.755 127.735 175.845 ;
        RECT 123.765 174.235 124.975 174.755 ;
        RECT 125.145 174.065 126.355 174.585 ;
        RECT 126.525 174.215 127.045 174.755 ;
        RECT 122.015 173.465 122.185 173.845 ;
        RECT 122.365 173.295 122.695 173.675 ;
        RECT 122.875 173.465 123.135 173.970 ;
        RECT 123.765 173.295 126.355 174.065 ;
        RECT 127.215 174.045 127.735 174.585 ;
        RECT 126.525 173.295 127.735 174.045 ;
        RECT 14.660 173.125 127.820 173.295 ;
        RECT 14.745 172.375 15.955 173.125 ;
        RECT 16.590 172.580 21.935 173.125 ;
        RECT 14.745 171.835 15.265 172.375 ;
        RECT 15.435 171.665 15.955 172.205 ;
        RECT 14.745 170.575 15.955 171.665 ;
        RECT 18.180 171.010 18.530 172.260 ;
        RECT 20.010 171.750 20.350 172.580 ;
        RECT 22.145 172.305 22.375 173.125 ;
        RECT 22.545 172.325 22.875 172.955 ;
        RECT 22.125 171.885 22.455 172.135 ;
        RECT 22.625 171.725 22.875 172.325 ;
        RECT 23.045 172.305 23.255 173.125 ;
        RECT 23.490 172.415 23.745 172.945 ;
        RECT 23.915 172.665 24.220 173.125 ;
        RECT 24.465 172.745 25.535 172.915 ;
        RECT 16.590 170.575 21.935 171.010 ;
        RECT 22.145 170.575 22.375 171.715 ;
        RECT 22.545 170.745 22.875 171.725 ;
        RECT 23.490 171.765 23.700 172.415 ;
        RECT 24.465 172.390 24.785 172.745 ;
        RECT 24.460 172.215 24.785 172.390 ;
        RECT 23.870 171.915 24.785 172.215 ;
        RECT 24.955 172.175 25.195 172.575 ;
        RECT 25.365 172.515 25.535 172.745 ;
        RECT 25.705 172.685 25.895 173.125 ;
        RECT 26.065 172.675 27.015 172.955 ;
        RECT 27.235 172.765 27.585 172.935 ;
        RECT 25.365 172.345 25.895 172.515 ;
        RECT 23.870 171.885 24.610 171.915 ;
        RECT 23.045 170.575 23.255 171.715 ;
        RECT 23.490 170.885 23.745 171.765 ;
        RECT 23.915 170.575 24.220 171.715 ;
        RECT 24.440 171.295 24.610 171.885 ;
        RECT 24.955 171.805 25.495 172.175 ;
        RECT 25.675 172.065 25.895 172.345 ;
        RECT 26.065 171.895 26.235 172.675 ;
        RECT 25.830 171.725 26.235 171.895 ;
        RECT 26.405 171.885 26.755 172.505 ;
        RECT 25.830 171.635 26.000 171.725 ;
        RECT 26.925 171.715 27.135 172.505 ;
        RECT 24.780 171.465 26.000 171.635 ;
        RECT 26.460 171.555 27.135 171.715 ;
        RECT 24.440 171.125 25.240 171.295 ;
        RECT 24.560 170.575 24.890 170.955 ;
        RECT 25.070 170.835 25.240 171.125 ;
        RECT 25.830 171.085 26.000 171.465 ;
        RECT 26.170 171.545 27.135 171.555 ;
        RECT 27.325 172.375 27.585 172.765 ;
        RECT 27.795 172.665 28.125 173.125 ;
        RECT 29.000 172.735 29.855 172.905 ;
        RECT 30.060 172.735 30.555 172.905 ;
        RECT 30.725 172.765 31.055 173.125 ;
        RECT 27.325 171.685 27.495 172.375 ;
        RECT 27.665 172.025 27.835 172.205 ;
        RECT 28.005 172.195 28.795 172.445 ;
        RECT 29.000 172.025 29.170 172.735 ;
        RECT 29.340 172.225 29.695 172.445 ;
        RECT 27.665 171.855 29.355 172.025 ;
        RECT 26.170 171.255 26.630 171.545 ;
        RECT 27.325 171.515 28.825 171.685 ;
        RECT 27.325 171.375 27.495 171.515 ;
        RECT 26.935 171.205 27.495 171.375 ;
        RECT 25.410 170.575 25.660 171.035 ;
        RECT 25.830 170.745 26.700 171.085 ;
        RECT 26.935 170.745 27.105 171.205 ;
        RECT 27.940 171.175 29.015 171.345 ;
        RECT 27.275 170.575 27.645 171.035 ;
        RECT 27.940 170.835 28.110 171.175 ;
        RECT 28.280 170.575 28.610 171.005 ;
        RECT 28.845 170.835 29.015 171.175 ;
        RECT 29.185 171.075 29.355 171.855 ;
        RECT 29.525 171.635 29.695 172.225 ;
        RECT 29.865 171.825 30.215 172.445 ;
        RECT 29.525 171.245 29.990 171.635 ;
        RECT 30.385 171.375 30.555 172.735 ;
        RECT 30.725 171.545 31.185 172.595 ;
        RECT 30.160 171.205 30.555 171.375 ;
        RECT 30.160 171.075 30.330 171.205 ;
        RECT 29.185 170.745 29.865 171.075 ;
        RECT 30.080 170.745 30.330 171.075 ;
        RECT 30.500 170.575 30.750 171.035 ;
        RECT 30.920 170.760 31.245 171.545 ;
        RECT 31.415 170.745 31.585 172.865 ;
        RECT 31.755 172.745 32.085 173.125 ;
        RECT 32.255 172.575 32.510 172.865 ;
        RECT 31.760 172.405 32.510 172.575 ;
        RECT 32.685 172.450 32.945 172.955 ;
        RECT 33.125 172.745 33.455 173.125 ;
        RECT 33.635 172.575 33.805 172.955 ;
        RECT 31.760 171.415 31.990 172.405 ;
        RECT 32.160 171.585 32.510 172.235 ;
        RECT 32.685 171.650 32.855 172.450 ;
        RECT 33.140 172.405 33.805 172.575 ;
        RECT 33.140 172.150 33.310 172.405 ;
        RECT 34.065 172.355 35.735 173.125 ;
        RECT 35.995 172.575 36.165 172.955 ;
        RECT 36.345 172.745 36.675 173.125 ;
        RECT 35.995 172.405 36.660 172.575 ;
        RECT 36.855 172.450 37.115 172.955 ;
        RECT 33.025 171.820 33.310 172.150 ;
        RECT 33.545 171.855 33.875 172.225 ;
        RECT 33.140 171.675 33.310 171.820 ;
        RECT 31.760 171.245 32.510 171.415 ;
        RECT 31.755 170.575 32.085 171.075 ;
        RECT 32.255 170.745 32.510 171.245 ;
        RECT 32.685 170.745 32.955 171.650 ;
        RECT 33.140 171.505 33.805 171.675 ;
        RECT 33.125 170.575 33.455 171.335 ;
        RECT 33.635 170.745 33.805 171.505 ;
        RECT 34.065 171.665 34.815 172.185 ;
        RECT 34.985 171.835 35.735 172.355 ;
        RECT 35.925 171.855 36.255 172.225 ;
        RECT 36.490 172.150 36.660 172.405 ;
        RECT 36.490 171.820 36.775 172.150 ;
        RECT 36.490 171.675 36.660 171.820 ;
        RECT 34.065 170.575 35.735 171.665 ;
        RECT 35.995 171.505 36.660 171.675 ;
        RECT 36.945 171.650 37.115 172.450 ;
        RECT 37.285 172.400 37.575 173.125 ;
        RECT 37.750 172.385 38.005 172.955 ;
        RECT 38.175 172.725 38.505 173.125 ;
        RECT 38.930 172.590 39.460 172.955 ;
        RECT 38.930 172.555 39.105 172.590 ;
        RECT 38.175 172.385 39.105 172.555 ;
        RECT 35.995 170.745 36.165 171.505 ;
        RECT 36.345 170.575 36.675 171.335 ;
        RECT 36.845 170.745 37.115 171.650 ;
        RECT 37.285 170.575 37.575 171.740 ;
        RECT 37.750 171.715 37.920 172.385 ;
        RECT 38.175 172.215 38.345 172.385 ;
        RECT 38.090 171.885 38.345 172.215 ;
        RECT 38.570 171.885 38.765 172.215 ;
        RECT 37.750 170.745 38.085 171.715 ;
        RECT 38.255 170.575 38.425 171.715 ;
        RECT 38.595 170.915 38.765 171.885 ;
        RECT 38.935 171.255 39.105 172.385 ;
        RECT 39.275 171.595 39.445 172.395 ;
        RECT 39.650 172.105 39.925 172.955 ;
        RECT 39.645 171.935 39.925 172.105 ;
        RECT 39.650 171.795 39.925 171.935 ;
        RECT 40.095 171.595 40.285 172.955 ;
        RECT 40.465 172.590 40.975 173.125 ;
        RECT 41.195 172.315 41.440 172.920 ;
        RECT 41.975 172.645 42.275 173.125 ;
        RECT 42.445 172.475 42.705 172.930 ;
        RECT 42.875 172.645 43.135 173.125 ;
        RECT 43.315 172.475 43.575 172.930 ;
        RECT 43.745 172.645 43.995 173.125 ;
        RECT 44.175 172.475 44.435 172.930 ;
        RECT 44.605 172.645 44.855 173.125 ;
        RECT 45.035 172.475 45.295 172.930 ;
        RECT 45.465 172.645 45.710 173.125 ;
        RECT 45.880 172.475 46.155 172.930 ;
        RECT 46.325 172.645 46.570 173.125 ;
        RECT 46.740 172.475 47.000 172.930 ;
        RECT 47.170 172.645 47.430 173.125 ;
        RECT 47.600 172.475 47.860 172.930 ;
        RECT 48.030 172.645 48.290 173.125 ;
        RECT 48.460 172.475 48.720 172.930 ;
        RECT 48.890 172.565 49.150 173.125 ;
        RECT 40.485 172.145 41.715 172.315 ;
        RECT 39.275 171.425 40.285 171.595 ;
        RECT 40.455 171.580 41.205 171.770 ;
        RECT 38.935 171.085 40.060 171.255 ;
        RECT 40.455 170.915 40.625 171.580 ;
        RECT 41.375 171.335 41.715 172.145 ;
        RECT 41.975 172.305 48.720 172.475 ;
        RECT 41.975 171.715 43.140 172.305 ;
        RECT 49.320 172.135 49.570 172.945 ;
        RECT 49.750 172.600 50.010 173.125 ;
        RECT 50.180 172.135 50.430 172.945 ;
        RECT 50.610 172.615 50.915 173.125 ;
        RECT 43.310 171.885 50.430 172.135 ;
        RECT 50.600 171.885 50.915 172.445 ;
        RECT 51.755 172.435 52.085 173.125 ;
        RECT 52.545 172.530 53.165 172.955 ;
        RECT 53.335 172.635 53.665 173.125 ;
        RECT 52.805 172.195 53.165 172.530 ;
        RECT 51.745 171.915 53.165 172.195 ;
        RECT 41.975 171.490 48.720 171.715 ;
        RECT 38.595 170.745 40.625 170.915 ;
        RECT 40.795 170.575 40.965 171.335 ;
        RECT 41.200 170.925 41.715 171.335 ;
        RECT 41.975 170.575 42.245 171.320 ;
        RECT 42.415 170.750 42.705 171.490 ;
        RECT 43.315 171.475 48.720 171.490 ;
        RECT 42.875 170.580 43.130 171.305 ;
        RECT 43.315 170.750 43.575 171.475 ;
        RECT 43.745 170.580 43.990 171.305 ;
        RECT 44.175 170.750 44.435 171.475 ;
        RECT 44.605 170.580 44.850 171.305 ;
        RECT 45.035 170.750 45.295 171.475 ;
        RECT 45.465 170.580 45.710 171.305 ;
        RECT 45.880 170.750 46.140 171.475 ;
        RECT 46.310 170.580 46.570 171.305 ;
        RECT 46.740 170.750 47.000 171.475 ;
        RECT 47.170 170.580 47.430 171.305 ;
        RECT 47.600 170.750 47.860 171.475 ;
        RECT 48.030 170.580 48.290 171.305 ;
        RECT 48.460 170.750 48.720 171.475 ;
        RECT 48.890 170.580 49.150 171.375 ;
        RECT 49.320 170.750 49.570 171.885 ;
        RECT 42.875 170.575 49.150 170.580 ;
        RECT 49.750 170.575 50.010 171.385 ;
        RECT 50.185 170.745 50.430 171.885 ;
        RECT 50.610 170.575 50.905 171.385 ;
        RECT 51.215 170.575 51.545 171.745 ;
        RECT 51.745 170.745 52.075 171.915 ;
        RECT 52.275 170.575 52.605 171.745 ;
        RECT 52.805 170.745 53.165 171.915 ;
        RECT 53.335 171.885 53.675 172.465 ;
        RECT 54.305 172.355 56.895 173.125 ;
        RECT 57.125 172.645 57.405 173.125 ;
        RECT 57.575 172.475 57.835 172.865 ;
        RECT 58.010 172.645 58.265 173.125 ;
        RECT 58.435 172.475 58.730 172.865 ;
        RECT 58.910 172.645 59.185 173.125 ;
        RECT 59.355 172.625 59.655 172.955 ;
        RECT 53.335 170.575 53.665 171.715 ;
        RECT 54.305 171.665 55.515 172.185 ;
        RECT 55.685 171.835 56.895 172.355 ;
        RECT 57.080 172.305 58.730 172.475 ;
        RECT 57.080 171.795 57.485 172.305 ;
        RECT 57.655 171.965 58.795 172.135 ;
        RECT 54.305 170.575 56.895 171.665 ;
        RECT 57.080 171.625 57.835 171.795 ;
        RECT 57.120 170.575 57.405 171.445 ;
        RECT 57.575 171.375 57.835 171.625 ;
        RECT 58.625 171.715 58.795 171.965 ;
        RECT 58.965 171.885 59.315 172.455 ;
        RECT 59.485 171.715 59.655 172.625 ;
        RECT 60.285 172.355 62.875 173.125 ;
        RECT 63.045 172.400 63.335 173.125 ;
        RECT 58.625 171.545 59.655 171.715 ;
        RECT 57.575 171.205 58.695 171.375 ;
        RECT 57.575 170.745 57.835 171.205 ;
        RECT 58.010 170.575 58.265 171.035 ;
        RECT 58.435 170.745 58.695 171.205 ;
        RECT 58.865 170.575 59.175 171.375 ;
        RECT 59.345 170.745 59.655 171.545 ;
        RECT 60.285 171.665 61.495 172.185 ;
        RECT 61.665 171.835 62.875 172.355 ;
        RECT 64.430 172.285 64.690 173.125 ;
        RECT 64.865 172.380 65.120 172.955 ;
        RECT 65.290 172.745 65.620 173.125 ;
        RECT 65.835 172.575 66.005 172.955 ;
        RECT 65.290 172.405 66.005 172.575 ;
        RECT 66.355 172.575 66.525 172.955 ;
        RECT 66.740 172.745 67.070 173.125 ;
        RECT 66.355 172.405 67.070 172.575 ;
        RECT 60.285 170.575 62.875 171.665 ;
        RECT 63.045 170.575 63.335 171.740 ;
        RECT 64.430 170.575 64.690 171.725 ;
        RECT 64.865 171.650 65.035 172.380 ;
        RECT 65.290 172.215 65.460 172.405 ;
        RECT 65.205 171.885 65.460 172.215 ;
        RECT 65.290 171.675 65.460 171.885 ;
        RECT 65.740 171.855 66.095 172.225 ;
        RECT 66.265 171.855 66.620 172.225 ;
        RECT 66.900 172.215 67.070 172.405 ;
        RECT 67.240 172.380 67.495 172.955 ;
        RECT 66.900 171.885 67.155 172.215 ;
        RECT 66.900 171.675 67.070 171.885 ;
        RECT 64.865 170.745 65.120 171.650 ;
        RECT 65.290 171.505 66.005 171.675 ;
        RECT 65.290 170.575 65.620 171.335 ;
        RECT 65.835 170.745 66.005 171.505 ;
        RECT 66.355 171.505 67.070 171.675 ;
        RECT 67.325 171.650 67.495 172.380 ;
        RECT 67.670 172.285 67.930 173.125 ;
        RECT 68.565 172.355 70.235 173.125 ;
        RECT 66.355 170.745 66.525 171.505 ;
        RECT 66.740 170.575 67.070 171.335 ;
        RECT 67.240 170.745 67.495 171.650 ;
        RECT 67.670 170.575 67.930 171.725 ;
        RECT 68.565 171.665 69.315 172.185 ;
        RECT 69.485 171.835 70.235 172.355 ;
        RECT 70.445 172.305 70.675 173.125 ;
        RECT 70.845 172.325 71.175 172.955 ;
        RECT 70.425 171.885 70.755 172.135 ;
        RECT 70.925 171.725 71.175 172.325 ;
        RECT 71.345 172.305 71.555 173.125 ;
        RECT 72.055 172.730 72.385 173.125 ;
        RECT 72.555 172.555 72.755 172.910 ;
        RECT 72.925 172.725 73.255 173.125 ;
        RECT 73.425 172.555 73.625 172.900 ;
        RECT 71.785 172.385 73.625 172.555 ;
        RECT 73.795 172.385 74.125 173.125 ;
        RECT 74.360 172.555 74.530 172.805 ;
        RECT 74.360 172.385 74.835 172.555 ;
        RECT 68.565 170.575 70.235 171.665 ;
        RECT 70.445 170.575 70.675 171.715 ;
        RECT 70.845 170.745 71.175 171.725 ;
        RECT 71.345 170.575 71.555 171.715 ;
        RECT 71.785 170.760 72.045 172.385 ;
        RECT 72.225 171.415 72.445 172.215 ;
        RECT 72.685 171.595 72.985 172.215 ;
        RECT 73.155 171.595 73.485 172.215 ;
        RECT 73.655 171.595 73.975 172.215 ;
        RECT 74.145 171.595 74.495 172.215 ;
        RECT 74.665 171.415 74.835 172.385 ;
        RECT 75.005 172.375 76.215 173.125 ;
        RECT 72.225 171.205 74.835 171.415 ;
        RECT 75.005 171.665 75.525 172.205 ;
        RECT 75.695 171.835 76.215 172.375 ;
        RECT 76.385 172.625 76.685 172.955 ;
        RECT 76.855 172.645 77.130 173.125 ;
        RECT 76.385 171.715 76.555 172.625 ;
        RECT 77.310 172.475 77.605 172.865 ;
        RECT 77.775 172.645 78.030 173.125 ;
        RECT 78.205 172.475 78.465 172.865 ;
        RECT 78.635 172.645 78.915 173.125 ;
        RECT 76.725 171.885 77.075 172.455 ;
        RECT 77.310 172.305 78.960 172.475 ;
        RECT 77.245 171.965 78.385 172.135 ;
        RECT 77.245 171.715 77.415 171.965 ;
        RECT 78.555 171.795 78.960 172.305 ;
        RECT 73.795 170.575 74.125 171.025 ;
        RECT 75.005 170.575 76.215 171.665 ;
        RECT 76.385 171.545 77.415 171.715 ;
        RECT 78.205 171.625 78.960 171.795 ;
        RECT 79.520 172.415 79.775 172.945 ;
        RECT 79.955 172.665 80.240 173.125 ;
        RECT 76.385 170.745 76.695 171.545 ;
        RECT 78.205 171.375 78.465 171.625 ;
        RECT 79.520 171.555 79.700 172.415 ;
        RECT 80.420 172.215 80.670 172.865 ;
        RECT 79.870 171.885 80.670 172.215 ;
        RECT 76.865 170.575 77.175 171.375 ;
        RECT 77.345 171.205 78.465 171.375 ;
        RECT 77.345 170.745 77.605 171.205 ;
        RECT 77.775 170.575 78.030 171.035 ;
        RECT 78.205 170.745 78.465 171.205 ;
        RECT 78.635 170.575 78.920 171.445 ;
        RECT 79.520 171.085 79.775 171.555 ;
        RECT 79.435 170.915 79.775 171.085 ;
        RECT 79.520 170.885 79.775 170.915 ;
        RECT 79.955 170.575 80.240 171.375 ;
        RECT 80.420 171.295 80.670 171.885 ;
        RECT 80.870 172.530 81.190 172.860 ;
        RECT 81.370 172.645 82.030 173.125 ;
        RECT 82.230 172.735 83.080 172.905 ;
        RECT 80.870 171.635 81.060 172.530 ;
        RECT 81.380 172.205 82.040 172.475 ;
        RECT 81.710 172.145 82.040 172.205 ;
        RECT 81.230 171.975 81.560 172.035 ;
        RECT 82.230 171.975 82.400 172.735 ;
        RECT 83.640 172.665 83.960 173.125 ;
        RECT 84.160 172.485 84.410 172.915 ;
        RECT 84.700 172.685 85.110 173.125 ;
        RECT 85.280 172.745 86.295 172.945 ;
        RECT 82.570 172.315 83.820 172.485 ;
        RECT 82.570 172.195 82.900 172.315 ;
        RECT 81.230 171.805 83.130 171.975 ;
        RECT 80.870 171.465 82.790 171.635 ;
        RECT 80.870 171.445 81.190 171.465 ;
        RECT 80.420 170.785 80.750 171.295 ;
        RECT 81.020 170.835 81.190 171.445 ;
        RECT 82.960 171.295 83.130 171.805 ;
        RECT 83.300 171.735 83.480 172.145 ;
        RECT 83.650 171.555 83.820 172.315 ;
        RECT 81.360 170.575 81.690 171.265 ;
        RECT 81.920 171.125 83.130 171.295 ;
        RECT 83.300 171.245 83.820 171.555 ;
        RECT 83.990 172.145 84.410 172.485 ;
        RECT 84.700 172.145 85.110 172.475 ;
        RECT 83.990 171.375 84.180 172.145 ;
        RECT 85.280 172.015 85.450 172.745 ;
        RECT 86.595 172.575 86.765 172.905 ;
        RECT 86.935 172.745 87.265 173.125 ;
        RECT 85.620 172.195 85.970 172.565 ;
        RECT 85.280 171.975 85.700 172.015 ;
        RECT 84.350 171.805 85.700 171.975 ;
        RECT 84.350 171.645 84.600 171.805 ;
        RECT 85.110 171.375 85.360 171.635 ;
        RECT 83.990 171.125 85.360 171.375 ;
        RECT 81.920 170.835 82.160 171.125 ;
        RECT 82.960 171.045 83.130 171.125 ;
        RECT 82.360 170.575 82.780 170.955 ;
        RECT 82.960 170.795 83.590 171.045 ;
        RECT 84.060 170.575 84.390 170.955 ;
        RECT 84.560 170.835 84.730 171.125 ;
        RECT 85.530 170.960 85.700 171.805 ;
        RECT 86.150 171.635 86.370 172.505 ;
        RECT 86.595 172.385 87.290 172.575 ;
        RECT 85.870 171.255 86.370 171.635 ;
        RECT 86.540 171.585 86.950 172.205 ;
        RECT 87.120 171.415 87.290 172.385 ;
        RECT 86.595 171.245 87.290 171.415 ;
        RECT 84.910 170.575 85.290 170.955 ;
        RECT 85.530 170.790 86.360 170.960 ;
        RECT 86.595 170.745 86.765 171.245 ;
        RECT 86.935 170.575 87.265 171.075 ;
        RECT 87.480 170.745 87.705 172.865 ;
        RECT 87.875 172.745 88.205 173.125 ;
        RECT 88.375 172.575 88.545 172.865 ;
        RECT 87.880 172.405 88.545 172.575 ;
        RECT 87.880 171.415 88.110 172.405 ;
        RECT 88.805 172.400 89.095 173.125 ;
        RECT 89.725 172.355 91.395 173.125 ;
        RECT 91.570 172.580 96.915 173.125 ;
        RECT 88.280 171.585 88.630 172.235 ;
        RECT 87.880 171.245 88.545 171.415 ;
        RECT 87.875 170.575 88.205 171.075 ;
        RECT 88.375 170.745 88.545 171.245 ;
        RECT 88.805 170.575 89.095 171.740 ;
        RECT 89.725 171.665 90.475 172.185 ;
        RECT 90.645 171.835 91.395 172.355 ;
        RECT 89.725 170.575 91.395 171.665 ;
        RECT 93.160 171.010 93.510 172.260 ;
        RECT 94.990 171.750 95.330 172.580 ;
        RECT 97.360 172.315 97.605 172.920 ;
        RECT 97.825 172.590 98.335 173.125 ;
        RECT 97.085 172.145 98.315 172.315 ;
        RECT 97.085 171.335 97.425 172.145 ;
        RECT 97.595 171.580 98.345 171.770 ;
        RECT 91.570 170.575 96.915 171.010 ;
        RECT 97.085 170.925 97.600 171.335 ;
        RECT 97.835 170.575 98.005 171.335 ;
        RECT 98.175 170.915 98.345 171.580 ;
        RECT 98.515 171.595 98.705 172.955 ;
        RECT 98.875 172.105 99.150 172.955 ;
        RECT 99.340 172.590 99.870 172.955 ;
        RECT 100.295 172.725 100.625 173.125 ;
        RECT 99.695 172.555 99.870 172.590 ;
        RECT 98.875 171.935 99.155 172.105 ;
        RECT 98.875 171.795 99.150 171.935 ;
        RECT 99.355 171.595 99.525 172.395 ;
        RECT 98.515 171.425 99.525 171.595 ;
        RECT 99.695 172.385 100.625 172.555 ;
        RECT 100.795 172.385 101.050 172.955 ;
        RECT 99.695 171.255 99.865 172.385 ;
        RECT 100.455 172.215 100.625 172.385 ;
        RECT 98.740 171.085 99.865 171.255 ;
        RECT 100.035 171.885 100.230 172.215 ;
        RECT 100.455 171.885 100.710 172.215 ;
        RECT 100.035 170.915 100.205 171.885 ;
        RECT 100.880 171.715 101.050 172.385 ;
        RECT 98.175 170.745 100.205 170.915 ;
        RECT 100.375 170.575 100.545 171.715 ;
        RECT 100.715 170.745 101.050 171.715 ;
        RECT 102.145 172.450 102.405 172.955 ;
        RECT 102.585 172.745 102.915 173.125 ;
        RECT 103.095 172.575 103.265 172.955 ;
        RECT 103.530 172.580 108.875 173.125 ;
        RECT 102.145 171.650 102.315 172.450 ;
        RECT 102.600 172.405 103.265 172.575 ;
        RECT 102.600 172.150 102.770 172.405 ;
        RECT 102.485 171.820 102.770 172.150 ;
        RECT 103.005 171.855 103.335 172.225 ;
        RECT 102.600 171.675 102.770 171.820 ;
        RECT 102.145 170.745 102.415 171.650 ;
        RECT 102.600 171.505 103.265 171.675 ;
        RECT 102.585 170.575 102.915 171.335 ;
        RECT 103.095 170.745 103.265 171.505 ;
        RECT 105.120 171.010 105.470 172.260 ;
        RECT 106.950 171.750 107.290 172.580 ;
        RECT 109.045 172.325 109.385 172.955 ;
        RECT 109.555 172.325 109.805 173.125 ;
        RECT 109.995 172.475 110.325 172.955 ;
        RECT 110.495 172.665 110.720 173.125 ;
        RECT 110.890 172.475 111.220 172.955 ;
        RECT 109.045 171.715 109.220 172.325 ;
        RECT 109.995 172.305 111.220 172.475 ;
        RECT 111.850 172.345 112.350 172.955 ;
        RECT 112.725 172.355 114.395 173.125 ;
        RECT 114.565 172.400 114.855 173.125 ;
        RECT 115.575 172.575 115.745 172.955 ;
        RECT 115.925 172.745 116.255 173.125 ;
        RECT 115.575 172.405 116.240 172.575 ;
        RECT 116.435 172.450 116.695 172.955 ;
        RECT 109.390 171.965 110.085 172.135 ;
        RECT 109.915 171.715 110.085 171.965 ;
        RECT 110.260 171.935 110.680 172.135 ;
        RECT 110.850 171.935 111.180 172.135 ;
        RECT 111.350 171.935 111.680 172.135 ;
        RECT 111.850 171.715 112.020 172.345 ;
        RECT 112.205 171.885 112.555 172.135 ;
        RECT 103.530 170.575 108.875 171.010 ;
        RECT 109.045 170.745 109.385 171.715 ;
        RECT 109.555 170.575 109.725 171.715 ;
        RECT 109.915 171.545 112.350 171.715 ;
        RECT 109.995 170.575 110.245 171.375 ;
        RECT 110.890 170.745 111.220 171.545 ;
        RECT 111.520 170.575 111.850 171.375 ;
        RECT 112.020 170.745 112.350 171.545 ;
        RECT 112.725 171.665 113.475 172.185 ;
        RECT 113.645 171.835 114.395 172.355 ;
        RECT 115.505 171.855 115.835 172.225 ;
        RECT 116.070 172.150 116.240 172.405 ;
        RECT 116.070 171.820 116.355 172.150 ;
        RECT 112.725 170.575 114.395 171.665 ;
        RECT 114.565 170.575 114.855 171.740 ;
        RECT 116.070 171.675 116.240 171.820 ;
        RECT 115.575 171.505 116.240 171.675 ;
        RECT 116.525 171.650 116.695 172.450 ;
        RECT 115.575 170.745 115.745 171.505 ;
        RECT 115.925 170.575 116.255 171.335 ;
        RECT 116.425 170.745 116.695 171.650 ;
        RECT 116.870 172.415 117.125 172.945 ;
        RECT 117.295 172.665 117.600 173.125 ;
        RECT 117.845 172.745 118.915 172.915 ;
        RECT 116.870 171.765 117.080 172.415 ;
        RECT 117.845 172.390 118.165 172.745 ;
        RECT 117.840 172.215 118.165 172.390 ;
        RECT 117.250 171.915 118.165 172.215 ;
        RECT 118.335 172.175 118.575 172.575 ;
        RECT 118.745 172.515 118.915 172.745 ;
        RECT 119.085 172.685 119.275 173.125 ;
        RECT 119.445 172.675 120.395 172.955 ;
        RECT 120.615 172.765 120.965 172.935 ;
        RECT 118.745 172.345 119.275 172.515 ;
        RECT 117.250 171.885 117.990 171.915 ;
        RECT 116.870 170.885 117.125 171.765 ;
        RECT 117.295 170.575 117.600 171.715 ;
        RECT 117.820 171.295 117.990 171.885 ;
        RECT 118.335 171.805 118.875 172.175 ;
        RECT 119.055 172.065 119.275 172.345 ;
        RECT 119.445 171.895 119.615 172.675 ;
        RECT 119.210 171.725 119.615 171.895 ;
        RECT 119.785 171.885 120.135 172.505 ;
        RECT 119.210 171.635 119.380 171.725 ;
        RECT 120.305 171.715 120.515 172.505 ;
        RECT 118.160 171.465 119.380 171.635 ;
        RECT 119.840 171.555 120.515 171.715 ;
        RECT 117.820 171.125 118.620 171.295 ;
        RECT 117.940 170.575 118.270 170.955 ;
        RECT 118.450 170.835 118.620 171.125 ;
        RECT 119.210 171.085 119.380 171.465 ;
        RECT 119.550 171.545 120.515 171.555 ;
        RECT 120.705 172.375 120.965 172.765 ;
        RECT 121.175 172.665 121.505 173.125 ;
        RECT 122.380 172.735 123.235 172.905 ;
        RECT 123.440 172.735 123.935 172.905 ;
        RECT 124.105 172.765 124.435 173.125 ;
        RECT 120.705 171.685 120.875 172.375 ;
        RECT 121.045 172.025 121.215 172.205 ;
        RECT 121.385 172.195 122.175 172.445 ;
        RECT 122.380 172.025 122.550 172.735 ;
        RECT 122.720 172.225 123.075 172.445 ;
        RECT 121.045 171.855 122.735 172.025 ;
        RECT 119.550 171.255 120.010 171.545 ;
        RECT 120.705 171.515 122.205 171.685 ;
        RECT 120.705 171.375 120.875 171.515 ;
        RECT 120.315 171.205 120.875 171.375 ;
        RECT 118.790 170.575 119.040 171.035 ;
        RECT 119.210 170.745 120.080 171.085 ;
        RECT 120.315 170.745 120.485 171.205 ;
        RECT 121.320 171.175 122.395 171.345 ;
        RECT 120.655 170.575 121.025 171.035 ;
        RECT 121.320 170.835 121.490 171.175 ;
        RECT 121.660 170.575 121.990 171.005 ;
        RECT 122.225 170.835 122.395 171.175 ;
        RECT 122.565 171.075 122.735 171.855 ;
        RECT 122.905 171.635 123.075 172.225 ;
        RECT 123.245 171.825 123.595 172.445 ;
        RECT 122.905 171.245 123.370 171.635 ;
        RECT 123.765 171.375 123.935 172.735 ;
        RECT 124.105 171.545 124.565 172.595 ;
        RECT 123.540 171.205 123.935 171.375 ;
        RECT 123.540 171.075 123.710 171.205 ;
        RECT 122.565 170.745 123.245 171.075 ;
        RECT 123.460 170.745 123.710 171.075 ;
        RECT 123.880 170.575 124.130 171.035 ;
        RECT 124.300 170.760 124.625 171.545 ;
        RECT 124.795 170.745 124.965 172.865 ;
        RECT 125.135 172.745 125.465 173.125 ;
        RECT 125.635 172.575 125.890 172.865 ;
        RECT 125.140 172.405 125.890 172.575 ;
        RECT 125.140 171.415 125.370 172.405 ;
        RECT 126.525 172.375 127.735 173.125 ;
        RECT 125.540 171.585 125.890 172.235 ;
        RECT 126.525 171.665 127.045 172.205 ;
        RECT 127.215 171.835 127.735 172.375 ;
        RECT 125.140 171.245 125.890 171.415 ;
        RECT 125.135 170.575 125.465 171.075 ;
        RECT 125.635 170.745 125.890 171.245 ;
        RECT 126.525 170.575 127.735 171.665 ;
        RECT 14.660 170.405 127.820 170.575 ;
        RECT 14.745 169.315 15.955 170.405 ;
        RECT 16.130 169.970 21.475 170.405 ;
        RECT 14.745 168.605 15.265 169.145 ;
        RECT 15.435 168.775 15.955 169.315 ;
        RECT 17.720 168.720 18.070 169.970 ;
        RECT 21.705 169.265 21.915 170.405 ;
        RECT 22.085 169.255 22.415 170.235 ;
        RECT 22.585 169.265 22.815 170.405 ;
        RECT 23.025 169.315 24.235 170.405 ;
        RECT 14.745 167.855 15.955 168.605 ;
        RECT 19.550 168.400 19.890 169.230 ;
        RECT 16.130 167.855 21.475 168.400 ;
        RECT 21.705 167.855 21.915 168.675 ;
        RECT 22.085 168.655 22.335 169.255 ;
        RECT 22.505 168.845 22.835 169.095 ;
        RECT 23.025 168.775 23.545 169.315 ;
        RECT 24.405 169.240 24.695 170.405 ;
        RECT 25.325 169.315 27.915 170.405 ;
        RECT 28.090 169.970 33.435 170.405 ;
        RECT 33.610 169.970 38.955 170.405 ;
        RECT 22.085 168.025 22.415 168.655 ;
        RECT 22.585 167.855 22.815 168.675 ;
        RECT 23.715 168.605 24.235 169.145 ;
        RECT 25.325 168.795 26.535 169.315 ;
        RECT 26.705 168.625 27.915 169.145 ;
        RECT 29.680 168.720 30.030 169.970 ;
        RECT 23.025 167.855 24.235 168.605 ;
        RECT 24.405 167.855 24.695 168.580 ;
        RECT 25.325 167.855 27.915 168.625 ;
        RECT 31.510 168.400 31.850 169.230 ;
        RECT 35.200 168.720 35.550 169.970 ;
        RECT 39.275 169.255 39.605 170.405 ;
        RECT 39.775 169.385 39.945 170.235 ;
        RECT 40.115 169.605 40.445 170.405 ;
        RECT 40.615 169.385 40.785 170.235 ;
        RECT 40.965 169.605 41.205 170.405 ;
        RECT 41.375 169.425 41.705 170.235 ;
        RECT 37.030 168.400 37.370 169.230 ;
        RECT 39.775 169.215 40.785 169.385 ;
        RECT 40.990 169.255 41.705 169.425 ;
        RECT 43.010 169.435 43.340 170.235 ;
        RECT 43.510 169.605 43.840 170.405 ;
        RECT 44.140 169.435 44.470 170.235 ;
        RECT 45.115 169.605 45.365 170.405 ;
        RECT 43.010 169.265 45.445 169.435 ;
        RECT 45.635 169.265 45.805 170.405 ;
        RECT 45.975 169.265 46.315 170.235 ;
        RECT 39.775 168.675 40.270 169.215 ;
        RECT 40.990 169.015 41.160 169.255 ;
        RECT 40.660 168.845 41.160 169.015 ;
        RECT 41.330 168.845 41.710 169.085 ;
        RECT 42.805 168.845 43.155 169.095 ;
        RECT 40.990 168.675 41.160 168.845 ;
        RECT 28.090 167.855 33.435 168.400 ;
        RECT 33.610 167.855 38.955 168.400 ;
        RECT 39.275 167.855 39.605 168.655 ;
        RECT 39.775 168.505 40.785 168.675 ;
        RECT 40.990 168.505 41.625 168.675 ;
        RECT 43.340 168.635 43.510 169.265 ;
        RECT 43.680 168.845 44.010 169.045 ;
        RECT 44.180 168.845 44.510 169.045 ;
        RECT 44.680 168.845 45.100 169.045 ;
        RECT 45.275 169.015 45.445 169.265 ;
        RECT 45.275 168.845 45.970 169.015 ;
        RECT 39.775 168.025 39.945 168.505 ;
        RECT 40.115 167.855 40.445 168.335 ;
        RECT 40.615 168.025 40.785 168.505 ;
        RECT 41.035 167.855 41.275 168.335 ;
        RECT 41.455 168.025 41.625 168.505 ;
        RECT 43.010 168.025 43.510 168.635 ;
        RECT 44.140 168.505 45.365 168.675 ;
        RECT 46.140 168.655 46.315 169.265 ;
        RECT 44.140 168.025 44.470 168.505 ;
        RECT 44.640 167.855 44.865 168.315 ;
        RECT 45.035 168.025 45.365 168.505 ;
        RECT 45.555 167.855 45.805 168.655 ;
        RECT 45.975 168.025 46.315 168.655 ;
        RECT 46.485 169.265 46.825 170.235 ;
        RECT 46.995 169.265 47.165 170.405 ;
        RECT 47.435 169.605 47.685 170.405 ;
        RECT 48.330 169.435 48.660 170.235 ;
        RECT 48.960 169.605 49.290 170.405 ;
        RECT 49.460 169.435 49.790 170.235 ;
        RECT 47.355 169.265 49.790 169.435 ;
        RECT 46.485 168.655 46.660 169.265 ;
        RECT 47.355 169.015 47.525 169.265 ;
        RECT 46.830 168.845 47.525 169.015 ;
        RECT 47.700 168.845 48.120 169.045 ;
        RECT 48.290 168.845 48.620 169.045 ;
        RECT 48.790 168.845 49.120 169.045 ;
        RECT 46.485 168.025 46.825 168.655 ;
        RECT 46.995 167.855 47.245 168.655 ;
        RECT 47.435 168.505 48.660 168.675 ;
        RECT 47.435 168.025 47.765 168.505 ;
        RECT 47.935 167.855 48.160 168.315 ;
        RECT 48.330 168.025 48.660 168.505 ;
        RECT 49.290 168.635 49.460 169.265 ;
        RECT 50.165 169.240 50.455 170.405 ;
        RECT 50.625 169.315 51.835 170.405 ;
        RECT 49.645 168.845 49.995 169.095 ;
        RECT 50.625 168.775 51.145 169.315 ;
        RECT 52.005 169.265 52.345 170.235 ;
        RECT 52.515 169.265 52.685 170.405 ;
        RECT 52.955 169.605 53.205 170.405 ;
        RECT 53.850 169.435 54.180 170.235 ;
        RECT 54.480 169.605 54.810 170.405 ;
        RECT 54.980 169.435 55.310 170.235 ;
        RECT 56.150 169.970 61.495 170.405 ;
        RECT 52.875 169.265 55.310 169.435 ;
        RECT 49.290 168.025 49.790 168.635 ;
        RECT 51.315 168.605 51.835 169.145 ;
        RECT 50.165 167.855 50.455 168.580 ;
        RECT 50.625 167.855 51.835 168.605 ;
        RECT 52.005 168.655 52.180 169.265 ;
        RECT 52.875 169.015 53.045 169.265 ;
        RECT 52.350 168.845 53.045 169.015 ;
        RECT 53.220 168.845 53.640 169.045 ;
        RECT 53.810 168.845 54.140 169.045 ;
        RECT 54.310 168.845 54.640 169.045 ;
        RECT 52.005 168.025 52.345 168.655 ;
        RECT 52.515 167.855 52.765 168.655 ;
        RECT 52.955 168.505 54.180 168.675 ;
        RECT 52.955 168.025 53.285 168.505 ;
        RECT 53.455 167.855 53.680 168.315 ;
        RECT 53.850 168.025 54.180 168.505 ;
        RECT 54.810 168.635 54.980 169.265 ;
        RECT 55.165 168.845 55.515 169.095 ;
        RECT 57.740 168.720 58.090 169.970 ;
        RECT 61.720 169.535 62.005 170.405 ;
        RECT 62.175 169.775 62.435 170.235 ;
        RECT 62.610 169.945 62.865 170.405 ;
        RECT 63.035 169.775 63.295 170.235 ;
        RECT 62.175 169.605 63.295 169.775 ;
        RECT 63.465 169.605 63.775 170.405 ;
        RECT 62.175 169.355 62.435 169.605 ;
        RECT 63.945 169.435 64.255 170.235 ;
        RECT 54.810 168.025 55.310 168.635 ;
        RECT 59.570 168.400 59.910 169.230 ;
        RECT 61.680 169.185 62.435 169.355 ;
        RECT 63.225 169.265 64.255 169.435 ;
        RECT 61.680 168.675 62.085 169.185 ;
        RECT 63.225 169.015 63.395 169.265 ;
        RECT 62.255 168.845 63.395 169.015 ;
        RECT 61.680 168.505 63.330 168.675 ;
        RECT 63.565 168.525 63.915 169.095 ;
        RECT 56.150 167.855 61.495 168.400 ;
        RECT 61.725 167.855 62.005 168.335 ;
        RECT 62.175 168.115 62.435 168.505 ;
        RECT 62.610 167.855 62.865 168.335 ;
        RECT 63.035 168.115 63.330 168.505 ;
        RECT 64.085 168.355 64.255 169.265 ;
        RECT 64.425 169.315 65.635 170.405 ;
        RECT 65.895 169.475 66.065 170.235 ;
        RECT 66.280 169.645 66.610 170.405 ;
        RECT 64.425 168.775 64.945 169.315 ;
        RECT 65.895 169.305 66.610 169.475 ;
        RECT 66.780 169.330 67.035 170.235 ;
        RECT 65.115 168.605 65.635 169.145 ;
        RECT 65.805 168.755 66.160 169.125 ;
        RECT 66.440 169.095 66.610 169.305 ;
        RECT 66.440 168.765 66.695 169.095 ;
        RECT 63.510 167.855 63.785 168.335 ;
        RECT 63.955 168.025 64.255 168.355 ;
        RECT 64.425 167.855 65.635 168.605 ;
        RECT 66.440 168.575 66.610 168.765 ;
        RECT 66.865 168.600 67.035 169.330 ;
        RECT 67.210 169.255 67.470 170.405 ;
        RECT 68.575 169.345 68.905 170.405 ;
        RECT 69.085 169.095 69.255 170.020 ;
        RECT 69.425 169.815 69.755 170.215 ;
        RECT 69.925 170.045 70.255 170.405 ;
        RECT 70.455 169.815 71.155 170.235 ;
        RECT 69.425 169.585 71.155 169.815 ;
        RECT 69.425 169.365 69.755 169.585 ;
        RECT 69.950 169.095 70.275 169.385 ;
        RECT 68.565 168.765 68.875 169.095 ;
        RECT 69.085 168.765 69.460 169.095 ;
        RECT 69.780 168.765 70.275 169.095 ;
        RECT 70.450 168.845 70.780 169.385 ;
        RECT 65.895 168.405 66.610 168.575 ;
        RECT 65.895 168.025 66.065 168.405 ;
        RECT 66.280 167.855 66.610 168.235 ;
        RECT 66.780 168.025 67.035 168.600 ;
        RECT 67.210 167.855 67.470 168.695 ;
        RECT 70.950 168.615 71.155 169.585 ;
        RECT 71.395 169.465 71.655 170.235 ;
        RECT 71.825 169.635 72.155 170.405 ;
        RECT 72.325 170.065 73.445 170.235 ;
        RECT 72.325 169.465 72.515 170.065 ;
        RECT 71.395 169.295 72.515 169.465 ;
        RECT 72.685 169.480 73.015 169.895 ;
        RECT 73.185 169.870 73.445 170.065 ;
        RECT 73.675 169.685 74.005 170.405 ;
        RECT 74.175 169.480 74.365 170.235 ;
        RECT 74.535 169.685 74.865 170.405 ;
        RECT 75.035 169.480 75.295 170.235 ;
        RECT 75.465 169.945 75.725 170.405 ;
        RECT 72.685 169.310 75.295 169.480 ;
        RECT 68.575 168.385 69.935 168.595 ;
        RECT 68.575 168.025 68.905 168.385 ;
        RECT 69.075 167.855 69.405 168.215 ;
        RECT 69.605 168.025 69.935 168.385 ;
        RECT 70.445 168.025 71.155 168.615 ;
        RECT 71.385 169.015 72.280 169.065 ;
        RECT 71.385 168.845 72.335 169.015 ;
        RECT 72.505 168.845 73.475 169.125 ;
        RECT 73.935 168.845 74.795 169.135 ;
        RECT 71.385 168.535 71.725 168.845 ;
        RECT 71.895 168.405 74.435 168.615 ;
        RECT 71.895 168.285 72.085 168.405 ;
        RECT 74.605 168.235 74.795 168.660 ;
        RECT 74.965 168.440 75.295 169.310 ;
        RECT 75.465 168.765 75.755 169.740 ;
        RECT 75.925 169.240 76.215 170.405 ;
        RECT 76.385 169.315 78.055 170.405 ;
        RECT 78.230 169.970 83.575 170.405 ;
        RECT 76.385 168.795 77.135 169.315 ;
        RECT 77.305 168.625 78.055 169.145 ;
        RECT 79.820 168.720 80.170 169.970 ;
        RECT 83.745 169.645 84.260 170.055 ;
        RECT 84.495 169.645 84.665 170.405 ;
        RECT 84.835 170.065 86.865 170.235 ;
        RECT 73.675 168.215 74.795 168.235 ;
        RECT 71.395 167.855 71.725 168.215 ;
        RECT 72.255 167.855 72.585 168.215 ;
        RECT 73.115 167.855 73.445 168.215 ;
        RECT 73.675 168.025 75.745 168.215 ;
        RECT 75.925 167.855 76.215 168.580 ;
        RECT 76.385 167.855 78.055 168.625 ;
        RECT 81.650 168.400 81.990 169.230 ;
        RECT 83.745 168.835 84.085 169.645 ;
        RECT 84.835 169.400 85.005 170.065 ;
        RECT 85.400 169.725 86.525 169.895 ;
        RECT 84.255 169.210 85.005 169.400 ;
        RECT 85.175 169.385 86.185 169.555 ;
        RECT 83.745 168.665 84.975 168.835 ;
        RECT 78.230 167.855 83.575 168.400 ;
        RECT 84.020 168.060 84.265 168.665 ;
        RECT 84.485 167.855 84.995 168.390 ;
        RECT 85.175 168.025 85.365 169.385 ;
        RECT 85.535 168.365 85.810 169.185 ;
        RECT 86.015 168.585 86.185 169.385 ;
        RECT 86.355 168.595 86.525 169.725 ;
        RECT 86.695 169.095 86.865 170.065 ;
        RECT 87.035 169.265 87.205 170.405 ;
        RECT 87.375 169.265 87.710 170.235 ;
        RECT 87.945 169.265 88.155 170.405 ;
        RECT 86.695 168.765 86.890 169.095 ;
        RECT 87.115 168.765 87.370 169.095 ;
        RECT 87.115 168.595 87.285 168.765 ;
        RECT 87.540 168.595 87.710 169.265 ;
        RECT 88.325 169.255 88.655 170.235 ;
        RECT 88.825 169.265 89.055 170.405 ;
        RECT 89.265 169.330 89.535 170.235 ;
        RECT 89.705 169.645 90.035 170.405 ;
        RECT 90.215 169.475 90.385 170.235 ;
        RECT 86.355 168.425 87.285 168.595 ;
        RECT 86.355 168.390 86.530 168.425 ;
        RECT 85.535 168.195 85.815 168.365 ;
        RECT 85.535 168.025 85.810 168.195 ;
        RECT 86.000 168.025 86.530 168.390 ;
        RECT 86.955 167.855 87.285 168.255 ;
        RECT 87.455 168.025 87.710 168.595 ;
        RECT 87.945 167.855 88.155 168.675 ;
        RECT 88.325 168.655 88.575 169.255 ;
        RECT 88.745 168.845 89.075 169.095 ;
        RECT 88.325 168.025 88.655 168.655 ;
        RECT 88.825 167.855 89.055 168.675 ;
        RECT 89.265 168.530 89.435 169.330 ;
        RECT 89.720 169.305 90.385 169.475 ;
        RECT 90.645 169.315 91.855 170.405 ;
        RECT 92.030 169.970 97.375 170.405 ;
        RECT 89.720 169.160 89.890 169.305 ;
        RECT 89.605 168.830 89.890 169.160 ;
        RECT 89.720 168.575 89.890 168.830 ;
        RECT 90.125 168.755 90.455 169.125 ;
        RECT 90.645 168.775 91.165 169.315 ;
        RECT 91.335 168.605 91.855 169.145 ;
        RECT 93.620 168.720 93.970 169.970 ;
        RECT 97.545 169.645 98.060 170.055 ;
        RECT 98.295 169.645 98.465 170.405 ;
        RECT 98.635 170.065 100.665 170.235 ;
        RECT 89.265 168.025 89.525 168.530 ;
        RECT 89.720 168.405 90.385 168.575 ;
        RECT 89.705 167.855 90.035 168.235 ;
        RECT 90.215 168.025 90.385 168.405 ;
        RECT 90.645 167.855 91.855 168.605 ;
        RECT 95.450 168.400 95.790 169.230 ;
        RECT 97.545 168.835 97.885 169.645 ;
        RECT 98.635 169.400 98.805 170.065 ;
        RECT 99.200 169.725 100.325 169.895 ;
        RECT 98.055 169.210 98.805 169.400 ;
        RECT 98.975 169.385 99.985 169.555 ;
        RECT 97.545 168.665 98.775 168.835 ;
        RECT 92.030 167.855 97.375 168.400 ;
        RECT 97.820 168.060 98.065 168.665 ;
        RECT 98.285 167.855 98.795 168.390 ;
        RECT 98.975 168.025 99.165 169.385 ;
        RECT 99.335 168.365 99.610 169.185 ;
        RECT 99.815 168.585 99.985 169.385 ;
        RECT 100.155 168.595 100.325 169.725 ;
        RECT 100.495 169.095 100.665 170.065 ;
        RECT 100.835 169.265 101.005 170.405 ;
        RECT 101.175 169.265 101.510 170.235 ;
        RECT 100.495 168.765 100.690 169.095 ;
        RECT 100.915 168.765 101.170 169.095 ;
        RECT 100.915 168.595 101.085 168.765 ;
        RECT 101.340 168.595 101.510 169.265 ;
        RECT 101.685 169.240 101.975 170.405 ;
        RECT 103.155 169.475 103.325 170.235 ;
        RECT 103.505 169.645 103.835 170.405 ;
        RECT 103.155 169.305 103.820 169.475 ;
        RECT 104.005 169.330 104.275 170.235 ;
        RECT 103.650 169.160 103.820 169.305 ;
        RECT 103.085 168.755 103.415 169.125 ;
        RECT 103.650 168.830 103.935 169.160 ;
        RECT 100.155 168.425 101.085 168.595 ;
        RECT 100.155 168.390 100.330 168.425 ;
        RECT 99.335 168.195 99.615 168.365 ;
        RECT 99.335 168.025 99.610 168.195 ;
        RECT 99.800 168.025 100.330 168.390 ;
        RECT 100.755 167.855 101.085 168.255 ;
        RECT 101.255 168.025 101.510 168.595 ;
        RECT 101.685 167.855 101.975 168.580 ;
        RECT 103.650 168.575 103.820 168.830 ;
        RECT 103.155 168.405 103.820 168.575 ;
        RECT 104.105 168.530 104.275 169.330 ;
        RECT 103.155 168.025 103.325 168.405 ;
        RECT 103.505 167.855 103.835 168.235 ;
        RECT 104.015 168.025 104.275 168.530 ;
        RECT 104.905 169.265 105.245 170.235 ;
        RECT 105.415 169.265 105.585 170.405 ;
        RECT 105.855 169.605 106.105 170.405 ;
        RECT 106.750 169.435 107.080 170.235 ;
        RECT 107.380 169.605 107.710 170.405 ;
        RECT 107.880 169.435 108.210 170.235 ;
        RECT 105.775 169.265 108.210 169.435 ;
        RECT 108.585 169.315 110.255 170.405 ;
        RECT 110.425 169.645 110.940 170.055 ;
        RECT 111.175 169.645 111.345 170.405 ;
        RECT 111.515 170.065 113.545 170.235 ;
        RECT 104.905 168.655 105.080 169.265 ;
        RECT 105.775 169.015 105.945 169.265 ;
        RECT 105.250 168.845 105.945 169.015 ;
        RECT 106.120 168.845 106.540 169.045 ;
        RECT 106.710 168.845 107.040 169.045 ;
        RECT 107.210 168.845 107.540 169.045 ;
        RECT 104.905 168.025 105.245 168.655 ;
        RECT 105.415 167.855 105.665 168.655 ;
        RECT 105.855 168.505 107.080 168.675 ;
        RECT 105.855 168.025 106.185 168.505 ;
        RECT 106.355 167.855 106.580 168.315 ;
        RECT 106.750 168.025 107.080 168.505 ;
        RECT 107.710 168.635 107.880 169.265 ;
        RECT 108.065 168.845 108.415 169.095 ;
        RECT 108.585 168.795 109.335 169.315 ;
        RECT 107.710 168.025 108.210 168.635 ;
        RECT 109.505 168.625 110.255 169.145 ;
        RECT 110.425 168.835 110.765 169.645 ;
        RECT 111.515 169.400 111.685 170.065 ;
        RECT 112.080 169.725 113.205 169.895 ;
        RECT 110.935 169.210 111.685 169.400 ;
        RECT 111.855 169.385 112.865 169.555 ;
        RECT 110.425 168.665 111.655 168.835 ;
        RECT 108.585 167.855 110.255 168.625 ;
        RECT 110.700 168.060 110.945 168.665 ;
        RECT 111.165 167.855 111.675 168.390 ;
        RECT 111.855 168.025 112.045 169.385 ;
        RECT 112.215 168.365 112.490 169.185 ;
        RECT 112.695 168.585 112.865 169.385 ;
        RECT 113.035 168.595 113.205 169.725 ;
        RECT 113.375 169.095 113.545 170.065 ;
        RECT 113.715 169.265 113.885 170.405 ;
        RECT 114.055 169.265 114.390 170.235 ;
        RECT 113.375 168.765 113.570 169.095 ;
        RECT 113.795 168.765 114.050 169.095 ;
        RECT 113.795 168.595 113.965 168.765 ;
        RECT 114.220 168.595 114.390 169.265 ;
        RECT 114.940 169.425 115.195 170.095 ;
        RECT 115.375 169.605 115.660 170.405 ;
        RECT 115.840 169.685 116.170 170.195 ;
        RECT 114.940 168.705 115.120 169.425 ;
        RECT 115.840 169.095 116.090 169.685 ;
        RECT 116.440 169.535 116.610 170.145 ;
        RECT 116.780 169.715 117.110 170.405 ;
        RECT 117.340 169.855 117.580 170.145 ;
        RECT 117.780 170.025 118.200 170.405 ;
        RECT 118.380 169.935 119.010 170.185 ;
        RECT 119.480 170.025 119.810 170.405 ;
        RECT 118.380 169.855 118.550 169.935 ;
        RECT 119.980 169.855 120.150 170.145 ;
        RECT 120.330 170.025 120.710 170.405 ;
        RECT 120.950 170.020 121.780 170.190 ;
        RECT 117.340 169.685 118.550 169.855 ;
        RECT 115.290 168.765 116.090 169.095 ;
        RECT 113.035 168.425 113.965 168.595 ;
        RECT 113.035 168.390 113.210 168.425 ;
        RECT 112.215 168.195 112.495 168.365 ;
        RECT 112.215 168.025 112.490 168.195 ;
        RECT 112.680 168.025 113.210 168.390 ;
        RECT 113.635 167.855 113.965 168.255 ;
        RECT 114.135 168.025 114.390 168.595 ;
        RECT 114.855 168.565 115.120 168.705 ;
        RECT 114.855 168.535 115.195 168.565 ;
        RECT 114.940 168.035 115.195 168.535 ;
        RECT 115.375 167.855 115.660 168.315 ;
        RECT 115.840 168.115 116.090 168.765 ;
        RECT 116.290 169.515 116.610 169.535 ;
        RECT 116.290 169.345 118.210 169.515 ;
        RECT 116.290 168.450 116.480 169.345 ;
        RECT 118.380 169.175 118.550 169.685 ;
        RECT 118.720 169.425 119.240 169.735 ;
        RECT 116.650 169.005 118.550 169.175 ;
        RECT 116.650 168.945 116.980 169.005 ;
        RECT 117.130 168.775 117.460 168.835 ;
        RECT 116.800 168.505 117.460 168.775 ;
        RECT 116.290 168.120 116.610 168.450 ;
        RECT 116.790 167.855 117.450 168.335 ;
        RECT 117.650 168.245 117.820 169.005 ;
        RECT 118.720 168.835 118.900 169.245 ;
        RECT 117.990 168.665 118.320 168.785 ;
        RECT 119.070 168.665 119.240 169.425 ;
        RECT 117.990 168.495 119.240 168.665 ;
        RECT 119.410 169.605 120.780 169.855 ;
        RECT 119.410 168.835 119.600 169.605 ;
        RECT 120.530 169.345 120.780 169.605 ;
        RECT 119.770 169.175 120.020 169.335 ;
        RECT 120.950 169.175 121.120 170.020 ;
        RECT 122.015 169.735 122.185 170.235 ;
        RECT 122.355 169.905 122.685 170.405 ;
        RECT 121.290 169.345 121.790 169.725 ;
        RECT 122.015 169.565 122.710 169.735 ;
        RECT 119.770 169.005 121.120 169.175 ;
        RECT 120.700 168.965 121.120 169.005 ;
        RECT 119.410 168.495 119.830 168.835 ;
        RECT 120.120 168.505 120.530 168.835 ;
        RECT 117.650 168.075 118.500 168.245 ;
        RECT 119.060 167.855 119.380 168.315 ;
        RECT 119.580 168.065 119.830 168.495 ;
        RECT 120.120 167.855 120.530 168.295 ;
        RECT 120.700 168.235 120.870 168.965 ;
        RECT 121.040 168.415 121.390 168.785 ;
        RECT 121.570 168.475 121.790 169.345 ;
        RECT 121.960 168.775 122.370 169.395 ;
        RECT 122.540 168.595 122.710 169.565 ;
        RECT 122.015 168.405 122.710 168.595 ;
        RECT 120.700 168.035 121.715 168.235 ;
        RECT 122.015 168.075 122.185 168.405 ;
        RECT 122.355 167.855 122.685 168.235 ;
        RECT 122.900 168.115 123.125 170.235 ;
        RECT 123.295 169.905 123.625 170.405 ;
        RECT 123.795 169.735 123.965 170.235 ;
        RECT 124.230 169.980 124.565 170.405 ;
        RECT 124.735 169.800 124.920 170.205 ;
        RECT 123.300 169.565 123.965 169.735 ;
        RECT 124.255 169.625 124.920 169.800 ;
        RECT 125.125 169.625 125.455 170.405 ;
        RECT 123.300 168.575 123.530 169.565 ;
        RECT 123.700 168.745 124.050 169.395 ;
        RECT 124.255 168.595 124.595 169.625 ;
        RECT 125.625 169.435 125.895 170.205 ;
        RECT 124.765 169.265 125.895 169.435 ;
        RECT 124.765 168.765 125.015 169.265 ;
        RECT 123.300 168.405 123.965 168.575 ;
        RECT 124.255 168.425 124.940 168.595 ;
        RECT 125.195 168.515 125.555 169.095 ;
        RECT 123.295 167.855 123.625 168.235 ;
        RECT 123.795 168.115 123.965 168.405 ;
        RECT 124.230 167.855 124.565 168.255 ;
        RECT 124.735 168.025 124.940 168.425 ;
        RECT 125.725 168.355 125.895 169.265 ;
        RECT 126.525 169.315 127.735 170.405 ;
        RECT 126.525 168.775 127.045 169.315 ;
        RECT 127.215 168.605 127.735 169.145 ;
        RECT 125.150 167.855 125.425 168.335 ;
        RECT 125.635 168.025 125.895 168.355 ;
        RECT 126.525 167.855 127.735 168.605 ;
        RECT 14.660 167.685 127.820 167.855 ;
        RECT 14.745 166.935 15.955 167.685 ;
        RECT 14.745 166.395 15.265 166.935 ;
        RECT 16.125 166.915 17.795 167.685 ;
        RECT 15.435 166.225 15.955 166.765 ;
        RECT 14.745 165.135 15.955 166.225 ;
        RECT 16.125 166.225 16.875 166.745 ;
        RECT 17.045 166.395 17.795 166.915 ;
        RECT 17.970 166.975 18.225 167.505 ;
        RECT 18.395 167.225 18.700 167.685 ;
        RECT 18.945 167.305 20.015 167.475 ;
        RECT 17.970 166.325 18.180 166.975 ;
        RECT 18.945 166.950 19.265 167.305 ;
        RECT 18.940 166.775 19.265 166.950 ;
        RECT 18.350 166.475 19.265 166.775 ;
        RECT 19.435 166.735 19.675 167.135 ;
        RECT 19.845 167.075 20.015 167.305 ;
        RECT 20.185 167.245 20.375 167.685 ;
        RECT 20.545 167.235 21.495 167.515 ;
        RECT 21.715 167.325 22.065 167.495 ;
        RECT 19.845 166.905 20.375 167.075 ;
        RECT 18.350 166.445 19.090 166.475 ;
        RECT 16.125 165.135 17.795 166.225 ;
        RECT 17.970 165.445 18.225 166.325 ;
        RECT 18.395 165.135 18.700 166.275 ;
        RECT 18.920 165.855 19.090 166.445 ;
        RECT 19.435 166.365 19.975 166.735 ;
        RECT 20.155 166.625 20.375 166.905 ;
        RECT 20.545 166.455 20.715 167.235 ;
        RECT 20.310 166.285 20.715 166.455 ;
        RECT 20.885 166.445 21.235 167.065 ;
        RECT 20.310 166.195 20.480 166.285 ;
        RECT 21.405 166.275 21.615 167.065 ;
        RECT 19.260 166.025 20.480 166.195 ;
        RECT 20.940 166.115 21.615 166.275 ;
        RECT 18.920 165.685 19.720 165.855 ;
        RECT 19.040 165.135 19.370 165.515 ;
        RECT 19.550 165.395 19.720 165.685 ;
        RECT 20.310 165.645 20.480 166.025 ;
        RECT 20.650 166.105 21.615 166.115 ;
        RECT 21.805 166.935 22.065 167.325 ;
        RECT 22.275 167.225 22.605 167.685 ;
        RECT 23.480 167.295 24.335 167.465 ;
        RECT 24.540 167.295 25.035 167.465 ;
        RECT 25.205 167.325 25.535 167.685 ;
        RECT 21.805 166.245 21.975 166.935 ;
        RECT 22.145 166.585 22.315 166.765 ;
        RECT 22.485 166.755 23.275 167.005 ;
        RECT 23.480 166.585 23.650 167.295 ;
        RECT 23.820 166.785 24.175 167.005 ;
        RECT 22.145 166.415 23.835 166.585 ;
        RECT 20.650 165.815 21.110 166.105 ;
        RECT 21.805 166.075 23.305 166.245 ;
        RECT 21.805 165.935 21.975 166.075 ;
        RECT 21.415 165.765 21.975 165.935 ;
        RECT 19.890 165.135 20.140 165.595 ;
        RECT 20.310 165.305 21.180 165.645 ;
        RECT 21.415 165.305 21.585 165.765 ;
        RECT 22.420 165.735 23.495 165.905 ;
        RECT 21.755 165.135 22.125 165.595 ;
        RECT 22.420 165.395 22.590 165.735 ;
        RECT 22.760 165.135 23.090 165.565 ;
        RECT 23.325 165.395 23.495 165.735 ;
        RECT 23.665 165.635 23.835 166.415 ;
        RECT 24.005 166.195 24.175 166.785 ;
        RECT 24.345 166.385 24.695 167.005 ;
        RECT 24.005 165.805 24.470 166.195 ;
        RECT 24.865 165.935 25.035 167.295 ;
        RECT 25.205 166.105 25.665 167.155 ;
        RECT 24.640 165.765 25.035 165.935 ;
        RECT 24.640 165.635 24.810 165.765 ;
        RECT 23.665 165.305 24.345 165.635 ;
        RECT 24.560 165.305 24.810 165.635 ;
        RECT 24.980 165.135 25.230 165.595 ;
        RECT 25.400 165.320 25.725 166.105 ;
        RECT 25.895 165.305 26.065 167.425 ;
        RECT 26.235 167.305 26.565 167.685 ;
        RECT 26.735 167.135 26.990 167.425 ;
        RECT 26.240 166.965 26.990 167.135 ;
        RECT 26.240 165.975 26.470 166.965 ;
        RECT 27.165 166.915 28.835 167.685 ;
        RECT 29.010 167.140 34.355 167.685 ;
        RECT 34.585 167.205 34.865 167.685 ;
        RECT 26.640 166.145 26.990 166.795 ;
        RECT 27.165 166.225 27.915 166.745 ;
        RECT 28.085 166.395 28.835 166.915 ;
        RECT 26.240 165.805 26.990 165.975 ;
        RECT 26.235 165.135 26.565 165.635 ;
        RECT 26.735 165.305 26.990 165.805 ;
        RECT 27.165 165.135 28.835 166.225 ;
        RECT 30.600 165.570 30.950 166.820 ;
        RECT 32.430 166.310 32.770 167.140 ;
        RECT 35.035 167.035 35.295 167.425 ;
        RECT 35.470 167.205 35.725 167.685 ;
        RECT 35.895 167.035 36.190 167.425 ;
        RECT 36.370 167.205 36.645 167.685 ;
        RECT 36.815 167.185 37.115 167.515 ;
        RECT 34.540 166.865 36.190 167.035 ;
        RECT 34.540 166.355 34.945 166.865 ;
        RECT 35.115 166.525 36.255 166.695 ;
        RECT 34.540 166.185 35.295 166.355 ;
        RECT 29.010 165.135 34.355 165.570 ;
        RECT 34.580 165.135 34.865 166.005 ;
        RECT 35.035 165.935 35.295 166.185 ;
        RECT 36.085 166.275 36.255 166.525 ;
        RECT 36.425 166.445 36.775 167.015 ;
        RECT 36.945 166.275 37.115 167.185 ;
        RECT 37.285 166.960 37.575 167.685 ;
        RECT 37.835 167.135 38.005 167.515 ;
        RECT 38.185 167.305 38.515 167.685 ;
        RECT 37.835 166.965 38.500 167.135 ;
        RECT 38.695 167.010 38.955 167.515 ;
        RECT 37.765 166.415 38.095 166.785 ;
        RECT 38.330 166.710 38.500 166.965 ;
        RECT 38.330 166.380 38.615 166.710 ;
        RECT 36.085 166.105 37.115 166.275 ;
        RECT 35.035 165.765 36.155 165.935 ;
        RECT 35.035 165.305 35.295 165.765 ;
        RECT 35.470 165.135 35.725 165.595 ;
        RECT 35.895 165.305 36.155 165.765 ;
        RECT 36.325 165.135 36.635 165.935 ;
        RECT 36.805 165.305 37.115 166.105 ;
        RECT 37.285 165.135 37.575 166.300 ;
        RECT 38.330 166.235 38.500 166.380 ;
        RECT 37.835 166.065 38.500 166.235 ;
        RECT 38.785 166.210 38.955 167.010 ;
        RECT 40.250 166.905 40.750 167.515 ;
        RECT 40.045 166.445 40.395 166.695 ;
        RECT 40.580 166.275 40.750 166.905 ;
        RECT 41.380 167.035 41.710 167.515 ;
        RECT 41.880 167.225 42.105 167.685 ;
        RECT 42.275 167.035 42.605 167.515 ;
        RECT 41.380 166.865 42.605 167.035 ;
        RECT 42.795 166.885 43.045 167.685 ;
        RECT 43.215 166.885 43.555 167.515 ;
        RECT 43.930 166.905 44.430 167.515 ;
        RECT 40.920 166.495 41.250 166.695 ;
        RECT 41.420 166.495 41.750 166.695 ;
        RECT 41.920 166.495 42.340 166.695 ;
        RECT 42.515 166.525 43.210 166.695 ;
        RECT 42.515 166.275 42.685 166.525 ;
        RECT 43.380 166.275 43.555 166.885 ;
        RECT 43.725 166.445 44.075 166.695 ;
        RECT 44.260 166.275 44.430 166.905 ;
        RECT 45.060 167.035 45.390 167.515 ;
        RECT 45.560 167.225 45.785 167.685 ;
        RECT 45.955 167.035 46.285 167.515 ;
        RECT 45.060 166.865 46.285 167.035 ;
        RECT 46.475 166.885 46.725 167.685 ;
        RECT 46.895 166.885 47.235 167.515 ;
        RECT 47.610 166.905 48.110 167.515 ;
        RECT 44.600 166.495 44.930 166.695 ;
        RECT 45.100 166.495 45.430 166.695 ;
        RECT 45.600 166.495 46.020 166.695 ;
        RECT 46.195 166.525 46.890 166.695 ;
        RECT 46.195 166.275 46.365 166.525 ;
        RECT 47.060 166.275 47.235 166.885 ;
        RECT 47.405 166.445 47.755 166.695 ;
        RECT 47.940 166.275 48.110 166.905 ;
        RECT 48.740 167.035 49.070 167.515 ;
        RECT 49.240 167.225 49.465 167.685 ;
        RECT 49.635 167.035 49.965 167.515 ;
        RECT 48.740 166.865 49.965 167.035 ;
        RECT 50.155 166.885 50.405 167.685 ;
        RECT 50.575 166.885 50.915 167.515 ;
        RECT 48.280 166.495 48.610 166.695 ;
        RECT 48.780 166.495 49.110 166.695 ;
        RECT 49.280 166.495 49.700 166.695 ;
        RECT 49.875 166.525 50.570 166.695 ;
        RECT 49.875 166.275 50.045 166.525 ;
        RECT 50.740 166.325 50.915 166.885 ;
        RECT 50.685 166.275 50.915 166.325 ;
        RECT 37.835 165.305 38.005 166.065 ;
        RECT 38.185 165.135 38.515 165.895 ;
        RECT 38.685 165.305 38.955 166.210 ;
        RECT 40.250 166.105 42.685 166.275 ;
        RECT 40.250 165.305 40.580 166.105 ;
        RECT 40.750 165.135 41.080 165.935 ;
        RECT 41.380 165.305 41.710 166.105 ;
        RECT 42.355 165.135 42.605 165.935 ;
        RECT 42.875 165.135 43.045 166.275 ;
        RECT 43.215 165.305 43.555 166.275 ;
        RECT 43.930 166.105 46.365 166.275 ;
        RECT 43.930 165.305 44.260 166.105 ;
        RECT 44.430 165.135 44.760 165.935 ;
        RECT 45.060 165.305 45.390 166.105 ;
        RECT 46.035 165.135 46.285 165.935 ;
        RECT 46.555 165.135 46.725 166.275 ;
        RECT 46.895 165.305 47.235 166.275 ;
        RECT 47.610 166.105 50.045 166.275 ;
        RECT 47.610 165.305 47.940 166.105 ;
        RECT 48.110 165.135 48.440 165.935 ;
        RECT 48.740 165.305 49.070 166.105 ;
        RECT 49.715 165.135 49.965 165.935 ;
        RECT 50.235 165.135 50.405 166.275 ;
        RECT 50.575 165.305 50.915 166.275 ;
        RECT 51.085 166.885 51.425 167.515 ;
        RECT 51.595 166.885 51.845 167.685 ;
        RECT 52.035 167.035 52.365 167.515 ;
        RECT 52.535 167.225 52.760 167.685 ;
        RECT 52.930 167.035 53.260 167.515 ;
        RECT 51.085 166.275 51.260 166.885 ;
        RECT 52.035 166.865 53.260 167.035 ;
        RECT 53.890 166.905 54.390 167.515 ;
        RECT 51.430 166.525 52.125 166.695 ;
        RECT 51.955 166.275 52.125 166.525 ;
        RECT 52.300 166.495 52.720 166.695 ;
        RECT 52.890 166.495 53.220 166.695 ;
        RECT 53.390 166.495 53.720 166.695 ;
        RECT 53.890 166.275 54.060 166.905 ;
        RECT 54.915 166.885 55.245 167.685 ;
        RECT 55.415 167.035 55.585 167.515 ;
        RECT 55.755 167.205 56.085 167.685 ;
        RECT 56.255 167.035 56.425 167.515 ;
        RECT 56.675 167.205 56.915 167.685 ;
        RECT 57.095 167.035 57.265 167.515 ;
        RECT 55.415 166.865 56.425 167.035 ;
        RECT 56.630 166.865 57.265 167.035 ;
        RECT 57.985 166.915 61.495 167.685 ;
        RECT 54.245 166.445 54.595 166.695 ;
        RECT 55.415 166.665 55.910 166.865 ;
        RECT 56.630 166.695 56.800 166.865 ;
        RECT 55.415 166.495 55.915 166.665 ;
        RECT 56.300 166.525 56.800 166.695 ;
        RECT 55.415 166.325 55.910 166.495 ;
        RECT 51.085 165.305 51.425 166.275 ;
        RECT 51.595 165.135 51.765 166.275 ;
        RECT 51.955 166.105 54.390 166.275 ;
        RECT 52.035 165.135 52.285 165.935 ;
        RECT 52.930 165.305 53.260 166.105 ;
        RECT 53.560 165.135 53.890 165.935 ;
        RECT 54.060 165.305 54.390 166.105 ;
        RECT 54.915 165.135 55.245 166.285 ;
        RECT 55.415 166.155 56.425 166.325 ;
        RECT 55.415 165.305 55.585 166.155 ;
        RECT 55.755 165.135 56.085 165.935 ;
        RECT 56.255 165.305 56.425 166.155 ;
        RECT 56.630 166.285 56.800 166.525 ;
        RECT 56.970 166.455 57.350 166.695 ;
        RECT 56.630 166.115 57.345 166.285 ;
        RECT 56.605 165.135 56.845 165.935 ;
        RECT 57.015 165.305 57.345 166.115 ;
        RECT 57.985 166.225 59.675 166.745 ;
        RECT 59.845 166.395 61.495 166.915 ;
        RECT 61.705 166.865 61.935 167.685 ;
        RECT 62.105 166.885 62.435 167.515 ;
        RECT 61.685 166.445 62.015 166.695 ;
        RECT 62.185 166.285 62.435 166.885 ;
        RECT 62.605 166.865 62.815 167.685 ;
        RECT 63.045 166.960 63.335 167.685 ;
        RECT 63.965 166.915 65.635 167.685 ;
        RECT 65.895 167.135 66.065 167.515 ;
        RECT 66.280 167.305 66.610 167.685 ;
        RECT 65.895 166.965 66.610 167.135 ;
        RECT 57.985 165.135 61.495 166.225 ;
        RECT 61.705 165.135 61.935 166.275 ;
        RECT 62.105 165.305 62.435 166.285 ;
        RECT 62.605 165.135 62.815 166.275 ;
        RECT 63.045 165.135 63.335 166.300 ;
        RECT 63.965 166.225 64.715 166.745 ;
        RECT 64.885 166.395 65.635 166.915 ;
        RECT 65.805 166.415 66.160 166.785 ;
        RECT 66.440 166.775 66.610 166.965 ;
        RECT 66.780 166.940 67.035 167.515 ;
        RECT 66.440 166.445 66.695 166.775 ;
        RECT 66.440 166.235 66.610 166.445 ;
        RECT 63.965 165.135 65.635 166.225 ;
        RECT 65.895 166.065 66.610 166.235 ;
        RECT 66.865 166.210 67.035 166.940 ;
        RECT 67.210 166.845 67.470 167.685 ;
        RECT 68.570 167.140 73.915 167.685 ;
        RECT 65.895 165.305 66.065 166.065 ;
        RECT 66.280 165.135 66.610 165.895 ;
        RECT 66.780 165.305 67.035 166.210 ;
        RECT 67.210 165.135 67.470 166.285 ;
        RECT 70.160 165.570 70.510 166.820 ;
        RECT 71.990 166.310 72.330 167.140 ;
        RECT 74.090 166.845 74.350 167.685 ;
        RECT 74.525 166.940 74.780 167.515 ;
        RECT 74.950 167.305 75.280 167.685 ;
        RECT 75.495 167.135 75.665 167.515 ;
        RECT 74.950 166.965 75.665 167.135 ;
        RECT 68.570 165.135 73.915 165.570 ;
        RECT 74.090 165.135 74.350 166.285 ;
        RECT 74.525 166.210 74.695 166.940 ;
        RECT 74.950 166.775 75.120 166.965 ;
        RECT 76.590 166.905 77.090 167.515 ;
        RECT 74.865 166.445 75.120 166.775 ;
        RECT 74.950 166.235 75.120 166.445 ;
        RECT 75.400 166.415 75.755 166.785 ;
        RECT 76.385 166.445 76.735 166.695 ;
        RECT 76.920 166.275 77.090 166.905 ;
        RECT 77.720 167.035 78.050 167.515 ;
        RECT 78.220 167.225 78.445 167.685 ;
        RECT 78.615 167.035 78.945 167.515 ;
        RECT 77.720 166.865 78.945 167.035 ;
        RECT 79.135 166.885 79.385 167.685 ;
        RECT 79.555 166.885 79.895 167.515 ;
        RECT 80.270 166.905 80.770 167.515 ;
        RECT 77.260 166.495 77.590 166.695 ;
        RECT 77.760 166.495 78.090 166.695 ;
        RECT 78.260 166.495 78.680 166.695 ;
        RECT 78.855 166.525 79.550 166.695 ;
        RECT 78.855 166.275 79.025 166.525 ;
        RECT 79.720 166.275 79.895 166.885 ;
        RECT 80.065 166.445 80.415 166.695 ;
        RECT 80.600 166.275 80.770 166.905 ;
        RECT 81.400 167.035 81.730 167.515 ;
        RECT 81.900 167.225 82.125 167.685 ;
        RECT 82.295 167.035 82.625 167.515 ;
        RECT 81.400 166.865 82.625 167.035 ;
        RECT 82.815 166.885 83.065 167.685 ;
        RECT 83.235 166.885 83.575 167.515 ;
        RECT 80.940 166.495 81.270 166.695 ;
        RECT 81.440 166.495 81.770 166.695 ;
        RECT 81.940 166.495 82.360 166.695 ;
        RECT 82.535 166.525 83.230 166.695 ;
        RECT 82.535 166.275 82.705 166.525 ;
        RECT 83.400 166.275 83.575 166.885 ;
        RECT 74.525 165.305 74.780 166.210 ;
        RECT 74.950 166.065 75.665 166.235 ;
        RECT 74.950 165.135 75.280 165.895 ;
        RECT 75.495 165.305 75.665 166.065 ;
        RECT 76.590 166.105 79.025 166.275 ;
        RECT 76.590 165.305 76.920 166.105 ;
        RECT 77.090 165.135 77.420 165.935 ;
        RECT 77.720 165.305 78.050 166.105 ;
        RECT 78.695 165.135 78.945 165.935 ;
        RECT 79.215 165.135 79.385 166.275 ;
        RECT 79.555 165.305 79.895 166.275 ;
        RECT 80.270 166.105 82.705 166.275 ;
        RECT 80.270 165.305 80.600 166.105 ;
        RECT 80.770 165.135 81.100 165.935 ;
        RECT 81.400 165.305 81.730 166.105 ;
        RECT 82.375 165.135 82.625 165.935 ;
        RECT 82.895 165.135 83.065 166.275 ;
        RECT 83.235 165.305 83.575 166.275 ;
        RECT 84.210 166.945 84.465 167.515 ;
        RECT 84.635 167.285 84.965 167.685 ;
        RECT 85.390 167.150 85.920 167.515 ;
        RECT 85.390 167.115 85.565 167.150 ;
        RECT 84.635 166.945 85.565 167.115 ;
        RECT 84.210 166.275 84.380 166.945 ;
        RECT 84.635 166.775 84.805 166.945 ;
        RECT 84.550 166.445 84.805 166.775 ;
        RECT 85.030 166.445 85.225 166.775 ;
        RECT 84.210 165.305 84.545 166.275 ;
        RECT 84.715 165.135 84.885 166.275 ;
        RECT 85.055 165.475 85.225 166.445 ;
        RECT 85.395 165.815 85.565 166.945 ;
        RECT 85.735 166.155 85.905 166.955 ;
        RECT 86.110 166.665 86.385 167.515 ;
        RECT 86.105 166.495 86.385 166.665 ;
        RECT 86.110 166.355 86.385 166.495 ;
        RECT 86.555 166.155 86.745 167.515 ;
        RECT 86.925 167.150 87.435 167.685 ;
        RECT 87.655 166.875 87.900 167.480 ;
        RECT 88.805 166.960 89.095 167.685 ;
        RECT 89.265 166.915 92.775 167.685 ;
        RECT 93.035 167.135 93.205 167.515 ;
        RECT 93.385 167.305 93.715 167.685 ;
        RECT 93.035 166.965 93.700 167.135 ;
        RECT 93.895 167.010 94.155 167.515 ;
        RECT 86.945 166.705 88.175 166.875 ;
        RECT 85.735 165.985 86.745 166.155 ;
        RECT 86.915 166.140 87.665 166.330 ;
        RECT 85.395 165.645 86.520 165.815 ;
        RECT 86.915 165.475 87.085 166.140 ;
        RECT 87.835 165.895 88.175 166.705 ;
        RECT 85.055 165.305 87.085 165.475 ;
        RECT 87.255 165.135 87.425 165.895 ;
        RECT 87.660 165.485 88.175 165.895 ;
        RECT 88.805 165.135 89.095 166.300 ;
        RECT 89.265 166.225 90.955 166.745 ;
        RECT 91.125 166.395 92.775 166.915 ;
        RECT 92.965 166.415 93.295 166.785 ;
        RECT 93.530 166.710 93.700 166.965 ;
        RECT 93.530 166.380 93.815 166.710 ;
        RECT 93.530 166.235 93.700 166.380 ;
        RECT 89.265 165.135 92.775 166.225 ;
        RECT 93.035 166.065 93.700 166.235 ;
        RECT 93.985 166.210 94.155 167.010 ;
        RECT 95.285 166.865 95.515 167.685 ;
        RECT 95.685 166.885 96.015 167.515 ;
        RECT 95.265 166.445 95.595 166.695 ;
        RECT 95.765 166.285 96.015 166.885 ;
        RECT 96.185 166.865 96.395 167.685 ;
        RECT 97.000 166.975 97.255 167.505 ;
        RECT 97.435 167.225 97.720 167.685 ;
        RECT 97.000 166.325 97.180 166.975 ;
        RECT 97.900 166.775 98.150 167.425 ;
        RECT 97.350 166.445 98.150 166.775 ;
        RECT 93.035 165.305 93.205 166.065 ;
        RECT 93.385 165.135 93.715 165.895 ;
        RECT 93.885 165.305 94.155 166.210 ;
        RECT 95.285 165.135 95.515 166.275 ;
        RECT 95.685 165.305 96.015 166.285 ;
        RECT 96.185 165.135 96.395 166.275 ;
        RECT 96.915 166.155 97.180 166.325 ;
        RECT 97.000 166.115 97.180 166.155 ;
        RECT 97.000 165.445 97.255 166.115 ;
        RECT 97.435 165.135 97.720 165.935 ;
        RECT 97.900 165.855 98.150 166.445 ;
        RECT 98.350 167.090 98.670 167.420 ;
        RECT 98.850 167.205 99.510 167.685 ;
        RECT 99.710 167.295 100.560 167.465 ;
        RECT 98.350 166.195 98.540 167.090 ;
        RECT 98.860 166.765 99.520 167.035 ;
        RECT 99.190 166.705 99.520 166.765 ;
        RECT 98.710 166.535 99.040 166.595 ;
        RECT 99.710 166.535 99.880 167.295 ;
        RECT 101.120 167.225 101.440 167.685 ;
        RECT 101.640 167.045 101.890 167.475 ;
        RECT 102.180 167.245 102.590 167.685 ;
        RECT 102.760 167.305 103.775 167.505 ;
        RECT 100.050 166.875 101.300 167.045 ;
        RECT 100.050 166.755 100.380 166.875 ;
        RECT 98.710 166.365 100.610 166.535 ;
        RECT 98.350 166.025 100.270 166.195 ;
        RECT 98.350 166.005 98.670 166.025 ;
        RECT 97.900 165.345 98.230 165.855 ;
        RECT 98.500 165.395 98.670 166.005 ;
        RECT 100.440 165.855 100.610 166.365 ;
        RECT 100.780 166.295 100.960 166.705 ;
        RECT 101.130 166.115 101.300 166.875 ;
        RECT 98.840 165.135 99.170 165.825 ;
        RECT 99.400 165.685 100.610 165.855 ;
        RECT 100.780 165.805 101.300 166.115 ;
        RECT 101.470 166.705 101.890 167.045 ;
        RECT 102.180 166.705 102.590 167.035 ;
        RECT 101.470 165.935 101.660 166.705 ;
        RECT 102.760 166.575 102.930 167.305 ;
        RECT 104.075 167.135 104.245 167.465 ;
        RECT 104.415 167.305 104.745 167.685 ;
        RECT 103.100 166.755 103.450 167.125 ;
        RECT 102.760 166.535 103.180 166.575 ;
        RECT 101.830 166.365 103.180 166.535 ;
        RECT 101.830 166.205 102.080 166.365 ;
        RECT 102.590 165.935 102.840 166.195 ;
        RECT 101.470 165.685 102.840 165.935 ;
        RECT 99.400 165.395 99.640 165.685 ;
        RECT 100.440 165.605 100.610 165.685 ;
        RECT 99.840 165.135 100.260 165.515 ;
        RECT 100.440 165.355 101.070 165.605 ;
        RECT 101.540 165.135 101.870 165.515 ;
        RECT 102.040 165.395 102.210 165.685 ;
        RECT 103.010 165.520 103.180 166.365 ;
        RECT 103.630 166.195 103.850 167.065 ;
        RECT 104.075 166.945 104.770 167.135 ;
        RECT 103.350 165.815 103.850 166.195 ;
        RECT 104.020 166.145 104.430 166.765 ;
        RECT 104.600 165.975 104.770 166.945 ;
        RECT 104.075 165.805 104.770 165.975 ;
        RECT 102.390 165.135 102.770 165.515 ;
        RECT 103.010 165.350 103.840 165.520 ;
        RECT 104.075 165.305 104.245 165.805 ;
        RECT 104.415 165.135 104.745 165.635 ;
        RECT 104.960 165.305 105.185 167.425 ;
        RECT 105.355 167.305 105.685 167.685 ;
        RECT 105.855 167.135 106.025 167.425 ;
        RECT 105.360 166.965 106.025 167.135 ;
        RECT 105.360 165.975 105.590 166.965 ;
        RECT 106.285 166.915 107.955 167.685 ;
        RECT 105.760 166.145 106.110 166.795 ;
        RECT 106.285 166.225 107.035 166.745 ;
        RECT 107.205 166.395 107.955 166.915 ;
        RECT 108.125 166.885 108.465 167.515 ;
        RECT 108.635 166.885 108.885 167.685 ;
        RECT 109.075 167.035 109.405 167.515 ;
        RECT 109.575 167.225 109.800 167.685 ;
        RECT 109.970 167.035 110.300 167.515 ;
        RECT 108.125 166.275 108.300 166.885 ;
        RECT 109.075 166.865 110.300 167.035 ;
        RECT 110.930 166.905 111.430 167.515 ;
        RECT 111.805 166.915 114.395 167.685 ;
        RECT 114.565 166.960 114.855 167.685 ;
        RECT 108.470 166.525 109.165 166.695 ;
        RECT 108.995 166.275 109.165 166.525 ;
        RECT 109.340 166.495 109.760 166.695 ;
        RECT 109.930 166.495 110.260 166.695 ;
        RECT 110.430 166.495 110.760 166.695 ;
        RECT 110.930 166.275 111.100 166.905 ;
        RECT 111.285 166.445 111.635 166.695 ;
        RECT 105.360 165.805 106.025 165.975 ;
        RECT 105.355 165.135 105.685 165.635 ;
        RECT 105.855 165.305 106.025 165.805 ;
        RECT 106.285 165.135 107.955 166.225 ;
        RECT 108.125 165.305 108.465 166.275 ;
        RECT 108.635 165.135 108.805 166.275 ;
        RECT 108.995 166.105 111.430 166.275 ;
        RECT 109.075 165.135 109.325 165.935 ;
        RECT 109.970 165.305 110.300 166.105 ;
        RECT 110.600 165.135 110.930 165.935 ;
        RECT 111.100 165.305 111.430 166.105 ;
        RECT 111.805 166.225 113.015 166.745 ;
        RECT 113.185 166.395 114.395 166.915 ;
        RECT 115.985 166.865 116.215 167.685 ;
        RECT 116.385 166.885 116.715 167.515 ;
        RECT 115.965 166.445 116.295 166.695 ;
        RECT 111.805 165.135 114.395 166.225 ;
        RECT 114.565 165.135 114.855 166.300 ;
        RECT 116.465 166.285 116.715 166.885 ;
        RECT 116.885 166.865 117.095 167.685 ;
        RECT 117.475 166.885 117.805 167.685 ;
        RECT 117.975 167.035 118.145 167.515 ;
        RECT 118.315 167.205 118.645 167.685 ;
        RECT 118.815 167.035 118.985 167.515 ;
        RECT 119.235 167.205 119.475 167.685 ;
        RECT 119.655 167.035 119.825 167.515 ;
        RECT 121.010 167.140 126.355 167.685 ;
        RECT 117.975 166.865 118.985 167.035 ;
        RECT 119.190 166.865 119.825 167.035 ;
        RECT 117.975 166.665 118.470 166.865 ;
        RECT 119.190 166.695 119.360 166.865 ;
        RECT 117.975 166.495 118.475 166.665 ;
        RECT 118.860 166.525 119.360 166.695 ;
        RECT 117.975 166.325 118.470 166.495 ;
        RECT 115.985 165.135 116.215 166.275 ;
        RECT 116.385 165.305 116.715 166.285 ;
        RECT 116.885 165.135 117.095 166.275 ;
        RECT 117.475 165.135 117.805 166.285 ;
        RECT 117.975 166.155 118.985 166.325 ;
        RECT 117.975 165.305 118.145 166.155 ;
        RECT 118.315 165.135 118.645 165.935 ;
        RECT 118.815 165.305 118.985 166.155 ;
        RECT 119.190 166.285 119.360 166.525 ;
        RECT 119.530 166.455 119.910 166.695 ;
        RECT 119.190 166.115 119.905 166.285 ;
        RECT 119.165 165.135 119.405 165.935 ;
        RECT 119.575 165.305 119.905 166.115 ;
        RECT 122.600 165.570 122.950 166.820 ;
        RECT 124.430 166.310 124.770 167.140 ;
        RECT 126.525 166.935 127.735 167.685 ;
        RECT 126.525 166.225 127.045 166.765 ;
        RECT 127.215 166.395 127.735 166.935 ;
        RECT 121.010 165.135 126.355 165.570 ;
        RECT 126.525 165.135 127.735 166.225 ;
        RECT 14.660 164.965 127.820 165.135 ;
        RECT 14.745 163.875 15.955 164.965 ;
        RECT 14.745 163.165 15.265 163.705 ;
        RECT 15.435 163.335 15.955 163.875 ;
        RECT 16.585 163.875 20.095 164.965 ;
        RECT 20.265 164.205 20.780 164.615 ;
        RECT 21.015 164.205 21.185 164.965 ;
        RECT 21.355 164.625 23.385 164.795 ;
        RECT 16.585 163.355 18.275 163.875 ;
        RECT 18.445 163.185 20.095 163.705 ;
        RECT 20.265 163.395 20.605 164.205 ;
        RECT 21.355 163.960 21.525 164.625 ;
        RECT 21.920 164.285 23.045 164.455 ;
        RECT 20.775 163.770 21.525 163.960 ;
        RECT 21.695 163.945 22.705 164.115 ;
        RECT 20.265 163.225 21.495 163.395 ;
        RECT 14.745 162.415 15.955 163.165 ;
        RECT 16.585 162.415 20.095 163.185 ;
        RECT 20.540 162.620 20.785 163.225 ;
        RECT 21.005 162.415 21.515 162.950 ;
        RECT 21.695 162.585 21.885 163.945 ;
        RECT 22.055 162.925 22.330 163.745 ;
        RECT 22.535 163.145 22.705 163.945 ;
        RECT 22.875 163.155 23.045 164.285 ;
        RECT 23.215 163.655 23.385 164.625 ;
        RECT 23.555 163.825 23.725 164.965 ;
        RECT 23.895 163.825 24.230 164.795 ;
        RECT 23.215 163.325 23.410 163.655 ;
        RECT 23.635 163.325 23.890 163.655 ;
        RECT 23.635 163.155 23.805 163.325 ;
        RECT 24.060 163.155 24.230 163.825 ;
        RECT 24.405 163.800 24.695 164.965 ;
        RECT 24.955 164.035 25.125 164.795 ;
        RECT 25.305 164.205 25.635 164.965 ;
        RECT 24.955 163.865 25.620 164.035 ;
        RECT 25.805 163.890 26.075 164.795 ;
        RECT 25.450 163.720 25.620 163.865 ;
        RECT 24.885 163.315 25.215 163.685 ;
        RECT 25.450 163.390 25.735 163.720 ;
        RECT 22.875 162.985 23.805 163.155 ;
        RECT 22.875 162.950 23.050 162.985 ;
        RECT 22.055 162.755 22.335 162.925 ;
        RECT 22.055 162.585 22.330 162.755 ;
        RECT 22.520 162.585 23.050 162.950 ;
        RECT 23.475 162.415 23.805 162.815 ;
        RECT 23.975 162.585 24.230 163.155 ;
        RECT 24.405 162.415 24.695 163.140 ;
        RECT 25.450 163.135 25.620 163.390 ;
        RECT 24.955 162.965 25.620 163.135 ;
        RECT 25.905 163.090 26.075 163.890 ;
        RECT 26.705 163.875 28.375 164.965 ;
        RECT 26.705 163.355 27.455 163.875 ;
        RECT 28.585 163.825 28.815 164.965 ;
        RECT 28.985 163.815 29.315 164.795 ;
        RECT 29.485 163.825 29.695 164.965 ;
        RECT 29.965 163.825 30.195 164.965 ;
        RECT 30.365 163.815 30.695 164.795 ;
        RECT 30.865 163.825 31.075 164.965 ;
        RECT 27.625 163.185 28.375 163.705 ;
        RECT 28.565 163.405 28.895 163.655 ;
        RECT 24.955 162.585 25.125 162.965 ;
        RECT 25.305 162.415 25.635 162.795 ;
        RECT 25.815 162.585 26.075 163.090 ;
        RECT 26.705 162.415 28.375 163.185 ;
        RECT 28.585 162.415 28.815 163.235 ;
        RECT 29.065 163.215 29.315 163.815 ;
        RECT 29.945 163.405 30.275 163.655 ;
        RECT 28.985 162.585 29.315 163.215 ;
        RECT 29.485 162.415 29.695 163.235 ;
        RECT 29.965 162.415 30.195 163.235 ;
        RECT 30.445 163.215 30.695 163.815 ;
        RECT 31.310 163.775 31.565 164.655 ;
        RECT 31.735 163.825 32.040 164.965 ;
        RECT 32.380 164.585 32.710 164.965 ;
        RECT 32.890 164.415 33.060 164.705 ;
        RECT 33.230 164.505 33.480 164.965 ;
        RECT 32.260 164.245 33.060 164.415 ;
        RECT 33.650 164.455 34.520 164.795 ;
        RECT 30.365 162.585 30.695 163.215 ;
        RECT 30.865 162.415 31.075 163.235 ;
        RECT 31.310 163.125 31.520 163.775 ;
        RECT 32.260 163.655 32.430 164.245 ;
        RECT 33.650 164.075 33.820 164.455 ;
        RECT 34.755 164.335 34.925 164.795 ;
        RECT 35.095 164.505 35.465 164.965 ;
        RECT 35.760 164.365 35.930 164.705 ;
        RECT 36.100 164.535 36.430 164.965 ;
        RECT 36.665 164.365 36.835 164.705 ;
        RECT 32.600 163.905 33.820 164.075 ;
        RECT 33.990 163.995 34.450 164.285 ;
        RECT 34.755 164.165 35.315 164.335 ;
        RECT 35.760 164.195 36.835 164.365 ;
        RECT 37.005 164.465 37.685 164.795 ;
        RECT 37.900 164.465 38.150 164.795 ;
        RECT 38.320 164.505 38.570 164.965 ;
        RECT 35.145 164.025 35.315 164.165 ;
        RECT 33.990 163.985 34.955 163.995 ;
        RECT 33.650 163.815 33.820 163.905 ;
        RECT 34.280 163.825 34.955 163.985 ;
        RECT 31.690 163.625 32.430 163.655 ;
        RECT 31.690 163.325 32.605 163.625 ;
        RECT 32.280 163.150 32.605 163.325 ;
        RECT 31.310 162.595 31.565 163.125 ;
        RECT 31.735 162.415 32.040 162.875 ;
        RECT 32.285 162.795 32.605 163.150 ;
        RECT 32.775 163.365 33.315 163.735 ;
        RECT 33.650 163.645 34.055 163.815 ;
        RECT 32.775 162.965 33.015 163.365 ;
        RECT 33.495 163.195 33.715 163.475 ;
        RECT 33.185 163.025 33.715 163.195 ;
        RECT 33.185 162.795 33.355 163.025 ;
        RECT 33.885 162.865 34.055 163.645 ;
        RECT 34.225 163.035 34.575 163.655 ;
        RECT 34.745 163.035 34.955 163.825 ;
        RECT 35.145 163.855 36.645 164.025 ;
        RECT 35.145 163.165 35.315 163.855 ;
        RECT 37.005 163.685 37.175 164.465 ;
        RECT 37.980 164.335 38.150 164.465 ;
        RECT 35.485 163.515 37.175 163.685 ;
        RECT 37.345 163.905 37.810 164.295 ;
        RECT 37.980 164.165 38.375 164.335 ;
        RECT 35.485 163.335 35.655 163.515 ;
        RECT 32.285 162.625 33.355 162.795 ;
        RECT 33.525 162.415 33.715 162.855 ;
        RECT 33.885 162.585 34.835 162.865 ;
        RECT 35.145 162.775 35.405 163.165 ;
        RECT 35.825 163.095 36.615 163.345 ;
        RECT 35.055 162.605 35.405 162.775 ;
        RECT 35.615 162.415 35.945 162.875 ;
        RECT 36.820 162.805 36.990 163.515 ;
        RECT 37.345 163.315 37.515 163.905 ;
        RECT 37.160 163.095 37.515 163.315 ;
        RECT 37.685 163.095 38.035 163.715 ;
        RECT 38.205 162.805 38.375 164.165 ;
        RECT 38.740 163.995 39.065 164.780 ;
        RECT 38.545 162.945 39.005 163.995 ;
        RECT 36.820 162.635 37.675 162.805 ;
        RECT 37.880 162.635 38.375 162.805 ;
        RECT 38.545 162.415 38.875 162.775 ;
        RECT 39.235 162.675 39.405 164.795 ;
        RECT 39.575 164.465 39.905 164.965 ;
        RECT 40.075 164.295 40.330 164.795 ;
        RECT 39.580 164.125 40.330 164.295 ;
        RECT 39.580 163.135 39.810 164.125 ;
        RECT 41.170 163.995 41.500 164.795 ;
        RECT 41.670 164.165 42.000 164.965 ;
        RECT 42.300 163.995 42.630 164.795 ;
        RECT 43.275 164.165 43.525 164.965 ;
        RECT 39.980 163.305 40.330 163.955 ;
        RECT 41.170 163.825 43.605 163.995 ;
        RECT 43.795 163.825 43.965 164.965 ;
        RECT 44.135 163.825 44.475 164.795 ;
        RECT 44.850 163.995 45.180 164.795 ;
        RECT 45.350 164.165 45.680 164.965 ;
        RECT 45.980 163.995 46.310 164.795 ;
        RECT 46.955 164.165 47.205 164.965 ;
        RECT 44.850 163.825 47.285 163.995 ;
        RECT 47.475 163.825 47.645 164.965 ;
        RECT 47.815 163.825 48.155 164.795 ;
        RECT 40.965 163.405 41.315 163.655 ;
        RECT 41.500 163.195 41.670 163.825 ;
        RECT 41.840 163.405 42.170 163.605 ;
        RECT 42.340 163.405 42.670 163.605 ;
        RECT 42.840 163.405 43.260 163.605 ;
        RECT 43.435 163.575 43.605 163.825 ;
        RECT 43.435 163.405 44.130 163.575 ;
        RECT 39.580 162.965 40.330 163.135 ;
        RECT 39.575 162.415 39.905 162.795 ;
        RECT 40.075 162.675 40.330 162.965 ;
        RECT 41.170 162.585 41.670 163.195 ;
        RECT 42.300 163.065 43.525 163.235 ;
        RECT 44.300 163.215 44.475 163.825 ;
        RECT 44.645 163.405 44.995 163.655 ;
        RECT 42.300 162.585 42.630 163.065 ;
        RECT 42.800 162.415 43.025 162.875 ;
        RECT 43.195 162.585 43.525 163.065 ;
        RECT 43.715 162.415 43.965 163.215 ;
        RECT 44.135 162.585 44.475 163.215 ;
        RECT 45.180 163.195 45.350 163.825 ;
        RECT 45.520 163.405 45.850 163.605 ;
        RECT 46.020 163.405 46.350 163.605 ;
        RECT 46.520 163.405 46.940 163.605 ;
        RECT 47.115 163.575 47.285 163.825 ;
        RECT 47.115 163.405 47.810 163.575 ;
        RECT 44.850 162.585 45.350 163.195 ;
        RECT 45.980 163.065 47.205 163.235 ;
        RECT 47.980 163.215 48.155 163.825 ;
        RECT 48.325 163.875 49.995 164.965 ;
        RECT 48.325 163.355 49.075 163.875 ;
        RECT 50.165 163.800 50.455 164.965 ;
        RECT 50.625 163.875 54.135 164.965 ;
        RECT 54.310 164.530 59.655 164.965 ;
        RECT 45.980 162.585 46.310 163.065 ;
        RECT 46.480 162.415 46.705 162.875 ;
        RECT 46.875 162.585 47.205 163.065 ;
        RECT 47.395 162.415 47.645 163.215 ;
        RECT 47.815 162.585 48.155 163.215 ;
        RECT 49.245 163.185 49.995 163.705 ;
        RECT 50.625 163.355 52.315 163.875 ;
        RECT 52.485 163.185 54.135 163.705 ;
        RECT 55.900 163.280 56.250 164.530 ;
        RECT 60.200 163.985 60.455 164.655 ;
        RECT 60.635 164.165 60.920 164.965 ;
        RECT 61.100 164.245 61.430 164.755 ;
        RECT 48.325 162.415 49.995 163.185 ;
        RECT 50.165 162.415 50.455 163.140 ;
        RECT 50.625 162.415 54.135 163.185 ;
        RECT 57.730 162.960 58.070 163.790 ;
        RECT 60.200 163.125 60.380 163.985 ;
        RECT 61.100 163.655 61.350 164.245 ;
        RECT 61.700 164.095 61.870 164.705 ;
        RECT 62.040 164.275 62.370 164.965 ;
        RECT 62.600 164.415 62.840 164.705 ;
        RECT 63.040 164.585 63.460 164.965 ;
        RECT 63.640 164.495 64.270 164.745 ;
        RECT 64.740 164.585 65.070 164.965 ;
        RECT 63.640 164.415 63.810 164.495 ;
        RECT 65.240 164.415 65.410 164.705 ;
        RECT 65.590 164.585 65.970 164.965 ;
        RECT 66.210 164.580 67.040 164.750 ;
        RECT 62.600 164.245 63.810 164.415 ;
        RECT 60.550 163.325 61.350 163.655 ;
        RECT 54.310 162.415 59.655 162.960 ;
        RECT 60.200 162.925 60.455 163.125 ;
        RECT 60.115 162.755 60.455 162.925 ;
        RECT 60.200 162.595 60.455 162.755 ;
        RECT 60.635 162.415 60.920 162.875 ;
        RECT 61.100 162.675 61.350 163.325 ;
        RECT 61.550 164.075 61.870 164.095 ;
        RECT 61.550 163.905 63.470 164.075 ;
        RECT 61.550 163.010 61.740 163.905 ;
        RECT 63.640 163.735 63.810 164.245 ;
        RECT 63.980 163.985 64.500 164.295 ;
        RECT 61.910 163.565 63.810 163.735 ;
        RECT 61.910 163.505 62.240 163.565 ;
        RECT 62.390 163.335 62.720 163.395 ;
        RECT 62.060 163.065 62.720 163.335 ;
        RECT 61.550 162.680 61.870 163.010 ;
        RECT 62.050 162.415 62.710 162.895 ;
        RECT 62.910 162.805 63.080 163.565 ;
        RECT 63.980 163.395 64.160 163.805 ;
        RECT 63.250 163.225 63.580 163.345 ;
        RECT 64.330 163.225 64.500 163.985 ;
        RECT 63.250 163.055 64.500 163.225 ;
        RECT 64.670 164.165 66.040 164.415 ;
        RECT 64.670 163.395 64.860 164.165 ;
        RECT 65.790 163.905 66.040 164.165 ;
        RECT 65.030 163.735 65.280 163.895 ;
        RECT 66.210 163.735 66.380 164.580 ;
        RECT 67.275 164.295 67.445 164.795 ;
        RECT 67.615 164.465 67.945 164.965 ;
        RECT 66.550 163.905 67.050 164.285 ;
        RECT 67.275 164.125 67.970 164.295 ;
        RECT 65.030 163.565 66.380 163.735 ;
        RECT 65.960 163.525 66.380 163.565 ;
        RECT 64.670 163.055 65.090 163.395 ;
        RECT 65.380 163.065 65.790 163.395 ;
        RECT 62.910 162.635 63.760 162.805 ;
        RECT 64.320 162.415 64.640 162.875 ;
        RECT 64.840 162.625 65.090 163.055 ;
        RECT 65.380 162.415 65.790 162.855 ;
        RECT 65.960 162.795 66.130 163.525 ;
        RECT 66.300 162.975 66.650 163.345 ;
        RECT 66.830 163.035 67.050 163.905 ;
        RECT 67.220 163.335 67.630 163.955 ;
        RECT 67.800 163.155 67.970 164.125 ;
        RECT 67.275 162.965 67.970 163.155 ;
        RECT 65.960 162.595 66.975 162.795 ;
        RECT 67.275 162.635 67.445 162.965 ;
        RECT 67.615 162.415 67.945 162.795 ;
        RECT 68.160 162.675 68.385 164.795 ;
        RECT 68.555 164.465 68.885 164.965 ;
        RECT 69.055 164.295 69.225 164.795 ;
        RECT 68.560 164.125 69.225 164.295 ;
        RECT 68.560 163.135 68.790 164.125 ;
        RECT 68.960 163.305 69.310 163.955 ;
        RECT 70.405 163.875 73.915 164.965 ;
        RECT 70.405 163.355 72.095 163.875 ;
        RECT 74.090 163.815 74.350 164.965 ;
        RECT 74.525 163.890 74.780 164.795 ;
        RECT 74.950 164.205 75.280 164.965 ;
        RECT 75.495 164.035 75.665 164.795 ;
        RECT 72.265 163.185 73.915 163.705 ;
        RECT 68.560 162.965 69.225 163.135 ;
        RECT 68.555 162.415 68.885 162.795 ;
        RECT 69.055 162.675 69.225 162.965 ;
        RECT 70.405 162.415 73.915 163.185 ;
        RECT 74.090 162.415 74.350 163.255 ;
        RECT 74.525 163.160 74.695 163.890 ;
        RECT 74.950 163.865 75.665 164.035 ;
        RECT 74.950 163.655 75.120 163.865 ;
        RECT 75.925 163.800 76.215 164.965 ;
        RECT 76.385 163.875 78.975 164.965 ;
        RECT 74.865 163.325 75.120 163.655 ;
        RECT 74.525 162.585 74.780 163.160 ;
        RECT 74.950 163.135 75.120 163.325 ;
        RECT 75.400 163.315 75.755 163.685 ;
        RECT 76.385 163.355 77.595 163.875 ;
        RECT 79.145 163.825 79.485 164.795 ;
        RECT 79.655 163.825 79.825 164.965 ;
        RECT 80.095 164.165 80.345 164.965 ;
        RECT 80.990 163.995 81.320 164.795 ;
        RECT 81.620 164.165 81.950 164.965 ;
        RECT 82.120 163.995 82.450 164.795 ;
        RECT 80.015 163.825 82.450 163.995 ;
        RECT 83.660 163.985 83.915 164.655 ;
        RECT 84.095 164.165 84.380 164.965 ;
        RECT 84.560 164.245 84.890 164.755 ;
        RECT 83.660 163.945 83.840 163.985 ;
        RECT 77.765 163.185 78.975 163.705 ;
        RECT 74.950 162.965 75.665 163.135 ;
        RECT 74.950 162.415 75.280 162.795 ;
        RECT 75.495 162.585 75.665 162.965 ;
        RECT 75.925 162.415 76.215 163.140 ;
        RECT 76.385 162.415 78.975 163.185 ;
        RECT 79.145 163.215 79.320 163.825 ;
        RECT 80.015 163.575 80.185 163.825 ;
        RECT 79.490 163.405 80.185 163.575 ;
        RECT 80.360 163.405 80.780 163.605 ;
        RECT 80.950 163.405 81.280 163.605 ;
        RECT 81.450 163.405 81.780 163.605 ;
        RECT 79.145 162.585 79.485 163.215 ;
        RECT 79.655 162.415 79.905 163.215 ;
        RECT 80.095 163.065 81.320 163.235 ;
        RECT 80.095 162.585 80.425 163.065 ;
        RECT 80.595 162.415 80.820 162.875 ;
        RECT 80.990 162.585 81.320 163.065 ;
        RECT 81.950 163.195 82.120 163.825 ;
        RECT 83.575 163.775 83.840 163.945 ;
        RECT 82.305 163.405 82.655 163.655 ;
        RECT 81.950 162.585 82.450 163.195 ;
        RECT 83.660 163.125 83.840 163.775 ;
        RECT 84.560 163.655 84.810 164.245 ;
        RECT 85.160 164.095 85.330 164.705 ;
        RECT 85.500 164.275 85.830 164.965 ;
        RECT 86.060 164.415 86.300 164.705 ;
        RECT 86.500 164.585 86.920 164.965 ;
        RECT 87.100 164.495 87.730 164.745 ;
        RECT 88.200 164.585 88.530 164.965 ;
        RECT 87.100 164.415 87.270 164.495 ;
        RECT 88.700 164.415 88.870 164.705 ;
        RECT 89.050 164.585 89.430 164.965 ;
        RECT 89.670 164.580 90.500 164.750 ;
        RECT 86.060 164.245 87.270 164.415 ;
        RECT 84.010 163.325 84.810 163.655 ;
        RECT 83.660 162.595 83.915 163.125 ;
        RECT 84.095 162.415 84.380 162.875 ;
        RECT 84.560 162.675 84.810 163.325 ;
        RECT 85.010 164.075 85.330 164.095 ;
        RECT 85.010 163.905 86.930 164.075 ;
        RECT 85.010 163.010 85.200 163.905 ;
        RECT 87.100 163.735 87.270 164.245 ;
        RECT 87.440 163.985 87.960 164.295 ;
        RECT 85.370 163.565 87.270 163.735 ;
        RECT 85.370 163.505 85.700 163.565 ;
        RECT 85.850 163.335 86.180 163.395 ;
        RECT 85.520 163.065 86.180 163.335 ;
        RECT 85.010 162.680 85.330 163.010 ;
        RECT 85.510 162.415 86.170 162.895 ;
        RECT 86.370 162.805 86.540 163.565 ;
        RECT 87.440 163.395 87.620 163.805 ;
        RECT 86.710 163.225 87.040 163.345 ;
        RECT 87.790 163.225 87.960 163.985 ;
        RECT 86.710 163.055 87.960 163.225 ;
        RECT 88.130 164.165 89.500 164.415 ;
        RECT 88.130 163.395 88.320 164.165 ;
        RECT 89.250 163.905 89.500 164.165 ;
        RECT 88.490 163.735 88.740 163.895 ;
        RECT 89.670 163.735 89.840 164.580 ;
        RECT 90.735 164.295 90.905 164.795 ;
        RECT 91.075 164.465 91.405 164.965 ;
        RECT 90.010 163.905 90.510 164.285 ;
        RECT 90.735 164.125 91.430 164.295 ;
        RECT 88.490 163.565 89.840 163.735 ;
        RECT 89.420 163.525 89.840 163.565 ;
        RECT 88.130 163.055 88.550 163.395 ;
        RECT 88.840 163.065 89.250 163.395 ;
        RECT 86.370 162.635 87.220 162.805 ;
        RECT 87.780 162.415 88.100 162.875 ;
        RECT 88.300 162.625 88.550 163.055 ;
        RECT 88.840 162.415 89.250 162.855 ;
        RECT 89.420 162.795 89.590 163.525 ;
        RECT 89.760 162.975 90.110 163.345 ;
        RECT 90.290 163.035 90.510 163.905 ;
        RECT 90.680 163.335 91.090 163.955 ;
        RECT 91.260 163.155 91.430 164.125 ;
        RECT 90.735 162.965 91.430 163.155 ;
        RECT 89.420 162.595 90.435 162.795 ;
        RECT 90.735 162.635 90.905 162.965 ;
        RECT 91.075 162.415 91.405 162.795 ;
        RECT 91.620 162.675 91.845 164.795 ;
        RECT 92.015 164.465 92.345 164.965 ;
        RECT 92.515 164.295 92.685 164.795 ;
        RECT 92.020 164.125 92.685 164.295 ;
        RECT 92.020 163.135 92.250 164.125 ;
        RECT 92.420 163.305 92.770 163.955 ;
        RECT 92.950 163.825 93.285 164.795 ;
        RECT 93.455 163.825 93.625 164.965 ;
        RECT 93.795 164.625 95.825 164.795 ;
        RECT 92.950 163.155 93.120 163.825 ;
        RECT 93.795 163.655 93.965 164.625 ;
        RECT 93.290 163.325 93.545 163.655 ;
        RECT 93.770 163.325 93.965 163.655 ;
        RECT 94.135 164.285 95.260 164.455 ;
        RECT 93.375 163.155 93.545 163.325 ;
        RECT 94.135 163.155 94.305 164.285 ;
        RECT 92.020 162.965 92.685 163.135 ;
        RECT 92.015 162.415 92.345 162.795 ;
        RECT 92.515 162.675 92.685 162.965 ;
        RECT 92.950 162.585 93.205 163.155 ;
        RECT 93.375 162.985 94.305 163.155 ;
        RECT 94.475 163.945 95.485 164.115 ;
        RECT 94.475 163.145 94.645 163.945 ;
        RECT 94.850 163.605 95.125 163.745 ;
        RECT 94.845 163.435 95.125 163.605 ;
        RECT 94.130 162.950 94.305 162.985 ;
        RECT 93.375 162.415 93.705 162.815 ;
        RECT 94.130 162.585 94.660 162.950 ;
        RECT 94.850 162.585 95.125 163.435 ;
        RECT 95.295 162.585 95.485 163.945 ;
        RECT 95.655 163.960 95.825 164.625 ;
        RECT 95.995 164.205 96.165 164.965 ;
        RECT 96.400 164.205 96.915 164.615 ;
        RECT 95.655 163.770 96.405 163.960 ;
        RECT 96.575 163.395 96.915 164.205 ;
        RECT 95.685 163.225 96.915 163.395 ;
        RECT 98.005 163.825 98.345 164.795 ;
        RECT 98.515 163.825 98.685 164.965 ;
        RECT 98.955 164.165 99.205 164.965 ;
        RECT 99.850 163.995 100.180 164.795 ;
        RECT 100.480 164.165 100.810 164.965 ;
        RECT 100.980 163.995 101.310 164.795 ;
        RECT 98.875 163.825 101.310 163.995 ;
        RECT 95.665 162.415 96.175 162.950 ;
        RECT 96.395 162.620 96.640 163.225 ;
        RECT 98.005 163.215 98.180 163.825 ;
        RECT 98.875 163.575 99.045 163.825 ;
        RECT 98.350 163.405 99.045 163.575 ;
        RECT 99.220 163.405 99.640 163.605 ;
        RECT 99.810 163.405 100.140 163.605 ;
        RECT 100.310 163.405 100.640 163.605 ;
        RECT 98.005 162.585 98.345 163.215 ;
        RECT 98.515 162.415 98.765 163.215 ;
        RECT 98.955 163.065 100.180 163.235 ;
        RECT 98.955 162.585 99.285 163.065 ;
        RECT 99.455 162.415 99.680 162.875 ;
        RECT 99.850 162.585 100.180 163.065 ;
        RECT 100.810 163.195 100.980 163.825 ;
        RECT 101.685 163.800 101.975 164.965 ;
        RECT 102.610 164.530 107.955 164.965 ;
        RECT 101.165 163.405 101.515 163.655 ;
        RECT 104.200 163.280 104.550 164.530 ;
        RECT 108.125 163.825 108.465 164.795 ;
        RECT 108.635 163.825 108.805 164.965 ;
        RECT 109.075 164.165 109.325 164.965 ;
        RECT 109.970 163.995 110.300 164.795 ;
        RECT 110.600 164.165 110.930 164.965 ;
        RECT 111.100 163.995 111.430 164.795 ;
        RECT 108.995 163.825 111.430 163.995 ;
        RECT 111.805 163.825 112.145 164.795 ;
        RECT 112.315 163.825 112.485 164.965 ;
        RECT 112.755 164.165 113.005 164.965 ;
        RECT 113.650 163.995 113.980 164.795 ;
        RECT 114.280 164.165 114.610 164.965 ;
        RECT 114.780 163.995 115.110 164.795 ;
        RECT 115.490 164.530 120.835 164.965 ;
        RECT 121.010 164.530 126.355 164.965 ;
        RECT 112.675 163.825 115.110 163.995 ;
        RECT 100.810 162.585 101.310 163.195 ;
        RECT 101.685 162.415 101.975 163.140 ;
        RECT 106.030 162.960 106.370 163.790 ;
        RECT 108.125 163.215 108.300 163.825 ;
        RECT 108.995 163.575 109.165 163.825 ;
        RECT 108.470 163.405 109.165 163.575 ;
        RECT 109.340 163.405 109.760 163.605 ;
        RECT 109.930 163.405 110.260 163.605 ;
        RECT 110.430 163.405 110.760 163.605 ;
        RECT 102.610 162.415 107.955 162.960 ;
        RECT 108.125 162.585 108.465 163.215 ;
        RECT 108.635 162.415 108.885 163.215 ;
        RECT 109.075 163.065 110.300 163.235 ;
        RECT 109.075 162.585 109.405 163.065 ;
        RECT 109.575 162.415 109.800 162.875 ;
        RECT 109.970 162.585 110.300 163.065 ;
        RECT 110.930 163.195 111.100 163.825 ;
        RECT 111.285 163.405 111.635 163.655 ;
        RECT 111.805 163.215 111.980 163.825 ;
        RECT 112.675 163.575 112.845 163.825 ;
        RECT 112.150 163.405 112.845 163.575 ;
        RECT 113.020 163.405 113.440 163.605 ;
        RECT 113.610 163.405 113.940 163.605 ;
        RECT 114.110 163.405 114.440 163.605 ;
        RECT 110.930 162.585 111.430 163.195 ;
        RECT 111.805 162.585 112.145 163.215 ;
        RECT 112.315 162.415 112.565 163.215 ;
        RECT 112.755 163.065 113.980 163.235 ;
        RECT 112.755 162.585 113.085 163.065 ;
        RECT 113.255 162.415 113.480 162.875 ;
        RECT 113.650 162.585 113.980 163.065 ;
        RECT 114.610 163.195 114.780 163.825 ;
        RECT 114.965 163.405 115.315 163.655 ;
        RECT 117.080 163.280 117.430 164.530 ;
        RECT 114.610 162.585 115.110 163.195 ;
        RECT 118.910 162.960 119.250 163.790 ;
        RECT 122.600 163.280 122.950 164.530 ;
        RECT 126.525 163.875 127.735 164.965 ;
        RECT 124.430 162.960 124.770 163.790 ;
        RECT 126.525 163.335 127.045 163.875 ;
        RECT 127.215 163.165 127.735 163.705 ;
        RECT 115.490 162.415 120.835 162.960 ;
        RECT 121.010 162.415 126.355 162.960 ;
        RECT 126.525 162.415 127.735 163.165 ;
        RECT 14.660 162.245 127.820 162.415 ;
        RECT 14.745 161.495 15.955 162.245 ;
        RECT 17.050 161.535 17.305 162.065 ;
        RECT 17.475 161.785 17.780 162.245 ;
        RECT 18.025 161.865 19.095 162.035 ;
        RECT 14.745 160.955 15.265 161.495 ;
        RECT 15.435 160.785 15.955 161.325 ;
        RECT 14.745 159.695 15.955 160.785 ;
        RECT 17.050 160.885 17.260 161.535 ;
        RECT 18.025 161.510 18.345 161.865 ;
        RECT 18.020 161.335 18.345 161.510 ;
        RECT 17.430 161.035 18.345 161.335 ;
        RECT 18.515 161.295 18.755 161.695 ;
        RECT 18.925 161.635 19.095 161.865 ;
        RECT 19.265 161.805 19.455 162.245 ;
        RECT 19.625 161.795 20.575 162.075 ;
        RECT 20.795 161.885 21.145 162.055 ;
        RECT 18.925 161.465 19.455 161.635 ;
        RECT 17.430 161.005 18.170 161.035 ;
        RECT 17.050 160.005 17.305 160.885 ;
        RECT 17.475 159.695 17.780 160.835 ;
        RECT 18.000 160.415 18.170 161.005 ;
        RECT 18.515 160.925 19.055 161.295 ;
        RECT 19.235 161.185 19.455 161.465 ;
        RECT 19.625 161.015 19.795 161.795 ;
        RECT 19.390 160.845 19.795 161.015 ;
        RECT 19.965 161.005 20.315 161.625 ;
        RECT 19.390 160.755 19.560 160.845 ;
        RECT 20.485 160.835 20.695 161.625 ;
        RECT 18.340 160.585 19.560 160.755 ;
        RECT 20.020 160.675 20.695 160.835 ;
        RECT 18.000 160.245 18.800 160.415 ;
        RECT 18.120 159.695 18.450 160.075 ;
        RECT 18.630 159.955 18.800 160.245 ;
        RECT 19.390 160.205 19.560 160.585 ;
        RECT 19.730 160.665 20.695 160.675 ;
        RECT 20.885 161.495 21.145 161.885 ;
        RECT 21.355 161.785 21.685 162.245 ;
        RECT 22.560 161.855 23.415 162.025 ;
        RECT 23.620 161.855 24.115 162.025 ;
        RECT 24.285 161.885 24.615 162.245 ;
        RECT 20.885 160.805 21.055 161.495 ;
        RECT 21.225 161.145 21.395 161.325 ;
        RECT 21.565 161.315 22.355 161.565 ;
        RECT 22.560 161.145 22.730 161.855 ;
        RECT 22.900 161.345 23.255 161.565 ;
        RECT 21.225 160.975 22.915 161.145 ;
        RECT 19.730 160.375 20.190 160.665 ;
        RECT 20.885 160.635 22.385 160.805 ;
        RECT 20.885 160.495 21.055 160.635 ;
        RECT 20.495 160.325 21.055 160.495 ;
        RECT 18.970 159.695 19.220 160.155 ;
        RECT 19.390 159.865 20.260 160.205 ;
        RECT 20.495 159.865 20.665 160.325 ;
        RECT 21.500 160.295 22.575 160.465 ;
        RECT 20.835 159.695 21.205 160.155 ;
        RECT 21.500 159.955 21.670 160.295 ;
        RECT 21.840 159.695 22.170 160.125 ;
        RECT 22.405 159.955 22.575 160.295 ;
        RECT 22.745 160.195 22.915 160.975 ;
        RECT 23.085 160.755 23.255 161.345 ;
        RECT 23.425 160.945 23.775 161.565 ;
        RECT 23.085 160.365 23.550 160.755 ;
        RECT 23.945 160.495 24.115 161.855 ;
        RECT 24.285 160.665 24.745 161.715 ;
        RECT 23.720 160.325 24.115 160.495 ;
        RECT 23.720 160.195 23.890 160.325 ;
        RECT 22.745 159.865 23.425 160.195 ;
        RECT 23.640 159.865 23.890 160.195 ;
        RECT 24.060 159.695 24.310 160.155 ;
        RECT 24.480 159.880 24.805 160.665 ;
        RECT 24.975 159.865 25.145 161.985 ;
        RECT 25.315 161.865 25.645 162.245 ;
        RECT 25.815 161.695 26.070 161.985 ;
        RECT 26.335 161.765 26.635 162.245 ;
        RECT 25.320 161.525 26.070 161.695 ;
        RECT 26.805 161.595 27.065 162.050 ;
        RECT 27.235 161.765 27.495 162.245 ;
        RECT 27.675 161.595 27.935 162.050 ;
        RECT 28.105 161.765 28.355 162.245 ;
        RECT 28.535 161.595 28.795 162.050 ;
        RECT 28.965 161.765 29.215 162.245 ;
        RECT 29.395 161.595 29.655 162.050 ;
        RECT 29.825 161.765 30.070 162.245 ;
        RECT 30.240 161.595 30.515 162.050 ;
        RECT 30.685 161.765 30.930 162.245 ;
        RECT 31.100 161.595 31.360 162.050 ;
        RECT 31.530 161.765 31.790 162.245 ;
        RECT 31.960 161.595 32.220 162.050 ;
        RECT 32.390 161.765 32.650 162.245 ;
        RECT 32.820 161.595 33.080 162.050 ;
        RECT 33.250 161.685 33.510 162.245 ;
        RECT 25.320 160.535 25.550 161.525 ;
        RECT 26.335 161.425 33.080 161.595 ;
        RECT 25.720 160.705 26.070 161.355 ;
        RECT 26.335 160.835 27.500 161.425 ;
        RECT 33.680 161.255 33.930 162.065 ;
        RECT 34.110 161.720 34.370 162.245 ;
        RECT 34.540 161.255 34.790 162.065 ;
        RECT 34.970 161.735 35.275 162.245 ;
        RECT 35.450 161.775 35.780 162.245 ;
        RECT 35.950 161.605 36.175 162.050 ;
        RECT 36.345 161.720 36.640 162.245 ;
        RECT 27.670 161.005 34.790 161.255 ;
        RECT 34.960 161.005 35.275 161.565 ;
        RECT 35.445 161.435 36.175 161.605 ;
        RECT 37.285 161.520 37.575 162.245 ;
        RECT 37.750 161.505 38.005 162.075 ;
        RECT 38.175 161.845 38.505 162.245 ;
        RECT 38.930 161.710 39.460 162.075 ;
        RECT 39.650 161.905 39.925 162.075 ;
        RECT 39.645 161.735 39.925 161.905 ;
        RECT 38.930 161.675 39.105 161.710 ;
        RECT 38.175 161.505 39.105 161.675 ;
        RECT 26.335 160.610 33.080 160.835 ;
        RECT 25.320 160.365 26.070 160.535 ;
        RECT 25.315 159.695 25.645 160.195 ;
        RECT 25.815 159.865 26.070 160.365 ;
        RECT 26.335 159.695 26.605 160.440 ;
        RECT 26.775 159.870 27.065 160.610 ;
        RECT 27.675 160.595 33.080 160.610 ;
        RECT 27.235 159.700 27.490 160.425 ;
        RECT 27.675 159.870 27.935 160.595 ;
        RECT 28.105 159.700 28.350 160.425 ;
        RECT 28.535 159.870 28.795 160.595 ;
        RECT 28.965 159.700 29.210 160.425 ;
        RECT 29.395 159.870 29.655 160.595 ;
        RECT 29.825 159.700 30.070 160.425 ;
        RECT 30.240 159.870 30.500 160.595 ;
        RECT 30.670 159.700 30.930 160.425 ;
        RECT 31.100 159.870 31.360 160.595 ;
        RECT 31.530 159.700 31.790 160.425 ;
        RECT 31.960 159.870 32.220 160.595 ;
        RECT 32.390 159.700 32.650 160.425 ;
        RECT 32.820 159.870 33.080 160.595 ;
        RECT 33.250 159.700 33.510 160.495 ;
        RECT 33.680 159.870 33.930 161.005 ;
        RECT 27.235 159.695 33.510 159.700 ;
        RECT 34.110 159.695 34.370 160.505 ;
        RECT 34.545 159.865 34.790 161.005 ;
        RECT 35.445 160.870 35.725 161.435 ;
        RECT 35.895 161.040 37.115 161.265 ;
        RECT 35.445 160.700 37.045 160.870 ;
        RECT 34.970 159.695 35.265 160.505 ;
        RECT 35.505 159.695 35.760 160.530 ;
        RECT 35.930 159.895 36.190 160.700 ;
        RECT 36.360 159.695 36.620 160.530 ;
        RECT 36.790 159.895 37.045 160.700 ;
        RECT 37.285 159.695 37.575 160.860 ;
        RECT 37.750 160.835 37.920 161.505 ;
        RECT 38.175 161.335 38.345 161.505 ;
        RECT 38.090 161.005 38.345 161.335 ;
        RECT 38.570 161.005 38.765 161.335 ;
        RECT 37.750 159.865 38.085 160.835 ;
        RECT 38.255 159.695 38.425 160.835 ;
        RECT 38.595 160.035 38.765 161.005 ;
        RECT 38.935 160.375 39.105 161.505 ;
        RECT 39.275 160.715 39.445 161.515 ;
        RECT 39.650 160.915 39.925 161.735 ;
        RECT 40.095 160.715 40.285 162.075 ;
        RECT 40.465 161.710 40.975 162.245 ;
        RECT 41.195 161.435 41.440 162.040 ;
        RECT 42.810 161.700 48.155 162.245 ;
        RECT 40.485 161.265 41.715 161.435 ;
        RECT 39.275 160.545 40.285 160.715 ;
        RECT 40.455 160.700 41.205 160.890 ;
        RECT 38.935 160.205 40.060 160.375 ;
        RECT 40.455 160.035 40.625 160.700 ;
        RECT 41.375 160.455 41.715 161.265 ;
        RECT 38.595 159.865 40.625 160.035 ;
        RECT 40.795 159.695 40.965 160.455 ;
        RECT 41.200 160.045 41.715 160.455 ;
        RECT 44.400 160.130 44.750 161.380 ;
        RECT 46.230 160.870 46.570 161.700 ;
        RECT 48.325 161.445 48.665 162.075 ;
        RECT 48.835 161.445 49.085 162.245 ;
        RECT 49.275 161.595 49.605 162.075 ;
        RECT 49.775 161.785 50.000 162.245 ;
        RECT 50.170 161.595 50.500 162.075 ;
        RECT 48.325 160.835 48.500 161.445 ;
        RECT 49.275 161.425 50.500 161.595 ;
        RECT 51.130 161.465 51.630 162.075 ;
        RECT 52.010 161.700 57.355 162.245 ;
        RECT 48.670 161.085 49.365 161.255 ;
        RECT 49.195 160.835 49.365 161.085 ;
        RECT 49.540 161.055 49.960 161.255 ;
        RECT 50.130 161.055 50.460 161.255 ;
        RECT 50.630 161.055 50.960 161.255 ;
        RECT 51.130 160.835 51.300 161.465 ;
        RECT 51.485 161.005 51.835 161.255 ;
        RECT 42.810 159.695 48.155 160.130 ;
        RECT 48.325 159.865 48.665 160.835 ;
        RECT 48.835 159.695 49.005 160.835 ;
        RECT 49.195 160.665 51.630 160.835 ;
        RECT 49.275 159.695 49.525 160.495 ;
        RECT 50.170 159.865 50.500 160.665 ;
        RECT 50.800 159.695 51.130 160.495 ;
        RECT 51.300 159.865 51.630 160.665 ;
        RECT 53.600 160.130 53.950 161.380 ;
        RECT 55.430 160.870 55.770 161.700 ;
        RECT 57.585 161.425 57.795 162.245 ;
        RECT 57.965 161.445 58.295 162.075 ;
        RECT 57.965 160.845 58.215 161.445 ;
        RECT 58.465 161.425 58.695 162.245 ;
        RECT 59.180 161.435 59.425 162.040 ;
        RECT 59.645 161.710 60.155 162.245 ;
        RECT 58.905 161.265 60.135 161.435 ;
        RECT 58.385 161.005 58.715 161.255 ;
        RECT 52.010 159.695 57.355 160.130 ;
        RECT 57.585 159.695 57.795 160.835 ;
        RECT 57.965 159.865 58.295 160.845 ;
        RECT 58.465 159.695 58.695 160.835 ;
        RECT 58.905 160.455 59.245 161.265 ;
        RECT 59.415 160.700 60.165 160.890 ;
        RECT 58.905 160.045 59.420 160.455 ;
        RECT 59.655 159.695 59.825 160.455 ;
        RECT 59.995 160.035 60.165 160.700 ;
        RECT 60.335 160.715 60.525 162.075 ;
        RECT 60.695 161.225 60.970 162.075 ;
        RECT 61.160 161.710 61.690 162.075 ;
        RECT 62.115 161.845 62.445 162.245 ;
        RECT 61.515 161.675 61.690 161.710 ;
        RECT 60.695 161.055 60.975 161.225 ;
        RECT 60.695 160.915 60.970 161.055 ;
        RECT 61.175 160.715 61.345 161.515 ;
        RECT 60.335 160.545 61.345 160.715 ;
        RECT 61.515 161.505 62.445 161.675 ;
        RECT 62.615 161.505 62.870 162.075 ;
        RECT 63.045 161.520 63.335 162.245 ;
        RECT 64.055 161.695 64.225 162.075 ;
        RECT 64.405 161.865 64.735 162.245 ;
        RECT 64.055 161.525 64.720 161.695 ;
        RECT 64.915 161.570 65.175 162.075 ;
        RECT 61.515 160.375 61.685 161.505 ;
        RECT 62.275 161.335 62.445 161.505 ;
        RECT 60.560 160.205 61.685 160.375 ;
        RECT 61.855 161.005 62.050 161.335 ;
        RECT 62.275 161.005 62.530 161.335 ;
        RECT 61.855 160.035 62.025 161.005 ;
        RECT 62.700 160.835 62.870 161.505 ;
        RECT 63.985 160.975 64.315 161.345 ;
        RECT 64.550 161.270 64.720 161.525 ;
        RECT 64.550 160.940 64.835 161.270 ;
        RECT 59.995 159.865 62.025 160.035 ;
        RECT 62.195 159.695 62.365 160.835 ;
        RECT 62.535 159.865 62.870 160.835 ;
        RECT 63.045 159.695 63.335 160.860 ;
        RECT 64.550 160.795 64.720 160.940 ;
        RECT 64.055 160.625 64.720 160.795 ;
        RECT 65.005 160.770 65.175 161.570 ;
        RECT 64.055 159.865 64.225 160.625 ;
        RECT 64.405 159.695 64.735 160.455 ;
        RECT 64.905 159.865 65.175 160.770 ;
        RECT 65.345 161.745 65.605 162.075 ;
        RECT 65.775 161.885 66.105 162.245 ;
        RECT 66.360 161.865 67.660 162.075 ;
        RECT 65.345 160.545 65.515 161.745 ;
        RECT 66.360 161.715 66.530 161.865 ;
        RECT 65.775 161.590 66.530 161.715 ;
        RECT 65.685 161.545 66.530 161.590 ;
        RECT 65.685 161.425 65.955 161.545 ;
        RECT 65.685 160.850 65.855 161.425 ;
        RECT 66.085 160.985 66.495 161.290 ;
        RECT 66.785 161.255 66.995 161.655 ;
        RECT 66.665 161.045 66.995 161.255 ;
        RECT 67.240 161.255 67.460 161.655 ;
        RECT 67.935 161.480 68.390 162.245 ;
        RECT 69.485 161.475 72.995 162.245 ;
        RECT 67.240 161.045 67.715 161.255 ;
        RECT 67.905 161.055 68.395 161.255 ;
        RECT 65.685 160.815 65.885 160.850 ;
        RECT 67.215 160.815 68.390 160.875 ;
        RECT 65.685 160.705 68.390 160.815 ;
        RECT 65.745 160.645 67.545 160.705 ;
        RECT 67.215 160.615 67.545 160.645 ;
        RECT 65.345 159.865 65.605 160.545 ;
        RECT 65.775 159.695 66.025 160.475 ;
        RECT 66.275 160.445 67.110 160.455 ;
        RECT 67.700 160.445 67.885 160.535 ;
        RECT 66.275 160.245 67.885 160.445 ;
        RECT 66.275 159.865 66.525 160.245 ;
        RECT 67.655 160.205 67.885 160.245 ;
        RECT 68.135 160.085 68.390 160.705 ;
        RECT 66.695 159.695 67.050 160.075 ;
        RECT 68.055 159.865 68.390 160.085 ;
        RECT 69.485 160.785 71.175 161.305 ;
        RECT 71.345 160.955 72.995 161.475 ;
        RECT 73.170 161.405 73.430 162.245 ;
        RECT 73.605 161.500 73.860 162.075 ;
        RECT 74.030 161.865 74.360 162.245 ;
        RECT 74.575 161.695 74.745 162.075 ;
        RECT 74.030 161.525 74.745 161.695 ;
        RECT 69.485 159.695 72.995 160.785 ;
        RECT 73.170 159.695 73.430 160.845 ;
        RECT 73.605 160.770 73.775 161.500 ;
        RECT 74.030 161.335 74.200 161.525 ;
        RECT 75.005 161.495 76.215 162.245 ;
        RECT 73.945 161.005 74.200 161.335 ;
        RECT 74.030 160.795 74.200 161.005 ;
        RECT 74.480 160.975 74.835 161.345 ;
        RECT 73.605 159.865 73.860 160.770 ;
        RECT 74.030 160.625 74.745 160.795 ;
        RECT 74.030 159.695 74.360 160.455 ;
        RECT 74.575 159.865 74.745 160.625 ;
        RECT 75.005 160.785 75.525 161.325 ;
        RECT 75.695 160.955 76.215 161.495 ;
        RECT 76.385 161.475 79.895 162.245 ;
        RECT 76.385 160.785 78.075 161.305 ;
        RECT 78.245 160.955 79.895 161.475 ;
        RECT 80.270 161.465 80.770 162.075 ;
        RECT 80.065 161.005 80.415 161.255 ;
        RECT 80.600 160.835 80.770 161.465 ;
        RECT 81.400 161.595 81.730 162.075 ;
        RECT 81.900 161.785 82.125 162.245 ;
        RECT 82.295 161.595 82.625 162.075 ;
        RECT 81.400 161.425 82.625 161.595 ;
        RECT 82.815 161.445 83.065 162.245 ;
        RECT 83.235 161.445 83.575 162.075 ;
        RECT 84.755 161.695 84.925 162.075 ;
        RECT 85.105 161.865 85.435 162.245 ;
        RECT 84.755 161.525 85.420 161.695 ;
        RECT 85.615 161.570 85.875 162.075 ;
        RECT 80.940 161.055 81.270 161.255 ;
        RECT 81.440 161.055 81.770 161.255 ;
        RECT 81.940 161.055 82.360 161.255 ;
        RECT 82.535 161.085 83.230 161.255 ;
        RECT 82.535 160.835 82.705 161.085 ;
        RECT 83.400 160.885 83.575 161.445 ;
        RECT 84.685 160.975 85.015 161.345 ;
        RECT 85.250 161.270 85.420 161.525 ;
        RECT 83.345 160.835 83.575 160.885 ;
        RECT 75.005 159.695 76.215 160.785 ;
        RECT 76.385 159.695 79.895 160.785 ;
        RECT 80.270 160.665 82.705 160.835 ;
        RECT 80.270 159.865 80.600 160.665 ;
        RECT 80.770 159.695 81.100 160.495 ;
        RECT 81.400 159.865 81.730 160.665 ;
        RECT 82.375 159.695 82.625 160.495 ;
        RECT 82.895 159.695 83.065 160.835 ;
        RECT 83.235 159.865 83.575 160.835 ;
        RECT 85.250 160.940 85.535 161.270 ;
        RECT 85.250 160.795 85.420 160.940 ;
        RECT 84.755 160.625 85.420 160.795 ;
        RECT 85.705 160.770 85.875 161.570 ;
        RECT 86.105 161.425 86.315 162.245 ;
        RECT 86.485 161.445 86.815 162.075 ;
        RECT 86.485 160.845 86.735 161.445 ;
        RECT 86.985 161.425 87.215 162.245 ;
        RECT 87.465 161.425 87.695 162.245 ;
        RECT 87.865 161.445 88.195 162.075 ;
        RECT 86.905 161.005 87.235 161.255 ;
        RECT 87.445 161.005 87.775 161.255 ;
        RECT 87.945 160.845 88.195 161.445 ;
        RECT 88.365 161.425 88.575 162.245 ;
        RECT 88.805 161.520 89.095 162.245 ;
        RECT 89.640 161.535 89.895 162.065 ;
        RECT 90.075 161.785 90.360 162.245 ;
        RECT 84.755 159.865 84.925 160.625 ;
        RECT 85.105 159.695 85.435 160.455 ;
        RECT 85.605 159.865 85.875 160.770 ;
        RECT 86.105 159.695 86.315 160.835 ;
        RECT 86.485 159.865 86.815 160.845 ;
        RECT 86.985 159.695 87.215 160.835 ;
        RECT 87.465 159.695 87.695 160.835 ;
        RECT 87.865 159.865 88.195 160.845 ;
        RECT 88.365 159.695 88.575 160.835 ;
        RECT 88.805 159.695 89.095 160.860 ;
        RECT 89.640 160.675 89.820 161.535 ;
        RECT 90.540 161.335 90.790 161.985 ;
        RECT 89.990 161.005 90.790 161.335 ;
        RECT 89.640 160.545 89.895 160.675 ;
        RECT 89.555 160.375 89.895 160.545 ;
        RECT 89.640 160.005 89.895 160.375 ;
        RECT 90.075 159.695 90.360 160.495 ;
        RECT 90.540 160.415 90.790 161.005 ;
        RECT 90.990 161.650 91.310 161.980 ;
        RECT 91.490 161.765 92.150 162.245 ;
        RECT 92.350 161.855 93.200 162.025 ;
        RECT 90.990 160.755 91.180 161.650 ;
        RECT 91.500 161.325 92.160 161.595 ;
        RECT 91.830 161.265 92.160 161.325 ;
        RECT 91.350 161.095 91.680 161.155 ;
        RECT 92.350 161.095 92.520 161.855 ;
        RECT 93.760 161.785 94.080 162.245 ;
        RECT 94.280 161.605 94.530 162.035 ;
        RECT 94.820 161.805 95.230 162.245 ;
        RECT 95.400 161.865 96.415 162.065 ;
        RECT 92.690 161.435 93.940 161.605 ;
        RECT 92.690 161.315 93.020 161.435 ;
        RECT 91.350 160.925 93.250 161.095 ;
        RECT 90.990 160.585 92.910 160.755 ;
        RECT 90.990 160.565 91.310 160.585 ;
        RECT 90.540 159.905 90.870 160.415 ;
        RECT 91.140 159.955 91.310 160.565 ;
        RECT 93.080 160.415 93.250 160.925 ;
        RECT 93.420 160.855 93.600 161.265 ;
        RECT 93.770 160.675 93.940 161.435 ;
        RECT 91.480 159.695 91.810 160.385 ;
        RECT 92.040 160.245 93.250 160.415 ;
        RECT 93.420 160.365 93.940 160.675 ;
        RECT 94.110 161.265 94.530 161.605 ;
        RECT 94.820 161.265 95.230 161.595 ;
        RECT 94.110 160.495 94.300 161.265 ;
        RECT 95.400 161.135 95.570 161.865 ;
        RECT 96.715 161.695 96.885 162.025 ;
        RECT 97.055 161.865 97.385 162.245 ;
        RECT 95.740 161.315 96.090 161.685 ;
        RECT 95.400 161.095 95.820 161.135 ;
        RECT 94.470 160.925 95.820 161.095 ;
        RECT 94.470 160.765 94.720 160.925 ;
        RECT 95.230 160.495 95.480 160.755 ;
        RECT 94.110 160.245 95.480 160.495 ;
        RECT 92.040 159.955 92.280 160.245 ;
        RECT 93.080 160.165 93.250 160.245 ;
        RECT 92.480 159.695 92.900 160.075 ;
        RECT 93.080 159.915 93.710 160.165 ;
        RECT 94.180 159.695 94.510 160.075 ;
        RECT 94.680 159.955 94.850 160.245 ;
        RECT 95.650 160.080 95.820 160.925 ;
        RECT 96.270 160.755 96.490 161.625 ;
        RECT 96.715 161.505 97.410 161.695 ;
        RECT 95.990 160.375 96.490 160.755 ;
        RECT 96.660 160.705 97.070 161.325 ;
        RECT 97.240 160.535 97.410 161.505 ;
        RECT 96.715 160.365 97.410 160.535 ;
        RECT 95.030 159.695 95.410 160.075 ;
        RECT 95.650 159.910 96.480 160.080 ;
        RECT 96.715 159.865 96.885 160.365 ;
        RECT 97.055 159.695 97.385 160.195 ;
        RECT 97.600 159.865 97.825 161.985 ;
        RECT 97.995 161.865 98.325 162.245 ;
        RECT 98.495 161.695 98.665 161.985 ;
        RECT 98.000 161.525 98.665 161.695 ;
        RECT 98.000 160.535 98.230 161.525 ;
        RECT 98.925 161.475 102.435 162.245 ;
        RECT 98.400 160.705 98.750 161.355 ;
        RECT 98.925 160.785 100.615 161.305 ;
        RECT 100.785 160.955 102.435 161.475 ;
        RECT 102.810 161.465 103.310 162.075 ;
        RECT 102.605 161.005 102.955 161.255 ;
        RECT 103.140 160.835 103.310 161.465 ;
        RECT 103.940 161.595 104.270 162.075 ;
        RECT 104.440 161.785 104.665 162.245 ;
        RECT 104.835 161.595 105.165 162.075 ;
        RECT 103.940 161.425 105.165 161.595 ;
        RECT 105.355 161.445 105.605 162.245 ;
        RECT 105.775 161.445 106.115 162.075 ;
        RECT 106.285 161.475 108.875 162.245 ;
        RECT 109.050 161.700 114.395 162.245 ;
        RECT 103.480 161.055 103.810 161.255 ;
        RECT 103.980 161.055 104.310 161.255 ;
        RECT 104.480 161.055 104.900 161.255 ;
        RECT 105.075 161.085 105.770 161.255 ;
        RECT 105.075 160.835 105.245 161.085 ;
        RECT 105.940 160.835 106.115 161.445 ;
        RECT 98.000 160.365 98.665 160.535 ;
        RECT 97.995 159.695 98.325 160.195 ;
        RECT 98.495 159.865 98.665 160.365 ;
        RECT 98.925 159.695 102.435 160.785 ;
        RECT 102.810 160.665 105.245 160.835 ;
        RECT 102.810 159.865 103.140 160.665 ;
        RECT 103.310 159.695 103.640 160.495 ;
        RECT 103.940 159.865 104.270 160.665 ;
        RECT 104.915 159.695 105.165 160.495 ;
        RECT 105.435 159.695 105.605 160.835 ;
        RECT 105.775 159.865 106.115 160.835 ;
        RECT 106.285 160.785 107.495 161.305 ;
        RECT 107.665 160.955 108.875 161.475 ;
        RECT 106.285 159.695 108.875 160.785 ;
        RECT 110.640 160.130 110.990 161.380 ;
        RECT 112.470 160.870 112.810 161.700 ;
        RECT 114.565 161.520 114.855 162.245 ;
        RECT 115.025 161.475 118.535 162.245 ;
        RECT 109.050 159.695 114.395 160.130 ;
        RECT 114.565 159.695 114.855 160.860 ;
        RECT 115.025 160.785 116.715 161.305 ;
        RECT 116.885 160.955 118.535 161.475 ;
        RECT 118.745 161.425 118.975 162.245 ;
        RECT 119.145 161.445 119.475 162.075 ;
        RECT 118.725 161.005 119.055 161.255 ;
        RECT 119.225 160.845 119.475 161.445 ;
        RECT 119.645 161.425 119.855 162.245 ;
        RECT 121.010 161.700 126.355 162.245 ;
        RECT 115.025 159.695 118.535 160.785 ;
        RECT 118.745 159.695 118.975 160.835 ;
        RECT 119.145 159.865 119.475 160.845 ;
        RECT 119.645 159.695 119.855 160.835 ;
        RECT 122.600 160.130 122.950 161.380 ;
        RECT 124.430 160.870 124.770 161.700 ;
        RECT 126.525 161.495 127.735 162.245 ;
        RECT 126.525 160.785 127.045 161.325 ;
        RECT 127.215 160.955 127.735 161.495 ;
        RECT 121.010 159.695 126.355 160.130 ;
        RECT 126.525 159.695 127.735 160.785 ;
        RECT 14.660 159.525 127.820 159.695 ;
        RECT 14.745 158.435 15.955 159.525 ;
        RECT 14.745 157.725 15.265 158.265 ;
        RECT 15.435 157.895 15.955 158.435 ;
        RECT 16.125 158.435 17.335 159.525 ;
        RECT 16.125 157.895 16.645 158.435 ;
        RECT 17.565 158.385 17.775 159.525 ;
        RECT 17.945 158.375 18.275 159.355 ;
        RECT 18.445 158.385 18.675 159.525 ;
        RECT 18.925 158.385 19.155 159.525 ;
        RECT 19.325 158.375 19.655 159.355 ;
        RECT 19.825 158.385 20.035 159.525 ;
        RECT 20.265 158.765 20.780 159.175 ;
        RECT 21.015 158.765 21.185 159.525 ;
        RECT 21.355 159.185 23.385 159.355 ;
        RECT 16.815 157.725 17.335 158.265 ;
        RECT 14.745 156.975 15.955 157.725 ;
        RECT 16.125 156.975 17.335 157.725 ;
        RECT 17.565 156.975 17.775 157.795 ;
        RECT 17.945 157.775 18.195 158.375 ;
        RECT 18.365 157.965 18.695 158.215 ;
        RECT 18.905 157.965 19.235 158.215 ;
        RECT 17.945 157.145 18.275 157.775 ;
        RECT 18.445 156.975 18.675 157.795 ;
        RECT 18.925 156.975 19.155 157.795 ;
        RECT 19.405 157.775 19.655 158.375 ;
        RECT 20.265 157.955 20.605 158.765 ;
        RECT 21.355 158.520 21.525 159.185 ;
        RECT 21.920 158.845 23.045 159.015 ;
        RECT 20.775 158.330 21.525 158.520 ;
        RECT 21.695 158.505 22.705 158.675 ;
        RECT 19.325 157.145 19.655 157.775 ;
        RECT 19.825 156.975 20.035 157.795 ;
        RECT 20.265 157.785 21.495 157.955 ;
        RECT 20.540 157.180 20.785 157.785 ;
        RECT 21.005 156.975 21.515 157.510 ;
        RECT 21.695 157.145 21.885 158.505 ;
        RECT 22.055 157.485 22.330 158.305 ;
        RECT 22.535 157.705 22.705 158.505 ;
        RECT 22.875 157.715 23.045 158.845 ;
        RECT 23.215 158.215 23.385 159.185 ;
        RECT 23.555 158.385 23.725 159.525 ;
        RECT 23.895 158.385 24.230 159.355 ;
        RECT 23.215 157.885 23.410 158.215 ;
        RECT 23.635 157.885 23.890 158.215 ;
        RECT 23.635 157.715 23.805 157.885 ;
        RECT 24.060 157.715 24.230 158.385 ;
        RECT 24.405 158.360 24.695 159.525 ;
        RECT 24.865 158.450 25.135 159.355 ;
        RECT 25.305 158.765 25.635 159.525 ;
        RECT 25.815 158.595 25.985 159.355 ;
        RECT 22.875 157.545 23.805 157.715 ;
        RECT 22.875 157.510 23.050 157.545 ;
        RECT 22.055 157.315 22.335 157.485 ;
        RECT 22.055 157.145 22.330 157.315 ;
        RECT 22.520 157.145 23.050 157.510 ;
        RECT 23.475 156.975 23.805 157.375 ;
        RECT 23.975 157.145 24.230 157.715 ;
        RECT 24.405 156.975 24.695 157.700 ;
        RECT 24.865 157.650 25.035 158.450 ;
        RECT 25.320 158.425 25.985 158.595 ;
        RECT 26.705 158.435 30.215 159.525 ;
        RECT 30.760 158.545 31.015 159.215 ;
        RECT 31.195 158.725 31.480 159.525 ;
        RECT 31.660 158.805 31.990 159.315 ;
        RECT 30.760 158.505 30.940 158.545 ;
        RECT 25.320 158.280 25.490 158.425 ;
        RECT 25.205 157.950 25.490 158.280 ;
        RECT 25.320 157.695 25.490 157.950 ;
        RECT 25.725 157.875 26.055 158.245 ;
        RECT 26.705 157.915 28.395 158.435 ;
        RECT 30.675 158.335 30.940 158.505 ;
        RECT 28.565 157.745 30.215 158.265 ;
        RECT 24.865 157.145 25.125 157.650 ;
        RECT 25.320 157.525 25.985 157.695 ;
        RECT 25.305 156.975 25.635 157.355 ;
        RECT 25.815 157.145 25.985 157.525 ;
        RECT 26.705 156.975 30.215 157.745 ;
        RECT 30.760 157.685 30.940 158.335 ;
        RECT 31.660 158.215 31.910 158.805 ;
        RECT 32.260 158.655 32.430 159.265 ;
        RECT 32.600 158.835 32.930 159.525 ;
        RECT 33.160 158.975 33.400 159.265 ;
        RECT 33.600 159.145 34.020 159.525 ;
        RECT 34.200 159.055 34.830 159.305 ;
        RECT 35.300 159.145 35.630 159.525 ;
        RECT 34.200 158.975 34.370 159.055 ;
        RECT 35.800 158.975 35.970 159.265 ;
        RECT 36.150 159.145 36.530 159.525 ;
        RECT 36.770 159.140 37.600 159.310 ;
        RECT 33.160 158.805 34.370 158.975 ;
        RECT 31.110 157.885 31.910 158.215 ;
        RECT 30.760 157.155 31.015 157.685 ;
        RECT 31.195 156.975 31.480 157.435 ;
        RECT 31.660 157.235 31.910 157.885 ;
        RECT 32.110 158.635 32.430 158.655 ;
        RECT 32.110 158.465 34.030 158.635 ;
        RECT 32.110 157.570 32.300 158.465 ;
        RECT 34.200 158.295 34.370 158.805 ;
        RECT 34.540 158.545 35.060 158.855 ;
        RECT 32.470 158.125 34.370 158.295 ;
        RECT 32.470 158.065 32.800 158.125 ;
        RECT 32.950 157.895 33.280 157.955 ;
        RECT 32.620 157.625 33.280 157.895 ;
        RECT 32.110 157.240 32.430 157.570 ;
        RECT 32.610 156.975 33.270 157.455 ;
        RECT 33.470 157.365 33.640 158.125 ;
        RECT 34.540 157.955 34.720 158.365 ;
        RECT 33.810 157.785 34.140 157.905 ;
        RECT 34.890 157.785 35.060 158.545 ;
        RECT 33.810 157.615 35.060 157.785 ;
        RECT 35.230 158.725 36.600 158.975 ;
        RECT 35.230 157.955 35.420 158.725 ;
        RECT 36.350 158.465 36.600 158.725 ;
        RECT 35.590 158.295 35.840 158.455 ;
        RECT 36.770 158.295 36.940 159.140 ;
        RECT 37.835 158.855 38.005 159.355 ;
        RECT 38.175 159.025 38.505 159.525 ;
        RECT 37.110 158.465 37.610 158.845 ;
        RECT 37.835 158.685 38.530 158.855 ;
        RECT 35.590 158.125 36.940 158.295 ;
        RECT 36.520 158.085 36.940 158.125 ;
        RECT 35.230 157.615 35.650 157.955 ;
        RECT 35.940 157.625 36.350 157.955 ;
        RECT 33.470 157.195 34.320 157.365 ;
        RECT 34.880 156.975 35.200 157.435 ;
        RECT 35.400 157.185 35.650 157.615 ;
        RECT 35.940 156.975 36.350 157.415 ;
        RECT 36.520 157.355 36.690 158.085 ;
        RECT 36.860 157.535 37.210 157.905 ;
        RECT 37.390 157.595 37.610 158.465 ;
        RECT 37.780 157.895 38.190 158.515 ;
        RECT 38.360 157.715 38.530 158.685 ;
        RECT 37.835 157.525 38.530 157.715 ;
        RECT 36.520 157.155 37.535 157.355 ;
        RECT 37.835 157.195 38.005 157.525 ;
        RECT 38.175 156.975 38.505 157.355 ;
        RECT 38.720 157.235 38.945 159.355 ;
        RECT 39.115 159.025 39.445 159.525 ;
        RECT 39.615 158.855 39.785 159.355 ;
        RECT 39.120 158.685 39.785 158.855 ;
        RECT 39.120 157.695 39.350 158.685 ;
        RECT 39.520 157.865 39.870 158.515 ;
        RECT 40.045 158.450 40.315 159.355 ;
        RECT 40.485 158.765 40.815 159.525 ;
        RECT 40.995 158.595 41.165 159.355 ;
        RECT 39.120 157.525 39.785 157.695 ;
        RECT 39.115 156.975 39.445 157.355 ;
        RECT 39.615 157.235 39.785 157.525 ;
        RECT 40.045 157.650 40.215 158.450 ;
        RECT 40.500 158.425 41.165 158.595 ;
        RECT 41.425 158.435 42.635 159.525 ;
        RECT 42.805 158.435 46.315 159.525 ;
        RECT 40.500 158.280 40.670 158.425 ;
        RECT 40.385 157.950 40.670 158.280 ;
        RECT 40.500 157.695 40.670 157.950 ;
        RECT 40.905 157.875 41.235 158.245 ;
        RECT 41.425 157.895 41.945 158.435 ;
        RECT 42.115 157.725 42.635 158.265 ;
        RECT 42.805 157.915 44.495 158.435 ;
        RECT 46.485 158.385 46.825 159.355 ;
        RECT 46.995 158.385 47.165 159.525 ;
        RECT 47.435 158.725 47.685 159.525 ;
        RECT 48.330 158.555 48.660 159.355 ;
        RECT 48.960 158.725 49.290 159.525 ;
        RECT 49.460 158.555 49.790 159.355 ;
        RECT 47.355 158.385 49.790 158.555 ;
        RECT 44.665 157.745 46.315 158.265 ;
        RECT 40.045 157.145 40.305 157.650 ;
        RECT 40.500 157.525 41.165 157.695 ;
        RECT 40.485 156.975 40.815 157.355 ;
        RECT 40.995 157.145 41.165 157.525 ;
        RECT 41.425 156.975 42.635 157.725 ;
        RECT 42.805 156.975 46.315 157.745 ;
        RECT 46.485 157.775 46.660 158.385 ;
        RECT 47.355 158.135 47.525 158.385 ;
        RECT 46.830 157.965 47.525 158.135 ;
        RECT 47.700 157.965 48.120 158.165 ;
        RECT 48.290 157.965 48.620 158.165 ;
        RECT 48.790 157.965 49.120 158.165 ;
        RECT 46.485 157.145 46.825 157.775 ;
        RECT 46.995 156.975 47.245 157.775 ;
        RECT 47.435 157.625 48.660 157.795 ;
        RECT 47.435 157.145 47.765 157.625 ;
        RECT 47.935 156.975 48.160 157.435 ;
        RECT 48.330 157.145 48.660 157.625 ;
        RECT 49.290 157.755 49.460 158.385 ;
        RECT 50.165 158.360 50.455 159.525 ;
        RECT 51.085 158.435 52.755 159.525 ;
        RECT 52.930 159.090 58.275 159.525 ;
        RECT 58.820 159.185 59.075 159.215 ;
        RECT 49.645 157.965 49.995 158.215 ;
        RECT 51.085 157.915 51.835 158.435 ;
        RECT 49.290 157.145 49.790 157.755 ;
        RECT 52.005 157.745 52.755 158.265 ;
        RECT 54.520 157.840 54.870 159.090 ;
        RECT 58.735 159.015 59.075 159.185 ;
        RECT 58.820 158.545 59.075 159.015 ;
        RECT 59.255 158.725 59.540 159.525 ;
        RECT 59.720 158.805 60.050 159.315 ;
        RECT 50.165 156.975 50.455 157.700 ;
        RECT 51.085 156.975 52.755 157.745 ;
        RECT 56.350 157.520 56.690 158.350 ;
        RECT 58.820 157.685 59.000 158.545 ;
        RECT 59.720 158.215 59.970 158.805 ;
        RECT 60.320 158.655 60.490 159.265 ;
        RECT 60.660 158.835 60.990 159.525 ;
        RECT 61.220 158.975 61.460 159.265 ;
        RECT 61.660 159.145 62.080 159.525 ;
        RECT 62.260 159.055 62.890 159.305 ;
        RECT 63.360 159.145 63.690 159.525 ;
        RECT 62.260 158.975 62.430 159.055 ;
        RECT 63.860 158.975 64.030 159.265 ;
        RECT 64.210 159.145 64.590 159.525 ;
        RECT 64.830 159.140 65.660 159.310 ;
        RECT 61.220 158.805 62.430 158.975 ;
        RECT 59.170 157.885 59.970 158.215 ;
        RECT 52.930 156.975 58.275 157.520 ;
        RECT 58.820 157.155 59.075 157.685 ;
        RECT 59.255 156.975 59.540 157.435 ;
        RECT 59.720 157.235 59.970 157.885 ;
        RECT 60.170 158.635 60.490 158.655 ;
        RECT 60.170 158.465 62.090 158.635 ;
        RECT 60.170 157.570 60.360 158.465 ;
        RECT 62.260 158.295 62.430 158.805 ;
        RECT 62.600 158.545 63.120 158.855 ;
        RECT 60.530 158.125 62.430 158.295 ;
        RECT 60.530 158.065 60.860 158.125 ;
        RECT 61.010 157.895 61.340 157.955 ;
        RECT 60.680 157.625 61.340 157.895 ;
        RECT 60.170 157.240 60.490 157.570 ;
        RECT 60.670 156.975 61.330 157.455 ;
        RECT 61.530 157.365 61.700 158.125 ;
        RECT 62.600 157.955 62.780 158.365 ;
        RECT 61.870 157.785 62.200 157.905 ;
        RECT 62.950 157.785 63.120 158.545 ;
        RECT 61.870 157.615 63.120 157.785 ;
        RECT 63.290 158.725 64.660 158.975 ;
        RECT 63.290 157.955 63.480 158.725 ;
        RECT 64.410 158.465 64.660 158.725 ;
        RECT 63.650 158.295 63.900 158.455 ;
        RECT 64.830 158.295 65.000 159.140 ;
        RECT 65.895 158.855 66.065 159.355 ;
        RECT 66.235 159.025 66.565 159.525 ;
        RECT 65.170 158.465 65.670 158.845 ;
        RECT 65.895 158.685 66.590 158.855 ;
        RECT 63.650 158.125 65.000 158.295 ;
        RECT 64.580 158.085 65.000 158.125 ;
        RECT 63.290 157.615 63.710 157.955 ;
        RECT 64.000 157.625 64.410 157.955 ;
        RECT 61.530 157.195 62.380 157.365 ;
        RECT 62.940 156.975 63.260 157.435 ;
        RECT 63.460 157.185 63.710 157.615 ;
        RECT 64.000 156.975 64.410 157.415 ;
        RECT 64.580 157.355 64.750 158.085 ;
        RECT 64.920 157.535 65.270 157.905 ;
        RECT 65.450 157.595 65.670 158.465 ;
        RECT 65.840 157.895 66.250 158.515 ;
        RECT 66.420 157.715 66.590 158.685 ;
        RECT 65.895 157.525 66.590 157.715 ;
        RECT 64.580 157.155 65.595 157.355 ;
        RECT 65.895 157.195 66.065 157.525 ;
        RECT 66.235 156.975 66.565 157.355 ;
        RECT 66.780 157.235 67.005 159.355 ;
        RECT 67.175 159.025 67.505 159.525 ;
        RECT 67.675 158.855 67.845 159.355 ;
        RECT 67.180 158.685 67.845 158.855 ;
        RECT 67.180 157.695 67.410 158.685 ;
        RECT 67.580 157.865 67.930 158.515 ;
        RECT 69.030 158.375 69.290 159.525 ;
        RECT 69.465 158.450 69.720 159.355 ;
        RECT 69.890 158.765 70.220 159.525 ;
        RECT 70.435 158.595 70.605 159.355 ;
        RECT 67.180 157.525 67.845 157.695 ;
        RECT 67.175 156.975 67.505 157.355 ;
        RECT 67.675 157.235 67.845 157.525 ;
        RECT 69.030 156.975 69.290 157.815 ;
        RECT 69.465 157.720 69.635 158.450 ;
        RECT 69.890 158.425 70.605 158.595 ;
        RECT 69.890 158.215 70.060 158.425 ;
        RECT 70.870 158.375 71.130 159.525 ;
        RECT 71.305 158.450 71.560 159.355 ;
        RECT 71.730 158.765 72.060 159.525 ;
        RECT 72.275 158.595 72.445 159.355 ;
        RECT 69.805 157.885 70.060 158.215 ;
        RECT 69.465 157.145 69.720 157.720 ;
        RECT 69.890 157.695 70.060 157.885 ;
        RECT 70.340 157.875 70.695 158.245 ;
        RECT 69.890 157.525 70.605 157.695 ;
        RECT 69.890 156.975 70.220 157.355 ;
        RECT 70.435 157.145 70.605 157.525 ;
        RECT 70.870 156.975 71.130 157.815 ;
        RECT 71.305 157.720 71.475 158.450 ;
        RECT 71.730 158.425 72.445 158.595 ;
        RECT 72.795 158.595 72.965 159.355 ;
        RECT 73.180 158.765 73.510 159.525 ;
        RECT 72.795 158.425 73.510 158.595 ;
        RECT 73.680 158.450 73.935 159.355 ;
        RECT 71.730 158.215 71.900 158.425 ;
        RECT 71.645 157.885 71.900 158.215 ;
        RECT 71.305 157.145 71.560 157.720 ;
        RECT 71.730 157.695 71.900 157.885 ;
        RECT 72.180 157.875 72.535 158.245 ;
        RECT 72.705 157.875 73.060 158.245 ;
        RECT 73.340 158.215 73.510 158.425 ;
        RECT 73.340 157.885 73.595 158.215 ;
        RECT 73.340 157.695 73.510 157.885 ;
        RECT 73.765 157.720 73.935 158.450 ;
        RECT 74.110 158.375 74.370 159.525 ;
        RECT 74.545 158.435 75.755 159.525 ;
        RECT 74.545 157.895 75.065 158.435 ;
        RECT 75.925 158.360 76.215 159.525 ;
        RECT 76.475 158.595 76.645 159.355 ;
        RECT 76.860 158.765 77.190 159.525 ;
        RECT 76.475 158.425 77.190 158.595 ;
        RECT 77.360 158.450 77.615 159.355 ;
        RECT 71.730 157.525 72.445 157.695 ;
        RECT 71.730 156.975 72.060 157.355 ;
        RECT 72.275 157.145 72.445 157.525 ;
        RECT 72.795 157.525 73.510 157.695 ;
        RECT 72.795 157.145 72.965 157.525 ;
        RECT 73.180 156.975 73.510 157.355 ;
        RECT 73.680 157.145 73.935 157.720 ;
        RECT 74.110 156.975 74.370 157.815 ;
        RECT 75.235 157.725 75.755 158.265 ;
        RECT 76.385 157.875 76.740 158.245 ;
        RECT 77.020 158.215 77.190 158.425 ;
        RECT 77.020 157.885 77.275 158.215 ;
        RECT 74.545 156.975 75.755 157.725 ;
        RECT 75.925 156.975 76.215 157.700 ;
        RECT 77.020 157.695 77.190 157.885 ;
        RECT 77.445 157.720 77.615 158.450 ;
        RECT 77.790 158.375 78.050 159.525 ;
        RECT 78.225 158.435 79.435 159.525 ;
        RECT 79.610 159.090 84.955 159.525 ;
        RECT 85.130 159.090 90.475 159.525 ;
        RECT 90.650 159.090 95.995 159.525 ;
        RECT 96.170 159.090 101.515 159.525 ;
        RECT 78.225 157.895 78.745 158.435 ;
        RECT 76.475 157.525 77.190 157.695 ;
        RECT 76.475 157.145 76.645 157.525 ;
        RECT 76.860 156.975 77.190 157.355 ;
        RECT 77.360 157.145 77.615 157.720 ;
        RECT 77.790 156.975 78.050 157.815 ;
        RECT 78.915 157.725 79.435 158.265 ;
        RECT 81.200 157.840 81.550 159.090 ;
        RECT 78.225 156.975 79.435 157.725 ;
        RECT 83.030 157.520 83.370 158.350 ;
        RECT 86.720 157.840 87.070 159.090 ;
        RECT 88.550 157.520 88.890 158.350 ;
        RECT 92.240 157.840 92.590 159.090 ;
        RECT 94.070 157.520 94.410 158.350 ;
        RECT 97.760 157.840 98.110 159.090 ;
        RECT 101.685 158.360 101.975 159.525 ;
        RECT 103.270 158.555 103.600 159.355 ;
        RECT 103.770 158.725 104.100 159.525 ;
        RECT 104.400 158.555 104.730 159.355 ;
        RECT 105.375 158.725 105.625 159.525 ;
        RECT 103.270 158.385 105.705 158.555 ;
        RECT 105.895 158.385 106.065 159.525 ;
        RECT 106.235 158.385 106.575 159.355 ;
        RECT 99.590 157.520 99.930 158.350 ;
        RECT 103.065 157.965 103.415 158.215 ;
        RECT 103.600 157.755 103.770 158.385 ;
        RECT 103.940 157.965 104.270 158.165 ;
        RECT 104.440 157.965 104.770 158.165 ;
        RECT 104.940 157.965 105.360 158.165 ;
        RECT 105.535 158.135 105.705 158.385 ;
        RECT 105.535 157.965 106.230 158.135 ;
        RECT 79.610 156.975 84.955 157.520 ;
        RECT 85.130 156.975 90.475 157.520 ;
        RECT 90.650 156.975 95.995 157.520 ;
        RECT 96.170 156.975 101.515 157.520 ;
        RECT 101.685 156.975 101.975 157.700 ;
        RECT 103.270 157.145 103.770 157.755 ;
        RECT 104.400 157.625 105.625 157.795 ;
        RECT 106.400 157.775 106.575 158.385 ;
        RECT 104.400 157.145 104.730 157.625 ;
        RECT 104.900 156.975 105.125 157.435 ;
        RECT 105.295 157.145 105.625 157.625 ;
        RECT 105.815 156.975 106.065 157.775 ;
        RECT 106.235 157.145 106.575 157.775 ;
        RECT 107.665 158.385 107.935 159.355 ;
        RECT 108.145 158.725 108.425 159.525 ;
        RECT 108.595 159.015 110.250 159.305 ;
        RECT 108.660 158.675 110.250 158.845 ;
        RECT 108.660 158.555 108.830 158.675 ;
        RECT 108.105 158.385 108.830 158.555 ;
        RECT 107.665 157.650 107.835 158.385 ;
        RECT 108.105 158.215 108.275 158.385 ;
        RECT 109.020 158.335 109.735 158.505 ;
        RECT 109.930 158.385 110.250 158.675 ;
        RECT 110.425 158.385 110.765 159.355 ;
        RECT 110.935 158.385 111.105 159.525 ;
        RECT 111.375 158.725 111.625 159.525 ;
        RECT 112.270 158.555 112.600 159.355 ;
        RECT 112.900 158.725 113.230 159.525 ;
        RECT 113.400 158.555 113.730 159.355 ;
        RECT 111.295 158.385 113.730 158.555 ;
        RECT 114.105 158.435 115.315 159.525 ;
        RECT 108.005 157.885 108.275 158.215 ;
        RECT 108.445 157.885 108.850 158.215 ;
        RECT 109.020 157.885 109.730 158.335 ;
        RECT 108.105 157.715 108.275 157.885 ;
        RECT 107.665 157.305 107.935 157.650 ;
        RECT 108.105 157.545 109.715 157.715 ;
        RECT 109.900 157.645 110.250 158.215 ;
        RECT 110.425 157.825 110.600 158.385 ;
        RECT 111.295 158.135 111.465 158.385 ;
        RECT 110.770 157.965 111.465 158.135 ;
        RECT 111.640 157.965 112.060 158.165 ;
        RECT 112.230 157.965 112.560 158.165 ;
        RECT 112.730 157.965 113.060 158.165 ;
        RECT 110.425 157.775 110.655 157.825 ;
        RECT 108.125 156.975 108.505 157.375 ;
        RECT 108.675 157.195 108.845 157.545 ;
        RECT 109.015 156.975 109.345 157.375 ;
        RECT 109.545 157.195 109.715 157.545 ;
        RECT 109.915 156.975 110.245 157.475 ;
        RECT 110.425 157.145 110.765 157.775 ;
        RECT 110.935 156.975 111.185 157.775 ;
        RECT 111.375 157.625 112.600 157.795 ;
        RECT 111.375 157.145 111.705 157.625 ;
        RECT 111.875 156.975 112.100 157.435 ;
        RECT 112.270 157.145 112.600 157.625 ;
        RECT 113.230 157.755 113.400 158.385 ;
        RECT 113.585 157.965 113.935 158.215 ;
        RECT 114.105 157.895 114.625 158.435 ;
        RECT 115.490 158.335 115.745 159.215 ;
        RECT 115.915 158.385 116.220 159.525 ;
        RECT 116.560 159.145 116.890 159.525 ;
        RECT 117.070 158.975 117.240 159.265 ;
        RECT 117.410 159.065 117.660 159.525 ;
        RECT 116.440 158.805 117.240 158.975 ;
        RECT 117.830 159.015 118.700 159.355 ;
        RECT 113.230 157.145 113.730 157.755 ;
        RECT 114.795 157.725 115.315 158.265 ;
        RECT 114.105 156.975 115.315 157.725 ;
        RECT 115.490 157.685 115.700 158.335 ;
        RECT 116.440 158.215 116.610 158.805 ;
        RECT 117.830 158.635 118.000 159.015 ;
        RECT 118.935 158.895 119.105 159.355 ;
        RECT 119.275 159.065 119.645 159.525 ;
        RECT 119.940 158.925 120.110 159.265 ;
        RECT 120.280 159.095 120.610 159.525 ;
        RECT 120.845 158.925 121.015 159.265 ;
        RECT 116.780 158.465 118.000 158.635 ;
        RECT 118.170 158.555 118.630 158.845 ;
        RECT 118.935 158.725 119.495 158.895 ;
        RECT 119.940 158.755 121.015 158.925 ;
        RECT 121.185 159.025 121.865 159.355 ;
        RECT 122.080 159.025 122.330 159.355 ;
        RECT 122.500 159.065 122.750 159.525 ;
        RECT 119.325 158.585 119.495 158.725 ;
        RECT 118.170 158.545 119.135 158.555 ;
        RECT 117.830 158.375 118.000 158.465 ;
        RECT 118.460 158.385 119.135 158.545 ;
        RECT 115.870 158.185 116.610 158.215 ;
        RECT 115.870 157.885 116.785 158.185 ;
        RECT 116.460 157.710 116.785 157.885 ;
        RECT 115.490 157.155 115.745 157.685 ;
        RECT 115.915 156.975 116.220 157.435 ;
        RECT 116.465 157.355 116.785 157.710 ;
        RECT 116.955 157.925 117.495 158.295 ;
        RECT 117.830 158.205 118.235 158.375 ;
        RECT 116.955 157.525 117.195 157.925 ;
        RECT 117.675 157.755 117.895 158.035 ;
        RECT 117.365 157.585 117.895 157.755 ;
        RECT 117.365 157.355 117.535 157.585 ;
        RECT 118.065 157.425 118.235 158.205 ;
        RECT 118.405 157.595 118.755 158.215 ;
        RECT 118.925 157.595 119.135 158.385 ;
        RECT 119.325 158.415 120.825 158.585 ;
        RECT 119.325 157.725 119.495 158.415 ;
        RECT 121.185 158.245 121.355 159.025 ;
        RECT 122.160 158.895 122.330 159.025 ;
        RECT 119.665 158.075 121.355 158.245 ;
        RECT 121.525 158.465 121.990 158.855 ;
        RECT 122.160 158.725 122.555 158.895 ;
        RECT 119.665 157.895 119.835 158.075 ;
        RECT 116.465 157.185 117.535 157.355 ;
        RECT 117.705 156.975 117.895 157.415 ;
        RECT 118.065 157.145 119.015 157.425 ;
        RECT 119.325 157.335 119.585 157.725 ;
        RECT 120.005 157.655 120.795 157.905 ;
        RECT 119.235 157.165 119.585 157.335 ;
        RECT 119.795 156.975 120.125 157.435 ;
        RECT 121.000 157.365 121.170 158.075 ;
        RECT 121.525 157.875 121.695 158.465 ;
        RECT 121.340 157.655 121.695 157.875 ;
        RECT 121.865 157.655 122.215 158.275 ;
        RECT 122.385 157.365 122.555 158.725 ;
        RECT 122.920 158.555 123.245 159.340 ;
        RECT 122.725 157.505 123.185 158.555 ;
        RECT 121.000 157.195 121.855 157.365 ;
        RECT 122.060 157.195 122.555 157.365 ;
        RECT 122.725 156.975 123.055 157.335 ;
        RECT 123.415 157.235 123.585 159.355 ;
        RECT 123.755 159.025 124.085 159.525 ;
        RECT 124.255 158.855 124.510 159.355 ;
        RECT 123.760 158.685 124.510 158.855 ;
        RECT 123.760 157.695 123.990 158.685 ;
        RECT 124.160 157.865 124.510 158.515 ;
        RECT 124.685 158.435 126.355 159.525 ;
        RECT 126.525 158.435 127.735 159.525 ;
        RECT 124.685 157.915 125.435 158.435 ;
        RECT 125.605 157.745 126.355 158.265 ;
        RECT 126.525 157.895 127.045 158.435 ;
        RECT 123.760 157.525 124.510 157.695 ;
        RECT 123.755 156.975 124.085 157.355 ;
        RECT 124.255 157.235 124.510 157.525 ;
        RECT 124.685 156.975 126.355 157.745 ;
        RECT 127.215 157.725 127.735 158.265 ;
        RECT 126.525 156.975 127.735 157.725 ;
        RECT 14.660 156.805 127.820 156.975 ;
        RECT 14.745 156.055 15.955 156.805 ;
        RECT 14.745 155.515 15.265 156.055 ;
        RECT 16.125 156.035 17.795 156.805 ;
        RECT 15.435 155.345 15.955 155.885 ;
        RECT 14.745 154.255 15.955 155.345 ;
        RECT 16.125 155.345 16.875 155.865 ;
        RECT 17.045 155.515 17.795 156.035 ;
        RECT 17.970 156.095 18.225 156.625 ;
        RECT 18.395 156.345 18.700 156.805 ;
        RECT 18.945 156.425 20.015 156.595 ;
        RECT 17.970 155.445 18.180 156.095 ;
        RECT 18.945 156.070 19.265 156.425 ;
        RECT 18.940 155.895 19.265 156.070 ;
        RECT 18.350 155.595 19.265 155.895 ;
        RECT 19.435 155.855 19.675 156.255 ;
        RECT 19.845 156.195 20.015 156.425 ;
        RECT 20.185 156.365 20.375 156.805 ;
        RECT 20.545 156.355 21.495 156.635 ;
        RECT 21.715 156.445 22.065 156.615 ;
        RECT 19.845 156.025 20.375 156.195 ;
        RECT 18.350 155.565 19.090 155.595 ;
        RECT 16.125 154.255 17.795 155.345 ;
        RECT 17.970 154.565 18.225 155.445 ;
        RECT 18.395 154.255 18.700 155.395 ;
        RECT 18.920 154.975 19.090 155.565 ;
        RECT 19.435 155.485 19.975 155.855 ;
        RECT 20.155 155.745 20.375 156.025 ;
        RECT 20.545 155.575 20.715 156.355 ;
        RECT 20.310 155.405 20.715 155.575 ;
        RECT 20.885 155.565 21.235 156.185 ;
        RECT 20.310 155.315 20.480 155.405 ;
        RECT 21.405 155.395 21.615 156.185 ;
        RECT 19.260 155.145 20.480 155.315 ;
        RECT 20.940 155.235 21.615 155.395 ;
        RECT 18.920 154.805 19.720 154.975 ;
        RECT 19.040 154.255 19.370 154.635 ;
        RECT 19.550 154.515 19.720 154.805 ;
        RECT 20.310 154.765 20.480 155.145 ;
        RECT 20.650 155.225 21.615 155.235 ;
        RECT 21.805 156.055 22.065 156.445 ;
        RECT 22.275 156.345 22.605 156.805 ;
        RECT 23.480 156.415 24.335 156.585 ;
        RECT 24.540 156.415 25.035 156.585 ;
        RECT 25.205 156.445 25.535 156.805 ;
        RECT 21.805 155.365 21.975 156.055 ;
        RECT 22.145 155.705 22.315 155.885 ;
        RECT 22.485 155.875 23.275 156.125 ;
        RECT 23.480 155.705 23.650 156.415 ;
        RECT 23.820 155.905 24.175 156.125 ;
        RECT 22.145 155.535 23.835 155.705 ;
        RECT 20.650 154.935 21.110 155.225 ;
        RECT 21.805 155.195 23.305 155.365 ;
        RECT 21.805 155.055 21.975 155.195 ;
        RECT 21.415 154.885 21.975 155.055 ;
        RECT 19.890 154.255 20.140 154.715 ;
        RECT 20.310 154.425 21.180 154.765 ;
        RECT 21.415 154.425 21.585 154.885 ;
        RECT 22.420 154.855 23.495 155.025 ;
        RECT 21.755 154.255 22.125 154.715 ;
        RECT 22.420 154.515 22.590 154.855 ;
        RECT 22.760 154.255 23.090 154.685 ;
        RECT 23.325 154.515 23.495 154.855 ;
        RECT 23.665 154.755 23.835 155.535 ;
        RECT 24.005 155.315 24.175 155.905 ;
        RECT 24.345 155.505 24.695 156.125 ;
        RECT 24.005 154.925 24.470 155.315 ;
        RECT 24.865 155.055 25.035 156.415 ;
        RECT 25.205 155.225 25.665 156.275 ;
        RECT 24.640 154.885 25.035 155.055 ;
        RECT 24.640 154.755 24.810 154.885 ;
        RECT 23.665 154.425 24.345 154.755 ;
        RECT 24.560 154.425 24.810 154.755 ;
        RECT 24.980 154.255 25.230 154.715 ;
        RECT 25.400 154.440 25.725 155.225 ;
        RECT 25.895 154.425 26.065 156.545 ;
        RECT 26.235 156.425 26.565 156.805 ;
        RECT 26.735 156.255 26.990 156.545 ;
        RECT 26.240 156.085 26.990 156.255 ;
        RECT 27.165 156.130 27.425 156.635 ;
        RECT 27.605 156.425 27.935 156.805 ;
        RECT 28.115 156.255 28.285 156.635 ;
        RECT 26.240 155.095 26.470 156.085 ;
        RECT 26.640 155.265 26.990 155.915 ;
        RECT 27.165 155.330 27.335 156.130 ;
        RECT 27.620 156.085 28.285 156.255 ;
        RECT 27.620 155.830 27.790 156.085 ;
        RECT 29.465 156.035 32.975 156.805 ;
        RECT 27.505 155.500 27.790 155.830 ;
        RECT 28.025 155.535 28.355 155.905 ;
        RECT 27.620 155.355 27.790 155.500 ;
        RECT 26.240 154.925 26.990 155.095 ;
        RECT 26.235 154.255 26.565 154.755 ;
        RECT 26.735 154.425 26.990 154.925 ;
        RECT 27.165 154.425 27.435 155.330 ;
        RECT 27.620 155.185 28.285 155.355 ;
        RECT 27.605 154.255 27.935 155.015 ;
        RECT 28.115 154.425 28.285 155.185 ;
        RECT 29.465 155.345 31.155 155.865 ;
        RECT 31.325 155.515 32.975 156.035 ;
        RECT 33.420 155.995 33.665 156.600 ;
        RECT 33.885 156.270 34.395 156.805 ;
        RECT 33.145 155.825 34.375 155.995 ;
        RECT 29.465 154.255 32.975 155.345 ;
        RECT 33.145 155.015 33.485 155.825 ;
        RECT 33.655 155.260 34.405 155.450 ;
        RECT 33.145 154.605 33.660 155.015 ;
        RECT 33.895 154.255 34.065 155.015 ;
        RECT 34.235 154.595 34.405 155.260 ;
        RECT 34.575 155.275 34.765 156.635 ;
        RECT 34.935 156.125 35.210 156.635 ;
        RECT 35.400 156.270 35.930 156.635 ;
        RECT 36.355 156.405 36.685 156.805 ;
        RECT 35.755 156.235 35.930 156.270 ;
        RECT 34.935 155.955 35.215 156.125 ;
        RECT 34.935 155.475 35.210 155.955 ;
        RECT 35.415 155.275 35.585 156.075 ;
        RECT 34.575 155.105 35.585 155.275 ;
        RECT 35.755 156.065 36.685 156.235 ;
        RECT 36.855 156.065 37.110 156.635 ;
        RECT 37.285 156.080 37.575 156.805 ;
        RECT 35.755 154.935 35.925 156.065 ;
        RECT 36.515 155.895 36.685 156.065 ;
        RECT 34.800 154.765 35.925 154.935 ;
        RECT 36.095 155.565 36.290 155.895 ;
        RECT 36.515 155.565 36.770 155.895 ;
        RECT 36.095 154.595 36.265 155.565 ;
        RECT 36.940 155.395 37.110 156.065 ;
        RECT 37.745 156.055 38.955 156.805 ;
        RECT 34.235 154.425 36.265 154.595 ;
        RECT 36.435 154.255 36.605 155.395 ;
        RECT 36.775 154.425 37.110 155.395 ;
        RECT 37.285 154.255 37.575 155.420 ;
        RECT 37.745 155.345 38.265 155.885 ;
        RECT 38.435 155.515 38.955 156.055 ;
        RECT 39.125 156.035 42.635 156.805 ;
        RECT 39.125 155.345 40.815 155.865 ;
        RECT 40.985 155.515 42.635 156.035 ;
        RECT 42.805 156.130 43.075 156.475 ;
        RECT 43.265 156.405 43.645 156.805 ;
        RECT 43.815 156.235 43.985 156.585 ;
        RECT 44.155 156.405 44.485 156.805 ;
        RECT 44.685 156.235 44.855 156.585 ;
        RECT 45.055 156.305 45.385 156.805 ;
        RECT 42.805 155.395 42.975 156.130 ;
        RECT 43.245 156.065 44.855 156.235 ;
        RECT 43.245 155.895 43.415 156.065 ;
        RECT 43.145 155.565 43.415 155.895 ;
        RECT 43.585 155.565 43.990 155.895 ;
        RECT 43.245 155.395 43.415 155.565 ;
        RECT 44.160 155.445 44.870 155.895 ;
        RECT 45.040 155.565 45.390 156.135 ;
        RECT 45.565 156.005 45.905 156.635 ;
        RECT 46.075 156.005 46.325 156.805 ;
        RECT 46.515 156.155 46.845 156.635 ;
        RECT 47.015 156.345 47.240 156.805 ;
        RECT 47.410 156.155 47.740 156.635 ;
        RECT 45.565 155.955 45.795 156.005 ;
        RECT 46.515 155.985 47.740 156.155 ;
        RECT 48.370 156.025 48.870 156.635 ;
        RECT 49.450 156.025 49.950 156.635 ;
        RECT 37.745 154.255 38.955 155.345 ;
        RECT 39.125 154.255 42.635 155.345 ;
        RECT 42.805 154.425 43.075 155.395 ;
        RECT 43.245 155.225 43.970 155.395 ;
        RECT 44.160 155.275 44.875 155.445 ;
        RECT 45.565 155.395 45.740 155.955 ;
        RECT 45.910 155.645 46.605 155.815 ;
        RECT 46.435 155.395 46.605 155.645 ;
        RECT 46.780 155.615 47.200 155.815 ;
        RECT 47.370 155.615 47.700 155.815 ;
        RECT 47.870 155.615 48.200 155.815 ;
        RECT 48.370 155.395 48.540 156.025 ;
        RECT 48.725 155.565 49.075 155.815 ;
        RECT 49.245 155.565 49.595 155.815 ;
        RECT 49.780 155.395 49.950 156.025 ;
        RECT 50.580 156.155 50.910 156.635 ;
        RECT 51.080 156.345 51.305 156.805 ;
        RECT 51.475 156.155 51.805 156.635 ;
        RECT 50.580 155.985 51.805 156.155 ;
        RECT 51.995 156.005 52.245 156.805 ;
        RECT 52.415 156.005 52.755 156.635 ;
        RECT 53.850 156.260 59.195 156.805 ;
        RECT 50.120 155.615 50.450 155.815 ;
        RECT 50.620 155.615 50.950 155.815 ;
        RECT 51.120 155.615 51.540 155.815 ;
        RECT 51.715 155.645 52.410 155.815 ;
        RECT 51.715 155.395 51.885 155.645 ;
        RECT 52.580 155.395 52.755 156.005 ;
        RECT 43.800 155.105 43.970 155.225 ;
        RECT 45.070 155.105 45.390 155.395 ;
        RECT 43.285 154.255 43.565 155.055 ;
        RECT 43.800 154.935 45.390 155.105 ;
        RECT 43.735 154.475 45.390 154.765 ;
        RECT 45.565 154.425 45.905 155.395 ;
        RECT 46.075 154.255 46.245 155.395 ;
        RECT 46.435 155.225 48.870 155.395 ;
        RECT 46.515 154.255 46.765 155.055 ;
        RECT 47.410 154.425 47.740 155.225 ;
        RECT 48.040 154.255 48.370 155.055 ;
        RECT 48.540 154.425 48.870 155.225 ;
        RECT 49.450 155.225 51.885 155.395 ;
        RECT 49.450 154.425 49.780 155.225 ;
        RECT 49.950 154.255 50.280 155.055 ;
        RECT 50.580 154.425 50.910 155.225 ;
        RECT 51.555 154.255 51.805 155.055 ;
        RECT 52.075 154.255 52.245 155.395 ;
        RECT 52.415 154.425 52.755 155.395 ;
        RECT 55.440 154.690 55.790 155.940 ;
        RECT 57.270 155.430 57.610 156.260 ;
        RECT 59.570 156.025 60.070 156.635 ;
        RECT 59.365 155.565 59.715 155.815 ;
        RECT 59.900 155.395 60.070 156.025 ;
        RECT 60.700 156.155 61.030 156.635 ;
        RECT 61.200 156.345 61.425 156.805 ;
        RECT 61.595 156.155 61.925 156.635 ;
        RECT 60.700 155.985 61.925 156.155 ;
        RECT 62.115 156.005 62.365 156.805 ;
        RECT 62.535 156.005 62.875 156.635 ;
        RECT 63.045 156.080 63.335 156.805 ;
        RECT 63.505 156.055 64.715 156.805 ;
        RECT 60.240 155.615 60.570 155.815 ;
        RECT 60.740 155.615 61.070 155.815 ;
        RECT 61.240 155.615 61.660 155.815 ;
        RECT 61.835 155.645 62.530 155.815 ;
        RECT 61.835 155.395 62.005 155.645 ;
        RECT 62.700 155.445 62.875 156.005 ;
        RECT 62.645 155.395 62.875 155.445 ;
        RECT 59.570 155.225 62.005 155.395 ;
        RECT 53.850 154.255 59.195 154.690 ;
        RECT 59.570 154.425 59.900 155.225 ;
        RECT 60.070 154.255 60.400 155.055 ;
        RECT 60.700 154.425 61.030 155.225 ;
        RECT 61.675 154.255 61.925 155.055 ;
        RECT 62.195 154.255 62.365 155.395 ;
        RECT 62.535 154.425 62.875 155.395 ;
        RECT 63.045 154.255 63.335 155.420 ;
        RECT 63.505 155.345 64.025 155.885 ;
        RECT 64.195 155.515 64.715 156.055 ;
        RECT 64.925 155.985 65.155 156.805 ;
        RECT 65.325 156.005 65.655 156.635 ;
        RECT 64.905 155.565 65.235 155.815 ;
        RECT 65.405 155.405 65.655 156.005 ;
        RECT 65.825 155.985 66.035 156.805 ;
        RECT 66.640 156.095 66.895 156.625 ;
        RECT 67.075 156.345 67.360 156.805 ;
        RECT 63.505 154.255 64.715 155.345 ;
        RECT 64.925 154.255 65.155 155.395 ;
        RECT 65.325 154.425 65.655 155.405 ;
        RECT 65.825 154.255 66.035 155.395 ;
        RECT 66.640 155.235 66.820 156.095 ;
        RECT 67.540 155.895 67.790 156.545 ;
        RECT 66.990 155.565 67.790 155.895 ;
        RECT 66.640 155.105 66.895 155.235 ;
        RECT 66.555 154.935 66.895 155.105 ;
        RECT 66.640 154.565 66.895 154.935 ;
        RECT 67.075 154.255 67.360 155.055 ;
        RECT 67.540 154.975 67.790 155.565 ;
        RECT 67.990 156.210 68.310 156.540 ;
        RECT 68.490 156.325 69.150 156.805 ;
        RECT 69.350 156.415 70.200 156.585 ;
        RECT 67.990 155.315 68.180 156.210 ;
        RECT 68.500 155.885 69.160 156.155 ;
        RECT 68.830 155.825 69.160 155.885 ;
        RECT 68.350 155.655 68.680 155.715 ;
        RECT 69.350 155.655 69.520 156.415 ;
        RECT 70.760 156.345 71.080 156.805 ;
        RECT 71.280 156.165 71.530 156.595 ;
        RECT 71.820 156.365 72.230 156.805 ;
        RECT 72.400 156.425 73.415 156.625 ;
        RECT 69.690 155.995 70.940 156.165 ;
        RECT 69.690 155.875 70.020 155.995 ;
        RECT 68.350 155.485 70.250 155.655 ;
        RECT 67.990 155.145 69.910 155.315 ;
        RECT 67.990 155.125 68.310 155.145 ;
        RECT 67.540 154.465 67.870 154.975 ;
        RECT 68.140 154.515 68.310 155.125 ;
        RECT 70.080 154.975 70.250 155.485 ;
        RECT 70.420 155.415 70.600 155.825 ;
        RECT 70.770 155.235 70.940 155.995 ;
        RECT 68.480 154.255 68.810 154.945 ;
        RECT 69.040 154.805 70.250 154.975 ;
        RECT 70.420 154.925 70.940 155.235 ;
        RECT 71.110 155.825 71.530 156.165 ;
        RECT 71.820 155.825 72.230 156.155 ;
        RECT 71.110 155.055 71.300 155.825 ;
        RECT 72.400 155.695 72.570 156.425 ;
        RECT 73.715 156.255 73.885 156.585 ;
        RECT 74.055 156.425 74.385 156.805 ;
        RECT 72.740 155.875 73.090 156.245 ;
        RECT 72.400 155.655 72.820 155.695 ;
        RECT 71.470 155.485 72.820 155.655 ;
        RECT 71.470 155.325 71.720 155.485 ;
        RECT 72.230 155.055 72.480 155.315 ;
        RECT 71.110 154.805 72.480 155.055 ;
        RECT 69.040 154.515 69.280 154.805 ;
        RECT 70.080 154.725 70.250 154.805 ;
        RECT 69.480 154.255 69.900 154.635 ;
        RECT 70.080 154.475 70.710 154.725 ;
        RECT 71.180 154.255 71.510 154.635 ;
        RECT 71.680 154.515 71.850 154.805 ;
        RECT 72.650 154.640 72.820 155.485 ;
        RECT 73.270 155.315 73.490 156.185 ;
        RECT 73.715 156.065 74.410 156.255 ;
        RECT 72.990 154.935 73.490 155.315 ;
        RECT 73.660 155.265 74.070 155.885 ;
        RECT 74.240 155.095 74.410 156.065 ;
        RECT 73.715 154.925 74.410 155.095 ;
        RECT 72.030 154.255 72.410 154.635 ;
        RECT 72.650 154.470 73.480 154.640 ;
        RECT 73.715 154.425 73.885 154.925 ;
        RECT 74.055 154.255 74.385 154.755 ;
        RECT 74.600 154.425 74.825 156.545 ;
        RECT 74.995 156.425 75.325 156.805 ;
        RECT 75.495 156.255 75.665 156.545 ;
        RECT 75.000 156.085 75.665 156.255 ;
        RECT 75.000 155.095 75.230 156.085 ;
        RECT 75.930 155.965 76.190 156.805 ;
        RECT 76.365 156.060 76.620 156.635 ;
        RECT 76.790 156.425 77.120 156.805 ;
        RECT 77.335 156.255 77.505 156.635 ;
        RECT 77.770 156.260 83.115 156.805 ;
        RECT 83.290 156.260 88.635 156.805 ;
        RECT 76.790 156.085 77.505 156.255 ;
        RECT 75.400 155.265 75.750 155.915 ;
        RECT 75.000 154.925 75.665 155.095 ;
        RECT 74.995 154.255 75.325 154.755 ;
        RECT 75.495 154.425 75.665 154.925 ;
        RECT 75.930 154.255 76.190 155.405 ;
        RECT 76.365 155.330 76.535 156.060 ;
        RECT 76.790 155.895 76.960 156.085 ;
        RECT 76.705 155.565 76.960 155.895 ;
        RECT 76.790 155.355 76.960 155.565 ;
        RECT 77.240 155.535 77.595 155.905 ;
        RECT 76.365 154.425 76.620 155.330 ;
        RECT 76.790 155.185 77.505 155.355 ;
        RECT 76.790 154.255 77.120 155.015 ;
        RECT 77.335 154.425 77.505 155.185 ;
        RECT 79.360 154.690 79.710 155.940 ;
        RECT 81.190 155.430 81.530 156.260 ;
        RECT 84.880 154.690 85.230 155.940 ;
        RECT 86.710 155.430 87.050 156.260 ;
        RECT 88.805 156.080 89.095 156.805 ;
        RECT 90.185 156.035 93.695 156.805 ;
        RECT 93.955 156.255 94.125 156.635 ;
        RECT 94.305 156.425 94.635 156.805 ;
        RECT 93.955 156.085 94.620 156.255 ;
        RECT 94.815 156.130 95.075 156.635 ;
        RECT 77.770 154.255 83.115 154.690 ;
        RECT 83.290 154.255 88.635 154.690 ;
        RECT 88.805 154.255 89.095 155.420 ;
        RECT 90.185 155.345 91.875 155.865 ;
        RECT 92.045 155.515 93.695 156.035 ;
        RECT 93.885 155.535 94.215 155.905 ;
        RECT 94.450 155.830 94.620 156.085 ;
        RECT 94.450 155.500 94.735 155.830 ;
        RECT 94.450 155.355 94.620 155.500 ;
        RECT 90.185 154.255 93.695 155.345 ;
        RECT 93.955 155.185 94.620 155.355 ;
        RECT 94.905 155.330 95.075 156.130 ;
        RECT 95.705 156.035 97.375 156.805 ;
        RECT 93.955 154.425 94.125 155.185 ;
        RECT 94.305 154.255 94.635 155.015 ;
        RECT 94.805 154.425 95.075 155.330 ;
        RECT 95.705 155.345 96.455 155.865 ;
        RECT 96.625 155.515 97.375 156.035 ;
        RECT 97.545 156.005 97.885 156.635 ;
        RECT 98.055 156.005 98.305 156.805 ;
        RECT 98.495 156.155 98.825 156.635 ;
        RECT 98.995 156.345 99.220 156.805 ;
        RECT 99.390 156.155 99.720 156.635 ;
        RECT 97.545 155.395 97.720 156.005 ;
        RECT 98.495 155.985 99.720 156.155 ;
        RECT 100.350 156.025 100.850 156.635 ;
        RECT 101.890 156.025 102.390 156.635 ;
        RECT 97.890 155.645 98.585 155.815 ;
        RECT 98.415 155.395 98.585 155.645 ;
        RECT 98.760 155.615 99.180 155.815 ;
        RECT 99.350 155.615 99.680 155.815 ;
        RECT 99.850 155.615 100.180 155.815 ;
        RECT 100.350 155.395 100.520 156.025 ;
        RECT 100.705 155.565 101.055 155.815 ;
        RECT 101.685 155.565 102.035 155.815 ;
        RECT 102.220 155.395 102.390 156.025 ;
        RECT 103.020 156.155 103.350 156.635 ;
        RECT 103.520 156.345 103.745 156.805 ;
        RECT 103.915 156.155 104.245 156.635 ;
        RECT 103.020 155.985 104.245 156.155 ;
        RECT 104.435 156.005 104.685 156.805 ;
        RECT 104.855 156.005 105.195 156.635 ;
        RECT 105.570 156.025 106.070 156.635 ;
        RECT 102.560 155.615 102.890 155.815 ;
        RECT 103.060 155.615 103.390 155.815 ;
        RECT 103.560 155.615 103.980 155.815 ;
        RECT 104.155 155.645 104.850 155.815 ;
        RECT 104.155 155.395 104.325 155.645 ;
        RECT 105.020 155.395 105.195 156.005 ;
        RECT 105.365 155.565 105.715 155.815 ;
        RECT 105.900 155.395 106.070 156.025 ;
        RECT 106.700 156.155 107.030 156.635 ;
        RECT 107.200 156.345 107.425 156.805 ;
        RECT 107.595 156.155 107.925 156.635 ;
        RECT 106.700 155.985 107.925 156.155 ;
        RECT 108.115 156.005 108.365 156.805 ;
        RECT 108.535 156.005 108.875 156.635 ;
        RECT 109.045 156.055 110.255 156.805 ;
        RECT 106.240 155.615 106.570 155.815 ;
        RECT 106.740 155.615 107.070 155.815 ;
        RECT 107.240 155.615 107.660 155.815 ;
        RECT 107.835 155.645 108.530 155.815 ;
        RECT 107.835 155.395 108.005 155.645 ;
        RECT 108.700 155.395 108.875 156.005 ;
        RECT 95.705 154.255 97.375 155.345 ;
        RECT 97.545 154.425 97.885 155.395 ;
        RECT 98.055 154.255 98.225 155.395 ;
        RECT 98.415 155.225 100.850 155.395 ;
        RECT 98.495 154.255 98.745 155.055 ;
        RECT 99.390 154.425 99.720 155.225 ;
        RECT 100.020 154.255 100.350 155.055 ;
        RECT 100.520 154.425 100.850 155.225 ;
        RECT 101.890 155.225 104.325 155.395 ;
        RECT 101.890 154.425 102.220 155.225 ;
        RECT 102.390 154.255 102.720 155.055 ;
        RECT 103.020 154.425 103.350 155.225 ;
        RECT 103.995 154.255 104.245 155.055 ;
        RECT 104.515 154.255 104.685 155.395 ;
        RECT 104.855 154.425 105.195 155.395 ;
        RECT 105.570 155.225 108.005 155.395 ;
        RECT 105.570 154.425 105.900 155.225 ;
        RECT 106.070 154.255 106.400 155.055 ;
        RECT 106.700 154.425 107.030 155.225 ;
        RECT 107.675 154.255 107.925 155.055 ;
        RECT 108.195 154.255 108.365 155.395 ;
        RECT 108.535 154.425 108.875 155.395 ;
        RECT 109.045 155.345 109.565 155.885 ;
        RECT 109.735 155.515 110.255 156.055 ;
        RECT 110.700 155.995 110.945 156.600 ;
        RECT 111.165 156.270 111.675 156.805 ;
        RECT 110.425 155.825 111.655 155.995 ;
        RECT 109.045 154.255 110.255 155.345 ;
        RECT 110.425 155.015 110.765 155.825 ;
        RECT 110.935 155.260 111.685 155.450 ;
        RECT 110.425 154.605 110.940 155.015 ;
        RECT 111.175 154.255 111.345 155.015 ;
        RECT 111.515 154.595 111.685 155.260 ;
        RECT 111.855 155.275 112.045 156.635 ;
        RECT 112.215 155.785 112.490 156.635 ;
        RECT 112.680 156.270 113.210 156.635 ;
        RECT 113.635 156.405 113.965 156.805 ;
        RECT 113.035 156.235 113.210 156.270 ;
        RECT 112.215 155.615 112.495 155.785 ;
        RECT 112.215 155.475 112.490 155.615 ;
        RECT 112.695 155.275 112.865 156.075 ;
        RECT 111.855 155.105 112.865 155.275 ;
        RECT 113.035 156.065 113.965 156.235 ;
        RECT 114.135 156.065 114.390 156.635 ;
        RECT 114.565 156.080 114.855 156.805 ;
        RECT 113.035 154.935 113.205 156.065 ;
        RECT 113.795 155.895 113.965 156.065 ;
        RECT 112.080 154.765 113.205 154.935 ;
        RECT 113.375 155.565 113.570 155.895 ;
        RECT 113.795 155.565 114.050 155.895 ;
        RECT 113.375 154.595 113.545 155.565 ;
        RECT 114.220 155.395 114.390 156.065 ;
        RECT 115.525 155.985 115.755 156.805 ;
        RECT 115.925 156.005 116.255 156.635 ;
        RECT 115.505 155.565 115.835 155.815 ;
        RECT 111.515 154.425 113.545 154.595 ;
        RECT 113.715 154.255 113.885 155.395 ;
        RECT 114.055 154.425 114.390 155.395 ;
        RECT 114.565 154.255 114.855 155.420 ;
        RECT 116.005 155.405 116.255 156.005 ;
        RECT 116.425 155.985 116.635 156.805 ;
        RECT 117.240 156.095 117.495 156.625 ;
        RECT 117.675 156.345 117.960 156.805 ;
        RECT 115.525 154.255 115.755 155.395 ;
        RECT 115.925 154.425 116.255 155.405 ;
        RECT 116.425 154.255 116.635 155.395 ;
        RECT 117.240 155.235 117.420 156.095 ;
        RECT 118.140 155.895 118.390 156.545 ;
        RECT 117.590 155.565 118.390 155.895 ;
        RECT 117.240 155.105 117.495 155.235 ;
        RECT 117.155 154.935 117.495 155.105 ;
        RECT 117.240 154.565 117.495 154.935 ;
        RECT 117.675 154.255 117.960 155.055 ;
        RECT 118.140 154.975 118.390 155.565 ;
        RECT 118.590 156.210 118.910 156.540 ;
        RECT 119.090 156.325 119.750 156.805 ;
        RECT 119.950 156.415 120.800 156.585 ;
        RECT 118.590 155.315 118.780 156.210 ;
        RECT 119.100 155.885 119.760 156.155 ;
        RECT 119.430 155.825 119.760 155.885 ;
        RECT 118.950 155.655 119.280 155.715 ;
        RECT 119.950 155.655 120.120 156.415 ;
        RECT 121.360 156.345 121.680 156.805 ;
        RECT 121.880 156.165 122.130 156.595 ;
        RECT 122.420 156.365 122.830 156.805 ;
        RECT 123.000 156.425 124.015 156.625 ;
        RECT 120.290 155.995 121.540 156.165 ;
        RECT 120.290 155.875 120.620 155.995 ;
        RECT 118.950 155.485 120.850 155.655 ;
        RECT 118.590 155.145 120.510 155.315 ;
        RECT 118.590 155.125 118.910 155.145 ;
        RECT 118.140 154.465 118.470 154.975 ;
        RECT 118.740 154.515 118.910 155.125 ;
        RECT 120.680 154.975 120.850 155.485 ;
        RECT 121.020 155.415 121.200 155.825 ;
        RECT 121.370 155.235 121.540 155.995 ;
        RECT 119.080 154.255 119.410 154.945 ;
        RECT 119.640 154.805 120.850 154.975 ;
        RECT 121.020 154.925 121.540 155.235 ;
        RECT 121.710 155.825 122.130 156.165 ;
        RECT 122.420 155.825 122.830 156.155 ;
        RECT 121.710 155.055 121.900 155.825 ;
        RECT 123.000 155.695 123.170 156.425 ;
        RECT 124.315 156.255 124.485 156.585 ;
        RECT 124.655 156.425 124.985 156.805 ;
        RECT 123.340 155.875 123.690 156.245 ;
        RECT 123.000 155.655 123.420 155.695 ;
        RECT 122.070 155.485 123.420 155.655 ;
        RECT 122.070 155.325 122.320 155.485 ;
        RECT 122.830 155.055 123.080 155.315 ;
        RECT 121.710 154.805 123.080 155.055 ;
        RECT 119.640 154.515 119.880 154.805 ;
        RECT 120.680 154.725 120.850 154.805 ;
        RECT 120.080 154.255 120.500 154.635 ;
        RECT 120.680 154.475 121.310 154.725 ;
        RECT 121.780 154.255 122.110 154.635 ;
        RECT 122.280 154.515 122.450 154.805 ;
        RECT 123.250 154.640 123.420 155.485 ;
        RECT 123.870 155.315 124.090 156.185 ;
        RECT 124.315 156.065 125.010 156.255 ;
        RECT 123.590 154.935 124.090 155.315 ;
        RECT 124.260 155.265 124.670 155.885 ;
        RECT 124.840 155.095 125.010 156.065 ;
        RECT 124.315 154.925 125.010 155.095 ;
        RECT 122.630 154.255 123.010 154.635 ;
        RECT 123.250 154.470 124.080 154.640 ;
        RECT 124.315 154.425 124.485 154.925 ;
        RECT 124.655 154.255 124.985 154.755 ;
        RECT 125.200 154.425 125.425 156.545 ;
        RECT 125.595 156.425 125.925 156.805 ;
        RECT 126.095 156.255 126.265 156.545 ;
        RECT 125.600 156.085 126.265 156.255 ;
        RECT 125.600 155.095 125.830 156.085 ;
        RECT 126.525 156.055 127.735 156.805 ;
        RECT 126.000 155.265 126.350 155.915 ;
        RECT 126.525 155.345 127.045 155.885 ;
        RECT 127.215 155.515 127.735 156.055 ;
        RECT 125.600 154.925 126.265 155.095 ;
        RECT 125.595 154.255 125.925 154.755 ;
        RECT 126.095 154.425 126.265 154.925 ;
        RECT 126.525 154.255 127.735 155.345 ;
        RECT 14.660 154.085 127.820 154.255 ;
        RECT 14.745 152.995 15.955 154.085 ;
        RECT 14.745 152.285 15.265 152.825 ;
        RECT 15.435 152.455 15.955 152.995 ;
        RECT 16.585 152.995 20.095 154.085 ;
        RECT 20.265 153.325 20.780 153.735 ;
        RECT 21.015 153.325 21.185 154.085 ;
        RECT 21.355 153.745 23.385 153.915 ;
        RECT 16.585 152.475 18.275 152.995 ;
        RECT 18.445 152.305 20.095 152.825 ;
        RECT 20.265 152.515 20.605 153.325 ;
        RECT 21.355 153.080 21.525 153.745 ;
        RECT 21.920 153.405 23.045 153.575 ;
        RECT 20.775 152.890 21.525 153.080 ;
        RECT 21.695 153.065 22.705 153.235 ;
        RECT 20.265 152.345 21.495 152.515 ;
        RECT 14.745 151.535 15.955 152.285 ;
        RECT 16.585 151.535 20.095 152.305 ;
        RECT 20.540 151.740 20.785 152.345 ;
        RECT 21.005 151.535 21.515 152.070 ;
        RECT 21.695 151.705 21.885 153.065 ;
        RECT 22.055 152.045 22.330 152.865 ;
        RECT 22.535 152.265 22.705 153.065 ;
        RECT 22.875 152.275 23.045 153.405 ;
        RECT 23.215 152.775 23.385 153.745 ;
        RECT 23.555 152.945 23.725 154.085 ;
        RECT 23.895 152.945 24.230 153.915 ;
        RECT 23.215 152.445 23.410 152.775 ;
        RECT 23.635 152.445 23.890 152.775 ;
        RECT 23.635 152.275 23.805 152.445 ;
        RECT 24.060 152.275 24.230 152.945 ;
        RECT 24.405 152.920 24.695 154.085 ;
        RECT 24.865 152.995 26.075 154.085 ;
        RECT 26.245 152.995 29.755 154.085 ;
        RECT 29.930 153.650 35.275 154.085 ;
        RECT 24.865 152.455 25.385 152.995 ;
        RECT 25.555 152.285 26.075 152.825 ;
        RECT 26.245 152.475 27.935 152.995 ;
        RECT 28.105 152.305 29.755 152.825 ;
        RECT 31.520 152.400 31.870 153.650 ;
        RECT 35.445 153.325 35.960 153.735 ;
        RECT 36.195 153.325 36.365 154.085 ;
        RECT 36.535 153.745 38.565 153.915 ;
        RECT 22.875 152.105 23.805 152.275 ;
        RECT 22.875 152.070 23.050 152.105 ;
        RECT 22.055 151.875 22.335 152.045 ;
        RECT 22.055 151.705 22.330 151.875 ;
        RECT 22.520 151.705 23.050 152.070 ;
        RECT 23.475 151.535 23.805 151.935 ;
        RECT 23.975 151.705 24.230 152.275 ;
        RECT 24.405 151.535 24.695 152.260 ;
        RECT 24.865 151.535 26.075 152.285 ;
        RECT 26.245 151.535 29.755 152.305 ;
        RECT 33.350 152.080 33.690 152.910 ;
        RECT 35.445 152.515 35.785 153.325 ;
        RECT 36.535 153.080 36.705 153.745 ;
        RECT 37.100 153.405 38.225 153.575 ;
        RECT 35.955 152.890 36.705 153.080 ;
        RECT 36.875 153.065 37.885 153.235 ;
        RECT 35.445 152.345 36.675 152.515 ;
        RECT 29.930 151.535 35.275 152.080 ;
        RECT 35.720 151.740 35.965 152.345 ;
        RECT 36.185 151.535 36.695 152.070 ;
        RECT 36.875 151.705 37.065 153.065 ;
        RECT 37.235 152.045 37.510 152.865 ;
        RECT 37.715 152.265 37.885 153.065 ;
        RECT 38.055 152.275 38.225 153.405 ;
        RECT 38.395 152.775 38.565 153.745 ;
        RECT 38.735 152.945 38.905 154.085 ;
        RECT 39.075 152.945 39.410 153.915 ;
        RECT 38.395 152.445 38.590 152.775 ;
        RECT 38.815 152.445 39.070 152.775 ;
        RECT 38.815 152.275 38.985 152.445 ;
        RECT 39.240 152.275 39.410 152.945 ;
        RECT 40.045 152.995 43.555 154.085 ;
        RECT 40.045 152.475 41.735 152.995 ;
        RECT 43.725 152.945 43.995 153.915 ;
        RECT 44.205 153.285 44.485 154.085 ;
        RECT 44.655 153.575 46.310 153.865 ;
        RECT 44.720 153.235 46.310 153.405 ;
        RECT 44.720 153.115 44.890 153.235 ;
        RECT 44.165 152.945 44.890 153.115 ;
        RECT 41.905 152.305 43.555 152.825 ;
        RECT 38.055 152.105 38.985 152.275 ;
        RECT 38.055 152.070 38.230 152.105 ;
        RECT 37.235 151.875 37.515 152.045 ;
        RECT 37.235 151.705 37.510 151.875 ;
        RECT 37.700 151.705 38.230 152.070 ;
        RECT 38.655 151.535 38.985 151.935 ;
        RECT 39.155 151.705 39.410 152.275 ;
        RECT 40.045 151.535 43.555 152.305 ;
        RECT 43.725 152.210 43.895 152.945 ;
        RECT 44.165 152.775 44.335 152.945 ;
        RECT 45.080 152.895 45.795 153.065 ;
        RECT 45.990 152.945 46.310 153.235 ;
        RECT 46.690 153.115 47.020 153.915 ;
        RECT 47.190 153.285 47.520 154.085 ;
        RECT 47.820 153.115 48.150 153.915 ;
        RECT 48.795 153.285 49.045 154.085 ;
        RECT 46.690 152.945 49.125 153.115 ;
        RECT 49.315 152.945 49.485 154.085 ;
        RECT 49.655 152.945 49.995 153.915 ;
        RECT 44.065 152.445 44.335 152.775 ;
        RECT 44.505 152.445 44.910 152.775 ;
        RECT 45.080 152.445 45.790 152.895 ;
        RECT 44.165 152.275 44.335 152.445 ;
        RECT 43.725 151.865 43.995 152.210 ;
        RECT 44.165 152.105 45.775 152.275 ;
        RECT 45.960 152.205 46.310 152.775 ;
        RECT 46.485 152.525 46.835 152.775 ;
        RECT 47.020 152.315 47.190 152.945 ;
        RECT 47.360 152.525 47.690 152.725 ;
        RECT 47.860 152.525 48.190 152.725 ;
        RECT 48.360 152.525 48.780 152.725 ;
        RECT 48.955 152.695 49.125 152.945 ;
        RECT 48.955 152.525 49.650 152.695 ;
        RECT 44.185 151.535 44.565 151.935 ;
        RECT 44.735 151.755 44.905 152.105 ;
        RECT 45.075 151.535 45.405 151.935 ;
        RECT 45.605 151.755 45.775 152.105 ;
        RECT 45.975 151.535 46.305 152.035 ;
        RECT 46.690 151.705 47.190 152.315 ;
        RECT 47.820 152.185 49.045 152.355 ;
        RECT 49.820 152.335 49.995 152.945 ;
        RECT 50.165 152.920 50.455 154.085 ;
        RECT 50.625 152.945 50.965 153.915 ;
        RECT 51.135 152.945 51.305 154.085 ;
        RECT 51.575 153.285 51.825 154.085 ;
        RECT 52.470 153.115 52.800 153.915 ;
        RECT 53.100 153.285 53.430 154.085 ;
        RECT 53.600 153.115 53.930 153.915 ;
        RECT 51.495 152.945 53.930 153.115 ;
        RECT 54.765 152.995 58.275 154.085 ;
        RECT 47.820 151.705 48.150 152.185 ;
        RECT 48.320 151.535 48.545 151.995 ;
        RECT 48.715 151.705 49.045 152.185 ;
        RECT 49.235 151.535 49.485 152.335 ;
        RECT 49.655 151.705 49.995 152.335 ;
        RECT 50.625 152.335 50.800 152.945 ;
        RECT 51.495 152.695 51.665 152.945 ;
        RECT 50.970 152.525 51.665 152.695 ;
        RECT 51.840 152.525 52.260 152.725 ;
        RECT 52.430 152.525 52.760 152.725 ;
        RECT 52.930 152.525 53.260 152.725 ;
        RECT 50.165 151.535 50.455 152.260 ;
        RECT 50.625 151.705 50.965 152.335 ;
        RECT 51.135 151.535 51.385 152.335 ;
        RECT 51.575 152.185 52.800 152.355 ;
        RECT 51.575 151.705 51.905 152.185 ;
        RECT 52.075 151.535 52.300 151.995 ;
        RECT 52.470 151.705 52.800 152.185 ;
        RECT 53.430 152.315 53.600 152.945 ;
        RECT 53.785 152.525 54.135 152.775 ;
        RECT 54.765 152.475 56.455 152.995 ;
        RECT 58.445 152.945 58.785 153.915 ;
        RECT 58.955 152.945 59.125 154.085 ;
        RECT 59.395 153.285 59.645 154.085 ;
        RECT 60.290 153.115 60.620 153.915 ;
        RECT 60.920 153.285 61.250 154.085 ;
        RECT 61.420 153.115 61.750 153.915 ;
        RECT 59.315 152.945 61.750 153.115 ;
        RECT 62.585 152.995 65.175 154.085 ;
        RECT 65.345 153.325 65.860 153.735 ;
        RECT 66.095 153.325 66.265 154.085 ;
        RECT 66.435 153.745 68.465 153.915 ;
        RECT 58.445 152.895 58.675 152.945 ;
        RECT 53.430 151.705 53.930 152.315 ;
        RECT 56.625 152.305 58.275 152.825 ;
        RECT 54.765 151.535 58.275 152.305 ;
        RECT 58.445 152.335 58.620 152.895 ;
        RECT 59.315 152.695 59.485 152.945 ;
        RECT 58.790 152.525 59.485 152.695 ;
        RECT 59.660 152.525 60.080 152.725 ;
        RECT 60.250 152.525 60.580 152.725 ;
        RECT 60.750 152.525 61.080 152.725 ;
        RECT 58.445 151.705 58.785 152.335 ;
        RECT 58.955 151.535 59.205 152.335 ;
        RECT 59.395 152.185 60.620 152.355 ;
        RECT 59.395 151.705 59.725 152.185 ;
        RECT 59.895 151.535 60.120 151.995 ;
        RECT 60.290 151.705 60.620 152.185 ;
        RECT 61.250 152.315 61.420 152.945 ;
        RECT 61.605 152.525 61.955 152.775 ;
        RECT 62.585 152.475 63.795 152.995 ;
        RECT 61.250 151.705 61.750 152.315 ;
        RECT 63.965 152.305 65.175 152.825 ;
        RECT 65.345 152.515 65.685 153.325 ;
        RECT 66.435 153.080 66.605 153.745 ;
        RECT 67.000 153.405 68.125 153.575 ;
        RECT 65.855 152.890 66.605 153.080 ;
        RECT 66.775 153.065 67.785 153.235 ;
        RECT 65.345 152.345 66.575 152.515 ;
        RECT 62.585 151.535 65.175 152.305 ;
        RECT 65.620 151.740 65.865 152.345 ;
        RECT 66.085 151.535 66.595 152.070 ;
        RECT 66.775 151.705 66.965 153.065 ;
        RECT 67.135 152.045 67.410 152.865 ;
        RECT 67.615 152.265 67.785 153.065 ;
        RECT 67.955 152.275 68.125 153.405 ;
        RECT 68.295 152.775 68.465 153.745 ;
        RECT 68.635 152.945 68.805 154.085 ;
        RECT 68.975 152.945 69.310 153.915 ;
        RECT 69.575 153.155 69.745 153.915 ;
        RECT 69.925 153.325 70.255 154.085 ;
        RECT 69.575 152.985 70.240 153.155 ;
        RECT 70.425 153.010 70.695 153.915 ;
        RECT 70.920 153.215 71.205 154.085 ;
        RECT 71.375 153.455 71.635 153.915 ;
        RECT 71.810 153.625 72.065 154.085 ;
        RECT 72.235 153.455 72.495 153.915 ;
        RECT 71.375 153.285 72.495 153.455 ;
        RECT 72.665 153.285 72.975 154.085 ;
        RECT 71.375 153.035 71.635 153.285 ;
        RECT 73.145 153.115 73.455 153.915 ;
        RECT 68.295 152.445 68.490 152.775 ;
        RECT 68.715 152.445 68.970 152.775 ;
        RECT 68.715 152.275 68.885 152.445 ;
        RECT 69.140 152.275 69.310 152.945 ;
        RECT 70.070 152.840 70.240 152.985 ;
        RECT 69.505 152.435 69.835 152.805 ;
        RECT 70.070 152.510 70.355 152.840 ;
        RECT 67.955 152.105 68.885 152.275 ;
        RECT 67.955 152.070 68.130 152.105 ;
        RECT 67.135 151.875 67.415 152.045 ;
        RECT 67.135 151.705 67.410 151.875 ;
        RECT 67.600 151.705 68.130 152.070 ;
        RECT 68.555 151.535 68.885 151.935 ;
        RECT 69.055 151.705 69.310 152.275 ;
        RECT 70.070 152.255 70.240 152.510 ;
        RECT 69.575 152.085 70.240 152.255 ;
        RECT 70.525 152.210 70.695 153.010 ;
        RECT 69.575 151.705 69.745 152.085 ;
        RECT 69.925 151.535 70.255 151.915 ;
        RECT 70.435 151.705 70.695 152.210 ;
        RECT 70.880 152.865 71.635 153.035 ;
        RECT 72.425 152.945 73.455 153.115 ;
        RECT 74.175 153.155 74.345 153.915 ;
        RECT 74.560 153.325 74.890 154.085 ;
        RECT 74.175 152.985 74.890 153.155 ;
        RECT 75.060 153.010 75.315 153.915 ;
        RECT 70.880 152.355 71.285 152.865 ;
        RECT 72.425 152.695 72.595 152.945 ;
        RECT 71.455 152.525 72.595 152.695 ;
        RECT 70.880 152.185 72.530 152.355 ;
        RECT 72.765 152.205 73.115 152.775 ;
        RECT 70.925 151.535 71.205 152.015 ;
        RECT 71.375 151.795 71.635 152.185 ;
        RECT 71.810 151.535 72.065 152.015 ;
        RECT 72.235 151.795 72.530 152.185 ;
        RECT 73.285 152.035 73.455 152.945 ;
        RECT 74.085 152.435 74.440 152.805 ;
        RECT 74.720 152.775 74.890 152.985 ;
        RECT 74.720 152.445 74.975 152.775 ;
        RECT 74.720 152.255 74.890 152.445 ;
        RECT 75.145 152.280 75.315 153.010 ;
        RECT 75.490 152.935 75.750 154.085 ;
        RECT 75.925 152.920 76.215 154.085 ;
        RECT 76.395 153.025 76.725 154.085 ;
        RECT 76.905 152.775 77.075 153.745 ;
        RECT 77.245 153.495 77.575 153.895 ;
        RECT 77.745 153.725 78.075 154.085 ;
        RECT 78.275 153.495 78.975 153.915 ;
        RECT 77.245 153.265 78.975 153.495 ;
        RECT 77.245 153.045 77.575 153.265 ;
        RECT 77.770 152.775 78.095 153.065 ;
        RECT 76.385 152.445 76.695 152.775 ;
        RECT 76.905 152.445 77.280 152.775 ;
        RECT 77.600 152.445 78.095 152.775 ;
        RECT 78.270 152.525 78.600 153.065 ;
        RECT 78.770 152.385 78.975 153.265 ;
        RECT 79.145 152.995 81.735 154.085 ;
        RECT 81.905 153.115 82.215 153.915 ;
        RECT 82.385 153.285 82.695 154.085 ;
        RECT 82.865 153.455 83.125 153.915 ;
        RECT 83.295 153.625 83.550 154.085 ;
        RECT 83.725 153.455 83.985 153.915 ;
        RECT 82.865 153.285 83.985 153.455 ;
        RECT 79.145 152.475 80.355 152.995 ;
        RECT 81.905 152.945 82.935 153.115 ;
        RECT 72.710 151.535 72.985 152.015 ;
        RECT 73.155 151.705 73.455 152.035 ;
        RECT 74.175 152.085 74.890 152.255 ;
        RECT 74.175 151.705 74.345 152.085 ;
        RECT 74.560 151.535 74.890 151.915 ;
        RECT 75.060 151.705 75.315 152.280 ;
        RECT 75.490 151.535 75.750 152.375 ;
        RECT 78.745 152.295 78.975 152.385 ;
        RECT 80.525 152.305 81.735 152.825 ;
        RECT 75.925 151.535 76.215 152.260 ;
        RECT 76.395 152.065 77.755 152.275 ;
        RECT 76.395 151.705 76.725 152.065 ;
        RECT 76.895 151.535 77.225 151.895 ;
        RECT 77.425 151.705 77.755 152.065 ;
        RECT 78.265 151.705 78.975 152.295 ;
        RECT 79.145 151.535 81.735 152.305 ;
        RECT 81.905 152.035 82.075 152.945 ;
        RECT 82.245 152.205 82.595 152.775 ;
        RECT 82.765 152.695 82.935 152.945 ;
        RECT 83.725 153.035 83.985 153.285 ;
        RECT 84.155 153.215 84.440 154.085 ;
        RECT 83.725 152.865 84.480 153.035 ;
        RECT 82.765 152.525 83.905 152.695 ;
        RECT 84.075 152.355 84.480 152.865 ;
        RECT 85.125 152.995 86.795 154.085 ;
        RECT 85.125 152.475 85.875 152.995 ;
        RECT 87.005 152.945 87.235 154.085 ;
        RECT 87.405 152.935 87.735 153.915 ;
        RECT 87.905 152.945 88.115 154.085 ;
        RECT 82.830 152.185 84.480 152.355 ;
        RECT 86.045 152.305 86.795 152.825 ;
        RECT 86.985 152.525 87.315 152.775 ;
        RECT 81.905 151.705 82.205 152.035 ;
        RECT 82.375 151.535 82.650 152.015 ;
        RECT 82.830 151.795 83.125 152.185 ;
        RECT 83.295 151.535 83.550 152.015 ;
        RECT 83.725 151.795 83.985 152.185 ;
        RECT 84.155 151.535 84.435 152.015 ;
        RECT 85.125 151.535 86.795 152.305 ;
        RECT 87.005 151.535 87.235 152.355 ;
        RECT 87.485 152.335 87.735 152.935 ;
        RECT 88.350 152.895 88.605 153.775 ;
        RECT 88.775 152.945 89.080 154.085 ;
        RECT 89.420 153.705 89.750 154.085 ;
        RECT 89.930 153.535 90.100 153.825 ;
        RECT 90.270 153.625 90.520 154.085 ;
        RECT 89.300 153.365 90.100 153.535 ;
        RECT 90.690 153.575 91.560 153.915 ;
        RECT 87.405 151.705 87.735 152.335 ;
        RECT 87.905 151.535 88.115 152.355 ;
        RECT 88.350 152.245 88.560 152.895 ;
        RECT 89.300 152.775 89.470 153.365 ;
        RECT 90.690 153.195 90.860 153.575 ;
        RECT 91.795 153.455 91.965 153.915 ;
        RECT 92.135 153.625 92.505 154.085 ;
        RECT 92.800 153.485 92.970 153.825 ;
        RECT 93.140 153.655 93.470 154.085 ;
        RECT 93.705 153.485 93.875 153.825 ;
        RECT 89.640 153.025 90.860 153.195 ;
        RECT 91.030 153.115 91.490 153.405 ;
        RECT 91.795 153.285 92.355 153.455 ;
        RECT 92.800 153.315 93.875 153.485 ;
        RECT 94.045 153.585 94.725 153.915 ;
        RECT 94.940 153.585 95.190 153.915 ;
        RECT 95.360 153.625 95.610 154.085 ;
        RECT 92.185 153.145 92.355 153.285 ;
        RECT 91.030 153.105 91.995 153.115 ;
        RECT 90.690 152.935 90.860 153.025 ;
        RECT 91.320 152.945 91.995 153.105 ;
        RECT 88.730 152.745 89.470 152.775 ;
        RECT 88.730 152.445 89.645 152.745 ;
        RECT 89.320 152.270 89.645 152.445 ;
        RECT 88.350 151.715 88.605 152.245 ;
        RECT 88.775 151.535 89.080 151.995 ;
        RECT 89.325 151.915 89.645 152.270 ;
        RECT 89.815 152.485 90.355 152.855 ;
        RECT 90.690 152.765 91.095 152.935 ;
        RECT 89.815 152.085 90.055 152.485 ;
        RECT 90.535 152.315 90.755 152.595 ;
        RECT 90.225 152.145 90.755 152.315 ;
        RECT 90.225 151.915 90.395 152.145 ;
        RECT 90.925 151.985 91.095 152.765 ;
        RECT 91.265 152.155 91.615 152.775 ;
        RECT 91.785 152.155 91.995 152.945 ;
        RECT 92.185 152.975 93.685 153.145 ;
        RECT 92.185 152.285 92.355 152.975 ;
        RECT 94.045 152.805 94.215 153.585 ;
        RECT 95.020 153.455 95.190 153.585 ;
        RECT 92.525 152.635 94.215 152.805 ;
        RECT 94.385 153.025 94.850 153.415 ;
        RECT 95.020 153.285 95.415 153.455 ;
        RECT 92.525 152.455 92.695 152.635 ;
        RECT 89.325 151.745 90.395 151.915 ;
        RECT 90.565 151.535 90.755 151.975 ;
        RECT 90.925 151.705 91.875 151.985 ;
        RECT 92.185 151.895 92.445 152.285 ;
        RECT 92.865 152.215 93.655 152.465 ;
        RECT 92.095 151.725 92.445 151.895 ;
        RECT 92.655 151.535 92.985 151.995 ;
        RECT 93.860 151.925 94.030 152.635 ;
        RECT 94.385 152.435 94.555 153.025 ;
        RECT 94.200 152.215 94.555 152.435 ;
        RECT 94.725 152.215 95.075 152.835 ;
        RECT 95.245 151.925 95.415 153.285 ;
        RECT 95.780 153.115 96.105 153.900 ;
        RECT 95.585 152.065 96.045 153.115 ;
        RECT 93.860 151.755 94.715 151.925 ;
        RECT 94.920 151.755 95.415 151.925 ;
        RECT 95.585 151.535 95.915 151.895 ;
        RECT 96.275 151.795 96.445 153.915 ;
        RECT 96.615 153.585 96.945 154.085 ;
        RECT 97.115 153.415 97.370 153.915 ;
        RECT 96.620 153.245 97.370 153.415 ;
        RECT 96.620 152.255 96.850 153.245 ;
        RECT 97.020 152.425 97.370 153.075 ;
        RECT 98.005 152.995 101.515 154.085 ;
        RECT 98.005 152.475 99.695 152.995 ;
        RECT 101.685 152.920 101.975 154.085 ;
        RECT 102.810 153.115 103.140 153.915 ;
        RECT 103.310 153.285 103.640 154.085 ;
        RECT 103.940 153.115 104.270 153.915 ;
        RECT 104.915 153.285 105.165 154.085 ;
        RECT 102.810 152.945 105.245 153.115 ;
        RECT 105.435 152.945 105.605 154.085 ;
        RECT 105.775 152.945 106.115 153.915 ;
        RECT 99.865 152.305 101.515 152.825 ;
        RECT 102.605 152.525 102.955 152.775 ;
        RECT 103.140 152.315 103.310 152.945 ;
        RECT 103.480 152.525 103.810 152.725 ;
        RECT 103.980 152.525 104.310 152.725 ;
        RECT 104.480 152.525 104.900 152.725 ;
        RECT 105.075 152.695 105.245 152.945 ;
        RECT 105.075 152.525 105.770 152.695 ;
        RECT 105.940 152.385 106.115 152.945 ;
        RECT 96.620 152.085 97.370 152.255 ;
        RECT 96.615 151.535 96.945 151.915 ;
        RECT 97.115 151.795 97.370 152.085 ;
        RECT 98.005 151.535 101.515 152.305 ;
        RECT 101.685 151.535 101.975 152.260 ;
        RECT 102.810 151.705 103.310 152.315 ;
        RECT 103.940 152.185 105.165 152.355 ;
        RECT 105.885 152.335 106.115 152.385 ;
        RECT 103.940 151.705 104.270 152.185 ;
        RECT 104.440 151.535 104.665 151.995 ;
        RECT 104.835 151.705 105.165 152.185 ;
        RECT 105.355 151.535 105.605 152.335 ;
        RECT 105.775 151.705 106.115 152.335 ;
        RECT 106.285 152.945 106.625 153.915 ;
        RECT 106.795 152.945 106.965 154.085 ;
        RECT 107.235 153.285 107.485 154.085 ;
        RECT 108.130 153.115 108.460 153.915 ;
        RECT 108.760 153.285 109.090 154.085 ;
        RECT 109.260 153.115 109.590 153.915 ;
        RECT 107.155 152.945 109.590 153.115 ;
        RECT 111.090 153.115 111.420 153.915 ;
        RECT 111.590 153.285 111.920 154.085 ;
        RECT 112.220 153.115 112.550 153.915 ;
        RECT 113.195 153.285 113.445 154.085 ;
        RECT 111.090 152.945 113.525 153.115 ;
        RECT 113.715 152.945 113.885 154.085 ;
        RECT 114.055 152.945 114.395 153.915 ;
        RECT 106.285 152.335 106.460 152.945 ;
        RECT 107.155 152.695 107.325 152.945 ;
        RECT 106.630 152.525 107.325 152.695 ;
        RECT 107.500 152.525 107.920 152.725 ;
        RECT 108.090 152.525 108.420 152.725 ;
        RECT 108.590 152.525 108.920 152.725 ;
        RECT 106.285 151.705 106.625 152.335 ;
        RECT 106.795 151.535 107.045 152.335 ;
        RECT 107.235 152.185 108.460 152.355 ;
        RECT 107.235 151.705 107.565 152.185 ;
        RECT 107.735 151.535 107.960 151.995 ;
        RECT 108.130 151.705 108.460 152.185 ;
        RECT 109.090 152.315 109.260 152.945 ;
        RECT 109.445 152.525 109.795 152.775 ;
        RECT 110.885 152.525 111.235 152.775 ;
        RECT 111.420 152.315 111.590 152.945 ;
        RECT 111.760 152.525 112.090 152.725 ;
        RECT 112.260 152.525 112.590 152.725 ;
        RECT 112.760 152.525 113.180 152.725 ;
        RECT 113.355 152.695 113.525 152.945 ;
        RECT 113.355 152.525 114.050 152.695 ;
        RECT 109.090 151.705 109.590 152.315 ;
        RECT 111.090 151.705 111.590 152.315 ;
        RECT 112.220 152.185 113.445 152.355 ;
        RECT 114.220 152.335 114.395 152.945 ;
        RECT 114.565 152.995 116.235 154.085 ;
        RECT 116.405 153.325 116.920 153.735 ;
        RECT 117.155 153.325 117.325 154.085 ;
        RECT 117.495 153.745 119.525 153.915 ;
        RECT 114.565 152.475 115.315 152.995 ;
        RECT 112.220 151.705 112.550 152.185 ;
        RECT 112.720 151.535 112.945 151.995 ;
        RECT 113.115 151.705 113.445 152.185 ;
        RECT 113.635 151.535 113.885 152.335 ;
        RECT 114.055 151.705 114.395 152.335 ;
        RECT 115.485 152.305 116.235 152.825 ;
        RECT 116.405 152.515 116.745 153.325 ;
        RECT 117.495 153.080 117.665 153.745 ;
        RECT 118.060 153.405 119.185 153.575 ;
        RECT 116.915 152.890 117.665 153.080 ;
        RECT 117.835 153.065 118.845 153.235 ;
        RECT 116.405 152.345 117.635 152.515 ;
        RECT 114.565 151.535 116.235 152.305 ;
        RECT 116.680 151.740 116.925 152.345 ;
        RECT 117.145 151.535 117.655 152.070 ;
        RECT 117.835 151.705 118.025 153.065 ;
        RECT 118.195 152.725 118.470 152.865 ;
        RECT 118.195 152.555 118.475 152.725 ;
        RECT 118.195 151.705 118.470 152.555 ;
        RECT 118.675 152.265 118.845 153.065 ;
        RECT 119.015 152.275 119.185 153.405 ;
        RECT 119.355 152.775 119.525 153.745 ;
        RECT 119.695 152.945 119.865 154.085 ;
        RECT 120.035 152.945 120.370 153.915 ;
        RECT 120.635 153.155 120.805 153.915 ;
        RECT 120.985 153.325 121.315 154.085 ;
        RECT 120.635 152.985 121.300 153.155 ;
        RECT 121.485 153.010 121.755 153.915 ;
        RECT 119.355 152.445 119.550 152.775 ;
        RECT 119.775 152.445 120.030 152.775 ;
        RECT 119.775 152.275 119.945 152.445 ;
        RECT 120.200 152.275 120.370 152.945 ;
        RECT 121.130 152.840 121.300 152.985 ;
        RECT 120.565 152.435 120.895 152.805 ;
        RECT 121.130 152.510 121.415 152.840 ;
        RECT 119.015 152.105 119.945 152.275 ;
        RECT 119.015 152.070 119.190 152.105 ;
        RECT 118.660 151.705 119.190 152.070 ;
        RECT 119.615 151.535 119.945 151.935 ;
        RECT 120.115 151.705 120.370 152.275 ;
        RECT 121.130 152.255 121.300 152.510 ;
        RECT 120.635 152.085 121.300 152.255 ;
        RECT 121.585 152.210 121.755 153.010 ;
        RECT 122.015 153.155 122.185 153.915 ;
        RECT 122.365 153.325 122.695 154.085 ;
        RECT 122.015 152.985 122.680 153.155 ;
        RECT 122.865 153.010 123.135 153.915 ;
        RECT 122.510 152.840 122.680 152.985 ;
        RECT 121.945 152.435 122.275 152.805 ;
        RECT 122.510 152.510 122.795 152.840 ;
        RECT 122.510 152.255 122.680 152.510 ;
        RECT 120.635 151.705 120.805 152.085 ;
        RECT 120.985 151.535 121.315 151.915 ;
        RECT 121.495 151.705 121.755 152.210 ;
        RECT 122.015 152.085 122.680 152.255 ;
        RECT 122.965 152.210 123.135 153.010 ;
        RECT 123.765 152.995 126.355 154.085 ;
        RECT 126.525 152.995 127.735 154.085 ;
        RECT 123.765 152.475 124.975 152.995 ;
        RECT 125.145 152.305 126.355 152.825 ;
        RECT 126.525 152.455 127.045 152.995 ;
        RECT 122.015 151.705 122.185 152.085 ;
        RECT 122.365 151.535 122.695 151.915 ;
        RECT 122.875 151.705 123.135 152.210 ;
        RECT 123.765 151.535 126.355 152.305 ;
        RECT 127.215 152.285 127.735 152.825 ;
        RECT 126.525 151.535 127.735 152.285 ;
        RECT 14.660 151.365 127.820 151.535 ;
        RECT 14.745 150.615 15.955 151.365 ;
        RECT 16.590 150.655 16.845 151.185 ;
        RECT 17.015 150.905 17.320 151.365 ;
        RECT 17.565 150.985 18.635 151.155 ;
        RECT 14.745 150.075 15.265 150.615 ;
        RECT 15.435 149.905 15.955 150.445 ;
        RECT 14.745 148.815 15.955 149.905 ;
        RECT 16.590 150.005 16.800 150.655 ;
        RECT 17.565 150.630 17.885 150.985 ;
        RECT 17.560 150.455 17.885 150.630 ;
        RECT 16.970 150.155 17.885 150.455 ;
        RECT 18.055 150.415 18.295 150.815 ;
        RECT 18.465 150.755 18.635 150.985 ;
        RECT 18.805 150.925 18.995 151.365 ;
        RECT 19.165 150.915 20.115 151.195 ;
        RECT 20.335 151.005 20.685 151.175 ;
        RECT 18.465 150.585 18.995 150.755 ;
        RECT 16.970 150.125 17.710 150.155 ;
        RECT 16.590 149.125 16.845 150.005 ;
        RECT 17.015 148.815 17.320 149.955 ;
        RECT 17.540 149.535 17.710 150.125 ;
        RECT 18.055 150.045 18.595 150.415 ;
        RECT 18.775 150.305 18.995 150.585 ;
        RECT 19.165 150.135 19.335 150.915 ;
        RECT 18.930 149.965 19.335 150.135 ;
        RECT 19.505 150.125 19.855 150.745 ;
        RECT 18.930 149.875 19.100 149.965 ;
        RECT 20.025 149.955 20.235 150.745 ;
        RECT 17.880 149.705 19.100 149.875 ;
        RECT 19.560 149.795 20.235 149.955 ;
        RECT 17.540 149.365 18.340 149.535 ;
        RECT 17.660 148.815 17.990 149.195 ;
        RECT 18.170 149.075 18.340 149.365 ;
        RECT 18.930 149.325 19.100 149.705 ;
        RECT 19.270 149.785 20.235 149.795 ;
        RECT 20.425 150.615 20.685 151.005 ;
        RECT 20.895 150.905 21.225 151.365 ;
        RECT 22.100 150.975 22.955 151.145 ;
        RECT 23.160 150.975 23.655 151.145 ;
        RECT 23.825 151.005 24.155 151.365 ;
        RECT 20.425 149.925 20.595 150.615 ;
        RECT 20.765 150.265 20.935 150.445 ;
        RECT 21.105 150.435 21.895 150.685 ;
        RECT 22.100 150.265 22.270 150.975 ;
        RECT 22.440 150.465 22.795 150.685 ;
        RECT 20.765 150.095 22.455 150.265 ;
        RECT 19.270 149.495 19.730 149.785 ;
        RECT 20.425 149.755 21.925 149.925 ;
        RECT 20.425 149.615 20.595 149.755 ;
        RECT 20.035 149.445 20.595 149.615 ;
        RECT 18.510 148.815 18.760 149.275 ;
        RECT 18.930 148.985 19.800 149.325 ;
        RECT 20.035 148.985 20.205 149.445 ;
        RECT 21.040 149.415 22.115 149.585 ;
        RECT 20.375 148.815 20.745 149.275 ;
        RECT 21.040 149.075 21.210 149.415 ;
        RECT 21.380 148.815 21.710 149.245 ;
        RECT 21.945 149.075 22.115 149.415 ;
        RECT 22.285 149.315 22.455 150.095 ;
        RECT 22.625 149.875 22.795 150.465 ;
        RECT 22.965 150.065 23.315 150.685 ;
        RECT 22.625 149.485 23.090 149.875 ;
        RECT 23.485 149.615 23.655 150.975 ;
        RECT 23.825 149.785 24.285 150.835 ;
        RECT 23.260 149.445 23.655 149.615 ;
        RECT 23.260 149.315 23.430 149.445 ;
        RECT 22.285 148.985 22.965 149.315 ;
        RECT 23.180 148.985 23.430 149.315 ;
        RECT 23.600 148.815 23.850 149.275 ;
        RECT 24.020 149.000 24.345 149.785 ;
        RECT 24.515 148.985 24.685 151.105 ;
        RECT 24.855 150.985 25.185 151.365 ;
        RECT 25.355 150.815 25.610 151.105 ;
        RECT 24.860 150.645 25.610 150.815 ;
        RECT 24.860 149.655 25.090 150.645 ;
        RECT 26.245 150.595 27.915 151.365 ;
        RECT 28.090 150.815 28.345 151.105 ;
        RECT 28.515 150.985 28.845 151.365 ;
        RECT 28.090 150.645 28.840 150.815 ;
        RECT 25.260 149.825 25.610 150.475 ;
        RECT 26.245 149.905 26.995 150.425 ;
        RECT 27.165 150.075 27.915 150.595 ;
        RECT 24.860 149.485 25.610 149.655 ;
        RECT 24.855 148.815 25.185 149.315 ;
        RECT 25.355 148.985 25.610 149.485 ;
        RECT 26.245 148.815 27.915 149.905 ;
        RECT 28.090 149.825 28.440 150.475 ;
        RECT 28.610 149.655 28.840 150.645 ;
        RECT 28.090 149.485 28.840 149.655 ;
        RECT 28.090 148.985 28.345 149.485 ;
        RECT 28.515 148.815 28.845 149.315 ;
        RECT 29.015 148.985 29.185 151.105 ;
        RECT 29.545 151.005 29.875 151.365 ;
        RECT 30.045 150.975 30.540 151.145 ;
        RECT 30.745 150.975 31.600 151.145 ;
        RECT 29.415 149.785 29.875 150.835 ;
        RECT 29.355 149.000 29.680 149.785 ;
        RECT 30.045 149.615 30.215 150.975 ;
        RECT 30.385 150.065 30.735 150.685 ;
        RECT 30.905 150.465 31.260 150.685 ;
        RECT 30.905 149.875 31.075 150.465 ;
        RECT 31.430 150.265 31.600 150.975 ;
        RECT 32.475 150.905 32.805 151.365 ;
        RECT 33.015 151.005 33.365 151.175 ;
        RECT 31.805 150.435 32.595 150.685 ;
        RECT 33.015 150.615 33.275 151.005 ;
        RECT 33.585 150.915 34.535 151.195 ;
        RECT 34.705 150.925 34.895 151.365 ;
        RECT 35.065 150.985 36.135 151.155 ;
        RECT 32.765 150.265 32.935 150.445 ;
        RECT 30.045 149.445 30.440 149.615 ;
        RECT 30.610 149.485 31.075 149.875 ;
        RECT 31.245 150.095 32.935 150.265 ;
        RECT 30.270 149.315 30.440 149.445 ;
        RECT 31.245 149.315 31.415 150.095 ;
        RECT 33.105 149.925 33.275 150.615 ;
        RECT 31.775 149.755 33.275 149.925 ;
        RECT 33.465 149.955 33.675 150.745 ;
        RECT 33.845 150.125 34.195 150.745 ;
        RECT 34.365 150.135 34.535 150.915 ;
        RECT 35.065 150.755 35.235 150.985 ;
        RECT 34.705 150.585 35.235 150.755 ;
        RECT 34.705 150.305 34.925 150.585 ;
        RECT 35.405 150.415 35.645 150.815 ;
        RECT 34.365 149.965 34.770 150.135 ;
        RECT 35.105 150.045 35.645 150.415 ;
        RECT 35.815 150.630 36.135 150.985 ;
        RECT 36.380 150.905 36.685 151.365 ;
        RECT 36.855 150.655 37.110 151.185 ;
        RECT 35.815 150.455 36.140 150.630 ;
        RECT 35.815 150.155 36.730 150.455 ;
        RECT 35.990 150.125 36.730 150.155 ;
        RECT 33.465 149.795 34.140 149.955 ;
        RECT 34.600 149.875 34.770 149.965 ;
        RECT 33.465 149.785 34.430 149.795 ;
        RECT 33.105 149.615 33.275 149.755 ;
        RECT 29.850 148.815 30.100 149.275 ;
        RECT 30.270 148.985 30.520 149.315 ;
        RECT 30.735 148.985 31.415 149.315 ;
        RECT 31.585 149.415 32.660 149.585 ;
        RECT 33.105 149.445 33.665 149.615 ;
        RECT 33.970 149.495 34.430 149.785 ;
        RECT 34.600 149.705 35.820 149.875 ;
        RECT 31.585 149.075 31.755 149.415 ;
        RECT 31.990 148.815 32.320 149.245 ;
        RECT 32.490 149.075 32.660 149.415 ;
        RECT 32.955 148.815 33.325 149.275 ;
        RECT 33.495 148.985 33.665 149.445 ;
        RECT 34.600 149.325 34.770 149.705 ;
        RECT 35.990 149.535 36.160 150.125 ;
        RECT 36.900 150.005 37.110 150.655 ;
        RECT 37.285 150.640 37.575 151.365 ;
        RECT 38.665 150.690 38.925 151.195 ;
        RECT 39.105 150.985 39.435 151.365 ;
        RECT 39.615 150.815 39.785 151.195 ;
        RECT 40.970 150.820 46.315 151.365 ;
        RECT 33.900 148.985 34.770 149.325 ;
        RECT 35.360 149.365 36.160 149.535 ;
        RECT 34.940 148.815 35.190 149.275 ;
        RECT 35.360 149.075 35.530 149.365 ;
        RECT 35.710 148.815 36.040 149.195 ;
        RECT 36.380 148.815 36.685 149.955 ;
        RECT 36.855 149.125 37.110 150.005 ;
        RECT 37.285 148.815 37.575 149.980 ;
        RECT 38.665 149.890 38.835 150.690 ;
        RECT 39.120 150.645 39.785 150.815 ;
        RECT 39.120 150.390 39.290 150.645 ;
        RECT 39.005 150.060 39.290 150.390 ;
        RECT 39.525 150.095 39.855 150.465 ;
        RECT 39.120 149.915 39.290 150.060 ;
        RECT 38.665 148.985 38.935 149.890 ;
        RECT 39.120 149.745 39.785 149.915 ;
        RECT 39.105 148.815 39.435 149.575 ;
        RECT 39.615 148.985 39.785 149.745 ;
        RECT 42.560 149.250 42.910 150.500 ;
        RECT 44.390 149.990 44.730 150.820 ;
        RECT 46.485 150.690 46.755 151.035 ;
        RECT 46.945 150.965 47.325 151.365 ;
        RECT 47.495 150.795 47.665 151.145 ;
        RECT 47.835 150.965 48.165 151.365 ;
        RECT 48.365 150.795 48.535 151.145 ;
        RECT 48.735 150.865 49.065 151.365 ;
        RECT 46.485 149.955 46.655 150.690 ;
        RECT 46.925 150.625 48.535 150.795 ;
        RECT 46.925 150.455 47.095 150.625 ;
        RECT 46.825 150.125 47.095 150.455 ;
        RECT 47.265 150.125 47.670 150.455 ;
        RECT 46.925 149.955 47.095 150.125 ;
        RECT 47.840 150.005 48.550 150.455 ;
        RECT 48.720 150.125 49.070 150.695 ;
        RECT 49.245 150.690 49.515 151.035 ;
        RECT 49.705 150.965 50.085 151.365 ;
        RECT 50.255 150.795 50.425 151.145 ;
        RECT 50.595 150.965 50.925 151.365 ;
        RECT 51.125 150.795 51.295 151.145 ;
        RECT 51.495 150.865 51.825 151.365 ;
        RECT 40.970 148.815 46.315 149.250 ;
        RECT 46.485 148.985 46.755 149.955 ;
        RECT 46.925 149.785 47.650 149.955 ;
        RECT 47.840 149.835 48.555 150.005 ;
        RECT 49.245 149.955 49.415 150.690 ;
        RECT 49.685 150.625 51.295 150.795 ;
        RECT 49.685 150.455 49.855 150.625 ;
        RECT 49.585 150.125 49.855 150.455 ;
        RECT 50.025 150.125 50.430 150.455 ;
        RECT 49.685 149.955 49.855 150.125 ;
        RECT 50.600 150.005 51.310 150.455 ;
        RECT 51.480 150.125 51.830 150.695 ;
        RECT 52.005 150.595 54.595 151.365 ;
        RECT 47.480 149.665 47.650 149.785 ;
        RECT 48.750 149.665 49.070 149.955 ;
        RECT 46.965 148.815 47.245 149.615 ;
        RECT 47.480 149.495 49.070 149.665 ;
        RECT 47.415 149.035 49.070 149.325 ;
        RECT 49.245 148.985 49.515 149.955 ;
        RECT 49.685 149.785 50.410 149.955 ;
        RECT 50.600 149.835 51.315 150.005 ;
        RECT 50.240 149.665 50.410 149.785 ;
        RECT 51.510 149.665 51.830 149.955 ;
        RECT 49.725 148.815 50.005 149.615 ;
        RECT 50.240 149.495 51.830 149.665 ;
        RECT 52.005 149.905 53.215 150.425 ;
        RECT 53.385 150.075 54.595 150.595 ;
        RECT 54.765 150.565 55.105 151.195 ;
        RECT 55.275 150.565 55.525 151.365 ;
        RECT 55.715 150.715 56.045 151.195 ;
        RECT 56.215 150.905 56.440 151.365 ;
        RECT 56.610 150.715 56.940 151.195 ;
        RECT 54.765 149.955 54.940 150.565 ;
        RECT 55.715 150.545 56.940 150.715 ;
        RECT 57.570 150.585 58.070 151.195 ;
        RECT 55.110 150.205 55.805 150.375 ;
        RECT 55.635 149.955 55.805 150.205 ;
        RECT 55.980 150.175 56.400 150.375 ;
        RECT 56.570 150.175 56.900 150.375 ;
        RECT 57.070 150.175 57.400 150.375 ;
        RECT 57.570 149.955 57.740 150.585 ;
        RECT 58.445 150.565 58.785 151.195 ;
        RECT 58.955 150.565 59.205 151.365 ;
        RECT 59.395 150.715 59.725 151.195 ;
        RECT 59.895 150.905 60.120 151.365 ;
        RECT 60.290 150.715 60.620 151.195 ;
        RECT 58.445 150.515 58.675 150.565 ;
        RECT 59.395 150.545 60.620 150.715 ;
        RECT 61.250 150.585 61.750 151.195 ;
        RECT 63.045 150.640 63.335 151.365 ;
        RECT 63.595 150.885 63.895 151.365 ;
        RECT 64.065 150.715 64.325 151.170 ;
        RECT 64.495 150.885 64.755 151.365 ;
        RECT 64.935 150.715 65.195 151.170 ;
        RECT 65.365 150.885 65.615 151.365 ;
        RECT 65.795 150.715 66.055 151.170 ;
        RECT 66.225 150.885 66.475 151.365 ;
        RECT 66.655 150.715 66.915 151.170 ;
        RECT 67.085 150.885 67.330 151.365 ;
        RECT 67.500 150.715 67.775 151.170 ;
        RECT 67.945 150.885 68.190 151.365 ;
        RECT 68.360 150.715 68.620 151.170 ;
        RECT 68.790 150.885 69.050 151.365 ;
        RECT 69.220 150.715 69.480 151.170 ;
        RECT 69.650 150.885 69.910 151.365 ;
        RECT 70.080 150.715 70.340 151.170 ;
        RECT 70.510 150.805 70.770 151.365 ;
        RECT 57.925 150.125 58.275 150.375 ;
        RECT 58.445 149.955 58.620 150.515 ;
        RECT 58.790 150.205 59.485 150.375 ;
        RECT 59.315 149.955 59.485 150.205 ;
        RECT 59.660 150.175 60.080 150.375 ;
        RECT 60.250 150.175 60.580 150.375 ;
        RECT 60.750 150.175 61.080 150.375 ;
        RECT 61.250 149.955 61.420 150.585 ;
        RECT 63.595 150.545 70.340 150.715 ;
        RECT 61.605 150.125 61.955 150.375 ;
        RECT 50.175 149.035 51.830 149.325 ;
        RECT 52.005 148.815 54.595 149.905 ;
        RECT 54.765 148.985 55.105 149.955 ;
        RECT 55.275 148.815 55.445 149.955 ;
        RECT 55.635 149.785 58.070 149.955 ;
        RECT 55.715 148.815 55.965 149.615 ;
        RECT 56.610 148.985 56.940 149.785 ;
        RECT 57.240 148.815 57.570 149.615 ;
        RECT 57.740 148.985 58.070 149.785 ;
        RECT 58.445 148.985 58.785 149.955 ;
        RECT 58.955 148.815 59.125 149.955 ;
        RECT 59.315 149.785 61.750 149.955 ;
        RECT 59.395 148.815 59.645 149.615 ;
        RECT 60.290 148.985 60.620 149.785 ;
        RECT 60.920 148.815 61.250 149.615 ;
        RECT 61.420 148.985 61.750 149.785 ;
        RECT 63.045 148.815 63.335 149.980 ;
        RECT 63.595 149.955 64.760 150.545 ;
        RECT 70.940 150.375 71.190 151.185 ;
        RECT 71.370 150.840 71.630 151.365 ;
        RECT 71.800 150.375 72.050 151.185 ;
        RECT 72.230 150.855 72.535 151.365 ;
        RECT 64.930 150.125 72.050 150.375 ;
        RECT 72.220 150.125 72.535 150.685 ;
        RECT 72.710 150.525 72.970 151.365 ;
        RECT 73.145 150.620 73.400 151.195 ;
        RECT 73.570 150.985 73.900 151.365 ;
        RECT 74.115 150.815 74.285 151.195 ;
        RECT 73.570 150.645 74.285 150.815 ;
        RECT 63.595 149.730 70.340 149.955 ;
        RECT 63.595 148.815 63.865 149.560 ;
        RECT 64.035 148.990 64.325 149.730 ;
        RECT 64.935 149.715 70.340 149.730 ;
        RECT 64.495 148.820 64.750 149.545 ;
        RECT 64.935 148.990 65.195 149.715 ;
        RECT 65.365 148.820 65.610 149.545 ;
        RECT 65.795 148.990 66.055 149.715 ;
        RECT 66.225 148.820 66.470 149.545 ;
        RECT 66.655 148.990 66.915 149.715 ;
        RECT 67.085 148.820 67.330 149.545 ;
        RECT 67.500 148.990 67.760 149.715 ;
        RECT 67.930 148.820 68.190 149.545 ;
        RECT 68.360 148.990 68.620 149.715 ;
        RECT 68.790 148.820 69.050 149.545 ;
        RECT 69.220 148.990 69.480 149.715 ;
        RECT 69.650 148.820 69.910 149.545 ;
        RECT 70.080 148.990 70.340 149.715 ;
        RECT 70.510 148.820 70.770 149.615 ;
        RECT 70.940 148.990 71.190 150.125 ;
        RECT 64.495 148.815 70.770 148.820 ;
        RECT 71.370 148.815 71.630 149.625 ;
        RECT 71.805 148.985 72.050 150.125 ;
        RECT 72.230 148.815 72.525 149.625 ;
        RECT 72.710 148.815 72.970 149.965 ;
        RECT 73.145 149.890 73.315 150.620 ;
        RECT 73.570 150.455 73.740 150.645 ;
        RECT 74.550 150.525 74.810 151.365 ;
        RECT 74.985 150.620 75.240 151.195 ;
        RECT 75.410 150.985 75.740 151.365 ;
        RECT 75.955 150.815 76.125 151.195 ;
        RECT 75.410 150.645 76.125 150.815 ;
        RECT 73.485 150.125 73.740 150.455 ;
        RECT 73.570 149.915 73.740 150.125 ;
        RECT 74.020 150.095 74.375 150.465 ;
        RECT 73.145 148.985 73.400 149.890 ;
        RECT 73.570 149.745 74.285 149.915 ;
        RECT 73.570 148.815 73.900 149.575 ;
        RECT 74.115 148.985 74.285 149.745 ;
        RECT 74.550 148.815 74.810 149.965 ;
        RECT 74.985 149.890 75.155 150.620 ;
        RECT 75.410 150.455 75.580 150.645 ;
        RECT 77.050 150.585 77.550 151.195 ;
        RECT 75.325 150.125 75.580 150.455 ;
        RECT 75.410 149.915 75.580 150.125 ;
        RECT 75.860 150.095 76.215 150.465 ;
        RECT 76.845 150.125 77.195 150.375 ;
        RECT 77.380 149.955 77.550 150.585 ;
        RECT 78.180 150.715 78.510 151.195 ;
        RECT 78.680 150.905 78.905 151.365 ;
        RECT 79.075 150.715 79.405 151.195 ;
        RECT 78.180 150.545 79.405 150.715 ;
        RECT 79.595 150.565 79.845 151.365 ;
        RECT 80.015 150.565 80.355 151.195 ;
        RECT 77.720 150.175 78.050 150.375 ;
        RECT 78.220 150.175 78.550 150.375 ;
        RECT 78.720 150.175 79.140 150.375 ;
        RECT 79.315 150.205 80.010 150.375 ;
        RECT 79.315 149.955 79.485 150.205 ;
        RECT 80.180 149.955 80.355 150.565 ;
        RECT 74.985 148.985 75.240 149.890 ;
        RECT 75.410 149.745 76.125 149.915 ;
        RECT 75.410 148.815 75.740 149.575 ;
        RECT 75.955 148.985 76.125 149.745 ;
        RECT 77.050 149.785 79.485 149.955 ;
        RECT 77.050 148.985 77.380 149.785 ;
        RECT 77.550 148.815 77.880 149.615 ;
        RECT 78.180 148.985 78.510 149.785 ;
        RECT 79.155 148.815 79.405 149.615 ;
        RECT 79.675 148.815 79.845 149.955 ;
        RECT 80.015 148.985 80.355 149.955 ;
        RECT 80.525 150.565 80.865 151.195 ;
        RECT 81.035 150.565 81.285 151.365 ;
        RECT 81.475 150.715 81.805 151.195 ;
        RECT 81.975 150.905 82.200 151.365 ;
        RECT 82.370 150.715 82.700 151.195 ;
        RECT 80.525 149.955 80.700 150.565 ;
        RECT 81.475 150.545 82.700 150.715 ;
        RECT 83.330 150.585 83.830 151.195 ;
        RECT 85.125 150.595 88.635 151.365 ;
        RECT 88.805 150.640 89.095 151.365 ;
        RECT 80.870 150.205 81.565 150.375 ;
        RECT 81.395 149.955 81.565 150.205 ;
        RECT 81.740 150.175 82.160 150.375 ;
        RECT 82.330 150.175 82.660 150.375 ;
        RECT 82.830 150.175 83.160 150.375 ;
        RECT 83.330 149.955 83.500 150.585 ;
        RECT 83.685 150.125 84.035 150.375 ;
        RECT 80.525 148.985 80.865 149.955 ;
        RECT 81.035 148.815 81.205 149.955 ;
        RECT 81.395 149.785 83.830 149.955 ;
        RECT 81.475 148.815 81.725 149.615 ;
        RECT 82.370 148.985 82.700 149.785 ;
        RECT 83.000 148.815 83.330 149.615 ;
        RECT 83.500 148.985 83.830 149.785 ;
        RECT 85.125 149.905 86.815 150.425 ;
        RECT 86.985 150.075 88.635 150.595 ;
        RECT 89.540 150.555 89.785 151.160 ;
        RECT 90.005 150.830 90.515 151.365 ;
        RECT 89.265 150.385 90.495 150.555 ;
        RECT 85.125 148.815 88.635 149.905 ;
        RECT 88.805 148.815 89.095 149.980 ;
        RECT 89.265 149.575 89.605 150.385 ;
        RECT 89.775 149.820 90.525 150.010 ;
        RECT 89.265 149.165 89.780 149.575 ;
        RECT 90.015 148.815 90.185 149.575 ;
        RECT 90.355 149.155 90.525 149.820 ;
        RECT 90.695 149.835 90.885 151.195 ;
        RECT 91.055 150.345 91.330 151.195 ;
        RECT 91.520 150.830 92.050 151.195 ;
        RECT 92.475 150.965 92.805 151.365 ;
        RECT 91.875 150.795 92.050 150.830 ;
        RECT 91.055 150.175 91.335 150.345 ;
        RECT 91.055 150.035 91.330 150.175 ;
        RECT 91.535 149.835 91.705 150.635 ;
        RECT 90.695 149.665 91.705 149.835 ;
        RECT 91.875 150.625 92.805 150.795 ;
        RECT 92.975 150.625 93.230 151.195 ;
        RECT 91.875 149.495 92.045 150.625 ;
        RECT 92.635 150.455 92.805 150.625 ;
        RECT 90.920 149.325 92.045 149.495 ;
        RECT 92.215 150.125 92.410 150.455 ;
        RECT 92.635 150.125 92.890 150.455 ;
        RECT 92.215 149.155 92.385 150.125 ;
        RECT 93.060 149.955 93.230 150.625 ;
        RECT 93.405 150.615 94.615 151.365 ;
        RECT 90.355 148.985 92.385 149.155 ;
        RECT 92.555 148.815 92.725 149.955 ;
        RECT 92.895 148.985 93.230 149.955 ;
        RECT 93.405 149.905 93.925 150.445 ;
        RECT 94.095 150.075 94.615 150.615 ;
        RECT 94.785 150.595 98.295 151.365 ;
        RECT 98.470 150.820 103.815 151.365 ;
        RECT 103.995 150.865 104.325 151.365 ;
        RECT 94.785 149.905 96.475 150.425 ;
        RECT 96.645 150.075 98.295 150.595 ;
        RECT 93.405 148.815 94.615 149.905 ;
        RECT 94.785 148.815 98.295 149.905 ;
        RECT 100.060 149.250 100.410 150.500 ;
        RECT 101.890 149.990 102.230 150.820 ;
        RECT 104.525 150.795 104.695 151.145 ;
        RECT 104.895 150.965 105.225 151.365 ;
        RECT 105.395 150.795 105.565 151.145 ;
        RECT 105.735 150.965 106.115 151.365 ;
        RECT 103.990 150.125 104.340 150.695 ;
        RECT 104.525 150.625 106.135 150.795 ;
        RECT 106.305 150.690 106.575 151.035 ;
        RECT 105.965 150.455 106.135 150.625 ;
        RECT 104.510 150.005 105.220 150.455 ;
        RECT 105.390 150.125 105.795 150.455 ;
        RECT 105.965 150.125 106.235 150.455 ;
        RECT 103.990 149.665 104.310 149.955 ;
        RECT 104.505 149.835 105.220 150.005 ;
        RECT 105.965 149.955 106.135 150.125 ;
        RECT 106.405 149.955 106.575 150.690 ;
        RECT 106.745 150.595 109.335 151.365 ;
        RECT 109.515 150.865 109.845 151.365 ;
        RECT 110.045 150.795 110.215 151.145 ;
        RECT 110.415 150.965 110.745 151.365 ;
        RECT 110.915 150.795 111.085 151.145 ;
        RECT 111.255 150.965 111.635 151.365 ;
        RECT 105.410 149.785 106.135 149.955 ;
        RECT 105.410 149.665 105.580 149.785 ;
        RECT 103.990 149.495 105.580 149.665 ;
        RECT 98.470 148.815 103.815 149.250 ;
        RECT 103.990 149.035 105.645 149.325 ;
        RECT 105.815 148.815 106.095 149.615 ;
        RECT 106.305 148.985 106.575 149.955 ;
        RECT 106.745 149.905 107.955 150.425 ;
        RECT 108.125 150.075 109.335 150.595 ;
        RECT 109.510 150.125 109.860 150.695 ;
        RECT 110.045 150.625 111.655 150.795 ;
        RECT 111.825 150.690 112.095 151.035 ;
        RECT 111.485 150.455 111.655 150.625 ;
        RECT 106.745 148.815 109.335 149.905 ;
        RECT 109.510 149.665 109.830 149.955 ;
        RECT 110.030 149.835 110.740 150.455 ;
        RECT 110.910 150.125 111.315 150.455 ;
        RECT 111.485 150.125 111.755 150.455 ;
        RECT 111.485 149.955 111.655 150.125 ;
        RECT 111.925 149.955 112.095 150.690 ;
        RECT 112.725 150.595 114.395 151.365 ;
        RECT 114.565 150.640 114.855 151.365 ;
        RECT 115.490 150.820 120.835 151.365 ;
        RECT 121.010 150.820 126.355 151.365 ;
        RECT 110.930 149.785 111.655 149.955 ;
        RECT 110.930 149.665 111.100 149.785 ;
        RECT 109.510 149.495 111.100 149.665 ;
        RECT 109.510 149.035 111.165 149.325 ;
        RECT 111.335 148.815 111.615 149.615 ;
        RECT 111.825 148.985 112.095 149.955 ;
        RECT 112.725 149.905 113.475 150.425 ;
        RECT 113.645 150.075 114.395 150.595 ;
        RECT 112.725 148.815 114.395 149.905 ;
        RECT 114.565 148.815 114.855 149.980 ;
        RECT 117.080 149.250 117.430 150.500 ;
        RECT 118.910 149.990 119.250 150.820 ;
        RECT 122.600 149.250 122.950 150.500 ;
        RECT 124.430 149.990 124.770 150.820 ;
        RECT 126.525 150.615 127.735 151.365 ;
        RECT 126.525 149.905 127.045 150.445 ;
        RECT 127.215 150.075 127.735 150.615 ;
        RECT 115.490 148.815 120.835 149.250 ;
        RECT 121.010 148.815 126.355 149.250 ;
        RECT 126.525 148.815 127.735 149.905 ;
        RECT 14.660 148.645 127.820 148.815 ;
        RECT 14.745 147.555 15.955 148.645 ;
        RECT 14.745 146.845 15.265 147.385 ;
        RECT 15.435 147.015 15.955 147.555 ;
        RECT 16.125 147.555 18.715 148.645 ;
        RECT 16.125 147.035 17.335 147.555 ;
        RECT 18.945 147.505 19.155 148.645 ;
        RECT 19.325 147.495 19.655 148.475 ;
        RECT 19.825 147.505 20.055 148.645 ;
        RECT 20.265 147.885 20.780 148.295 ;
        RECT 21.015 147.885 21.185 148.645 ;
        RECT 21.355 148.305 23.385 148.475 ;
        RECT 17.505 146.865 18.715 147.385 ;
        RECT 14.745 146.095 15.955 146.845 ;
        RECT 16.125 146.095 18.715 146.865 ;
        RECT 18.945 146.095 19.155 146.915 ;
        RECT 19.325 146.895 19.575 147.495 ;
        RECT 19.745 147.085 20.075 147.335 ;
        RECT 20.265 147.075 20.605 147.885 ;
        RECT 21.355 147.640 21.525 148.305 ;
        RECT 21.920 147.965 23.045 148.135 ;
        RECT 20.775 147.450 21.525 147.640 ;
        RECT 21.695 147.625 22.705 147.795 ;
        RECT 19.325 146.265 19.655 146.895 ;
        RECT 19.825 146.095 20.055 146.915 ;
        RECT 20.265 146.905 21.495 147.075 ;
        RECT 20.540 146.300 20.785 146.905 ;
        RECT 21.005 146.095 21.515 146.630 ;
        RECT 21.695 146.265 21.885 147.625 ;
        RECT 22.055 146.945 22.330 147.425 ;
        RECT 22.055 146.775 22.335 146.945 ;
        RECT 22.535 146.825 22.705 147.625 ;
        RECT 22.875 146.835 23.045 147.965 ;
        RECT 23.215 147.335 23.385 148.305 ;
        RECT 23.555 147.505 23.725 148.645 ;
        RECT 23.895 147.505 24.230 148.475 ;
        RECT 23.215 147.005 23.410 147.335 ;
        RECT 23.635 147.005 23.890 147.335 ;
        RECT 23.635 146.835 23.805 147.005 ;
        RECT 24.060 146.835 24.230 147.505 ;
        RECT 24.405 147.480 24.695 148.645 ;
        RECT 25.325 147.555 26.995 148.645 ;
        RECT 27.170 148.210 32.515 148.645 ;
        RECT 25.325 147.035 26.075 147.555 ;
        RECT 26.245 146.865 26.995 147.385 ;
        RECT 28.760 146.960 29.110 148.210 ;
        RECT 32.725 147.505 32.955 148.645 ;
        RECT 33.125 147.495 33.455 148.475 ;
        RECT 33.625 147.505 33.835 148.645 ;
        RECT 34.155 147.715 34.325 148.475 ;
        RECT 34.505 147.885 34.835 148.645 ;
        RECT 34.155 147.545 34.820 147.715 ;
        RECT 35.005 147.570 35.275 148.475 ;
        RECT 36.370 148.210 41.715 148.645 ;
        RECT 22.055 146.265 22.330 146.775 ;
        RECT 22.875 146.665 23.805 146.835 ;
        RECT 22.875 146.630 23.050 146.665 ;
        RECT 22.520 146.265 23.050 146.630 ;
        RECT 23.475 146.095 23.805 146.495 ;
        RECT 23.975 146.265 24.230 146.835 ;
        RECT 24.405 146.095 24.695 146.820 ;
        RECT 25.325 146.095 26.995 146.865 ;
        RECT 30.590 146.640 30.930 147.470 ;
        RECT 32.705 147.085 33.035 147.335 ;
        RECT 27.170 146.095 32.515 146.640 ;
        RECT 32.725 146.095 32.955 146.915 ;
        RECT 33.205 146.895 33.455 147.495 ;
        RECT 34.650 147.400 34.820 147.545 ;
        RECT 34.085 146.995 34.415 147.365 ;
        RECT 34.650 147.070 34.935 147.400 ;
        RECT 33.125 146.265 33.455 146.895 ;
        RECT 33.625 146.095 33.835 146.915 ;
        RECT 34.650 146.815 34.820 147.070 ;
        RECT 34.155 146.645 34.820 146.815 ;
        RECT 35.105 146.770 35.275 147.570 ;
        RECT 37.960 146.960 38.310 148.210 ;
        RECT 41.895 147.665 42.225 148.475 ;
        RECT 42.395 147.845 42.635 148.645 ;
        RECT 41.895 147.495 42.610 147.665 ;
        RECT 34.155 146.265 34.325 146.645 ;
        RECT 34.505 146.095 34.835 146.475 ;
        RECT 35.015 146.265 35.275 146.770 ;
        RECT 39.790 146.640 40.130 147.470 ;
        RECT 41.890 147.085 42.270 147.325 ;
        RECT 42.440 147.255 42.610 147.495 ;
        RECT 42.815 147.625 42.985 148.475 ;
        RECT 43.155 147.845 43.485 148.645 ;
        RECT 43.655 147.625 43.825 148.475 ;
        RECT 42.815 147.455 43.825 147.625 ;
        RECT 43.995 147.495 44.325 148.645 ;
        RECT 44.650 148.210 49.995 148.645 ;
        RECT 42.440 147.085 42.940 147.255 ;
        RECT 42.440 146.915 42.610 147.085 ;
        RECT 43.330 146.945 43.825 147.455 ;
        RECT 46.240 146.960 46.590 148.210 ;
        RECT 50.165 147.480 50.455 148.645 ;
        RECT 51.085 147.555 54.595 148.645 ;
        RECT 54.770 148.210 60.115 148.645 ;
        RECT 43.325 146.915 43.825 146.945 ;
        RECT 41.975 146.745 42.610 146.915 ;
        RECT 42.815 146.745 43.825 146.915 ;
        RECT 36.370 146.095 41.715 146.640 ;
        RECT 41.975 146.265 42.145 146.745 ;
        RECT 42.325 146.095 42.565 146.575 ;
        RECT 42.815 146.265 42.985 146.745 ;
        RECT 43.155 146.095 43.485 146.575 ;
        RECT 43.655 146.265 43.825 146.745 ;
        RECT 43.995 146.095 44.325 146.895 ;
        RECT 48.070 146.640 48.410 147.470 ;
        RECT 51.085 147.035 52.775 147.555 ;
        RECT 52.945 146.865 54.595 147.385 ;
        RECT 56.360 146.960 56.710 148.210 ;
        RECT 60.345 147.505 60.555 148.645 ;
        RECT 60.725 147.495 61.055 148.475 ;
        RECT 61.225 147.505 61.455 148.645 ;
        RECT 62.125 147.555 64.715 148.645 ;
        RECT 64.885 147.570 65.155 148.475 ;
        RECT 65.325 147.885 65.655 148.645 ;
        RECT 65.835 147.715 66.005 148.475 ;
        RECT 44.650 146.095 49.995 146.640 ;
        RECT 50.165 146.095 50.455 146.820 ;
        RECT 51.085 146.095 54.595 146.865 ;
        RECT 58.190 146.640 58.530 147.470 ;
        RECT 54.770 146.095 60.115 146.640 ;
        RECT 60.345 146.095 60.555 146.915 ;
        RECT 60.725 146.895 60.975 147.495 ;
        RECT 61.145 147.085 61.475 147.335 ;
        RECT 62.125 147.035 63.335 147.555 ;
        RECT 60.725 146.265 61.055 146.895 ;
        RECT 61.225 146.095 61.455 146.915 ;
        RECT 63.505 146.865 64.715 147.385 ;
        RECT 62.125 146.095 64.715 146.865 ;
        RECT 64.885 146.770 65.055 147.570 ;
        RECT 65.340 147.545 66.005 147.715 ;
        RECT 66.265 147.555 67.475 148.645 ;
        RECT 67.645 147.555 71.155 148.645 ;
        RECT 71.415 147.715 71.585 148.475 ;
        RECT 71.800 147.885 72.130 148.645 ;
        RECT 65.340 147.400 65.510 147.545 ;
        RECT 65.225 147.070 65.510 147.400 ;
        RECT 65.340 146.815 65.510 147.070 ;
        RECT 65.745 146.995 66.075 147.365 ;
        RECT 66.265 147.015 66.785 147.555 ;
        RECT 66.955 146.845 67.475 147.385 ;
        RECT 67.645 147.035 69.335 147.555 ;
        RECT 71.415 147.545 72.130 147.715 ;
        RECT 72.300 147.570 72.555 148.475 ;
        RECT 69.505 146.865 71.155 147.385 ;
        RECT 71.325 146.995 71.680 147.365 ;
        RECT 71.960 147.335 72.130 147.545 ;
        RECT 71.960 147.005 72.215 147.335 ;
        RECT 64.885 146.265 65.145 146.770 ;
        RECT 65.340 146.645 66.005 146.815 ;
        RECT 65.325 146.095 65.655 146.475 ;
        RECT 65.835 146.265 66.005 146.645 ;
        RECT 66.265 146.095 67.475 146.845 ;
        RECT 67.645 146.095 71.155 146.865 ;
        RECT 71.960 146.815 72.130 147.005 ;
        RECT 72.385 146.840 72.555 147.570 ;
        RECT 72.730 147.495 72.990 148.645 ;
        RECT 73.715 147.715 73.885 148.475 ;
        RECT 74.100 147.885 74.430 148.645 ;
        RECT 73.715 147.545 74.430 147.715 ;
        RECT 74.600 147.570 74.855 148.475 ;
        RECT 73.625 146.995 73.980 147.365 ;
        RECT 74.260 147.335 74.430 147.545 ;
        RECT 74.260 147.005 74.515 147.335 ;
        RECT 71.415 146.645 72.130 146.815 ;
        RECT 71.415 146.265 71.585 146.645 ;
        RECT 71.800 146.095 72.130 146.475 ;
        RECT 72.300 146.265 72.555 146.840 ;
        RECT 72.730 146.095 72.990 146.935 ;
        RECT 74.260 146.815 74.430 147.005 ;
        RECT 74.685 146.840 74.855 147.570 ;
        RECT 75.030 147.495 75.290 148.645 ;
        RECT 75.925 147.480 76.215 148.645 ;
        RECT 76.475 147.715 76.645 148.475 ;
        RECT 76.860 147.885 77.190 148.645 ;
        RECT 76.475 147.545 77.190 147.715 ;
        RECT 77.360 147.570 77.615 148.475 ;
        RECT 76.385 146.995 76.740 147.365 ;
        RECT 77.020 147.335 77.190 147.545 ;
        RECT 77.020 147.005 77.275 147.335 ;
        RECT 73.715 146.645 74.430 146.815 ;
        RECT 73.715 146.265 73.885 146.645 ;
        RECT 74.100 146.095 74.430 146.475 ;
        RECT 74.600 146.265 74.855 146.840 ;
        RECT 75.030 146.095 75.290 146.935 ;
        RECT 75.925 146.095 76.215 146.820 ;
        RECT 77.020 146.815 77.190 147.005 ;
        RECT 77.445 146.840 77.615 147.570 ;
        RECT 77.790 147.495 78.050 148.645 ;
        RECT 78.890 147.675 79.220 148.475 ;
        RECT 79.390 147.845 79.720 148.645 ;
        RECT 80.020 147.675 80.350 148.475 ;
        RECT 80.995 147.845 81.245 148.645 ;
        RECT 78.890 147.505 81.325 147.675 ;
        RECT 81.515 147.505 81.685 148.645 ;
        RECT 81.855 147.505 82.195 148.475 ;
        RECT 78.685 147.085 79.035 147.335 ;
        RECT 76.475 146.645 77.190 146.815 ;
        RECT 76.475 146.265 76.645 146.645 ;
        RECT 76.860 146.095 77.190 146.475 ;
        RECT 77.360 146.265 77.615 146.840 ;
        RECT 77.790 146.095 78.050 146.935 ;
        RECT 79.220 146.875 79.390 147.505 ;
        RECT 79.560 147.085 79.890 147.285 ;
        RECT 80.060 147.085 80.390 147.285 ;
        RECT 80.560 147.085 80.980 147.285 ;
        RECT 81.155 147.255 81.325 147.505 ;
        RECT 81.155 147.085 81.850 147.255 ;
        RECT 78.890 146.265 79.390 146.875 ;
        RECT 80.020 146.745 81.245 146.915 ;
        RECT 82.020 146.895 82.195 147.505 ;
        RECT 80.020 146.265 80.350 146.745 ;
        RECT 80.520 146.095 80.745 146.555 ;
        RECT 80.915 146.265 81.245 146.745 ;
        RECT 81.435 146.095 81.685 146.895 ;
        RECT 81.855 146.265 82.195 146.895 ;
        RECT 82.365 147.505 82.705 148.475 ;
        RECT 82.875 147.505 83.045 148.645 ;
        RECT 83.315 147.845 83.565 148.645 ;
        RECT 84.210 147.675 84.540 148.475 ;
        RECT 84.840 147.845 85.170 148.645 ;
        RECT 85.340 147.675 85.670 148.475 ;
        RECT 86.970 148.210 92.315 148.645 ;
        RECT 83.235 147.505 85.670 147.675 ;
        RECT 82.365 146.895 82.540 147.505 ;
        RECT 83.235 147.255 83.405 147.505 ;
        RECT 82.710 147.085 83.405 147.255 ;
        RECT 83.580 147.085 84.000 147.285 ;
        RECT 84.170 147.085 84.500 147.285 ;
        RECT 84.670 147.085 85.000 147.285 ;
        RECT 82.365 146.265 82.705 146.895 ;
        RECT 82.875 146.095 83.125 146.895 ;
        RECT 83.315 146.745 84.540 146.915 ;
        RECT 83.315 146.265 83.645 146.745 ;
        RECT 83.815 146.095 84.040 146.555 ;
        RECT 84.210 146.265 84.540 146.745 ;
        RECT 85.170 146.875 85.340 147.505 ;
        RECT 85.525 147.085 85.875 147.335 ;
        RECT 88.560 146.960 88.910 148.210 ;
        RECT 92.545 147.505 92.755 148.645 ;
        RECT 92.925 147.495 93.255 148.475 ;
        RECT 93.425 147.505 93.655 148.645 ;
        RECT 93.865 147.555 95.075 148.645 ;
        RECT 85.170 146.265 85.670 146.875 ;
        RECT 90.390 146.640 90.730 147.470 ;
        RECT 86.970 146.095 92.315 146.640 ;
        RECT 92.545 146.095 92.755 146.915 ;
        RECT 92.925 146.895 93.175 147.495 ;
        RECT 93.345 147.085 93.675 147.335 ;
        RECT 93.865 147.015 94.385 147.555 ;
        RECT 95.245 147.505 95.515 148.475 ;
        RECT 95.725 147.845 96.005 148.645 ;
        RECT 96.175 148.135 97.830 148.425 ;
        RECT 96.240 147.795 97.830 147.965 ;
        RECT 96.240 147.675 96.410 147.795 ;
        RECT 95.685 147.505 96.410 147.675 ;
        RECT 92.925 146.265 93.255 146.895 ;
        RECT 93.425 146.095 93.655 146.915 ;
        RECT 94.555 146.845 95.075 147.385 ;
        RECT 93.865 146.095 95.075 146.845 ;
        RECT 95.245 146.770 95.415 147.505 ;
        RECT 95.685 147.335 95.855 147.505 ;
        RECT 96.600 147.455 97.315 147.625 ;
        RECT 97.510 147.505 97.830 147.795 ;
        RECT 98.005 147.505 98.345 148.475 ;
        RECT 98.515 147.505 98.685 148.645 ;
        RECT 98.955 147.845 99.205 148.645 ;
        RECT 99.850 147.675 100.180 148.475 ;
        RECT 100.480 147.845 100.810 148.645 ;
        RECT 100.980 147.675 101.310 148.475 ;
        RECT 98.875 147.505 101.310 147.675 ;
        RECT 95.585 147.005 95.855 147.335 ;
        RECT 96.025 147.005 96.430 147.335 ;
        RECT 96.600 147.005 97.310 147.455 ;
        RECT 95.685 146.835 95.855 147.005 ;
        RECT 95.245 146.425 95.515 146.770 ;
        RECT 95.685 146.665 97.295 146.835 ;
        RECT 97.480 146.765 97.830 147.335 ;
        RECT 98.005 146.945 98.180 147.505 ;
        RECT 98.875 147.255 99.045 147.505 ;
        RECT 98.350 147.085 99.045 147.255 ;
        RECT 99.220 147.085 99.640 147.285 ;
        RECT 99.810 147.085 100.140 147.285 ;
        RECT 100.310 147.085 100.640 147.285 ;
        RECT 98.005 146.895 98.235 146.945 ;
        RECT 95.705 146.095 96.085 146.495 ;
        RECT 96.255 146.315 96.425 146.665 ;
        RECT 96.595 146.095 96.925 146.495 ;
        RECT 97.125 146.315 97.295 146.665 ;
        RECT 97.495 146.095 97.825 146.595 ;
        RECT 98.005 146.265 98.345 146.895 ;
        RECT 98.515 146.095 98.765 146.895 ;
        RECT 98.955 146.745 100.180 146.915 ;
        RECT 98.955 146.265 99.285 146.745 ;
        RECT 99.455 146.095 99.680 146.555 ;
        RECT 99.850 146.265 100.180 146.745 ;
        RECT 100.810 146.875 100.980 147.505 ;
        RECT 101.685 147.480 101.975 148.645 ;
        RECT 102.150 148.210 107.495 148.645 ;
        RECT 101.165 147.085 101.515 147.335 ;
        RECT 103.740 146.960 104.090 148.210 ;
        RECT 107.670 148.135 109.325 148.425 ;
        RECT 107.670 147.795 109.260 147.965 ;
        RECT 109.495 147.845 109.775 148.645 ;
        RECT 107.670 147.505 107.990 147.795 ;
        RECT 109.090 147.675 109.260 147.795 ;
        RECT 100.810 146.265 101.310 146.875 ;
        RECT 101.685 146.095 101.975 146.820 ;
        RECT 105.570 146.640 105.910 147.470 ;
        RECT 108.185 147.455 108.900 147.625 ;
        RECT 109.090 147.505 109.815 147.675 ;
        RECT 109.985 147.505 110.255 148.475 ;
        RECT 107.670 146.765 108.020 147.335 ;
        RECT 108.190 147.005 108.900 147.455 ;
        RECT 109.645 147.335 109.815 147.505 ;
        RECT 109.070 147.005 109.475 147.335 ;
        RECT 109.645 147.005 109.915 147.335 ;
        RECT 109.645 146.835 109.815 147.005 ;
        RECT 108.205 146.665 109.815 146.835 ;
        RECT 110.085 146.770 110.255 147.505 ;
        RECT 102.150 146.095 107.495 146.640 ;
        RECT 107.675 146.095 108.005 146.595 ;
        RECT 108.205 146.315 108.375 146.665 ;
        RECT 108.575 146.095 108.905 146.495 ;
        RECT 109.075 146.315 109.245 146.665 ;
        RECT 109.415 146.095 109.795 146.495 ;
        RECT 109.985 146.425 110.255 146.770 ;
        RECT 110.425 147.505 110.765 148.475 ;
        RECT 110.935 147.505 111.105 148.645 ;
        RECT 111.375 147.845 111.625 148.645 ;
        RECT 112.270 147.675 112.600 148.475 ;
        RECT 112.900 147.845 113.230 148.645 ;
        RECT 113.400 147.675 113.730 148.475 ;
        RECT 111.295 147.505 113.730 147.675 ;
        RECT 114.565 147.555 116.235 148.645 ;
        RECT 116.405 147.885 116.920 148.295 ;
        RECT 117.155 147.885 117.325 148.645 ;
        RECT 117.495 148.305 119.525 148.475 ;
        RECT 110.425 146.945 110.600 147.505 ;
        RECT 111.295 147.255 111.465 147.505 ;
        RECT 110.770 147.085 111.465 147.255 ;
        RECT 111.640 147.085 112.060 147.285 ;
        RECT 112.230 147.085 112.560 147.285 ;
        RECT 112.730 147.085 113.060 147.285 ;
        RECT 110.425 146.895 110.655 146.945 ;
        RECT 110.425 146.265 110.765 146.895 ;
        RECT 110.935 146.095 111.185 146.895 ;
        RECT 111.375 146.745 112.600 146.915 ;
        RECT 111.375 146.265 111.705 146.745 ;
        RECT 111.875 146.095 112.100 146.555 ;
        RECT 112.270 146.265 112.600 146.745 ;
        RECT 113.230 146.875 113.400 147.505 ;
        RECT 113.585 147.085 113.935 147.335 ;
        RECT 114.565 147.035 115.315 147.555 ;
        RECT 113.230 146.265 113.730 146.875 ;
        RECT 115.485 146.865 116.235 147.385 ;
        RECT 116.405 147.075 116.745 147.885 ;
        RECT 117.495 147.640 117.665 148.305 ;
        RECT 118.060 147.965 119.185 148.135 ;
        RECT 116.915 147.450 117.665 147.640 ;
        RECT 117.835 147.625 118.845 147.795 ;
        RECT 116.405 146.905 117.635 147.075 ;
        RECT 114.565 146.095 116.235 146.865 ;
        RECT 116.680 146.300 116.925 146.905 ;
        RECT 117.145 146.095 117.655 146.630 ;
        RECT 117.835 146.265 118.025 147.625 ;
        RECT 118.195 147.285 118.470 147.425 ;
        RECT 118.195 147.115 118.475 147.285 ;
        RECT 118.195 146.265 118.470 147.115 ;
        RECT 118.675 146.825 118.845 147.625 ;
        RECT 119.015 146.835 119.185 147.965 ;
        RECT 119.355 147.335 119.525 148.305 ;
        RECT 119.695 147.505 119.865 148.645 ;
        RECT 120.035 147.505 120.370 148.475 ;
        RECT 119.355 147.005 119.550 147.335 ;
        RECT 119.775 147.005 120.030 147.335 ;
        RECT 119.775 146.835 119.945 147.005 ;
        RECT 120.200 146.835 120.370 147.505 ;
        RECT 120.545 147.555 121.755 148.645 ;
        RECT 122.015 147.715 122.185 148.475 ;
        RECT 122.365 147.885 122.695 148.645 ;
        RECT 120.545 147.015 121.065 147.555 ;
        RECT 122.015 147.545 122.680 147.715 ;
        RECT 122.865 147.570 123.135 148.475 ;
        RECT 122.510 147.400 122.680 147.545 ;
        RECT 121.235 146.845 121.755 147.385 ;
        RECT 121.945 146.995 122.275 147.365 ;
        RECT 122.510 147.070 122.795 147.400 ;
        RECT 119.015 146.665 119.945 146.835 ;
        RECT 119.015 146.630 119.190 146.665 ;
        RECT 118.660 146.265 119.190 146.630 ;
        RECT 119.615 146.095 119.945 146.495 ;
        RECT 120.115 146.265 120.370 146.835 ;
        RECT 120.545 146.095 121.755 146.845 ;
        RECT 122.510 146.815 122.680 147.070 ;
        RECT 122.015 146.645 122.680 146.815 ;
        RECT 122.965 146.770 123.135 147.570 ;
        RECT 123.765 147.555 126.355 148.645 ;
        RECT 126.525 147.555 127.735 148.645 ;
        RECT 123.765 147.035 124.975 147.555 ;
        RECT 125.145 146.865 126.355 147.385 ;
        RECT 126.525 147.015 127.045 147.555 ;
        RECT 122.015 146.265 122.185 146.645 ;
        RECT 122.365 146.095 122.695 146.475 ;
        RECT 122.875 146.265 123.135 146.770 ;
        RECT 123.765 146.095 126.355 146.865 ;
        RECT 127.215 146.845 127.735 147.385 ;
        RECT 126.525 146.095 127.735 146.845 ;
        RECT 14.660 145.925 127.820 146.095 ;
        RECT 14.745 145.175 15.955 145.925 ;
        RECT 17.135 145.375 17.305 145.755 ;
        RECT 17.485 145.545 17.815 145.925 ;
        RECT 17.135 145.205 17.800 145.375 ;
        RECT 17.995 145.250 18.255 145.755 ;
        RECT 14.745 144.635 15.265 145.175 ;
        RECT 15.435 144.465 15.955 145.005 ;
        RECT 17.065 144.655 17.395 145.025 ;
        RECT 17.630 144.950 17.800 145.205 ;
        RECT 17.630 144.620 17.915 144.950 ;
        RECT 17.630 144.475 17.800 144.620 ;
        RECT 14.745 143.375 15.955 144.465 ;
        RECT 17.135 144.305 17.800 144.475 ;
        RECT 18.085 144.450 18.255 145.250 ;
        RECT 17.135 143.545 17.305 144.305 ;
        RECT 17.485 143.375 17.815 144.135 ;
        RECT 17.985 143.545 18.255 144.450 ;
        RECT 18.430 145.215 18.685 145.745 ;
        RECT 18.855 145.465 19.160 145.925 ;
        RECT 19.405 145.545 20.475 145.715 ;
        RECT 18.430 144.565 18.640 145.215 ;
        RECT 19.405 145.190 19.725 145.545 ;
        RECT 19.400 145.015 19.725 145.190 ;
        RECT 18.810 144.715 19.725 145.015 ;
        RECT 19.895 144.975 20.135 145.375 ;
        RECT 20.305 145.315 20.475 145.545 ;
        RECT 20.645 145.485 20.835 145.925 ;
        RECT 21.005 145.475 21.955 145.755 ;
        RECT 22.175 145.565 22.525 145.735 ;
        RECT 20.305 145.145 20.835 145.315 ;
        RECT 18.810 144.685 19.550 144.715 ;
        RECT 18.430 143.685 18.685 144.565 ;
        RECT 18.855 143.375 19.160 144.515 ;
        RECT 19.380 144.095 19.550 144.685 ;
        RECT 19.895 144.605 20.435 144.975 ;
        RECT 20.615 144.865 20.835 145.145 ;
        RECT 21.005 144.695 21.175 145.475 ;
        RECT 20.770 144.525 21.175 144.695 ;
        RECT 21.345 144.685 21.695 145.305 ;
        RECT 20.770 144.435 20.940 144.525 ;
        RECT 21.865 144.515 22.075 145.305 ;
        RECT 19.720 144.265 20.940 144.435 ;
        RECT 21.400 144.355 22.075 144.515 ;
        RECT 19.380 143.925 20.180 144.095 ;
        RECT 19.500 143.375 19.830 143.755 ;
        RECT 20.010 143.635 20.180 143.925 ;
        RECT 20.770 143.885 20.940 144.265 ;
        RECT 21.110 144.345 22.075 144.355 ;
        RECT 22.265 145.175 22.525 145.565 ;
        RECT 22.735 145.465 23.065 145.925 ;
        RECT 23.940 145.535 24.795 145.705 ;
        RECT 25.000 145.535 25.495 145.705 ;
        RECT 25.665 145.565 25.995 145.925 ;
        RECT 22.265 144.485 22.435 145.175 ;
        RECT 22.605 144.825 22.775 145.005 ;
        RECT 22.945 144.995 23.735 145.245 ;
        RECT 23.940 144.825 24.110 145.535 ;
        RECT 24.280 145.025 24.635 145.245 ;
        RECT 22.605 144.655 24.295 144.825 ;
        RECT 21.110 144.055 21.570 144.345 ;
        RECT 22.265 144.315 23.765 144.485 ;
        RECT 22.265 144.175 22.435 144.315 ;
        RECT 21.875 144.005 22.435 144.175 ;
        RECT 20.350 143.375 20.600 143.835 ;
        RECT 20.770 143.545 21.640 143.885 ;
        RECT 21.875 143.545 22.045 144.005 ;
        RECT 22.880 143.975 23.955 144.145 ;
        RECT 22.215 143.375 22.585 143.835 ;
        RECT 22.880 143.635 23.050 143.975 ;
        RECT 23.220 143.375 23.550 143.805 ;
        RECT 23.785 143.635 23.955 143.975 ;
        RECT 24.125 143.875 24.295 144.655 ;
        RECT 24.465 144.435 24.635 145.025 ;
        RECT 24.805 144.625 25.155 145.245 ;
        RECT 24.465 144.045 24.930 144.435 ;
        RECT 25.325 144.175 25.495 145.535 ;
        RECT 25.665 144.345 26.125 145.395 ;
        RECT 25.100 144.005 25.495 144.175 ;
        RECT 25.100 143.875 25.270 144.005 ;
        RECT 24.125 143.545 24.805 143.875 ;
        RECT 25.020 143.545 25.270 143.875 ;
        RECT 25.440 143.375 25.690 143.835 ;
        RECT 25.860 143.560 26.185 144.345 ;
        RECT 26.355 143.545 26.525 145.665 ;
        RECT 26.695 145.545 27.025 145.925 ;
        RECT 27.195 145.375 27.450 145.665 ;
        RECT 26.700 145.205 27.450 145.375 ;
        RECT 27.630 145.215 27.885 145.745 ;
        RECT 28.055 145.465 28.360 145.925 ;
        RECT 28.605 145.545 29.675 145.715 ;
        RECT 26.700 144.215 26.930 145.205 ;
        RECT 27.100 144.385 27.450 145.035 ;
        RECT 27.630 144.565 27.840 145.215 ;
        RECT 28.605 145.190 28.925 145.545 ;
        RECT 28.600 145.015 28.925 145.190 ;
        RECT 28.010 144.715 28.925 145.015 ;
        RECT 29.095 144.975 29.335 145.375 ;
        RECT 29.505 145.315 29.675 145.545 ;
        RECT 29.845 145.485 30.035 145.925 ;
        RECT 30.205 145.475 31.155 145.755 ;
        RECT 31.375 145.565 31.725 145.735 ;
        RECT 29.505 145.145 30.035 145.315 ;
        RECT 28.010 144.685 28.750 144.715 ;
        RECT 26.700 144.045 27.450 144.215 ;
        RECT 26.695 143.375 27.025 143.875 ;
        RECT 27.195 143.545 27.450 144.045 ;
        RECT 27.630 143.685 27.885 144.565 ;
        RECT 28.055 143.375 28.360 144.515 ;
        RECT 28.580 144.095 28.750 144.685 ;
        RECT 29.095 144.605 29.635 144.975 ;
        RECT 29.815 144.865 30.035 145.145 ;
        RECT 30.205 144.695 30.375 145.475 ;
        RECT 29.970 144.525 30.375 144.695 ;
        RECT 30.545 144.685 30.895 145.305 ;
        RECT 29.970 144.435 30.140 144.525 ;
        RECT 31.065 144.515 31.275 145.305 ;
        RECT 28.920 144.265 30.140 144.435 ;
        RECT 30.600 144.355 31.275 144.515 ;
        RECT 28.580 143.925 29.380 144.095 ;
        RECT 28.700 143.375 29.030 143.755 ;
        RECT 29.210 143.635 29.380 143.925 ;
        RECT 29.970 143.885 30.140 144.265 ;
        RECT 30.310 144.345 31.275 144.355 ;
        RECT 31.465 145.175 31.725 145.565 ;
        RECT 31.935 145.465 32.265 145.925 ;
        RECT 33.140 145.535 33.995 145.705 ;
        RECT 34.200 145.535 34.695 145.705 ;
        RECT 34.865 145.565 35.195 145.925 ;
        RECT 31.465 144.485 31.635 145.175 ;
        RECT 31.805 144.825 31.975 145.005 ;
        RECT 32.145 144.995 32.935 145.245 ;
        RECT 33.140 144.825 33.310 145.535 ;
        RECT 33.480 145.025 33.835 145.245 ;
        RECT 31.805 144.655 33.495 144.825 ;
        RECT 30.310 144.055 30.770 144.345 ;
        RECT 31.465 144.315 32.965 144.485 ;
        RECT 31.465 144.175 31.635 144.315 ;
        RECT 31.075 144.005 31.635 144.175 ;
        RECT 29.550 143.375 29.800 143.835 ;
        RECT 29.970 143.545 30.840 143.885 ;
        RECT 31.075 143.545 31.245 144.005 ;
        RECT 32.080 143.975 33.155 144.145 ;
        RECT 31.415 143.375 31.785 143.835 ;
        RECT 32.080 143.635 32.250 143.975 ;
        RECT 32.420 143.375 32.750 143.805 ;
        RECT 32.985 143.635 33.155 143.975 ;
        RECT 33.325 143.875 33.495 144.655 ;
        RECT 33.665 144.435 33.835 145.025 ;
        RECT 34.005 144.625 34.355 145.245 ;
        RECT 33.665 144.045 34.130 144.435 ;
        RECT 34.525 144.175 34.695 145.535 ;
        RECT 34.865 144.345 35.325 145.395 ;
        RECT 34.300 144.005 34.695 144.175 ;
        RECT 34.300 143.875 34.470 144.005 ;
        RECT 33.325 143.545 34.005 143.875 ;
        RECT 34.220 143.545 34.470 143.875 ;
        RECT 34.640 143.375 34.890 143.835 ;
        RECT 35.060 143.560 35.385 144.345 ;
        RECT 35.555 143.545 35.725 145.665 ;
        RECT 35.895 145.545 36.225 145.925 ;
        RECT 36.395 145.375 36.650 145.665 ;
        RECT 35.900 145.205 36.650 145.375 ;
        RECT 35.900 144.215 36.130 145.205 ;
        RECT 37.285 145.200 37.575 145.925 ;
        RECT 38.020 145.115 38.265 145.720 ;
        RECT 38.485 145.390 38.995 145.925 ;
        RECT 36.300 144.385 36.650 145.035 ;
        RECT 37.745 144.945 38.975 145.115 ;
        RECT 35.900 144.045 36.650 144.215 ;
        RECT 35.895 143.375 36.225 143.875 ;
        RECT 36.395 143.545 36.650 144.045 ;
        RECT 37.285 143.375 37.575 144.540 ;
        RECT 37.745 144.135 38.085 144.945 ;
        RECT 38.255 144.380 39.005 144.570 ;
        RECT 37.745 143.725 38.260 144.135 ;
        RECT 38.495 143.375 38.665 144.135 ;
        RECT 38.835 143.715 39.005 144.380 ;
        RECT 39.175 144.395 39.365 145.755 ;
        RECT 39.535 145.245 39.810 145.755 ;
        RECT 40.000 145.390 40.530 145.755 ;
        RECT 40.955 145.525 41.285 145.925 ;
        RECT 40.355 145.355 40.530 145.390 ;
        RECT 39.535 145.075 39.815 145.245 ;
        RECT 39.535 144.595 39.810 145.075 ;
        RECT 40.015 144.395 40.185 145.195 ;
        RECT 39.175 144.225 40.185 144.395 ;
        RECT 40.355 145.185 41.285 145.355 ;
        RECT 41.455 145.185 41.710 145.755 ;
        RECT 40.355 144.055 40.525 145.185 ;
        RECT 41.115 145.015 41.285 145.185 ;
        RECT 39.400 143.885 40.525 144.055 ;
        RECT 40.695 144.685 40.890 145.015 ;
        RECT 41.115 144.685 41.370 145.015 ;
        RECT 40.695 143.715 40.865 144.685 ;
        RECT 41.540 144.515 41.710 145.185 ;
        RECT 42.550 145.145 43.050 145.755 ;
        RECT 42.345 144.685 42.695 144.935 ;
        RECT 42.880 144.515 43.050 145.145 ;
        RECT 43.680 145.275 44.010 145.755 ;
        RECT 44.180 145.465 44.405 145.925 ;
        RECT 44.575 145.275 44.905 145.755 ;
        RECT 43.680 145.105 44.905 145.275 ;
        RECT 45.095 145.125 45.345 145.925 ;
        RECT 45.515 145.125 45.855 145.755 ;
        RECT 43.220 144.735 43.550 144.935 ;
        RECT 43.720 144.735 44.050 144.935 ;
        RECT 44.220 144.735 44.640 144.935 ;
        RECT 44.815 144.765 45.510 144.935 ;
        RECT 44.815 144.515 44.985 144.765 ;
        RECT 45.680 144.515 45.855 145.125 ;
        RECT 38.835 143.545 40.865 143.715 ;
        RECT 41.035 143.375 41.205 144.515 ;
        RECT 41.375 143.545 41.710 144.515 ;
        RECT 42.550 144.345 44.985 144.515 ;
        RECT 42.550 143.545 42.880 144.345 ;
        RECT 43.050 143.375 43.380 144.175 ;
        RECT 43.680 143.545 44.010 144.345 ;
        RECT 44.655 143.375 44.905 144.175 ;
        RECT 45.175 143.375 45.345 144.515 ;
        RECT 45.515 143.545 45.855 144.515 ;
        RECT 46.025 145.125 46.365 145.755 ;
        RECT 46.535 145.125 46.785 145.925 ;
        RECT 46.975 145.275 47.305 145.755 ;
        RECT 47.475 145.465 47.700 145.925 ;
        RECT 47.870 145.275 48.200 145.755 ;
        RECT 46.025 145.075 46.255 145.125 ;
        RECT 46.975 145.105 48.200 145.275 ;
        RECT 48.830 145.145 49.330 145.755 ;
        RECT 50.165 145.155 53.675 145.925 ;
        RECT 46.025 144.515 46.200 145.075 ;
        RECT 46.370 144.765 47.065 144.935 ;
        RECT 46.895 144.515 47.065 144.765 ;
        RECT 47.240 144.735 47.660 144.935 ;
        RECT 47.830 144.735 48.160 144.935 ;
        RECT 48.330 144.735 48.660 144.935 ;
        RECT 48.830 144.515 49.000 145.145 ;
        RECT 49.185 144.685 49.535 144.935 ;
        RECT 46.025 143.545 46.365 144.515 ;
        RECT 46.535 143.375 46.705 144.515 ;
        RECT 46.895 144.345 49.330 144.515 ;
        RECT 46.975 143.375 47.225 144.175 ;
        RECT 47.870 143.545 48.200 144.345 ;
        RECT 48.500 143.375 48.830 144.175 ;
        RECT 49.000 143.545 49.330 144.345 ;
        RECT 50.165 144.465 51.855 144.985 ;
        RECT 52.025 144.635 53.675 145.155 ;
        RECT 53.850 145.215 54.105 145.745 ;
        RECT 54.275 145.465 54.580 145.925 ;
        RECT 54.825 145.545 55.895 145.715 ;
        RECT 53.850 144.565 54.060 145.215 ;
        RECT 54.825 145.190 55.145 145.545 ;
        RECT 54.820 145.015 55.145 145.190 ;
        RECT 54.230 144.715 55.145 145.015 ;
        RECT 55.315 144.975 55.555 145.375 ;
        RECT 55.725 145.315 55.895 145.545 ;
        RECT 56.065 145.485 56.255 145.925 ;
        RECT 56.425 145.475 57.375 145.755 ;
        RECT 57.595 145.565 57.945 145.735 ;
        RECT 55.725 145.145 56.255 145.315 ;
        RECT 54.230 144.685 54.970 144.715 ;
        RECT 50.165 143.375 53.675 144.465 ;
        RECT 53.850 143.685 54.105 144.565 ;
        RECT 54.275 143.375 54.580 144.515 ;
        RECT 54.800 144.095 54.970 144.685 ;
        RECT 55.315 144.605 55.855 144.975 ;
        RECT 56.035 144.865 56.255 145.145 ;
        RECT 56.425 144.695 56.595 145.475 ;
        RECT 56.190 144.525 56.595 144.695 ;
        RECT 56.765 144.685 57.115 145.305 ;
        RECT 56.190 144.435 56.360 144.525 ;
        RECT 57.285 144.515 57.495 145.305 ;
        RECT 55.140 144.265 56.360 144.435 ;
        RECT 56.820 144.355 57.495 144.515 ;
        RECT 54.800 143.925 55.600 144.095 ;
        RECT 54.920 143.375 55.250 143.755 ;
        RECT 55.430 143.635 55.600 143.925 ;
        RECT 56.190 143.885 56.360 144.265 ;
        RECT 56.530 144.345 57.495 144.355 ;
        RECT 57.685 145.175 57.945 145.565 ;
        RECT 58.155 145.465 58.485 145.925 ;
        RECT 59.360 145.535 60.215 145.705 ;
        RECT 60.420 145.535 60.915 145.705 ;
        RECT 61.085 145.565 61.415 145.925 ;
        RECT 57.685 144.485 57.855 145.175 ;
        RECT 58.025 144.825 58.195 145.005 ;
        RECT 58.365 144.995 59.155 145.245 ;
        RECT 59.360 144.825 59.530 145.535 ;
        RECT 59.700 145.025 60.055 145.245 ;
        RECT 58.025 144.655 59.715 144.825 ;
        RECT 56.530 144.055 56.990 144.345 ;
        RECT 57.685 144.315 59.185 144.485 ;
        RECT 57.685 144.175 57.855 144.315 ;
        RECT 57.295 144.005 57.855 144.175 ;
        RECT 55.770 143.375 56.020 143.835 ;
        RECT 56.190 143.545 57.060 143.885 ;
        RECT 57.295 143.545 57.465 144.005 ;
        RECT 58.300 143.975 59.375 144.145 ;
        RECT 57.635 143.375 58.005 143.835 ;
        RECT 58.300 143.635 58.470 143.975 ;
        RECT 58.640 143.375 58.970 143.805 ;
        RECT 59.205 143.635 59.375 143.975 ;
        RECT 59.545 143.875 59.715 144.655 ;
        RECT 59.885 144.435 60.055 145.025 ;
        RECT 60.225 144.625 60.575 145.245 ;
        RECT 59.885 144.045 60.350 144.435 ;
        RECT 60.745 144.175 60.915 145.535 ;
        RECT 61.085 144.345 61.545 145.395 ;
        RECT 60.520 144.005 60.915 144.175 ;
        RECT 60.520 143.875 60.690 144.005 ;
        RECT 59.545 143.545 60.225 143.875 ;
        RECT 60.440 143.545 60.690 143.875 ;
        RECT 60.860 143.375 61.110 143.835 ;
        RECT 61.280 143.560 61.605 144.345 ;
        RECT 61.775 143.545 61.945 145.665 ;
        RECT 62.115 145.545 62.445 145.925 ;
        RECT 62.615 145.375 62.870 145.665 ;
        RECT 62.120 145.205 62.870 145.375 ;
        RECT 62.120 144.215 62.350 145.205 ;
        RECT 63.045 145.200 63.335 145.925 ;
        RECT 63.510 145.185 63.765 145.755 ;
        RECT 63.935 145.525 64.265 145.925 ;
        RECT 64.690 145.390 65.220 145.755 ;
        RECT 65.410 145.585 65.685 145.755 ;
        RECT 65.405 145.415 65.685 145.585 ;
        RECT 64.690 145.355 64.865 145.390 ;
        RECT 63.935 145.185 64.865 145.355 ;
        RECT 62.520 144.385 62.870 145.035 ;
        RECT 62.120 144.045 62.870 144.215 ;
        RECT 62.115 143.375 62.445 143.875 ;
        RECT 62.615 143.545 62.870 144.045 ;
        RECT 63.045 143.375 63.335 144.540 ;
        RECT 63.510 144.515 63.680 145.185 ;
        RECT 63.935 145.015 64.105 145.185 ;
        RECT 63.850 144.685 64.105 145.015 ;
        RECT 64.330 144.685 64.525 145.015 ;
        RECT 63.510 143.545 63.845 144.515 ;
        RECT 64.015 143.375 64.185 144.515 ;
        RECT 64.355 143.715 64.525 144.685 ;
        RECT 64.695 144.055 64.865 145.185 ;
        RECT 65.035 144.395 65.205 145.195 ;
        RECT 65.410 144.595 65.685 145.415 ;
        RECT 65.855 144.395 66.045 145.755 ;
        RECT 66.225 145.390 66.735 145.925 ;
        RECT 66.955 145.115 67.200 145.720 ;
        RECT 66.245 144.945 67.475 145.115 ;
        RECT 67.685 145.105 67.915 145.925 ;
        RECT 68.085 145.125 68.415 145.755 ;
        RECT 65.035 144.225 66.045 144.395 ;
        RECT 66.215 144.380 66.965 144.570 ;
        RECT 64.695 143.885 65.820 144.055 ;
        RECT 66.215 143.715 66.385 144.380 ;
        RECT 67.135 144.135 67.475 144.945 ;
        RECT 67.665 144.685 67.995 144.935 ;
        RECT 68.165 144.525 68.415 145.125 ;
        RECT 68.585 145.105 68.795 145.925 ;
        RECT 69.575 145.375 69.745 145.755 ;
        RECT 69.925 145.545 70.255 145.925 ;
        RECT 69.575 145.205 70.240 145.375 ;
        RECT 70.435 145.250 70.695 145.755 ;
        RECT 69.505 144.655 69.835 145.025 ;
        RECT 70.070 144.950 70.240 145.205 ;
        RECT 64.355 143.545 66.385 143.715 ;
        RECT 66.555 143.375 66.725 144.135 ;
        RECT 66.960 143.725 67.475 144.135 ;
        RECT 67.685 143.375 67.915 144.515 ;
        RECT 68.085 143.545 68.415 144.525 ;
        RECT 70.070 144.620 70.355 144.950 ;
        RECT 68.585 143.375 68.795 144.515 ;
        RECT 70.070 144.475 70.240 144.620 ;
        RECT 69.575 144.305 70.240 144.475 ;
        RECT 70.525 144.450 70.695 145.250 ;
        RECT 70.865 145.155 74.375 145.925 ;
        RECT 74.550 145.380 79.895 145.925 ;
        RECT 69.575 143.545 69.745 144.305 ;
        RECT 69.925 143.375 70.255 144.135 ;
        RECT 70.425 143.545 70.695 144.450 ;
        RECT 70.865 144.465 72.555 144.985 ;
        RECT 72.725 144.635 74.375 145.155 ;
        RECT 70.865 143.375 74.375 144.465 ;
        RECT 76.140 143.810 76.490 145.060 ;
        RECT 77.970 144.550 78.310 145.380 ;
        RECT 80.065 145.125 80.405 145.755 ;
        RECT 80.575 145.125 80.825 145.925 ;
        RECT 81.015 145.275 81.345 145.755 ;
        RECT 81.515 145.465 81.740 145.925 ;
        RECT 81.910 145.275 82.240 145.755 ;
        RECT 80.065 144.515 80.240 145.125 ;
        RECT 81.015 145.105 82.240 145.275 ;
        RECT 82.870 145.145 83.370 145.755 ;
        RECT 80.410 144.765 81.105 144.935 ;
        RECT 80.935 144.515 81.105 144.765 ;
        RECT 81.280 144.735 81.700 144.935 ;
        RECT 81.870 144.735 82.200 144.935 ;
        RECT 82.370 144.735 82.700 144.935 ;
        RECT 82.870 144.515 83.040 145.145 ;
        RECT 84.940 145.115 85.185 145.720 ;
        RECT 85.405 145.390 85.915 145.925 ;
        RECT 84.665 144.945 85.895 145.115 ;
        RECT 83.225 144.685 83.575 144.935 ;
        RECT 74.550 143.375 79.895 143.810 ;
        RECT 80.065 143.545 80.405 144.515 ;
        RECT 80.575 143.375 80.745 144.515 ;
        RECT 80.935 144.345 83.370 144.515 ;
        RECT 81.015 143.375 81.265 144.175 ;
        RECT 81.910 143.545 82.240 144.345 ;
        RECT 82.540 143.375 82.870 144.175 ;
        RECT 83.040 143.545 83.370 144.345 ;
        RECT 84.665 144.135 85.005 144.945 ;
        RECT 85.175 144.380 85.925 144.570 ;
        RECT 84.665 143.725 85.180 144.135 ;
        RECT 85.415 143.375 85.585 144.135 ;
        RECT 85.755 143.715 85.925 144.380 ;
        RECT 86.095 144.395 86.285 145.755 ;
        RECT 86.455 144.905 86.730 145.755 ;
        RECT 86.920 145.390 87.450 145.755 ;
        RECT 87.875 145.525 88.205 145.925 ;
        RECT 87.275 145.355 87.450 145.390 ;
        RECT 86.455 144.735 86.735 144.905 ;
        RECT 86.455 144.595 86.730 144.735 ;
        RECT 86.935 144.395 87.105 145.195 ;
        RECT 86.095 144.225 87.105 144.395 ;
        RECT 87.275 145.185 88.205 145.355 ;
        RECT 88.375 145.185 88.630 145.755 ;
        RECT 88.805 145.200 89.095 145.925 ;
        RECT 89.640 145.215 89.895 145.745 ;
        RECT 90.075 145.465 90.360 145.925 ;
        RECT 87.275 144.055 87.445 145.185 ;
        RECT 88.035 145.015 88.205 145.185 ;
        RECT 86.320 143.885 87.445 144.055 ;
        RECT 87.615 144.685 87.810 145.015 ;
        RECT 88.035 144.685 88.290 145.015 ;
        RECT 87.615 143.715 87.785 144.685 ;
        RECT 88.460 144.515 88.630 145.185 ;
        RECT 89.640 144.565 89.820 145.215 ;
        RECT 90.540 145.015 90.790 145.665 ;
        RECT 89.990 144.685 90.790 145.015 ;
        RECT 85.755 143.545 87.785 143.715 ;
        RECT 87.955 143.375 88.125 144.515 ;
        RECT 88.295 143.545 88.630 144.515 ;
        RECT 88.805 143.375 89.095 144.540 ;
        RECT 89.555 144.395 89.820 144.565 ;
        RECT 89.640 144.355 89.820 144.395 ;
        RECT 89.640 143.685 89.895 144.355 ;
        RECT 90.075 143.375 90.360 144.175 ;
        RECT 90.540 144.095 90.790 144.685 ;
        RECT 90.990 145.330 91.310 145.660 ;
        RECT 91.490 145.445 92.150 145.925 ;
        RECT 92.350 145.535 93.200 145.705 ;
        RECT 90.990 144.435 91.180 145.330 ;
        RECT 91.500 145.005 92.160 145.275 ;
        RECT 91.830 144.945 92.160 145.005 ;
        RECT 91.350 144.775 91.680 144.835 ;
        RECT 92.350 144.775 92.520 145.535 ;
        RECT 93.760 145.465 94.080 145.925 ;
        RECT 94.280 145.285 94.530 145.715 ;
        RECT 94.820 145.485 95.230 145.925 ;
        RECT 95.400 145.545 96.415 145.745 ;
        RECT 92.690 145.115 93.940 145.285 ;
        RECT 92.690 144.995 93.020 145.115 ;
        RECT 91.350 144.605 93.250 144.775 ;
        RECT 90.990 144.265 92.910 144.435 ;
        RECT 90.990 144.245 91.310 144.265 ;
        RECT 90.540 143.585 90.870 144.095 ;
        RECT 91.140 143.635 91.310 144.245 ;
        RECT 93.080 144.095 93.250 144.605 ;
        RECT 93.420 144.535 93.600 144.945 ;
        RECT 93.770 144.355 93.940 145.115 ;
        RECT 91.480 143.375 91.810 144.065 ;
        RECT 92.040 143.925 93.250 144.095 ;
        RECT 93.420 144.045 93.940 144.355 ;
        RECT 94.110 144.945 94.530 145.285 ;
        RECT 94.820 144.945 95.230 145.275 ;
        RECT 94.110 144.175 94.300 144.945 ;
        RECT 95.400 144.815 95.570 145.545 ;
        RECT 96.715 145.375 96.885 145.705 ;
        RECT 97.055 145.545 97.385 145.925 ;
        RECT 95.740 144.995 96.090 145.365 ;
        RECT 95.400 144.775 95.820 144.815 ;
        RECT 94.470 144.605 95.820 144.775 ;
        RECT 94.470 144.445 94.720 144.605 ;
        RECT 95.230 144.175 95.480 144.435 ;
        RECT 94.110 143.925 95.480 144.175 ;
        RECT 92.040 143.635 92.280 143.925 ;
        RECT 93.080 143.845 93.250 143.925 ;
        RECT 92.480 143.375 92.900 143.755 ;
        RECT 93.080 143.595 93.710 143.845 ;
        RECT 94.180 143.375 94.510 143.755 ;
        RECT 94.680 143.635 94.850 143.925 ;
        RECT 95.650 143.760 95.820 144.605 ;
        RECT 96.270 144.435 96.490 145.305 ;
        RECT 96.715 145.185 97.410 145.375 ;
        RECT 95.990 144.055 96.490 144.435 ;
        RECT 96.660 144.385 97.070 145.005 ;
        RECT 97.240 144.215 97.410 145.185 ;
        RECT 96.715 144.045 97.410 144.215 ;
        RECT 95.030 143.375 95.410 143.755 ;
        RECT 95.650 143.590 96.480 143.760 ;
        RECT 96.715 143.545 96.885 144.045 ;
        RECT 97.055 143.375 97.385 143.875 ;
        RECT 97.600 143.545 97.825 145.665 ;
        RECT 97.995 145.545 98.325 145.925 ;
        RECT 98.495 145.375 98.665 145.665 ;
        RECT 99.390 145.380 104.735 145.925 ;
        RECT 104.915 145.425 105.245 145.925 ;
        RECT 98.000 145.205 98.665 145.375 ;
        RECT 98.000 144.215 98.230 145.205 ;
        RECT 98.400 144.385 98.750 145.035 ;
        RECT 98.000 144.045 98.665 144.215 ;
        RECT 97.995 143.375 98.325 143.875 ;
        RECT 98.495 143.545 98.665 144.045 ;
        RECT 100.980 143.810 101.330 145.060 ;
        RECT 102.810 144.550 103.150 145.380 ;
        RECT 105.445 145.355 105.615 145.705 ;
        RECT 105.815 145.525 106.145 145.925 ;
        RECT 106.315 145.355 106.485 145.705 ;
        RECT 106.655 145.525 107.035 145.925 ;
        RECT 104.910 144.685 105.260 145.255 ;
        RECT 105.445 145.185 107.055 145.355 ;
        RECT 107.225 145.250 107.495 145.595 ;
        RECT 106.885 145.015 107.055 145.185 ;
        RECT 105.430 144.565 106.140 145.015 ;
        RECT 106.310 144.685 106.715 145.015 ;
        RECT 106.885 144.685 107.155 145.015 ;
        RECT 104.910 144.225 105.230 144.515 ;
        RECT 105.425 144.395 106.140 144.565 ;
        RECT 106.885 144.515 107.055 144.685 ;
        RECT 107.325 144.515 107.495 145.250 ;
        RECT 106.330 144.345 107.055 144.515 ;
        RECT 106.330 144.225 106.500 144.345 ;
        RECT 104.910 144.055 106.500 144.225 ;
        RECT 99.390 143.375 104.735 143.810 ;
        RECT 104.910 143.595 106.565 143.885 ;
        RECT 106.735 143.375 107.015 144.175 ;
        RECT 107.225 143.545 107.495 144.515 ;
        RECT 107.665 145.125 108.005 145.755 ;
        RECT 108.175 145.125 108.425 145.925 ;
        RECT 108.615 145.275 108.945 145.755 ;
        RECT 109.115 145.465 109.340 145.925 ;
        RECT 109.510 145.275 109.840 145.755 ;
        RECT 107.665 145.075 107.895 145.125 ;
        RECT 108.615 145.105 109.840 145.275 ;
        RECT 110.470 145.145 110.970 145.755 ;
        RECT 111.895 145.275 112.065 145.755 ;
        RECT 112.245 145.445 112.485 145.925 ;
        RECT 112.735 145.275 112.905 145.755 ;
        RECT 113.075 145.445 113.405 145.925 ;
        RECT 113.575 145.275 113.745 145.755 ;
        RECT 107.665 144.515 107.840 145.075 ;
        RECT 108.010 144.765 108.705 144.935 ;
        RECT 108.535 144.515 108.705 144.765 ;
        RECT 108.880 144.735 109.300 144.935 ;
        RECT 109.470 144.735 109.800 144.935 ;
        RECT 109.970 144.735 110.300 144.935 ;
        RECT 110.470 144.515 110.640 145.145 ;
        RECT 111.895 145.105 112.530 145.275 ;
        RECT 112.735 145.105 113.745 145.275 ;
        RECT 113.915 145.125 114.245 145.925 ;
        RECT 114.565 145.200 114.855 145.925 ;
        RECT 115.525 145.105 115.755 145.925 ;
        RECT 115.925 145.125 116.255 145.755 ;
        RECT 112.360 144.935 112.530 145.105 ;
        RECT 110.825 144.685 111.175 144.935 ;
        RECT 111.810 144.695 112.190 144.935 ;
        RECT 112.360 144.765 112.860 144.935 ;
        RECT 113.250 144.905 113.745 145.105 ;
        RECT 112.360 144.525 112.530 144.765 ;
        RECT 113.245 144.735 113.745 144.905 ;
        RECT 113.250 144.565 113.745 144.735 ;
        RECT 115.505 144.685 115.835 144.935 ;
        RECT 107.665 143.545 108.005 144.515 ;
        RECT 108.175 143.375 108.345 144.515 ;
        RECT 108.535 144.345 110.970 144.515 ;
        RECT 108.615 143.375 108.865 144.175 ;
        RECT 109.510 143.545 109.840 144.345 ;
        RECT 110.140 143.375 110.470 144.175 ;
        RECT 110.640 143.545 110.970 144.345 ;
        RECT 111.815 144.355 112.530 144.525 ;
        RECT 112.735 144.395 113.745 144.565 ;
        RECT 111.815 143.545 112.145 144.355 ;
        RECT 112.315 143.375 112.555 144.175 ;
        RECT 112.735 143.545 112.905 144.395 ;
        RECT 113.075 143.375 113.405 144.175 ;
        RECT 113.575 143.545 113.745 144.395 ;
        RECT 113.915 143.375 114.245 144.525 ;
        RECT 114.565 143.375 114.855 144.540 ;
        RECT 116.005 144.525 116.255 145.125 ;
        RECT 116.425 145.105 116.635 145.925 ;
        RECT 117.240 145.215 117.495 145.745 ;
        RECT 117.675 145.465 117.960 145.925 ;
        RECT 117.240 144.905 117.420 145.215 ;
        RECT 118.140 145.015 118.390 145.665 ;
        RECT 117.155 144.735 117.420 144.905 ;
        RECT 115.525 143.375 115.755 144.515 ;
        RECT 115.925 143.545 116.255 144.525 ;
        RECT 116.425 143.375 116.635 144.515 ;
        RECT 117.240 144.355 117.420 144.735 ;
        RECT 117.590 144.685 118.390 145.015 ;
        RECT 117.240 143.685 117.495 144.355 ;
        RECT 117.675 143.375 117.960 144.175 ;
        RECT 118.140 144.095 118.390 144.685 ;
        RECT 118.590 145.330 118.910 145.660 ;
        RECT 119.090 145.445 119.750 145.925 ;
        RECT 119.950 145.535 120.800 145.705 ;
        RECT 118.590 144.435 118.780 145.330 ;
        RECT 119.100 145.005 119.760 145.275 ;
        RECT 119.430 144.945 119.760 145.005 ;
        RECT 118.950 144.775 119.280 144.835 ;
        RECT 119.950 144.775 120.120 145.535 ;
        RECT 121.360 145.465 121.680 145.925 ;
        RECT 121.880 145.285 122.130 145.715 ;
        RECT 122.420 145.485 122.830 145.925 ;
        RECT 123.000 145.545 124.015 145.745 ;
        RECT 120.290 145.115 121.540 145.285 ;
        RECT 120.290 144.995 120.620 145.115 ;
        RECT 118.950 144.605 120.850 144.775 ;
        RECT 118.590 144.265 120.510 144.435 ;
        RECT 118.590 144.245 118.910 144.265 ;
        RECT 118.140 143.585 118.470 144.095 ;
        RECT 118.740 143.635 118.910 144.245 ;
        RECT 120.680 144.095 120.850 144.605 ;
        RECT 121.020 144.535 121.200 144.945 ;
        RECT 121.370 144.355 121.540 145.115 ;
        RECT 119.080 143.375 119.410 144.065 ;
        RECT 119.640 143.925 120.850 144.095 ;
        RECT 121.020 144.045 121.540 144.355 ;
        RECT 121.710 144.945 122.130 145.285 ;
        RECT 122.420 144.945 122.830 145.275 ;
        RECT 121.710 144.175 121.900 144.945 ;
        RECT 123.000 144.815 123.170 145.545 ;
        RECT 124.315 145.375 124.485 145.705 ;
        RECT 124.655 145.545 124.985 145.925 ;
        RECT 123.340 144.995 123.690 145.365 ;
        RECT 123.000 144.775 123.420 144.815 ;
        RECT 122.070 144.605 123.420 144.775 ;
        RECT 122.070 144.445 122.320 144.605 ;
        RECT 122.830 144.175 123.080 144.435 ;
        RECT 121.710 143.925 123.080 144.175 ;
        RECT 119.640 143.635 119.880 143.925 ;
        RECT 120.680 143.845 120.850 143.925 ;
        RECT 120.080 143.375 120.500 143.755 ;
        RECT 120.680 143.595 121.310 143.845 ;
        RECT 121.780 143.375 122.110 143.755 ;
        RECT 122.280 143.635 122.450 143.925 ;
        RECT 123.250 143.760 123.420 144.605 ;
        RECT 123.870 144.435 124.090 145.305 ;
        RECT 124.315 145.185 125.010 145.375 ;
        RECT 123.590 144.055 124.090 144.435 ;
        RECT 124.260 144.385 124.670 145.005 ;
        RECT 124.840 144.215 125.010 145.185 ;
        RECT 124.315 144.045 125.010 144.215 ;
        RECT 122.630 143.375 123.010 143.755 ;
        RECT 123.250 143.590 124.080 143.760 ;
        RECT 124.315 143.545 124.485 144.045 ;
        RECT 124.655 143.375 124.985 143.875 ;
        RECT 125.200 143.545 125.425 145.665 ;
        RECT 125.595 145.545 125.925 145.925 ;
        RECT 126.095 145.375 126.265 145.665 ;
        RECT 125.600 145.205 126.265 145.375 ;
        RECT 125.600 144.215 125.830 145.205 ;
        RECT 126.525 145.175 127.735 145.925 ;
        RECT 126.000 144.385 126.350 145.035 ;
        RECT 126.525 144.465 127.045 145.005 ;
        RECT 127.215 144.635 127.735 145.175 ;
        RECT 125.600 144.045 126.265 144.215 ;
        RECT 125.595 143.375 125.925 143.875 ;
        RECT 126.095 143.545 126.265 144.045 ;
        RECT 126.525 143.375 127.735 144.465 ;
        RECT 14.660 143.205 127.820 143.375 ;
        RECT 14.745 142.115 15.955 143.205 ;
        RECT 14.745 141.405 15.265 141.945 ;
        RECT 15.435 141.575 15.955 142.115 ;
        RECT 16.125 142.115 18.715 143.205 ;
        RECT 16.125 141.595 17.335 142.115 ;
        RECT 18.945 142.065 19.155 143.205 ;
        RECT 19.325 142.055 19.655 143.035 ;
        RECT 19.825 142.065 20.055 143.205 ;
        RECT 20.270 142.065 20.605 143.035 ;
        RECT 20.775 142.065 20.945 143.205 ;
        RECT 21.115 142.865 23.145 143.035 ;
        RECT 17.505 141.425 18.715 141.945 ;
        RECT 14.745 140.655 15.955 141.405 ;
        RECT 16.125 140.655 18.715 141.425 ;
        RECT 18.945 140.655 19.155 141.475 ;
        RECT 19.325 141.455 19.575 142.055 ;
        RECT 19.745 141.645 20.075 141.895 ;
        RECT 19.325 140.825 19.655 141.455 ;
        RECT 19.825 140.655 20.055 141.475 ;
        RECT 20.270 141.395 20.440 142.065 ;
        RECT 21.115 141.895 21.285 142.865 ;
        RECT 20.610 141.565 20.865 141.895 ;
        RECT 21.090 141.565 21.285 141.895 ;
        RECT 21.455 142.525 22.580 142.695 ;
        RECT 20.695 141.395 20.865 141.565 ;
        RECT 21.455 141.395 21.625 142.525 ;
        RECT 20.270 140.825 20.525 141.395 ;
        RECT 20.695 141.225 21.625 141.395 ;
        RECT 21.795 142.185 22.805 142.355 ;
        RECT 21.795 141.385 21.965 142.185 ;
        RECT 21.450 141.190 21.625 141.225 ;
        RECT 20.695 140.655 21.025 141.055 ;
        RECT 21.450 140.825 21.980 141.190 ;
        RECT 22.170 141.165 22.445 141.985 ;
        RECT 22.165 140.995 22.445 141.165 ;
        RECT 22.170 140.825 22.445 140.995 ;
        RECT 22.615 140.825 22.805 142.185 ;
        RECT 22.975 142.200 23.145 142.865 ;
        RECT 23.315 142.445 23.485 143.205 ;
        RECT 23.720 142.445 24.235 142.855 ;
        RECT 22.975 142.010 23.725 142.200 ;
        RECT 23.895 141.635 24.235 142.445 ;
        RECT 24.405 142.040 24.695 143.205 ;
        RECT 25.415 142.275 25.585 143.035 ;
        RECT 25.765 142.445 26.095 143.205 ;
        RECT 25.415 142.105 26.080 142.275 ;
        RECT 26.265 142.130 26.535 143.035 ;
        RECT 25.910 141.960 26.080 142.105 ;
        RECT 23.005 141.465 24.235 141.635 ;
        RECT 25.345 141.555 25.675 141.925 ;
        RECT 25.910 141.630 26.195 141.960 ;
        RECT 22.985 140.655 23.495 141.190 ;
        RECT 23.715 140.860 23.960 141.465 ;
        RECT 24.405 140.655 24.695 141.380 ;
        RECT 25.910 141.375 26.080 141.630 ;
        RECT 25.415 141.205 26.080 141.375 ;
        RECT 26.365 141.330 26.535 142.130 ;
        RECT 26.705 142.115 29.295 143.205 ;
        RECT 26.705 141.595 27.915 142.115 ;
        RECT 29.505 142.065 29.735 143.205 ;
        RECT 29.905 142.055 30.235 143.035 ;
        RECT 30.405 142.065 30.615 143.205 ;
        RECT 30.885 142.065 31.115 143.205 ;
        RECT 31.285 142.055 31.615 143.035 ;
        RECT 31.785 142.065 31.995 143.205 ;
        RECT 28.085 141.425 29.295 141.945 ;
        RECT 29.485 141.645 29.815 141.895 ;
        RECT 25.415 140.825 25.585 141.205 ;
        RECT 25.765 140.655 26.095 141.035 ;
        RECT 26.275 140.825 26.535 141.330 ;
        RECT 26.705 140.655 29.295 141.425 ;
        RECT 29.505 140.655 29.735 141.475 ;
        RECT 29.985 141.455 30.235 142.055 ;
        RECT 30.865 141.645 31.195 141.895 ;
        RECT 29.905 140.825 30.235 141.455 ;
        RECT 30.405 140.655 30.615 141.475 ;
        RECT 30.885 140.655 31.115 141.475 ;
        RECT 31.365 141.455 31.615 142.055 ;
        RECT 32.230 142.015 32.485 142.895 ;
        RECT 32.655 142.065 32.960 143.205 ;
        RECT 33.300 142.825 33.630 143.205 ;
        RECT 33.810 142.655 33.980 142.945 ;
        RECT 34.150 142.745 34.400 143.205 ;
        RECT 33.180 142.485 33.980 142.655 ;
        RECT 34.570 142.695 35.440 143.035 ;
        RECT 31.285 140.825 31.615 141.455 ;
        RECT 31.785 140.655 31.995 141.475 ;
        RECT 32.230 141.365 32.440 142.015 ;
        RECT 33.180 141.895 33.350 142.485 ;
        RECT 34.570 142.315 34.740 142.695 ;
        RECT 35.675 142.575 35.845 143.035 ;
        RECT 36.015 142.745 36.385 143.205 ;
        RECT 36.680 142.605 36.850 142.945 ;
        RECT 37.020 142.775 37.350 143.205 ;
        RECT 37.585 142.605 37.755 142.945 ;
        RECT 33.520 142.145 34.740 142.315 ;
        RECT 34.910 142.235 35.370 142.525 ;
        RECT 35.675 142.405 36.235 142.575 ;
        RECT 36.680 142.435 37.755 142.605 ;
        RECT 37.925 142.705 38.605 143.035 ;
        RECT 38.820 142.705 39.070 143.035 ;
        RECT 39.240 142.745 39.490 143.205 ;
        RECT 36.065 142.265 36.235 142.405 ;
        RECT 34.910 142.225 35.875 142.235 ;
        RECT 34.570 142.055 34.740 142.145 ;
        RECT 35.200 142.065 35.875 142.225 ;
        RECT 32.610 141.865 33.350 141.895 ;
        RECT 32.610 141.565 33.525 141.865 ;
        RECT 33.200 141.390 33.525 141.565 ;
        RECT 32.230 140.835 32.485 141.365 ;
        RECT 32.655 140.655 32.960 141.115 ;
        RECT 33.205 141.035 33.525 141.390 ;
        RECT 33.695 141.605 34.235 141.975 ;
        RECT 34.570 141.885 34.975 142.055 ;
        RECT 33.695 141.205 33.935 141.605 ;
        RECT 34.415 141.435 34.635 141.715 ;
        RECT 34.105 141.265 34.635 141.435 ;
        RECT 34.105 141.035 34.275 141.265 ;
        RECT 34.805 141.105 34.975 141.885 ;
        RECT 35.145 141.275 35.495 141.895 ;
        RECT 35.665 141.275 35.875 142.065 ;
        RECT 36.065 142.095 37.565 142.265 ;
        RECT 36.065 141.405 36.235 142.095 ;
        RECT 37.925 141.925 38.095 142.705 ;
        RECT 38.900 142.575 39.070 142.705 ;
        RECT 36.405 141.755 38.095 141.925 ;
        RECT 38.265 142.145 38.730 142.535 ;
        RECT 38.900 142.405 39.295 142.575 ;
        RECT 36.405 141.575 36.575 141.755 ;
        RECT 33.205 140.865 34.275 141.035 ;
        RECT 34.445 140.655 34.635 141.095 ;
        RECT 34.805 140.825 35.755 141.105 ;
        RECT 36.065 141.015 36.325 141.405 ;
        RECT 36.745 141.335 37.535 141.585 ;
        RECT 35.975 140.845 36.325 141.015 ;
        RECT 36.535 140.655 36.865 141.115 ;
        RECT 37.740 141.045 37.910 141.755 ;
        RECT 38.265 141.555 38.435 142.145 ;
        RECT 38.080 141.335 38.435 141.555 ;
        RECT 38.605 141.335 38.955 141.955 ;
        RECT 39.125 141.045 39.295 142.405 ;
        RECT 39.660 142.235 39.985 143.020 ;
        RECT 39.465 141.185 39.925 142.235 ;
        RECT 37.740 140.875 38.595 141.045 ;
        RECT 38.800 140.875 39.295 141.045 ;
        RECT 39.465 140.655 39.795 141.015 ;
        RECT 40.155 140.915 40.325 143.035 ;
        RECT 40.495 142.705 40.825 143.205 ;
        RECT 40.995 142.535 41.250 143.035 ;
        RECT 40.500 142.365 41.250 142.535 ;
        RECT 40.500 141.375 40.730 142.365 ;
        RECT 40.900 141.545 41.250 142.195 ;
        RECT 41.425 142.130 41.695 143.035 ;
        RECT 41.865 142.445 42.195 143.205 ;
        RECT 42.375 142.275 42.545 143.035 ;
        RECT 40.500 141.205 41.250 141.375 ;
        RECT 40.495 140.655 40.825 141.035 ;
        RECT 40.995 140.915 41.250 141.205 ;
        RECT 41.425 141.330 41.595 142.130 ;
        RECT 41.880 142.105 42.545 142.275 ;
        RECT 43.010 142.235 43.340 143.035 ;
        RECT 43.510 142.405 43.840 143.205 ;
        RECT 44.140 142.235 44.470 143.035 ;
        RECT 45.115 142.405 45.365 143.205 ;
        RECT 41.880 141.960 42.050 142.105 ;
        RECT 43.010 142.065 45.445 142.235 ;
        RECT 45.635 142.065 45.805 143.205 ;
        RECT 45.975 142.065 46.315 143.035 ;
        RECT 46.690 142.235 47.020 143.035 ;
        RECT 47.190 142.405 47.520 143.205 ;
        RECT 47.820 142.235 48.150 143.035 ;
        RECT 48.795 142.405 49.045 143.205 ;
        RECT 46.690 142.065 49.125 142.235 ;
        RECT 49.315 142.065 49.485 143.205 ;
        RECT 49.655 142.065 49.995 143.035 ;
        RECT 41.765 141.630 42.050 141.960 ;
        RECT 41.880 141.375 42.050 141.630 ;
        RECT 42.285 141.555 42.615 141.925 ;
        RECT 42.805 141.645 43.155 141.895 ;
        RECT 43.340 141.435 43.510 142.065 ;
        RECT 43.680 141.645 44.010 141.845 ;
        RECT 44.180 141.645 44.510 141.845 ;
        RECT 44.680 141.645 45.100 141.845 ;
        RECT 45.275 141.815 45.445 142.065 ;
        RECT 45.275 141.645 45.970 141.815 ;
        RECT 41.425 140.825 41.685 141.330 ;
        RECT 41.880 141.205 42.545 141.375 ;
        RECT 41.865 140.655 42.195 141.035 ;
        RECT 42.375 140.825 42.545 141.205 ;
        RECT 43.010 140.825 43.510 141.435 ;
        RECT 44.140 141.305 45.365 141.475 ;
        RECT 46.140 141.455 46.315 142.065 ;
        RECT 46.485 141.645 46.835 141.895 ;
        RECT 44.140 140.825 44.470 141.305 ;
        RECT 44.640 140.655 44.865 141.115 ;
        RECT 45.035 140.825 45.365 141.305 ;
        RECT 45.555 140.655 45.805 141.455 ;
        RECT 45.975 140.825 46.315 141.455 ;
        RECT 47.020 141.435 47.190 142.065 ;
        RECT 47.360 141.645 47.690 141.845 ;
        RECT 47.860 141.645 48.190 141.845 ;
        RECT 48.360 141.645 48.780 141.845 ;
        RECT 48.955 141.815 49.125 142.065 ;
        RECT 48.955 141.645 49.650 141.815 ;
        RECT 46.690 140.825 47.190 141.435 ;
        RECT 47.820 141.305 49.045 141.475 ;
        RECT 49.820 141.455 49.995 142.065 ;
        RECT 50.165 142.040 50.455 143.205 ;
        RECT 50.630 142.695 52.285 142.985 ;
        RECT 50.630 142.355 52.220 142.525 ;
        RECT 52.455 142.405 52.735 143.205 ;
        RECT 50.630 142.065 50.950 142.355 ;
        RECT 52.050 142.235 52.220 142.355 ;
        RECT 51.145 142.015 51.860 142.185 ;
        RECT 52.050 142.065 52.775 142.235 ;
        RECT 52.945 142.065 53.215 143.035 ;
        RECT 47.820 140.825 48.150 141.305 ;
        RECT 48.320 140.655 48.545 141.115 ;
        RECT 48.715 140.825 49.045 141.305 ;
        RECT 49.235 140.655 49.485 141.455 ;
        RECT 49.655 140.825 49.995 141.455 ;
        RECT 50.165 140.655 50.455 141.380 ;
        RECT 50.630 141.325 50.980 141.895 ;
        RECT 51.150 141.565 51.860 142.015 ;
        RECT 52.605 141.895 52.775 142.065 ;
        RECT 52.030 141.565 52.435 141.895 ;
        RECT 52.605 141.565 52.875 141.895 ;
        RECT 52.605 141.395 52.775 141.565 ;
        RECT 51.165 141.225 52.775 141.395 ;
        RECT 53.045 141.330 53.215 142.065 ;
        RECT 53.385 142.115 55.975 143.205 ;
        RECT 53.385 141.595 54.595 142.115 ;
        RECT 56.145 142.065 56.485 143.035 ;
        RECT 56.655 142.065 56.825 143.205 ;
        RECT 57.095 142.405 57.345 143.205 ;
        RECT 57.990 142.235 58.320 143.035 ;
        RECT 58.620 142.405 58.950 143.205 ;
        RECT 59.120 142.235 59.450 143.035 ;
        RECT 57.015 142.065 59.450 142.235 ;
        RECT 60.745 142.445 61.260 142.855 ;
        RECT 61.495 142.445 61.665 143.205 ;
        RECT 61.835 142.865 63.865 143.035 ;
        RECT 54.765 141.425 55.975 141.945 ;
        RECT 50.635 140.655 50.965 141.155 ;
        RECT 51.165 140.875 51.335 141.225 ;
        RECT 51.535 140.655 51.865 141.055 ;
        RECT 52.035 140.875 52.205 141.225 ;
        RECT 52.375 140.655 52.755 141.055 ;
        RECT 52.945 140.985 53.215 141.330 ;
        RECT 53.385 140.655 55.975 141.425 ;
        RECT 56.145 141.505 56.320 142.065 ;
        RECT 57.015 141.815 57.185 142.065 ;
        RECT 56.490 141.645 57.185 141.815 ;
        RECT 57.360 141.645 57.780 141.845 ;
        RECT 57.950 141.645 58.280 141.845 ;
        RECT 58.450 141.645 58.780 141.845 ;
        RECT 56.145 141.455 56.375 141.505 ;
        RECT 56.145 140.825 56.485 141.455 ;
        RECT 56.655 140.655 56.905 141.455 ;
        RECT 57.095 141.305 58.320 141.475 ;
        RECT 57.095 140.825 57.425 141.305 ;
        RECT 57.595 140.655 57.820 141.115 ;
        RECT 57.990 140.825 58.320 141.305 ;
        RECT 58.950 141.435 59.120 142.065 ;
        RECT 59.305 141.645 59.655 141.895 ;
        RECT 60.745 141.635 61.085 142.445 ;
        RECT 61.835 142.200 62.005 142.865 ;
        RECT 62.400 142.525 63.525 142.695 ;
        RECT 61.255 142.010 62.005 142.200 ;
        RECT 62.175 142.185 63.185 142.355 ;
        RECT 60.745 141.465 61.975 141.635 ;
        RECT 58.950 140.825 59.450 141.435 ;
        RECT 61.020 140.860 61.265 141.465 ;
        RECT 61.485 140.655 61.995 141.190 ;
        RECT 62.175 140.825 62.365 142.185 ;
        RECT 62.535 141.505 62.810 141.985 ;
        RECT 62.535 141.335 62.815 141.505 ;
        RECT 63.015 141.385 63.185 142.185 ;
        RECT 63.355 141.395 63.525 142.525 ;
        RECT 63.695 141.895 63.865 142.865 ;
        RECT 64.035 142.065 64.205 143.205 ;
        RECT 64.375 142.065 64.710 143.035 ;
        RECT 63.695 141.565 63.890 141.895 ;
        RECT 64.115 141.565 64.370 141.895 ;
        RECT 64.115 141.395 64.285 141.565 ;
        RECT 64.540 141.395 64.710 142.065 ;
        RECT 62.535 140.825 62.810 141.335 ;
        RECT 63.355 141.225 64.285 141.395 ;
        RECT 63.355 141.190 63.530 141.225 ;
        RECT 63.000 140.825 63.530 141.190 ;
        RECT 63.955 140.655 64.285 141.055 ;
        RECT 64.455 140.825 64.710 141.395 ;
        RECT 65.260 142.225 65.515 142.895 ;
        RECT 65.695 142.405 65.980 143.205 ;
        RECT 66.160 142.485 66.490 142.995 ;
        RECT 65.260 141.365 65.440 142.225 ;
        RECT 66.160 141.895 66.410 142.485 ;
        RECT 66.760 142.335 66.930 142.945 ;
        RECT 67.100 142.515 67.430 143.205 ;
        RECT 67.660 142.655 67.900 142.945 ;
        RECT 68.100 142.825 68.520 143.205 ;
        RECT 68.700 142.735 69.330 142.985 ;
        RECT 69.800 142.825 70.130 143.205 ;
        RECT 68.700 142.655 68.870 142.735 ;
        RECT 70.300 142.655 70.470 142.945 ;
        RECT 70.650 142.825 71.030 143.205 ;
        RECT 71.270 142.820 72.100 142.990 ;
        RECT 67.660 142.485 68.870 142.655 ;
        RECT 65.610 141.565 66.410 141.895 ;
        RECT 65.260 141.165 65.515 141.365 ;
        RECT 65.175 140.995 65.515 141.165 ;
        RECT 65.260 140.835 65.515 140.995 ;
        RECT 65.695 140.655 65.980 141.115 ;
        RECT 66.160 140.915 66.410 141.565 ;
        RECT 66.610 142.315 66.930 142.335 ;
        RECT 66.610 142.145 68.530 142.315 ;
        RECT 66.610 141.250 66.800 142.145 ;
        RECT 68.700 141.975 68.870 142.485 ;
        RECT 69.040 142.225 69.560 142.535 ;
        RECT 66.970 141.805 68.870 141.975 ;
        RECT 66.970 141.745 67.300 141.805 ;
        RECT 67.450 141.575 67.780 141.635 ;
        RECT 67.120 141.305 67.780 141.575 ;
        RECT 66.610 140.920 66.930 141.250 ;
        RECT 67.110 140.655 67.770 141.135 ;
        RECT 67.970 141.045 68.140 141.805 ;
        RECT 69.040 141.635 69.220 142.045 ;
        RECT 68.310 141.465 68.640 141.585 ;
        RECT 69.390 141.465 69.560 142.225 ;
        RECT 68.310 141.295 69.560 141.465 ;
        RECT 69.730 142.405 71.100 142.655 ;
        RECT 69.730 141.635 69.920 142.405 ;
        RECT 70.850 142.145 71.100 142.405 ;
        RECT 70.090 141.975 70.340 142.135 ;
        RECT 71.270 141.975 71.440 142.820 ;
        RECT 72.335 142.535 72.505 143.035 ;
        RECT 72.675 142.705 73.005 143.205 ;
        RECT 71.610 142.145 72.110 142.525 ;
        RECT 72.335 142.365 73.030 142.535 ;
        RECT 70.090 141.805 71.440 141.975 ;
        RECT 71.020 141.765 71.440 141.805 ;
        RECT 69.730 141.295 70.150 141.635 ;
        RECT 70.440 141.305 70.850 141.635 ;
        RECT 67.970 140.875 68.820 141.045 ;
        RECT 69.380 140.655 69.700 141.115 ;
        RECT 69.900 140.865 70.150 141.295 ;
        RECT 70.440 140.655 70.850 141.095 ;
        RECT 71.020 141.035 71.190 141.765 ;
        RECT 71.360 141.215 71.710 141.585 ;
        RECT 71.890 141.275 72.110 142.145 ;
        RECT 72.280 141.575 72.690 142.195 ;
        RECT 72.860 141.395 73.030 142.365 ;
        RECT 72.335 141.205 73.030 141.395 ;
        RECT 71.020 140.835 72.035 141.035 ;
        RECT 72.335 140.875 72.505 141.205 ;
        RECT 72.675 140.655 73.005 141.035 ;
        RECT 73.220 140.915 73.445 143.035 ;
        RECT 73.615 142.705 73.945 143.205 ;
        RECT 74.115 142.535 74.285 143.035 ;
        RECT 73.620 142.365 74.285 142.535 ;
        RECT 73.620 141.375 73.850 142.365 ;
        RECT 74.020 141.545 74.370 142.195 ;
        RECT 74.545 142.115 75.755 143.205 ;
        RECT 74.545 141.575 75.065 142.115 ;
        RECT 75.925 142.040 76.215 143.205 ;
        RECT 76.385 142.065 76.655 143.035 ;
        RECT 76.865 142.405 77.145 143.205 ;
        RECT 77.315 142.695 78.970 142.985 ;
        RECT 77.380 142.355 78.970 142.525 ;
        RECT 77.380 142.235 77.550 142.355 ;
        RECT 76.825 142.065 77.550 142.235 ;
        RECT 75.235 141.405 75.755 141.945 ;
        RECT 73.620 141.205 74.285 141.375 ;
        RECT 73.615 140.655 73.945 141.035 ;
        RECT 74.115 140.915 74.285 141.205 ;
        RECT 74.545 140.655 75.755 141.405 ;
        RECT 75.925 140.655 76.215 141.380 ;
        RECT 76.385 141.330 76.555 142.065 ;
        RECT 76.825 141.895 76.995 142.065 ;
        RECT 77.740 142.015 78.455 142.185 ;
        RECT 78.650 142.065 78.970 142.355 ;
        RECT 79.145 142.065 79.415 143.035 ;
        RECT 79.625 142.405 79.905 143.205 ;
        RECT 80.075 142.695 81.730 142.985 ;
        RECT 80.140 142.355 81.730 142.525 ;
        RECT 80.140 142.235 80.310 142.355 ;
        RECT 79.585 142.065 80.310 142.235 ;
        RECT 76.725 141.565 76.995 141.895 ;
        RECT 77.165 141.565 77.570 141.895 ;
        RECT 77.740 141.565 78.450 142.015 ;
        RECT 76.825 141.395 76.995 141.565 ;
        RECT 76.385 140.985 76.655 141.330 ;
        RECT 76.825 141.225 78.435 141.395 ;
        RECT 78.620 141.325 78.970 141.895 ;
        RECT 79.145 141.330 79.315 142.065 ;
        RECT 79.585 141.895 79.755 142.065 ;
        RECT 79.485 141.565 79.755 141.895 ;
        RECT 79.925 141.565 80.330 141.895 ;
        RECT 80.500 141.565 81.210 142.185 ;
        RECT 81.410 142.065 81.730 142.355 ;
        RECT 81.905 142.065 82.245 143.035 ;
        RECT 82.415 142.065 82.585 143.205 ;
        RECT 82.855 142.405 83.105 143.205 ;
        RECT 83.750 142.235 84.080 143.035 ;
        RECT 84.380 142.405 84.710 143.205 ;
        RECT 84.880 142.235 85.210 143.035 ;
        RECT 86.050 142.770 91.395 143.205 ;
        RECT 82.775 142.065 85.210 142.235 ;
        RECT 79.585 141.395 79.755 141.565 ;
        RECT 76.845 140.655 77.225 141.055 ;
        RECT 77.395 140.875 77.565 141.225 ;
        RECT 77.735 140.655 78.065 141.055 ;
        RECT 78.265 140.875 78.435 141.225 ;
        RECT 78.635 140.655 78.965 141.155 ;
        RECT 79.145 140.985 79.415 141.330 ;
        RECT 79.585 141.225 81.195 141.395 ;
        RECT 81.380 141.325 81.730 141.895 ;
        RECT 81.905 141.505 82.080 142.065 ;
        RECT 82.775 141.815 82.945 142.065 ;
        RECT 82.250 141.645 82.945 141.815 ;
        RECT 83.120 141.645 83.540 141.845 ;
        RECT 83.710 141.645 84.040 141.845 ;
        RECT 84.210 141.645 84.540 141.845 ;
        RECT 81.905 141.455 82.135 141.505 ;
        RECT 79.605 140.655 79.985 141.055 ;
        RECT 80.155 140.875 80.325 141.225 ;
        RECT 80.495 140.655 80.825 141.055 ;
        RECT 81.025 140.875 81.195 141.225 ;
        RECT 81.395 140.655 81.725 141.155 ;
        RECT 81.905 140.825 82.245 141.455 ;
        RECT 82.415 140.655 82.665 141.455 ;
        RECT 82.855 141.305 84.080 141.475 ;
        RECT 82.855 140.825 83.185 141.305 ;
        RECT 83.355 140.655 83.580 141.115 ;
        RECT 83.750 140.825 84.080 141.305 ;
        RECT 84.710 141.435 84.880 142.065 ;
        RECT 85.065 141.645 85.415 141.895 ;
        RECT 87.640 141.520 87.990 142.770 ;
        RECT 91.655 142.275 91.825 143.035 ;
        RECT 92.005 142.445 92.335 143.205 ;
        RECT 91.655 142.105 92.320 142.275 ;
        RECT 92.505 142.130 92.775 143.035 ;
        RECT 84.710 140.825 85.210 141.435 ;
        RECT 89.470 141.200 89.810 142.030 ;
        RECT 92.150 141.960 92.320 142.105 ;
        RECT 91.585 141.555 91.915 141.925 ;
        RECT 92.150 141.630 92.435 141.960 ;
        RECT 92.150 141.375 92.320 141.630 ;
        RECT 91.655 141.205 92.320 141.375 ;
        RECT 92.605 141.330 92.775 142.130 ;
        RECT 93.035 142.275 93.205 143.035 ;
        RECT 93.385 142.445 93.715 143.205 ;
        RECT 93.035 142.105 93.700 142.275 ;
        RECT 93.885 142.130 94.155 143.035 ;
        RECT 93.530 141.960 93.700 142.105 ;
        RECT 92.965 141.555 93.295 141.925 ;
        RECT 93.530 141.630 93.815 141.960 ;
        RECT 93.530 141.375 93.700 141.630 ;
        RECT 86.050 140.655 91.395 141.200 ;
        RECT 91.655 140.825 91.825 141.205 ;
        RECT 92.005 140.655 92.335 141.035 ;
        RECT 92.515 140.825 92.775 141.330 ;
        RECT 93.035 141.205 93.700 141.375 ;
        RECT 93.985 141.330 94.155 142.130 ;
        RECT 94.325 142.115 95.995 143.205 ;
        RECT 96.170 142.770 101.515 143.205 ;
        RECT 94.325 141.595 95.075 142.115 ;
        RECT 95.245 141.425 95.995 141.945 ;
        RECT 97.760 141.520 98.110 142.770 ;
        RECT 101.685 142.040 101.975 143.205 ;
        RECT 102.145 142.115 103.355 143.205 ;
        RECT 103.525 142.115 107.035 143.205 ;
        RECT 107.205 142.445 107.720 142.855 ;
        RECT 107.955 142.445 108.125 143.205 ;
        RECT 108.295 142.865 110.325 143.035 ;
        RECT 93.035 140.825 93.205 141.205 ;
        RECT 93.385 140.655 93.715 141.035 ;
        RECT 93.895 140.825 94.155 141.330 ;
        RECT 94.325 140.655 95.995 141.425 ;
        RECT 99.590 141.200 99.930 142.030 ;
        RECT 102.145 141.575 102.665 142.115 ;
        RECT 102.835 141.405 103.355 141.945 ;
        RECT 103.525 141.595 105.215 142.115 ;
        RECT 105.385 141.425 107.035 141.945 ;
        RECT 107.205 141.635 107.545 142.445 ;
        RECT 108.295 142.200 108.465 142.865 ;
        RECT 108.860 142.525 109.985 142.695 ;
        RECT 107.715 142.010 108.465 142.200 ;
        RECT 108.635 142.185 109.645 142.355 ;
        RECT 107.205 141.465 108.435 141.635 ;
        RECT 96.170 140.655 101.515 141.200 ;
        RECT 101.685 140.655 101.975 141.380 ;
        RECT 102.145 140.655 103.355 141.405 ;
        RECT 103.525 140.655 107.035 141.425 ;
        RECT 107.480 140.860 107.725 141.465 ;
        RECT 107.945 140.655 108.455 141.190 ;
        RECT 108.635 140.825 108.825 142.185 ;
        RECT 108.995 141.845 109.270 141.985 ;
        RECT 108.995 141.675 109.275 141.845 ;
        RECT 108.995 140.825 109.270 141.675 ;
        RECT 109.475 141.385 109.645 142.185 ;
        RECT 109.815 141.395 109.985 142.525 ;
        RECT 110.155 141.895 110.325 142.865 ;
        RECT 110.495 142.065 110.665 143.205 ;
        RECT 110.835 142.065 111.170 143.035 ;
        RECT 110.155 141.565 110.350 141.895 ;
        RECT 110.575 141.565 110.830 141.895 ;
        RECT 110.575 141.395 110.745 141.565 ;
        RECT 111.000 141.395 111.170 142.065 ;
        RECT 111.805 142.115 113.475 143.205 ;
        RECT 111.805 141.595 112.555 142.115 ;
        RECT 113.685 142.065 113.915 143.205 ;
        RECT 114.085 142.055 114.415 143.035 ;
        RECT 114.585 142.065 114.795 143.205 ;
        RECT 115.400 142.525 115.655 142.895 ;
        RECT 115.315 142.355 115.655 142.525 ;
        RECT 115.835 142.405 116.120 143.205 ;
        RECT 116.300 142.485 116.630 142.995 ;
        RECT 115.400 142.225 115.655 142.355 ;
        RECT 112.725 141.425 113.475 141.945 ;
        RECT 113.665 141.645 113.995 141.895 ;
        RECT 109.815 141.225 110.745 141.395 ;
        RECT 109.815 141.190 109.990 141.225 ;
        RECT 109.460 140.825 109.990 141.190 ;
        RECT 110.415 140.655 110.745 141.055 ;
        RECT 110.915 140.825 111.170 141.395 ;
        RECT 111.805 140.655 113.475 141.425 ;
        RECT 113.685 140.655 113.915 141.475 ;
        RECT 114.165 141.455 114.415 142.055 ;
        RECT 114.085 140.825 114.415 141.455 ;
        RECT 114.585 140.655 114.795 141.475 ;
        RECT 115.400 141.365 115.580 142.225 ;
        RECT 116.300 141.895 116.550 142.485 ;
        RECT 116.900 142.335 117.070 142.945 ;
        RECT 117.240 142.515 117.570 143.205 ;
        RECT 117.800 142.655 118.040 142.945 ;
        RECT 118.240 142.825 118.660 143.205 ;
        RECT 118.840 142.735 119.470 142.985 ;
        RECT 119.940 142.825 120.270 143.205 ;
        RECT 118.840 142.655 119.010 142.735 ;
        RECT 120.440 142.655 120.610 142.945 ;
        RECT 120.790 142.825 121.170 143.205 ;
        RECT 121.410 142.820 122.240 142.990 ;
        RECT 117.800 142.485 119.010 142.655 ;
        RECT 115.750 141.565 116.550 141.895 ;
        RECT 115.400 140.835 115.655 141.365 ;
        RECT 115.835 140.655 116.120 141.115 ;
        RECT 116.300 140.915 116.550 141.565 ;
        RECT 116.750 142.315 117.070 142.335 ;
        RECT 116.750 142.145 118.670 142.315 ;
        RECT 116.750 141.250 116.940 142.145 ;
        RECT 118.840 141.975 119.010 142.485 ;
        RECT 119.180 142.225 119.700 142.535 ;
        RECT 117.110 141.805 119.010 141.975 ;
        RECT 117.110 141.745 117.440 141.805 ;
        RECT 117.590 141.575 117.920 141.635 ;
        RECT 117.260 141.305 117.920 141.575 ;
        RECT 116.750 140.920 117.070 141.250 ;
        RECT 117.250 140.655 117.910 141.135 ;
        RECT 118.110 141.045 118.280 141.805 ;
        RECT 119.180 141.635 119.360 142.045 ;
        RECT 118.450 141.465 118.780 141.585 ;
        RECT 119.530 141.465 119.700 142.225 ;
        RECT 118.450 141.295 119.700 141.465 ;
        RECT 119.870 142.405 121.240 142.655 ;
        RECT 119.870 141.635 120.060 142.405 ;
        RECT 120.990 142.145 121.240 142.405 ;
        RECT 120.230 141.975 120.480 142.135 ;
        RECT 121.410 141.975 121.580 142.820 ;
        RECT 122.475 142.535 122.645 143.035 ;
        RECT 122.815 142.705 123.145 143.205 ;
        RECT 121.750 142.145 122.250 142.525 ;
        RECT 122.475 142.365 123.170 142.535 ;
        RECT 120.230 141.805 121.580 141.975 ;
        RECT 121.160 141.765 121.580 141.805 ;
        RECT 119.870 141.295 120.290 141.635 ;
        RECT 120.580 141.305 120.990 141.635 ;
        RECT 118.110 140.875 118.960 141.045 ;
        RECT 119.520 140.655 119.840 141.115 ;
        RECT 120.040 140.865 120.290 141.295 ;
        RECT 120.580 140.655 120.990 141.095 ;
        RECT 121.160 141.035 121.330 141.765 ;
        RECT 121.500 141.215 121.850 141.585 ;
        RECT 122.030 141.275 122.250 142.145 ;
        RECT 122.420 141.575 122.830 142.195 ;
        RECT 123.000 141.395 123.170 142.365 ;
        RECT 122.475 141.205 123.170 141.395 ;
        RECT 121.160 140.835 122.175 141.035 ;
        RECT 122.475 140.875 122.645 141.205 ;
        RECT 122.815 140.655 123.145 141.035 ;
        RECT 123.360 140.915 123.585 143.035 ;
        RECT 123.755 142.705 124.085 143.205 ;
        RECT 124.255 142.535 124.425 143.035 ;
        RECT 123.760 142.365 124.425 142.535 ;
        RECT 123.760 141.375 123.990 142.365 ;
        RECT 124.160 141.545 124.510 142.195 ;
        RECT 124.685 142.115 126.355 143.205 ;
        RECT 126.525 142.115 127.735 143.205 ;
        RECT 124.685 141.595 125.435 142.115 ;
        RECT 125.605 141.425 126.355 141.945 ;
        RECT 126.525 141.575 127.045 142.115 ;
        RECT 123.760 141.205 124.425 141.375 ;
        RECT 123.755 140.655 124.085 141.035 ;
        RECT 124.255 140.915 124.425 141.205 ;
        RECT 124.685 140.655 126.355 141.425 ;
        RECT 127.215 141.405 127.735 141.945 ;
        RECT 126.525 140.655 127.735 141.405 ;
        RECT 14.660 140.485 127.820 140.655 ;
        RECT 14.745 139.735 15.955 140.485 ;
        RECT 16.590 139.940 21.935 140.485 ;
        RECT 22.110 139.940 27.455 140.485 ;
        RECT 27.630 139.940 32.975 140.485 ;
        RECT 14.745 139.195 15.265 139.735 ;
        RECT 15.435 139.025 15.955 139.565 ;
        RECT 14.745 137.935 15.955 139.025 ;
        RECT 18.180 138.370 18.530 139.620 ;
        RECT 20.010 139.110 20.350 139.940 ;
        RECT 23.700 138.370 24.050 139.620 ;
        RECT 25.530 139.110 25.870 139.940 ;
        RECT 29.220 138.370 29.570 139.620 ;
        RECT 31.050 139.110 31.390 139.940 ;
        RECT 33.150 139.745 33.405 140.315 ;
        RECT 33.575 140.085 33.905 140.485 ;
        RECT 34.330 139.950 34.860 140.315 ;
        RECT 34.330 139.915 34.505 139.950 ;
        RECT 33.575 139.745 34.505 139.915 ;
        RECT 33.150 139.075 33.320 139.745 ;
        RECT 33.575 139.575 33.745 139.745 ;
        RECT 33.490 139.245 33.745 139.575 ;
        RECT 33.970 139.245 34.165 139.575 ;
        RECT 16.590 137.935 21.935 138.370 ;
        RECT 22.110 137.935 27.455 138.370 ;
        RECT 27.630 137.935 32.975 138.370 ;
        RECT 33.150 138.105 33.485 139.075 ;
        RECT 33.655 137.935 33.825 139.075 ;
        RECT 33.995 138.275 34.165 139.245 ;
        RECT 34.335 138.615 34.505 139.745 ;
        RECT 34.675 138.955 34.845 139.755 ;
        RECT 35.050 139.465 35.325 140.315 ;
        RECT 35.045 139.295 35.325 139.465 ;
        RECT 35.050 139.155 35.325 139.295 ;
        RECT 35.495 138.955 35.685 140.315 ;
        RECT 35.865 139.950 36.375 140.485 ;
        RECT 36.595 139.675 36.840 140.280 ;
        RECT 37.285 139.760 37.575 140.485 ;
        RECT 37.750 139.940 43.095 140.485 ;
        RECT 35.885 139.505 37.115 139.675 ;
        RECT 34.675 138.785 35.685 138.955 ;
        RECT 35.855 138.940 36.605 139.130 ;
        RECT 34.335 138.445 35.460 138.615 ;
        RECT 35.855 138.275 36.025 138.940 ;
        RECT 36.775 138.695 37.115 139.505 ;
        RECT 33.995 138.105 36.025 138.275 ;
        RECT 36.195 137.935 36.365 138.695 ;
        RECT 36.600 138.285 37.115 138.695 ;
        RECT 37.285 137.935 37.575 139.100 ;
        RECT 39.340 138.370 39.690 139.620 ;
        RECT 41.170 139.110 41.510 139.940 ;
        RECT 43.265 139.810 43.535 140.155 ;
        RECT 43.725 140.085 44.105 140.485 ;
        RECT 44.275 139.915 44.445 140.265 ;
        RECT 44.615 140.085 44.945 140.485 ;
        RECT 45.145 139.915 45.315 140.265 ;
        RECT 45.515 139.985 45.845 140.485 ;
        RECT 43.265 139.075 43.435 139.810 ;
        RECT 43.705 139.745 45.315 139.915 ;
        RECT 43.705 139.575 43.875 139.745 ;
        RECT 43.605 139.245 43.875 139.575 ;
        RECT 44.045 139.245 44.450 139.575 ;
        RECT 43.705 139.075 43.875 139.245 ;
        RECT 44.620 139.125 45.330 139.575 ;
        RECT 45.500 139.245 45.850 139.815 ;
        RECT 46.025 139.685 46.365 140.315 ;
        RECT 46.535 139.685 46.785 140.485 ;
        RECT 46.975 139.835 47.305 140.315 ;
        RECT 47.475 140.025 47.700 140.485 ;
        RECT 47.870 139.835 48.200 140.315 ;
        RECT 46.025 139.125 46.200 139.685 ;
        RECT 46.975 139.665 48.200 139.835 ;
        RECT 48.830 139.705 49.330 140.315 ;
        RECT 50.165 139.715 51.835 140.485 ;
        RECT 52.010 139.940 57.355 140.485 ;
        RECT 46.370 139.325 47.065 139.495 ;
        RECT 37.750 137.935 43.095 138.370 ;
        RECT 43.265 138.105 43.535 139.075 ;
        RECT 43.705 138.905 44.430 139.075 ;
        RECT 44.620 138.955 45.335 139.125 ;
        RECT 46.025 139.075 46.255 139.125 ;
        RECT 46.895 139.075 47.065 139.325 ;
        RECT 47.240 139.295 47.660 139.495 ;
        RECT 47.830 139.295 48.160 139.495 ;
        RECT 48.330 139.295 48.660 139.495 ;
        RECT 48.830 139.075 49.000 139.705 ;
        RECT 49.185 139.245 49.535 139.495 ;
        RECT 44.260 138.785 44.430 138.905 ;
        RECT 45.530 138.785 45.850 139.075 ;
        RECT 43.745 137.935 44.025 138.735 ;
        RECT 44.260 138.615 45.850 138.785 ;
        RECT 44.195 138.155 45.850 138.445 ;
        RECT 46.025 138.105 46.365 139.075 ;
        RECT 46.535 137.935 46.705 139.075 ;
        RECT 46.895 138.905 49.330 139.075 ;
        RECT 46.975 137.935 47.225 138.735 ;
        RECT 47.870 138.105 48.200 138.905 ;
        RECT 48.500 137.935 48.830 138.735 ;
        RECT 49.000 138.105 49.330 138.905 ;
        RECT 50.165 139.025 50.915 139.545 ;
        RECT 51.085 139.195 51.835 139.715 ;
        RECT 50.165 137.935 51.835 139.025 ;
        RECT 53.600 138.370 53.950 139.620 ;
        RECT 55.430 139.110 55.770 139.940 ;
        RECT 57.525 139.685 57.865 140.315 ;
        RECT 58.035 139.685 58.285 140.485 ;
        RECT 58.475 139.835 58.805 140.315 ;
        RECT 58.975 140.025 59.200 140.485 ;
        RECT 59.370 139.835 59.700 140.315 ;
        RECT 57.525 139.635 57.755 139.685 ;
        RECT 58.475 139.665 59.700 139.835 ;
        RECT 60.330 139.705 60.830 140.315 ;
        RECT 61.205 139.715 62.875 140.485 ;
        RECT 63.045 139.760 63.335 140.485 ;
        RECT 63.505 139.735 64.715 140.485 ;
        RECT 57.525 139.075 57.700 139.635 ;
        RECT 57.870 139.325 58.565 139.495 ;
        RECT 58.395 139.075 58.565 139.325 ;
        RECT 58.740 139.295 59.160 139.495 ;
        RECT 59.330 139.295 59.660 139.495 ;
        RECT 59.830 139.295 60.160 139.495 ;
        RECT 60.330 139.075 60.500 139.705 ;
        RECT 60.685 139.245 61.035 139.495 ;
        RECT 52.010 137.935 57.355 138.370 ;
        RECT 57.525 138.105 57.865 139.075 ;
        RECT 58.035 137.935 58.205 139.075 ;
        RECT 58.395 138.905 60.830 139.075 ;
        RECT 58.475 137.935 58.725 138.735 ;
        RECT 59.370 138.105 59.700 138.905 ;
        RECT 60.000 137.935 60.330 138.735 ;
        RECT 60.500 138.105 60.830 138.905 ;
        RECT 61.205 139.025 61.955 139.545 ;
        RECT 62.125 139.195 62.875 139.715 ;
        RECT 61.205 137.935 62.875 139.025 ;
        RECT 63.045 137.935 63.335 139.100 ;
        RECT 63.505 139.025 64.025 139.565 ;
        RECT 64.195 139.195 64.715 139.735 ;
        RECT 64.885 139.715 68.395 140.485 ;
        RECT 64.885 139.025 66.575 139.545 ;
        RECT 66.745 139.195 68.395 139.715 ;
        RECT 68.605 139.665 68.835 140.485 ;
        RECT 69.005 139.685 69.335 140.315 ;
        RECT 68.585 139.245 68.915 139.495 ;
        RECT 69.085 139.085 69.335 139.685 ;
        RECT 69.505 139.665 69.715 140.485 ;
        RECT 69.945 139.735 71.155 140.485 ;
        RECT 71.415 139.935 71.585 140.315 ;
        RECT 71.765 140.105 72.095 140.485 ;
        RECT 71.415 139.765 72.080 139.935 ;
        RECT 72.275 139.810 72.535 140.315 ;
        RECT 63.505 137.935 64.715 139.025 ;
        RECT 64.885 137.935 68.395 139.025 ;
        RECT 68.605 137.935 68.835 139.075 ;
        RECT 69.005 138.105 69.335 139.085 ;
        RECT 69.505 137.935 69.715 139.075 ;
        RECT 69.945 139.025 70.465 139.565 ;
        RECT 70.635 139.195 71.155 139.735 ;
        RECT 71.345 139.215 71.675 139.585 ;
        RECT 71.910 139.510 72.080 139.765 ;
        RECT 71.910 139.180 72.195 139.510 ;
        RECT 71.910 139.035 72.080 139.180 ;
        RECT 69.945 137.935 71.155 139.025 ;
        RECT 71.415 138.865 72.080 139.035 ;
        RECT 72.365 139.010 72.535 139.810 ;
        RECT 72.705 139.735 73.915 140.485 ;
        RECT 71.415 138.105 71.585 138.865 ;
        RECT 71.765 137.935 72.095 138.695 ;
        RECT 72.265 138.105 72.535 139.010 ;
        RECT 72.705 139.025 73.225 139.565 ;
        RECT 73.395 139.195 73.915 139.735 ;
        RECT 74.085 139.715 77.595 140.485 ;
        RECT 77.770 139.940 83.115 140.485 ;
        RECT 83.290 139.940 88.635 140.485 ;
        RECT 74.085 139.025 75.775 139.545 ;
        RECT 75.945 139.195 77.595 139.715 ;
        RECT 72.705 137.935 73.915 139.025 ;
        RECT 74.085 137.935 77.595 139.025 ;
        RECT 79.360 138.370 79.710 139.620 ;
        RECT 81.190 139.110 81.530 139.940 ;
        RECT 84.880 138.370 85.230 139.620 ;
        RECT 86.710 139.110 87.050 139.940 ;
        RECT 88.805 139.760 89.095 140.485 ;
        RECT 89.640 140.145 89.895 140.305 ;
        RECT 89.555 139.975 89.895 140.145 ;
        RECT 90.075 140.025 90.360 140.485 ;
        RECT 89.640 139.775 89.895 139.975 ;
        RECT 77.770 137.935 83.115 138.370 ;
        RECT 83.290 137.935 88.635 138.370 ;
        RECT 88.805 137.935 89.095 139.100 ;
        RECT 89.640 138.915 89.820 139.775 ;
        RECT 90.540 139.575 90.790 140.225 ;
        RECT 89.990 139.245 90.790 139.575 ;
        RECT 89.640 138.245 89.895 138.915 ;
        RECT 90.075 137.935 90.360 138.735 ;
        RECT 90.540 138.655 90.790 139.245 ;
        RECT 90.990 139.890 91.310 140.220 ;
        RECT 91.490 140.005 92.150 140.485 ;
        RECT 92.350 140.095 93.200 140.265 ;
        RECT 90.990 138.995 91.180 139.890 ;
        RECT 91.500 139.565 92.160 139.835 ;
        RECT 91.830 139.505 92.160 139.565 ;
        RECT 91.350 139.335 91.680 139.395 ;
        RECT 92.350 139.335 92.520 140.095 ;
        RECT 93.760 140.025 94.080 140.485 ;
        RECT 94.280 139.845 94.530 140.275 ;
        RECT 94.820 140.045 95.230 140.485 ;
        RECT 95.400 140.105 96.415 140.305 ;
        RECT 92.690 139.675 93.940 139.845 ;
        RECT 92.690 139.555 93.020 139.675 ;
        RECT 91.350 139.165 93.250 139.335 ;
        RECT 90.990 138.825 92.910 138.995 ;
        RECT 90.990 138.805 91.310 138.825 ;
        RECT 90.540 138.145 90.870 138.655 ;
        RECT 91.140 138.195 91.310 138.805 ;
        RECT 93.080 138.655 93.250 139.165 ;
        RECT 93.420 139.095 93.600 139.505 ;
        RECT 93.770 138.915 93.940 139.675 ;
        RECT 91.480 137.935 91.810 138.625 ;
        RECT 92.040 138.485 93.250 138.655 ;
        RECT 93.420 138.605 93.940 138.915 ;
        RECT 94.110 139.505 94.530 139.845 ;
        RECT 94.820 139.505 95.230 139.835 ;
        RECT 94.110 138.735 94.300 139.505 ;
        RECT 95.400 139.375 95.570 140.105 ;
        RECT 96.715 139.935 96.885 140.265 ;
        RECT 97.055 140.105 97.385 140.485 ;
        RECT 95.740 139.555 96.090 139.925 ;
        RECT 95.400 139.335 95.820 139.375 ;
        RECT 94.470 139.165 95.820 139.335 ;
        RECT 94.470 139.005 94.720 139.165 ;
        RECT 95.230 138.735 95.480 138.995 ;
        RECT 94.110 138.485 95.480 138.735 ;
        RECT 92.040 138.195 92.280 138.485 ;
        RECT 93.080 138.405 93.250 138.485 ;
        RECT 92.480 137.935 92.900 138.315 ;
        RECT 93.080 138.155 93.710 138.405 ;
        RECT 94.180 137.935 94.510 138.315 ;
        RECT 94.680 138.195 94.850 138.485 ;
        RECT 95.650 138.320 95.820 139.165 ;
        RECT 96.270 138.995 96.490 139.865 ;
        RECT 96.715 139.745 97.410 139.935 ;
        RECT 95.990 138.615 96.490 138.995 ;
        RECT 96.660 138.945 97.070 139.565 ;
        RECT 97.240 138.775 97.410 139.745 ;
        RECT 96.715 138.605 97.410 138.775 ;
        RECT 95.030 137.935 95.410 138.315 ;
        RECT 95.650 138.150 96.480 138.320 ;
        RECT 96.715 138.105 96.885 138.605 ;
        RECT 97.055 137.935 97.385 138.435 ;
        RECT 97.600 138.105 97.825 140.225 ;
        RECT 97.995 140.105 98.325 140.485 ;
        RECT 98.495 139.935 98.665 140.225 ;
        RECT 98.000 139.765 98.665 139.935 ;
        RECT 98.000 138.775 98.230 139.765 ;
        RECT 99.845 139.715 103.355 140.485 ;
        RECT 98.400 138.945 98.750 139.595 ;
        RECT 99.845 139.025 101.535 139.545 ;
        RECT 101.705 139.195 103.355 139.715 ;
        RECT 103.900 139.775 104.155 140.305 ;
        RECT 104.335 140.025 104.620 140.485 ;
        RECT 98.000 138.605 98.665 138.775 ;
        RECT 97.995 137.935 98.325 138.435 ;
        RECT 98.495 138.105 98.665 138.605 ;
        RECT 99.845 137.935 103.355 139.025 ;
        RECT 103.900 138.915 104.080 139.775 ;
        RECT 104.800 139.575 105.050 140.225 ;
        RECT 104.250 139.245 105.050 139.575 ;
        RECT 103.900 138.445 104.155 138.915 ;
        RECT 103.815 138.275 104.155 138.445 ;
        RECT 103.900 138.245 104.155 138.275 ;
        RECT 104.335 137.935 104.620 138.735 ;
        RECT 104.800 138.655 105.050 139.245 ;
        RECT 105.250 139.890 105.570 140.220 ;
        RECT 105.750 140.005 106.410 140.485 ;
        RECT 106.610 140.095 107.460 140.265 ;
        RECT 105.250 138.995 105.440 139.890 ;
        RECT 105.760 139.565 106.420 139.835 ;
        RECT 106.090 139.505 106.420 139.565 ;
        RECT 105.610 139.335 105.940 139.395 ;
        RECT 106.610 139.335 106.780 140.095 ;
        RECT 108.020 140.025 108.340 140.485 ;
        RECT 108.540 139.845 108.790 140.275 ;
        RECT 109.080 140.045 109.490 140.485 ;
        RECT 109.660 140.105 110.675 140.305 ;
        RECT 106.950 139.675 108.200 139.845 ;
        RECT 106.950 139.555 107.280 139.675 ;
        RECT 105.610 139.165 107.510 139.335 ;
        RECT 105.250 138.825 107.170 138.995 ;
        RECT 105.250 138.805 105.570 138.825 ;
        RECT 104.800 138.145 105.130 138.655 ;
        RECT 105.400 138.195 105.570 138.805 ;
        RECT 107.340 138.655 107.510 139.165 ;
        RECT 107.680 139.095 107.860 139.505 ;
        RECT 108.030 138.915 108.200 139.675 ;
        RECT 105.740 137.935 106.070 138.625 ;
        RECT 106.300 138.485 107.510 138.655 ;
        RECT 107.680 138.605 108.200 138.915 ;
        RECT 108.370 139.505 108.790 139.845 ;
        RECT 109.080 139.505 109.490 139.835 ;
        RECT 108.370 138.735 108.560 139.505 ;
        RECT 109.660 139.375 109.830 140.105 ;
        RECT 110.975 139.935 111.145 140.265 ;
        RECT 111.315 140.105 111.645 140.485 ;
        RECT 110.000 139.555 110.350 139.925 ;
        RECT 109.660 139.335 110.080 139.375 ;
        RECT 108.730 139.165 110.080 139.335 ;
        RECT 108.730 139.005 108.980 139.165 ;
        RECT 109.490 138.735 109.740 138.995 ;
        RECT 108.370 138.485 109.740 138.735 ;
        RECT 106.300 138.195 106.540 138.485 ;
        RECT 107.340 138.405 107.510 138.485 ;
        RECT 106.740 137.935 107.160 138.315 ;
        RECT 107.340 138.155 107.970 138.405 ;
        RECT 108.440 137.935 108.770 138.315 ;
        RECT 108.940 138.195 109.110 138.485 ;
        RECT 109.910 138.320 110.080 139.165 ;
        RECT 110.530 138.995 110.750 139.865 ;
        RECT 110.975 139.745 111.670 139.935 ;
        RECT 110.250 138.615 110.750 138.995 ;
        RECT 110.920 138.945 111.330 139.565 ;
        RECT 111.500 138.775 111.670 139.745 ;
        RECT 110.975 138.605 111.670 138.775 ;
        RECT 109.290 137.935 109.670 138.315 ;
        RECT 109.910 138.150 110.740 138.320 ;
        RECT 110.975 138.105 111.145 138.605 ;
        RECT 111.315 137.935 111.645 138.435 ;
        RECT 111.860 138.105 112.085 140.225 ;
        RECT 112.255 140.105 112.585 140.485 ;
        RECT 112.755 139.935 112.925 140.225 ;
        RECT 112.260 139.765 112.925 139.935 ;
        RECT 112.260 138.775 112.490 139.765 ;
        RECT 113.185 139.735 114.395 140.485 ;
        RECT 114.565 139.760 114.855 140.485 ;
        RECT 112.660 138.945 113.010 139.595 ;
        RECT 113.185 139.025 113.705 139.565 ;
        RECT 113.875 139.195 114.395 139.735 ;
        RECT 115.760 139.675 116.005 140.280 ;
        RECT 116.225 139.950 116.735 140.485 ;
        RECT 115.485 139.505 116.715 139.675 ;
        RECT 112.260 138.605 112.925 138.775 ;
        RECT 112.255 137.935 112.585 138.435 ;
        RECT 112.755 138.105 112.925 138.605 ;
        RECT 113.185 137.935 114.395 139.025 ;
        RECT 114.565 137.935 114.855 139.100 ;
        RECT 115.485 138.695 115.825 139.505 ;
        RECT 115.995 138.940 116.745 139.130 ;
        RECT 115.485 138.285 116.000 138.695 ;
        RECT 116.235 137.935 116.405 138.695 ;
        RECT 116.575 138.275 116.745 138.940 ;
        RECT 116.915 138.955 117.105 140.315 ;
        RECT 117.275 140.145 117.550 140.315 ;
        RECT 117.275 139.975 117.555 140.145 ;
        RECT 117.275 139.155 117.550 139.975 ;
        RECT 117.740 139.950 118.270 140.315 ;
        RECT 118.695 140.085 119.025 140.485 ;
        RECT 118.095 139.915 118.270 139.950 ;
        RECT 117.755 138.955 117.925 139.755 ;
        RECT 116.915 138.785 117.925 138.955 ;
        RECT 118.095 139.745 119.025 139.915 ;
        RECT 119.195 139.745 119.450 140.315 ;
        RECT 120.175 139.935 120.345 140.315 ;
        RECT 120.525 140.105 120.855 140.485 ;
        RECT 120.175 139.765 120.840 139.935 ;
        RECT 121.035 139.810 121.295 140.315 ;
        RECT 118.095 138.615 118.265 139.745 ;
        RECT 118.855 139.575 119.025 139.745 ;
        RECT 117.140 138.445 118.265 138.615 ;
        RECT 118.435 139.245 118.630 139.575 ;
        RECT 118.855 139.245 119.110 139.575 ;
        RECT 118.435 138.275 118.605 139.245 ;
        RECT 119.280 139.075 119.450 139.745 ;
        RECT 120.105 139.215 120.435 139.585 ;
        RECT 120.670 139.510 120.840 139.765 ;
        RECT 116.575 138.105 118.605 138.275 ;
        RECT 118.775 137.935 118.945 139.075 ;
        RECT 119.115 138.105 119.450 139.075 ;
        RECT 120.670 139.180 120.955 139.510 ;
        RECT 120.670 139.035 120.840 139.180 ;
        RECT 120.175 138.865 120.840 139.035 ;
        RECT 121.125 139.010 121.295 139.810 ;
        RECT 121.465 139.735 122.675 140.485 ;
        RECT 120.175 138.105 120.345 138.865 ;
        RECT 120.525 137.935 120.855 138.695 ;
        RECT 121.025 138.105 121.295 139.010 ;
        RECT 121.465 139.025 121.985 139.565 ;
        RECT 122.155 139.195 122.675 139.735 ;
        RECT 122.845 139.715 126.355 140.485 ;
        RECT 126.525 139.735 127.735 140.485 ;
        RECT 122.845 139.025 124.535 139.545 ;
        RECT 124.705 139.195 126.355 139.715 ;
        RECT 126.525 139.025 127.045 139.565 ;
        RECT 127.215 139.195 127.735 139.735 ;
        RECT 121.465 137.935 122.675 139.025 ;
        RECT 122.845 137.935 126.355 139.025 ;
        RECT 126.525 137.935 127.735 139.025 ;
        RECT 14.660 137.765 127.820 137.935 ;
        RECT 14.745 136.675 15.955 137.765 ;
        RECT 14.745 135.965 15.265 136.505 ;
        RECT 15.435 136.135 15.955 136.675 ;
        RECT 16.125 136.675 18.715 137.765 ;
        RECT 18.890 137.330 24.235 137.765 ;
        RECT 16.125 136.155 17.335 136.675 ;
        RECT 17.505 135.985 18.715 136.505 ;
        RECT 20.480 136.080 20.830 137.330 ;
        RECT 24.405 136.600 24.695 137.765 ;
        RECT 25.330 137.330 30.675 137.765 ;
        RECT 30.850 137.330 36.195 137.765 ;
        RECT 36.370 137.330 41.715 137.765 ;
        RECT 41.890 137.330 47.235 137.765 ;
        RECT 14.745 135.215 15.955 135.965 ;
        RECT 16.125 135.215 18.715 135.985 ;
        RECT 22.310 135.760 22.650 136.590 ;
        RECT 26.920 136.080 27.270 137.330 ;
        RECT 18.890 135.215 24.235 135.760 ;
        RECT 24.405 135.215 24.695 135.940 ;
        RECT 28.750 135.760 29.090 136.590 ;
        RECT 32.440 136.080 32.790 137.330 ;
        RECT 34.270 135.760 34.610 136.590 ;
        RECT 37.960 136.080 38.310 137.330 ;
        RECT 39.790 135.760 40.130 136.590 ;
        RECT 43.480 136.080 43.830 137.330 ;
        RECT 47.605 137.095 47.885 137.765 ;
        RECT 48.055 136.875 48.355 137.425 ;
        RECT 48.555 137.045 48.885 137.765 ;
        RECT 49.075 137.045 49.535 137.595 ;
        RECT 45.310 135.760 45.650 136.590 ;
        RECT 47.420 136.455 47.685 136.815 ;
        RECT 48.055 136.705 48.995 136.875 ;
        RECT 48.825 136.455 48.995 136.705 ;
        RECT 47.420 136.205 48.095 136.455 ;
        RECT 48.315 136.205 48.655 136.455 ;
        RECT 48.825 136.125 49.115 136.455 ;
        RECT 48.825 136.035 48.995 136.125 ;
        RECT 47.605 135.845 48.995 136.035 ;
        RECT 25.330 135.215 30.675 135.760 ;
        RECT 30.850 135.215 36.195 135.760 ;
        RECT 36.370 135.215 41.715 135.760 ;
        RECT 41.890 135.215 47.235 135.760 ;
        RECT 47.605 135.485 47.935 135.845 ;
        RECT 49.285 135.675 49.535 137.045 ;
        RECT 50.165 136.600 50.455 137.765 ;
        RECT 51.090 137.330 56.435 137.765 ;
        RECT 56.610 137.330 61.955 137.765 ;
        RECT 52.680 136.080 53.030 137.330 ;
        RECT 48.555 135.215 48.805 135.675 ;
        RECT 48.975 135.385 49.535 135.675 ;
        RECT 50.165 135.215 50.455 135.940 ;
        RECT 54.510 135.760 54.850 136.590 ;
        RECT 58.200 136.080 58.550 137.330 ;
        RECT 62.125 137.005 62.640 137.415 ;
        RECT 62.875 137.005 63.045 137.765 ;
        RECT 63.215 137.425 65.245 137.595 ;
        RECT 60.030 135.760 60.370 136.590 ;
        RECT 62.125 136.195 62.465 137.005 ;
        RECT 63.215 136.760 63.385 137.425 ;
        RECT 63.780 137.085 64.905 137.255 ;
        RECT 62.635 136.570 63.385 136.760 ;
        RECT 63.555 136.745 64.565 136.915 ;
        RECT 62.125 136.025 63.355 136.195 ;
        RECT 51.090 135.215 56.435 135.760 ;
        RECT 56.610 135.215 61.955 135.760 ;
        RECT 62.400 135.420 62.645 136.025 ;
        RECT 62.865 135.215 63.375 135.750 ;
        RECT 63.555 135.385 63.745 136.745 ;
        RECT 63.915 136.405 64.190 136.545 ;
        RECT 63.915 136.235 64.195 136.405 ;
        RECT 63.915 135.385 64.190 136.235 ;
        RECT 64.395 135.945 64.565 136.745 ;
        RECT 64.735 135.955 64.905 137.085 ;
        RECT 65.075 136.455 65.245 137.425 ;
        RECT 65.415 136.625 65.585 137.765 ;
        RECT 65.755 136.625 66.090 137.595 ;
        RECT 65.075 136.125 65.270 136.455 ;
        RECT 65.495 136.125 65.750 136.455 ;
        RECT 65.495 135.955 65.665 136.125 ;
        RECT 65.920 135.955 66.090 136.625 ;
        RECT 64.735 135.785 65.665 135.955 ;
        RECT 64.735 135.750 64.910 135.785 ;
        RECT 64.380 135.385 64.910 135.750 ;
        RECT 65.335 135.215 65.665 135.615 ;
        RECT 65.835 135.385 66.090 135.955 ;
        RECT 66.640 136.785 66.895 137.455 ;
        RECT 67.075 136.965 67.360 137.765 ;
        RECT 67.540 137.045 67.870 137.555 ;
        RECT 66.640 135.925 66.820 136.785 ;
        RECT 67.540 136.455 67.790 137.045 ;
        RECT 68.140 136.895 68.310 137.505 ;
        RECT 68.480 137.075 68.810 137.765 ;
        RECT 69.040 137.215 69.280 137.505 ;
        RECT 69.480 137.385 69.900 137.765 ;
        RECT 70.080 137.295 70.710 137.545 ;
        RECT 71.180 137.385 71.510 137.765 ;
        RECT 70.080 137.215 70.250 137.295 ;
        RECT 71.680 137.215 71.850 137.505 ;
        RECT 72.030 137.385 72.410 137.765 ;
        RECT 72.650 137.380 73.480 137.550 ;
        RECT 69.040 137.045 70.250 137.215 ;
        RECT 66.990 136.125 67.790 136.455 ;
        RECT 66.640 135.725 66.895 135.925 ;
        RECT 66.555 135.555 66.895 135.725 ;
        RECT 66.640 135.395 66.895 135.555 ;
        RECT 67.075 135.215 67.360 135.675 ;
        RECT 67.540 135.475 67.790 136.125 ;
        RECT 67.990 136.875 68.310 136.895 ;
        RECT 67.990 136.705 69.910 136.875 ;
        RECT 67.990 135.810 68.180 136.705 ;
        RECT 70.080 136.535 70.250 137.045 ;
        RECT 70.420 136.785 70.940 137.095 ;
        RECT 68.350 136.365 70.250 136.535 ;
        RECT 68.350 136.305 68.680 136.365 ;
        RECT 68.830 136.135 69.160 136.195 ;
        RECT 68.500 135.865 69.160 136.135 ;
        RECT 67.990 135.480 68.310 135.810 ;
        RECT 68.490 135.215 69.150 135.695 ;
        RECT 69.350 135.605 69.520 136.365 ;
        RECT 70.420 136.195 70.600 136.605 ;
        RECT 69.690 136.025 70.020 136.145 ;
        RECT 70.770 136.025 70.940 136.785 ;
        RECT 69.690 135.855 70.940 136.025 ;
        RECT 71.110 136.965 72.480 137.215 ;
        RECT 71.110 136.195 71.300 136.965 ;
        RECT 72.230 136.705 72.480 136.965 ;
        RECT 71.470 136.535 71.720 136.695 ;
        RECT 72.650 136.535 72.820 137.380 ;
        RECT 73.715 137.095 73.885 137.595 ;
        RECT 74.055 137.265 74.385 137.765 ;
        RECT 72.990 136.705 73.490 137.085 ;
        RECT 73.715 136.925 74.410 137.095 ;
        RECT 71.470 136.365 72.820 136.535 ;
        RECT 72.400 136.325 72.820 136.365 ;
        RECT 71.110 135.855 71.530 136.195 ;
        RECT 71.820 135.865 72.230 136.195 ;
        RECT 69.350 135.435 70.200 135.605 ;
        RECT 70.760 135.215 71.080 135.675 ;
        RECT 71.280 135.425 71.530 135.855 ;
        RECT 71.820 135.215 72.230 135.655 ;
        RECT 72.400 135.595 72.570 136.325 ;
        RECT 72.740 135.775 73.090 136.145 ;
        RECT 73.270 135.835 73.490 136.705 ;
        RECT 73.660 136.135 74.070 136.755 ;
        RECT 74.240 135.955 74.410 136.925 ;
        RECT 73.715 135.765 74.410 135.955 ;
        RECT 72.400 135.395 73.415 135.595 ;
        RECT 73.715 135.435 73.885 135.765 ;
        RECT 74.055 135.215 74.385 135.595 ;
        RECT 74.600 135.475 74.825 137.595 ;
        RECT 74.995 137.265 75.325 137.765 ;
        RECT 75.495 137.095 75.665 137.595 ;
        RECT 75.000 136.925 75.665 137.095 ;
        RECT 75.000 135.935 75.230 136.925 ;
        RECT 75.400 136.105 75.750 136.755 ;
        RECT 75.925 136.600 76.215 137.765 ;
        RECT 77.305 136.675 80.815 137.765 ;
        RECT 80.990 137.255 82.645 137.545 ;
        RECT 80.990 136.915 82.580 137.085 ;
        RECT 82.815 136.965 83.095 137.765 ;
        RECT 77.305 136.155 78.995 136.675 ;
        RECT 80.990 136.625 81.310 136.915 ;
        RECT 82.410 136.795 82.580 136.915 ;
        RECT 81.505 136.575 82.220 136.745 ;
        RECT 82.410 136.625 83.135 136.795 ;
        RECT 83.305 136.625 83.575 137.595 ;
        RECT 79.165 135.985 80.815 136.505 ;
        RECT 75.000 135.765 75.665 135.935 ;
        RECT 74.995 135.215 75.325 135.595 ;
        RECT 75.495 135.475 75.665 135.765 ;
        RECT 75.925 135.215 76.215 135.940 ;
        RECT 77.305 135.215 80.815 135.985 ;
        RECT 80.990 135.885 81.340 136.455 ;
        RECT 81.510 136.125 82.220 136.575 ;
        RECT 82.965 136.455 83.135 136.625 ;
        RECT 82.390 136.125 82.795 136.455 ;
        RECT 82.965 136.125 83.235 136.455 ;
        RECT 82.965 135.955 83.135 136.125 ;
        RECT 81.525 135.785 83.135 135.955 ;
        RECT 83.405 135.890 83.575 136.625 ;
        RECT 84.665 136.675 88.175 137.765 ;
        RECT 88.345 137.005 88.860 137.415 ;
        RECT 89.095 137.005 89.265 137.765 ;
        RECT 89.435 137.425 91.465 137.595 ;
        RECT 84.665 136.155 86.355 136.675 ;
        RECT 86.525 135.985 88.175 136.505 ;
        RECT 88.345 136.195 88.685 137.005 ;
        RECT 89.435 136.760 89.605 137.425 ;
        RECT 90.000 137.085 91.125 137.255 ;
        RECT 88.855 136.570 89.605 136.760 ;
        RECT 89.775 136.745 90.785 136.915 ;
        RECT 88.345 136.025 89.575 136.195 ;
        RECT 80.995 135.215 81.325 135.715 ;
        RECT 81.525 135.435 81.695 135.785 ;
        RECT 81.895 135.215 82.225 135.615 ;
        RECT 82.395 135.435 82.565 135.785 ;
        RECT 82.735 135.215 83.115 135.615 ;
        RECT 83.305 135.545 83.575 135.890 ;
        RECT 84.665 135.215 88.175 135.985 ;
        RECT 88.620 135.420 88.865 136.025 ;
        RECT 89.085 135.215 89.595 135.750 ;
        RECT 89.775 135.385 89.965 136.745 ;
        RECT 90.135 135.725 90.410 136.545 ;
        RECT 90.615 135.945 90.785 136.745 ;
        RECT 90.955 135.955 91.125 137.085 ;
        RECT 91.295 136.455 91.465 137.425 ;
        RECT 91.635 136.625 91.805 137.765 ;
        RECT 91.975 136.625 92.310 137.595 ;
        RECT 92.545 136.625 92.755 137.765 ;
        RECT 91.295 136.125 91.490 136.455 ;
        RECT 91.715 136.125 91.970 136.455 ;
        RECT 91.715 135.955 91.885 136.125 ;
        RECT 92.140 135.955 92.310 136.625 ;
        RECT 92.925 136.615 93.255 137.595 ;
        RECT 93.425 136.625 93.655 137.765 ;
        RECT 93.865 136.675 97.375 137.765 ;
        RECT 97.545 137.005 98.060 137.415 ;
        RECT 98.295 137.005 98.465 137.765 ;
        RECT 98.635 137.425 100.665 137.595 ;
        RECT 90.955 135.785 91.885 135.955 ;
        RECT 90.955 135.750 91.130 135.785 ;
        RECT 90.135 135.555 90.415 135.725 ;
        RECT 90.135 135.385 90.410 135.555 ;
        RECT 90.600 135.385 91.130 135.750 ;
        RECT 91.555 135.215 91.885 135.615 ;
        RECT 92.055 135.385 92.310 135.955 ;
        RECT 92.545 135.215 92.755 136.035 ;
        RECT 92.925 136.015 93.175 136.615 ;
        RECT 93.345 136.205 93.675 136.455 ;
        RECT 93.865 136.155 95.555 136.675 ;
        RECT 92.925 135.385 93.255 136.015 ;
        RECT 93.425 135.215 93.655 136.035 ;
        RECT 95.725 135.985 97.375 136.505 ;
        RECT 97.545 136.195 97.885 137.005 ;
        RECT 98.635 136.760 98.805 137.425 ;
        RECT 99.200 137.085 100.325 137.255 ;
        RECT 98.055 136.570 98.805 136.760 ;
        RECT 98.975 136.745 99.985 136.915 ;
        RECT 97.545 136.025 98.775 136.195 ;
        RECT 93.865 135.215 97.375 135.985 ;
        RECT 97.820 135.420 98.065 136.025 ;
        RECT 98.285 135.215 98.795 135.750 ;
        RECT 98.975 135.385 99.165 136.745 ;
        RECT 99.335 136.405 99.610 136.545 ;
        RECT 99.335 136.235 99.615 136.405 ;
        RECT 99.335 135.385 99.610 136.235 ;
        RECT 99.815 135.945 99.985 136.745 ;
        RECT 100.155 135.955 100.325 137.085 ;
        RECT 100.495 136.455 100.665 137.425 ;
        RECT 100.835 136.625 101.005 137.765 ;
        RECT 101.175 136.625 101.510 137.595 ;
        RECT 100.495 136.125 100.690 136.455 ;
        RECT 100.915 136.125 101.170 136.455 ;
        RECT 100.915 135.955 101.085 136.125 ;
        RECT 101.340 135.955 101.510 136.625 ;
        RECT 101.685 136.600 101.975 137.765 ;
        RECT 102.145 136.675 103.815 137.765 ;
        RECT 104.075 136.835 104.245 137.595 ;
        RECT 104.425 137.005 104.755 137.765 ;
        RECT 102.145 136.155 102.895 136.675 ;
        RECT 104.075 136.665 104.740 136.835 ;
        RECT 104.925 136.690 105.195 137.595 ;
        RECT 104.570 136.520 104.740 136.665 ;
        RECT 103.065 135.985 103.815 136.505 ;
        RECT 104.005 136.115 104.335 136.485 ;
        RECT 104.570 136.190 104.855 136.520 ;
        RECT 100.155 135.785 101.085 135.955 ;
        RECT 100.155 135.750 100.330 135.785 ;
        RECT 99.800 135.385 100.330 135.750 ;
        RECT 100.755 135.215 101.085 135.615 ;
        RECT 101.255 135.385 101.510 135.955 ;
        RECT 101.685 135.215 101.975 135.940 ;
        RECT 102.145 135.215 103.815 135.985 ;
        RECT 104.570 135.935 104.740 136.190 ;
        RECT 104.075 135.765 104.740 135.935 ;
        RECT 105.025 135.890 105.195 136.690 ;
        RECT 105.365 136.675 106.575 137.765 ;
        RECT 105.365 136.135 105.885 136.675 ;
        RECT 106.785 136.625 107.015 137.765 ;
        RECT 107.185 136.615 107.515 137.595 ;
        RECT 107.685 136.625 107.895 137.765 ;
        RECT 108.125 136.675 109.795 137.765 ;
        RECT 110.055 136.835 110.225 137.595 ;
        RECT 110.405 137.005 110.735 137.765 ;
        RECT 106.055 135.965 106.575 136.505 ;
        RECT 106.765 136.205 107.095 136.455 ;
        RECT 104.075 135.385 104.245 135.765 ;
        RECT 104.425 135.215 104.755 135.595 ;
        RECT 104.935 135.385 105.195 135.890 ;
        RECT 105.365 135.215 106.575 135.965 ;
        RECT 106.785 135.215 107.015 136.035 ;
        RECT 107.265 136.015 107.515 136.615 ;
        RECT 108.125 136.155 108.875 136.675 ;
        RECT 110.055 136.665 110.720 136.835 ;
        RECT 110.905 136.690 111.175 137.595 ;
        RECT 110.550 136.520 110.720 136.665 ;
        RECT 107.185 135.385 107.515 136.015 ;
        RECT 107.685 135.215 107.895 136.035 ;
        RECT 109.045 135.985 109.795 136.505 ;
        RECT 109.985 136.115 110.315 136.485 ;
        RECT 110.550 136.190 110.835 136.520 ;
        RECT 108.125 135.215 109.795 135.985 ;
        RECT 110.550 135.935 110.720 136.190 ;
        RECT 110.055 135.765 110.720 135.935 ;
        RECT 111.005 135.890 111.175 136.690 ;
        RECT 111.805 136.675 115.315 137.765 ;
        RECT 115.490 137.330 120.835 137.765 ;
        RECT 121.010 137.330 126.355 137.765 ;
        RECT 111.805 136.155 113.495 136.675 ;
        RECT 113.665 135.985 115.315 136.505 ;
        RECT 117.080 136.080 117.430 137.330 ;
        RECT 110.055 135.385 110.225 135.765 ;
        RECT 110.405 135.215 110.735 135.595 ;
        RECT 110.915 135.385 111.175 135.890 ;
        RECT 111.805 135.215 115.315 135.985 ;
        RECT 118.910 135.760 119.250 136.590 ;
        RECT 122.600 136.080 122.950 137.330 ;
        RECT 126.525 136.675 127.735 137.765 ;
        RECT 124.430 135.760 124.770 136.590 ;
        RECT 126.525 136.135 127.045 136.675 ;
        RECT 127.215 135.965 127.735 136.505 ;
        RECT 115.490 135.215 120.835 135.760 ;
        RECT 121.010 135.215 126.355 135.760 ;
        RECT 126.525 135.215 127.735 135.965 ;
        RECT 14.660 135.045 127.820 135.215 ;
        RECT 14.745 134.295 15.955 135.045 ;
        RECT 14.745 133.755 15.265 134.295 ;
        RECT 16.585 134.275 18.255 135.045 ;
        RECT 18.430 134.500 23.775 135.045 ;
        RECT 15.435 133.585 15.955 134.125 ;
        RECT 14.745 132.495 15.955 133.585 ;
        RECT 16.585 133.585 17.335 134.105 ;
        RECT 17.505 133.755 18.255 134.275 ;
        RECT 16.585 132.495 18.255 133.585 ;
        RECT 20.020 132.930 20.370 134.180 ;
        RECT 21.850 133.670 22.190 134.500 ;
        RECT 24.320 134.335 24.575 134.865 ;
        RECT 24.755 134.585 25.040 135.045 ;
        RECT 24.320 133.685 24.500 134.335 ;
        RECT 25.220 134.135 25.470 134.785 ;
        RECT 24.670 133.805 25.470 134.135 ;
        RECT 24.235 133.515 24.500 133.685 ;
        RECT 24.320 133.475 24.500 133.515 ;
        RECT 18.430 132.495 23.775 132.930 ;
        RECT 24.320 132.805 24.575 133.475 ;
        RECT 24.755 132.495 25.040 133.295 ;
        RECT 25.220 133.215 25.470 133.805 ;
        RECT 25.670 134.450 25.990 134.780 ;
        RECT 26.170 134.565 26.830 135.045 ;
        RECT 27.030 134.655 27.880 134.825 ;
        RECT 25.670 133.555 25.860 134.450 ;
        RECT 26.180 134.125 26.840 134.395 ;
        RECT 26.510 134.065 26.840 134.125 ;
        RECT 26.030 133.895 26.360 133.955 ;
        RECT 27.030 133.895 27.200 134.655 ;
        RECT 28.440 134.585 28.760 135.045 ;
        RECT 28.960 134.405 29.210 134.835 ;
        RECT 29.500 134.605 29.910 135.045 ;
        RECT 30.080 134.665 31.095 134.865 ;
        RECT 27.370 134.235 28.620 134.405 ;
        RECT 27.370 134.115 27.700 134.235 ;
        RECT 26.030 133.725 27.930 133.895 ;
        RECT 25.670 133.385 27.590 133.555 ;
        RECT 25.670 133.365 25.990 133.385 ;
        RECT 25.220 132.705 25.550 133.215 ;
        RECT 25.820 132.755 25.990 133.365 ;
        RECT 27.760 133.215 27.930 133.725 ;
        RECT 28.100 133.655 28.280 134.065 ;
        RECT 28.450 133.475 28.620 134.235 ;
        RECT 26.160 132.495 26.490 133.185 ;
        RECT 26.720 133.045 27.930 133.215 ;
        RECT 28.100 133.165 28.620 133.475 ;
        RECT 28.790 134.065 29.210 134.405 ;
        RECT 29.500 134.065 29.910 134.395 ;
        RECT 28.790 133.295 28.980 134.065 ;
        RECT 30.080 133.935 30.250 134.665 ;
        RECT 31.395 134.495 31.565 134.825 ;
        RECT 31.735 134.665 32.065 135.045 ;
        RECT 30.420 134.115 30.770 134.485 ;
        RECT 30.080 133.895 30.500 133.935 ;
        RECT 29.150 133.725 30.500 133.895 ;
        RECT 29.150 133.565 29.400 133.725 ;
        RECT 29.910 133.295 30.160 133.555 ;
        RECT 28.790 133.045 30.160 133.295 ;
        RECT 26.720 132.755 26.960 133.045 ;
        RECT 27.760 132.965 27.930 133.045 ;
        RECT 27.160 132.495 27.580 132.875 ;
        RECT 27.760 132.715 28.390 132.965 ;
        RECT 28.860 132.495 29.190 132.875 ;
        RECT 29.360 132.755 29.530 133.045 ;
        RECT 30.330 132.880 30.500 133.725 ;
        RECT 30.950 133.555 31.170 134.425 ;
        RECT 31.395 134.305 32.090 134.495 ;
        RECT 30.670 133.175 31.170 133.555 ;
        RECT 31.340 133.505 31.750 134.125 ;
        RECT 31.920 133.335 32.090 134.305 ;
        RECT 31.395 133.165 32.090 133.335 ;
        RECT 29.710 132.495 30.090 132.875 ;
        RECT 30.330 132.710 31.160 132.880 ;
        RECT 31.395 132.665 31.565 133.165 ;
        RECT 31.735 132.495 32.065 132.995 ;
        RECT 32.280 132.665 32.505 134.785 ;
        RECT 32.675 134.665 33.005 135.045 ;
        RECT 33.175 134.495 33.345 134.785 ;
        RECT 32.680 134.325 33.345 134.495 ;
        RECT 32.680 133.335 32.910 134.325 ;
        RECT 33.605 134.295 34.815 135.045 ;
        RECT 33.080 133.505 33.430 134.155 ;
        RECT 33.605 133.585 34.125 134.125 ;
        RECT 34.295 133.755 34.815 134.295 ;
        RECT 35.025 134.225 35.255 135.045 ;
        RECT 35.425 134.245 35.755 134.875 ;
        RECT 35.005 133.805 35.335 134.055 ;
        RECT 35.505 133.645 35.755 134.245 ;
        RECT 35.925 134.225 36.135 135.045 ;
        RECT 37.285 134.320 37.575 135.045 ;
        RECT 37.745 134.275 40.335 135.045 ;
        RECT 32.680 133.165 33.345 133.335 ;
        RECT 32.675 132.495 33.005 132.995 ;
        RECT 33.175 132.665 33.345 133.165 ;
        RECT 33.605 132.495 34.815 133.585 ;
        RECT 35.025 132.495 35.255 133.635 ;
        RECT 35.425 132.665 35.755 133.645 ;
        RECT 35.925 132.495 36.135 133.635 ;
        RECT 37.285 132.495 37.575 133.660 ;
        RECT 37.745 133.585 38.955 134.105 ;
        RECT 39.125 133.755 40.335 134.275 ;
        RECT 40.705 134.415 41.035 134.775 ;
        RECT 41.655 134.585 41.905 135.045 ;
        RECT 42.075 134.585 42.635 134.875 ;
        RECT 40.705 134.225 42.095 134.415 ;
        RECT 41.925 134.135 42.095 134.225 ;
        RECT 40.520 133.805 41.195 134.055 ;
        RECT 41.415 133.805 41.755 134.055 ;
        RECT 41.925 133.805 42.215 134.135 ;
        RECT 37.745 132.495 40.335 133.585 ;
        RECT 40.520 133.445 40.785 133.805 ;
        RECT 41.925 133.555 42.095 133.805 ;
        RECT 41.155 133.385 42.095 133.555 ;
        RECT 40.705 132.495 40.985 133.165 ;
        RECT 41.155 132.835 41.455 133.385 ;
        RECT 42.385 133.215 42.635 134.585 ;
        RECT 43.005 134.415 43.335 134.775 ;
        RECT 43.955 134.585 44.205 135.045 ;
        RECT 44.375 134.585 44.935 134.875 ;
        RECT 43.005 134.225 44.395 134.415 ;
        RECT 44.225 134.135 44.395 134.225 ;
        RECT 42.820 133.805 43.495 134.055 ;
        RECT 43.715 133.805 44.055 134.055 ;
        RECT 44.225 133.805 44.515 134.135 ;
        RECT 42.820 133.445 43.085 133.805 ;
        RECT 44.225 133.555 44.395 133.805 ;
        RECT 41.655 132.495 41.985 133.215 ;
        RECT 42.175 132.665 42.635 133.215 ;
        RECT 43.455 133.385 44.395 133.555 ;
        RECT 43.005 132.495 43.285 133.165 ;
        RECT 43.455 132.835 43.755 133.385 ;
        RECT 44.685 133.215 44.935 134.585 ;
        RECT 43.955 132.495 44.285 133.215 ;
        RECT 44.475 132.665 44.935 133.215 ;
        RECT 45.105 134.585 45.665 134.875 ;
        RECT 45.835 134.585 46.085 135.045 ;
        RECT 45.105 133.215 45.355 134.585 ;
        RECT 46.705 134.415 47.035 134.775 ;
        RECT 47.415 134.545 47.745 135.045 ;
        RECT 45.645 134.225 47.035 134.415 ;
        RECT 47.945 134.475 48.115 134.825 ;
        RECT 48.315 134.645 48.645 135.045 ;
        RECT 48.815 134.475 48.985 134.825 ;
        RECT 49.155 134.645 49.535 135.045 ;
        RECT 45.645 134.135 45.815 134.225 ;
        RECT 45.525 133.805 45.815 134.135 ;
        RECT 45.985 133.805 46.325 134.055 ;
        RECT 46.545 133.805 47.220 134.055 ;
        RECT 47.410 133.805 47.760 134.375 ;
        RECT 47.945 134.305 49.555 134.475 ;
        RECT 49.725 134.370 49.995 134.715 ;
        RECT 49.385 134.135 49.555 134.305 ;
        RECT 45.645 133.555 45.815 133.805 ;
        RECT 45.645 133.385 46.585 133.555 ;
        RECT 46.955 133.445 47.220 133.805 ;
        RECT 47.930 133.685 48.640 134.135 ;
        RECT 48.810 133.805 49.215 134.135 ;
        RECT 49.385 133.805 49.655 134.135 ;
        RECT 45.105 132.665 45.565 133.215 ;
        RECT 45.755 132.495 46.085 133.215 ;
        RECT 46.285 132.835 46.585 133.385 ;
        RECT 47.410 133.345 47.730 133.635 ;
        RECT 47.925 133.515 48.640 133.685 ;
        RECT 49.385 133.635 49.555 133.805 ;
        RECT 49.825 133.635 49.995 134.370 ;
        RECT 50.165 134.275 51.835 135.045 ;
        RECT 52.010 134.500 57.355 135.045 ;
        RECT 48.830 133.465 49.555 133.635 ;
        RECT 48.830 133.345 49.000 133.465 ;
        RECT 47.410 133.175 49.000 133.345 ;
        RECT 46.755 132.495 47.035 133.165 ;
        RECT 47.410 132.715 49.065 133.005 ;
        RECT 49.235 132.495 49.515 133.295 ;
        RECT 49.725 132.665 49.995 133.635 ;
        RECT 50.165 133.585 50.915 134.105 ;
        RECT 51.085 133.755 51.835 134.275 ;
        RECT 50.165 132.495 51.835 133.585 ;
        RECT 53.600 132.930 53.950 134.180 ;
        RECT 55.430 133.670 55.770 134.500 ;
        RECT 57.525 134.245 57.865 134.875 ;
        RECT 58.035 134.245 58.285 135.045 ;
        RECT 58.475 134.395 58.805 134.875 ;
        RECT 58.975 134.585 59.200 135.045 ;
        RECT 59.370 134.395 59.700 134.875 ;
        RECT 57.525 134.195 57.755 134.245 ;
        RECT 58.475 134.225 59.700 134.395 ;
        RECT 60.330 134.265 60.830 134.875 ;
        RECT 61.205 134.275 62.875 135.045 ;
        RECT 63.045 134.320 63.335 135.045 ;
        RECT 64.425 134.275 67.935 135.045 ;
        RECT 68.110 134.500 73.455 135.045 ;
        RECT 73.630 134.500 78.975 135.045 ;
        RECT 57.525 133.635 57.700 134.195 ;
        RECT 57.870 133.885 58.565 134.055 ;
        RECT 58.395 133.635 58.565 133.885 ;
        RECT 58.740 133.855 59.160 134.055 ;
        RECT 59.330 133.855 59.660 134.055 ;
        RECT 59.830 133.855 60.160 134.055 ;
        RECT 60.330 133.635 60.500 134.265 ;
        RECT 60.685 133.805 61.035 134.055 ;
        RECT 52.010 132.495 57.355 132.930 ;
        RECT 57.525 132.665 57.865 133.635 ;
        RECT 58.035 132.495 58.205 133.635 ;
        RECT 58.395 133.465 60.830 133.635 ;
        RECT 58.475 132.495 58.725 133.295 ;
        RECT 59.370 132.665 59.700 133.465 ;
        RECT 60.000 132.495 60.330 133.295 ;
        RECT 60.500 132.665 60.830 133.465 ;
        RECT 61.205 133.585 61.955 134.105 ;
        RECT 62.125 133.755 62.875 134.275 ;
        RECT 61.205 132.495 62.875 133.585 ;
        RECT 63.045 132.495 63.335 133.660 ;
        RECT 64.425 133.585 66.115 134.105 ;
        RECT 66.285 133.755 67.935 134.275 ;
        RECT 64.425 132.495 67.935 133.585 ;
        RECT 69.700 132.930 70.050 134.180 ;
        RECT 71.530 133.670 71.870 134.500 ;
        RECT 75.220 132.930 75.570 134.180 ;
        RECT 77.050 133.670 77.390 134.500 ;
        RECT 79.350 134.265 79.850 134.875 ;
        RECT 79.145 133.805 79.495 134.055 ;
        RECT 79.680 133.635 79.850 134.265 ;
        RECT 80.480 134.395 80.810 134.875 ;
        RECT 80.980 134.585 81.205 135.045 ;
        RECT 81.375 134.395 81.705 134.875 ;
        RECT 80.480 134.225 81.705 134.395 ;
        RECT 81.895 134.245 82.145 135.045 ;
        RECT 82.315 134.245 82.655 134.875 ;
        RECT 80.020 133.855 80.350 134.055 ;
        RECT 80.520 133.855 80.850 134.055 ;
        RECT 81.020 133.855 81.440 134.055 ;
        RECT 81.615 133.885 82.310 134.055 ;
        RECT 81.615 133.635 81.785 133.885 ;
        RECT 82.480 133.635 82.655 134.245 ;
        RECT 79.350 133.465 81.785 133.635 ;
        RECT 68.110 132.495 73.455 132.930 ;
        RECT 73.630 132.495 78.975 132.930 ;
        RECT 79.350 132.665 79.680 133.465 ;
        RECT 79.850 132.495 80.180 133.295 ;
        RECT 80.480 132.665 80.810 133.465 ;
        RECT 81.455 132.495 81.705 133.295 ;
        RECT 81.975 132.495 82.145 133.635 ;
        RECT 82.315 132.665 82.655 133.635 ;
        RECT 82.825 134.245 83.165 134.875 ;
        RECT 83.335 134.245 83.585 135.045 ;
        RECT 83.775 134.395 84.105 134.875 ;
        RECT 84.275 134.585 84.500 135.045 ;
        RECT 84.670 134.395 85.000 134.875 ;
        RECT 82.825 133.635 83.000 134.245 ;
        RECT 83.775 134.225 85.000 134.395 ;
        RECT 85.630 134.265 86.130 134.875 ;
        RECT 86.965 134.275 88.635 135.045 ;
        RECT 88.805 134.320 89.095 135.045 ;
        RECT 83.170 133.885 83.865 134.055 ;
        RECT 83.695 133.635 83.865 133.885 ;
        RECT 84.040 133.855 84.460 134.055 ;
        RECT 84.630 133.855 84.960 134.055 ;
        RECT 85.130 133.855 85.460 134.055 ;
        RECT 85.630 133.635 85.800 134.265 ;
        RECT 85.985 133.805 86.335 134.055 ;
        RECT 82.825 132.665 83.165 133.635 ;
        RECT 83.335 132.495 83.505 133.635 ;
        RECT 83.695 133.465 86.130 133.635 ;
        RECT 83.775 132.495 84.025 133.295 ;
        RECT 84.670 132.665 85.000 133.465 ;
        RECT 85.300 132.495 85.630 133.295 ;
        RECT 85.800 132.665 86.130 133.465 ;
        RECT 86.965 133.585 87.715 134.105 ;
        RECT 87.885 133.755 88.635 134.275 ;
        RECT 89.540 134.235 89.785 134.840 ;
        RECT 90.005 134.510 90.515 135.045 ;
        RECT 89.265 134.065 90.495 134.235 ;
        RECT 86.965 132.495 88.635 133.585 ;
        RECT 88.805 132.495 89.095 133.660 ;
        RECT 89.265 133.255 89.605 134.065 ;
        RECT 89.775 133.500 90.525 133.690 ;
        RECT 89.265 132.845 89.780 133.255 ;
        RECT 90.015 132.495 90.185 133.255 ;
        RECT 90.355 132.835 90.525 133.500 ;
        RECT 90.695 133.515 90.885 134.875 ;
        RECT 91.055 134.365 91.330 134.875 ;
        RECT 91.520 134.510 92.050 134.875 ;
        RECT 92.475 134.645 92.805 135.045 ;
        RECT 91.875 134.475 92.050 134.510 ;
        RECT 91.055 134.195 91.335 134.365 ;
        RECT 91.055 133.715 91.330 134.195 ;
        RECT 91.535 133.515 91.705 134.315 ;
        RECT 90.695 133.345 91.705 133.515 ;
        RECT 91.875 134.305 92.805 134.475 ;
        RECT 92.975 134.305 93.230 134.875 ;
        RECT 93.495 134.495 93.665 134.875 ;
        RECT 93.845 134.665 94.175 135.045 ;
        RECT 93.495 134.325 94.160 134.495 ;
        RECT 94.355 134.370 94.615 134.875 ;
        RECT 91.875 133.175 92.045 134.305 ;
        RECT 92.635 134.135 92.805 134.305 ;
        RECT 90.920 133.005 92.045 133.175 ;
        RECT 92.215 133.805 92.410 134.135 ;
        RECT 92.635 133.805 92.890 134.135 ;
        RECT 92.215 132.835 92.385 133.805 ;
        RECT 93.060 133.635 93.230 134.305 ;
        RECT 93.425 133.775 93.755 134.145 ;
        RECT 93.990 134.070 94.160 134.325 ;
        RECT 90.355 132.665 92.385 132.835 ;
        RECT 92.555 132.495 92.725 133.635 ;
        RECT 92.895 132.665 93.230 133.635 ;
        RECT 93.990 133.740 94.275 134.070 ;
        RECT 93.990 133.595 94.160 133.740 ;
        RECT 93.495 133.425 94.160 133.595 ;
        RECT 94.445 133.570 94.615 134.370 ;
        RECT 95.245 134.275 96.915 135.045 ;
        RECT 97.460 134.365 97.715 134.865 ;
        RECT 97.895 134.585 98.180 135.045 ;
        RECT 93.495 132.665 93.665 133.425 ;
        RECT 93.845 132.495 94.175 133.255 ;
        RECT 94.345 132.665 94.615 133.570 ;
        RECT 95.245 133.585 95.995 134.105 ;
        RECT 96.165 133.755 96.915 134.275 ;
        RECT 97.375 134.335 97.715 134.365 ;
        RECT 97.375 134.195 97.640 134.335 ;
        RECT 95.245 132.495 96.915 133.585 ;
        RECT 97.460 133.475 97.640 134.195 ;
        RECT 98.360 134.135 98.610 134.785 ;
        RECT 97.810 133.805 98.610 134.135 ;
        RECT 97.460 132.805 97.715 133.475 ;
        RECT 97.895 132.495 98.180 133.295 ;
        RECT 98.360 133.215 98.610 133.805 ;
        RECT 98.810 134.450 99.130 134.780 ;
        RECT 99.310 134.565 99.970 135.045 ;
        RECT 100.170 134.655 101.020 134.825 ;
        RECT 98.810 133.555 99.000 134.450 ;
        RECT 99.320 134.125 99.980 134.395 ;
        RECT 99.650 134.065 99.980 134.125 ;
        RECT 99.170 133.895 99.500 133.955 ;
        RECT 100.170 133.895 100.340 134.655 ;
        RECT 101.580 134.585 101.900 135.045 ;
        RECT 102.100 134.405 102.350 134.835 ;
        RECT 102.640 134.605 103.050 135.045 ;
        RECT 103.220 134.665 104.235 134.865 ;
        RECT 100.510 134.235 101.760 134.405 ;
        RECT 100.510 134.115 100.840 134.235 ;
        RECT 99.170 133.725 101.070 133.895 ;
        RECT 98.810 133.385 100.730 133.555 ;
        RECT 98.810 133.365 99.130 133.385 ;
        RECT 98.360 132.705 98.690 133.215 ;
        RECT 98.960 132.755 99.130 133.365 ;
        RECT 100.900 133.215 101.070 133.725 ;
        RECT 101.240 133.655 101.420 134.065 ;
        RECT 101.590 133.475 101.760 134.235 ;
        RECT 99.300 132.495 99.630 133.185 ;
        RECT 99.860 133.045 101.070 133.215 ;
        RECT 101.240 133.165 101.760 133.475 ;
        RECT 101.930 134.065 102.350 134.405 ;
        RECT 102.640 134.065 103.050 134.395 ;
        RECT 101.930 133.295 102.120 134.065 ;
        RECT 103.220 133.935 103.390 134.665 ;
        RECT 104.535 134.495 104.705 134.825 ;
        RECT 104.875 134.665 105.205 135.045 ;
        RECT 103.560 134.115 103.910 134.485 ;
        RECT 103.220 133.895 103.640 133.935 ;
        RECT 102.290 133.725 103.640 133.895 ;
        RECT 102.290 133.565 102.540 133.725 ;
        RECT 103.050 133.295 103.300 133.555 ;
        RECT 101.930 133.045 103.300 133.295 ;
        RECT 99.860 132.755 100.100 133.045 ;
        RECT 100.900 132.965 101.070 133.045 ;
        RECT 100.300 132.495 100.720 132.875 ;
        RECT 100.900 132.715 101.530 132.965 ;
        RECT 102.000 132.495 102.330 132.875 ;
        RECT 102.500 132.755 102.670 133.045 ;
        RECT 103.470 132.880 103.640 133.725 ;
        RECT 104.090 133.555 104.310 134.425 ;
        RECT 104.535 134.305 105.230 134.495 ;
        RECT 103.810 133.175 104.310 133.555 ;
        RECT 104.480 133.505 104.890 134.125 ;
        RECT 105.060 133.335 105.230 134.305 ;
        RECT 104.535 133.165 105.230 133.335 ;
        RECT 102.850 132.495 103.230 132.875 ;
        RECT 103.470 132.710 104.300 132.880 ;
        RECT 104.535 132.665 104.705 133.165 ;
        RECT 104.875 132.495 105.205 132.995 ;
        RECT 105.420 132.665 105.645 134.785 ;
        RECT 105.815 134.665 106.145 135.045 ;
        RECT 106.315 134.495 106.485 134.785 ;
        RECT 105.820 134.325 106.485 134.495 ;
        RECT 105.820 133.335 106.050 134.325 ;
        RECT 106.745 134.275 109.335 135.045 ;
        RECT 106.220 133.505 106.570 134.155 ;
        RECT 106.745 133.585 107.955 134.105 ;
        RECT 108.125 133.755 109.335 134.275 ;
        RECT 109.505 134.585 110.065 134.875 ;
        RECT 110.235 134.585 110.485 135.045 ;
        RECT 105.820 133.165 106.485 133.335 ;
        RECT 105.815 132.495 106.145 132.995 ;
        RECT 106.315 132.665 106.485 133.165 ;
        RECT 106.745 132.495 109.335 133.585 ;
        RECT 109.505 133.215 109.755 134.585 ;
        RECT 111.105 134.415 111.435 134.775 ;
        RECT 110.045 134.225 111.435 134.415 ;
        RECT 111.805 134.585 112.365 134.875 ;
        RECT 112.535 134.585 112.785 135.045 ;
        RECT 110.045 134.135 110.215 134.225 ;
        RECT 109.925 133.805 110.215 134.135 ;
        RECT 110.385 133.805 110.725 134.055 ;
        RECT 110.945 133.805 111.620 134.055 ;
        RECT 110.045 133.555 110.215 133.805 ;
        RECT 110.045 133.385 110.985 133.555 ;
        RECT 111.355 133.445 111.620 133.805 ;
        RECT 109.505 132.665 109.965 133.215 ;
        RECT 110.155 132.495 110.485 133.215 ;
        RECT 110.685 132.835 110.985 133.385 ;
        RECT 111.805 133.215 112.055 134.585 ;
        RECT 113.405 134.415 113.735 134.775 ;
        RECT 112.345 134.225 113.735 134.415 ;
        RECT 114.565 134.320 114.855 135.045 ;
        RECT 115.490 134.500 120.835 135.045 ;
        RECT 121.010 134.500 126.355 135.045 ;
        RECT 112.345 134.135 112.515 134.225 ;
        RECT 112.225 133.805 112.515 134.135 ;
        RECT 112.685 133.805 113.025 134.055 ;
        RECT 113.245 133.805 113.920 134.055 ;
        RECT 112.345 133.555 112.515 133.805 ;
        RECT 112.345 133.385 113.285 133.555 ;
        RECT 113.655 133.445 113.920 133.805 ;
        RECT 111.155 132.495 111.435 133.165 ;
        RECT 111.805 132.665 112.265 133.215 ;
        RECT 112.455 132.495 112.785 133.215 ;
        RECT 112.985 132.835 113.285 133.385 ;
        RECT 113.455 132.495 113.735 133.165 ;
        RECT 114.565 132.495 114.855 133.660 ;
        RECT 117.080 132.930 117.430 134.180 ;
        RECT 118.910 133.670 119.250 134.500 ;
        RECT 122.600 132.930 122.950 134.180 ;
        RECT 124.430 133.670 124.770 134.500 ;
        RECT 126.525 134.295 127.735 135.045 ;
        RECT 126.525 133.585 127.045 134.125 ;
        RECT 127.215 133.755 127.735 134.295 ;
        RECT 115.490 132.495 120.835 132.930 ;
        RECT 121.010 132.495 126.355 132.930 ;
        RECT 126.525 132.495 127.735 133.585 ;
        RECT 14.660 132.325 127.820 132.495 ;
        RECT 14.745 131.235 15.955 132.325 ;
        RECT 14.745 130.525 15.265 131.065 ;
        RECT 15.435 130.695 15.955 131.235 ;
        RECT 16.125 131.235 18.715 132.325 ;
        RECT 16.125 130.715 17.335 131.235 ;
        RECT 18.945 131.185 19.155 132.325 ;
        RECT 19.325 131.175 19.655 132.155 ;
        RECT 19.825 131.185 20.055 132.325 ;
        RECT 20.265 131.565 20.780 131.975 ;
        RECT 21.015 131.565 21.185 132.325 ;
        RECT 21.355 131.985 23.385 132.155 ;
        RECT 17.505 130.545 18.715 131.065 ;
        RECT 14.745 129.775 15.955 130.525 ;
        RECT 16.125 129.775 18.715 130.545 ;
        RECT 18.945 129.775 19.155 130.595 ;
        RECT 19.325 130.575 19.575 131.175 ;
        RECT 19.745 130.765 20.075 131.015 ;
        RECT 20.265 130.755 20.605 131.565 ;
        RECT 21.355 131.320 21.525 131.985 ;
        RECT 21.920 131.645 23.045 131.815 ;
        RECT 20.775 131.130 21.525 131.320 ;
        RECT 21.695 131.305 22.705 131.475 ;
        RECT 19.325 129.945 19.655 130.575 ;
        RECT 19.825 129.775 20.055 130.595 ;
        RECT 20.265 130.585 21.495 130.755 ;
        RECT 20.540 129.980 20.785 130.585 ;
        RECT 21.005 129.775 21.515 130.310 ;
        RECT 21.695 129.945 21.885 131.305 ;
        RECT 22.055 130.285 22.330 131.105 ;
        RECT 22.535 130.505 22.705 131.305 ;
        RECT 22.875 130.515 23.045 131.645 ;
        RECT 23.215 131.015 23.385 131.985 ;
        RECT 23.555 131.185 23.725 132.325 ;
        RECT 23.895 131.185 24.230 132.155 ;
        RECT 23.215 130.685 23.410 131.015 ;
        RECT 23.635 130.685 23.890 131.015 ;
        RECT 23.635 130.515 23.805 130.685 ;
        RECT 24.060 130.515 24.230 131.185 ;
        RECT 24.405 131.160 24.695 132.325 ;
        RECT 24.865 131.250 25.135 132.155 ;
        RECT 25.305 131.565 25.635 132.325 ;
        RECT 25.815 131.395 25.985 132.155 ;
        RECT 22.875 130.345 23.805 130.515 ;
        RECT 22.875 130.310 23.050 130.345 ;
        RECT 22.055 130.115 22.335 130.285 ;
        RECT 22.055 129.945 22.330 130.115 ;
        RECT 22.520 129.945 23.050 130.310 ;
        RECT 23.475 129.775 23.805 130.175 ;
        RECT 23.975 129.945 24.230 130.515 ;
        RECT 24.405 129.775 24.695 130.500 ;
        RECT 24.865 130.450 25.035 131.250 ;
        RECT 25.320 131.225 25.985 131.395 ;
        RECT 25.320 131.080 25.490 131.225 ;
        RECT 26.285 131.185 26.515 132.325 ;
        RECT 26.685 131.175 27.015 132.155 ;
        RECT 27.185 131.185 27.395 132.325 ;
        RECT 27.625 131.565 28.140 131.975 ;
        RECT 28.375 131.565 28.545 132.325 ;
        RECT 28.715 131.985 30.745 132.155 ;
        RECT 25.205 130.750 25.490 131.080 ;
        RECT 25.320 130.495 25.490 130.750 ;
        RECT 25.725 130.675 26.055 131.045 ;
        RECT 26.265 130.765 26.595 131.015 ;
        RECT 24.865 129.945 25.125 130.450 ;
        RECT 25.320 130.325 25.985 130.495 ;
        RECT 25.305 129.775 25.635 130.155 ;
        RECT 25.815 129.945 25.985 130.325 ;
        RECT 26.285 129.775 26.515 130.595 ;
        RECT 26.765 130.575 27.015 131.175 ;
        RECT 27.625 130.755 27.965 131.565 ;
        RECT 28.715 131.320 28.885 131.985 ;
        RECT 29.280 131.645 30.405 131.815 ;
        RECT 28.135 131.130 28.885 131.320 ;
        RECT 29.055 131.305 30.065 131.475 ;
        RECT 26.685 129.945 27.015 130.575 ;
        RECT 27.185 129.775 27.395 130.595 ;
        RECT 27.625 130.585 28.855 130.755 ;
        RECT 27.900 129.980 28.145 130.585 ;
        RECT 28.365 129.775 28.875 130.310 ;
        RECT 29.055 129.945 29.245 131.305 ;
        RECT 29.415 130.965 29.690 131.105 ;
        RECT 29.415 130.795 29.695 130.965 ;
        RECT 29.415 129.945 29.690 130.795 ;
        RECT 29.895 130.505 30.065 131.305 ;
        RECT 30.235 130.515 30.405 131.645 ;
        RECT 30.575 131.015 30.745 131.985 ;
        RECT 30.915 131.185 31.085 132.325 ;
        RECT 31.255 131.185 31.590 132.155 ;
        RECT 32.140 131.345 32.395 132.015 ;
        RECT 32.575 131.525 32.860 132.325 ;
        RECT 33.040 131.605 33.370 132.115 ;
        RECT 32.140 131.305 32.320 131.345 ;
        RECT 30.575 130.685 30.770 131.015 ;
        RECT 30.995 130.685 31.250 131.015 ;
        RECT 30.995 130.515 31.165 130.685 ;
        RECT 31.420 130.515 31.590 131.185 ;
        RECT 32.055 131.135 32.320 131.305 ;
        RECT 30.235 130.345 31.165 130.515 ;
        RECT 30.235 130.310 30.410 130.345 ;
        RECT 29.880 129.945 30.410 130.310 ;
        RECT 30.835 129.775 31.165 130.175 ;
        RECT 31.335 129.945 31.590 130.515 ;
        RECT 32.140 130.485 32.320 131.135 ;
        RECT 33.040 131.015 33.290 131.605 ;
        RECT 33.640 131.455 33.810 132.065 ;
        RECT 33.980 131.635 34.310 132.325 ;
        RECT 34.540 131.775 34.780 132.065 ;
        RECT 34.980 131.945 35.400 132.325 ;
        RECT 35.580 131.855 36.210 132.105 ;
        RECT 36.680 131.945 37.010 132.325 ;
        RECT 35.580 131.775 35.750 131.855 ;
        RECT 37.180 131.775 37.350 132.065 ;
        RECT 37.530 131.945 37.910 132.325 ;
        RECT 38.150 131.940 38.980 132.110 ;
        RECT 34.540 131.605 35.750 131.775 ;
        RECT 32.490 130.685 33.290 131.015 ;
        RECT 32.140 129.955 32.395 130.485 ;
        RECT 32.575 129.775 32.860 130.235 ;
        RECT 33.040 130.035 33.290 130.685 ;
        RECT 33.490 131.435 33.810 131.455 ;
        RECT 33.490 131.265 35.410 131.435 ;
        RECT 33.490 130.370 33.680 131.265 ;
        RECT 35.580 131.095 35.750 131.605 ;
        RECT 35.920 131.345 36.440 131.655 ;
        RECT 33.850 130.925 35.750 131.095 ;
        RECT 33.850 130.865 34.180 130.925 ;
        RECT 34.330 130.695 34.660 130.755 ;
        RECT 34.000 130.425 34.660 130.695 ;
        RECT 33.490 130.040 33.810 130.370 ;
        RECT 33.990 129.775 34.650 130.255 ;
        RECT 34.850 130.165 35.020 130.925 ;
        RECT 35.920 130.755 36.100 131.165 ;
        RECT 35.190 130.585 35.520 130.705 ;
        RECT 36.270 130.585 36.440 131.345 ;
        RECT 35.190 130.415 36.440 130.585 ;
        RECT 36.610 131.525 37.980 131.775 ;
        RECT 36.610 130.755 36.800 131.525 ;
        RECT 37.730 131.265 37.980 131.525 ;
        RECT 36.970 131.095 37.220 131.255 ;
        RECT 38.150 131.095 38.320 131.940 ;
        RECT 39.215 131.655 39.385 132.155 ;
        RECT 39.555 131.825 39.885 132.325 ;
        RECT 38.490 131.265 38.990 131.645 ;
        RECT 39.215 131.485 39.910 131.655 ;
        RECT 36.970 130.925 38.320 131.095 ;
        RECT 37.900 130.885 38.320 130.925 ;
        RECT 36.610 130.415 37.030 130.755 ;
        RECT 37.320 130.425 37.730 130.755 ;
        RECT 34.850 129.995 35.700 130.165 ;
        RECT 36.260 129.775 36.580 130.235 ;
        RECT 36.780 129.985 37.030 130.415 ;
        RECT 37.320 129.775 37.730 130.215 ;
        RECT 37.900 130.155 38.070 130.885 ;
        RECT 38.240 130.335 38.590 130.705 ;
        RECT 38.770 130.395 38.990 131.265 ;
        RECT 39.160 130.695 39.570 131.315 ;
        RECT 39.740 130.515 39.910 131.485 ;
        RECT 39.215 130.325 39.910 130.515 ;
        RECT 37.900 129.955 38.915 130.155 ;
        RECT 39.215 129.995 39.385 130.325 ;
        RECT 39.555 129.775 39.885 130.155 ;
        RECT 40.100 130.035 40.325 132.155 ;
        RECT 40.495 131.825 40.825 132.325 ;
        RECT 40.995 131.655 41.165 132.155 ;
        RECT 40.500 131.485 41.165 131.655 ;
        RECT 40.500 130.495 40.730 131.485 ;
        RECT 40.900 130.665 41.250 131.315 ;
        RECT 42.350 131.185 42.685 132.155 ;
        RECT 42.855 131.185 43.025 132.325 ;
        RECT 43.195 131.985 45.225 132.155 ;
        RECT 42.350 130.515 42.520 131.185 ;
        RECT 43.195 131.015 43.365 131.985 ;
        RECT 42.690 130.685 42.945 131.015 ;
        RECT 43.170 130.685 43.365 131.015 ;
        RECT 43.535 131.645 44.660 131.815 ;
        RECT 42.775 130.515 42.945 130.685 ;
        RECT 43.535 130.515 43.705 131.645 ;
        RECT 40.500 130.325 41.165 130.495 ;
        RECT 40.495 129.775 40.825 130.155 ;
        RECT 40.995 130.035 41.165 130.325 ;
        RECT 42.350 129.945 42.605 130.515 ;
        RECT 42.775 130.345 43.705 130.515 ;
        RECT 43.875 131.305 44.885 131.475 ;
        RECT 43.875 130.505 44.045 131.305 ;
        RECT 44.250 130.625 44.525 131.105 ;
        RECT 44.245 130.455 44.525 130.625 ;
        RECT 43.530 130.310 43.705 130.345 ;
        RECT 42.775 129.775 43.105 130.175 ;
        RECT 43.530 129.945 44.060 130.310 ;
        RECT 44.250 129.945 44.525 130.455 ;
        RECT 44.695 129.945 44.885 131.305 ;
        RECT 45.055 131.320 45.225 131.985 ;
        RECT 45.395 131.565 45.565 132.325 ;
        RECT 45.800 131.565 46.315 131.975 ;
        RECT 45.055 131.130 45.805 131.320 ;
        RECT 45.975 130.755 46.315 131.565 ;
        RECT 45.085 130.585 46.315 130.755 ;
        RECT 46.945 131.185 47.215 132.155 ;
        RECT 47.425 131.525 47.705 132.325 ;
        RECT 47.875 131.815 49.530 132.105 ;
        RECT 47.940 131.475 49.530 131.645 ;
        RECT 47.940 131.355 48.110 131.475 ;
        RECT 47.385 131.185 48.110 131.355 ;
        RECT 45.065 129.775 45.575 130.310 ;
        RECT 45.795 129.980 46.040 130.585 ;
        RECT 46.945 130.450 47.115 131.185 ;
        RECT 47.385 131.015 47.555 131.185 ;
        RECT 48.300 131.135 49.015 131.305 ;
        RECT 49.210 131.185 49.530 131.475 ;
        RECT 50.165 131.160 50.455 132.325 ;
        RECT 50.625 131.605 51.085 132.155 ;
        RECT 51.275 131.605 51.605 132.325 ;
        RECT 47.285 130.685 47.555 131.015 ;
        RECT 47.725 130.685 48.130 131.015 ;
        RECT 48.300 130.685 49.010 131.135 ;
        RECT 47.385 130.515 47.555 130.685 ;
        RECT 46.945 130.105 47.215 130.450 ;
        RECT 47.385 130.345 48.995 130.515 ;
        RECT 49.180 130.445 49.530 131.015 ;
        RECT 47.405 129.775 47.785 130.175 ;
        RECT 47.955 129.995 48.125 130.345 ;
        RECT 48.295 129.775 48.625 130.175 ;
        RECT 48.825 129.995 48.995 130.345 ;
        RECT 49.195 129.775 49.525 130.275 ;
        RECT 50.165 129.775 50.455 130.500 ;
        RECT 50.625 130.235 50.875 131.605 ;
        RECT 51.805 131.435 52.105 131.985 ;
        RECT 52.275 131.655 52.555 132.325 ;
        RECT 51.165 131.265 52.105 131.435 ;
        RECT 51.165 131.015 51.335 131.265 ;
        RECT 52.475 131.015 52.740 131.375 ;
        RECT 51.045 130.685 51.335 131.015 ;
        RECT 51.505 130.765 51.845 131.015 ;
        RECT 52.065 130.765 52.740 131.015 ;
        RECT 53.845 131.185 54.185 132.155 ;
        RECT 54.355 131.185 54.525 132.325 ;
        RECT 54.795 131.525 55.045 132.325 ;
        RECT 55.690 131.355 56.020 132.155 ;
        RECT 56.320 131.525 56.650 132.325 ;
        RECT 56.820 131.355 57.150 132.155 ;
        RECT 54.715 131.185 57.150 131.355 ;
        RECT 57.525 131.185 57.865 132.155 ;
        RECT 58.035 131.185 58.205 132.325 ;
        RECT 58.475 131.525 58.725 132.325 ;
        RECT 59.370 131.355 59.700 132.155 ;
        RECT 60.000 131.525 60.330 132.325 ;
        RECT 60.500 131.355 60.830 132.155 ;
        RECT 58.395 131.185 60.830 131.355 ;
        RECT 61.665 131.235 65.175 132.325 ;
        RECT 65.345 131.565 65.860 131.975 ;
        RECT 66.095 131.565 66.265 132.325 ;
        RECT 66.435 131.985 68.465 132.155 ;
        RECT 51.165 130.595 51.335 130.685 ;
        RECT 51.165 130.405 52.555 130.595 ;
        RECT 50.625 129.945 51.185 130.235 ;
        RECT 51.355 129.775 51.605 130.235 ;
        RECT 52.225 130.045 52.555 130.405 ;
        RECT 53.845 130.575 54.020 131.185 ;
        RECT 54.715 130.935 54.885 131.185 ;
        RECT 54.190 130.765 54.885 130.935 ;
        RECT 55.060 130.765 55.480 130.965 ;
        RECT 55.650 130.765 55.980 130.965 ;
        RECT 56.150 130.765 56.480 130.965 ;
        RECT 53.845 129.945 54.185 130.575 ;
        RECT 54.355 129.775 54.605 130.575 ;
        RECT 54.795 130.425 56.020 130.595 ;
        RECT 54.795 129.945 55.125 130.425 ;
        RECT 55.295 129.775 55.520 130.235 ;
        RECT 55.690 129.945 56.020 130.425 ;
        RECT 56.650 130.555 56.820 131.185 ;
        RECT 57.005 130.765 57.355 131.015 ;
        RECT 57.525 130.625 57.700 131.185 ;
        RECT 58.395 130.935 58.565 131.185 ;
        RECT 57.870 130.765 58.565 130.935 ;
        RECT 58.740 130.765 59.160 130.965 ;
        RECT 59.330 130.765 59.660 130.965 ;
        RECT 59.830 130.765 60.160 130.965 ;
        RECT 57.525 130.575 57.755 130.625 ;
        RECT 56.650 129.945 57.150 130.555 ;
        RECT 57.525 129.945 57.865 130.575 ;
        RECT 58.035 129.775 58.285 130.575 ;
        RECT 58.475 130.425 59.700 130.595 ;
        RECT 58.475 129.945 58.805 130.425 ;
        RECT 58.975 129.775 59.200 130.235 ;
        RECT 59.370 129.945 59.700 130.425 ;
        RECT 60.330 130.555 60.500 131.185 ;
        RECT 60.685 130.765 61.035 131.015 ;
        RECT 61.665 130.715 63.355 131.235 ;
        RECT 60.330 129.945 60.830 130.555 ;
        RECT 63.525 130.545 65.175 131.065 ;
        RECT 65.345 130.755 65.685 131.565 ;
        RECT 66.435 131.320 66.605 131.985 ;
        RECT 67.000 131.645 68.125 131.815 ;
        RECT 65.855 131.130 66.605 131.320 ;
        RECT 66.775 131.305 67.785 131.475 ;
        RECT 65.345 130.585 66.575 130.755 ;
        RECT 61.665 129.775 65.175 130.545 ;
        RECT 65.620 129.980 65.865 130.585 ;
        RECT 66.085 129.775 66.595 130.310 ;
        RECT 66.775 129.945 66.965 131.305 ;
        RECT 67.135 130.965 67.410 131.105 ;
        RECT 67.135 130.795 67.415 130.965 ;
        RECT 67.135 129.945 67.410 130.795 ;
        RECT 67.615 130.505 67.785 131.305 ;
        RECT 67.955 130.515 68.125 131.645 ;
        RECT 68.295 131.015 68.465 131.985 ;
        RECT 68.635 131.185 68.805 132.325 ;
        RECT 68.975 131.185 69.310 132.155 ;
        RECT 69.575 131.395 69.745 132.155 ;
        RECT 69.925 131.565 70.255 132.325 ;
        RECT 69.575 131.225 70.240 131.395 ;
        RECT 70.425 131.250 70.695 132.155 ;
        RECT 70.870 131.900 71.205 132.325 ;
        RECT 71.375 131.720 71.560 132.125 ;
        RECT 68.295 130.685 68.490 131.015 ;
        RECT 68.715 130.685 68.970 131.015 ;
        RECT 68.715 130.515 68.885 130.685 ;
        RECT 69.140 130.515 69.310 131.185 ;
        RECT 70.070 131.080 70.240 131.225 ;
        RECT 69.505 130.675 69.835 131.045 ;
        RECT 70.070 130.750 70.355 131.080 ;
        RECT 67.955 130.345 68.885 130.515 ;
        RECT 67.955 130.310 68.130 130.345 ;
        RECT 67.600 129.945 68.130 130.310 ;
        RECT 68.555 129.775 68.885 130.175 ;
        RECT 69.055 129.945 69.310 130.515 ;
        RECT 70.070 130.495 70.240 130.750 ;
        RECT 69.575 130.325 70.240 130.495 ;
        RECT 70.525 130.450 70.695 131.250 ;
        RECT 69.575 129.945 69.745 130.325 ;
        RECT 69.925 129.775 70.255 130.155 ;
        RECT 70.435 129.945 70.695 130.450 ;
        RECT 70.895 131.545 71.560 131.720 ;
        RECT 71.765 131.545 72.095 132.325 ;
        RECT 70.895 130.515 71.235 131.545 ;
        RECT 72.265 131.355 72.535 132.125 ;
        RECT 72.710 131.900 73.045 132.325 ;
        RECT 73.215 131.720 73.400 132.125 ;
        RECT 71.405 131.185 72.535 131.355 ;
        RECT 71.405 130.685 71.655 131.185 ;
        RECT 70.895 130.345 71.580 130.515 ;
        RECT 71.835 130.435 72.195 131.015 ;
        RECT 70.870 129.775 71.205 130.175 ;
        RECT 71.375 129.945 71.580 130.345 ;
        RECT 72.365 130.275 72.535 131.185 ;
        RECT 72.735 131.545 73.400 131.720 ;
        RECT 73.605 131.545 73.935 132.325 ;
        RECT 72.735 130.515 73.075 131.545 ;
        RECT 74.105 131.355 74.375 132.125 ;
        RECT 73.245 131.185 74.375 131.355 ;
        RECT 73.245 130.685 73.495 131.185 ;
        RECT 72.735 130.345 73.420 130.515 ;
        RECT 73.675 130.435 74.035 131.015 ;
        RECT 71.790 129.775 72.065 130.255 ;
        RECT 72.275 129.945 72.535 130.275 ;
        RECT 72.710 129.775 73.045 130.175 ;
        RECT 73.215 129.945 73.420 130.345 ;
        RECT 74.205 130.275 74.375 131.185 ;
        RECT 74.545 131.235 75.755 132.325 ;
        RECT 74.545 130.695 75.065 131.235 ;
        RECT 75.925 131.160 76.215 132.325 ;
        RECT 76.385 131.235 79.895 132.325 ;
        RECT 75.235 130.525 75.755 131.065 ;
        RECT 76.385 130.715 78.075 131.235 ;
        RECT 80.065 131.185 80.335 132.155 ;
        RECT 80.545 131.525 80.825 132.325 ;
        RECT 80.995 131.815 82.650 132.105 ;
        RECT 81.060 131.475 82.650 131.645 ;
        RECT 81.060 131.355 81.230 131.475 ;
        RECT 80.505 131.185 81.230 131.355 ;
        RECT 78.245 130.545 79.895 131.065 ;
        RECT 73.630 129.775 73.905 130.255 ;
        RECT 74.115 129.945 74.375 130.275 ;
        RECT 74.545 129.775 75.755 130.525 ;
        RECT 75.925 129.775 76.215 130.500 ;
        RECT 76.385 129.775 79.895 130.545 ;
        RECT 80.065 130.450 80.235 131.185 ;
        RECT 80.505 131.015 80.675 131.185 ;
        RECT 80.405 130.685 80.675 131.015 ;
        RECT 80.845 130.685 81.250 131.015 ;
        RECT 81.420 130.685 82.130 131.305 ;
        RECT 82.330 131.185 82.650 131.475 ;
        RECT 82.825 131.235 84.035 132.325 ;
        RECT 84.205 131.235 87.715 132.325 ;
        RECT 88.260 131.985 88.515 132.015 ;
        RECT 88.175 131.815 88.515 131.985 ;
        RECT 88.260 131.345 88.515 131.815 ;
        RECT 88.695 131.525 88.980 132.325 ;
        RECT 89.160 131.605 89.490 132.115 ;
        RECT 80.505 130.515 80.675 130.685 ;
        RECT 80.065 130.105 80.335 130.450 ;
        RECT 80.505 130.345 82.115 130.515 ;
        RECT 82.300 130.445 82.650 131.015 ;
        RECT 82.825 130.695 83.345 131.235 ;
        RECT 83.515 130.525 84.035 131.065 ;
        RECT 84.205 130.715 85.895 131.235 ;
        RECT 86.065 130.545 87.715 131.065 ;
        RECT 80.525 129.775 80.905 130.175 ;
        RECT 81.075 129.995 81.245 130.345 ;
        RECT 81.415 129.775 81.745 130.175 ;
        RECT 81.945 129.995 82.115 130.345 ;
        RECT 82.315 129.775 82.645 130.275 ;
        RECT 82.825 129.775 84.035 130.525 ;
        RECT 84.205 129.775 87.715 130.545 ;
        RECT 88.260 130.485 88.440 131.345 ;
        RECT 89.160 131.015 89.410 131.605 ;
        RECT 89.760 131.455 89.930 132.065 ;
        RECT 90.100 131.635 90.430 132.325 ;
        RECT 90.660 131.775 90.900 132.065 ;
        RECT 91.100 131.945 91.520 132.325 ;
        RECT 91.700 131.855 92.330 132.105 ;
        RECT 92.800 131.945 93.130 132.325 ;
        RECT 91.700 131.775 91.870 131.855 ;
        RECT 93.300 131.775 93.470 132.065 ;
        RECT 93.650 131.945 94.030 132.325 ;
        RECT 94.270 131.940 95.100 132.110 ;
        RECT 90.660 131.605 91.870 131.775 ;
        RECT 88.610 130.685 89.410 131.015 ;
        RECT 88.260 129.955 88.515 130.485 ;
        RECT 88.695 129.775 88.980 130.235 ;
        RECT 89.160 130.035 89.410 130.685 ;
        RECT 89.610 131.435 89.930 131.455 ;
        RECT 89.610 131.265 91.530 131.435 ;
        RECT 89.610 130.370 89.800 131.265 ;
        RECT 91.700 131.095 91.870 131.605 ;
        RECT 92.040 131.345 92.560 131.655 ;
        RECT 89.970 130.925 91.870 131.095 ;
        RECT 89.970 130.865 90.300 130.925 ;
        RECT 90.450 130.695 90.780 130.755 ;
        RECT 90.120 130.425 90.780 130.695 ;
        RECT 89.610 130.040 89.930 130.370 ;
        RECT 90.110 129.775 90.770 130.255 ;
        RECT 90.970 130.165 91.140 130.925 ;
        RECT 92.040 130.755 92.220 131.165 ;
        RECT 91.310 130.585 91.640 130.705 ;
        RECT 92.390 130.585 92.560 131.345 ;
        RECT 91.310 130.415 92.560 130.585 ;
        RECT 92.730 131.525 94.100 131.775 ;
        RECT 92.730 130.755 92.920 131.525 ;
        RECT 93.850 131.265 94.100 131.525 ;
        RECT 93.090 131.095 93.340 131.255 ;
        RECT 94.270 131.095 94.440 131.940 ;
        RECT 95.335 131.655 95.505 132.155 ;
        RECT 95.675 131.825 96.005 132.325 ;
        RECT 94.610 131.265 95.110 131.645 ;
        RECT 95.335 131.485 96.030 131.655 ;
        RECT 93.090 130.925 94.440 131.095 ;
        RECT 94.020 130.885 94.440 130.925 ;
        RECT 92.730 130.415 93.150 130.755 ;
        RECT 93.440 130.425 93.850 130.755 ;
        RECT 90.970 129.995 91.820 130.165 ;
        RECT 92.380 129.775 92.700 130.235 ;
        RECT 92.900 129.985 93.150 130.415 ;
        RECT 93.440 129.775 93.850 130.215 ;
        RECT 94.020 130.155 94.190 130.885 ;
        RECT 94.360 130.335 94.710 130.705 ;
        RECT 94.890 130.395 95.110 131.265 ;
        RECT 95.280 130.695 95.690 131.315 ;
        RECT 95.860 130.515 96.030 131.485 ;
        RECT 95.335 130.325 96.030 130.515 ;
        RECT 94.020 129.955 95.035 130.155 ;
        RECT 95.335 129.995 95.505 130.325 ;
        RECT 95.675 129.775 96.005 130.155 ;
        RECT 96.220 130.035 96.445 132.155 ;
        RECT 96.615 131.825 96.945 132.325 ;
        RECT 97.115 131.655 97.285 132.155 ;
        RECT 96.620 131.485 97.285 131.655 ;
        RECT 96.620 130.495 96.850 131.485 ;
        RECT 97.020 130.665 97.370 131.315 ;
        RECT 97.545 131.235 100.135 132.325 ;
        RECT 97.545 130.715 98.755 131.235 ;
        RECT 100.345 131.185 100.575 132.325 ;
        RECT 100.745 131.175 101.075 132.155 ;
        RECT 101.245 131.185 101.455 132.325 ;
        RECT 98.925 130.545 100.135 131.065 ;
        RECT 100.325 130.765 100.655 131.015 ;
        RECT 96.620 130.325 97.285 130.495 ;
        RECT 96.615 129.775 96.945 130.155 ;
        RECT 97.115 130.035 97.285 130.325 ;
        RECT 97.545 129.775 100.135 130.545 ;
        RECT 100.345 129.775 100.575 130.595 ;
        RECT 100.825 130.575 101.075 131.175 ;
        RECT 101.685 131.160 101.975 132.325 ;
        RECT 102.145 131.235 103.815 132.325 ;
        RECT 103.985 131.605 104.445 132.155 ;
        RECT 104.635 131.605 104.965 132.325 ;
        RECT 102.145 130.715 102.895 131.235 ;
        RECT 100.745 129.945 101.075 130.575 ;
        RECT 101.245 129.775 101.455 130.595 ;
        RECT 103.065 130.545 103.815 131.065 ;
        RECT 101.685 129.775 101.975 130.500 ;
        RECT 102.145 129.775 103.815 130.545 ;
        RECT 103.985 130.235 104.235 131.605 ;
        RECT 105.165 131.435 105.465 131.985 ;
        RECT 105.635 131.655 105.915 132.325 ;
        RECT 104.525 131.265 105.465 131.435 ;
        RECT 106.285 131.605 106.745 132.155 ;
        RECT 106.935 131.605 107.265 132.325 ;
        RECT 104.525 131.015 104.695 131.265 ;
        RECT 105.835 131.015 106.100 131.375 ;
        RECT 104.405 130.685 104.695 131.015 ;
        RECT 104.865 130.765 105.205 131.015 ;
        RECT 105.425 130.765 106.100 131.015 ;
        RECT 104.525 130.595 104.695 130.685 ;
        RECT 104.525 130.405 105.915 130.595 ;
        RECT 103.985 129.945 104.545 130.235 ;
        RECT 104.715 129.775 104.965 130.235 ;
        RECT 105.585 130.045 105.915 130.405 ;
        RECT 106.285 130.235 106.535 131.605 ;
        RECT 107.465 131.435 107.765 131.985 ;
        RECT 107.935 131.655 108.215 132.325 ;
        RECT 106.825 131.265 107.765 131.435 ;
        RECT 108.585 131.565 109.100 131.975 ;
        RECT 109.335 131.565 109.505 132.325 ;
        RECT 109.675 131.985 111.705 132.155 ;
        RECT 106.825 131.015 106.995 131.265 ;
        RECT 108.135 131.015 108.400 131.375 ;
        RECT 106.705 130.685 106.995 131.015 ;
        RECT 107.165 130.765 107.505 131.015 ;
        RECT 107.725 130.765 108.400 131.015 ;
        RECT 106.825 130.595 106.995 130.685 ;
        RECT 108.585 130.755 108.925 131.565 ;
        RECT 109.675 131.320 109.845 131.985 ;
        RECT 110.240 131.645 111.365 131.815 ;
        RECT 109.095 131.130 109.845 131.320 ;
        RECT 110.015 131.305 111.025 131.475 ;
        RECT 106.825 130.405 108.215 130.595 ;
        RECT 108.585 130.585 109.815 130.755 ;
        RECT 106.285 129.945 106.845 130.235 ;
        RECT 107.015 129.775 107.265 130.235 ;
        RECT 107.885 130.045 108.215 130.405 ;
        RECT 108.860 129.980 109.105 130.585 ;
        RECT 109.325 129.775 109.835 130.310 ;
        RECT 110.015 129.945 110.205 131.305 ;
        RECT 110.375 130.965 110.650 131.105 ;
        RECT 110.375 130.795 110.655 130.965 ;
        RECT 110.375 129.945 110.650 130.795 ;
        RECT 110.855 130.505 111.025 131.305 ;
        RECT 111.195 130.515 111.365 131.645 ;
        RECT 111.535 131.015 111.705 131.985 ;
        RECT 111.875 131.185 112.045 132.325 ;
        RECT 112.215 131.185 112.550 132.155 ;
        RECT 111.535 130.685 111.730 131.015 ;
        RECT 111.955 130.685 112.210 131.015 ;
        RECT 111.955 130.515 112.125 130.685 ;
        RECT 112.380 130.515 112.550 131.185 ;
        RECT 111.195 130.345 112.125 130.515 ;
        RECT 111.195 130.310 111.370 130.345 ;
        RECT 110.840 129.945 111.370 130.310 ;
        RECT 111.795 129.775 112.125 130.175 ;
        RECT 112.295 129.945 112.550 130.515 ;
        RECT 112.725 131.605 113.185 132.155 ;
        RECT 113.375 131.605 113.705 132.325 ;
        RECT 112.725 130.235 112.975 131.605 ;
        RECT 113.905 131.435 114.205 131.985 ;
        RECT 114.375 131.655 114.655 132.325 ;
        RECT 113.265 131.265 114.205 131.435 ;
        RECT 115.485 131.565 116.000 131.975 ;
        RECT 116.235 131.565 116.405 132.325 ;
        RECT 116.575 131.985 118.605 132.155 ;
        RECT 113.265 131.015 113.435 131.265 ;
        RECT 114.575 131.015 114.840 131.375 ;
        RECT 113.145 130.685 113.435 131.015 ;
        RECT 113.605 130.765 113.945 131.015 ;
        RECT 114.165 130.765 114.840 131.015 ;
        RECT 113.265 130.595 113.435 130.685 ;
        RECT 115.485 130.755 115.825 131.565 ;
        RECT 116.575 131.320 116.745 131.985 ;
        RECT 117.140 131.645 118.265 131.815 ;
        RECT 115.995 131.130 116.745 131.320 ;
        RECT 116.915 131.305 117.925 131.475 ;
        RECT 113.265 130.405 114.655 130.595 ;
        RECT 115.485 130.585 116.715 130.755 ;
        RECT 112.725 129.945 113.285 130.235 ;
        RECT 113.455 129.775 113.705 130.235 ;
        RECT 114.325 130.045 114.655 130.405 ;
        RECT 115.760 129.980 116.005 130.585 ;
        RECT 116.225 129.775 116.735 130.310 ;
        RECT 116.915 129.945 117.105 131.305 ;
        RECT 117.275 130.285 117.550 131.105 ;
        RECT 117.755 130.505 117.925 131.305 ;
        RECT 118.095 130.515 118.265 131.645 ;
        RECT 118.435 131.015 118.605 131.985 ;
        RECT 118.775 131.185 118.945 132.325 ;
        RECT 119.115 131.185 119.450 132.155 ;
        RECT 118.435 130.685 118.630 131.015 ;
        RECT 118.855 130.685 119.110 131.015 ;
        RECT 118.855 130.515 119.025 130.685 ;
        RECT 119.280 130.515 119.450 131.185 ;
        RECT 119.625 131.235 120.835 132.325 ;
        RECT 121.010 131.890 126.355 132.325 ;
        RECT 119.625 130.695 120.145 131.235 ;
        RECT 120.315 130.525 120.835 131.065 ;
        RECT 122.600 130.640 122.950 131.890 ;
        RECT 126.525 131.235 127.735 132.325 ;
        RECT 118.095 130.345 119.025 130.515 ;
        RECT 118.095 130.310 118.270 130.345 ;
        RECT 117.275 130.115 117.555 130.285 ;
        RECT 117.275 129.945 117.550 130.115 ;
        RECT 117.740 129.945 118.270 130.310 ;
        RECT 118.695 129.775 119.025 130.175 ;
        RECT 119.195 129.945 119.450 130.515 ;
        RECT 119.625 129.775 120.835 130.525 ;
        RECT 124.430 130.320 124.770 131.150 ;
        RECT 126.525 130.695 127.045 131.235 ;
        RECT 127.215 130.525 127.735 131.065 ;
        RECT 121.010 129.775 126.355 130.320 ;
        RECT 126.525 129.775 127.735 130.525 ;
        RECT 14.660 129.605 127.820 129.775 ;
        RECT 14.745 128.855 15.955 129.605 ;
        RECT 16.960 129.265 17.215 129.425 ;
        RECT 16.875 129.095 17.215 129.265 ;
        RECT 17.395 129.145 17.680 129.605 ;
        RECT 16.960 128.895 17.215 129.095 ;
        RECT 14.745 128.315 15.265 128.855 ;
        RECT 15.435 128.145 15.955 128.685 ;
        RECT 14.745 127.055 15.955 128.145 ;
        RECT 16.960 128.035 17.140 128.895 ;
        RECT 17.860 128.695 18.110 129.345 ;
        RECT 17.310 128.365 18.110 128.695 ;
        RECT 16.960 127.365 17.215 128.035 ;
        RECT 17.395 127.055 17.680 127.855 ;
        RECT 17.860 127.775 18.110 128.365 ;
        RECT 18.310 129.010 18.630 129.340 ;
        RECT 18.810 129.125 19.470 129.605 ;
        RECT 19.670 129.215 20.520 129.385 ;
        RECT 18.310 128.115 18.500 129.010 ;
        RECT 18.820 128.685 19.480 128.955 ;
        RECT 19.150 128.625 19.480 128.685 ;
        RECT 18.670 128.455 19.000 128.515 ;
        RECT 19.670 128.455 19.840 129.215 ;
        RECT 21.080 129.145 21.400 129.605 ;
        RECT 21.600 128.965 21.850 129.395 ;
        RECT 22.140 129.165 22.550 129.605 ;
        RECT 22.720 129.225 23.735 129.425 ;
        RECT 20.010 128.795 21.260 128.965 ;
        RECT 20.010 128.675 20.340 128.795 ;
        RECT 18.670 128.285 20.570 128.455 ;
        RECT 18.310 127.945 20.230 128.115 ;
        RECT 18.310 127.925 18.630 127.945 ;
        RECT 17.860 127.265 18.190 127.775 ;
        RECT 18.460 127.315 18.630 127.925 ;
        RECT 20.400 127.775 20.570 128.285 ;
        RECT 20.740 128.215 20.920 128.625 ;
        RECT 21.090 128.035 21.260 128.795 ;
        RECT 18.800 127.055 19.130 127.745 ;
        RECT 19.360 127.605 20.570 127.775 ;
        RECT 20.740 127.725 21.260 128.035 ;
        RECT 21.430 128.625 21.850 128.965 ;
        RECT 22.140 128.625 22.550 128.955 ;
        RECT 21.430 127.855 21.620 128.625 ;
        RECT 22.720 128.495 22.890 129.225 ;
        RECT 24.035 129.055 24.205 129.385 ;
        RECT 24.375 129.225 24.705 129.605 ;
        RECT 23.060 128.675 23.410 129.045 ;
        RECT 22.720 128.455 23.140 128.495 ;
        RECT 21.790 128.285 23.140 128.455 ;
        RECT 21.790 128.125 22.040 128.285 ;
        RECT 22.550 127.855 22.800 128.115 ;
        RECT 21.430 127.605 22.800 127.855 ;
        RECT 19.360 127.315 19.600 127.605 ;
        RECT 20.400 127.525 20.570 127.605 ;
        RECT 19.800 127.055 20.220 127.435 ;
        RECT 20.400 127.275 21.030 127.525 ;
        RECT 21.500 127.055 21.830 127.435 ;
        RECT 22.000 127.315 22.170 127.605 ;
        RECT 22.970 127.440 23.140 128.285 ;
        RECT 23.590 128.115 23.810 128.985 ;
        RECT 24.035 128.865 24.730 129.055 ;
        RECT 23.310 127.735 23.810 128.115 ;
        RECT 23.980 128.065 24.390 128.685 ;
        RECT 24.560 127.895 24.730 128.865 ;
        RECT 24.035 127.725 24.730 127.895 ;
        RECT 22.350 127.055 22.730 127.435 ;
        RECT 22.970 127.270 23.800 127.440 ;
        RECT 24.035 127.225 24.205 127.725 ;
        RECT 24.375 127.055 24.705 127.555 ;
        RECT 24.920 127.225 25.145 129.345 ;
        RECT 25.315 129.225 25.645 129.605 ;
        RECT 25.815 129.055 25.985 129.345 ;
        RECT 26.710 129.060 32.055 129.605 ;
        RECT 25.320 128.885 25.985 129.055 ;
        RECT 25.320 127.895 25.550 128.885 ;
        RECT 25.720 128.065 26.070 128.715 ;
        RECT 25.320 127.725 25.985 127.895 ;
        RECT 25.315 127.055 25.645 127.555 ;
        RECT 25.815 127.225 25.985 127.725 ;
        RECT 28.300 127.490 28.650 128.740 ;
        RECT 30.130 128.230 30.470 129.060 ;
        RECT 32.225 128.930 32.485 129.435 ;
        RECT 32.665 129.225 32.995 129.605 ;
        RECT 33.175 129.055 33.345 129.435 ;
        RECT 32.225 128.130 32.395 128.930 ;
        RECT 32.680 128.885 33.345 129.055 ;
        RECT 32.680 128.630 32.850 128.885 ;
        RECT 33.605 128.835 37.115 129.605 ;
        RECT 37.285 128.880 37.575 129.605 ;
        RECT 37.745 128.835 41.255 129.605 ;
        RECT 32.565 128.300 32.850 128.630 ;
        RECT 33.085 128.335 33.415 128.705 ;
        RECT 32.680 128.155 32.850 128.300 ;
        RECT 26.710 127.055 32.055 127.490 ;
        RECT 32.225 127.225 32.495 128.130 ;
        RECT 32.680 127.985 33.345 128.155 ;
        RECT 32.665 127.055 32.995 127.815 ;
        RECT 33.175 127.225 33.345 127.985 ;
        RECT 33.605 128.145 35.295 128.665 ;
        RECT 35.465 128.315 37.115 128.835 ;
        RECT 33.605 127.055 37.115 128.145 ;
        RECT 37.285 127.055 37.575 128.220 ;
        RECT 37.745 128.145 39.435 128.665 ;
        RECT 39.605 128.315 41.255 128.835 ;
        RECT 41.425 128.930 41.685 129.435 ;
        RECT 41.865 129.225 42.195 129.605 ;
        RECT 42.375 129.055 42.545 129.435 ;
        RECT 37.745 127.055 41.255 128.145 ;
        RECT 41.425 128.130 41.595 128.930 ;
        RECT 41.880 128.885 42.545 129.055 ;
        RECT 43.005 128.975 43.335 129.335 ;
        RECT 43.955 129.145 44.205 129.605 ;
        RECT 44.375 129.145 44.935 129.435 ;
        RECT 41.880 128.630 42.050 128.885 ;
        RECT 43.005 128.785 44.395 128.975 ;
        RECT 41.765 128.300 42.050 128.630 ;
        RECT 42.285 128.335 42.615 128.705 ;
        RECT 44.225 128.695 44.395 128.785 ;
        RECT 42.820 128.365 43.495 128.615 ;
        RECT 43.715 128.365 44.055 128.615 ;
        RECT 44.225 128.365 44.515 128.695 ;
        RECT 41.880 128.155 42.050 128.300 ;
        RECT 41.425 127.225 41.695 128.130 ;
        RECT 41.880 127.985 42.545 128.155 ;
        RECT 42.820 128.005 43.085 128.365 ;
        RECT 44.225 128.115 44.395 128.365 ;
        RECT 41.865 127.055 42.195 127.815 ;
        RECT 42.375 127.225 42.545 127.985 ;
        RECT 43.455 127.945 44.395 128.115 ;
        RECT 43.005 127.055 43.285 127.725 ;
        RECT 43.455 127.395 43.755 127.945 ;
        RECT 44.685 127.775 44.935 129.145 ;
        RECT 43.955 127.055 44.285 127.775 ;
        RECT 44.475 127.225 44.935 127.775 ;
        RECT 45.105 128.930 45.375 129.275 ;
        RECT 45.565 129.205 45.945 129.605 ;
        RECT 46.115 129.035 46.285 129.385 ;
        RECT 46.455 129.205 46.785 129.605 ;
        RECT 46.985 129.035 47.155 129.385 ;
        RECT 47.355 129.105 47.685 129.605 ;
        RECT 45.105 128.195 45.275 128.930 ;
        RECT 45.545 128.865 47.155 129.035 ;
        RECT 45.545 128.695 45.715 128.865 ;
        RECT 45.445 128.365 45.715 128.695 ;
        RECT 45.885 128.365 46.290 128.695 ;
        RECT 45.545 128.195 45.715 128.365 ;
        RECT 45.105 127.225 45.375 128.195 ;
        RECT 45.545 128.025 46.270 128.195 ;
        RECT 46.460 128.075 47.170 128.695 ;
        RECT 47.340 128.365 47.690 128.935 ;
        RECT 47.865 128.835 49.535 129.605 ;
        RECT 46.100 127.905 46.270 128.025 ;
        RECT 47.370 127.905 47.690 128.195 ;
        RECT 45.585 127.055 45.865 127.855 ;
        RECT 46.100 127.735 47.690 127.905 ;
        RECT 47.865 128.145 48.615 128.665 ;
        RECT 48.785 128.315 49.535 128.835 ;
        RECT 49.705 128.930 49.975 129.275 ;
        RECT 50.165 129.205 50.545 129.605 ;
        RECT 50.715 129.035 50.885 129.385 ;
        RECT 51.055 129.205 51.385 129.605 ;
        RECT 51.585 129.035 51.755 129.385 ;
        RECT 51.955 129.105 52.285 129.605 ;
        RECT 49.705 128.195 49.875 128.930 ;
        RECT 50.145 128.865 51.755 129.035 ;
        RECT 50.145 128.695 50.315 128.865 ;
        RECT 50.045 128.365 50.315 128.695 ;
        RECT 50.485 128.365 50.890 128.695 ;
        RECT 50.145 128.195 50.315 128.365 ;
        RECT 51.060 128.245 51.770 128.695 ;
        RECT 51.940 128.365 52.290 128.935 ;
        RECT 52.465 128.855 53.675 129.605 ;
        RECT 53.905 129.125 54.185 129.605 ;
        RECT 54.355 128.955 54.615 129.345 ;
        RECT 54.790 129.125 55.045 129.605 ;
        RECT 55.215 128.955 55.510 129.345 ;
        RECT 55.690 129.125 55.965 129.605 ;
        RECT 56.135 129.105 56.435 129.435 ;
        RECT 46.035 127.275 47.690 127.565 ;
        RECT 47.865 127.055 49.535 128.145 ;
        RECT 49.705 127.225 49.975 128.195 ;
        RECT 50.145 128.025 50.870 128.195 ;
        RECT 51.060 128.075 51.775 128.245 ;
        RECT 50.700 127.905 50.870 128.025 ;
        RECT 51.970 127.905 52.290 128.195 ;
        RECT 50.185 127.055 50.465 127.855 ;
        RECT 50.700 127.735 52.290 127.905 ;
        RECT 52.465 128.145 52.985 128.685 ;
        RECT 53.155 128.315 53.675 128.855 ;
        RECT 53.860 128.785 55.510 128.955 ;
        RECT 53.860 128.275 54.265 128.785 ;
        RECT 54.435 128.445 55.575 128.615 ;
        RECT 50.635 127.275 52.290 127.565 ;
        RECT 52.465 127.055 53.675 128.145 ;
        RECT 53.860 128.105 54.615 128.275 ;
        RECT 53.900 127.055 54.185 127.925 ;
        RECT 54.355 127.855 54.615 128.105 ;
        RECT 55.405 128.195 55.575 128.445 ;
        RECT 55.745 128.365 56.095 128.935 ;
        RECT 56.265 128.195 56.435 129.105 ;
        RECT 55.405 128.025 56.435 128.195 ;
        RECT 54.355 127.685 55.475 127.855 ;
        RECT 54.355 127.225 54.615 127.685 ;
        RECT 54.790 127.055 55.045 127.515 ;
        RECT 55.215 127.225 55.475 127.685 ;
        RECT 55.645 127.055 55.955 127.855 ;
        RECT 56.125 127.225 56.435 128.025 ;
        RECT 57.065 128.805 57.405 129.435 ;
        RECT 57.575 128.805 57.825 129.605 ;
        RECT 58.015 128.955 58.345 129.435 ;
        RECT 58.515 129.145 58.740 129.605 ;
        RECT 58.910 128.955 59.240 129.435 ;
        RECT 57.065 128.245 57.240 128.805 ;
        RECT 58.015 128.785 59.240 128.955 ;
        RECT 59.870 128.825 60.370 129.435 ;
        RECT 57.410 128.445 58.105 128.615 ;
        RECT 57.065 128.195 57.295 128.245 ;
        RECT 57.935 128.195 58.105 128.445 ;
        RECT 58.280 128.415 58.700 128.615 ;
        RECT 58.870 128.415 59.200 128.615 ;
        RECT 59.370 128.415 59.700 128.615 ;
        RECT 59.870 128.195 60.040 128.825 ;
        RECT 61.705 128.785 61.935 129.605 ;
        RECT 62.105 128.805 62.435 129.435 ;
        RECT 60.225 128.365 60.575 128.615 ;
        RECT 61.685 128.365 62.015 128.615 ;
        RECT 62.185 128.205 62.435 128.805 ;
        RECT 62.605 128.785 62.815 129.605 ;
        RECT 63.045 128.880 63.335 129.605 ;
        RECT 63.545 128.785 63.775 129.605 ;
        RECT 63.945 128.805 64.275 129.435 ;
        RECT 63.525 128.365 63.855 128.615 ;
        RECT 57.065 127.225 57.405 128.195 ;
        RECT 57.575 127.055 57.745 128.195 ;
        RECT 57.935 128.025 60.370 128.195 ;
        RECT 58.015 127.055 58.265 127.855 ;
        RECT 58.910 127.225 59.240 128.025 ;
        RECT 59.540 127.055 59.870 127.855 ;
        RECT 60.040 127.225 60.370 128.025 ;
        RECT 61.705 127.055 61.935 128.195 ;
        RECT 62.105 127.225 62.435 128.205 ;
        RECT 62.605 127.055 62.815 128.195 ;
        RECT 63.045 127.055 63.335 128.220 ;
        RECT 64.025 128.205 64.275 128.805 ;
        RECT 64.445 128.785 64.655 129.605 ;
        RECT 65.260 128.895 65.515 129.425 ;
        RECT 65.695 129.145 65.980 129.605 ;
        RECT 65.260 128.585 65.440 128.895 ;
        RECT 66.160 128.695 66.410 129.345 ;
        RECT 65.175 128.415 65.440 128.585 ;
        RECT 63.545 127.055 63.775 128.195 ;
        RECT 63.945 127.225 64.275 128.205 ;
        RECT 64.445 127.055 64.655 128.195 ;
        RECT 65.260 128.035 65.440 128.415 ;
        RECT 65.610 128.365 66.410 128.695 ;
        RECT 65.260 127.365 65.515 128.035 ;
        RECT 65.695 127.055 65.980 127.855 ;
        RECT 66.160 127.775 66.410 128.365 ;
        RECT 66.610 129.010 66.930 129.340 ;
        RECT 67.110 129.125 67.770 129.605 ;
        RECT 67.970 129.215 68.820 129.385 ;
        RECT 66.610 128.115 66.800 129.010 ;
        RECT 67.120 128.685 67.780 128.955 ;
        RECT 67.450 128.625 67.780 128.685 ;
        RECT 66.970 128.455 67.300 128.515 ;
        RECT 67.970 128.455 68.140 129.215 ;
        RECT 69.380 129.145 69.700 129.605 ;
        RECT 69.900 128.965 70.150 129.395 ;
        RECT 70.440 129.165 70.850 129.605 ;
        RECT 71.020 129.225 72.035 129.425 ;
        RECT 68.310 128.795 69.560 128.965 ;
        RECT 68.310 128.675 68.640 128.795 ;
        RECT 66.970 128.285 68.870 128.455 ;
        RECT 66.610 127.945 68.530 128.115 ;
        RECT 66.610 127.925 66.930 127.945 ;
        RECT 66.160 127.265 66.490 127.775 ;
        RECT 66.760 127.315 66.930 127.925 ;
        RECT 68.700 127.775 68.870 128.285 ;
        RECT 69.040 128.215 69.220 128.625 ;
        RECT 69.390 128.035 69.560 128.795 ;
        RECT 67.100 127.055 67.430 127.745 ;
        RECT 67.660 127.605 68.870 127.775 ;
        RECT 69.040 127.725 69.560 128.035 ;
        RECT 69.730 128.625 70.150 128.965 ;
        RECT 70.440 128.625 70.850 128.955 ;
        RECT 69.730 127.855 69.920 128.625 ;
        RECT 71.020 128.495 71.190 129.225 ;
        RECT 72.335 129.055 72.505 129.385 ;
        RECT 72.675 129.225 73.005 129.605 ;
        RECT 71.360 128.675 71.710 129.045 ;
        RECT 71.020 128.455 71.440 128.495 ;
        RECT 70.090 128.285 71.440 128.455 ;
        RECT 70.090 128.125 70.340 128.285 ;
        RECT 70.850 127.855 71.100 128.115 ;
        RECT 69.730 127.605 71.100 127.855 ;
        RECT 67.660 127.315 67.900 127.605 ;
        RECT 68.700 127.525 68.870 127.605 ;
        RECT 68.100 127.055 68.520 127.435 ;
        RECT 68.700 127.275 69.330 127.525 ;
        RECT 69.800 127.055 70.130 127.435 ;
        RECT 70.300 127.315 70.470 127.605 ;
        RECT 71.270 127.440 71.440 128.285 ;
        RECT 71.890 128.115 72.110 128.985 ;
        RECT 72.335 128.865 73.030 129.055 ;
        RECT 71.610 127.735 72.110 128.115 ;
        RECT 72.280 128.065 72.690 128.685 ;
        RECT 72.860 127.895 73.030 128.865 ;
        RECT 72.335 127.725 73.030 127.895 ;
        RECT 70.650 127.055 71.030 127.435 ;
        RECT 71.270 127.270 72.100 127.440 ;
        RECT 72.335 127.225 72.505 127.725 ;
        RECT 72.675 127.055 73.005 127.555 ;
        RECT 73.220 127.225 73.445 129.345 ;
        RECT 73.615 129.225 73.945 129.605 ;
        RECT 74.115 129.055 74.285 129.345 ;
        RECT 73.620 128.885 74.285 129.055 ;
        RECT 74.545 129.145 75.105 129.435 ;
        RECT 75.275 129.145 75.525 129.605 ;
        RECT 73.620 127.895 73.850 128.885 ;
        RECT 74.020 128.065 74.370 128.715 ;
        RECT 73.620 127.725 74.285 127.895 ;
        RECT 73.615 127.055 73.945 127.555 ;
        RECT 74.115 127.225 74.285 127.725 ;
        RECT 74.545 127.775 74.795 129.145 ;
        RECT 76.145 128.975 76.475 129.335 ;
        RECT 76.850 129.060 82.195 129.605 ;
        RECT 82.365 129.145 82.925 129.435 ;
        RECT 83.095 129.145 83.345 129.605 ;
        RECT 75.085 128.785 76.475 128.975 ;
        RECT 75.085 128.695 75.255 128.785 ;
        RECT 74.965 128.365 75.255 128.695 ;
        RECT 75.425 128.365 75.765 128.615 ;
        RECT 75.985 128.365 76.660 128.615 ;
        RECT 75.085 128.115 75.255 128.365 ;
        RECT 75.085 127.945 76.025 128.115 ;
        RECT 76.395 128.005 76.660 128.365 ;
        RECT 74.545 127.225 75.005 127.775 ;
        RECT 75.195 127.055 75.525 127.775 ;
        RECT 75.725 127.395 76.025 127.945 ;
        RECT 76.195 127.055 76.475 127.725 ;
        RECT 78.440 127.490 78.790 128.740 ;
        RECT 80.270 128.230 80.610 129.060 ;
        RECT 82.365 127.775 82.615 129.145 ;
        RECT 83.965 128.975 84.295 129.335 ;
        RECT 82.905 128.785 84.295 128.975 ;
        RECT 85.125 128.835 88.635 129.605 ;
        RECT 88.805 128.880 89.095 129.605 ;
        RECT 89.725 128.835 92.315 129.605 ;
        RECT 82.905 128.695 83.075 128.785 ;
        RECT 82.785 128.365 83.075 128.695 ;
        RECT 83.245 128.365 83.585 128.615 ;
        RECT 83.805 128.365 84.480 128.615 ;
        RECT 82.905 128.115 83.075 128.365 ;
        RECT 82.905 127.945 83.845 128.115 ;
        RECT 84.215 128.005 84.480 128.365 ;
        RECT 85.125 128.145 86.815 128.665 ;
        RECT 86.985 128.315 88.635 128.835 ;
        RECT 76.850 127.055 82.195 127.490 ;
        RECT 82.365 127.225 82.825 127.775 ;
        RECT 83.015 127.055 83.345 127.775 ;
        RECT 83.545 127.395 83.845 127.945 ;
        RECT 84.015 127.055 84.295 127.725 ;
        RECT 85.125 127.055 88.635 128.145 ;
        RECT 88.805 127.055 89.095 128.220 ;
        RECT 89.725 128.145 90.935 128.665 ;
        RECT 91.105 128.315 92.315 128.835 ;
        RECT 92.545 128.785 92.755 129.605 ;
        RECT 92.925 128.805 93.255 129.435 ;
        RECT 92.925 128.205 93.175 128.805 ;
        RECT 93.425 128.785 93.655 129.605 ;
        RECT 93.870 129.060 99.215 129.605 ;
        RECT 99.385 129.145 99.945 129.435 ;
        RECT 100.115 129.145 100.365 129.605 ;
        RECT 93.345 128.365 93.675 128.615 ;
        RECT 89.725 127.055 92.315 128.145 ;
        RECT 92.545 127.055 92.755 128.195 ;
        RECT 92.925 127.225 93.255 128.205 ;
        RECT 93.425 127.055 93.655 128.195 ;
        RECT 95.460 127.490 95.810 128.740 ;
        RECT 97.290 128.230 97.630 129.060 ;
        RECT 99.385 127.775 99.635 129.145 ;
        RECT 100.985 128.975 101.315 129.335 ;
        RECT 99.925 128.785 101.315 128.975 ;
        RECT 101.685 128.835 103.355 129.605 ;
        RECT 103.525 129.095 103.830 129.605 ;
        RECT 99.925 128.695 100.095 128.785 ;
        RECT 99.805 128.365 100.095 128.695 ;
        RECT 100.265 128.365 100.605 128.615 ;
        RECT 100.825 128.365 101.500 128.615 ;
        RECT 99.925 128.115 100.095 128.365 ;
        RECT 99.925 127.945 100.865 128.115 ;
        RECT 101.235 128.005 101.500 128.365 ;
        RECT 101.685 128.145 102.435 128.665 ;
        RECT 102.605 128.315 103.355 128.835 ;
        RECT 103.525 128.365 103.840 128.925 ;
        RECT 104.010 128.615 104.260 129.425 ;
        RECT 104.430 129.080 104.690 129.605 ;
        RECT 104.870 128.615 105.120 129.425 ;
        RECT 105.290 129.045 105.550 129.605 ;
        RECT 105.720 128.955 105.980 129.410 ;
        RECT 106.150 129.125 106.410 129.605 ;
        RECT 106.580 128.955 106.840 129.410 ;
        RECT 107.010 129.125 107.270 129.605 ;
        RECT 107.440 128.955 107.700 129.410 ;
        RECT 107.870 129.125 108.115 129.605 ;
        RECT 108.285 128.955 108.560 129.410 ;
        RECT 108.730 129.125 108.975 129.605 ;
        RECT 109.145 128.955 109.405 129.410 ;
        RECT 109.585 129.125 109.835 129.605 ;
        RECT 110.005 128.955 110.265 129.410 ;
        RECT 110.445 129.125 110.695 129.605 ;
        RECT 110.865 128.955 111.125 129.410 ;
        RECT 111.305 129.125 111.565 129.605 ;
        RECT 111.735 128.955 111.995 129.410 ;
        RECT 112.165 129.125 112.465 129.605 ;
        RECT 105.720 128.925 112.465 128.955 ;
        RECT 105.720 128.785 112.495 128.925 ;
        RECT 113.225 128.785 113.455 129.605 ;
        RECT 113.625 128.805 113.955 129.435 ;
        RECT 111.300 128.755 112.495 128.785 ;
        RECT 104.010 128.365 111.130 128.615 ;
        RECT 93.870 127.055 99.215 127.490 ;
        RECT 99.385 127.225 99.845 127.775 ;
        RECT 100.035 127.055 100.365 127.775 ;
        RECT 100.565 127.395 100.865 127.945 ;
        RECT 101.035 127.055 101.315 127.725 ;
        RECT 101.685 127.055 103.355 128.145 ;
        RECT 103.535 127.055 103.830 127.865 ;
        RECT 104.010 127.225 104.255 128.365 ;
        RECT 104.430 127.055 104.690 127.865 ;
        RECT 104.870 127.230 105.120 128.365 ;
        RECT 111.300 128.195 112.465 128.755 ;
        RECT 113.205 128.365 113.535 128.615 ;
        RECT 113.705 128.205 113.955 128.805 ;
        RECT 114.125 128.785 114.335 129.605 ;
        RECT 114.565 128.880 114.855 129.605 ;
        RECT 115.065 128.785 115.295 129.605 ;
        RECT 115.465 128.805 115.795 129.435 ;
        RECT 115.045 128.365 115.375 128.615 ;
        RECT 105.720 127.970 112.465 128.195 ;
        RECT 105.720 127.955 111.125 127.970 ;
        RECT 105.290 127.060 105.550 127.855 ;
        RECT 105.720 127.230 105.980 127.955 ;
        RECT 106.150 127.060 106.410 127.785 ;
        RECT 106.580 127.230 106.840 127.955 ;
        RECT 107.010 127.060 107.270 127.785 ;
        RECT 107.440 127.230 107.700 127.955 ;
        RECT 107.870 127.060 108.130 127.785 ;
        RECT 108.300 127.230 108.560 127.955 ;
        RECT 108.730 127.060 108.975 127.785 ;
        RECT 109.145 127.230 109.405 127.955 ;
        RECT 109.590 127.060 109.835 127.785 ;
        RECT 110.005 127.230 110.265 127.955 ;
        RECT 110.450 127.060 110.695 127.785 ;
        RECT 110.865 127.230 111.125 127.955 ;
        RECT 111.310 127.060 111.565 127.785 ;
        RECT 111.735 127.230 112.025 127.970 ;
        RECT 105.290 127.055 111.565 127.060 ;
        RECT 112.195 127.055 112.465 127.800 ;
        RECT 113.225 127.055 113.455 128.195 ;
        RECT 113.625 127.225 113.955 128.205 ;
        RECT 114.125 127.055 114.335 128.195 ;
        RECT 114.565 127.055 114.855 128.220 ;
        RECT 115.545 128.205 115.795 128.805 ;
        RECT 115.965 128.785 116.175 129.605 ;
        RECT 116.780 129.265 117.035 129.425 ;
        RECT 116.695 129.095 117.035 129.265 ;
        RECT 117.215 129.145 117.500 129.605 ;
        RECT 116.780 128.895 117.035 129.095 ;
        RECT 115.065 127.055 115.295 128.195 ;
        RECT 115.465 127.225 115.795 128.205 ;
        RECT 115.965 127.055 116.175 128.195 ;
        RECT 116.780 128.035 116.960 128.895 ;
        RECT 117.680 128.695 117.930 129.345 ;
        RECT 117.130 128.365 117.930 128.695 ;
        RECT 116.780 127.365 117.035 128.035 ;
        RECT 117.215 127.055 117.500 127.855 ;
        RECT 117.680 127.775 117.930 128.365 ;
        RECT 118.130 129.010 118.450 129.340 ;
        RECT 118.630 129.125 119.290 129.605 ;
        RECT 119.490 129.215 120.340 129.385 ;
        RECT 118.130 128.115 118.320 129.010 ;
        RECT 118.640 128.685 119.300 128.955 ;
        RECT 118.970 128.625 119.300 128.685 ;
        RECT 118.490 128.455 118.820 128.515 ;
        RECT 119.490 128.455 119.660 129.215 ;
        RECT 120.900 129.145 121.220 129.605 ;
        RECT 121.420 128.965 121.670 129.395 ;
        RECT 121.960 129.165 122.370 129.605 ;
        RECT 122.540 129.225 123.555 129.425 ;
        RECT 119.830 128.795 121.080 128.965 ;
        RECT 119.830 128.675 120.160 128.795 ;
        RECT 118.490 128.285 120.390 128.455 ;
        RECT 118.130 127.945 120.050 128.115 ;
        RECT 118.130 127.925 118.450 127.945 ;
        RECT 117.680 127.265 118.010 127.775 ;
        RECT 118.280 127.315 118.450 127.925 ;
        RECT 120.220 127.775 120.390 128.285 ;
        RECT 120.560 128.215 120.740 128.625 ;
        RECT 120.910 128.035 121.080 128.795 ;
        RECT 118.620 127.055 118.950 127.745 ;
        RECT 119.180 127.605 120.390 127.775 ;
        RECT 120.560 127.725 121.080 128.035 ;
        RECT 121.250 128.625 121.670 128.965 ;
        RECT 121.960 128.625 122.370 128.955 ;
        RECT 121.250 127.855 121.440 128.625 ;
        RECT 122.540 128.495 122.710 129.225 ;
        RECT 123.855 129.055 124.025 129.385 ;
        RECT 124.195 129.225 124.525 129.605 ;
        RECT 122.880 128.675 123.230 129.045 ;
        RECT 122.540 128.455 122.960 128.495 ;
        RECT 121.610 128.285 122.960 128.455 ;
        RECT 121.610 128.125 121.860 128.285 ;
        RECT 122.370 127.855 122.620 128.115 ;
        RECT 121.250 127.605 122.620 127.855 ;
        RECT 119.180 127.315 119.420 127.605 ;
        RECT 120.220 127.525 120.390 127.605 ;
        RECT 119.620 127.055 120.040 127.435 ;
        RECT 120.220 127.275 120.850 127.525 ;
        RECT 121.320 127.055 121.650 127.435 ;
        RECT 121.820 127.315 121.990 127.605 ;
        RECT 122.790 127.440 122.960 128.285 ;
        RECT 123.410 128.115 123.630 128.985 ;
        RECT 123.855 128.865 124.550 129.055 ;
        RECT 123.130 127.735 123.630 128.115 ;
        RECT 123.800 128.065 124.210 128.685 ;
        RECT 124.380 127.895 124.550 128.865 ;
        RECT 123.855 127.725 124.550 127.895 ;
        RECT 122.170 127.055 122.550 127.435 ;
        RECT 122.790 127.270 123.620 127.440 ;
        RECT 123.855 127.225 124.025 127.725 ;
        RECT 124.195 127.055 124.525 127.555 ;
        RECT 124.740 127.225 124.965 129.345 ;
        RECT 125.135 129.225 125.465 129.605 ;
        RECT 125.635 129.055 125.805 129.345 ;
        RECT 125.140 128.885 125.805 129.055 ;
        RECT 125.140 127.895 125.370 128.885 ;
        RECT 126.525 128.855 127.735 129.605 ;
        RECT 125.540 128.065 125.890 128.715 ;
        RECT 126.525 128.145 127.045 128.685 ;
        RECT 127.215 128.315 127.735 128.855 ;
        RECT 125.140 127.725 125.805 127.895 ;
        RECT 125.135 127.055 125.465 127.555 ;
        RECT 125.635 127.225 125.805 127.725 ;
        RECT 126.525 127.055 127.735 128.145 ;
        RECT 14.660 126.885 127.820 127.055 ;
        RECT 14.745 125.795 15.955 126.885 ;
        RECT 14.745 125.085 15.265 125.625 ;
        RECT 15.435 125.255 15.955 125.795 ;
        RECT 16.125 125.795 18.715 126.885 ;
        RECT 18.975 125.955 19.145 126.715 ;
        RECT 19.325 126.125 19.655 126.885 ;
        RECT 16.125 125.275 17.335 125.795 ;
        RECT 18.975 125.785 19.640 125.955 ;
        RECT 19.825 125.810 20.095 126.715 ;
        RECT 19.470 125.640 19.640 125.785 ;
        RECT 17.505 125.105 18.715 125.625 ;
        RECT 18.905 125.235 19.235 125.605 ;
        RECT 19.470 125.310 19.755 125.640 ;
        RECT 14.745 124.335 15.955 125.085 ;
        RECT 16.125 124.335 18.715 125.105 ;
        RECT 19.470 125.055 19.640 125.310 ;
        RECT 18.975 124.885 19.640 125.055 ;
        RECT 19.925 125.010 20.095 125.810 ;
        RECT 18.975 124.505 19.145 124.885 ;
        RECT 19.325 124.335 19.655 124.715 ;
        RECT 19.835 124.505 20.095 125.010 ;
        RECT 20.270 125.745 20.605 126.715 ;
        RECT 20.775 125.745 20.945 126.885 ;
        RECT 21.115 126.545 23.145 126.715 ;
        RECT 20.270 125.075 20.440 125.745 ;
        RECT 21.115 125.575 21.285 126.545 ;
        RECT 20.610 125.245 20.865 125.575 ;
        RECT 21.090 125.245 21.285 125.575 ;
        RECT 21.455 126.205 22.580 126.375 ;
        RECT 20.695 125.075 20.865 125.245 ;
        RECT 21.455 125.075 21.625 126.205 ;
        RECT 20.270 124.505 20.525 125.075 ;
        RECT 20.695 124.905 21.625 125.075 ;
        RECT 21.795 125.865 22.805 126.035 ;
        RECT 21.795 125.065 21.965 125.865 ;
        RECT 22.170 125.525 22.445 125.665 ;
        RECT 22.165 125.355 22.445 125.525 ;
        RECT 21.450 124.870 21.625 124.905 ;
        RECT 20.695 124.335 21.025 124.735 ;
        RECT 21.450 124.505 21.980 124.870 ;
        RECT 22.170 124.505 22.445 125.355 ;
        RECT 22.615 124.505 22.805 125.865 ;
        RECT 22.975 125.880 23.145 126.545 ;
        RECT 23.315 126.125 23.485 126.885 ;
        RECT 23.720 126.125 24.235 126.535 ;
        RECT 22.975 125.690 23.725 125.880 ;
        RECT 23.895 125.315 24.235 126.125 ;
        RECT 24.405 125.720 24.695 126.885 ;
        RECT 25.790 125.745 26.125 126.715 ;
        RECT 26.295 125.745 26.465 126.885 ;
        RECT 26.635 126.545 28.665 126.715 ;
        RECT 23.005 125.145 24.235 125.315 ;
        RECT 22.985 124.335 23.495 124.870 ;
        RECT 23.715 124.540 23.960 125.145 ;
        RECT 25.790 125.075 25.960 125.745 ;
        RECT 26.635 125.575 26.805 126.545 ;
        RECT 26.130 125.245 26.385 125.575 ;
        RECT 26.610 125.245 26.805 125.575 ;
        RECT 26.975 126.205 28.100 126.375 ;
        RECT 26.215 125.075 26.385 125.245 ;
        RECT 26.975 125.075 27.145 126.205 ;
        RECT 24.405 124.335 24.695 125.060 ;
        RECT 25.790 124.505 26.045 125.075 ;
        RECT 26.215 124.905 27.145 125.075 ;
        RECT 27.315 125.865 28.325 126.035 ;
        RECT 27.315 125.065 27.485 125.865 ;
        RECT 26.970 124.870 27.145 124.905 ;
        RECT 26.215 124.335 26.545 124.735 ;
        RECT 26.970 124.505 27.500 124.870 ;
        RECT 27.690 124.845 27.965 125.665 ;
        RECT 27.685 124.675 27.965 124.845 ;
        RECT 27.690 124.505 27.965 124.675 ;
        RECT 28.135 124.505 28.325 125.865 ;
        RECT 28.495 125.880 28.665 126.545 ;
        RECT 28.835 126.125 29.005 126.885 ;
        RECT 29.240 126.125 29.755 126.535 ;
        RECT 28.495 125.690 29.245 125.880 ;
        RECT 29.415 125.315 29.755 126.125 ;
        RECT 28.525 125.145 29.755 125.315 ;
        RECT 30.385 125.795 32.975 126.885 ;
        RECT 33.145 126.125 33.660 126.535 ;
        RECT 33.895 126.125 34.065 126.885 ;
        RECT 34.235 126.545 36.265 126.715 ;
        RECT 30.385 125.275 31.595 125.795 ;
        RECT 28.505 124.335 29.015 124.870 ;
        RECT 29.235 124.540 29.480 125.145 ;
        RECT 31.765 125.105 32.975 125.625 ;
        RECT 33.145 125.315 33.485 126.125 ;
        RECT 34.235 125.880 34.405 126.545 ;
        RECT 34.800 126.205 35.925 126.375 ;
        RECT 33.655 125.690 34.405 125.880 ;
        RECT 34.575 125.865 35.585 126.035 ;
        RECT 33.145 125.145 34.375 125.315 ;
        RECT 30.385 124.335 32.975 125.105 ;
        RECT 33.420 124.540 33.665 125.145 ;
        RECT 33.885 124.335 34.395 124.870 ;
        RECT 34.575 124.505 34.765 125.865 ;
        RECT 34.935 124.845 35.210 125.665 ;
        RECT 35.415 125.065 35.585 125.865 ;
        RECT 35.755 125.075 35.925 126.205 ;
        RECT 36.095 125.575 36.265 126.545 ;
        RECT 36.435 125.745 36.605 126.885 ;
        RECT 36.775 125.745 37.110 126.715 ;
        RECT 36.095 125.245 36.290 125.575 ;
        RECT 36.515 125.245 36.770 125.575 ;
        RECT 36.515 125.075 36.685 125.245 ;
        RECT 36.940 125.075 37.110 125.745 ;
        RECT 37.745 125.795 39.415 126.885 ;
        RECT 39.785 126.215 40.065 126.885 ;
        RECT 40.235 125.995 40.535 126.545 ;
        RECT 40.735 126.165 41.065 126.885 ;
        RECT 41.255 126.165 41.715 126.715 ;
        RECT 42.085 126.215 42.365 126.885 ;
        RECT 37.745 125.275 38.495 125.795 ;
        RECT 38.665 125.105 39.415 125.625 ;
        RECT 39.600 125.575 39.865 125.935 ;
        RECT 40.235 125.825 41.175 125.995 ;
        RECT 41.005 125.575 41.175 125.825 ;
        RECT 39.600 125.325 40.275 125.575 ;
        RECT 40.495 125.325 40.835 125.575 ;
        RECT 41.005 125.245 41.295 125.575 ;
        RECT 41.005 125.155 41.175 125.245 ;
        RECT 35.755 124.905 36.685 125.075 ;
        RECT 35.755 124.870 35.930 124.905 ;
        RECT 34.935 124.675 35.215 124.845 ;
        RECT 34.935 124.505 35.210 124.675 ;
        RECT 35.400 124.505 35.930 124.870 ;
        RECT 36.355 124.335 36.685 124.735 ;
        RECT 36.855 124.505 37.110 125.075 ;
        RECT 37.745 124.335 39.415 125.105 ;
        RECT 39.785 124.965 41.175 125.155 ;
        RECT 39.785 124.605 40.115 124.965 ;
        RECT 41.465 124.795 41.715 126.165 ;
        RECT 42.535 125.995 42.835 126.545 ;
        RECT 43.035 126.165 43.365 126.885 ;
        RECT 43.555 126.165 44.015 126.715 ;
        RECT 44.385 126.215 44.665 126.885 ;
        RECT 41.900 125.575 42.165 125.935 ;
        RECT 42.535 125.825 43.475 125.995 ;
        RECT 43.305 125.575 43.475 125.825 ;
        RECT 41.900 125.325 42.575 125.575 ;
        RECT 42.795 125.325 43.135 125.575 ;
        RECT 43.305 125.245 43.595 125.575 ;
        RECT 43.305 125.155 43.475 125.245 ;
        RECT 40.735 124.335 40.985 124.795 ;
        RECT 41.155 124.505 41.715 124.795 ;
        RECT 42.085 124.965 43.475 125.155 ;
        RECT 42.085 124.605 42.415 124.965 ;
        RECT 43.765 124.795 44.015 126.165 ;
        RECT 44.835 125.995 45.135 126.545 ;
        RECT 45.335 126.165 45.665 126.885 ;
        RECT 45.855 126.165 46.315 126.715 ;
        RECT 44.200 125.575 44.465 125.935 ;
        RECT 44.835 125.825 45.775 125.995 ;
        RECT 45.605 125.575 45.775 125.825 ;
        RECT 44.200 125.325 44.875 125.575 ;
        RECT 45.095 125.325 45.435 125.575 ;
        RECT 45.605 125.245 45.895 125.575 ;
        RECT 45.605 125.155 45.775 125.245 ;
        RECT 43.035 124.335 43.285 124.795 ;
        RECT 43.455 124.505 44.015 124.795 ;
        RECT 44.385 124.965 45.775 125.155 ;
        RECT 44.385 124.605 44.715 124.965 ;
        RECT 46.065 124.795 46.315 126.165 ;
        RECT 46.485 125.795 47.695 126.885 ;
        RECT 48.065 126.215 48.345 126.885 ;
        RECT 48.515 125.995 48.815 126.545 ;
        RECT 49.015 126.165 49.345 126.885 ;
        RECT 49.535 126.165 49.995 126.715 ;
        RECT 46.485 125.255 47.005 125.795 ;
        RECT 47.175 125.085 47.695 125.625 ;
        RECT 47.880 125.575 48.145 125.935 ;
        RECT 48.515 125.825 49.455 125.995 ;
        RECT 49.285 125.575 49.455 125.825 ;
        RECT 47.880 125.325 48.555 125.575 ;
        RECT 48.775 125.325 49.115 125.575 ;
        RECT 49.285 125.245 49.575 125.575 ;
        RECT 49.285 125.155 49.455 125.245 ;
        RECT 45.335 124.335 45.585 124.795 ;
        RECT 45.755 124.505 46.315 124.795 ;
        RECT 46.485 124.335 47.695 125.085 ;
        RECT 48.065 124.965 49.455 125.155 ;
        RECT 48.065 124.605 48.395 124.965 ;
        RECT 49.745 124.795 49.995 126.165 ;
        RECT 50.165 125.720 50.455 126.885 ;
        RECT 50.625 125.795 51.835 126.885 ;
        RECT 52.005 125.795 55.515 126.885 ;
        RECT 55.690 126.450 61.035 126.885 ;
        RECT 50.625 125.255 51.145 125.795 ;
        RECT 51.315 125.085 51.835 125.625 ;
        RECT 52.005 125.275 53.695 125.795 ;
        RECT 53.865 125.105 55.515 125.625 ;
        RECT 57.280 125.200 57.630 126.450 ;
        RECT 61.580 125.905 61.835 126.575 ;
        RECT 62.015 126.085 62.300 126.885 ;
        RECT 62.480 126.165 62.810 126.675 ;
        RECT 49.015 124.335 49.265 124.795 ;
        RECT 49.435 124.505 49.995 124.795 ;
        RECT 50.165 124.335 50.455 125.060 ;
        RECT 50.625 124.335 51.835 125.085 ;
        RECT 52.005 124.335 55.515 125.105 ;
        RECT 59.110 124.880 59.450 125.710 ;
        RECT 61.580 125.185 61.760 125.905 ;
        RECT 62.480 125.575 62.730 126.165 ;
        RECT 63.080 126.015 63.250 126.625 ;
        RECT 63.420 126.195 63.750 126.885 ;
        RECT 63.980 126.335 64.220 126.625 ;
        RECT 64.420 126.505 64.840 126.885 ;
        RECT 65.020 126.415 65.650 126.665 ;
        RECT 66.120 126.505 66.450 126.885 ;
        RECT 65.020 126.335 65.190 126.415 ;
        RECT 66.620 126.335 66.790 126.625 ;
        RECT 66.970 126.505 67.350 126.885 ;
        RECT 67.590 126.500 68.420 126.670 ;
        RECT 63.980 126.165 65.190 126.335 ;
        RECT 61.930 125.245 62.730 125.575 ;
        RECT 61.495 125.045 61.760 125.185 ;
        RECT 61.495 125.015 61.835 125.045 ;
        RECT 55.690 124.335 61.035 124.880 ;
        RECT 61.580 124.515 61.835 125.015 ;
        RECT 62.015 124.335 62.300 124.795 ;
        RECT 62.480 124.595 62.730 125.245 ;
        RECT 62.930 125.995 63.250 126.015 ;
        RECT 62.930 125.825 64.850 125.995 ;
        RECT 62.930 124.930 63.120 125.825 ;
        RECT 65.020 125.655 65.190 126.165 ;
        RECT 65.360 125.905 65.880 126.215 ;
        RECT 63.290 125.485 65.190 125.655 ;
        RECT 63.290 125.425 63.620 125.485 ;
        RECT 63.770 125.255 64.100 125.315 ;
        RECT 63.440 124.985 64.100 125.255 ;
        RECT 62.930 124.600 63.250 124.930 ;
        RECT 63.430 124.335 64.090 124.815 ;
        RECT 64.290 124.725 64.460 125.485 ;
        RECT 65.360 125.315 65.540 125.725 ;
        RECT 64.630 125.145 64.960 125.265 ;
        RECT 65.710 125.145 65.880 125.905 ;
        RECT 64.630 124.975 65.880 125.145 ;
        RECT 66.050 126.085 67.420 126.335 ;
        RECT 66.050 125.315 66.240 126.085 ;
        RECT 67.170 125.825 67.420 126.085 ;
        RECT 66.410 125.655 66.660 125.815 ;
        RECT 67.590 125.655 67.760 126.500 ;
        RECT 68.655 126.215 68.825 126.715 ;
        RECT 68.995 126.385 69.325 126.885 ;
        RECT 67.930 125.825 68.430 126.205 ;
        RECT 68.655 126.045 69.350 126.215 ;
        RECT 66.410 125.485 67.760 125.655 ;
        RECT 67.340 125.445 67.760 125.485 ;
        RECT 66.050 124.975 66.470 125.315 ;
        RECT 66.760 124.985 67.170 125.315 ;
        RECT 64.290 124.555 65.140 124.725 ;
        RECT 65.700 124.335 66.020 124.795 ;
        RECT 66.220 124.545 66.470 124.975 ;
        RECT 66.760 124.335 67.170 124.775 ;
        RECT 67.340 124.715 67.510 125.445 ;
        RECT 67.680 124.895 68.030 125.265 ;
        RECT 68.210 124.955 68.430 125.825 ;
        RECT 68.600 125.255 69.010 125.875 ;
        RECT 69.180 125.075 69.350 126.045 ;
        RECT 68.655 124.885 69.350 125.075 ;
        RECT 67.340 124.515 68.355 124.715 ;
        RECT 68.655 124.555 68.825 124.885 ;
        RECT 68.995 124.335 69.325 124.715 ;
        RECT 69.540 124.595 69.765 126.715 ;
        RECT 69.935 126.385 70.265 126.885 ;
        RECT 70.435 126.215 70.605 126.715 ;
        RECT 69.940 126.045 70.605 126.215 ;
        RECT 69.940 125.055 70.170 126.045 ;
        RECT 70.340 125.225 70.690 125.875 ;
        RECT 70.865 125.810 71.135 126.715 ;
        RECT 71.305 126.125 71.635 126.885 ;
        RECT 71.815 125.955 71.985 126.715 ;
        RECT 69.940 124.885 70.605 125.055 ;
        RECT 69.935 124.335 70.265 124.715 ;
        RECT 70.435 124.595 70.605 124.885 ;
        RECT 70.865 125.010 71.035 125.810 ;
        RECT 71.320 125.785 71.985 125.955 ;
        RECT 73.165 125.915 73.475 126.715 ;
        RECT 73.645 126.085 73.955 126.885 ;
        RECT 74.125 126.255 74.385 126.715 ;
        RECT 74.555 126.425 74.810 126.885 ;
        RECT 74.985 126.255 75.245 126.715 ;
        RECT 74.125 126.085 75.245 126.255 ;
        RECT 71.320 125.640 71.490 125.785 ;
        RECT 71.205 125.310 71.490 125.640 ;
        RECT 73.165 125.745 74.195 125.915 ;
        RECT 71.320 125.055 71.490 125.310 ;
        RECT 71.725 125.235 72.055 125.605 ;
        RECT 70.865 124.505 71.125 125.010 ;
        RECT 71.320 124.885 71.985 125.055 ;
        RECT 71.305 124.335 71.635 124.715 ;
        RECT 71.815 124.505 71.985 124.885 ;
        RECT 73.165 124.835 73.335 125.745 ;
        RECT 73.505 125.005 73.855 125.575 ;
        RECT 74.025 125.495 74.195 125.745 ;
        RECT 74.985 125.835 75.245 126.085 ;
        RECT 75.415 126.015 75.700 126.885 ;
        RECT 74.985 125.665 75.740 125.835 ;
        RECT 75.925 125.720 76.215 126.885 ;
        RECT 76.385 125.795 78.055 126.885 ;
        RECT 78.225 126.165 78.685 126.715 ;
        RECT 78.875 126.165 79.205 126.885 ;
        RECT 74.025 125.325 75.165 125.495 ;
        RECT 75.335 125.155 75.740 125.665 ;
        RECT 76.385 125.275 77.135 125.795 ;
        RECT 74.090 124.985 75.740 125.155 ;
        RECT 77.305 125.105 78.055 125.625 ;
        RECT 73.165 124.505 73.465 124.835 ;
        RECT 73.635 124.335 73.910 124.815 ;
        RECT 74.090 124.595 74.385 124.985 ;
        RECT 74.555 124.335 74.810 124.815 ;
        RECT 74.985 124.595 75.245 124.985 ;
        RECT 75.415 124.335 75.695 124.815 ;
        RECT 75.925 124.335 76.215 125.060 ;
        RECT 76.385 124.335 78.055 125.105 ;
        RECT 78.225 124.795 78.475 126.165 ;
        RECT 79.405 125.995 79.705 126.545 ;
        RECT 79.875 126.215 80.155 126.885 ;
        RECT 80.725 126.215 81.005 126.885 ;
        RECT 78.765 125.825 79.705 125.995 ;
        RECT 81.175 125.995 81.475 126.545 ;
        RECT 81.675 126.165 82.005 126.885 ;
        RECT 82.195 126.165 82.655 126.715 ;
        RECT 78.765 125.575 78.935 125.825 ;
        RECT 80.075 125.575 80.340 125.935 ;
        RECT 78.645 125.245 78.935 125.575 ;
        RECT 79.105 125.325 79.445 125.575 ;
        RECT 79.665 125.325 80.340 125.575 ;
        RECT 80.540 125.575 80.805 125.935 ;
        RECT 81.175 125.825 82.115 125.995 ;
        RECT 81.945 125.575 82.115 125.825 ;
        RECT 80.540 125.325 81.215 125.575 ;
        RECT 81.435 125.325 81.775 125.575 ;
        RECT 78.765 125.155 78.935 125.245 ;
        RECT 81.945 125.245 82.235 125.575 ;
        RECT 81.945 125.155 82.115 125.245 ;
        RECT 78.765 124.965 80.155 125.155 ;
        RECT 78.225 124.505 78.785 124.795 ;
        RECT 78.955 124.335 79.205 124.795 ;
        RECT 79.825 124.605 80.155 124.965 ;
        RECT 80.725 124.965 82.115 125.155 ;
        RECT 80.725 124.605 81.055 124.965 ;
        RECT 82.405 124.795 82.655 126.165 ;
        RECT 81.675 124.335 81.925 124.795 ;
        RECT 82.095 124.505 82.655 124.795 ;
        RECT 82.825 126.165 83.285 126.715 ;
        RECT 83.475 126.165 83.805 126.885 ;
        RECT 82.825 124.795 83.075 126.165 ;
        RECT 84.005 125.995 84.305 126.545 ;
        RECT 84.475 126.215 84.755 126.885 ;
        RECT 85.590 126.450 90.935 126.885 ;
        RECT 91.110 126.450 96.455 126.885 ;
        RECT 83.365 125.825 84.305 125.995 ;
        RECT 83.365 125.575 83.535 125.825 ;
        RECT 84.675 125.575 84.940 125.935 ;
        RECT 83.245 125.245 83.535 125.575 ;
        RECT 83.705 125.325 84.045 125.575 ;
        RECT 84.265 125.325 84.940 125.575 ;
        RECT 83.365 125.155 83.535 125.245 ;
        RECT 87.180 125.200 87.530 126.450 ;
        RECT 83.365 124.965 84.755 125.155 ;
        RECT 82.825 124.505 83.385 124.795 ;
        RECT 83.555 124.335 83.805 124.795 ;
        RECT 84.425 124.605 84.755 124.965 ;
        RECT 89.010 124.880 89.350 125.710 ;
        RECT 92.700 125.200 93.050 126.450 ;
        RECT 96.715 125.955 96.885 126.715 ;
        RECT 97.065 126.125 97.395 126.885 ;
        RECT 96.715 125.785 97.380 125.955 ;
        RECT 97.565 125.810 97.835 126.715 ;
        RECT 94.530 124.880 94.870 125.710 ;
        RECT 97.210 125.640 97.380 125.785 ;
        RECT 96.645 125.235 96.975 125.605 ;
        RECT 97.210 125.310 97.495 125.640 ;
        RECT 97.210 125.055 97.380 125.310 ;
        RECT 96.715 124.885 97.380 125.055 ;
        RECT 97.665 125.010 97.835 125.810 ;
        RECT 98.005 125.795 101.515 126.885 ;
        RECT 98.005 125.275 99.695 125.795 ;
        RECT 101.685 125.720 101.975 126.885 ;
        RECT 102.645 125.745 102.875 126.885 ;
        RECT 103.045 125.735 103.375 126.715 ;
        RECT 103.545 125.745 103.755 126.885 ;
        RECT 104.360 125.905 104.615 126.575 ;
        RECT 104.795 126.085 105.080 126.885 ;
        RECT 105.260 126.165 105.590 126.675 ;
        RECT 99.865 125.105 101.515 125.625 ;
        RECT 102.625 125.325 102.955 125.575 ;
        RECT 85.590 124.335 90.935 124.880 ;
        RECT 91.110 124.335 96.455 124.880 ;
        RECT 96.715 124.505 96.885 124.885 ;
        RECT 97.065 124.335 97.395 124.715 ;
        RECT 97.575 124.505 97.835 125.010 ;
        RECT 98.005 124.335 101.515 125.105 ;
        RECT 101.685 124.335 101.975 125.060 ;
        RECT 102.645 124.335 102.875 125.155 ;
        RECT 103.125 125.135 103.375 125.735 ;
        RECT 103.045 124.505 103.375 125.135 ;
        RECT 103.545 124.335 103.755 125.155 ;
        RECT 104.360 125.045 104.540 125.905 ;
        RECT 105.260 125.575 105.510 126.165 ;
        RECT 105.860 126.015 106.030 126.625 ;
        RECT 106.200 126.195 106.530 126.885 ;
        RECT 106.760 126.335 107.000 126.625 ;
        RECT 107.200 126.505 107.620 126.885 ;
        RECT 107.800 126.415 108.430 126.665 ;
        RECT 108.900 126.505 109.230 126.885 ;
        RECT 107.800 126.335 107.970 126.415 ;
        RECT 109.400 126.335 109.570 126.625 ;
        RECT 109.750 126.505 110.130 126.885 ;
        RECT 110.370 126.500 111.200 126.670 ;
        RECT 106.760 126.165 107.970 126.335 ;
        RECT 104.710 125.245 105.510 125.575 ;
        RECT 104.360 124.845 104.615 125.045 ;
        RECT 104.275 124.675 104.615 124.845 ;
        RECT 104.360 124.515 104.615 124.675 ;
        RECT 104.795 124.335 105.080 124.795 ;
        RECT 105.260 124.595 105.510 125.245 ;
        RECT 105.710 125.995 106.030 126.015 ;
        RECT 105.710 125.825 107.630 125.995 ;
        RECT 105.710 124.930 105.900 125.825 ;
        RECT 107.800 125.655 107.970 126.165 ;
        RECT 108.140 125.905 108.660 126.215 ;
        RECT 106.070 125.485 107.970 125.655 ;
        RECT 106.070 125.425 106.400 125.485 ;
        RECT 106.550 125.255 106.880 125.315 ;
        RECT 106.220 124.985 106.880 125.255 ;
        RECT 105.710 124.600 106.030 124.930 ;
        RECT 106.210 124.335 106.870 124.815 ;
        RECT 107.070 124.725 107.240 125.485 ;
        RECT 108.140 125.315 108.320 125.725 ;
        RECT 107.410 125.145 107.740 125.265 ;
        RECT 108.490 125.145 108.660 125.905 ;
        RECT 107.410 124.975 108.660 125.145 ;
        RECT 108.830 126.085 110.200 126.335 ;
        RECT 108.830 125.315 109.020 126.085 ;
        RECT 109.950 125.825 110.200 126.085 ;
        RECT 109.190 125.655 109.440 125.815 ;
        RECT 110.370 125.655 110.540 126.500 ;
        RECT 111.435 126.215 111.605 126.715 ;
        RECT 111.775 126.385 112.105 126.885 ;
        RECT 110.710 125.825 111.210 126.205 ;
        RECT 111.435 126.045 112.130 126.215 ;
        RECT 109.190 125.485 110.540 125.655 ;
        RECT 110.120 125.445 110.540 125.485 ;
        RECT 108.830 124.975 109.250 125.315 ;
        RECT 109.540 124.985 109.950 125.315 ;
        RECT 107.070 124.555 107.920 124.725 ;
        RECT 108.480 124.335 108.800 124.795 ;
        RECT 109.000 124.545 109.250 124.975 ;
        RECT 109.540 124.335 109.950 124.775 ;
        RECT 110.120 124.715 110.290 125.445 ;
        RECT 110.460 124.895 110.810 125.265 ;
        RECT 110.990 124.955 111.210 125.825 ;
        RECT 111.380 125.255 111.790 125.875 ;
        RECT 111.960 125.075 112.130 126.045 ;
        RECT 111.435 124.885 112.130 125.075 ;
        RECT 110.120 124.515 111.135 124.715 ;
        RECT 111.435 124.555 111.605 124.885 ;
        RECT 111.775 124.335 112.105 124.715 ;
        RECT 112.320 124.595 112.545 126.715 ;
        RECT 112.715 126.385 113.045 126.885 ;
        RECT 113.215 126.215 113.385 126.715 ;
        RECT 112.720 126.045 113.385 126.215 ;
        RECT 112.720 125.055 112.950 126.045 ;
        RECT 113.120 125.225 113.470 125.875 ;
        RECT 113.645 125.810 113.915 126.715 ;
        RECT 114.085 126.125 114.415 126.885 ;
        RECT 114.595 125.955 114.765 126.715 ;
        RECT 112.720 124.885 113.385 125.055 ;
        RECT 112.715 124.335 113.045 124.715 ;
        RECT 113.215 124.595 113.385 124.885 ;
        RECT 113.645 125.010 113.815 125.810 ;
        RECT 114.100 125.785 114.765 125.955 ;
        RECT 115.860 125.905 116.115 126.575 ;
        RECT 116.295 126.085 116.580 126.885 ;
        RECT 116.760 126.165 117.090 126.675 ;
        RECT 115.860 125.865 116.040 125.905 ;
        RECT 114.100 125.640 114.270 125.785 ;
        RECT 115.775 125.695 116.040 125.865 ;
        RECT 113.985 125.310 114.270 125.640 ;
        RECT 114.100 125.055 114.270 125.310 ;
        RECT 114.505 125.235 114.835 125.605 ;
        RECT 113.645 124.505 113.905 125.010 ;
        RECT 114.100 124.885 114.765 125.055 ;
        RECT 114.085 124.335 114.415 124.715 ;
        RECT 114.595 124.505 114.765 124.885 ;
        RECT 115.860 125.045 116.040 125.695 ;
        RECT 116.760 125.575 117.010 126.165 ;
        RECT 117.360 126.015 117.530 126.625 ;
        RECT 117.700 126.195 118.030 126.885 ;
        RECT 118.260 126.335 118.500 126.625 ;
        RECT 118.700 126.505 119.120 126.885 ;
        RECT 119.300 126.415 119.930 126.665 ;
        RECT 120.400 126.505 120.730 126.885 ;
        RECT 119.300 126.335 119.470 126.415 ;
        RECT 120.900 126.335 121.070 126.625 ;
        RECT 121.250 126.505 121.630 126.885 ;
        RECT 121.870 126.500 122.700 126.670 ;
        RECT 118.260 126.165 119.470 126.335 ;
        RECT 116.210 125.245 117.010 125.575 ;
        RECT 115.860 124.515 116.115 125.045 ;
        RECT 116.295 124.335 116.580 124.795 ;
        RECT 116.760 124.595 117.010 125.245 ;
        RECT 117.210 125.995 117.530 126.015 ;
        RECT 117.210 125.825 119.130 125.995 ;
        RECT 117.210 124.930 117.400 125.825 ;
        RECT 119.300 125.655 119.470 126.165 ;
        RECT 119.640 125.905 120.160 126.215 ;
        RECT 117.570 125.485 119.470 125.655 ;
        RECT 117.570 125.425 117.900 125.485 ;
        RECT 118.050 125.255 118.380 125.315 ;
        RECT 117.720 124.985 118.380 125.255 ;
        RECT 117.210 124.600 117.530 124.930 ;
        RECT 117.710 124.335 118.370 124.815 ;
        RECT 118.570 124.725 118.740 125.485 ;
        RECT 119.640 125.315 119.820 125.725 ;
        RECT 118.910 125.145 119.240 125.265 ;
        RECT 119.990 125.145 120.160 125.905 ;
        RECT 118.910 124.975 120.160 125.145 ;
        RECT 120.330 126.085 121.700 126.335 ;
        RECT 120.330 125.315 120.520 126.085 ;
        RECT 121.450 125.825 121.700 126.085 ;
        RECT 120.690 125.655 120.940 125.815 ;
        RECT 121.870 125.655 122.040 126.500 ;
        RECT 122.935 126.215 123.105 126.715 ;
        RECT 123.275 126.385 123.605 126.885 ;
        RECT 122.210 125.825 122.710 126.205 ;
        RECT 122.935 126.045 123.630 126.215 ;
        RECT 120.690 125.485 122.040 125.655 ;
        RECT 121.620 125.445 122.040 125.485 ;
        RECT 120.330 124.975 120.750 125.315 ;
        RECT 121.040 124.985 121.450 125.315 ;
        RECT 118.570 124.555 119.420 124.725 ;
        RECT 119.980 124.335 120.300 124.795 ;
        RECT 120.500 124.545 120.750 124.975 ;
        RECT 121.040 124.335 121.450 124.775 ;
        RECT 121.620 124.715 121.790 125.445 ;
        RECT 121.960 124.895 122.310 125.265 ;
        RECT 122.490 124.955 122.710 125.825 ;
        RECT 122.880 125.255 123.290 125.875 ;
        RECT 123.460 125.075 123.630 126.045 ;
        RECT 122.935 124.885 123.630 125.075 ;
        RECT 121.620 124.515 122.635 124.715 ;
        RECT 122.935 124.555 123.105 124.885 ;
        RECT 123.275 124.335 123.605 124.715 ;
        RECT 123.820 124.595 124.045 126.715 ;
        RECT 124.215 126.385 124.545 126.885 ;
        RECT 124.715 126.215 124.885 126.715 ;
        RECT 124.220 126.045 124.885 126.215 ;
        RECT 124.220 125.055 124.450 126.045 ;
        RECT 124.620 125.225 124.970 125.875 ;
        RECT 125.145 125.810 125.415 126.715 ;
        RECT 125.585 126.125 125.915 126.885 ;
        RECT 126.095 125.955 126.265 126.715 ;
        RECT 124.220 124.885 124.885 125.055 ;
        RECT 124.215 124.335 124.545 124.715 ;
        RECT 124.715 124.595 124.885 124.885 ;
        RECT 125.145 125.010 125.315 125.810 ;
        RECT 125.600 125.785 126.265 125.955 ;
        RECT 126.525 125.795 127.735 126.885 ;
        RECT 125.600 125.640 125.770 125.785 ;
        RECT 125.485 125.310 125.770 125.640 ;
        RECT 125.600 125.055 125.770 125.310 ;
        RECT 126.005 125.235 126.335 125.605 ;
        RECT 126.525 125.255 127.045 125.795 ;
        RECT 127.215 125.085 127.735 125.625 ;
        RECT 125.145 124.505 125.405 125.010 ;
        RECT 125.600 124.885 126.265 125.055 ;
        RECT 125.585 124.335 125.915 124.715 ;
        RECT 126.095 124.505 126.265 124.885 ;
        RECT 126.525 124.335 127.735 125.085 ;
        RECT 14.660 124.165 127.820 124.335 ;
        RECT 14.745 123.415 15.955 124.165 ;
        RECT 16.500 123.825 16.755 123.985 ;
        RECT 16.415 123.655 16.755 123.825 ;
        RECT 16.935 123.705 17.220 124.165 ;
        RECT 16.500 123.455 16.755 123.655 ;
        RECT 14.745 122.875 15.265 123.415 ;
        RECT 15.435 122.705 15.955 123.245 ;
        RECT 14.745 121.615 15.955 122.705 ;
        RECT 16.500 122.595 16.680 123.455 ;
        RECT 17.400 123.255 17.650 123.905 ;
        RECT 16.850 122.925 17.650 123.255 ;
        RECT 16.500 121.925 16.755 122.595 ;
        RECT 16.935 121.615 17.220 122.415 ;
        RECT 17.400 122.335 17.650 122.925 ;
        RECT 17.850 123.570 18.170 123.900 ;
        RECT 18.350 123.685 19.010 124.165 ;
        RECT 19.210 123.775 20.060 123.945 ;
        RECT 17.850 122.675 18.040 123.570 ;
        RECT 18.360 123.245 19.020 123.515 ;
        RECT 18.690 123.185 19.020 123.245 ;
        RECT 18.210 123.015 18.540 123.075 ;
        RECT 19.210 123.015 19.380 123.775 ;
        RECT 20.620 123.705 20.940 124.165 ;
        RECT 21.140 123.525 21.390 123.955 ;
        RECT 21.680 123.725 22.090 124.165 ;
        RECT 22.260 123.785 23.275 123.985 ;
        RECT 19.550 123.355 20.800 123.525 ;
        RECT 19.550 123.235 19.880 123.355 ;
        RECT 18.210 122.845 20.110 123.015 ;
        RECT 17.850 122.505 19.770 122.675 ;
        RECT 17.850 122.485 18.170 122.505 ;
        RECT 17.400 121.825 17.730 122.335 ;
        RECT 18.000 121.875 18.170 122.485 ;
        RECT 19.940 122.335 20.110 122.845 ;
        RECT 20.280 122.775 20.460 123.185 ;
        RECT 20.630 122.595 20.800 123.355 ;
        RECT 18.340 121.615 18.670 122.305 ;
        RECT 18.900 122.165 20.110 122.335 ;
        RECT 20.280 122.285 20.800 122.595 ;
        RECT 20.970 123.185 21.390 123.525 ;
        RECT 21.680 123.185 22.090 123.515 ;
        RECT 20.970 122.415 21.160 123.185 ;
        RECT 22.260 123.055 22.430 123.785 ;
        RECT 23.575 123.615 23.745 123.945 ;
        RECT 23.915 123.785 24.245 124.165 ;
        RECT 22.600 123.235 22.950 123.605 ;
        RECT 22.260 123.015 22.680 123.055 ;
        RECT 21.330 122.845 22.680 123.015 ;
        RECT 21.330 122.685 21.580 122.845 ;
        RECT 22.090 122.415 22.340 122.675 ;
        RECT 20.970 122.165 22.340 122.415 ;
        RECT 18.900 121.875 19.140 122.165 ;
        RECT 19.940 122.085 20.110 122.165 ;
        RECT 19.340 121.615 19.760 121.995 ;
        RECT 19.940 121.835 20.570 122.085 ;
        RECT 21.040 121.615 21.370 121.995 ;
        RECT 21.540 121.875 21.710 122.165 ;
        RECT 22.510 122.000 22.680 122.845 ;
        RECT 23.130 122.675 23.350 123.545 ;
        RECT 23.575 123.425 24.270 123.615 ;
        RECT 22.850 122.295 23.350 122.675 ;
        RECT 23.520 122.625 23.930 123.245 ;
        RECT 24.100 122.455 24.270 123.425 ;
        RECT 23.575 122.285 24.270 122.455 ;
        RECT 21.890 121.615 22.270 121.995 ;
        RECT 22.510 121.830 23.340 122.000 ;
        RECT 23.575 121.785 23.745 122.285 ;
        RECT 23.915 121.615 24.245 122.115 ;
        RECT 24.460 121.785 24.685 123.905 ;
        RECT 24.855 123.785 25.185 124.165 ;
        RECT 25.355 123.615 25.525 123.905 ;
        RECT 24.860 123.445 25.525 123.615 ;
        RECT 24.860 122.455 25.090 123.445 ;
        RECT 26.245 123.395 27.915 124.165 ;
        RECT 28.175 123.685 28.475 124.165 ;
        RECT 28.645 123.515 28.905 123.970 ;
        RECT 29.075 123.685 29.335 124.165 ;
        RECT 29.515 123.515 29.775 123.970 ;
        RECT 29.945 123.685 30.195 124.165 ;
        RECT 30.375 123.515 30.635 123.970 ;
        RECT 30.805 123.685 31.055 124.165 ;
        RECT 31.235 123.515 31.495 123.970 ;
        RECT 31.665 123.685 31.910 124.165 ;
        RECT 32.080 123.515 32.355 123.970 ;
        RECT 32.525 123.685 32.770 124.165 ;
        RECT 32.940 123.515 33.200 123.970 ;
        RECT 33.370 123.685 33.630 124.165 ;
        RECT 33.800 123.515 34.060 123.970 ;
        RECT 34.230 123.685 34.490 124.165 ;
        RECT 34.660 123.515 34.920 123.970 ;
        RECT 35.090 123.605 35.350 124.165 ;
        RECT 25.260 122.625 25.610 123.275 ;
        RECT 26.245 122.705 26.995 123.225 ;
        RECT 27.165 122.875 27.915 123.395 ;
        RECT 28.175 123.345 34.920 123.515 ;
        RECT 28.175 122.755 29.340 123.345 ;
        RECT 35.520 123.175 35.770 123.985 ;
        RECT 35.950 123.640 36.210 124.165 ;
        RECT 36.380 123.175 36.630 123.985 ;
        RECT 36.810 123.655 37.115 124.165 ;
        RECT 29.510 122.925 36.630 123.175 ;
        RECT 36.800 122.925 37.115 123.485 ;
        RECT 37.285 123.440 37.575 124.165 ;
        RECT 38.205 123.395 39.875 124.165 ;
        RECT 40.050 123.620 45.395 124.165 ;
        RECT 45.570 123.620 50.915 124.165 ;
        RECT 24.860 122.285 25.525 122.455 ;
        RECT 24.855 121.615 25.185 122.115 ;
        RECT 25.355 121.785 25.525 122.285 ;
        RECT 26.245 121.615 27.915 122.705 ;
        RECT 28.175 122.530 34.920 122.755 ;
        RECT 28.175 121.615 28.445 122.360 ;
        RECT 28.615 121.790 28.905 122.530 ;
        RECT 29.515 122.515 34.920 122.530 ;
        RECT 29.075 121.620 29.330 122.345 ;
        RECT 29.515 121.790 29.775 122.515 ;
        RECT 29.945 121.620 30.190 122.345 ;
        RECT 30.375 121.790 30.635 122.515 ;
        RECT 30.805 121.620 31.050 122.345 ;
        RECT 31.235 121.790 31.495 122.515 ;
        RECT 31.665 121.620 31.910 122.345 ;
        RECT 32.080 121.790 32.340 122.515 ;
        RECT 32.510 121.620 32.770 122.345 ;
        RECT 32.940 121.790 33.200 122.515 ;
        RECT 33.370 121.620 33.630 122.345 ;
        RECT 33.800 121.790 34.060 122.515 ;
        RECT 34.230 121.620 34.490 122.345 ;
        RECT 34.660 121.790 34.920 122.515 ;
        RECT 35.090 121.620 35.350 122.415 ;
        RECT 35.520 121.790 35.770 122.925 ;
        RECT 29.075 121.615 35.350 121.620 ;
        RECT 35.950 121.615 36.210 122.425 ;
        RECT 36.385 121.785 36.630 122.925 ;
        RECT 36.810 121.615 37.105 122.425 ;
        RECT 37.285 121.615 37.575 122.780 ;
        RECT 38.205 122.705 38.955 123.225 ;
        RECT 39.125 122.875 39.875 123.395 ;
        RECT 38.205 121.615 39.875 122.705 ;
        RECT 41.640 122.050 41.990 123.300 ;
        RECT 43.470 122.790 43.810 123.620 ;
        RECT 47.160 122.050 47.510 123.300 ;
        RECT 48.990 122.790 49.330 123.620 ;
        RECT 51.360 123.355 51.605 123.960 ;
        RECT 51.825 123.630 52.335 124.165 ;
        RECT 51.085 123.185 52.315 123.355 ;
        RECT 51.085 122.375 51.425 123.185 ;
        RECT 51.595 122.620 52.345 122.810 ;
        RECT 40.050 121.615 45.395 122.050 ;
        RECT 45.570 121.615 50.915 122.050 ;
        RECT 51.085 121.965 51.600 122.375 ;
        RECT 51.835 121.615 52.005 122.375 ;
        RECT 52.175 121.955 52.345 122.620 ;
        RECT 52.515 122.635 52.705 123.995 ;
        RECT 52.875 123.145 53.150 123.995 ;
        RECT 53.340 123.630 53.870 123.995 ;
        RECT 54.295 123.765 54.625 124.165 ;
        RECT 53.695 123.595 53.870 123.630 ;
        RECT 52.875 122.975 53.155 123.145 ;
        RECT 52.875 122.835 53.150 122.975 ;
        RECT 53.355 122.635 53.525 123.435 ;
        RECT 52.515 122.465 53.525 122.635 ;
        RECT 53.695 123.425 54.625 123.595 ;
        RECT 54.795 123.425 55.050 123.995 ;
        RECT 53.695 122.295 53.865 123.425 ;
        RECT 54.455 123.255 54.625 123.425 ;
        RECT 52.740 122.125 53.865 122.295 ;
        RECT 54.035 122.925 54.230 123.255 ;
        RECT 54.455 122.925 54.710 123.255 ;
        RECT 54.035 121.955 54.205 122.925 ;
        RECT 54.880 122.755 55.050 123.425 ;
        RECT 56.295 123.365 56.625 124.165 ;
        RECT 56.795 123.515 56.965 123.995 ;
        RECT 57.135 123.685 57.465 124.165 ;
        RECT 57.635 123.515 57.805 123.995 ;
        RECT 58.055 123.685 58.295 124.165 ;
        RECT 58.475 123.515 58.645 123.995 ;
        RECT 56.795 123.345 57.805 123.515 ;
        RECT 58.010 123.345 58.645 123.515 ;
        RECT 60.035 123.475 60.365 124.165 ;
        RECT 60.825 123.570 61.445 123.995 ;
        RECT 61.615 123.675 61.945 124.165 ;
        RECT 56.795 122.805 57.290 123.345 ;
        RECT 58.010 123.175 58.180 123.345 ;
        RECT 61.085 123.235 61.445 123.570 ;
        RECT 57.680 123.005 58.180 123.175 ;
        RECT 52.175 121.785 54.205 121.955 ;
        RECT 54.375 121.615 54.545 122.755 ;
        RECT 54.715 121.785 55.050 122.755 ;
        RECT 56.295 121.615 56.625 122.765 ;
        RECT 56.795 122.635 57.805 122.805 ;
        RECT 56.795 121.785 56.965 122.635 ;
        RECT 57.135 121.615 57.465 122.415 ;
        RECT 57.635 121.785 57.805 122.635 ;
        RECT 58.010 122.765 58.180 123.005 ;
        RECT 58.350 122.935 58.730 123.175 ;
        RECT 60.025 122.955 61.445 123.235 ;
        RECT 58.010 122.595 58.725 122.765 ;
        RECT 57.985 121.615 58.225 122.415 ;
        RECT 58.395 121.785 58.725 122.595 ;
        RECT 59.495 121.615 59.825 122.785 ;
        RECT 60.025 121.785 60.355 122.955 ;
        RECT 60.555 121.615 60.885 122.785 ;
        RECT 61.085 121.785 61.445 122.955 ;
        RECT 61.615 122.925 61.955 123.505 ;
        RECT 63.045 123.440 63.335 124.165 ;
        RECT 63.780 123.355 64.025 123.960 ;
        RECT 64.245 123.630 64.755 124.165 ;
        RECT 63.505 123.185 64.735 123.355 ;
        RECT 61.615 121.615 61.945 122.755 ;
        RECT 63.045 121.615 63.335 122.780 ;
        RECT 63.505 122.375 63.845 123.185 ;
        RECT 64.015 122.620 64.765 122.810 ;
        RECT 63.505 121.965 64.020 122.375 ;
        RECT 64.255 121.615 64.425 122.375 ;
        RECT 64.595 121.955 64.765 122.620 ;
        RECT 64.935 122.635 65.125 123.995 ;
        RECT 65.295 123.825 65.570 123.995 ;
        RECT 65.295 123.655 65.575 123.825 ;
        RECT 65.295 122.835 65.570 123.655 ;
        RECT 65.760 123.630 66.290 123.995 ;
        RECT 66.715 123.765 67.045 124.165 ;
        RECT 66.115 123.595 66.290 123.630 ;
        RECT 65.775 122.635 65.945 123.435 ;
        RECT 64.935 122.465 65.945 122.635 ;
        RECT 66.115 123.425 67.045 123.595 ;
        RECT 67.215 123.425 67.470 123.995 ;
        RECT 66.115 122.295 66.285 123.425 ;
        RECT 66.875 123.255 67.045 123.425 ;
        RECT 65.160 122.125 66.285 122.295 ;
        RECT 66.455 122.925 66.650 123.255 ;
        RECT 66.875 122.925 67.130 123.255 ;
        RECT 66.455 121.955 66.625 122.925 ;
        RECT 67.300 122.755 67.470 123.425 ;
        RECT 67.645 123.415 68.855 124.165 ;
        RECT 64.595 121.785 66.625 121.955 ;
        RECT 66.795 121.615 66.965 122.755 ;
        RECT 67.135 121.785 67.470 122.755 ;
        RECT 67.645 122.705 68.165 123.245 ;
        RECT 68.335 122.875 68.855 123.415 ;
        RECT 69.025 123.395 72.535 124.165 ;
        RECT 72.710 123.620 78.055 124.165 ;
        RECT 69.025 122.705 70.715 123.225 ;
        RECT 70.885 122.875 72.535 123.395 ;
        RECT 67.645 121.615 68.855 122.705 ;
        RECT 69.025 121.615 72.535 122.705 ;
        RECT 74.300 122.050 74.650 123.300 ;
        RECT 76.130 122.790 76.470 123.620 ;
        RECT 78.500 123.355 78.745 123.960 ;
        RECT 78.965 123.630 79.475 124.165 ;
        RECT 78.225 123.185 79.455 123.355 ;
        RECT 78.225 122.375 78.565 123.185 ;
        RECT 78.735 122.620 79.485 122.810 ;
        RECT 72.710 121.615 78.055 122.050 ;
        RECT 78.225 121.965 78.740 122.375 ;
        RECT 78.975 121.615 79.145 122.375 ;
        RECT 79.315 121.955 79.485 122.620 ;
        RECT 79.655 122.635 79.845 123.995 ;
        RECT 80.015 123.485 80.290 123.995 ;
        RECT 80.480 123.630 81.010 123.995 ;
        RECT 81.435 123.765 81.765 124.165 ;
        RECT 80.835 123.595 81.010 123.630 ;
        RECT 80.015 123.315 80.295 123.485 ;
        RECT 80.015 122.835 80.290 123.315 ;
        RECT 80.495 122.635 80.665 123.435 ;
        RECT 79.655 122.465 80.665 122.635 ;
        RECT 80.835 123.425 81.765 123.595 ;
        RECT 81.935 123.425 82.190 123.995 ;
        RECT 80.835 122.295 81.005 123.425 ;
        RECT 81.595 123.255 81.765 123.425 ;
        RECT 79.880 122.125 81.005 122.295 ;
        RECT 81.175 122.925 81.370 123.255 ;
        RECT 81.595 122.925 81.850 123.255 ;
        RECT 81.175 121.955 81.345 122.925 ;
        RECT 82.020 122.755 82.190 123.425 ;
        RECT 82.640 123.355 82.885 123.960 ;
        RECT 83.105 123.630 83.615 124.165 ;
        RECT 79.315 121.785 81.345 121.955 ;
        RECT 81.515 121.615 81.685 122.755 ;
        RECT 81.855 121.785 82.190 122.755 ;
        RECT 82.365 123.185 83.595 123.355 ;
        RECT 82.365 122.375 82.705 123.185 ;
        RECT 82.875 122.620 83.625 122.810 ;
        RECT 82.365 121.965 82.880 122.375 ;
        RECT 83.115 121.615 83.285 122.375 ;
        RECT 83.455 121.955 83.625 122.620 ;
        RECT 83.795 122.635 83.985 123.995 ;
        RECT 84.155 123.145 84.430 123.995 ;
        RECT 84.620 123.630 85.150 123.995 ;
        RECT 85.575 123.765 85.905 124.165 ;
        RECT 84.975 123.595 85.150 123.630 ;
        RECT 84.155 122.975 84.435 123.145 ;
        RECT 84.155 122.835 84.430 122.975 ;
        RECT 84.635 122.635 84.805 123.435 ;
        RECT 83.795 122.465 84.805 122.635 ;
        RECT 84.975 123.425 85.905 123.595 ;
        RECT 86.075 123.425 86.330 123.995 ;
        RECT 84.975 122.295 85.145 123.425 ;
        RECT 85.735 123.255 85.905 123.425 ;
        RECT 84.020 122.125 85.145 122.295 ;
        RECT 85.315 122.925 85.510 123.255 ;
        RECT 85.735 122.925 85.990 123.255 ;
        RECT 85.315 121.955 85.485 122.925 ;
        RECT 86.160 122.755 86.330 123.425 ;
        RECT 86.965 123.395 88.635 124.165 ;
        RECT 88.805 123.440 89.095 124.165 ;
        RECT 89.265 123.415 90.475 124.165 ;
        RECT 83.455 121.785 85.485 121.955 ;
        RECT 85.655 121.615 85.825 122.755 ;
        RECT 85.995 121.785 86.330 122.755 ;
        RECT 86.965 122.705 87.715 123.225 ;
        RECT 87.885 122.875 88.635 123.395 ;
        RECT 86.965 121.615 88.635 122.705 ;
        RECT 88.805 121.615 89.095 122.780 ;
        RECT 89.265 122.705 89.785 123.245 ;
        RECT 89.955 122.875 90.475 123.415 ;
        RECT 90.685 123.345 90.915 124.165 ;
        RECT 91.085 123.365 91.415 123.995 ;
        RECT 90.665 122.925 90.995 123.175 ;
        RECT 91.165 122.765 91.415 123.365 ;
        RECT 91.585 123.345 91.795 124.165 ;
        RECT 92.300 123.355 92.545 123.960 ;
        RECT 92.765 123.630 93.275 124.165 ;
        RECT 89.265 121.615 90.475 122.705 ;
        RECT 90.685 121.615 90.915 122.755 ;
        RECT 91.085 121.785 91.415 122.765 ;
        RECT 92.025 123.185 93.255 123.355 ;
        RECT 91.585 121.615 91.795 122.755 ;
        RECT 92.025 122.375 92.365 123.185 ;
        RECT 92.535 122.620 93.285 122.810 ;
        RECT 92.025 121.965 92.540 122.375 ;
        RECT 92.775 121.615 92.945 122.375 ;
        RECT 93.115 121.955 93.285 122.620 ;
        RECT 93.455 122.635 93.645 123.995 ;
        RECT 93.815 123.825 94.090 123.995 ;
        RECT 93.815 123.655 94.095 123.825 ;
        RECT 93.815 122.835 94.090 123.655 ;
        RECT 94.280 123.630 94.810 123.995 ;
        RECT 95.235 123.765 95.565 124.165 ;
        RECT 94.635 123.595 94.810 123.630 ;
        RECT 94.295 122.635 94.465 123.435 ;
        RECT 93.455 122.465 94.465 122.635 ;
        RECT 94.635 123.425 95.565 123.595 ;
        RECT 95.735 123.425 95.990 123.995 ;
        RECT 94.635 122.295 94.805 123.425 ;
        RECT 95.395 123.255 95.565 123.425 ;
        RECT 93.680 122.125 94.805 122.295 ;
        RECT 94.975 122.925 95.170 123.255 ;
        RECT 95.395 122.925 95.650 123.255 ;
        RECT 94.975 121.955 95.145 122.925 ;
        RECT 95.820 122.755 95.990 123.425 ;
        RECT 96.540 123.455 96.795 123.985 ;
        RECT 96.975 123.705 97.260 124.165 ;
        RECT 96.540 123.145 96.720 123.455 ;
        RECT 97.440 123.255 97.690 123.905 ;
        RECT 96.455 122.975 96.720 123.145 ;
        RECT 93.115 121.785 95.145 121.955 ;
        RECT 95.315 121.615 95.485 122.755 ;
        RECT 95.655 121.785 95.990 122.755 ;
        RECT 96.540 122.595 96.720 122.975 ;
        RECT 96.890 122.925 97.690 123.255 ;
        RECT 96.540 121.925 96.795 122.595 ;
        RECT 96.975 121.615 97.260 122.415 ;
        RECT 97.440 122.335 97.690 122.925 ;
        RECT 97.890 123.570 98.210 123.900 ;
        RECT 98.390 123.685 99.050 124.165 ;
        RECT 99.250 123.775 100.100 123.945 ;
        RECT 97.890 122.675 98.080 123.570 ;
        RECT 98.400 123.245 99.060 123.515 ;
        RECT 98.730 123.185 99.060 123.245 ;
        RECT 98.250 123.015 98.580 123.075 ;
        RECT 99.250 123.015 99.420 123.775 ;
        RECT 100.660 123.705 100.980 124.165 ;
        RECT 101.180 123.525 101.430 123.955 ;
        RECT 101.720 123.725 102.130 124.165 ;
        RECT 102.300 123.785 103.315 123.985 ;
        RECT 99.590 123.355 100.840 123.525 ;
        RECT 99.590 123.235 99.920 123.355 ;
        RECT 98.250 122.845 100.150 123.015 ;
        RECT 97.890 122.505 99.810 122.675 ;
        RECT 97.890 122.485 98.210 122.505 ;
        RECT 97.440 121.825 97.770 122.335 ;
        RECT 98.040 121.875 98.210 122.485 ;
        RECT 99.980 122.335 100.150 122.845 ;
        RECT 100.320 122.775 100.500 123.185 ;
        RECT 100.670 122.595 100.840 123.355 ;
        RECT 98.380 121.615 98.710 122.305 ;
        RECT 98.940 122.165 100.150 122.335 ;
        RECT 100.320 122.285 100.840 122.595 ;
        RECT 101.010 123.185 101.430 123.525 ;
        RECT 101.720 123.185 102.130 123.515 ;
        RECT 101.010 122.415 101.200 123.185 ;
        RECT 102.300 123.055 102.470 123.785 ;
        RECT 103.615 123.615 103.785 123.945 ;
        RECT 103.955 123.785 104.285 124.165 ;
        RECT 102.640 123.235 102.990 123.605 ;
        RECT 102.300 123.015 102.720 123.055 ;
        RECT 101.370 122.845 102.720 123.015 ;
        RECT 101.370 122.685 101.620 122.845 ;
        RECT 102.130 122.415 102.380 122.675 ;
        RECT 101.010 122.165 102.380 122.415 ;
        RECT 98.940 121.875 99.180 122.165 ;
        RECT 99.980 122.085 100.150 122.165 ;
        RECT 99.380 121.615 99.800 121.995 ;
        RECT 99.980 121.835 100.610 122.085 ;
        RECT 101.080 121.615 101.410 121.995 ;
        RECT 101.580 121.875 101.750 122.165 ;
        RECT 102.550 122.000 102.720 122.845 ;
        RECT 103.170 122.675 103.390 123.545 ;
        RECT 103.615 123.425 104.310 123.615 ;
        RECT 102.890 122.295 103.390 122.675 ;
        RECT 103.560 122.625 103.970 123.245 ;
        RECT 104.140 122.455 104.310 123.425 ;
        RECT 103.615 122.285 104.310 122.455 ;
        RECT 101.930 121.615 102.310 121.995 ;
        RECT 102.550 121.830 103.380 122.000 ;
        RECT 103.615 121.785 103.785 122.285 ;
        RECT 103.955 121.615 104.285 122.115 ;
        RECT 104.500 121.785 104.725 123.905 ;
        RECT 104.895 123.785 105.225 124.165 ;
        RECT 105.395 123.615 105.565 123.905 ;
        RECT 104.900 123.445 105.565 123.615 ;
        RECT 104.900 122.455 105.130 123.445 ;
        RECT 105.830 123.425 106.085 123.995 ;
        RECT 106.255 123.765 106.585 124.165 ;
        RECT 107.010 123.630 107.540 123.995 ;
        RECT 107.730 123.825 108.005 123.995 ;
        RECT 107.725 123.655 108.005 123.825 ;
        RECT 107.010 123.595 107.185 123.630 ;
        RECT 106.255 123.425 107.185 123.595 ;
        RECT 105.300 122.625 105.650 123.275 ;
        RECT 105.830 122.755 106.000 123.425 ;
        RECT 106.255 123.255 106.425 123.425 ;
        RECT 106.170 122.925 106.425 123.255 ;
        RECT 106.650 122.925 106.845 123.255 ;
        RECT 104.900 122.285 105.565 122.455 ;
        RECT 104.895 121.615 105.225 122.115 ;
        RECT 105.395 121.785 105.565 122.285 ;
        RECT 105.830 121.785 106.165 122.755 ;
        RECT 106.335 121.615 106.505 122.755 ;
        RECT 106.675 121.955 106.845 122.925 ;
        RECT 107.015 122.295 107.185 123.425 ;
        RECT 107.355 122.635 107.525 123.435 ;
        RECT 107.730 122.835 108.005 123.655 ;
        RECT 108.175 122.635 108.365 123.995 ;
        RECT 108.545 123.630 109.055 124.165 ;
        RECT 109.275 123.355 109.520 123.960 ;
        RECT 110.890 123.695 111.220 124.165 ;
        RECT 111.390 123.525 111.615 123.970 ;
        RECT 111.785 123.640 112.080 124.165 ;
        RECT 110.885 123.355 111.615 123.525 ;
        RECT 112.725 123.395 114.395 124.165 ;
        RECT 114.565 123.440 114.855 124.165 ;
        RECT 108.565 123.185 109.795 123.355 ;
        RECT 107.355 122.465 108.365 122.635 ;
        RECT 108.535 122.620 109.285 122.810 ;
        RECT 107.015 122.125 108.140 122.295 ;
        RECT 108.535 121.955 108.705 122.620 ;
        RECT 109.455 122.375 109.795 123.185 ;
        RECT 110.885 122.790 111.165 123.355 ;
        RECT 111.335 122.960 112.555 123.185 ;
        RECT 110.885 122.620 112.485 122.790 ;
        RECT 106.675 121.785 108.705 121.955 ;
        RECT 108.875 121.615 109.045 122.375 ;
        RECT 109.280 121.965 109.795 122.375 ;
        RECT 110.945 121.615 111.200 122.450 ;
        RECT 111.370 121.815 111.630 122.620 ;
        RECT 111.800 121.615 112.060 122.450 ;
        RECT 112.230 121.815 112.485 122.620 ;
        RECT 112.725 122.705 113.475 123.225 ;
        RECT 113.645 122.875 114.395 123.395 ;
        RECT 115.760 123.355 116.005 123.960 ;
        RECT 116.225 123.630 116.735 124.165 ;
        RECT 115.485 123.185 116.715 123.355 ;
        RECT 112.725 121.615 114.395 122.705 ;
        RECT 114.565 121.615 114.855 122.780 ;
        RECT 115.485 122.375 115.825 123.185 ;
        RECT 115.995 122.620 116.745 122.810 ;
        RECT 115.485 121.965 116.000 122.375 ;
        RECT 116.235 121.615 116.405 122.375 ;
        RECT 116.575 121.955 116.745 122.620 ;
        RECT 116.915 122.635 117.105 123.995 ;
        RECT 117.275 123.825 117.550 123.995 ;
        RECT 117.275 123.655 117.555 123.825 ;
        RECT 117.275 122.835 117.550 123.655 ;
        RECT 117.740 123.630 118.270 123.995 ;
        RECT 118.695 123.765 119.025 124.165 ;
        RECT 118.095 123.595 118.270 123.630 ;
        RECT 117.755 122.635 117.925 123.435 ;
        RECT 116.915 122.465 117.925 122.635 ;
        RECT 118.095 123.425 119.025 123.595 ;
        RECT 119.195 123.425 119.450 123.995 ;
        RECT 118.095 122.295 118.265 123.425 ;
        RECT 118.855 123.255 119.025 123.425 ;
        RECT 117.140 122.125 118.265 122.295 ;
        RECT 118.435 122.925 118.630 123.255 ;
        RECT 118.855 122.925 119.110 123.255 ;
        RECT 118.435 121.955 118.605 122.925 ;
        RECT 119.280 122.755 119.450 123.425 ;
        RECT 119.625 123.415 120.835 124.165 ;
        RECT 121.095 123.615 121.265 123.995 ;
        RECT 121.445 123.785 121.775 124.165 ;
        RECT 121.095 123.445 121.760 123.615 ;
        RECT 121.955 123.490 122.215 123.995 ;
        RECT 116.575 121.785 118.605 121.955 ;
        RECT 118.775 121.615 118.945 122.755 ;
        RECT 119.115 121.785 119.450 122.755 ;
        RECT 119.625 122.705 120.145 123.245 ;
        RECT 120.315 122.875 120.835 123.415 ;
        RECT 121.025 122.895 121.355 123.265 ;
        RECT 121.590 123.190 121.760 123.445 ;
        RECT 121.590 122.860 121.875 123.190 ;
        RECT 121.590 122.715 121.760 122.860 ;
        RECT 119.625 121.615 120.835 122.705 ;
        RECT 121.095 122.545 121.760 122.715 ;
        RECT 122.045 122.690 122.215 123.490 ;
        RECT 122.845 123.395 126.355 124.165 ;
        RECT 126.525 123.415 127.735 124.165 ;
        RECT 121.095 121.785 121.265 122.545 ;
        RECT 121.445 121.615 121.775 122.375 ;
        RECT 121.945 121.785 122.215 122.690 ;
        RECT 122.845 122.705 124.535 123.225 ;
        RECT 124.705 122.875 126.355 123.395 ;
        RECT 126.525 122.705 127.045 123.245 ;
        RECT 127.215 122.875 127.735 123.415 ;
        RECT 122.845 121.615 126.355 122.705 ;
        RECT 126.525 121.615 127.735 122.705 ;
        RECT 14.660 121.445 127.820 121.615 ;
        RECT 14.745 120.355 15.955 121.445 ;
        RECT 14.745 119.645 15.265 120.185 ;
        RECT 15.435 119.815 15.955 120.355 ;
        RECT 16.585 120.355 19.175 121.445 ;
        RECT 16.585 119.835 17.795 120.355 ;
        RECT 19.405 120.305 19.615 121.445 ;
        RECT 19.785 120.295 20.115 121.275 ;
        RECT 20.285 120.305 20.515 121.445 ;
        RECT 21.185 120.355 22.855 121.445 ;
        RECT 23.115 120.515 23.285 121.275 ;
        RECT 23.465 120.685 23.795 121.445 ;
        RECT 17.965 119.665 19.175 120.185 ;
        RECT 14.745 118.895 15.955 119.645 ;
        RECT 16.585 118.895 19.175 119.665 ;
        RECT 19.405 118.895 19.615 119.715 ;
        RECT 19.785 119.695 20.035 120.295 ;
        RECT 20.205 119.885 20.535 120.135 ;
        RECT 21.185 119.835 21.935 120.355 ;
        RECT 23.115 120.345 23.780 120.515 ;
        RECT 23.965 120.370 24.235 121.275 ;
        RECT 23.610 120.200 23.780 120.345 ;
        RECT 19.785 119.065 20.115 119.695 ;
        RECT 20.285 118.895 20.515 119.715 ;
        RECT 22.105 119.665 22.855 120.185 ;
        RECT 23.045 119.795 23.375 120.165 ;
        RECT 23.610 119.870 23.895 120.200 ;
        RECT 21.185 118.895 22.855 119.665 ;
        RECT 23.610 119.615 23.780 119.870 ;
        RECT 23.115 119.445 23.780 119.615 ;
        RECT 24.065 119.570 24.235 120.370 ;
        RECT 24.405 120.280 24.695 121.445 ;
        RECT 24.955 120.775 25.125 121.275 ;
        RECT 25.295 120.945 25.625 121.445 ;
        RECT 24.955 120.605 25.620 120.775 ;
        RECT 24.870 119.785 25.220 120.435 ;
        RECT 23.115 119.065 23.285 119.445 ;
        RECT 23.465 118.895 23.795 119.275 ;
        RECT 23.975 119.065 24.235 119.570 ;
        RECT 24.405 118.895 24.695 119.620 ;
        RECT 25.390 119.615 25.620 120.605 ;
        RECT 24.955 119.445 25.620 119.615 ;
        RECT 24.955 119.155 25.125 119.445 ;
        RECT 25.295 118.895 25.625 119.275 ;
        RECT 25.795 119.155 26.020 121.275 ;
        RECT 26.235 120.945 26.565 121.445 ;
        RECT 26.735 120.775 26.905 121.275 ;
        RECT 27.140 121.060 27.970 121.230 ;
        RECT 28.210 121.065 28.590 121.445 ;
        RECT 26.210 120.605 26.905 120.775 ;
        RECT 26.210 119.635 26.380 120.605 ;
        RECT 26.550 119.815 26.960 120.435 ;
        RECT 27.130 120.385 27.630 120.765 ;
        RECT 26.210 119.445 26.905 119.635 ;
        RECT 27.130 119.515 27.350 120.385 ;
        RECT 27.800 120.215 27.970 121.060 ;
        RECT 28.770 120.895 28.940 121.185 ;
        RECT 29.110 121.065 29.440 121.445 ;
        RECT 29.910 120.975 30.540 121.225 ;
        RECT 30.720 121.065 31.140 121.445 ;
        RECT 30.370 120.895 30.540 120.975 ;
        RECT 31.340 120.895 31.580 121.185 ;
        RECT 28.140 120.645 29.510 120.895 ;
        RECT 28.140 120.385 28.390 120.645 ;
        RECT 28.900 120.215 29.150 120.375 ;
        RECT 27.800 120.045 29.150 120.215 ;
        RECT 27.800 120.005 28.220 120.045 ;
        RECT 27.530 119.455 27.880 119.825 ;
        RECT 26.235 118.895 26.565 119.275 ;
        RECT 26.735 119.115 26.905 119.445 ;
        RECT 28.050 119.275 28.220 120.005 ;
        RECT 29.320 119.875 29.510 120.645 ;
        RECT 28.390 119.545 28.800 119.875 ;
        RECT 29.090 119.535 29.510 119.875 ;
        RECT 29.680 120.465 30.200 120.775 ;
        RECT 30.370 120.725 31.580 120.895 ;
        RECT 31.810 120.755 32.140 121.445 ;
        RECT 29.680 119.705 29.850 120.465 ;
        RECT 30.020 119.875 30.200 120.285 ;
        RECT 30.370 120.215 30.540 120.725 ;
        RECT 32.310 120.575 32.480 121.185 ;
        RECT 32.750 120.725 33.080 121.235 ;
        RECT 32.310 120.555 32.630 120.575 ;
        RECT 30.710 120.385 32.630 120.555 ;
        RECT 30.370 120.045 32.270 120.215 ;
        RECT 30.600 119.705 30.930 119.825 ;
        RECT 29.680 119.535 30.930 119.705 ;
        RECT 27.205 119.075 28.220 119.275 ;
        RECT 28.390 118.895 28.800 119.335 ;
        RECT 29.090 119.105 29.340 119.535 ;
        RECT 29.540 118.895 29.860 119.355 ;
        RECT 31.100 119.285 31.270 120.045 ;
        RECT 31.940 119.985 32.270 120.045 ;
        RECT 31.460 119.815 31.790 119.875 ;
        RECT 31.460 119.545 32.120 119.815 ;
        RECT 32.440 119.490 32.630 120.385 ;
        RECT 30.420 119.115 31.270 119.285 ;
        RECT 31.470 118.895 32.130 119.375 ;
        RECT 32.310 119.160 32.630 119.490 ;
        RECT 32.830 120.135 33.080 120.725 ;
        RECT 33.260 120.645 33.545 121.445 ;
        RECT 33.725 120.465 33.980 121.135 ;
        RECT 33.800 120.425 33.980 120.465 ;
        RECT 33.800 120.255 34.065 120.425 ;
        RECT 34.565 120.305 34.795 121.445 ;
        RECT 34.965 120.295 35.295 121.275 ;
        RECT 35.465 120.305 35.675 121.445 ;
        RECT 36.280 121.105 36.535 121.135 ;
        RECT 36.195 120.935 36.535 121.105 ;
        RECT 36.280 120.465 36.535 120.935 ;
        RECT 36.715 120.645 37.000 121.445 ;
        RECT 37.180 120.725 37.510 121.235 ;
        RECT 32.830 119.805 33.630 120.135 ;
        RECT 32.830 119.155 33.080 119.805 ;
        RECT 33.800 119.605 33.980 120.255 ;
        RECT 34.545 119.885 34.875 120.135 ;
        RECT 33.260 118.895 33.545 119.355 ;
        RECT 33.725 119.075 33.980 119.605 ;
        RECT 34.565 118.895 34.795 119.715 ;
        RECT 35.045 119.695 35.295 120.295 ;
        RECT 34.965 119.065 35.295 119.695 ;
        RECT 35.465 118.895 35.675 119.715 ;
        RECT 36.280 119.605 36.460 120.465 ;
        RECT 37.180 120.135 37.430 120.725 ;
        RECT 37.780 120.575 37.950 121.185 ;
        RECT 38.120 120.755 38.450 121.445 ;
        RECT 38.680 120.895 38.920 121.185 ;
        RECT 39.120 121.065 39.540 121.445 ;
        RECT 39.720 120.975 40.350 121.225 ;
        RECT 40.820 121.065 41.150 121.445 ;
        RECT 39.720 120.895 39.890 120.975 ;
        RECT 41.320 120.895 41.490 121.185 ;
        RECT 41.670 121.065 42.050 121.445 ;
        RECT 42.290 121.060 43.120 121.230 ;
        RECT 38.680 120.725 39.890 120.895 ;
        RECT 36.630 119.805 37.430 120.135 ;
        RECT 36.280 119.075 36.535 119.605 ;
        RECT 36.715 118.895 37.000 119.355 ;
        RECT 37.180 119.155 37.430 119.805 ;
        RECT 37.630 120.555 37.950 120.575 ;
        RECT 37.630 120.385 39.550 120.555 ;
        RECT 37.630 119.490 37.820 120.385 ;
        RECT 39.720 120.215 39.890 120.725 ;
        RECT 40.060 120.465 40.580 120.775 ;
        RECT 37.990 120.045 39.890 120.215 ;
        RECT 37.990 119.985 38.320 120.045 ;
        RECT 38.470 119.815 38.800 119.875 ;
        RECT 38.140 119.545 38.800 119.815 ;
        RECT 37.630 119.160 37.950 119.490 ;
        RECT 38.130 118.895 38.790 119.375 ;
        RECT 38.990 119.285 39.160 120.045 ;
        RECT 40.060 119.875 40.240 120.285 ;
        RECT 39.330 119.705 39.660 119.825 ;
        RECT 40.410 119.705 40.580 120.465 ;
        RECT 39.330 119.535 40.580 119.705 ;
        RECT 40.750 120.645 42.120 120.895 ;
        RECT 40.750 119.875 40.940 120.645 ;
        RECT 41.870 120.385 42.120 120.645 ;
        RECT 41.110 120.215 41.360 120.375 ;
        RECT 42.290 120.215 42.460 121.060 ;
        RECT 43.355 120.775 43.525 121.275 ;
        RECT 43.695 120.945 44.025 121.445 ;
        RECT 42.630 120.385 43.130 120.765 ;
        RECT 43.355 120.605 44.050 120.775 ;
        RECT 41.110 120.045 42.460 120.215 ;
        RECT 42.040 120.005 42.460 120.045 ;
        RECT 40.750 119.535 41.170 119.875 ;
        RECT 41.460 119.545 41.870 119.875 ;
        RECT 38.990 119.115 39.840 119.285 ;
        RECT 40.400 118.895 40.720 119.355 ;
        RECT 40.920 119.105 41.170 119.535 ;
        RECT 41.460 118.895 41.870 119.335 ;
        RECT 42.040 119.275 42.210 120.005 ;
        RECT 42.380 119.455 42.730 119.825 ;
        RECT 42.910 119.515 43.130 120.385 ;
        RECT 43.300 119.815 43.710 120.435 ;
        RECT 43.880 119.635 44.050 120.605 ;
        RECT 43.355 119.445 44.050 119.635 ;
        RECT 42.040 119.075 43.055 119.275 ;
        RECT 43.355 119.115 43.525 119.445 ;
        RECT 43.695 118.895 44.025 119.275 ;
        RECT 44.240 119.155 44.465 121.275 ;
        RECT 44.635 120.945 44.965 121.445 ;
        RECT 45.135 120.775 45.305 121.275 ;
        RECT 44.640 120.605 45.305 120.775 ;
        RECT 46.025 120.685 46.540 121.095 ;
        RECT 46.775 120.685 46.945 121.445 ;
        RECT 47.115 121.105 49.145 121.275 ;
        RECT 44.640 119.615 44.870 120.605 ;
        RECT 45.040 119.785 45.390 120.435 ;
        RECT 46.025 119.875 46.365 120.685 ;
        RECT 47.115 120.440 47.285 121.105 ;
        RECT 47.680 120.765 48.805 120.935 ;
        RECT 46.535 120.250 47.285 120.440 ;
        RECT 47.455 120.425 48.465 120.595 ;
        RECT 46.025 119.705 47.255 119.875 ;
        RECT 44.640 119.445 45.305 119.615 ;
        RECT 44.635 118.895 44.965 119.275 ;
        RECT 45.135 119.155 45.305 119.445 ;
        RECT 46.300 119.100 46.545 119.705 ;
        RECT 46.765 118.895 47.275 119.430 ;
        RECT 47.455 119.065 47.645 120.425 ;
        RECT 47.815 119.405 48.090 120.225 ;
        RECT 48.295 119.625 48.465 120.425 ;
        RECT 48.635 119.635 48.805 120.765 ;
        RECT 48.975 120.135 49.145 121.105 ;
        RECT 49.315 120.305 49.485 121.445 ;
        RECT 49.655 120.305 49.990 121.275 ;
        RECT 48.975 119.805 49.170 120.135 ;
        RECT 49.395 119.805 49.650 120.135 ;
        RECT 49.395 119.635 49.565 119.805 ;
        RECT 49.820 119.635 49.990 120.305 ;
        RECT 50.165 120.280 50.455 121.445 ;
        RECT 51.085 120.355 52.755 121.445 ;
        RECT 52.935 120.635 53.230 121.445 ;
        RECT 51.085 119.835 51.835 120.355 ;
        RECT 52.005 119.665 52.755 120.185 ;
        RECT 53.410 120.135 53.655 121.275 ;
        RECT 53.830 120.635 54.090 121.445 ;
        RECT 54.690 121.440 60.965 121.445 ;
        RECT 54.270 120.135 54.520 121.270 ;
        RECT 54.690 120.645 54.950 121.440 ;
        RECT 55.120 120.545 55.380 121.270 ;
        RECT 55.550 120.715 55.810 121.440 ;
        RECT 55.980 120.545 56.240 121.270 ;
        RECT 56.410 120.715 56.670 121.440 ;
        RECT 56.840 120.545 57.100 121.270 ;
        RECT 57.270 120.715 57.530 121.440 ;
        RECT 57.700 120.545 57.960 121.270 ;
        RECT 58.130 120.715 58.375 121.440 ;
        RECT 58.545 120.545 58.805 121.270 ;
        RECT 58.990 120.715 59.235 121.440 ;
        RECT 59.405 120.545 59.665 121.270 ;
        RECT 59.850 120.715 60.095 121.440 ;
        RECT 60.265 120.545 60.525 121.270 ;
        RECT 60.710 120.715 60.965 121.440 ;
        RECT 55.120 120.530 60.525 120.545 ;
        RECT 61.135 120.530 61.425 121.270 ;
        RECT 61.595 120.700 61.865 121.445 ;
        RECT 55.120 120.305 61.865 120.530 ;
        RECT 48.635 119.465 49.565 119.635 ;
        RECT 48.635 119.430 48.810 119.465 ;
        RECT 47.815 119.235 48.095 119.405 ;
        RECT 47.815 119.065 48.090 119.235 ;
        RECT 48.280 119.065 48.810 119.430 ;
        RECT 49.235 118.895 49.565 119.295 ;
        RECT 49.735 119.065 49.990 119.635 ;
        RECT 50.165 118.895 50.455 119.620 ;
        RECT 51.085 118.895 52.755 119.665 ;
        RECT 52.925 119.575 53.240 120.135 ;
        RECT 53.410 119.885 60.530 120.135 ;
        RECT 52.925 118.895 53.230 119.405 ;
        RECT 53.410 119.075 53.660 119.885 ;
        RECT 53.830 118.895 54.090 119.420 ;
        RECT 54.270 119.075 54.520 119.885 ;
        RECT 60.700 119.715 61.865 120.305 ;
        RECT 62.125 120.355 63.335 121.445 ;
        RECT 63.505 120.685 64.020 121.095 ;
        RECT 64.255 120.685 64.425 121.445 ;
        RECT 64.595 121.105 66.625 121.275 ;
        RECT 62.125 119.815 62.645 120.355 ;
        RECT 55.120 119.545 61.865 119.715 ;
        RECT 62.815 119.645 63.335 120.185 ;
        RECT 63.505 119.875 63.845 120.685 ;
        RECT 64.595 120.440 64.765 121.105 ;
        RECT 65.160 120.765 66.285 120.935 ;
        RECT 64.015 120.250 64.765 120.440 ;
        RECT 64.935 120.425 65.945 120.595 ;
        RECT 63.505 119.705 64.735 119.875 ;
        RECT 54.690 118.895 54.950 119.455 ;
        RECT 55.120 119.090 55.380 119.545 ;
        RECT 55.550 118.895 55.810 119.375 ;
        RECT 55.980 119.090 56.240 119.545 ;
        RECT 56.410 118.895 56.670 119.375 ;
        RECT 56.840 119.090 57.100 119.545 ;
        RECT 57.270 118.895 57.515 119.375 ;
        RECT 57.685 119.090 57.960 119.545 ;
        RECT 58.130 118.895 58.375 119.375 ;
        RECT 58.545 119.090 58.805 119.545 ;
        RECT 58.985 118.895 59.235 119.375 ;
        RECT 59.405 119.090 59.665 119.545 ;
        RECT 59.845 118.895 60.095 119.375 ;
        RECT 60.265 119.090 60.525 119.545 ;
        RECT 60.705 118.895 60.965 119.375 ;
        RECT 61.135 119.090 61.395 119.545 ;
        RECT 61.565 118.895 61.865 119.375 ;
        RECT 62.125 118.895 63.335 119.645 ;
        RECT 63.780 119.100 64.025 119.705 ;
        RECT 64.245 118.895 64.755 119.430 ;
        RECT 64.935 119.065 65.125 120.425 ;
        RECT 65.295 120.085 65.570 120.225 ;
        RECT 65.295 119.915 65.575 120.085 ;
        RECT 65.295 119.065 65.570 119.915 ;
        RECT 65.775 119.625 65.945 120.425 ;
        RECT 66.115 119.635 66.285 120.765 ;
        RECT 66.455 120.135 66.625 121.105 ;
        RECT 66.795 120.305 66.965 121.445 ;
        RECT 67.135 120.305 67.470 121.275 ;
        RECT 68.195 120.515 68.365 121.275 ;
        RECT 68.545 120.685 68.875 121.445 ;
        RECT 68.195 120.345 68.860 120.515 ;
        RECT 69.045 120.370 69.315 121.275 ;
        RECT 70.410 121.010 75.755 121.445 ;
        RECT 66.455 119.805 66.650 120.135 ;
        RECT 66.875 119.805 67.130 120.135 ;
        RECT 66.875 119.635 67.045 119.805 ;
        RECT 67.300 119.635 67.470 120.305 ;
        RECT 68.690 120.200 68.860 120.345 ;
        RECT 68.125 119.795 68.455 120.165 ;
        RECT 68.690 119.870 68.975 120.200 ;
        RECT 66.115 119.465 67.045 119.635 ;
        RECT 66.115 119.430 66.290 119.465 ;
        RECT 65.760 119.065 66.290 119.430 ;
        RECT 66.715 118.895 67.045 119.295 ;
        RECT 67.215 119.065 67.470 119.635 ;
        RECT 68.690 119.615 68.860 119.870 ;
        RECT 68.195 119.445 68.860 119.615 ;
        RECT 69.145 119.570 69.315 120.370 ;
        RECT 72.000 119.760 72.350 121.010 ;
        RECT 75.925 120.280 76.215 121.445 ;
        RECT 76.885 120.305 77.115 121.445 ;
        RECT 77.285 120.295 77.615 121.275 ;
        RECT 77.785 120.305 77.995 121.445 ;
        RECT 78.600 121.105 78.855 121.135 ;
        RECT 78.515 120.935 78.855 121.105 ;
        RECT 78.600 120.465 78.855 120.935 ;
        RECT 79.035 120.645 79.320 121.445 ;
        RECT 79.500 120.725 79.830 121.235 ;
        RECT 68.195 119.065 68.365 119.445 ;
        RECT 68.545 118.895 68.875 119.275 ;
        RECT 69.055 119.065 69.315 119.570 ;
        RECT 73.830 119.440 74.170 120.270 ;
        RECT 76.865 119.885 77.195 120.135 ;
        RECT 70.410 118.895 75.755 119.440 ;
        RECT 75.925 118.895 76.215 119.620 ;
        RECT 76.885 118.895 77.115 119.715 ;
        RECT 77.365 119.695 77.615 120.295 ;
        RECT 77.285 119.065 77.615 119.695 ;
        RECT 77.785 118.895 77.995 119.715 ;
        RECT 78.600 119.605 78.780 120.465 ;
        RECT 79.500 120.135 79.750 120.725 ;
        RECT 80.100 120.575 80.270 121.185 ;
        RECT 80.440 120.755 80.770 121.445 ;
        RECT 81.000 120.895 81.240 121.185 ;
        RECT 81.440 121.065 81.860 121.445 ;
        RECT 82.040 120.975 82.670 121.225 ;
        RECT 83.140 121.065 83.470 121.445 ;
        RECT 82.040 120.895 82.210 120.975 ;
        RECT 83.640 120.895 83.810 121.185 ;
        RECT 83.990 121.065 84.370 121.445 ;
        RECT 84.610 121.060 85.440 121.230 ;
        RECT 81.000 120.725 82.210 120.895 ;
        RECT 78.950 119.805 79.750 120.135 ;
        RECT 78.600 119.075 78.855 119.605 ;
        RECT 79.035 118.895 79.320 119.355 ;
        RECT 79.500 119.155 79.750 119.805 ;
        RECT 79.950 120.555 80.270 120.575 ;
        RECT 79.950 120.385 81.870 120.555 ;
        RECT 79.950 119.490 80.140 120.385 ;
        RECT 82.040 120.215 82.210 120.725 ;
        RECT 82.380 120.465 82.900 120.775 ;
        RECT 80.310 120.045 82.210 120.215 ;
        RECT 80.310 119.985 80.640 120.045 ;
        RECT 80.790 119.815 81.120 119.875 ;
        RECT 80.460 119.545 81.120 119.815 ;
        RECT 79.950 119.160 80.270 119.490 ;
        RECT 80.450 118.895 81.110 119.375 ;
        RECT 81.310 119.285 81.480 120.045 ;
        RECT 82.380 119.875 82.560 120.285 ;
        RECT 81.650 119.705 81.980 119.825 ;
        RECT 82.730 119.705 82.900 120.465 ;
        RECT 81.650 119.535 82.900 119.705 ;
        RECT 83.070 120.645 84.440 120.895 ;
        RECT 83.070 119.875 83.260 120.645 ;
        RECT 84.190 120.385 84.440 120.645 ;
        RECT 83.430 120.215 83.680 120.375 ;
        RECT 84.610 120.215 84.780 121.060 ;
        RECT 85.675 120.775 85.845 121.275 ;
        RECT 86.015 120.945 86.345 121.445 ;
        RECT 84.950 120.385 85.450 120.765 ;
        RECT 85.675 120.605 86.370 120.775 ;
        RECT 83.430 120.045 84.780 120.215 ;
        RECT 84.360 120.005 84.780 120.045 ;
        RECT 83.070 119.535 83.490 119.875 ;
        RECT 83.780 119.545 84.190 119.875 ;
        RECT 81.310 119.115 82.160 119.285 ;
        RECT 82.720 118.895 83.040 119.355 ;
        RECT 83.240 119.105 83.490 119.535 ;
        RECT 83.780 118.895 84.190 119.335 ;
        RECT 84.360 119.275 84.530 120.005 ;
        RECT 84.700 119.455 85.050 119.825 ;
        RECT 85.230 119.515 85.450 120.385 ;
        RECT 85.620 119.815 86.030 120.435 ;
        RECT 86.200 119.635 86.370 120.605 ;
        RECT 85.675 119.445 86.370 119.635 ;
        RECT 84.360 119.075 85.375 119.275 ;
        RECT 85.675 119.115 85.845 119.445 ;
        RECT 86.015 118.895 86.345 119.275 ;
        RECT 86.560 119.155 86.785 121.275 ;
        RECT 86.955 120.945 87.285 121.445 ;
        RECT 87.455 120.775 87.625 121.275 ;
        RECT 86.960 120.605 87.625 120.775 ;
        RECT 86.960 119.615 87.190 120.605 ;
        RECT 87.360 119.785 87.710 120.435 ;
        RECT 87.885 120.370 88.155 121.275 ;
        RECT 88.325 120.685 88.655 121.445 ;
        RECT 88.835 120.515 89.005 121.275 ;
        RECT 90.100 121.105 90.355 121.135 ;
        RECT 90.015 120.935 90.355 121.105 ;
        RECT 86.960 119.445 87.625 119.615 ;
        RECT 86.955 118.895 87.285 119.275 ;
        RECT 87.455 119.155 87.625 119.445 ;
        RECT 87.885 119.570 88.055 120.370 ;
        RECT 88.340 120.345 89.005 120.515 ;
        RECT 90.100 120.465 90.355 120.935 ;
        RECT 90.535 120.645 90.820 121.445 ;
        RECT 91.000 120.725 91.330 121.235 ;
        RECT 88.340 120.200 88.510 120.345 ;
        RECT 88.225 119.870 88.510 120.200 ;
        RECT 88.340 119.615 88.510 119.870 ;
        RECT 88.745 119.795 89.075 120.165 ;
        RECT 87.885 119.065 88.145 119.570 ;
        RECT 88.340 119.445 89.005 119.615 ;
        RECT 88.325 118.895 88.655 119.275 ;
        RECT 88.835 119.065 89.005 119.445 ;
        RECT 90.100 119.605 90.280 120.465 ;
        RECT 91.000 120.135 91.250 120.725 ;
        RECT 91.600 120.575 91.770 121.185 ;
        RECT 91.940 120.755 92.270 121.445 ;
        RECT 92.500 120.895 92.740 121.185 ;
        RECT 92.940 121.065 93.360 121.445 ;
        RECT 93.540 120.975 94.170 121.225 ;
        RECT 94.640 121.065 94.970 121.445 ;
        RECT 93.540 120.895 93.710 120.975 ;
        RECT 95.140 120.895 95.310 121.185 ;
        RECT 95.490 121.065 95.870 121.445 ;
        RECT 96.110 121.060 96.940 121.230 ;
        RECT 92.500 120.725 93.710 120.895 ;
        RECT 90.450 119.805 91.250 120.135 ;
        RECT 90.100 119.075 90.355 119.605 ;
        RECT 90.535 118.895 90.820 119.355 ;
        RECT 91.000 119.155 91.250 119.805 ;
        RECT 91.450 120.555 91.770 120.575 ;
        RECT 91.450 120.385 93.370 120.555 ;
        RECT 91.450 119.490 91.640 120.385 ;
        RECT 93.540 120.215 93.710 120.725 ;
        RECT 93.880 120.465 94.400 120.775 ;
        RECT 91.810 120.045 93.710 120.215 ;
        RECT 91.810 119.985 92.140 120.045 ;
        RECT 92.290 119.815 92.620 119.875 ;
        RECT 91.960 119.545 92.620 119.815 ;
        RECT 91.450 119.160 91.770 119.490 ;
        RECT 91.950 118.895 92.610 119.375 ;
        RECT 92.810 119.285 92.980 120.045 ;
        RECT 93.880 119.875 94.060 120.285 ;
        RECT 93.150 119.705 93.480 119.825 ;
        RECT 94.230 119.705 94.400 120.465 ;
        RECT 93.150 119.535 94.400 119.705 ;
        RECT 94.570 120.645 95.940 120.895 ;
        RECT 94.570 119.875 94.760 120.645 ;
        RECT 95.690 120.385 95.940 120.645 ;
        RECT 94.930 120.215 95.180 120.375 ;
        RECT 96.110 120.215 96.280 121.060 ;
        RECT 97.175 120.775 97.345 121.275 ;
        RECT 97.515 120.945 97.845 121.445 ;
        RECT 96.450 120.385 96.950 120.765 ;
        RECT 97.175 120.605 97.870 120.775 ;
        RECT 94.930 120.045 96.280 120.215 ;
        RECT 95.860 120.005 96.280 120.045 ;
        RECT 94.570 119.535 94.990 119.875 ;
        RECT 95.280 119.545 95.690 119.875 ;
        RECT 92.810 119.115 93.660 119.285 ;
        RECT 94.220 118.895 94.540 119.355 ;
        RECT 94.740 119.105 94.990 119.535 ;
        RECT 95.280 118.895 95.690 119.335 ;
        RECT 95.860 119.275 96.030 120.005 ;
        RECT 96.200 119.455 96.550 119.825 ;
        RECT 96.730 119.515 96.950 120.385 ;
        RECT 97.120 119.815 97.530 120.435 ;
        RECT 97.700 119.635 97.870 120.605 ;
        RECT 97.175 119.445 97.870 119.635 ;
        RECT 95.860 119.075 96.875 119.275 ;
        RECT 97.175 119.115 97.345 119.445 ;
        RECT 97.515 118.895 97.845 119.275 ;
        RECT 98.060 119.155 98.285 121.275 ;
        RECT 98.455 120.945 98.785 121.445 ;
        RECT 98.955 120.775 99.125 121.275 ;
        RECT 98.460 120.605 99.125 120.775 ;
        RECT 98.460 119.615 98.690 120.605 ;
        RECT 99.385 120.475 99.665 121.445 ;
        RECT 98.860 119.785 99.210 120.435 ;
        RECT 99.835 120.100 100.165 121.275 ;
        RECT 100.335 120.475 100.595 121.445 ;
        RECT 101.685 120.280 101.975 121.445 ;
        RECT 102.145 120.355 103.815 121.445 ;
        RECT 103.985 120.370 104.255 121.275 ;
        RECT 104.425 120.685 104.755 121.445 ;
        RECT 104.935 120.515 105.105 121.275 ;
        RECT 98.460 119.445 99.125 119.615 ;
        RECT 99.385 119.570 100.165 120.100 ;
        RECT 98.455 118.895 98.785 119.275 ;
        RECT 98.955 119.155 99.125 119.445 ;
        RECT 99.385 118.895 99.670 119.400 ;
        RECT 99.840 119.065 100.165 119.570 ;
        RECT 100.355 119.185 100.595 120.135 ;
        RECT 102.145 119.835 102.895 120.355 ;
        RECT 103.065 119.665 103.815 120.185 ;
        RECT 101.685 118.895 101.975 119.620 ;
        RECT 102.145 118.895 103.815 119.665 ;
        RECT 103.985 119.570 104.155 120.370 ;
        RECT 104.440 120.345 105.105 120.515 ;
        RECT 105.365 120.355 107.035 121.445 ;
        RECT 107.210 121.010 112.555 121.445 ;
        RECT 112.730 121.010 118.075 121.445 ;
        RECT 104.440 120.200 104.610 120.345 ;
        RECT 104.325 119.870 104.610 120.200 ;
        RECT 104.440 119.615 104.610 119.870 ;
        RECT 104.845 119.795 105.175 120.165 ;
        RECT 105.365 119.835 106.115 120.355 ;
        RECT 106.285 119.665 107.035 120.185 ;
        RECT 108.800 119.760 109.150 121.010 ;
        RECT 103.985 119.065 104.245 119.570 ;
        RECT 104.440 119.445 105.105 119.615 ;
        RECT 104.425 118.895 104.755 119.275 ;
        RECT 104.935 119.065 105.105 119.445 ;
        RECT 105.365 118.895 107.035 119.665 ;
        RECT 110.630 119.440 110.970 120.270 ;
        RECT 114.320 119.760 114.670 121.010 ;
        RECT 118.285 120.305 118.515 121.445 ;
        RECT 118.685 120.295 119.015 121.275 ;
        RECT 119.185 120.305 119.395 121.445 ;
        RECT 119.715 120.515 119.885 121.275 ;
        RECT 120.065 120.685 120.395 121.445 ;
        RECT 119.715 120.345 120.380 120.515 ;
        RECT 120.565 120.370 120.835 121.275 ;
        RECT 121.010 121.010 126.355 121.445 ;
        RECT 116.150 119.440 116.490 120.270 ;
        RECT 118.265 119.885 118.595 120.135 ;
        RECT 107.210 118.895 112.555 119.440 ;
        RECT 112.730 118.895 118.075 119.440 ;
        RECT 118.285 118.895 118.515 119.715 ;
        RECT 118.765 119.695 119.015 120.295 ;
        RECT 120.210 120.200 120.380 120.345 ;
        RECT 119.645 119.795 119.975 120.165 ;
        RECT 120.210 119.870 120.495 120.200 ;
        RECT 118.685 119.065 119.015 119.695 ;
        RECT 119.185 118.895 119.395 119.715 ;
        RECT 120.210 119.615 120.380 119.870 ;
        RECT 119.715 119.445 120.380 119.615 ;
        RECT 120.665 119.570 120.835 120.370 ;
        RECT 122.600 119.760 122.950 121.010 ;
        RECT 126.525 120.355 127.735 121.445 ;
        RECT 119.715 119.065 119.885 119.445 ;
        RECT 120.065 118.895 120.395 119.275 ;
        RECT 120.575 119.065 120.835 119.570 ;
        RECT 124.430 119.440 124.770 120.270 ;
        RECT 126.525 119.815 127.045 120.355 ;
        RECT 127.215 119.645 127.735 120.185 ;
        RECT 121.010 118.895 126.355 119.440 ;
        RECT 126.525 118.895 127.735 119.645 ;
        RECT 14.660 118.725 127.820 118.895 ;
        RECT 14.745 117.975 15.955 118.725 ;
        RECT 14.745 117.435 15.265 117.975 ;
        RECT 16.125 117.955 17.795 118.725 ;
        RECT 15.435 117.265 15.955 117.805 ;
        RECT 14.745 116.175 15.955 117.265 ;
        RECT 16.125 117.265 16.875 117.785 ;
        RECT 17.045 117.435 17.795 117.955 ;
        RECT 18.240 117.915 18.485 118.520 ;
        RECT 18.705 118.190 19.215 118.725 ;
        RECT 17.965 117.745 19.195 117.915 ;
        RECT 16.125 116.175 17.795 117.265 ;
        RECT 17.965 116.935 18.305 117.745 ;
        RECT 18.475 117.180 19.225 117.370 ;
        RECT 17.965 116.525 18.480 116.935 ;
        RECT 18.715 116.175 18.885 116.935 ;
        RECT 19.055 116.515 19.225 117.180 ;
        RECT 19.395 117.195 19.585 118.555 ;
        RECT 19.755 118.385 20.030 118.555 ;
        RECT 19.755 118.215 20.035 118.385 ;
        RECT 19.755 117.395 20.030 118.215 ;
        RECT 20.220 118.190 20.750 118.555 ;
        RECT 21.175 118.325 21.505 118.725 ;
        RECT 20.575 118.155 20.750 118.190 ;
        RECT 20.235 117.195 20.405 117.995 ;
        RECT 19.395 117.025 20.405 117.195 ;
        RECT 20.575 117.985 21.505 118.155 ;
        RECT 21.675 117.985 21.930 118.555 ;
        RECT 22.195 118.175 22.365 118.465 ;
        RECT 22.535 118.345 22.865 118.725 ;
        RECT 22.195 118.005 22.860 118.175 ;
        RECT 20.575 116.855 20.745 117.985 ;
        RECT 21.335 117.815 21.505 117.985 ;
        RECT 19.620 116.685 20.745 116.855 ;
        RECT 20.915 117.485 21.110 117.815 ;
        RECT 21.335 117.485 21.590 117.815 ;
        RECT 20.915 116.515 21.085 117.485 ;
        RECT 21.760 117.315 21.930 117.985 ;
        RECT 19.055 116.345 21.085 116.515 ;
        RECT 21.255 116.175 21.425 117.315 ;
        RECT 21.595 116.345 21.930 117.315 ;
        RECT 22.110 117.185 22.460 117.835 ;
        RECT 22.630 117.015 22.860 118.005 ;
        RECT 22.195 116.845 22.860 117.015 ;
        RECT 22.195 116.345 22.365 116.845 ;
        RECT 22.535 116.175 22.865 116.675 ;
        RECT 23.035 116.345 23.260 118.465 ;
        RECT 23.475 118.345 23.805 118.725 ;
        RECT 23.975 118.175 24.145 118.505 ;
        RECT 24.445 118.345 25.460 118.545 ;
        RECT 23.450 117.985 24.145 118.175 ;
        RECT 23.450 117.015 23.620 117.985 ;
        RECT 23.790 117.185 24.200 117.805 ;
        RECT 24.370 117.235 24.590 118.105 ;
        RECT 24.770 117.795 25.120 118.165 ;
        RECT 25.290 117.615 25.460 118.345 ;
        RECT 25.630 118.285 26.040 118.725 ;
        RECT 26.330 118.085 26.580 118.515 ;
        RECT 26.780 118.265 27.100 118.725 ;
        RECT 27.660 118.335 28.510 118.505 ;
        RECT 25.630 117.745 26.040 118.075 ;
        RECT 26.330 117.745 26.750 118.085 ;
        RECT 25.040 117.575 25.460 117.615 ;
        RECT 25.040 117.405 26.390 117.575 ;
        RECT 23.450 116.845 24.145 117.015 ;
        RECT 24.370 116.855 24.870 117.235 ;
        RECT 23.475 116.175 23.805 116.675 ;
        RECT 23.975 116.345 24.145 116.845 ;
        RECT 25.040 116.560 25.210 117.405 ;
        RECT 26.140 117.245 26.390 117.405 ;
        RECT 25.380 116.975 25.630 117.235 ;
        RECT 26.560 116.975 26.750 117.745 ;
        RECT 25.380 116.725 26.750 116.975 ;
        RECT 26.920 117.915 28.170 118.085 ;
        RECT 26.920 117.155 27.090 117.915 ;
        RECT 27.840 117.795 28.170 117.915 ;
        RECT 27.260 117.335 27.440 117.745 ;
        RECT 28.340 117.575 28.510 118.335 ;
        RECT 28.710 118.245 29.370 118.725 ;
        RECT 29.550 118.130 29.870 118.460 ;
        RECT 28.700 117.805 29.360 118.075 ;
        RECT 28.700 117.745 29.030 117.805 ;
        RECT 29.180 117.575 29.510 117.635 ;
        RECT 27.610 117.405 29.510 117.575 ;
        RECT 26.920 116.845 27.440 117.155 ;
        RECT 27.610 116.895 27.780 117.405 ;
        RECT 29.680 117.235 29.870 118.130 ;
        RECT 27.950 117.065 29.870 117.235 ;
        RECT 29.550 117.045 29.870 117.065 ;
        RECT 30.070 117.815 30.320 118.465 ;
        RECT 30.500 118.265 30.785 118.725 ;
        RECT 30.965 118.015 31.220 118.545 ;
        RECT 30.070 117.485 30.870 117.815 ;
        RECT 31.040 117.705 31.220 118.015 ;
        RECT 31.805 117.905 32.035 118.725 ;
        RECT 32.205 117.925 32.535 118.555 ;
        RECT 31.040 117.535 31.305 117.705 ;
        RECT 27.610 116.725 28.820 116.895 ;
        RECT 24.380 116.390 25.210 116.560 ;
        RECT 25.450 116.175 25.830 116.555 ;
        RECT 26.010 116.435 26.180 116.725 ;
        RECT 27.610 116.645 27.780 116.725 ;
        RECT 26.350 116.175 26.680 116.555 ;
        RECT 27.150 116.395 27.780 116.645 ;
        RECT 27.960 116.175 28.380 116.555 ;
        RECT 28.580 116.435 28.820 116.725 ;
        RECT 29.050 116.175 29.380 116.865 ;
        RECT 29.550 116.435 29.720 117.045 ;
        RECT 30.070 116.895 30.320 117.485 ;
        RECT 31.040 117.155 31.220 117.535 ;
        RECT 31.785 117.485 32.115 117.735 ;
        RECT 32.285 117.325 32.535 117.925 ;
        RECT 32.705 117.905 32.915 118.725 ;
        RECT 33.420 117.915 33.665 118.520 ;
        RECT 33.885 118.190 34.395 118.725 ;
        RECT 29.990 116.385 30.320 116.895 ;
        RECT 30.500 116.175 30.785 116.975 ;
        RECT 30.965 116.485 31.220 117.155 ;
        RECT 31.805 116.175 32.035 117.315 ;
        RECT 32.205 116.345 32.535 117.325 ;
        RECT 33.145 117.745 34.375 117.915 ;
        RECT 32.705 116.175 32.915 117.315 ;
        RECT 33.145 116.935 33.485 117.745 ;
        RECT 33.655 117.180 34.405 117.370 ;
        RECT 33.145 116.525 33.660 116.935 ;
        RECT 33.895 116.175 34.065 116.935 ;
        RECT 34.235 116.515 34.405 117.180 ;
        RECT 34.575 117.195 34.765 118.555 ;
        RECT 34.935 118.385 35.210 118.555 ;
        RECT 34.935 118.215 35.215 118.385 ;
        RECT 34.935 117.395 35.210 118.215 ;
        RECT 35.400 118.190 35.930 118.555 ;
        RECT 36.355 118.325 36.685 118.725 ;
        RECT 35.755 118.155 35.930 118.190 ;
        RECT 35.415 117.195 35.585 117.995 ;
        RECT 34.575 117.025 35.585 117.195 ;
        RECT 35.755 117.985 36.685 118.155 ;
        RECT 36.855 117.985 37.110 118.555 ;
        RECT 37.285 118.000 37.575 118.725 ;
        RECT 37.835 118.175 38.005 118.555 ;
        RECT 38.185 118.345 38.515 118.725 ;
        RECT 37.835 118.005 38.500 118.175 ;
        RECT 38.695 118.050 38.955 118.555 ;
        RECT 35.755 116.855 35.925 117.985 ;
        RECT 36.515 117.815 36.685 117.985 ;
        RECT 34.800 116.685 35.925 116.855 ;
        RECT 36.095 117.485 36.290 117.815 ;
        RECT 36.515 117.485 36.770 117.815 ;
        RECT 36.095 116.515 36.265 117.485 ;
        RECT 36.940 117.315 37.110 117.985 ;
        RECT 37.765 117.455 38.095 117.825 ;
        RECT 38.330 117.750 38.500 118.005 ;
        RECT 38.330 117.420 38.615 117.750 ;
        RECT 34.235 116.345 36.265 116.515 ;
        RECT 36.435 116.175 36.605 117.315 ;
        RECT 36.775 116.345 37.110 117.315 ;
        RECT 37.285 116.175 37.575 117.340 ;
        RECT 38.330 117.275 38.500 117.420 ;
        RECT 37.835 117.105 38.500 117.275 ;
        RECT 38.785 117.250 38.955 118.050 ;
        RECT 39.215 118.175 39.385 118.555 ;
        RECT 39.565 118.345 39.895 118.725 ;
        RECT 39.215 118.005 39.880 118.175 ;
        RECT 40.075 118.050 40.335 118.555 ;
        RECT 40.880 118.385 41.135 118.545 ;
        RECT 40.795 118.215 41.135 118.385 ;
        RECT 41.315 118.265 41.600 118.725 ;
        RECT 39.145 117.455 39.475 117.825 ;
        RECT 39.710 117.750 39.880 118.005 ;
        RECT 39.710 117.420 39.995 117.750 ;
        RECT 39.710 117.275 39.880 117.420 ;
        RECT 37.835 116.345 38.005 117.105 ;
        RECT 38.185 116.175 38.515 116.935 ;
        RECT 38.685 116.345 38.955 117.250 ;
        RECT 39.215 117.105 39.880 117.275 ;
        RECT 40.165 117.250 40.335 118.050 ;
        RECT 39.215 116.345 39.385 117.105 ;
        RECT 39.565 116.175 39.895 116.935 ;
        RECT 40.065 116.345 40.335 117.250 ;
        RECT 40.880 118.015 41.135 118.215 ;
        RECT 40.880 117.155 41.060 118.015 ;
        RECT 41.780 117.815 42.030 118.465 ;
        RECT 41.230 117.485 42.030 117.815 ;
        RECT 40.880 116.485 41.135 117.155 ;
        RECT 41.315 116.175 41.600 116.975 ;
        RECT 41.780 116.895 42.030 117.485 ;
        RECT 42.230 118.130 42.550 118.460 ;
        RECT 42.730 118.245 43.390 118.725 ;
        RECT 43.590 118.335 44.440 118.505 ;
        RECT 42.230 117.235 42.420 118.130 ;
        RECT 42.740 117.805 43.400 118.075 ;
        RECT 43.070 117.745 43.400 117.805 ;
        RECT 42.590 117.575 42.920 117.635 ;
        RECT 43.590 117.575 43.760 118.335 ;
        RECT 45.000 118.265 45.320 118.725 ;
        RECT 45.520 118.085 45.770 118.515 ;
        RECT 46.060 118.285 46.470 118.725 ;
        RECT 46.640 118.345 47.655 118.545 ;
        RECT 43.930 117.915 45.180 118.085 ;
        RECT 43.930 117.795 44.260 117.915 ;
        RECT 42.590 117.405 44.490 117.575 ;
        RECT 42.230 117.065 44.150 117.235 ;
        RECT 42.230 117.045 42.550 117.065 ;
        RECT 41.780 116.385 42.110 116.895 ;
        RECT 42.380 116.435 42.550 117.045 ;
        RECT 44.320 116.895 44.490 117.405 ;
        RECT 44.660 117.335 44.840 117.745 ;
        RECT 45.010 117.155 45.180 117.915 ;
        RECT 42.720 116.175 43.050 116.865 ;
        RECT 43.280 116.725 44.490 116.895 ;
        RECT 44.660 116.845 45.180 117.155 ;
        RECT 45.350 117.745 45.770 118.085 ;
        RECT 46.060 117.745 46.470 118.075 ;
        RECT 45.350 116.975 45.540 117.745 ;
        RECT 46.640 117.615 46.810 118.345 ;
        RECT 47.955 118.175 48.125 118.505 ;
        RECT 48.295 118.345 48.625 118.725 ;
        RECT 46.980 117.795 47.330 118.165 ;
        RECT 46.640 117.575 47.060 117.615 ;
        RECT 45.710 117.405 47.060 117.575 ;
        RECT 45.710 117.245 45.960 117.405 ;
        RECT 46.470 116.975 46.720 117.235 ;
        RECT 45.350 116.725 46.720 116.975 ;
        RECT 43.280 116.435 43.520 116.725 ;
        RECT 44.320 116.645 44.490 116.725 ;
        RECT 43.720 116.175 44.140 116.555 ;
        RECT 44.320 116.395 44.950 116.645 ;
        RECT 45.420 116.175 45.750 116.555 ;
        RECT 45.920 116.435 46.090 116.725 ;
        RECT 46.890 116.560 47.060 117.405 ;
        RECT 47.510 117.235 47.730 118.105 ;
        RECT 47.955 117.985 48.650 118.175 ;
        RECT 47.230 116.855 47.730 117.235 ;
        RECT 47.900 117.185 48.310 117.805 ;
        RECT 48.480 117.015 48.650 117.985 ;
        RECT 47.955 116.845 48.650 117.015 ;
        RECT 46.270 116.175 46.650 116.555 ;
        RECT 46.890 116.390 47.720 116.560 ;
        RECT 47.955 116.345 48.125 116.845 ;
        RECT 48.295 116.175 48.625 116.675 ;
        RECT 48.840 116.345 49.065 118.465 ;
        RECT 49.235 118.345 49.565 118.725 ;
        RECT 49.735 118.175 49.905 118.465 ;
        RECT 49.240 118.005 49.905 118.175 ;
        RECT 50.540 118.015 50.795 118.545 ;
        RECT 50.975 118.265 51.260 118.725 ;
        RECT 49.240 117.015 49.470 118.005 ;
        RECT 49.640 117.185 49.990 117.835 ;
        RECT 50.540 117.365 50.720 118.015 ;
        RECT 51.440 117.815 51.690 118.465 ;
        RECT 50.890 117.485 51.690 117.815 ;
        RECT 50.455 117.195 50.720 117.365 ;
        RECT 50.540 117.155 50.720 117.195 ;
        RECT 49.240 116.845 49.905 117.015 ;
        RECT 49.235 116.175 49.565 116.675 ;
        RECT 49.735 116.345 49.905 116.845 ;
        RECT 50.540 116.485 50.795 117.155 ;
        RECT 50.975 116.175 51.260 116.975 ;
        RECT 51.440 116.895 51.690 117.485 ;
        RECT 51.890 118.130 52.210 118.460 ;
        RECT 52.390 118.245 53.050 118.725 ;
        RECT 53.250 118.335 54.100 118.505 ;
        RECT 51.890 117.235 52.080 118.130 ;
        RECT 52.400 117.805 53.060 118.075 ;
        RECT 52.730 117.745 53.060 117.805 ;
        RECT 52.250 117.575 52.580 117.635 ;
        RECT 53.250 117.575 53.420 118.335 ;
        RECT 54.660 118.265 54.980 118.725 ;
        RECT 55.180 118.085 55.430 118.515 ;
        RECT 55.720 118.285 56.130 118.725 ;
        RECT 56.300 118.345 57.315 118.545 ;
        RECT 53.590 117.915 54.840 118.085 ;
        RECT 53.590 117.795 53.920 117.915 ;
        RECT 52.250 117.405 54.150 117.575 ;
        RECT 51.890 117.065 53.810 117.235 ;
        RECT 51.890 117.045 52.210 117.065 ;
        RECT 51.440 116.385 51.770 116.895 ;
        RECT 52.040 116.435 52.210 117.045 ;
        RECT 53.980 116.895 54.150 117.405 ;
        RECT 54.320 117.335 54.500 117.745 ;
        RECT 54.670 117.155 54.840 117.915 ;
        RECT 52.380 116.175 52.710 116.865 ;
        RECT 52.940 116.725 54.150 116.895 ;
        RECT 54.320 116.845 54.840 117.155 ;
        RECT 55.010 117.745 55.430 118.085 ;
        RECT 55.720 117.745 56.130 118.075 ;
        RECT 55.010 116.975 55.200 117.745 ;
        RECT 56.300 117.615 56.470 118.345 ;
        RECT 57.615 118.175 57.785 118.505 ;
        RECT 57.955 118.345 58.285 118.725 ;
        RECT 56.640 117.795 56.990 118.165 ;
        RECT 56.300 117.575 56.720 117.615 ;
        RECT 55.370 117.405 56.720 117.575 ;
        RECT 55.370 117.245 55.620 117.405 ;
        RECT 56.130 116.975 56.380 117.235 ;
        RECT 55.010 116.725 56.380 116.975 ;
        RECT 52.940 116.435 53.180 116.725 ;
        RECT 53.980 116.645 54.150 116.725 ;
        RECT 53.380 116.175 53.800 116.555 ;
        RECT 53.980 116.395 54.610 116.645 ;
        RECT 55.080 116.175 55.410 116.555 ;
        RECT 55.580 116.435 55.750 116.725 ;
        RECT 56.550 116.560 56.720 117.405 ;
        RECT 57.170 117.235 57.390 118.105 ;
        RECT 57.615 117.985 58.310 118.175 ;
        RECT 56.890 116.855 57.390 117.235 ;
        RECT 57.560 117.185 57.970 117.805 ;
        RECT 58.140 117.015 58.310 117.985 ;
        RECT 57.615 116.845 58.310 117.015 ;
        RECT 55.930 116.175 56.310 116.555 ;
        RECT 56.550 116.390 57.380 116.560 ;
        RECT 57.615 116.345 57.785 116.845 ;
        RECT 57.955 116.175 58.285 116.675 ;
        RECT 58.500 116.345 58.725 118.465 ;
        RECT 58.895 118.345 59.225 118.725 ;
        RECT 59.395 118.175 59.565 118.465 ;
        RECT 58.900 118.005 59.565 118.175 ;
        RECT 58.900 117.015 59.130 118.005 ;
        RECT 60.285 117.955 62.875 118.725 ;
        RECT 63.045 118.000 63.335 118.725 ;
        RECT 64.800 118.015 65.055 118.545 ;
        RECT 65.235 118.265 65.520 118.725 ;
        RECT 59.300 117.185 59.650 117.835 ;
        RECT 60.285 117.265 61.495 117.785 ;
        RECT 61.665 117.435 62.875 117.955 ;
        RECT 58.900 116.845 59.565 117.015 ;
        RECT 58.895 116.175 59.225 116.675 ;
        RECT 59.395 116.345 59.565 116.845 ;
        RECT 60.285 116.175 62.875 117.265 ;
        RECT 63.045 116.175 63.335 117.340 ;
        RECT 64.800 117.155 64.980 118.015 ;
        RECT 65.700 117.815 65.950 118.465 ;
        RECT 65.150 117.485 65.950 117.815 ;
        RECT 64.800 116.685 65.055 117.155 ;
        RECT 64.715 116.515 65.055 116.685 ;
        RECT 64.800 116.485 65.055 116.515 ;
        RECT 65.235 116.175 65.520 116.975 ;
        RECT 65.700 116.895 65.950 117.485 ;
        RECT 66.150 118.130 66.470 118.460 ;
        RECT 66.650 118.245 67.310 118.725 ;
        RECT 67.510 118.335 68.360 118.505 ;
        RECT 66.150 117.235 66.340 118.130 ;
        RECT 66.660 117.805 67.320 118.075 ;
        RECT 66.990 117.745 67.320 117.805 ;
        RECT 66.510 117.575 66.840 117.635 ;
        RECT 67.510 117.575 67.680 118.335 ;
        RECT 68.920 118.265 69.240 118.725 ;
        RECT 69.440 118.085 69.690 118.515 ;
        RECT 69.980 118.285 70.390 118.725 ;
        RECT 70.560 118.345 71.575 118.545 ;
        RECT 67.850 117.915 69.100 118.085 ;
        RECT 67.850 117.795 68.180 117.915 ;
        RECT 66.510 117.405 68.410 117.575 ;
        RECT 66.150 117.065 68.070 117.235 ;
        RECT 66.150 117.045 66.470 117.065 ;
        RECT 65.700 116.385 66.030 116.895 ;
        RECT 66.300 116.435 66.470 117.045 ;
        RECT 68.240 116.895 68.410 117.405 ;
        RECT 68.580 117.335 68.760 117.745 ;
        RECT 68.930 117.155 69.100 117.915 ;
        RECT 66.640 116.175 66.970 116.865 ;
        RECT 67.200 116.725 68.410 116.895 ;
        RECT 68.580 116.845 69.100 117.155 ;
        RECT 69.270 117.745 69.690 118.085 ;
        RECT 69.980 117.745 70.390 118.075 ;
        RECT 69.270 116.975 69.460 117.745 ;
        RECT 70.560 117.615 70.730 118.345 ;
        RECT 71.875 118.175 72.045 118.505 ;
        RECT 72.215 118.345 72.545 118.725 ;
        RECT 70.900 117.795 71.250 118.165 ;
        RECT 70.560 117.575 70.980 117.615 ;
        RECT 69.630 117.405 70.980 117.575 ;
        RECT 69.630 117.245 69.880 117.405 ;
        RECT 70.390 116.975 70.640 117.235 ;
        RECT 69.270 116.725 70.640 116.975 ;
        RECT 67.200 116.435 67.440 116.725 ;
        RECT 68.240 116.645 68.410 116.725 ;
        RECT 67.640 116.175 68.060 116.555 ;
        RECT 68.240 116.395 68.870 116.645 ;
        RECT 69.340 116.175 69.670 116.555 ;
        RECT 69.840 116.435 70.010 116.725 ;
        RECT 70.810 116.560 70.980 117.405 ;
        RECT 71.430 117.235 71.650 118.105 ;
        RECT 71.875 117.985 72.570 118.175 ;
        RECT 71.150 116.855 71.650 117.235 ;
        RECT 71.820 117.185 72.230 117.805 ;
        RECT 72.400 117.015 72.570 117.985 ;
        RECT 71.875 116.845 72.570 117.015 ;
        RECT 70.190 116.175 70.570 116.555 ;
        RECT 70.810 116.390 71.640 116.560 ;
        RECT 71.875 116.345 72.045 116.845 ;
        RECT 72.215 116.175 72.545 116.675 ;
        RECT 72.760 116.345 72.985 118.465 ;
        RECT 73.155 118.345 73.485 118.725 ;
        RECT 73.655 118.175 73.825 118.465 ;
        RECT 73.160 118.005 73.825 118.175 ;
        RECT 73.160 117.015 73.390 118.005 ;
        RECT 74.545 117.955 76.215 118.725 ;
        RECT 73.560 117.185 73.910 117.835 ;
        RECT 74.545 117.265 75.295 117.785 ;
        RECT 75.465 117.435 76.215 117.955 ;
        RECT 76.760 118.015 77.015 118.545 ;
        RECT 77.195 118.265 77.480 118.725 ;
        RECT 73.160 116.845 73.825 117.015 ;
        RECT 73.155 116.175 73.485 116.675 ;
        RECT 73.655 116.345 73.825 116.845 ;
        RECT 74.545 116.175 76.215 117.265 ;
        RECT 76.760 117.155 76.940 118.015 ;
        RECT 77.660 117.815 77.910 118.465 ;
        RECT 77.110 117.485 77.910 117.815 ;
        RECT 76.760 116.685 77.015 117.155 ;
        RECT 76.675 116.515 77.015 116.685 ;
        RECT 76.760 116.485 77.015 116.515 ;
        RECT 77.195 116.175 77.480 116.975 ;
        RECT 77.660 116.895 77.910 117.485 ;
        RECT 78.110 118.130 78.430 118.460 ;
        RECT 78.610 118.245 79.270 118.725 ;
        RECT 79.470 118.335 80.320 118.505 ;
        RECT 78.110 117.235 78.300 118.130 ;
        RECT 78.620 117.805 79.280 118.075 ;
        RECT 78.950 117.745 79.280 117.805 ;
        RECT 78.470 117.575 78.800 117.635 ;
        RECT 79.470 117.575 79.640 118.335 ;
        RECT 80.880 118.265 81.200 118.725 ;
        RECT 81.400 118.085 81.650 118.515 ;
        RECT 81.940 118.285 82.350 118.725 ;
        RECT 82.520 118.345 83.535 118.545 ;
        RECT 79.810 117.915 81.060 118.085 ;
        RECT 79.810 117.795 80.140 117.915 ;
        RECT 78.470 117.405 80.370 117.575 ;
        RECT 78.110 117.065 80.030 117.235 ;
        RECT 78.110 117.045 78.430 117.065 ;
        RECT 77.660 116.385 77.990 116.895 ;
        RECT 78.260 116.435 78.430 117.045 ;
        RECT 80.200 116.895 80.370 117.405 ;
        RECT 80.540 117.335 80.720 117.745 ;
        RECT 80.890 117.155 81.060 117.915 ;
        RECT 78.600 116.175 78.930 116.865 ;
        RECT 79.160 116.725 80.370 116.895 ;
        RECT 80.540 116.845 81.060 117.155 ;
        RECT 81.230 117.745 81.650 118.085 ;
        RECT 81.940 117.745 82.350 118.075 ;
        RECT 81.230 116.975 81.420 117.745 ;
        RECT 82.520 117.615 82.690 118.345 ;
        RECT 83.835 118.175 84.005 118.505 ;
        RECT 84.175 118.345 84.505 118.725 ;
        RECT 82.860 117.795 83.210 118.165 ;
        RECT 82.520 117.575 82.940 117.615 ;
        RECT 81.590 117.405 82.940 117.575 ;
        RECT 81.590 117.245 81.840 117.405 ;
        RECT 82.350 116.975 82.600 117.235 ;
        RECT 81.230 116.725 82.600 116.975 ;
        RECT 79.160 116.435 79.400 116.725 ;
        RECT 80.200 116.645 80.370 116.725 ;
        RECT 79.600 116.175 80.020 116.555 ;
        RECT 80.200 116.395 80.830 116.645 ;
        RECT 81.300 116.175 81.630 116.555 ;
        RECT 81.800 116.435 81.970 116.725 ;
        RECT 82.770 116.560 82.940 117.405 ;
        RECT 83.390 117.235 83.610 118.105 ;
        RECT 83.835 117.985 84.530 118.175 ;
        RECT 83.110 116.855 83.610 117.235 ;
        RECT 83.780 117.185 84.190 117.805 ;
        RECT 84.360 117.015 84.530 117.985 ;
        RECT 83.835 116.845 84.530 117.015 ;
        RECT 82.150 116.175 82.530 116.555 ;
        RECT 82.770 116.390 83.600 116.560 ;
        RECT 83.835 116.345 84.005 116.845 ;
        RECT 84.175 116.175 84.505 116.675 ;
        RECT 84.720 116.345 84.945 118.465 ;
        RECT 85.115 118.345 85.445 118.725 ;
        RECT 85.615 118.175 85.785 118.465 ;
        RECT 85.120 118.005 85.785 118.175 ;
        RECT 85.120 117.015 85.350 118.005 ;
        RECT 86.045 117.975 87.255 118.725 ;
        RECT 85.520 117.185 85.870 117.835 ;
        RECT 86.045 117.265 86.565 117.805 ;
        RECT 86.735 117.435 87.255 117.975 ;
        RECT 87.465 117.905 87.695 118.725 ;
        RECT 87.865 117.925 88.195 118.555 ;
        RECT 87.445 117.485 87.775 117.735 ;
        RECT 87.945 117.325 88.195 117.925 ;
        RECT 88.365 117.905 88.575 118.725 ;
        RECT 88.805 118.000 89.095 118.725 ;
        RECT 89.265 118.215 89.570 118.725 ;
        RECT 89.265 117.485 89.580 118.045 ;
        RECT 89.750 117.735 90.000 118.545 ;
        RECT 90.170 118.200 90.430 118.725 ;
        RECT 90.610 117.735 90.860 118.545 ;
        RECT 91.030 118.165 91.290 118.725 ;
        RECT 91.460 118.075 91.720 118.530 ;
        RECT 91.890 118.245 92.150 118.725 ;
        RECT 92.320 118.075 92.580 118.530 ;
        RECT 92.750 118.245 93.010 118.725 ;
        RECT 93.180 118.075 93.440 118.530 ;
        RECT 93.610 118.245 93.855 118.725 ;
        RECT 94.025 118.075 94.300 118.530 ;
        RECT 94.470 118.245 94.715 118.725 ;
        RECT 94.885 118.075 95.145 118.530 ;
        RECT 95.325 118.245 95.575 118.725 ;
        RECT 95.745 118.075 96.005 118.530 ;
        RECT 96.185 118.245 96.435 118.725 ;
        RECT 96.605 118.075 96.865 118.530 ;
        RECT 97.045 118.245 97.305 118.725 ;
        RECT 97.475 118.075 97.735 118.530 ;
        RECT 97.905 118.245 98.205 118.725 ;
        RECT 91.460 118.045 98.205 118.075 ;
        RECT 91.460 117.905 98.235 118.045 ;
        RECT 98.505 117.905 98.735 118.725 ;
        RECT 98.905 117.925 99.235 118.555 ;
        RECT 97.040 117.875 98.235 117.905 ;
        RECT 89.750 117.485 96.870 117.735 ;
        RECT 85.120 116.845 85.785 117.015 ;
        RECT 85.115 116.175 85.445 116.675 ;
        RECT 85.615 116.345 85.785 116.845 ;
        RECT 86.045 116.175 87.255 117.265 ;
        RECT 87.465 116.175 87.695 117.315 ;
        RECT 87.865 116.345 88.195 117.325 ;
        RECT 88.365 116.175 88.575 117.315 ;
        RECT 88.805 116.175 89.095 117.340 ;
        RECT 89.275 116.175 89.570 116.985 ;
        RECT 89.750 116.345 89.995 117.485 ;
        RECT 90.170 116.175 90.430 116.985 ;
        RECT 90.610 116.350 90.860 117.485 ;
        RECT 97.040 117.315 98.205 117.875 ;
        RECT 98.485 117.485 98.815 117.735 ;
        RECT 98.985 117.325 99.235 117.925 ;
        RECT 99.405 117.905 99.615 118.725 ;
        RECT 99.845 117.955 103.355 118.725 ;
        RECT 91.460 117.090 98.205 117.315 ;
        RECT 91.460 117.075 96.865 117.090 ;
        RECT 91.030 116.180 91.290 116.975 ;
        RECT 91.460 116.350 91.720 117.075 ;
        RECT 91.890 116.180 92.150 116.905 ;
        RECT 92.320 116.350 92.580 117.075 ;
        RECT 92.750 116.180 93.010 116.905 ;
        RECT 93.180 116.350 93.440 117.075 ;
        RECT 93.610 116.180 93.870 116.905 ;
        RECT 94.040 116.350 94.300 117.075 ;
        RECT 94.470 116.180 94.715 116.905 ;
        RECT 94.885 116.350 95.145 117.075 ;
        RECT 95.330 116.180 95.575 116.905 ;
        RECT 95.745 116.350 96.005 117.075 ;
        RECT 96.190 116.180 96.435 116.905 ;
        RECT 96.605 116.350 96.865 117.075 ;
        RECT 97.050 116.180 97.305 116.905 ;
        RECT 97.475 116.350 97.765 117.090 ;
        RECT 91.030 116.175 97.305 116.180 ;
        RECT 97.935 116.175 98.205 116.920 ;
        RECT 98.505 116.175 98.735 117.315 ;
        RECT 98.905 116.345 99.235 117.325 ;
        RECT 99.405 116.175 99.615 117.315 ;
        RECT 99.845 117.265 101.535 117.785 ;
        RECT 101.705 117.435 103.355 117.955 ;
        RECT 103.565 117.905 103.795 118.725 ;
        RECT 103.965 117.925 104.295 118.555 ;
        RECT 103.545 117.485 103.875 117.735 ;
        RECT 104.045 117.325 104.295 117.925 ;
        RECT 104.465 117.905 104.675 118.725 ;
        RECT 105.180 117.915 105.425 118.520 ;
        RECT 105.645 118.190 106.155 118.725 ;
        RECT 99.845 116.175 103.355 117.265 ;
        RECT 103.565 116.175 103.795 117.315 ;
        RECT 103.965 116.345 104.295 117.325 ;
        RECT 104.905 117.745 106.135 117.915 ;
        RECT 104.465 116.175 104.675 117.315 ;
        RECT 104.905 116.935 105.245 117.745 ;
        RECT 105.415 117.180 106.165 117.370 ;
        RECT 104.905 116.525 105.420 116.935 ;
        RECT 105.655 116.175 105.825 116.935 ;
        RECT 105.995 116.515 106.165 117.180 ;
        RECT 106.335 117.195 106.525 118.555 ;
        RECT 106.695 118.385 106.970 118.555 ;
        RECT 106.695 118.215 106.975 118.385 ;
        RECT 106.695 117.395 106.970 118.215 ;
        RECT 107.160 118.190 107.690 118.555 ;
        RECT 108.115 118.325 108.445 118.725 ;
        RECT 107.515 118.155 107.690 118.190 ;
        RECT 107.175 117.195 107.345 117.995 ;
        RECT 106.335 117.025 107.345 117.195 ;
        RECT 107.515 117.985 108.445 118.155 ;
        RECT 108.615 117.985 108.870 118.555 ;
        RECT 107.515 116.855 107.685 117.985 ;
        RECT 108.275 117.815 108.445 117.985 ;
        RECT 106.560 116.685 107.685 116.855 ;
        RECT 107.855 117.485 108.050 117.815 ;
        RECT 108.275 117.485 108.530 117.815 ;
        RECT 107.855 116.515 108.025 117.485 ;
        RECT 108.700 117.315 108.870 117.985 ;
        RECT 109.045 117.975 110.255 118.725 ;
        RECT 105.995 116.345 108.025 116.515 ;
        RECT 108.195 116.175 108.365 117.315 ;
        RECT 108.535 116.345 108.870 117.315 ;
        RECT 109.045 117.265 109.565 117.805 ;
        RECT 109.735 117.435 110.255 117.975 ;
        RECT 110.700 117.915 110.945 118.520 ;
        RECT 111.165 118.190 111.675 118.725 ;
        RECT 110.425 117.745 111.655 117.915 ;
        RECT 109.045 116.175 110.255 117.265 ;
        RECT 110.425 116.935 110.765 117.745 ;
        RECT 110.935 117.180 111.685 117.370 ;
        RECT 110.425 116.525 110.940 116.935 ;
        RECT 111.175 116.175 111.345 116.935 ;
        RECT 111.515 116.515 111.685 117.180 ;
        RECT 111.855 117.195 112.045 118.555 ;
        RECT 112.215 118.045 112.490 118.555 ;
        RECT 112.680 118.190 113.210 118.555 ;
        RECT 113.635 118.325 113.965 118.725 ;
        RECT 113.035 118.155 113.210 118.190 ;
        RECT 112.215 117.875 112.495 118.045 ;
        RECT 112.215 117.395 112.490 117.875 ;
        RECT 112.695 117.195 112.865 117.995 ;
        RECT 111.855 117.025 112.865 117.195 ;
        RECT 113.035 117.985 113.965 118.155 ;
        RECT 114.135 117.985 114.390 118.555 ;
        RECT 114.565 118.000 114.855 118.725 ;
        RECT 115.400 118.385 115.655 118.545 ;
        RECT 115.315 118.215 115.655 118.385 ;
        RECT 115.835 118.265 116.120 118.725 ;
        RECT 115.400 118.015 115.655 118.215 ;
        RECT 113.035 116.855 113.205 117.985 ;
        RECT 113.795 117.815 113.965 117.985 ;
        RECT 112.080 116.685 113.205 116.855 ;
        RECT 113.375 117.485 113.570 117.815 ;
        RECT 113.795 117.485 114.050 117.815 ;
        RECT 113.375 116.515 113.545 117.485 ;
        RECT 114.220 117.315 114.390 117.985 ;
        RECT 111.515 116.345 113.545 116.515 ;
        RECT 113.715 116.175 113.885 117.315 ;
        RECT 114.055 116.345 114.390 117.315 ;
        RECT 114.565 116.175 114.855 117.340 ;
        RECT 115.400 117.155 115.580 118.015 ;
        RECT 116.300 117.815 116.550 118.465 ;
        RECT 115.750 117.485 116.550 117.815 ;
        RECT 115.400 116.485 115.655 117.155 ;
        RECT 115.835 116.175 116.120 116.975 ;
        RECT 116.300 116.895 116.550 117.485 ;
        RECT 116.750 118.130 117.070 118.460 ;
        RECT 117.250 118.245 117.910 118.725 ;
        RECT 118.110 118.335 118.960 118.505 ;
        RECT 116.750 117.235 116.940 118.130 ;
        RECT 117.260 117.805 117.920 118.075 ;
        RECT 117.590 117.745 117.920 117.805 ;
        RECT 117.110 117.575 117.440 117.635 ;
        RECT 118.110 117.575 118.280 118.335 ;
        RECT 119.520 118.265 119.840 118.725 ;
        RECT 120.040 118.085 120.290 118.515 ;
        RECT 120.580 118.285 120.990 118.725 ;
        RECT 121.160 118.345 122.175 118.545 ;
        RECT 118.450 117.915 119.700 118.085 ;
        RECT 118.450 117.795 118.780 117.915 ;
        RECT 117.110 117.405 119.010 117.575 ;
        RECT 116.750 117.065 118.670 117.235 ;
        RECT 116.750 117.045 117.070 117.065 ;
        RECT 116.300 116.385 116.630 116.895 ;
        RECT 116.900 116.435 117.070 117.045 ;
        RECT 118.840 116.895 119.010 117.405 ;
        RECT 119.180 117.335 119.360 117.745 ;
        RECT 119.530 117.155 119.700 117.915 ;
        RECT 117.240 116.175 117.570 116.865 ;
        RECT 117.800 116.725 119.010 116.895 ;
        RECT 119.180 116.845 119.700 117.155 ;
        RECT 119.870 117.745 120.290 118.085 ;
        RECT 120.580 117.745 120.990 118.075 ;
        RECT 119.870 116.975 120.060 117.745 ;
        RECT 121.160 117.615 121.330 118.345 ;
        RECT 122.475 118.175 122.645 118.505 ;
        RECT 122.815 118.345 123.145 118.725 ;
        RECT 121.500 117.795 121.850 118.165 ;
        RECT 121.160 117.575 121.580 117.615 ;
        RECT 120.230 117.405 121.580 117.575 ;
        RECT 120.230 117.245 120.480 117.405 ;
        RECT 120.990 116.975 121.240 117.235 ;
        RECT 119.870 116.725 121.240 116.975 ;
        RECT 117.800 116.435 118.040 116.725 ;
        RECT 118.840 116.645 119.010 116.725 ;
        RECT 118.240 116.175 118.660 116.555 ;
        RECT 118.840 116.395 119.470 116.645 ;
        RECT 119.940 116.175 120.270 116.555 ;
        RECT 120.440 116.435 120.610 116.725 ;
        RECT 121.410 116.560 121.580 117.405 ;
        RECT 122.030 117.235 122.250 118.105 ;
        RECT 122.475 117.985 123.170 118.175 ;
        RECT 121.750 116.855 122.250 117.235 ;
        RECT 122.420 117.185 122.830 117.805 ;
        RECT 123.000 117.015 123.170 117.985 ;
        RECT 122.475 116.845 123.170 117.015 ;
        RECT 120.790 116.175 121.170 116.555 ;
        RECT 121.410 116.390 122.240 116.560 ;
        RECT 122.475 116.345 122.645 116.845 ;
        RECT 122.815 116.175 123.145 116.675 ;
        RECT 123.360 116.345 123.585 118.465 ;
        RECT 123.755 118.345 124.085 118.725 ;
        RECT 124.255 118.175 124.425 118.465 ;
        RECT 123.760 118.005 124.425 118.175 ;
        RECT 123.760 117.015 123.990 118.005 ;
        RECT 124.685 117.955 126.355 118.725 ;
        RECT 126.525 117.975 127.735 118.725 ;
        RECT 124.160 117.185 124.510 117.835 ;
        RECT 124.685 117.265 125.435 117.785 ;
        RECT 125.605 117.435 126.355 117.955 ;
        RECT 126.525 117.265 127.045 117.805 ;
        RECT 127.215 117.435 127.735 117.975 ;
        RECT 123.760 116.845 124.425 117.015 ;
        RECT 123.755 116.175 124.085 116.675 ;
        RECT 124.255 116.345 124.425 116.845 ;
        RECT 124.685 116.175 126.355 117.265 ;
        RECT 126.525 116.175 127.735 117.265 ;
        RECT 14.660 116.005 127.820 116.175 ;
        RECT 14.745 114.915 15.955 116.005 ;
        RECT 17.050 115.570 22.395 116.005 ;
        RECT 14.745 114.205 15.265 114.745 ;
        RECT 15.435 114.375 15.955 114.915 ;
        RECT 18.640 114.320 18.990 115.570 ;
        RECT 22.605 114.865 22.835 116.005 ;
        RECT 23.005 114.855 23.335 115.835 ;
        RECT 23.505 114.865 23.715 116.005 ;
        RECT 14.745 113.455 15.955 114.205 ;
        RECT 20.470 114.000 20.810 114.830 ;
        RECT 22.585 114.445 22.915 114.695 ;
        RECT 17.050 113.455 22.395 114.000 ;
        RECT 22.605 113.455 22.835 114.275 ;
        RECT 23.085 114.255 23.335 114.855 ;
        RECT 24.405 114.840 24.695 116.005 ;
        RECT 24.905 114.865 25.135 116.005 ;
        RECT 25.305 114.855 25.635 115.835 ;
        RECT 25.805 114.865 26.015 116.005 ;
        RECT 26.705 114.930 26.975 115.835 ;
        RECT 27.145 115.245 27.475 116.005 ;
        RECT 27.655 115.075 27.825 115.835 ;
        RECT 24.885 114.445 25.215 114.695 ;
        RECT 23.005 113.625 23.335 114.255 ;
        RECT 23.505 113.455 23.715 114.275 ;
        RECT 24.405 113.455 24.695 114.180 ;
        RECT 24.905 113.455 25.135 114.275 ;
        RECT 25.385 114.255 25.635 114.855 ;
        RECT 25.305 113.625 25.635 114.255 ;
        RECT 25.805 113.455 26.015 114.275 ;
        RECT 26.705 114.130 26.875 114.930 ;
        RECT 27.160 114.905 27.825 115.075 ;
        RECT 28.545 114.915 32.055 116.005 ;
        RECT 32.600 115.665 32.855 115.695 ;
        RECT 32.515 115.495 32.855 115.665 ;
        RECT 32.600 115.025 32.855 115.495 ;
        RECT 33.035 115.205 33.320 116.005 ;
        RECT 33.500 115.285 33.830 115.795 ;
        RECT 27.160 114.760 27.330 114.905 ;
        RECT 27.045 114.430 27.330 114.760 ;
        RECT 27.160 114.175 27.330 114.430 ;
        RECT 27.565 114.355 27.895 114.725 ;
        RECT 28.545 114.395 30.235 114.915 ;
        RECT 30.405 114.225 32.055 114.745 ;
        RECT 26.705 113.625 26.965 114.130 ;
        RECT 27.160 114.005 27.825 114.175 ;
        RECT 27.145 113.455 27.475 113.835 ;
        RECT 27.655 113.625 27.825 114.005 ;
        RECT 28.545 113.455 32.055 114.225 ;
        RECT 32.600 114.165 32.780 115.025 ;
        RECT 33.500 114.695 33.750 115.285 ;
        RECT 34.100 115.135 34.270 115.745 ;
        RECT 34.440 115.315 34.770 116.005 ;
        RECT 35.000 115.455 35.240 115.745 ;
        RECT 35.440 115.625 35.860 116.005 ;
        RECT 36.040 115.535 36.670 115.785 ;
        RECT 37.140 115.625 37.470 116.005 ;
        RECT 36.040 115.455 36.210 115.535 ;
        RECT 37.640 115.455 37.810 115.745 ;
        RECT 37.990 115.625 38.370 116.005 ;
        RECT 38.610 115.620 39.440 115.790 ;
        RECT 35.000 115.285 36.210 115.455 ;
        RECT 32.950 114.365 33.750 114.695 ;
        RECT 32.600 113.635 32.855 114.165 ;
        RECT 33.035 113.455 33.320 113.915 ;
        RECT 33.500 113.715 33.750 114.365 ;
        RECT 33.950 115.115 34.270 115.135 ;
        RECT 33.950 114.945 35.870 115.115 ;
        RECT 33.950 114.050 34.140 114.945 ;
        RECT 36.040 114.775 36.210 115.285 ;
        RECT 36.380 115.025 36.900 115.335 ;
        RECT 34.310 114.605 36.210 114.775 ;
        RECT 34.310 114.545 34.640 114.605 ;
        RECT 34.790 114.375 35.120 114.435 ;
        RECT 34.460 114.105 35.120 114.375 ;
        RECT 33.950 113.720 34.270 114.050 ;
        RECT 34.450 113.455 35.110 113.935 ;
        RECT 35.310 113.845 35.480 114.605 ;
        RECT 36.380 114.435 36.560 114.845 ;
        RECT 35.650 114.265 35.980 114.385 ;
        RECT 36.730 114.265 36.900 115.025 ;
        RECT 35.650 114.095 36.900 114.265 ;
        RECT 37.070 115.205 38.440 115.455 ;
        RECT 37.070 114.435 37.260 115.205 ;
        RECT 38.190 114.945 38.440 115.205 ;
        RECT 37.430 114.775 37.680 114.935 ;
        RECT 38.610 114.775 38.780 115.620 ;
        RECT 39.675 115.335 39.845 115.835 ;
        RECT 40.015 115.505 40.345 116.005 ;
        RECT 38.950 114.945 39.450 115.325 ;
        RECT 39.675 115.165 40.370 115.335 ;
        RECT 37.430 114.605 38.780 114.775 ;
        RECT 38.360 114.565 38.780 114.605 ;
        RECT 37.070 114.095 37.490 114.435 ;
        RECT 37.780 114.105 38.190 114.435 ;
        RECT 35.310 113.675 36.160 113.845 ;
        RECT 36.720 113.455 37.040 113.915 ;
        RECT 37.240 113.665 37.490 114.095 ;
        RECT 37.780 113.455 38.190 113.895 ;
        RECT 38.360 113.835 38.530 114.565 ;
        RECT 38.700 114.015 39.050 114.385 ;
        RECT 39.230 114.075 39.450 114.945 ;
        RECT 39.620 114.375 40.030 114.995 ;
        RECT 40.200 114.195 40.370 115.165 ;
        RECT 39.675 114.005 40.370 114.195 ;
        RECT 38.360 113.635 39.375 113.835 ;
        RECT 39.675 113.675 39.845 114.005 ;
        RECT 40.015 113.455 40.345 113.835 ;
        RECT 40.560 113.715 40.785 115.835 ;
        RECT 40.955 115.505 41.285 116.005 ;
        RECT 41.455 115.335 41.625 115.835 ;
        RECT 40.960 115.165 41.625 115.335 ;
        RECT 40.960 114.175 41.190 115.165 ;
        RECT 41.360 114.345 41.710 114.995 ;
        RECT 41.885 114.915 44.475 116.005 ;
        RECT 44.650 115.570 49.995 116.005 ;
        RECT 41.885 114.395 43.095 114.915 ;
        RECT 43.265 114.225 44.475 114.745 ;
        RECT 46.240 114.320 46.590 115.570 ;
        RECT 50.165 114.840 50.455 116.005 ;
        RECT 51.145 114.865 51.355 116.005 ;
        RECT 51.525 114.855 51.855 115.835 ;
        RECT 52.025 114.865 52.255 116.005 ;
        RECT 52.505 114.865 52.735 116.005 ;
        RECT 52.905 114.855 53.235 115.835 ;
        RECT 53.405 114.865 53.615 116.005 ;
        RECT 53.845 114.930 54.115 115.835 ;
        RECT 54.285 115.245 54.615 116.005 ;
        RECT 54.795 115.075 54.965 115.835 ;
        RECT 40.960 114.005 41.625 114.175 ;
        RECT 40.955 113.455 41.285 113.835 ;
        RECT 41.455 113.715 41.625 114.005 ;
        RECT 41.885 113.455 44.475 114.225 ;
        RECT 48.070 114.000 48.410 114.830 ;
        RECT 44.650 113.455 49.995 114.000 ;
        RECT 50.165 113.455 50.455 114.180 ;
        RECT 51.145 113.455 51.355 114.275 ;
        RECT 51.525 114.255 51.775 114.855 ;
        RECT 51.945 114.445 52.275 114.695 ;
        RECT 52.485 114.445 52.815 114.695 ;
        RECT 51.525 113.625 51.855 114.255 ;
        RECT 52.025 113.455 52.255 114.275 ;
        RECT 52.505 113.455 52.735 114.275 ;
        RECT 52.985 114.255 53.235 114.855 ;
        RECT 52.905 113.625 53.235 114.255 ;
        RECT 53.405 113.455 53.615 114.275 ;
        RECT 53.845 114.130 54.015 114.930 ;
        RECT 54.300 114.905 54.965 115.075 ;
        RECT 55.775 115.075 55.945 115.835 ;
        RECT 56.125 115.245 56.455 116.005 ;
        RECT 55.775 114.905 56.440 115.075 ;
        RECT 56.625 114.930 56.895 115.835 ;
        RECT 54.300 114.760 54.470 114.905 ;
        RECT 54.185 114.430 54.470 114.760 ;
        RECT 56.270 114.760 56.440 114.905 ;
        RECT 54.300 114.175 54.470 114.430 ;
        RECT 54.705 114.355 55.035 114.725 ;
        RECT 55.705 114.355 56.035 114.725 ;
        RECT 56.270 114.430 56.555 114.760 ;
        RECT 56.270 114.175 56.440 114.430 ;
        RECT 53.845 113.625 54.105 114.130 ;
        RECT 54.300 114.005 54.965 114.175 ;
        RECT 54.285 113.455 54.615 113.835 ;
        RECT 54.795 113.625 54.965 114.005 ;
        RECT 55.775 114.005 56.440 114.175 ;
        RECT 56.725 114.130 56.895 114.930 ;
        RECT 57.525 114.915 61.035 116.005 ;
        RECT 57.525 114.395 59.215 114.915 ;
        RECT 61.245 114.865 61.475 116.005 ;
        RECT 61.645 114.855 61.975 115.835 ;
        RECT 62.145 114.865 62.355 116.005 ;
        RECT 62.960 115.665 63.215 115.695 ;
        RECT 62.875 115.495 63.215 115.665 ;
        RECT 62.960 115.025 63.215 115.495 ;
        RECT 63.395 115.205 63.680 116.005 ;
        RECT 63.860 115.285 64.190 115.795 ;
        RECT 59.385 114.225 61.035 114.745 ;
        RECT 61.225 114.445 61.555 114.695 ;
        RECT 55.775 113.625 55.945 114.005 ;
        RECT 56.125 113.455 56.455 113.835 ;
        RECT 56.635 113.625 56.895 114.130 ;
        RECT 57.525 113.455 61.035 114.225 ;
        RECT 61.245 113.455 61.475 114.275 ;
        RECT 61.725 114.255 61.975 114.855 ;
        RECT 61.645 113.625 61.975 114.255 ;
        RECT 62.145 113.455 62.355 114.275 ;
        RECT 62.960 114.165 63.140 115.025 ;
        RECT 63.860 114.695 64.110 115.285 ;
        RECT 64.460 115.135 64.630 115.745 ;
        RECT 64.800 115.315 65.130 116.005 ;
        RECT 65.360 115.455 65.600 115.745 ;
        RECT 65.800 115.625 66.220 116.005 ;
        RECT 66.400 115.535 67.030 115.785 ;
        RECT 67.500 115.625 67.830 116.005 ;
        RECT 66.400 115.455 66.570 115.535 ;
        RECT 68.000 115.455 68.170 115.745 ;
        RECT 68.350 115.625 68.730 116.005 ;
        RECT 68.970 115.620 69.800 115.790 ;
        RECT 65.360 115.285 66.570 115.455 ;
        RECT 63.310 114.365 64.110 114.695 ;
        RECT 62.960 113.635 63.215 114.165 ;
        RECT 63.395 113.455 63.680 113.915 ;
        RECT 63.860 113.715 64.110 114.365 ;
        RECT 64.310 115.115 64.630 115.135 ;
        RECT 64.310 114.945 66.230 115.115 ;
        RECT 64.310 114.050 64.500 114.945 ;
        RECT 66.400 114.775 66.570 115.285 ;
        RECT 66.740 115.025 67.260 115.335 ;
        RECT 64.670 114.605 66.570 114.775 ;
        RECT 64.670 114.545 65.000 114.605 ;
        RECT 65.150 114.375 65.480 114.435 ;
        RECT 64.820 114.105 65.480 114.375 ;
        RECT 64.310 113.720 64.630 114.050 ;
        RECT 64.810 113.455 65.470 113.935 ;
        RECT 65.670 113.845 65.840 114.605 ;
        RECT 66.740 114.435 66.920 114.845 ;
        RECT 66.010 114.265 66.340 114.385 ;
        RECT 67.090 114.265 67.260 115.025 ;
        RECT 66.010 114.095 67.260 114.265 ;
        RECT 67.430 115.205 68.800 115.455 ;
        RECT 67.430 114.435 67.620 115.205 ;
        RECT 68.550 114.945 68.800 115.205 ;
        RECT 67.790 114.775 68.040 114.935 ;
        RECT 68.970 114.775 69.140 115.620 ;
        RECT 70.035 115.335 70.205 115.835 ;
        RECT 70.375 115.505 70.705 116.005 ;
        RECT 69.310 114.945 69.810 115.325 ;
        RECT 70.035 115.165 70.730 115.335 ;
        RECT 67.790 114.605 69.140 114.775 ;
        RECT 68.720 114.565 69.140 114.605 ;
        RECT 67.430 114.095 67.850 114.435 ;
        RECT 68.140 114.105 68.550 114.435 ;
        RECT 65.670 113.675 66.520 113.845 ;
        RECT 67.080 113.455 67.400 113.915 ;
        RECT 67.600 113.665 67.850 114.095 ;
        RECT 68.140 113.455 68.550 113.895 ;
        RECT 68.720 113.835 68.890 114.565 ;
        RECT 69.060 114.015 69.410 114.385 ;
        RECT 69.590 114.075 69.810 114.945 ;
        RECT 69.980 114.375 70.390 114.995 ;
        RECT 70.560 114.195 70.730 115.165 ;
        RECT 70.035 114.005 70.730 114.195 ;
        RECT 68.720 113.635 69.735 113.835 ;
        RECT 70.035 113.675 70.205 114.005 ;
        RECT 70.375 113.455 70.705 113.835 ;
        RECT 70.920 113.715 71.145 115.835 ;
        RECT 71.315 115.505 71.645 116.005 ;
        RECT 71.815 115.335 71.985 115.835 ;
        RECT 71.320 115.165 71.985 115.335 ;
        RECT 71.320 114.175 71.550 115.165 ;
        RECT 71.720 114.345 72.070 114.995 ;
        RECT 72.305 114.865 72.515 116.005 ;
        RECT 72.685 114.855 73.015 115.835 ;
        RECT 73.185 114.865 73.415 116.005 ;
        RECT 74.085 114.915 75.755 116.005 ;
        RECT 71.320 114.005 71.985 114.175 ;
        RECT 71.315 113.455 71.645 113.835 ;
        RECT 71.815 113.715 71.985 114.005 ;
        RECT 72.305 113.455 72.515 114.275 ;
        RECT 72.685 114.255 72.935 114.855 ;
        RECT 73.105 114.445 73.435 114.695 ;
        RECT 74.085 114.395 74.835 114.915 ;
        RECT 75.925 114.840 76.215 116.005 ;
        RECT 76.845 114.915 79.435 116.005 ;
        RECT 72.685 113.625 73.015 114.255 ;
        RECT 73.185 113.455 73.415 114.275 ;
        RECT 75.005 114.225 75.755 114.745 ;
        RECT 76.845 114.395 78.055 114.915 ;
        RECT 79.645 114.865 79.875 116.005 ;
        RECT 80.045 114.855 80.375 115.835 ;
        RECT 80.545 114.865 80.755 116.005 ;
        RECT 80.985 114.915 82.655 116.005 ;
        RECT 82.915 115.075 83.085 115.835 ;
        RECT 83.265 115.245 83.595 116.005 ;
        RECT 78.225 114.225 79.435 114.745 ;
        RECT 79.625 114.445 79.955 114.695 ;
        RECT 74.085 113.455 75.755 114.225 ;
        RECT 75.925 113.455 76.215 114.180 ;
        RECT 76.845 113.455 79.435 114.225 ;
        RECT 79.645 113.455 79.875 114.275 ;
        RECT 80.125 114.255 80.375 114.855 ;
        RECT 80.985 114.395 81.735 114.915 ;
        RECT 82.915 114.905 83.580 115.075 ;
        RECT 83.765 114.930 84.035 115.835 ;
        RECT 83.410 114.760 83.580 114.905 ;
        RECT 80.045 113.625 80.375 114.255 ;
        RECT 80.545 113.455 80.755 114.275 ;
        RECT 81.905 114.225 82.655 114.745 ;
        RECT 82.845 114.355 83.175 114.725 ;
        RECT 83.410 114.430 83.695 114.760 ;
        RECT 80.985 113.455 82.655 114.225 ;
        RECT 83.410 114.175 83.580 114.430 ;
        RECT 82.915 114.005 83.580 114.175 ;
        RECT 83.865 114.130 84.035 114.930 ;
        RECT 84.205 114.915 87.715 116.005 ;
        RECT 88.260 115.665 88.515 115.695 ;
        RECT 88.175 115.495 88.515 115.665 ;
        RECT 88.260 115.025 88.515 115.495 ;
        RECT 88.695 115.205 88.980 116.005 ;
        RECT 89.160 115.285 89.490 115.795 ;
        RECT 84.205 114.395 85.895 114.915 ;
        RECT 86.065 114.225 87.715 114.745 ;
        RECT 82.915 113.625 83.085 114.005 ;
        RECT 83.265 113.455 83.595 113.835 ;
        RECT 83.775 113.625 84.035 114.130 ;
        RECT 84.205 113.455 87.715 114.225 ;
        RECT 88.260 114.165 88.440 115.025 ;
        RECT 89.160 114.695 89.410 115.285 ;
        RECT 89.760 115.135 89.930 115.745 ;
        RECT 90.100 115.315 90.430 116.005 ;
        RECT 90.660 115.455 90.900 115.745 ;
        RECT 91.100 115.625 91.520 116.005 ;
        RECT 91.700 115.535 92.330 115.785 ;
        RECT 92.800 115.625 93.130 116.005 ;
        RECT 91.700 115.455 91.870 115.535 ;
        RECT 93.300 115.455 93.470 115.745 ;
        RECT 93.650 115.625 94.030 116.005 ;
        RECT 94.270 115.620 95.100 115.790 ;
        RECT 90.660 115.285 91.870 115.455 ;
        RECT 88.610 114.365 89.410 114.695 ;
        RECT 88.260 113.635 88.515 114.165 ;
        RECT 88.695 113.455 88.980 113.915 ;
        RECT 89.160 113.715 89.410 114.365 ;
        RECT 89.610 115.115 89.930 115.135 ;
        RECT 89.610 114.945 91.530 115.115 ;
        RECT 89.610 114.050 89.800 114.945 ;
        RECT 91.700 114.775 91.870 115.285 ;
        RECT 92.040 115.025 92.560 115.335 ;
        RECT 89.970 114.605 91.870 114.775 ;
        RECT 89.970 114.545 90.300 114.605 ;
        RECT 90.450 114.375 90.780 114.435 ;
        RECT 90.120 114.105 90.780 114.375 ;
        RECT 89.610 113.720 89.930 114.050 ;
        RECT 90.110 113.455 90.770 113.935 ;
        RECT 90.970 113.845 91.140 114.605 ;
        RECT 92.040 114.435 92.220 114.845 ;
        RECT 91.310 114.265 91.640 114.385 ;
        RECT 92.390 114.265 92.560 115.025 ;
        RECT 91.310 114.095 92.560 114.265 ;
        RECT 92.730 115.205 94.100 115.455 ;
        RECT 92.730 114.435 92.920 115.205 ;
        RECT 93.850 114.945 94.100 115.205 ;
        RECT 93.090 114.775 93.340 114.935 ;
        RECT 94.270 114.775 94.440 115.620 ;
        RECT 95.335 115.335 95.505 115.835 ;
        RECT 95.675 115.505 96.005 116.005 ;
        RECT 94.610 114.945 95.110 115.325 ;
        RECT 95.335 115.165 96.030 115.335 ;
        RECT 93.090 114.605 94.440 114.775 ;
        RECT 94.020 114.565 94.440 114.605 ;
        RECT 92.730 114.095 93.150 114.435 ;
        RECT 93.440 114.105 93.850 114.435 ;
        RECT 90.970 113.675 91.820 113.845 ;
        RECT 92.380 113.455 92.700 113.915 ;
        RECT 92.900 113.665 93.150 114.095 ;
        RECT 93.440 113.455 93.850 113.895 ;
        RECT 94.020 113.835 94.190 114.565 ;
        RECT 94.360 114.015 94.710 114.385 ;
        RECT 94.890 114.075 95.110 114.945 ;
        RECT 95.280 114.375 95.690 114.995 ;
        RECT 95.860 114.195 96.030 115.165 ;
        RECT 95.335 114.005 96.030 114.195 ;
        RECT 94.020 113.635 95.035 113.835 ;
        RECT 95.335 113.675 95.505 114.005 ;
        RECT 95.675 113.455 96.005 113.835 ;
        RECT 96.220 113.715 96.445 115.835 ;
        RECT 96.615 115.505 96.945 116.005 ;
        RECT 97.115 115.335 97.285 115.835 ;
        RECT 96.620 115.165 97.285 115.335 ;
        RECT 96.620 114.175 96.850 115.165 ;
        RECT 97.020 114.345 97.370 114.995 ;
        RECT 98.005 114.915 101.515 116.005 ;
        RECT 98.005 114.395 99.695 114.915 ;
        RECT 101.685 114.840 101.975 116.005 ;
        RECT 102.605 114.915 104.275 116.005 ;
        RECT 104.820 115.665 105.075 115.695 ;
        RECT 104.735 115.495 105.075 115.665 ;
        RECT 104.820 115.025 105.075 115.495 ;
        RECT 105.255 115.205 105.540 116.005 ;
        RECT 105.720 115.285 106.050 115.795 ;
        RECT 99.865 114.225 101.515 114.745 ;
        RECT 102.605 114.395 103.355 114.915 ;
        RECT 103.525 114.225 104.275 114.745 ;
        RECT 96.620 114.005 97.285 114.175 ;
        RECT 96.615 113.455 96.945 113.835 ;
        RECT 97.115 113.715 97.285 114.005 ;
        RECT 98.005 113.455 101.515 114.225 ;
        RECT 101.685 113.455 101.975 114.180 ;
        RECT 102.605 113.455 104.275 114.225 ;
        RECT 104.820 114.165 105.000 115.025 ;
        RECT 105.720 114.695 105.970 115.285 ;
        RECT 106.320 115.135 106.490 115.745 ;
        RECT 106.660 115.315 106.990 116.005 ;
        RECT 107.220 115.455 107.460 115.745 ;
        RECT 107.660 115.625 108.080 116.005 ;
        RECT 108.260 115.535 108.890 115.785 ;
        RECT 109.360 115.625 109.690 116.005 ;
        RECT 108.260 115.455 108.430 115.535 ;
        RECT 109.860 115.455 110.030 115.745 ;
        RECT 110.210 115.625 110.590 116.005 ;
        RECT 110.830 115.620 111.660 115.790 ;
        RECT 107.220 115.285 108.430 115.455 ;
        RECT 105.170 114.365 105.970 114.695 ;
        RECT 104.820 113.635 105.075 114.165 ;
        RECT 105.255 113.455 105.540 113.915 ;
        RECT 105.720 113.715 105.970 114.365 ;
        RECT 106.170 115.115 106.490 115.135 ;
        RECT 106.170 114.945 108.090 115.115 ;
        RECT 106.170 114.050 106.360 114.945 ;
        RECT 108.260 114.775 108.430 115.285 ;
        RECT 108.600 115.025 109.120 115.335 ;
        RECT 106.530 114.605 108.430 114.775 ;
        RECT 106.530 114.545 106.860 114.605 ;
        RECT 107.010 114.375 107.340 114.435 ;
        RECT 106.680 114.105 107.340 114.375 ;
        RECT 106.170 113.720 106.490 114.050 ;
        RECT 106.670 113.455 107.330 113.935 ;
        RECT 107.530 113.845 107.700 114.605 ;
        RECT 108.600 114.435 108.780 114.845 ;
        RECT 107.870 114.265 108.200 114.385 ;
        RECT 108.950 114.265 109.120 115.025 ;
        RECT 107.870 114.095 109.120 114.265 ;
        RECT 109.290 115.205 110.660 115.455 ;
        RECT 109.290 114.435 109.480 115.205 ;
        RECT 110.410 114.945 110.660 115.205 ;
        RECT 109.650 114.775 109.900 114.935 ;
        RECT 110.830 114.775 111.000 115.620 ;
        RECT 111.895 115.335 112.065 115.835 ;
        RECT 112.235 115.505 112.565 116.005 ;
        RECT 111.170 114.945 111.670 115.325 ;
        RECT 111.895 115.165 112.590 115.335 ;
        RECT 109.650 114.605 111.000 114.775 ;
        RECT 110.580 114.565 111.000 114.605 ;
        RECT 109.290 114.095 109.710 114.435 ;
        RECT 110.000 114.105 110.410 114.435 ;
        RECT 107.530 113.675 108.380 113.845 ;
        RECT 108.940 113.455 109.260 113.915 ;
        RECT 109.460 113.665 109.710 114.095 ;
        RECT 110.000 113.455 110.410 113.895 ;
        RECT 110.580 113.835 110.750 114.565 ;
        RECT 110.920 114.015 111.270 114.385 ;
        RECT 111.450 114.075 111.670 114.945 ;
        RECT 111.840 114.375 112.250 114.995 ;
        RECT 112.420 114.195 112.590 115.165 ;
        RECT 111.895 114.005 112.590 114.195 ;
        RECT 110.580 113.635 111.595 113.835 ;
        RECT 111.895 113.675 112.065 114.005 ;
        RECT 112.235 113.455 112.565 113.835 ;
        RECT 112.780 113.715 113.005 115.835 ;
        RECT 113.175 115.505 113.505 116.005 ;
        RECT 113.675 115.335 113.845 115.835 ;
        RECT 113.180 115.165 113.845 115.335 ;
        RECT 113.180 114.175 113.410 115.165 ;
        RECT 113.580 114.345 113.930 114.995 ;
        RECT 114.105 114.915 115.315 116.005 ;
        RECT 115.490 115.570 120.835 116.005 ;
        RECT 121.010 115.570 126.355 116.005 ;
        RECT 114.105 114.375 114.625 114.915 ;
        RECT 114.795 114.205 115.315 114.745 ;
        RECT 117.080 114.320 117.430 115.570 ;
        RECT 113.180 114.005 113.845 114.175 ;
        RECT 113.175 113.455 113.505 113.835 ;
        RECT 113.675 113.715 113.845 114.005 ;
        RECT 114.105 113.455 115.315 114.205 ;
        RECT 118.910 114.000 119.250 114.830 ;
        RECT 122.600 114.320 122.950 115.570 ;
        RECT 126.525 114.915 127.735 116.005 ;
        RECT 124.430 114.000 124.770 114.830 ;
        RECT 126.525 114.375 127.045 114.915 ;
        RECT 127.215 114.205 127.735 114.745 ;
        RECT 115.490 113.455 120.835 114.000 ;
        RECT 121.010 113.455 126.355 114.000 ;
        RECT 126.525 113.455 127.735 114.205 ;
        RECT 14.660 113.285 127.820 113.455 ;
        RECT 14.745 112.535 15.955 113.285 ;
        RECT 14.745 111.995 15.265 112.535 ;
        RECT 16.585 112.515 18.255 113.285 ;
        RECT 18.735 112.815 18.905 113.285 ;
        RECT 19.075 112.635 19.405 113.115 ;
        RECT 19.575 112.815 19.745 113.285 ;
        RECT 19.915 112.635 20.245 113.115 ;
        RECT 15.435 111.825 15.955 112.365 ;
        RECT 14.745 110.735 15.955 111.825 ;
        RECT 16.585 111.825 17.335 112.345 ;
        RECT 17.505 111.995 18.255 112.515 ;
        RECT 18.480 112.465 20.245 112.635 ;
        RECT 20.415 112.475 20.585 113.285 ;
        RECT 20.785 112.905 21.855 113.075 ;
        RECT 20.785 112.550 21.105 112.905 ;
        RECT 18.480 111.915 18.890 112.465 ;
        RECT 20.780 112.295 21.105 112.550 ;
        RECT 19.075 112.085 21.105 112.295 ;
        RECT 20.760 112.075 21.105 112.085 ;
        RECT 21.275 112.335 21.515 112.735 ;
        RECT 21.685 112.675 21.855 112.905 ;
        RECT 22.025 112.845 22.215 113.285 ;
        RECT 22.385 112.835 23.335 113.115 ;
        RECT 23.555 112.925 23.905 113.095 ;
        RECT 21.685 112.505 22.215 112.675 ;
        RECT 16.585 110.735 18.255 111.825 ;
        RECT 18.480 111.745 20.205 111.915 ;
        RECT 18.735 110.735 18.905 111.575 ;
        RECT 19.115 110.905 19.365 111.745 ;
        RECT 19.575 110.735 19.745 111.575 ;
        RECT 19.915 110.905 20.205 111.745 ;
        RECT 20.415 110.735 20.585 111.795 ;
        RECT 20.760 111.455 20.930 112.075 ;
        RECT 21.275 111.965 21.815 112.335 ;
        RECT 21.995 112.225 22.215 112.505 ;
        RECT 22.385 112.055 22.555 112.835 ;
        RECT 22.150 111.885 22.555 112.055 ;
        RECT 22.725 112.045 23.075 112.665 ;
        RECT 22.150 111.795 22.320 111.885 ;
        RECT 23.245 111.875 23.455 112.665 ;
        RECT 21.100 111.625 22.320 111.795 ;
        RECT 22.780 111.715 23.455 111.875 ;
        RECT 20.760 111.285 21.560 111.455 ;
        RECT 20.880 110.735 21.210 111.115 ;
        RECT 21.390 110.995 21.560 111.285 ;
        RECT 22.150 111.245 22.320 111.625 ;
        RECT 22.490 111.705 23.455 111.715 ;
        RECT 23.645 112.535 23.905 112.925 ;
        RECT 24.115 112.825 24.445 113.285 ;
        RECT 25.320 112.895 26.175 113.065 ;
        RECT 26.380 112.895 26.875 113.065 ;
        RECT 27.045 112.925 27.375 113.285 ;
        RECT 23.645 111.845 23.815 112.535 ;
        RECT 23.985 112.185 24.155 112.365 ;
        RECT 24.325 112.355 25.115 112.605 ;
        RECT 25.320 112.185 25.490 112.895 ;
        RECT 25.660 112.385 26.015 112.605 ;
        RECT 23.985 112.015 25.675 112.185 ;
        RECT 22.490 111.415 22.950 111.705 ;
        RECT 23.645 111.675 25.145 111.845 ;
        RECT 23.645 111.535 23.815 111.675 ;
        RECT 23.255 111.365 23.815 111.535 ;
        RECT 21.730 110.735 21.980 111.195 ;
        RECT 22.150 110.905 23.020 111.245 ;
        RECT 23.255 110.905 23.425 111.365 ;
        RECT 24.260 111.335 25.335 111.505 ;
        RECT 23.595 110.735 23.965 111.195 ;
        RECT 24.260 110.995 24.430 111.335 ;
        RECT 24.600 110.735 24.930 111.165 ;
        RECT 25.165 110.995 25.335 111.335 ;
        RECT 25.505 111.235 25.675 112.015 ;
        RECT 25.845 111.795 26.015 112.385 ;
        RECT 26.185 111.985 26.535 112.605 ;
        RECT 25.845 111.405 26.310 111.795 ;
        RECT 26.705 111.535 26.875 112.895 ;
        RECT 27.045 111.705 27.505 112.755 ;
        RECT 26.480 111.365 26.875 111.535 ;
        RECT 26.480 111.235 26.650 111.365 ;
        RECT 25.505 110.905 26.185 111.235 ;
        RECT 26.400 110.905 26.650 111.235 ;
        RECT 26.820 110.735 27.070 111.195 ;
        RECT 27.240 110.920 27.565 111.705 ;
        RECT 27.735 110.905 27.905 113.025 ;
        RECT 28.075 112.905 28.405 113.285 ;
        RECT 28.575 112.735 28.830 113.025 ;
        RECT 28.080 112.565 28.830 112.735 ;
        RECT 28.080 111.575 28.310 112.565 ;
        RECT 29.005 112.535 30.215 113.285 ;
        RECT 28.480 111.745 28.830 112.395 ;
        RECT 29.005 111.825 29.525 112.365 ;
        RECT 29.695 111.995 30.215 112.535 ;
        RECT 30.385 112.515 33.895 113.285 ;
        RECT 30.385 111.825 32.075 112.345 ;
        RECT 32.245 111.995 33.895 112.515 ;
        RECT 34.125 112.465 34.335 113.285 ;
        RECT 34.505 112.485 34.835 113.115 ;
        RECT 34.505 111.885 34.755 112.485 ;
        RECT 35.005 112.465 35.235 113.285 ;
        RECT 35.905 112.610 36.165 113.115 ;
        RECT 36.345 112.905 36.675 113.285 ;
        RECT 36.855 112.735 37.025 113.115 ;
        RECT 34.925 112.045 35.255 112.295 ;
        RECT 28.080 111.405 28.830 111.575 ;
        RECT 28.075 110.735 28.405 111.235 ;
        RECT 28.575 110.905 28.830 111.405 ;
        RECT 29.005 110.735 30.215 111.825 ;
        RECT 30.385 110.735 33.895 111.825 ;
        RECT 34.125 110.735 34.335 111.875 ;
        RECT 34.505 110.905 34.835 111.885 ;
        RECT 35.005 110.735 35.235 111.875 ;
        RECT 35.905 111.810 36.075 112.610 ;
        RECT 36.360 112.565 37.025 112.735 ;
        RECT 36.360 112.310 36.530 112.565 ;
        RECT 37.285 112.560 37.575 113.285 ;
        RECT 37.750 112.740 43.095 113.285 ;
        RECT 36.245 111.980 36.530 112.310 ;
        RECT 36.765 112.015 37.095 112.385 ;
        RECT 36.360 111.835 36.530 111.980 ;
        RECT 35.905 110.905 36.175 111.810 ;
        RECT 36.360 111.665 37.025 111.835 ;
        RECT 36.345 110.735 36.675 111.495 ;
        RECT 36.855 110.905 37.025 111.665 ;
        RECT 37.285 110.735 37.575 111.900 ;
        RECT 39.340 111.170 39.690 112.420 ;
        RECT 41.170 111.910 41.510 112.740 ;
        RECT 43.265 112.610 43.525 113.115 ;
        RECT 43.705 112.905 44.035 113.285 ;
        RECT 44.215 112.735 44.385 113.115 ;
        RECT 43.265 111.810 43.435 112.610 ;
        RECT 43.720 112.565 44.385 112.735 ;
        RECT 45.655 112.735 45.825 113.115 ;
        RECT 46.005 112.905 46.335 113.285 ;
        RECT 45.655 112.565 46.320 112.735 ;
        RECT 46.515 112.610 46.775 113.115 ;
        RECT 43.720 112.310 43.890 112.565 ;
        RECT 43.605 111.980 43.890 112.310 ;
        RECT 44.125 112.015 44.455 112.385 ;
        RECT 45.585 112.015 45.915 112.385 ;
        RECT 46.150 112.310 46.320 112.565 ;
        RECT 43.720 111.835 43.890 111.980 ;
        RECT 46.150 111.980 46.435 112.310 ;
        RECT 46.150 111.835 46.320 111.980 ;
        RECT 37.750 110.735 43.095 111.170 ;
        RECT 43.265 110.905 43.535 111.810 ;
        RECT 43.720 111.665 44.385 111.835 ;
        RECT 43.705 110.735 44.035 111.495 ;
        RECT 44.215 110.905 44.385 111.665 ;
        RECT 45.655 111.665 46.320 111.835 ;
        RECT 46.605 111.810 46.775 112.610 ;
        RECT 46.945 112.535 48.155 113.285 ;
        RECT 45.655 110.905 45.825 111.665 ;
        RECT 46.005 110.735 46.335 111.495 ;
        RECT 46.505 110.905 46.775 111.810 ;
        RECT 46.945 111.825 47.465 112.365 ;
        RECT 47.635 111.995 48.155 112.535 ;
        RECT 48.325 112.515 51.835 113.285 ;
        RECT 52.010 112.740 57.355 113.285 ;
        RECT 57.530 112.740 62.875 113.285 ;
        RECT 48.325 111.825 50.015 112.345 ;
        RECT 50.185 111.995 51.835 112.515 ;
        RECT 46.945 110.735 48.155 111.825 ;
        RECT 48.325 110.735 51.835 111.825 ;
        RECT 53.600 111.170 53.950 112.420 ;
        RECT 55.430 111.910 55.770 112.740 ;
        RECT 59.120 111.170 59.470 112.420 ;
        RECT 60.950 111.910 61.290 112.740 ;
        RECT 63.045 112.560 63.335 113.285 ;
        RECT 63.505 112.535 64.715 113.285 ;
        RECT 52.010 110.735 57.355 111.170 ;
        RECT 57.530 110.735 62.875 111.170 ;
        RECT 63.045 110.735 63.335 111.900 ;
        RECT 63.505 111.825 64.025 112.365 ;
        RECT 64.195 111.995 64.715 112.535 ;
        RECT 65.160 112.475 65.405 113.080 ;
        RECT 65.625 112.750 66.135 113.285 ;
        RECT 64.885 112.305 66.115 112.475 ;
        RECT 63.505 110.735 64.715 111.825 ;
        RECT 64.885 111.495 65.225 112.305 ;
        RECT 65.395 111.740 66.145 111.930 ;
        RECT 64.885 111.085 65.400 111.495 ;
        RECT 65.635 110.735 65.805 111.495 ;
        RECT 65.975 111.075 66.145 111.740 ;
        RECT 66.315 111.755 66.505 113.115 ;
        RECT 66.675 112.605 66.950 113.115 ;
        RECT 67.140 112.750 67.670 113.115 ;
        RECT 68.095 112.885 68.425 113.285 ;
        RECT 67.495 112.715 67.670 112.750 ;
        RECT 66.675 112.435 66.955 112.605 ;
        RECT 66.675 111.955 66.950 112.435 ;
        RECT 67.155 111.755 67.325 112.555 ;
        RECT 66.315 111.585 67.325 111.755 ;
        RECT 67.495 112.545 68.425 112.715 ;
        RECT 68.595 112.545 68.850 113.115 ;
        RECT 69.575 112.735 69.745 113.115 ;
        RECT 69.925 112.905 70.255 113.285 ;
        RECT 69.575 112.565 70.240 112.735 ;
        RECT 70.435 112.610 70.695 113.115 ;
        RECT 67.495 111.415 67.665 112.545 ;
        RECT 68.255 112.375 68.425 112.545 ;
        RECT 66.540 111.245 67.665 111.415 ;
        RECT 67.835 112.045 68.030 112.375 ;
        RECT 68.255 112.045 68.510 112.375 ;
        RECT 67.835 111.075 68.005 112.045 ;
        RECT 68.680 111.875 68.850 112.545 ;
        RECT 69.505 112.015 69.835 112.385 ;
        RECT 70.070 112.310 70.240 112.565 ;
        RECT 65.975 110.905 68.005 111.075 ;
        RECT 68.175 110.735 68.345 111.875 ;
        RECT 68.515 110.905 68.850 111.875 ;
        RECT 70.070 111.980 70.355 112.310 ;
        RECT 70.070 111.835 70.240 111.980 ;
        RECT 69.575 111.665 70.240 111.835 ;
        RECT 70.525 111.810 70.695 112.610 ;
        RECT 71.325 112.515 73.915 113.285 ;
        RECT 74.090 112.740 79.435 113.285 ;
        RECT 69.575 110.905 69.745 111.665 ;
        RECT 69.925 110.735 70.255 111.495 ;
        RECT 70.425 110.905 70.695 111.810 ;
        RECT 71.325 111.825 72.535 112.345 ;
        RECT 72.705 111.995 73.915 112.515 ;
        RECT 71.325 110.735 73.915 111.825 ;
        RECT 75.680 111.170 76.030 112.420 ;
        RECT 77.510 111.910 77.850 112.740 ;
        RECT 79.665 112.465 79.875 113.285 ;
        RECT 80.045 112.485 80.375 113.115 ;
        RECT 80.045 111.885 80.295 112.485 ;
        RECT 80.545 112.465 80.775 113.285 ;
        RECT 81.445 112.515 83.115 113.285 ;
        RECT 83.290 112.740 88.635 113.285 ;
        RECT 80.465 112.045 80.795 112.295 ;
        RECT 74.090 110.735 79.435 111.170 ;
        RECT 79.665 110.735 79.875 111.875 ;
        RECT 80.045 110.905 80.375 111.885 ;
        RECT 80.545 110.735 80.775 111.875 ;
        RECT 81.445 111.825 82.195 112.345 ;
        RECT 82.365 111.995 83.115 112.515 ;
        RECT 81.445 110.735 83.115 111.825 ;
        RECT 84.880 111.170 85.230 112.420 ;
        RECT 86.710 111.910 87.050 112.740 ;
        RECT 88.805 112.560 89.095 113.285 ;
        RECT 89.540 112.475 89.785 113.080 ;
        RECT 90.005 112.750 90.515 113.285 ;
        RECT 89.265 112.305 90.495 112.475 ;
        RECT 83.290 110.735 88.635 111.170 ;
        RECT 88.805 110.735 89.095 111.900 ;
        RECT 89.265 111.495 89.605 112.305 ;
        RECT 89.775 111.740 90.525 111.930 ;
        RECT 89.265 111.085 89.780 111.495 ;
        RECT 90.015 110.735 90.185 111.495 ;
        RECT 90.355 111.075 90.525 111.740 ;
        RECT 90.695 111.755 90.885 113.115 ;
        RECT 91.055 112.605 91.330 113.115 ;
        RECT 91.520 112.750 92.050 113.115 ;
        RECT 92.475 112.885 92.805 113.285 ;
        RECT 91.875 112.715 92.050 112.750 ;
        RECT 91.055 112.435 91.335 112.605 ;
        RECT 91.055 111.955 91.330 112.435 ;
        RECT 91.535 111.755 91.705 112.555 ;
        RECT 90.695 111.585 91.705 111.755 ;
        RECT 91.875 112.545 92.805 112.715 ;
        RECT 92.975 112.545 93.230 113.115 ;
        RECT 93.495 112.735 93.665 113.115 ;
        RECT 93.845 112.905 94.175 113.285 ;
        RECT 93.495 112.565 94.160 112.735 ;
        RECT 94.355 112.610 94.615 113.115 ;
        RECT 91.875 111.415 92.045 112.545 ;
        RECT 92.635 112.375 92.805 112.545 ;
        RECT 90.920 111.245 92.045 111.415 ;
        RECT 92.215 112.045 92.410 112.375 ;
        RECT 92.635 112.045 92.890 112.375 ;
        RECT 92.215 111.075 92.385 112.045 ;
        RECT 93.060 111.875 93.230 112.545 ;
        RECT 93.425 112.015 93.755 112.385 ;
        RECT 93.990 112.310 94.160 112.565 ;
        RECT 90.355 110.905 92.385 111.075 ;
        RECT 92.555 110.735 92.725 111.875 ;
        RECT 92.895 110.905 93.230 111.875 ;
        RECT 93.990 111.980 94.275 112.310 ;
        RECT 93.990 111.835 94.160 111.980 ;
        RECT 93.495 111.665 94.160 111.835 ;
        RECT 94.445 111.810 94.615 112.610 ;
        RECT 94.785 112.515 98.295 113.285 ;
        RECT 98.470 112.740 103.815 113.285 ;
        RECT 103.990 112.740 109.335 113.285 ;
        RECT 93.495 110.905 93.665 111.665 ;
        RECT 93.845 110.735 94.175 111.495 ;
        RECT 94.345 110.905 94.615 111.810 ;
        RECT 94.785 111.825 96.475 112.345 ;
        RECT 96.645 111.995 98.295 112.515 ;
        RECT 94.785 110.735 98.295 111.825 ;
        RECT 100.060 111.170 100.410 112.420 ;
        RECT 101.890 111.910 102.230 112.740 ;
        RECT 105.580 111.170 105.930 112.420 ;
        RECT 107.410 111.910 107.750 112.740 ;
        RECT 109.595 112.735 109.765 113.115 ;
        RECT 109.945 112.905 110.275 113.285 ;
        RECT 109.595 112.565 110.260 112.735 ;
        RECT 110.455 112.610 110.715 113.115 ;
        RECT 109.525 112.015 109.855 112.385 ;
        RECT 110.090 112.310 110.260 112.565 ;
        RECT 110.090 111.980 110.375 112.310 ;
        RECT 110.090 111.835 110.260 111.980 ;
        RECT 109.595 111.665 110.260 111.835 ;
        RECT 110.545 111.810 110.715 112.610 ;
        RECT 110.885 112.515 114.395 113.285 ;
        RECT 114.565 112.560 114.855 113.285 ;
        RECT 115.485 112.515 118.995 113.285 ;
        RECT 98.470 110.735 103.815 111.170 ;
        RECT 103.990 110.735 109.335 111.170 ;
        RECT 109.595 110.905 109.765 111.665 ;
        RECT 109.945 110.735 110.275 111.495 ;
        RECT 110.445 110.905 110.715 111.810 ;
        RECT 110.885 111.825 112.575 112.345 ;
        RECT 112.745 111.995 114.395 112.515 ;
        RECT 110.885 110.735 114.395 111.825 ;
        RECT 114.565 110.735 114.855 111.900 ;
        RECT 115.485 111.825 117.175 112.345 ;
        RECT 117.345 111.995 118.995 112.515 ;
        RECT 119.205 112.465 119.435 113.285 ;
        RECT 119.605 112.485 119.935 113.115 ;
        RECT 119.185 112.045 119.515 112.295 ;
        RECT 119.685 111.885 119.935 112.485 ;
        RECT 120.105 112.465 120.315 113.285 ;
        RECT 120.635 112.735 120.805 113.115 ;
        RECT 120.985 112.905 121.315 113.285 ;
        RECT 120.635 112.565 121.300 112.735 ;
        RECT 121.495 112.610 121.755 113.115 ;
        RECT 120.565 112.015 120.895 112.385 ;
        RECT 121.130 112.310 121.300 112.565 ;
        RECT 115.485 110.735 118.995 111.825 ;
        RECT 119.205 110.735 119.435 111.875 ;
        RECT 119.605 110.905 119.935 111.885 ;
        RECT 121.130 111.980 121.415 112.310 ;
        RECT 120.105 110.735 120.315 111.875 ;
        RECT 121.130 111.835 121.300 111.980 ;
        RECT 120.635 111.665 121.300 111.835 ;
        RECT 121.585 111.810 121.755 112.610 ;
        RECT 120.635 110.905 120.805 111.665 ;
        RECT 120.985 110.735 121.315 111.495 ;
        RECT 121.485 110.905 121.755 111.810 ;
        RECT 121.925 112.610 122.185 113.115 ;
        RECT 122.365 112.905 122.695 113.285 ;
        RECT 122.875 112.735 123.045 113.115 ;
        RECT 121.925 111.810 122.095 112.610 ;
        RECT 122.380 112.565 123.045 112.735 ;
        RECT 122.380 112.310 122.550 112.565 ;
        RECT 123.765 112.515 126.355 113.285 ;
        RECT 126.525 112.535 127.735 113.285 ;
        RECT 122.265 111.980 122.550 112.310 ;
        RECT 122.785 112.015 123.115 112.385 ;
        RECT 122.380 111.835 122.550 111.980 ;
        RECT 121.925 110.905 122.195 111.810 ;
        RECT 122.380 111.665 123.045 111.835 ;
        RECT 122.365 110.735 122.695 111.495 ;
        RECT 122.875 110.905 123.045 111.665 ;
        RECT 123.765 111.825 124.975 112.345 ;
        RECT 125.145 111.995 126.355 112.515 ;
        RECT 126.525 111.825 127.045 112.365 ;
        RECT 127.215 111.995 127.735 112.535 ;
        RECT 123.765 110.735 126.355 111.825 ;
        RECT 126.525 110.735 127.735 111.825 ;
        RECT 14.660 110.565 127.820 110.735 ;
        RECT 14.745 109.475 15.955 110.565 ;
        RECT 14.745 108.765 15.265 109.305 ;
        RECT 15.435 108.935 15.955 109.475 ;
        RECT 16.125 109.475 17.335 110.565 ;
        RECT 17.510 110.130 22.855 110.565 ;
        RECT 16.125 108.935 16.645 109.475 ;
        RECT 16.815 108.765 17.335 109.305 ;
        RECT 19.100 108.880 19.450 110.130 ;
        RECT 23.115 109.635 23.285 110.395 ;
        RECT 23.465 109.805 23.795 110.565 ;
        RECT 23.115 109.465 23.780 109.635 ;
        RECT 23.965 109.490 24.235 110.395 ;
        RECT 14.745 108.015 15.955 108.765 ;
        RECT 16.125 108.015 17.335 108.765 ;
        RECT 20.930 108.560 21.270 109.390 ;
        RECT 23.610 109.320 23.780 109.465 ;
        RECT 23.045 108.915 23.375 109.285 ;
        RECT 23.610 108.990 23.895 109.320 ;
        RECT 23.610 108.735 23.780 108.990 ;
        RECT 23.115 108.565 23.780 108.735 ;
        RECT 24.065 108.690 24.235 109.490 ;
        RECT 24.405 109.400 24.695 110.565 ;
        RECT 25.175 109.725 25.345 110.565 ;
        RECT 25.555 109.555 25.805 110.395 ;
        RECT 26.015 109.725 26.185 110.565 ;
        RECT 26.355 109.555 26.645 110.395 ;
        RECT 24.920 109.385 26.645 109.555 ;
        RECT 26.855 109.505 27.025 110.565 ;
        RECT 27.320 110.185 27.650 110.565 ;
        RECT 27.830 110.015 28.000 110.305 ;
        RECT 28.170 110.105 28.420 110.565 ;
        RECT 27.200 109.845 28.000 110.015 ;
        RECT 28.590 110.055 29.460 110.395 ;
        RECT 24.920 108.835 25.330 109.385 ;
        RECT 27.200 109.225 27.370 109.845 ;
        RECT 28.590 109.675 28.760 110.055 ;
        RECT 29.695 109.935 29.865 110.395 ;
        RECT 30.035 110.105 30.405 110.565 ;
        RECT 30.700 109.965 30.870 110.305 ;
        RECT 31.040 110.135 31.370 110.565 ;
        RECT 31.605 109.965 31.775 110.305 ;
        RECT 27.540 109.505 28.760 109.675 ;
        RECT 28.930 109.595 29.390 109.885 ;
        RECT 29.695 109.765 30.255 109.935 ;
        RECT 30.700 109.795 31.775 109.965 ;
        RECT 31.945 110.065 32.625 110.395 ;
        RECT 32.840 110.065 33.090 110.395 ;
        RECT 33.260 110.105 33.510 110.565 ;
        RECT 30.085 109.625 30.255 109.765 ;
        RECT 28.930 109.585 29.895 109.595 ;
        RECT 28.590 109.415 28.760 109.505 ;
        RECT 29.220 109.425 29.895 109.585 ;
        RECT 27.200 109.215 27.545 109.225 ;
        RECT 25.515 109.005 27.545 109.215 ;
        RECT 17.510 108.015 22.855 108.560 ;
        RECT 23.115 108.185 23.285 108.565 ;
        RECT 23.465 108.015 23.795 108.395 ;
        RECT 23.975 108.185 24.235 108.690 ;
        RECT 24.405 108.015 24.695 108.740 ;
        RECT 24.920 108.665 26.685 108.835 ;
        RECT 25.175 108.015 25.345 108.485 ;
        RECT 25.515 108.185 25.845 108.665 ;
        RECT 26.015 108.015 26.185 108.485 ;
        RECT 26.355 108.185 26.685 108.665 ;
        RECT 26.855 108.015 27.025 108.825 ;
        RECT 27.220 108.750 27.545 109.005 ;
        RECT 27.225 108.395 27.545 108.750 ;
        RECT 27.715 108.965 28.255 109.335 ;
        RECT 28.590 109.245 28.995 109.415 ;
        RECT 27.715 108.565 27.955 108.965 ;
        RECT 28.435 108.795 28.655 109.075 ;
        RECT 28.125 108.625 28.655 108.795 ;
        RECT 28.125 108.395 28.295 108.625 ;
        RECT 28.825 108.465 28.995 109.245 ;
        RECT 29.165 108.635 29.515 109.255 ;
        RECT 29.685 108.635 29.895 109.425 ;
        RECT 30.085 109.455 31.585 109.625 ;
        RECT 30.085 108.765 30.255 109.455 ;
        RECT 31.945 109.285 32.115 110.065 ;
        RECT 32.920 109.935 33.090 110.065 ;
        RECT 30.425 109.115 32.115 109.285 ;
        RECT 32.285 109.505 32.750 109.895 ;
        RECT 32.920 109.765 33.315 109.935 ;
        RECT 30.425 108.935 30.595 109.115 ;
        RECT 27.225 108.225 28.295 108.395 ;
        RECT 28.465 108.015 28.655 108.455 ;
        RECT 28.825 108.185 29.775 108.465 ;
        RECT 30.085 108.375 30.345 108.765 ;
        RECT 30.765 108.695 31.555 108.945 ;
        RECT 29.995 108.205 30.345 108.375 ;
        RECT 30.555 108.015 30.885 108.475 ;
        RECT 31.760 108.405 31.930 109.115 ;
        RECT 32.285 108.915 32.455 109.505 ;
        RECT 32.100 108.695 32.455 108.915 ;
        RECT 32.625 108.695 32.975 109.315 ;
        RECT 33.145 108.405 33.315 109.765 ;
        RECT 33.680 109.595 34.005 110.380 ;
        RECT 33.485 108.545 33.945 109.595 ;
        RECT 31.760 108.235 32.615 108.405 ;
        RECT 32.820 108.235 33.315 108.405 ;
        RECT 33.485 108.015 33.815 108.375 ;
        RECT 34.175 108.275 34.345 110.395 ;
        RECT 34.515 110.065 34.845 110.565 ;
        RECT 35.015 109.895 35.270 110.395 ;
        RECT 34.520 109.725 35.270 109.895 ;
        RECT 36.675 109.725 36.845 110.565 ;
        RECT 34.520 108.735 34.750 109.725 ;
        RECT 37.055 109.555 37.305 110.395 ;
        RECT 37.515 109.725 37.685 110.565 ;
        RECT 37.855 109.555 38.145 110.395 ;
        RECT 34.920 108.905 35.270 109.555 ;
        RECT 36.420 109.385 38.145 109.555 ;
        RECT 38.355 109.505 38.525 110.565 ;
        RECT 38.820 110.185 39.150 110.565 ;
        RECT 39.330 110.015 39.500 110.305 ;
        RECT 39.670 110.105 39.920 110.565 ;
        RECT 38.700 109.845 39.500 110.015 ;
        RECT 40.090 110.055 40.960 110.395 ;
        RECT 36.420 108.835 36.830 109.385 ;
        RECT 38.700 109.225 38.870 109.845 ;
        RECT 40.090 109.675 40.260 110.055 ;
        RECT 41.195 109.935 41.365 110.395 ;
        RECT 41.535 110.105 41.905 110.565 ;
        RECT 42.200 109.965 42.370 110.305 ;
        RECT 42.540 110.135 42.870 110.565 ;
        RECT 43.105 109.965 43.275 110.305 ;
        RECT 39.040 109.505 40.260 109.675 ;
        RECT 40.430 109.595 40.890 109.885 ;
        RECT 41.195 109.765 41.755 109.935 ;
        RECT 42.200 109.795 43.275 109.965 ;
        RECT 43.445 110.065 44.125 110.395 ;
        RECT 44.340 110.065 44.590 110.395 ;
        RECT 44.760 110.105 45.010 110.565 ;
        RECT 41.585 109.625 41.755 109.765 ;
        RECT 40.430 109.585 41.395 109.595 ;
        RECT 40.090 109.415 40.260 109.505 ;
        RECT 40.720 109.425 41.395 109.585 ;
        RECT 38.700 109.215 39.045 109.225 ;
        RECT 37.015 109.005 39.045 109.215 ;
        RECT 34.520 108.565 35.270 108.735 ;
        RECT 36.420 108.665 38.185 108.835 ;
        RECT 34.515 108.015 34.845 108.395 ;
        RECT 35.015 108.275 35.270 108.565 ;
        RECT 36.675 108.015 36.845 108.485 ;
        RECT 37.015 108.185 37.345 108.665 ;
        RECT 37.515 108.015 37.685 108.485 ;
        RECT 37.855 108.185 38.185 108.665 ;
        RECT 38.355 108.015 38.525 108.825 ;
        RECT 38.720 108.750 39.045 109.005 ;
        RECT 38.725 108.395 39.045 108.750 ;
        RECT 39.215 108.965 39.755 109.335 ;
        RECT 40.090 109.245 40.495 109.415 ;
        RECT 39.215 108.565 39.455 108.965 ;
        RECT 39.935 108.795 40.155 109.075 ;
        RECT 39.625 108.625 40.155 108.795 ;
        RECT 39.625 108.395 39.795 108.625 ;
        RECT 40.325 108.465 40.495 109.245 ;
        RECT 40.665 108.635 41.015 109.255 ;
        RECT 41.185 108.635 41.395 109.425 ;
        RECT 41.585 109.455 43.085 109.625 ;
        RECT 41.585 108.765 41.755 109.455 ;
        RECT 43.445 109.285 43.615 110.065 ;
        RECT 44.420 109.935 44.590 110.065 ;
        RECT 41.925 109.115 43.615 109.285 ;
        RECT 43.785 109.505 44.250 109.895 ;
        RECT 44.420 109.765 44.815 109.935 ;
        RECT 41.925 108.935 42.095 109.115 ;
        RECT 38.725 108.225 39.795 108.395 ;
        RECT 39.965 108.015 40.155 108.455 ;
        RECT 40.325 108.185 41.275 108.465 ;
        RECT 41.585 108.375 41.845 108.765 ;
        RECT 42.265 108.695 43.055 108.945 ;
        RECT 41.495 108.205 41.845 108.375 ;
        RECT 42.055 108.015 42.385 108.475 ;
        RECT 43.260 108.405 43.430 109.115 ;
        RECT 43.785 108.915 43.955 109.505 ;
        RECT 43.600 108.695 43.955 108.915 ;
        RECT 44.125 108.695 44.475 109.315 ;
        RECT 44.645 108.405 44.815 109.765 ;
        RECT 45.180 109.595 45.505 110.380 ;
        RECT 44.985 108.545 45.445 109.595 ;
        RECT 43.260 108.235 44.115 108.405 ;
        RECT 44.320 108.235 44.815 108.405 ;
        RECT 44.985 108.015 45.315 108.375 ;
        RECT 45.675 108.275 45.845 110.395 ;
        RECT 46.015 110.065 46.345 110.565 ;
        RECT 46.515 109.895 46.770 110.395 ;
        RECT 46.020 109.725 46.770 109.895 ;
        RECT 46.020 108.735 46.250 109.725 ;
        RECT 46.420 108.905 46.770 109.555 ;
        RECT 46.945 109.490 47.215 110.395 ;
        RECT 47.385 109.805 47.715 110.565 ;
        RECT 47.895 109.635 48.065 110.395 ;
        RECT 46.020 108.565 46.770 108.735 ;
        RECT 46.015 108.015 46.345 108.395 ;
        RECT 46.515 108.275 46.770 108.565 ;
        RECT 46.945 108.690 47.115 109.490 ;
        RECT 47.400 109.465 48.065 109.635 ;
        RECT 48.325 109.475 49.995 110.565 ;
        RECT 47.400 109.320 47.570 109.465 ;
        RECT 47.285 108.990 47.570 109.320 ;
        RECT 47.400 108.735 47.570 108.990 ;
        RECT 47.805 108.915 48.135 109.285 ;
        RECT 48.325 108.955 49.075 109.475 ;
        RECT 50.165 109.400 50.455 110.565 ;
        RECT 51.545 109.475 55.055 110.565 ;
        RECT 55.315 109.635 55.485 110.395 ;
        RECT 55.665 109.805 55.995 110.565 ;
        RECT 49.245 108.785 49.995 109.305 ;
        RECT 51.545 108.955 53.235 109.475 ;
        RECT 55.315 109.465 55.980 109.635 ;
        RECT 56.165 109.490 56.435 110.395 ;
        RECT 55.810 109.320 55.980 109.465 ;
        RECT 53.405 108.785 55.055 109.305 ;
        RECT 55.245 108.915 55.575 109.285 ;
        RECT 55.810 108.990 56.095 109.320 ;
        RECT 46.945 108.185 47.205 108.690 ;
        RECT 47.400 108.565 48.065 108.735 ;
        RECT 47.385 108.015 47.715 108.395 ;
        RECT 47.895 108.185 48.065 108.565 ;
        RECT 48.325 108.015 49.995 108.785 ;
        RECT 50.165 108.015 50.455 108.740 ;
        RECT 51.545 108.015 55.055 108.785 ;
        RECT 55.810 108.735 55.980 108.990 ;
        RECT 55.315 108.565 55.980 108.735 ;
        RECT 56.265 108.690 56.435 109.490 ;
        RECT 56.605 109.475 60.115 110.565 ;
        RECT 60.295 109.585 60.625 110.395 ;
        RECT 60.795 109.765 61.035 110.565 ;
        RECT 56.605 108.955 58.295 109.475 ;
        RECT 60.295 109.415 61.010 109.585 ;
        RECT 58.465 108.785 60.115 109.305 ;
        RECT 60.290 109.005 60.670 109.245 ;
        RECT 60.840 109.175 61.010 109.415 ;
        RECT 61.215 109.545 61.385 110.395 ;
        RECT 61.555 109.765 61.885 110.565 ;
        RECT 62.055 109.545 62.225 110.395 ;
        RECT 61.215 109.375 62.225 109.545 ;
        RECT 62.395 109.415 62.725 110.565 ;
        RECT 63.595 109.635 63.765 110.395 ;
        RECT 63.945 109.805 64.275 110.565 ;
        RECT 63.595 109.465 64.260 109.635 ;
        RECT 64.445 109.490 64.715 110.395 ;
        RECT 60.840 109.005 61.340 109.175 ;
        RECT 60.840 108.835 61.010 109.005 ;
        RECT 61.730 108.865 62.225 109.375 ;
        RECT 64.090 109.320 64.260 109.465 ;
        RECT 63.525 108.915 63.855 109.285 ;
        RECT 64.090 108.990 64.375 109.320 ;
        RECT 61.725 108.835 62.225 108.865 ;
        RECT 55.315 108.185 55.485 108.565 ;
        RECT 55.665 108.015 55.995 108.395 ;
        RECT 56.175 108.185 56.435 108.690 ;
        RECT 56.605 108.015 60.115 108.785 ;
        RECT 60.375 108.665 61.010 108.835 ;
        RECT 61.215 108.665 62.225 108.835 ;
        RECT 60.375 108.185 60.545 108.665 ;
        RECT 60.725 108.015 60.965 108.495 ;
        RECT 61.215 108.185 61.385 108.665 ;
        RECT 61.555 108.015 61.885 108.495 ;
        RECT 62.055 108.185 62.225 108.665 ;
        RECT 62.395 108.015 62.725 108.815 ;
        RECT 64.090 108.735 64.260 108.990 ;
        RECT 63.595 108.565 64.260 108.735 ;
        RECT 64.545 108.690 64.715 109.490 ;
        RECT 65.345 109.475 67.935 110.565 ;
        RECT 68.195 109.635 68.365 110.395 ;
        RECT 68.545 109.805 68.875 110.565 ;
        RECT 65.345 108.955 66.555 109.475 ;
        RECT 68.195 109.465 68.860 109.635 ;
        RECT 69.045 109.490 69.315 110.395 ;
        RECT 68.690 109.320 68.860 109.465 ;
        RECT 66.725 108.785 67.935 109.305 ;
        RECT 68.125 108.915 68.455 109.285 ;
        RECT 68.690 108.990 68.975 109.320 ;
        RECT 63.595 108.185 63.765 108.565 ;
        RECT 63.945 108.015 64.275 108.395 ;
        RECT 64.455 108.185 64.715 108.690 ;
        RECT 65.345 108.015 67.935 108.785 ;
        RECT 68.690 108.735 68.860 108.990 ;
        RECT 68.195 108.565 68.860 108.735 ;
        RECT 69.145 108.690 69.315 109.490 ;
        RECT 69.485 109.475 70.695 110.565 ;
        RECT 70.865 109.475 74.375 110.565 ;
        RECT 69.485 108.935 70.005 109.475 ;
        RECT 70.175 108.765 70.695 109.305 ;
        RECT 70.865 108.955 72.555 109.475 ;
        RECT 74.605 109.425 74.815 110.565 ;
        RECT 74.985 109.415 75.315 110.395 ;
        RECT 75.485 109.425 75.715 110.565 ;
        RECT 72.725 108.785 74.375 109.305 ;
        RECT 68.195 108.185 68.365 108.565 ;
        RECT 68.545 108.015 68.875 108.395 ;
        RECT 69.055 108.185 69.315 108.690 ;
        RECT 69.485 108.015 70.695 108.765 ;
        RECT 70.865 108.015 74.375 108.785 ;
        RECT 74.605 108.015 74.815 108.835 ;
        RECT 74.985 108.815 75.235 109.415 ;
        RECT 75.925 109.400 76.215 110.565 ;
        RECT 76.905 109.425 77.115 110.565 ;
        RECT 77.285 109.415 77.615 110.395 ;
        RECT 77.785 109.425 78.015 110.565 ;
        RECT 78.235 109.585 78.565 110.395 ;
        RECT 78.735 109.765 78.975 110.565 ;
        RECT 78.235 109.415 78.950 109.585 ;
        RECT 75.405 109.005 75.735 109.255 ;
        RECT 74.985 108.185 75.315 108.815 ;
        RECT 75.485 108.015 75.715 108.835 ;
        RECT 75.925 108.015 76.215 108.740 ;
        RECT 76.905 108.015 77.115 108.835 ;
        RECT 77.285 108.815 77.535 109.415 ;
        RECT 77.705 109.005 78.035 109.255 ;
        RECT 78.230 109.005 78.610 109.245 ;
        RECT 78.780 109.175 78.950 109.415 ;
        RECT 79.155 109.545 79.325 110.395 ;
        RECT 79.495 109.765 79.825 110.565 ;
        RECT 79.995 109.545 80.165 110.395 ;
        RECT 79.155 109.375 80.165 109.545 ;
        RECT 80.335 109.415 80.665 110.565 ;
        RECT 81.075 109.635 81.245 110.395 ;
        RECT 81.425 109.805 81.755 110.565 ;
        RECT 81.075 109.465 81.740 109.635 ;
        RECT 81.925 109.490 82.195 110.395 ;
        RECT 79.670 109.205 80.165 109.375 ;
        RECT 81.570 109.320 81.740 109.465 ;
        RECT 78.780 109.005 79.280 109.175 ;
        RECT 79.665 109.035 80.165 109.205 ;
        RECT 78.780 108.835 78.950 109.005 ;
        RECT 79.670 108.835 80.165 109.035 ;
        RECT 81.005 108.915 81.335 109.285 ;
        RECT 81.570 108.990 81.855 109.320 ;
        RECT 77.285 108.185 77.615 108.815 ;
        RECT 77.785 108.015 78.015 108.835 ;
        RECT 78.315 108.665 78.950 108.835 ;
        RECT 79.155 108.665 80.165 108.835 ;
        RECT 78.315 108.185 78.485 108.665 ;
        RECT 78.665 108.015 78.905 108.495 ;
        RECT 79.155 108.185 79.325 108.665 ;
        RECT 79.495 108.015 79.825 108.495 ;
        RECT 79.995 108.185 80.165 108.665 ;
        RECT 80.335 108.015 80.665 108.815 ;
        RECT 81.570 108.735 81.740 108.990 ;
        RECT 81.075 108.565 81.740 108.735 ;
        RECT 82.025 108.690 82.195 109.490 ;
        RECT 82.455 109.635 82.625 110.395 ;
        RECT 82.805 109.805 83.135 110.565 ;
        RECT 82.455 109.465 83.120 109.635 ;
        RECT 83.305 109.490 83.575 110.395 ;
        RECT 82.950 109.320 83.120 109.465 ;
        RECT 82.385 108.915 82.715 109.285 ;
        RECT 82.950 108.990 83.235 109.320 ;
        RECT 82.950 108.735 83.120 108.990 ;
        RECT 81.075 108.185 81.245 108.565 ;
        RECT 81.425 108.015 81.755 108.395 ;
        RECT 81.935 108.185 82.195 108.690 ;
        RECT 82.455 108.565 83.120 108.735 ;
        RECT 83.405 108.690 83.575 109.490 ;
        RECT 84.665 109.475 88.175 110.565 ;
        RECT 84.665 108.955 86.355 109.475 ;
        RECT 88.385 109.425 88.615 110.565 ;
        RECT 88.785 109.415 89.115 110.395 ;
        RECT 89.285 109.425 89.495 110.565 ;
        RECT 89.815 109.635 89.985 110.395 ;
        RECT 90.165 109.805 90.495 110.565 ;
        RECT 89.815 109.465 90.480 109.635 ;
        RECT 90.665 109.490 90.935 110.395 ;
        RECT 91.415 109.725 91.585 110.565 ;
        RECT 91.795 109.555 92.045 110.395 ;
        RECT 92.255 109.725 92.425 110.565 ;
        RECT 92.595 109.555 92.885 110.395 ;
        RECT 86.525 108.785 88.175 109.305 ;
        RECT 88.365 109.005 88.695 109.255 ;
        RECT 82.455 108.185 82.625 108.565 ;
        RECT 82.805 108.015 83.135 108.395 ;
        RECT 83.315 108.185 83.575 108.690 ;
        RECT 84.665 108.015 88.175 108.785 ;
        RECT 88.385 108.015 88.615 108.835 ;
        RECT 88.865 108.815 89.115 109.415 ;
        RECT 90.310 109.320 90.480 109.465 ;
        RECT 89.745 108.915 90.075 109.285 ;
        RECT 90.310 108.990 90.595 109.320 ;
        RECT 88.785 108.185 89.115 108.815 ;
        RECT 89.285 108.015 89.495 108.835 ;
        RECT 90.310 108.735 90.480 108.990 ;
        RECT 89.815 108.565 90.480 108.735 ;
        RECT 90.765 108.690 90.935 109.490 ;
        RECT 89.815 108.185 89.985 108.565 ;
        RECT 90.165 108.015 90.495 108.395 ;
        RECT 90.675 108.185 90.935 108.690 ;
        RECT 91.160 109.385 92.885 109.555 ;
        RECT 93.095 109.505 93.265 110.565 ;
        RECT 93.560 110.185 93.890 110.565 ;
        RECT 94.070 110.015 94.240 110.305 ;
        RECT 94.410 110.105 94.660 110.565 ;
        RECT 93.440 109.845 94.240 110.015 ;
        RECT 94.830 110.055 95.700 110.395 ;
        RECT 91.160 108.835 91.570 109.385 ;
        RECT 93.440 109.225 93.610 109.845 ;
        RECT 94.830 109.675 95.000 110.055 ;
        RECT 95.935 109.935 96.105 110.395 ;
        RECT 96.275 110.105 96.645 110.565 ;
        RECT 96.940 109.965 97.110 110.305 ;
        RECT 97.280 110.135 97.610 110.565 ;
        RECT 97.845 109.965 98.015 110.305 ;
        RECT 93.780 109.505 95.000 109.675 ;
        RECT 95.170 109.595 95.630 109.885 ;
        RECT 95.935 109.765 96.495 109.935 ;
        RECT 96.940 109.795 98.015 109.965 ;
        RECT 98.185 110.065 98.865 110.395 ;
        RECT 99.080 110.065 99.330 110.395 ;
        RECT 99.500 110.105 99.750 110.565 ;
        RECT 96.325 109.625 96.495 109.765 ;
        RECT 95.170 109.585 96.135 109.595 ;
        RECT 94.830 109.415 95.000 109.505 ;
        RECT 95.460 109.425 96.135 109.585 ;
        RECT 93.440 109.215 93.785 109.225 ;
        RECT 91.755 109.005 93.785 109.215 ;
        RECT 91.160 108.665 92.925 108.835 ;
        RECT 91.415 108.015 91.585 108.485 ;
        RECT 91.755 108.185 92.085 108.665 ;
        RECT 92.255 108.015 92.425 108.485 ;
        RECT 92.595 108.185 92.925 108.665 ;
        RECT 93.095 108.015 93.265 108.825 ;
        RECT 93.460 108.750 93.785 109.005 ;
        RECT 93.465 108.395 93.785 108.750 ;
        RECT 93.955 108.965 94.495 109.335 ;
        RECT 94.830 109.245 95.235 109.415 ;
        RECT 93.955 108.565 94.195 108.965 ;
        RECT 94.675 108.795 94.895 109.075 ;
        RECT 94.365 108.625 94.895 108.795 ;
        RECT 94.365 108.395 94.535 108.625 ;
        RECT 95.065 108.465 95.235 109.245 ;
        RECT 95.405 108.635 95.755 109.255 ;
        RECT 95.925 108.635 96.135 109.425 ;
        RECT 96.325 109.455 97.825 109.625 ;
        RECT 96.325 108.765 96.495 109.455 ;
        RECT 98.185 109.285 98.355 110.065 ;
        RECT 99.160 109.935 99.330 110.065 ;
        RECT 96.665 109.115 98.355 109.285 ;
        RECT 98.525 109.505 98.990 109.895 ;
        RECT 99.160 109.765 99.555 109.935 ;
        RECT 96.665 108.935 96.835 109.115 ;
        RECT 93.465 108.225 94.535 108.395 ;
        RECT 94.705 108.015 94.895 108.455 ;
        RECT 95.065 108.185 96.015 108.465 ;
        RECT 96.325 108.375 96.585 108.765 ;
        RECT 97.005 108.695 97.795 108.945 ;
        RECT 96.235 108.205 96.585 108.375 ;
        RECT 96.795 108.015 97.125 108.475 ;
        RECT 98.000 108.405 98.170 109.115 ;
        RECT 98.525 108.915 98.695 109.505 ;
        RECT 98.340 108.695 98.695 108.915 ;
        RECT 98.865 108.695 99.215 109.315 ;
        RECT 99.385 108.405 99.555 109.765 ;
        RECT 99.920 109.595 100.245 110.380 ;
        RECT 99.725 108.545 100.185 109.595 ;
        RECT 98.000 108.235 98.855 108.405 ;
        RECT 99.060 108.235 99.555 108.405 ;
        RECT 99.725 108.015 100.055 108.375 ;
        RECT 100.415 108.275 100.585 110.395 ;
        RECT 100.755 110.065 101.085 110.565 ;
        RECT 101.255 109.895 101.510 110.395 ;
        RECT 100.760 109.725 101.510 109.895 ;
        RECT 100.760 108.735 100.990 109.725 ;
        RECT 101.160 108.905 101.510 109.555 ;
        RECT 101.685 109.400 101.975 110.565 ;
        RECT 102.145 109.490 102.415 110.395 ;
        RECT 102.585 109.805 102.915 110.565 ;
        RECT 103.095 109.635 103.265 110.395 ;
        RECT 100.760 108.565 101.510 108.735 ;
        RECT 100.755 108.015 101.085 108.395 ;
        RECT 101.255 108.275 101.510 108.565 ;
        RECT 101.685 108.015 101.975 108.740 ;
        RECT 102.145 108.690 102.315 109.490 ;
        RECT 102.600 109.465 103.265 109.635 ;
        RECT 102.600 109.320 102.770 109.465 ;
        RECT 104.505 109.425 104.715 110.565 ;
        RECT 102.485 108.990 102.770 109.320 ;
        RECT 104.885 109.415 105.215 110.395 ;
        RECT 105.385 109.425 105.615 110.565 ;
        RECT 106.835 109.635 107.005 110.395 ;
        RECT 107.185 109.805 107.515 110.565 ;
        RECT 106.835 109.465 107.500 109.635 ;
        RECT 107.685 109.490 107.955 110.395 ;
        RECT 102.600 108.735 102.770 108.990 ;
        RECT 103.005 108.915 103.335 109.285 ;
        RECT 102.145 108.185 102.405 108.690 ;
        RECT 102.600 108.565 103.265 108.735 ;
        RECT 102.585 108.015 102.915 108.395 ;
        RECT 103.095 108.185 103.265 108.565 ;
        RECT 104.505 108.015 104.715 108.835 ;
        RECT 104.885 108.815 105.135 109.415 ;
        RECT 107.330 109.320 107.500 109.465 ;
        RECT 105.305 109.005 105.635 109.255 ;
        RECT 106.765 108.915 107.095 109.285 ;
        RECT 107.330 108.990 107.615 109.320 ;
        RECT 104.885 108.185 105.215 108.815 ;
        RECT 105.385 108.015 105.615 108.835 ;
        RECT 107.330 108.735 107.500 108.990 ;
        RECT 106.835 108.565 107.500 108.735 ;
        RECT 107.785 108.690 107.955 109.490 ;
        RECT 108.125 109.475 109.335 110.565 ;
        RECT 109.505 109.490 109.775 110.395 ;
        RECT 109.945 109.805 110.275 110.565 ;
        RECT 110.455 109.635 110.625 110.395 ;
        RECT 108.125 108.935 108.645 109.475 ;
        RECT 108.815 108.765 109.335 109.305 ;
        RECT 106.835 108.185 107.005 108.565 ;
        RECT 107.185 108.015 107.515 108.395 ;
        RECT 107.695 108.185 107.955 108.690 ;
        RECT 108.125 108.015 109.335 108.765 ;
        RECT 109.505 108.690 109.675 109.490 ;
        RECT 109.960 109.465 110.625 109.635 ;
        RECT 110.885 109.475 114.395 110.565 ;
        RECT 114.655 109.635 114.825 110.395 ;
        RECT 115.005 109.805 115.335 110.565 ;
        RECT 109.960 109.320 110.130 109.465 ;
        RECT 109.845 108.990 110.130 109.320 ;
        RECT 109.960 108.735 110.130 108.990 ;
        RECT 110.365 108.915 110.695 109.285 ;
        RECT 110.885 108.955 112.575 109.475 ;
        RECT 114.655 109.465 115.320 109.635 ;
        RECT 115.505 109.490 115.775 110.395 ;
        RECT 115.950 109.895 116.205 110.395 ;
        RECT 116.375 110.065 116.705 110.565 ;
        RECT 115.950 109.725 116.700 109.895 ;
        RECT 115.150 109.320 115.320 109.465 ;
        RECT 112.745 108.785 114.395 109.305 ;
        RECT 114.585 108.915 114.915 109.285 ;
        RECT 115.150 108.990 115.435 109.320 ;
        RECT 109.505 108.185 109.765 108.690 ;
        RECT 109.960 108.565 110.625 108.735 ;
        RECT 109.945 108.015 110.275 108.395 ;
        RECT 110.455 108.185 110.625 108.565 ;
        RECT 110.885 108.015 114.395 108.785 ;
        RECT 115.150 108.735 115.320 108.990 ;
        RECT 114.655 108.565 115.320 108.735 ;
        RECT 115.605 108.690 115.775 109.490 ;
        RECT 115.950 108.905 116.300 109.555 ;
        RECT 116.470 108.735 116.700 109.725 ;
        RECT 114.655 108.185 114.825 108.565 ;
        RECT 115.005 108.015 115.335 108.395 ;
        RECT 115.515 108.185 115.775 108.690 ;
        RECT 115.950 108.565 116.700 108.735 ;
        RECT 115.950 108.275 116.205 108.565 ;
        RECT 116.375 108.015 116.705 108.395 ;
        RECT 116.875 108.275 117.045 110.395 ;
        RECT 117.215 109.595 117.540 110.380 ;
        RECT 117.710 110.105 117.960 110.565 ;
        RECT 118.130 110.065 118.380 110.395 ;
        RECT 118.595 110.065 119.275 110.395 ;
        RECT 118.130 109.935 118.300 110.065 ;
        RECT 117.905 109.765 118.300 109.935 ;
        RECT 117.275 108.545 117.735 109.595 ;
        RECT 117.905 108.405 118.075 109.765 ;
        RECT 118.470 109.505 118.935 109.895 ;
        RECT 118.245 108.695 118.595 109.315 ;
        RECT 118.765 108.915 118.935 109.505 ;
        RECT 119.105 109.285 119.275 110.065 ;
        RECT 119.445 109.965 119.615 110.305 ;
        RECT 119.850 110.135 120.180 110.565 ;
        RECT 120.350 109.965 120.520 110.305 ;
        RECT 120.815 110.105 121.185 110.565 ;
        RECT 119.445 109.795 120.520 109.965 ;
        RECT 121.355 109.935 121.525 110.395 ;
        RECT 121.760 110.055 122.630 110.395 ;
        RECT 122.800 110.105 123.050 110.565 ;
        RECT 120.965 109.765 121.525 109.935 ;
        RECT 120.965 109.625 121.135 109.765 ;
        RECT 119.635 109.455 121.135 109.625 ;
        RECT 121.830 109.595 122.290 109.885 ;
        RECT 119.105 109.115 120.795 109.285 ;
        RECT 118.765 108.695 119.120 108.915 ;
        RECT 119.290 108.405 119.460 109.115 ;
        RECT 119.665 108.695 120.455 108.945 ;
        RECT 120.625 108.935 120.795 109.115 ;
        RECT 120.965 108.765 121.135 109.455 ;
        RECT 117.405 108.015 117.735 108.375 ;
        RECT 117.905 108.235 118.400 108.405 ;
        RECT 118.605 108.235 119.460 108.405 ;
        RECT 120.335 108.015 120.665 108.475 ;
        RECT 120.875 108.375 121.135 108.765 ;
        RECT 121.325 109.585 122.290 109.595 ;
        RECT 122.460 109.675 122.630 110.055 ;
        RECT 123.220 110.015 123.390 110.305 ;
        RECT 123.570 110.185 123.900 110.565 ;
        RECT 123.220 109.845 124.020 110.015 ;
        RECT 121.325 109.425 122.000 109.585 ;
        RECT 122.460 109.505 123.680 109.675 ;
        RECT 121.325 108.635 121.535 109.425 ;
        RECT 122.460 109.415 122.630 109.505 ;
        RECT 121.705 108.635 122.055 109.255 ;
        RECT 122.225 109.245 122.630 109.415 ;
        RECT 122.225 108.465 122.395 109.245 ;
        RECT 122.565 108.795 122.785 109.075 ;
        RECT 122.965 108.965 123.505 109.335 ;
        RECT 123.850 109.225 124.020 109.845 ;
        RECT 124.195 109.505 124.365 110.565 ;
        RECT 124.575 109.555 124.865 110.395 ;
        RECT 125.035 109.725 125.205 110.565 ;
        RECT 125.415 109.555 125.665 110.395 ;
        RECT 125.875 109.725 126.045 110.565 ;
        RECT 124.575 109.385 126.300 109.555 ;
        RECT 122.565 108.625 123.095 108.795 ;
        RECT 120.875 108.205 121.225 108.375 ;
        RECT 121.445 108.185 122.395 108.465 ;
        RECT 122.565 108.015 122.755 108.455 ;
        RECT 122.925 108.395 123.095 108.625 ;
        RECT 123.265 108.565 123.505 108.965 ;
        RECT 123.675 109.215 124.020 109.225 ;
        RECT 123.675 109.005 125.705 109.215 ;
        RECT 123.675 108.750 124.000 109.005 ;
        RECT 125.890 108.835 126.300 109.385 ;
        RECT 126.525 109.475 127.735 110.565 ;
        RECT 126.525 108.935 127.045 109.475 ;
        RECT 123.675 108.395 123.995 108.750 ;
        RECT 122.925 108.225 123.995 108.395 ;
        RECT 124.195 108.015 124.365 108.825 ;
        RECT 124.535 108.665 126.300 108.835 ;
        RECT 127.215 108.765 127.735 109.305 ;
        RECT 124.535 108.185 124.865 108.665 ;
        RECT 125.035 108.015 125.205 108.485 ;
        RECT 125.375 108.185 125.705 108.665 ;
        RECT 125.875 108.015 126.045 108.485 ;
        RECT 126.525 108.015 127.735 108.765 ;
        RECT 14.660 107.845 127.820 108.015 ;
        RECT 14.745 107.095 15.955 107.845 ;
        RECT 14.745 106.555 15.265 107.095 ;
        RECT 16.585 107.075 20.095 107.845 ;
        RECT 15.435 106.385 15.955 106.925 ;
        RECT 14.745 105.295 15.955 106.385 ;
        RECT 16.585 106.385 18.275 106.905 ;
        RECT 18.445 106.555 20.095 107.075 ;
        RECT 20.325 107.025 20.535 107.845 ;
        RECT 20.705 107.045 21.035 107.675 ;
        RECT 20.705 106.445 20.955 107.045 ;
        RECT 21.205 107.025 21.435 107.845 ;
        RECT 22.625 107.025 22.835 107.845 ;
        RECT 23.005 107.045 23.335 107.675 ;
        RECT 21.125 106.605 21.455 106.855 ;
        RECT 23.005 106.445 23.255 107.045 ;
        RECT 23.505 107.025 23.735 107.845 ;
        RECT 24.255 107.375 24.425 107.845 ;
        RECT 24.595 107.195 24.925 107.675 ;
        RECT 25.095 107.375 25.265 107.845 ;
        RECT 25.435 107.195 25.765 107.675 ;
        RECT 24.000 107.025 25.765 107.195 ;
        RECT 25.935 107.035 26.105 107.845 ;
        RECT 26.305 107.465 27.375 107.635 ;
        RECT 26.305 107.110 26.625 107.465 ;
        RECT 23.425 106.605 23.755 106.855 ;
        RECT 24.000 106.475 24.410 107.025 ;
        RECT 26.300 106.855 26.625 107.110 ;
        RECT 24.595 106.645 26.625 106.855 ;
        RECT 26.280 106.635 26.625 106.645 ;
        RECT 26.795 106.895 27.035 107.295 ;
        RECT 27.205 107.235 27.375 107.465 ;
        RECT 27.545 107.405 27.735 107.845 ;
        RECT 27.905 107.395 28.855 107.675 ;
        RECT 29.075 107.485 29.425 107.655 ;
        RECT 27.205 107.065 27.735 107.235 ;
        RECT 16.585 105.295 20.095 106.385 ;
        RECT 20.325 105.295 20.535 106.435 ;
        RECT 20.705 105.465 21.035 106.445 ;
        RECT 21.205 105.295 21.435 106.435 ;
        RECT 22.625 105.295 22.835 106.435 ;
        RECT 23.005 105.465 23.335 106.445 ;
        RECT 23.505 105.295 23.735 106.435 ;
        RECT 24.000 106.305 25.725 106.475 ;
        RECT 24.255 105.295 24.425 106.135 ;
        RECT 24.635 105.465 24.885 106.305 ;
        RECT 25.095 105.295 25.265 106.135 ;
        RECT 25.435 105.465 25.725 106.305 ;
        RECT 25.935 105.295 26.105 106.355 ;
        RECT 26.280 106.015 26.450 106.635 ;
        RECT 26.795 106.525 27.335 106.895 ;
        RECT 27.515 106.785 27.735 107.065 ;
        RECT 27.905 106.615 28.075 107.395 ;
        RECT 27.670 106.445 28.075 106.615 ;
        RECT 28.245 106.605 28.595 107.225 ;
        RECT 27.670 106.355 27.840 106.445 ;
        RECT 28.765 106.435 28.975 107.225 ;
        RECT 26.620 106.185 27.840 106.355 ;
        RECT 28.300 106.275 28.975 106.435 ;
        RECT 26.280 105.845 27.080 106.015 ;
        RECT 26.400 105.295 26.730 105.675 ;
        RECT 26.910 105.555 27.080 105.845 ;
        RECT 27.670 105.805 27.840 106.185 ;
        RECT 28.010 106.265 28.975 106.275 ;
        RECT 29.165 107.095 29.425 107.485 ;
        RECT 29.635 107.385 29.965 107.845 ;
        RECT 30.840 107.455 31.695 107.625 ;
        RECT 31.900 107.455 32.395 107.625 ;
        RECT 32.565 107.485 32.895 107.845 ;
        RECT 29.165 106.405 29.335 107.095 ;
        RECT 29.505 106.745 29.675 106.925 ;
        RECT 29.845 106.915 30.635 107.165 ;
        RECT 30.840 106.745 31.010 107.455 ;
        RECT 31.180 106.945 31.535 107.165 ;
        RECT 29.505 106.575 31.195 106.745 ;
        RECT 28.010 105.975 28.470 106.265 ;
        RECT 29.165 106.235 30.665 106.405 ;
        RECT 29.165 106.095 29.335 106.235 ;
        RECT 28.775 105.925 29.335 106.095 ;
        RECT 27.250 105.295 27.500 105.755 ;
        RECT 27.670 105.465 28.540 105.805 ;
        RECT 28.775 105.465 28.945 105.925 ;
        RECT 29.780 105.895 30.855 106.065 ;
        RECT 29.115 105.295 29.485 105.755 ;
        RECT 29.780 105.555 29.950 105.895 ;
        RECT 30.120 105.295 30.450 105.725 ;
        RECT 30.685 105.555 30.855 105.895 ;
        RECT 31.025 105.795 31.195 106.575 ;
        RECT 31.365 106.355 31.535 106.945 ;
        RECT 31.705 106.545 32.055 107.165 ;
        RECT 31.365 105.965 31.830 106.355 ;
        RECT 32.225 106.095 32.395 107.455 ;
        RECT 32.565 106.265 33.025 107.315 ;
        RECT 32.000 105.925 32.395 106.095 ;
        RECT 32.000 105.795 32.170 105.925 ;
        RECT 31.025 105.465 31.705 105.795 ;
        RECT 31.920 105.465 32.170 105.795 ;
        RECT 32.340 105.295 32.590 105.755 ;
        RECT 32.760 105.480 33.085 106.265 ;
        RECT 33.255 105.465 33.425 107.585 ;
        RECT 33.595 107.465 33.925 107.845 ;
        RECT 34.095 107.295 34.350 107.585 ;
        RECT 33.600 107.125 34.350 107.295 ;
        RECT 33.600 106.135 33.830 107.125 ;
        RECT 34.565 107.025 34.795 107.845 ;
        RECT 34.965 107.045 35.295 107.675 ;
        RECT 34.000 106.305 34.350 106.955 ;
        RECT 34.545 106.605 34.875 106.855 ;
        RECT 35.045 106.445 35.295 107.045 ;
        RECT 35.465 107.025 35.675 107.845 ;
        RECT 35.945 107.025 36.175 107.845 ;
        RECT 36.345 107.045 36.675 107.675 ;
        RECT 35.925 106.605 36.255 106.855 ;
        RECT 36.425 106.445 36.675 107.045 ;
        RECT 36.845 107.025 37.055 107.845 ;
        RECT 37.285 107.120 37.575 107.845 ;
        RECT 38.515 107.375 38.685 107.845 ;
        RECT 38.855 107.195 39.185 107.675 ;
        RECT 39.355 107.375 39.525 107.845 ;
        RECT 39.695 107.195 40.025 107.675 ;
        RECT 38.260 107.025 40.025 107.195 ;
        RECT 40.195 107.035 40.365 107.845 ;
        RECT 40.565 107.465 41.635 107.635 ;
        RECT 40.565 107.110 40.885 107.465 ;
        RECT 38.260 106.475 38.670 107.025 ;
        RECT 40.560 106.855 40.885 107.110 ;
        RECT 38.855 106.645 40.885 106.855 ;
        RECT 40.540 106.635 40.885 106.645 ;
        RECT 41.055 106.895 41.295 107.295 ;
        RECT 41.465 107.235 41.635 107.465 ;
        RECT 41.805 107.405 41.995 107.845 ;
        RECT 42.165 107.395 43.115 107.675 ;
        RECT 43.335 107.485 43.685 107.655 ;
        RECT 41.465 107.065 41.995 107.235 ;
        RECT 33.600 105.965 34.350 106.135 ;
        RECT 33.595 105.295 33.925 105.795 ;
        RECT 34.095 105.465 34.350 105.965 ;
        RECT 34.565 105.295 34.795 106.435 ;
        RECT 34.965 105.465 35.295 106.445 ;
        RECT 35.465 105.295 35.675 106.435 ;
        RECT 35.945 105.295 36.175 106.435 ;
        RECT 36.345 105.465 36.675 106.445 ;
        RECT 36.845 105.295 37.055 106.435 ;
        RECT 37.285 105.295 37.575 106.460 ;
        RECT 38.260 106.305 39.985 106.475 ;
        RECT 38.515 105.295 38.685 106.135 ;
        RECT 38.895 105.465 39.145 106.305 ;
        RECT 39.355 105.295 39.525 106.135 ;
        RECT 39.695 105.465 39.985 106.305 ;
        RECT 40.195 105.295 40.365 106.355 ;
        RECT 40.540 106.015 40.710 106.635 ;
        RECT 41.055 106.525 41.595 106.895 ;
        RECT 41.775 106.785 41.995 107.065 ;
        RECT 42.165 106.615 42.335 107.395 ;
        RECT 41.930 106.445 42.335 106.615 ;
        RECT 42.505 106.605 42.855 107.225 ;
        RECT 41.930 106.355 42.100 106.445 ;
        RECT 43.025 106.435 43.235 107.225 ;
        RECT 40.880 106.185 42.100 106.355 ;
        RECT 42.560 106.275 43.235 106.435 ;
        RECT 40.540 105.845 41.340 106.015 ;
        RECT 40.660 105.295 40.990 105.675 ;
        RECT 41.170 105.555 41.340 105.845 ;
        RECT 41.930 105.805 42.100 106.185 ;
        RECT 42.270 106.265 43.235 106.275 ;
        RECT 43.425 107.095 43.685 107.485 ;
        RECT 43.895 107.385 44.225 107.845 ;
        RECT 45.100 107.455 45.955 107.625 ;
        RECT 46.160 107.455 46.655 107.625 ;
        RECT 46.825 107.485 47.155 107.845 ;
        RECT 43.425 106.405 43.595 107.095 ;
        RECT 43.765 106.745 43.935 106.925 ;
        RECT 44.105 106.915 44.895 107.165 ;
        RECT 45.100 106.745 45.270 107.455 ;
        RECT 45.440 106.945 45.795 107.165 ;
        RECT 43.765 106.575 45.455 106.745 ;
        RECT 42.270 105.975 42.730 106.265 ;
        RECT 43.425 106.235 44.925 106.405 ;
        RECT 43.425 106.095 43.595 106.235 ;
        RECT 43.035 105.925 43.595 106.095 ;
        RECT 41.510 105.295 41.760 105.755 ;
        RECT 41.930 105.465 42.800 105.805 ;
        RECT 43.035 105.465 43.205 105.925 ;
        RECT 44.040 105.895 45.115 106.065 ;
        RECT 43.375 105.295 43.745 105.755 ;
        RECT 44.040 105.555 44.210 105.895 ;
        RECT 44.380 105.295 44.710 105.725 ;
        RECT 44.945 105.555 45.115 105.895 ;
        RECT 45.285 105.795 45.455 106.575 ;
        RECT 45.625 106.355 45.795 106.945 ;
        RECT 45.965 106.545 46.315 107.165 ;
        RECT 45.625 105.965 46.090 106.355 ;
        RECT 46.485 106.095 46.655 107.455 ;
        RECT 46.825 106.265 47.285 107.315 ;
        RECT 46.260 105.925 46.655 106.095 ;
        RECT 46.260 105.795 46.430 105.925 ;
        RECT 45.285 105.465 45.965 105.795 ;
        RECT 46.180 105.465 46.430 105.795 ;
        RECT 46.600 105.295 46.850 105.755 ;
        RECT 47.020 105.480 47.345 106.265 ;
        RECT 47.515 105.465 47.685 107.585 ;
        RECT 47.855 107.465 48.185 107.845 ;
        RECT 48.355 107.295 48.610 107.585 ;
        RECT 47.860 107.125 48.610 107.295 ;
        RECT 47.860 106.135 48.090 107.125 ;
        RECT 48.845 107.025 49.055 107.845 ;
        RECT 49.225 107.045 49.555 107.675 ;
        RECT 48.260 106.305 48.610 106.955 ;
        RECT 49.225 106.445 49.475 107.045 ;
        RECT 49.725 107.025 49.955 107.845 ;
        RECT 50.165 107.170 50.425 107.675 ;
        RECT 50.605 107.465 50.935 107.845 ;
        RECT 51.115 107.295 51.285 107.675 ;
        RECT 51.855 107.375 52.025 107.845 ;
        RECT 49.645 106.605 49.975 106.855 ;
        RECT 47.860 105.965 48.610 106.135 ;
        RECT 47.855 105.295 48.185 105.795 ;
        RECT 48.355 105.465 48.610 105.965 ;
        RECT 48.845 105.295 49.055 106.435 ;
        RECT 49.225 105.465 49.555 106.445 ;
        RECT 49.725 105.295 49.955 106.435 ;
        RECT 50.165 106.370 50.335 107.170 ;
        RECT 50.620 107.125 51.285 107.295 ;
        RECT 52.195 107.195 52.525 107.675 ;
        RECT 52.695 107.375 52.865 107.845 ;
        RECT 53.035 107.195 53.365 107.675 ;
        RECT 50.620 106.870 50.790 107.125 ;
        RECT 51.600 107.025 53.365 107.195 ;
        RECT 53.535 107.035 53.705 107.845 ;
        RECT 53.905 107.465 54.975 107.635 ;
        RECT 53.905 107.110 54.225 107.465 ;
        RECT 50.505 106.540 50.790 106.870 ;
        RECT 51.025 106.575 51.355 106.945 ;
        RECT 50.620 106.395 50.790 106.540 ;
        RECT 51.600 106.475 52.010 107.025 ;
        RECT 53.900 106.855 54.225 107.110 ;
        RECT 52.195 106.645 54.225 106.855 ;
        RECT 53.880 106.635 54.225 106.645 ;
        RECT 54.395 106.895 54.635 107.295 ;
        RECT 54.805 107.235 54.975 107.465 ;
        RECT 55.145 107.405 55.335 107.845 ;
        RECT 55.505 107.395 56.455 107.675 ;
        RECT 56.675 107.485 57.025 107.655 ;
        RECT 54.805 107.065 55.335 107.235 ;
        RECT 50.165 105.465 50.435 106.370 ;
        RECT 50.620 106.225 51.285 106.395 ;
        RECT 51.600 106.305 53.325 106.475 ;
        RECT 50.605 105.295 50.935 106.055 ;
        RECT 51.115 105.465 51.285 106.225 ;
        RECT 51.855 105.295 52.025 106.135 ;
        RECT 52.235 105.465 52.485 106.305 ;
        RECT 52.695 105.295 52.865 106.135 ;
        RECT 53.035 105.465 53.325 106.305 ;
        RECT 53.535 105.295 53.705 106.355 ;
        RECT 53.880 106.015 54.050 106.635 ;
        RECT 54.395 106.525 54.935 106.895 ;
        RECT 55.115 106.785 55.335 107.065 ;
        RECT 55.505 106.615 55.675 107.395 ;
        RECT 55.270 106.445 55.675 106.615 ;
        RECT 55.845 106.605 56.195 107.225 ;
        RECT 55.270 106.355 55.440 106.445 ;
        RECT 56.365 106.435 56.575 107.225 ;
        RECT 54.220 106.185 55.440 106.355 ;
        RECT 55.900 106.275 56.575 106.435 ;
        RECT 53.880 105.845 54.680 106.015 ;
        RECT 54.000 105.295 54.330 105.675 ;
        RECT 54.510 105.555 54.680 105.845 ;
        RECT 55.270 105.805 55.440 106.185 ;
        RECT 55.610 106.265 56.575 106.275 ;
        RECT 56.765 107.095 57.025 107.485 ;
        RECT 57.235 107.385 57.565 107.845 ;
        RECT 58.440 107.455 59.295 107.625 ;
        RECT 59.500 107.455 59.995 107.625 ;
        RECT 60.165 107.485 60.495 107.845 ;
        RECT 56.765 106.405 56.935 107.095 ;
        RECT 57.105 106.745 57.275 106.925 ;
        RECT 57.445 106.915 58.235 107.165 ;
        RECT 58.440 106.745 58.610 107.455 ;
        RECT 58.780 106.945 59.135 107.165 ;
        RECT 57.105 106.575 58.795 106.745 ;
        RECT 55.610 105.975 56.070 106.265 ;
        RECT 56.765 106.235 58.265 106.405 ;
        RECT 56.765 106.095 56.935 106.235 ;
        RECT 56.375 105.925 56.935 106.095 ;
        RECT 54.850 105.295 55.100 105.755 ;
        RECT 55.270 105.465 56.140 105.805 ;
        RECT 56.375 105.465 56.545 105.925 ;
        RECT 57.380 105.895 58.455 106.065 ;
        RECT 56.715 105.295 57.085 105.755 ;
        RECT 57.380 105.555 57.550 105.895 ;
        RECT 57.720 105.295 58.050 105.725 ;
        RECT 58.285 105.555 58.455 105.895 ;
        RECT 58.625 105.795 58.795 106.575 ;
        RECT 58.965 106.355 59.135 106.945 ;
        RECT 59.305 106.545 59.655 107.165 ;
        RECT 58.965 105.965 59.430 106.355 ;
        RECT 59.825 106.095 59.995 107.455 ;
        RECT 60.165 106.265 60.625 107.315 ;
        RECT 59.600 105.925 59.995 106.095 ;
        RECT 59.600 105.795 59.770 105.925 ;
        RECT 58.625 105.465 59.305 105.795 ;
        RECT 59.520 105.465 59.770 105.795 ;
        RECT 59.940 105.295 60.190 105.755 ;
        RECT 60.360 105.480 60.685 106.265 ;
        RECT 60.855 105.465 61.025 107.585 ;
        RECT 61.195 107.465 61.525 107.845 ;
        RECT 61.695 107.295 61.950 107.585 ;
        RECT 61.200 107.125 61.950 107.295 ;
        RECT 61.200 106.135 61.430 107.125 ;
        RECT 63.045 107.120 63.335 107.845 ;
        RECT 63.815 107.375 63.985 107.845 ;
        RECT 64.155 107.195 64.485 107.675 ;
        RECT 64.655 107.375 64.825 107.845 ;
        RECT 64.995 107.195 65.325 107.675 ;
        RECT 63.560 107.025 65.325 107.195 ;
        RECT 65.495 107.035 65.665 107.845 ;
        RECT 65.865 107.465 66.935 107.635 ;
        RECT 65.865 107.110 66.185 107.465 ;
        RECT 61.600 106.305 61.950 106.955 ;
        RECT 63.560 106.475 63.970 107.025 ;
        RECT 65.860 106.855 66.185 107.110 ;
        RECT 64.155 106.645 66.185 106.855 ;
        RECT 65.840 106.635 66.185 106.645 ;
        RECT 66.355 106.895 66.595 107.295 ;
        RECT 66.765 107.235 66.935 107.465 ;
        RECT 67.105 107.405 67.295 107.845 ;
        RECT 67.465 107.395 68.415 107.675 ;
        RECT 68.635 107.485 68.985 107.655 ;
        RECT 66.765 107.065 67.295 107.235 ;
        RECT 61.200 105.965 61.950 106.135 ;
        RECT 61.195 105.295 61.525 105.795 ;
        RECT 61.695 105.465 61.950 105.965 ;
        RECT 63.045 105.295 63.335 106.460 ;
        RECT 63.560 106.305 65.285 106.475 ;
        RECT 63.815 105.295 63.985 106.135 ;
        RECT 64.195 105.465 64.445 106.305 ;
        RECT 64.655 105.295 64.825 106.135 ;
        RECT 64.995 105.465 65.285 106.305 ;
        RECT 65.495 105.295 65.665 106.355 ;
        RECT 65.840 106.015 66.010 106.635 ;
        RECT 66.355 106.525 66.895 106.895 ;
        RECT 67.075 106.785 67.295 107.065 ;
        RECT 67.465 106.615 67.635 107.395 ;
        RECT 67.230 106.445 67.635 106.615 ;
        RECT 67.805 106.605 68.155 107.225 ;
        RECT 67.230 106.355 67.400 106.445 ;
        RECT 68.325 106.435 68.535 107.225 ;
        RECT 66.180 106.185 67.400 106.355 ;
        RECT 67.860 106.275 68.535 106.435 ;
        RECT 65.840 105.845 66.640 106.015 ;
        RECT 65.960 105.295 66.290 105.675 ;
        RECT 66.470 105.555 66.640 105.845 ;
        RECT 67.230 105.805 67.400 106.185 ;
        RECT 67.570 106.265 68.535 106.275 ;
        RECT 68.725 107.095 68.985 107.485 ;
        RECT 69.195 107.385 69.525 107.845 ;
        RECT 70.400 107.455 71.255 107.625 ;
        RECT 71.460 107.455 71.955 107.625 ;
        RECT 72.125 107.485 72.455 107.845 ;
        RECT 68.725 106.405 68.895 107.095 ;
        RECT 69.065 106.745 69.235 106.925 ;
        RECT 69.405 106.915 70.195 107.165 ;
        RECT 70.400 106.745 70.570 107.455 ;
        RECT 70.740 106.945 71.095 107.165 ;
        RECT 69.065 106.575 70.755 106.745 ;
        RECT 67.570 105.975 68.030 106.265 ;
        RECT 68.725 106.235 70.225 106.405 ;
        RECT 68.725 106.095 68.895 106.235 ;
        RECT 68.335 105.925 68.895 106.095 ;
        RECT 66.810 105.295 67.060 105.755 ;
        RECT 67.230 105.465 68.100 105.805 ;
        RECT 68.335 105.465 68.505 105.925 ;
        RECT 69.340 105.895 70.415 106.065 ;
        RECT 68.675 105.295 69.045 105.755 ;
        RECT 69.340 105.555 69.510 105.895 ;
        RECT 69.680 105.295 70.010 105.725 ;
        RECT 70.245 105.555 70.415 105.895 ;
        RECT 70.585 105.795 70.755 106.575 ;
        RECT 70.925 106.355 71.095 106.945 ;
        RECT 71.265 106.545 71.615 107.165 ;
        RECT 70.925 105.965 71.390 106.355 ;
        RECT 71.785 106.095 71.955 107.455 ;
        RECT 72.125 106.265 72.585 107.315 ;
        RECT 71.560 105.925 71.955 106.095 ;
        RECT 71.560 105.795 71.730 105.925 ;
        RECT 70.585 105.465 71.265 105.795 ;
        RECT 71.480 105.465 71.730 105.795 ;
        RECT 71.900 105.295 72.150 105.755 ;
        RECT 72.320 105.480 72.645 106.265 ;
        RECT 72.815 105.465 72.985 107.585 ;
        RECT 73.155 107.465 73.485 107.845 ;
        RECT 73.655 107.295 73.910 107.585 ;
        RECT 75.315 107.375 75.485 107.845 ;
        RECT 73.160 107.125 73.910 107.295 ;
        RECT 75.655 107.195 75.985 107.675 ;
        RECT 76.155 107.375 76.325 107.845 ;
        RECT 76.495 107.195 76.825 107.675 ;
        RECT 73.160 106.135 73.390 107.125 ;
        RECT 75.060 107.025 76.825 107.195 ;
        RECT 76.995 107.035 77.165 107.845 ;
        RECT 77.365 107.465 78.435 107.635 ;
        RECT 77.365 107.110 77.685 107.465 ;
        RECT 73.560 106.305 73.910 106.955 ;
        RECT 75.060 106.475 75.470 107.025 ;
        RECT 77.360 106.855 77.685 107.110 ;
        RECT 75.655 106.645 77.685 106.855 ;
        RECT 77.340 106.635 77.685 106.645 ;
        RECT 77.855 106.895 78.095 107.295 ;
        RECT 78.265 107.235 78.435 107.465 ;
        RECT 78.605 107.405 78.795 107.845 ;
        RECT 78.965 107.395 79.915 107.675 ;
        RECT 80.135 107.485 80.485 107.655 ;
        RECT 78.265 107.065 78.795 107.235 ;
        RECT 75.060 106.305 76.785 106.475 ;
        RECT 73.160 105.965 73.910 106.135 ;
        RECT 73.155 105.295 73.485 105.795 ;
        RECT 73.655 105.465 73.910 105.965 ;
        RECT 75.315 105.295 75.485 106.135 ;
        RECT 75.695 105.465 75.945 106.305 ;
        RECT 76.155 105.295 76.325 106.135 ;
        RECT 76.495 105.465 76.785 106.305 ;
        RECT 76.995 105.295 77.165 106.355 ;
        RECT 77.340 106.015 77.510 106.635 ;
        RECT 77.855 106.525 78.395 106.895 ;
        RECT 78.575 106.785 78.795 107.065 ;
        RECT 78.965 106.615 79.135 107.395 ;
        RECT 78.730 106.445 79.135 106.615 ;
        RECT 79.305 106.605 79.655 107.225 ;
        RECT 78.730 106.355 78.900 106.445 ;
        RECT 79.825 106.435 80.035 107.225 ;
        RECT 77.680 106.185 78.900 106.355 ;
        RECT 79.360 106.275 80.035 106.435 ;
        RECT 77.340 105.845 78.140 106.015 ;
        RECT 77.460 105.295 77.790 105.675 ;
        RECT 77.970 105.555 78.140 105.845 ;
        RECT 78.730 105.805 78.900 106.185 ;
        RECT 79.070 106.265 80.035 106.275 ;
        RECT 80.225 107.095 80.485 107.485 ;
        RECT 80.695 107.385 81.025 107.845 ;
        RECT 81.900 107.455 82.755 107.625 ;
        RECT 82.960 107.455 83.455 107.625 ;
        RECT 83.625 107.485 83.955 107.845 ;
        RECT 80.225 106.405 80.395 107.095 ;
        RECT 80.565 106.745 80.735 106.925 ;
        RECT 80.905 106.915 81.695 107.165 ;
        RECT 81.900 106.745 82.070 107.455 ;
        RECT 82.240 106.945 82.595 107.165 ;
        RECT 80.565 106.575 82.255 106.745 ;
        RECT 79.070 105.975 79.530 106.265 ;
        RECT 80.225 106.235 81.725 106.405 ;
        RECT 80.225 106.095 80.395 106.235 ;
        RECT 79.835 105.925 80.395 106.095 ;
        RECT 78.310 105.295 78.560 105.755 ;
        RECT 78.730 105.465 79.600 105.805 ;
        RECT 79.835 105.465 80.005 105.925 ;
        RECT 80.840 105.895 81.915 106.065 ;
        RECT 80.175 105.295 80.545 105.755 ;
        RECT 80.840 105.555 81.010 105.895 ;
        RECT 81.180 105.295 81.510 105.725 ;
        RECT 81.745 105.555 81.915 105.895 ;
        RECT 82.085 105.795 82.255 106.575 ;
        RECT 82.425 106.355 82.595 106.945 ;
        RECT 82.765 106.545 83.115 107.165 ;
        RECT 82.425 105.965 82.890 106.355 ;
        RECT 83.285 106.095 83.455 107.455 ;
        RECT 83.625 106.265 84.085 107.315 ;
        RECT 83.060 105.925 83.455 106.095 ;
        RECT 83.060 105.795 83.230 105.925 ;
        RECT 82.085 105.465 82.765 105.795 ;
        RECT 82.980 105.465 83.230 105.795 ;
        RECT 83.400 105.295 83.650 105.755 ;
        RECT 83.820 105.480 84.145 106.265 ;
        RECT 84.315 105.465 84.485 107.585 ;
        RECT 84.655 107.465 84.985 107.845 ;
        RECT 85.155 107.295 85.410 107.585 ;
        RECT 84.660 107.125 85.410 107.295 ;
        RECT 84.660 106.135 84.890 107.125 ;
        RECT 85.625 107.025 85.855 107.845 ;
        RECT 86.025 107.045 86.355 107.675 ;
        RECT 85.060 106.305 85.410 106.955 ;
        RECT 85.605 106.605 85.935 106.855 ;
        RECT 86.105 106.445 86.355 107.045 ;
        RECT 86.525 107.025 86.735 107.845 ;
        RECT 87.055 107.295 87.225 107.675 ;
        RECT 87.405 107.465 87.735 107.845 ;
        RECT 87.055 107.125 87.720 107.295 ;
        RECT 87.915 107.170 88.175 107.675 ;
        RECT 86.985 106.575 87.315 106.945 ;
        RECT 87.550 106.870 87.720 107.125 ;
        RECT 84.660 105.965 85.410 106.135 ;
        RECT 84.655 105.295 84.985 105.795 ;
        RECT 85.155 105.465 85.410 105.965 ;
        RECT 85.625 105.295 85.855 106.435 ;
        RECT 86.025 105.465 86.355 106.445 ;
        RECT 87.550 106.540 87.835 106.870 ;
        RECT 86.525 105.295 86.735 106.435 ;
        RECT 87.550 106.395 87.720 106.540 ;
        RECT 87.055 106.225 87.720 106.395 ;
        RECT 88.005 106.370 88.175 107.170 ;
        RECT 88.805 107.120 89.095 107.845 ;
        RECT 89.270 107.295 89.525 107.585 ;
        RECT 89.695 107.465 90.025 107.845 ;
        RECT 89.270 107.125 90.020 107.295 ;
        RECT 87.055 105.465 87.225 106.225 ;
        RECT 87.405 105.295 87.735 106.055 ;
        RECT 87.905 105.465 88.175 106.370 ;
        RECT 88.805 105.295 89.095 106.460 ;
        RECT 89.270 106.305 89.620 106.955 ;
        RECT 89.790 106.135 90.020 107.125 ;
        RECT 89.270 105.965 90.020 106.135 ;
        RECT 89.270 105.465 89.525 105.965 ;
        RECT 89.695 105.295 90.025 105.795 ;
        RECT 90.195 105.465 90.365 107.585 ;
        RECT 90.725 107.485 91.055 107.845 ;
        RECT 91.225 107.455 91.720 107.625 ;
        RECT 91.925 107.455 92.780 107.625 ;
        RECT 90.595 106.265 91.055 107.315 ;
        RECT 90.535 105.480 90.860 106.265 ;
        RECT 91.225 106.095 91.395 107.455 ;
        RECT 91.565 106.545 91.915 107.165 ;
        RECT 92.085 106.945 92.440 107.165 ;
        RECT 92.085 106.355 92.255 106.945 ;
        RECT 92.610 106.745 92.780 107.455 ;
        RECT 93.655 107.385 93.985 107.845 ;
        RECT 94.195 107.485 94.545 107.655 ;
        RECT 92.985 106.915 93.775 107.165 ;
        RECT 94.195 107.095 94.455 107.485 ;
        RECT 94.765 107.395 95.715 107.675 ;
        RECT 95.885 107.405 96.075 107.845 ;
        RECT 96.245 107.465 97.315 107.635 ;
        RECT 93.945 106.745 94.115 106.925 ;
        RECT 91.225 105.925 91.620 106.095 ;
        RECT 91.790 105.965 92.255 106.355 ;
        RECT 92.425 106.575 94.115 106.745 ;
        RECT 91.450 105.795 91.620 105.925 ;
        RECT 92.425 105.795 92.595 106.575 ;
        RECT 94.285 106.405 94.455 107.095 ;
        RECT 92.955 106.235 94.455 106.405 ;
        RECT 94.645 106.435 94.855 107.225 ;
        RECT 95.025 106.605 95.375 107.225 ;
        RECT 95.545 106.615 95.715 107.395 ;
        RECT 96.245 107.235 96.415 107.465 ;
        RECT 95.885 107.065 96.415 107.235 ;
        RECT 95.885 106.785 96.105 107.065 ;
        RECT 96.585 106.895 96.825 107.295 ;
        RECT 95.545 106.445 95.950 106.615 ;
        RECT 96.285 106.525 96.825 106.895 ;
        RECT 96.995 107.110 97.315 107.465 ;
        RECT 96.995 106.855 97.320 107.110 ;
        RECT 97.515 107.035 97.685 107.845 ;
        RECT 97.855 107.195 98.185 107.675 ;
        RECT 98.355 107.375 98.525 107.845 ;
        RECT 98.695 107.195 99.025 107.675 ;
        RECT 99.195 107.375 99.365 107.845 ;
        RECT 100.615 107.375 100.785 107.845 ;
        RECT 100.955 107.195 101.285 107.675 ;
        RECT 101.455 107.375 101.625 107.845 ;
        RECT 101.795 107.195 102.125 107.675 ;
        RECT 97.855 107.025 99.620 107.195 ;
        RECT 96.995 106.645 99.025 106.855 ;
        RECT 96.995 106.635 97.340 106.645 ;
        RECT 94.645 106.275 95.320 106.435 ;
        RECT 95.780 106.355 95.950 106.445 ;
        RECT 94.645 106.265 95.610 106.275 ;
        RECT 94.285 106.095 94.455 106.235 ;
        RECT 91.030 105.295 91.280 105.755 ;
        RECT 91.450 105.465 91.700 105.795 ;
        RECT 91.915 105.465 92.595 105.795 ;
        RECT 92.765 105.895 93.840 106.065 ;
        RECT 94.285 105.925 94.845 106.095 ;
        RECT 95.150 105.975 95.610 106.265 ;
        RECT 95.780 106.185 97.000 106.355 ;
        RECT 92.765 105.555 92.935 105.895 ;
        RECT 93.170 105.295 93.500 105.725 ;
        RECT 93.670 105.555 93.840 105.895 ;
        RECT 94.135 105.295 94.505 105.755 ;
        RECT 94.675 105.465 94.845 105.925 ;
        RECT 95.780 105.805 95.950 106.185 ;
        RECT 97.170 106.015 97.340 106.635 ;
        RECT 99.210 106.475 99.620 107.025 ;
        RECT 95.080 105.465 95.950 105.805 ;
        RECT 96.540 105.845 97.340 106.015 ;
        RECT 96.120 105.295 96.370 105.755 ;
        RECT 96.540 105.555 96.710 105.845 ;
        RECT 96.890 105.295 97.220 105.675 ;
        RECT 97.515 105.295 97.685 106.355 ;
        RECT 97.895 106.305 99.620 106.475 ;
        RECT 100.360 107.025 102.125 107.195 ;
        RECT 102.295 107.035 102.465 107.845 ;
        RECT 102.665 107.465 103.735 107.635 ;
        RECT 102.665 107.110 102.985 107.465 ;
        RECT 100.360 106.475 100.770 107.025 ;
        RECT 102.660 106.855 102.985 107.110 ;
        RECT 100.955 106.645 102.985 106.855 ;
        RECT 102.640 106.635 102.985 106.645 ;
        RECT 103.155 106.895 103.395 107.295 ;
        RECT 103.565 107.235 103.735 107.465 ;
        RECT 103.905 107.405 104.095 107.845 ;
        RECT 104.265 107.395 105.215 107.675 ;
        RECT 105.435 107.485 105.785 107.655 ;
        RECT 103.565 107.065 104.095 107.235 ;
        RECT 100.360 106.305 102.085 106.475 ;
        RECT 97.895 105.465 98.185 106.305 ;
        RECT 98.355 105.295 98.525 106.135 ;
        RECT 98.735 105.465 98.985 106.305 ;
        RECT 99.195 105.295 99.365 106.135 ;
        RECT 100.615 105.295 100.785 106.135 ;
        RECT 100.995 105.465 101.245 106.305 ;
        RECT 101.455 105.295 101.625 106.135 ;
        RECT 101.795 105.465 102.085 106.305 ;
        RECT 102.295 105.295 102.465 106.355 ;
        RECT 102.640 106.015 102.810 106.635 ;
        RECT 103.155 106.525 103.695 106.895 ;
        RECT 103.875 106.785 104.095 107.065 ;
        RECT 104.265 106.615 104.435 107.395 ;
        RECT 104.030 106.445 104.435 106.615 ;
        RECT 104.605 106.605 104.955 107.225 ;
        RECT 104.030 106.355 104.200 106.445 ;
        RECT 105.125 106.435 105.335 107.225 ;
        RECT 102.980 106.185 104.200 106.355 ;
        RECT 104.660 106.275 105.335 106.435 ;
        RECT 102.640 105.845 103.440 106.015 ;
        RECT 102.760 105.295 103.090 105.675 ;
        RECT 103.270 105.555 103.440 105.845 ;
        RECT 104.030 105.805 104.200 106.185 ;
        RECT 104.370 106.265 105.335 106.275 ;
        RECT 105.525 107.095 105.785 107.485 ;
        RECT 105.995 107.385 106.325 107.845 ;
        RECT 107.200 107.455 108.055 107.625 ;
        RECT 108.260 107.455 108.755 107.625 ;
        RECT 108.925 107.485 109.255 107.845 ;
        RECT 105.525 106.405 105.695 107.095 ;
        RECT 105.865 106.745 106.035 106.925 ;
        RECT 106.205 106.915 106.995 107.165 ;
        RECT 107.200 106.745 107.370 107.455 ;
        RECT 107.540 106.945 107.895 107.165 ;
        RECT 105.865 106.575 107.555 106.745 ;
        RECT 104.370 105.975 104.830 106.265 ;
        RECT 105.525 106.235 107.025 106.405 ;
        RECT 105.525 106.095 105.695 106.235 ;
        RECT 105.135 105.925 105.695 106.095 ;
        RECT 103.610 105.295 103.860 105.755 ;
        RECT 104.030 105.465 104.900 105.805 ;
        RECT 105.135 105.465 105.305 105.925 ;
        RECT 106.140 105.895 107.215 106.065 ;
        RECT 105.475 105.295 105.845 105.755 ;
        RECT 106.140 105.555 106.310 105.895 ;
        RECT 106.480 105.295 106.810 105.725 ;
        RECT 107.045 105.555 107.215 105.895 ;
        RECT 107.385 105.795 107.555 106.575 ;
        RECT 107.725 106.355 107.895 106.945 ;
        RECT 108.065 106.545 108.415 107.165 ;
        RECT 107.725 105.965 108.190 106.355 ;
        RECT 108.585 106.095 108.755 107.455 ;
        RECT 108.925 106.265 109.385 107.315 ;
        RECT 108.360 105.925 108.755 106.095 ;
        RECT 108.360 105.795 108.530 105.925 ;
        RECT 107.385 105.465 108.065 105.795 ;
        RECT 108.280 105.465 108.530 105.795 ;
        RECT 108.700 105.295 108.950 105.755 ;
        RECT 109.120 105.480 109.445 106.265 ;
        RECT 109.615 105.465 109.785 107.585 ;
        RECT 109.955 107.465 110.285 107.845 ;
        RECT 110.455 107.295 110.710 107.585 ;
        RECT 109.960 107.125 110.710 107.295 ;
        RECT 109.960 106.135 110.190 107.125 ;
        RECT 110.945 107.025 111.155 107.845 ;
        RECT 111.325 107.045 111.655 107.675 ;
        RECT 110.360 106.305 110.710 106.955 ;
        RECT 111.325 106.445 111.575 107.045 ;
        RECT 111.825 107.025 112.055 107.845 ;
        RECT 113.225 107.025 113.455 107.845 ;
        RECT 113.625 107.045 113.955 107.675 ;
        RECT 111.745 106.605 112.075 106.855 ;
        RECT 113.205 106.605 113.535 106.855 ;
        RECT 113.705 106.445 113.955 107.045 ;
        RECT 114.125 107.025 114.335 107.845 ;
        RECT 114.565 107.120 114.855 107.845 ;
        RECT 116.255 107.375 116.425 107.845 ;
        RECT 116.595 107.195 116.925 107.675 ;
        RECT 117.095 107.375 117.265 107.845 ;
        RECT 117.435 107.195 117.765 107.675 ;
        RECT 116.000 107.025 117.765 107.195 ;
        RECT 117.935 107.035 118.105 107.845 ;
        RECT 118.305 107.465 119.375 107.635 ;
        RECT 118.305 107.110 118.625 107.465 ;
        RECT 116.000 106.475 116.410 107.025 ;
        RECT 118.300 106.855 118.625 107.110 ;
        RECT 116.595 106.645 118.625 106.855 ;
        RECT 118.280 106.635 118.625 106.645 ;
        RECT 118.795 106.895 119.035 107.295 ;
        RECT 119.205 107.235 119.375 107.465 ;
        RECT 119.545 107.405 119.735 107.845 ;
        RECT 119.905 107.395 120.855 107.675 ;
        RECT 121.075 107.485 121.425 107.655 ;
        RECT 119.205 107.065 119.735 107.235 ;
        RECT 109.960 105.965 110.710 106.135 ;
        RECT 109.955 105.295 110.285 105.795 ;
        RECT 110.455 105.465 110.710 105.965 ;
        RECT 110.945 105.295 111.155 106.435 ;
        RECT 111.325 105.465 111.655 106.445 ;
        RECT 111.825 105.295 112.055 106.435 ;
        RECT 113.225 105.295 113.455 106.435 ;
        RECT 113.625 105.465 113.955 106.445 ;
        RECT 114.125 105.295 114.335 106.435 ;
        RECT 114.565 105.295 114.855 106.460 ;
        RECT 116.000 106.305 117.725 106.475 ;
        RECT 116.255 105.295 116.425 106.135 ;
        RECT 116.635 105.465 116.885 106.305 ;
        RECT 117.095 105.295 117.265 106.135 ;
        RECT 117.435 105.465 117.725 106.305 ;
        RECT 117.935 105.295 118.105 106.355 ;
        RECT 118.280 106.015 118.450 106.635 ;
        RECT 118.795 106.525 119.335 106.895 ;
        RECT 119.515 106.785 119.735 107.065 ;
        RECT 119.905 106.615 120.075 107.395 ;
        RECT 119.670 106.445 120.075 106.615 ;
        RECT 120.245 106.605 120.595 107.225 ;
        RECT 119.670 106.355 119.840 106.445 ;
        RECT 120.765 106.435 120.975 107.225 ;
        RECT 118.620 106.185 119.840 106.355 ;
        RECT 120.300 106.275 120.975 106.435 ;
        RECT 118.280 105.845 119.080 106.015 ;
        RECT 118.400 105.295 118.730 105.675 ;
        RECT 118.910 105.555 119.080 105.845 ;
        RECT 119.670 105.805 119.840 106.185 ;
        RECT 120.010 106.265 120.975 106.275 ;
        RECT 121.165 107.095 121.425 107.485 ;
        RECT 121.635 107.385 121.965 107.845 ;
        RECT 122.840 107.455 123.695 107.625 ;
        RECT 123.900 107.455 124.395 107.625 ;
        RECT 124.565 107.485 124.895 107.845 ;
        RECT 121.165 106.405 121.335 107.095 ;
        RECT 121.505 106.745 121.675 106.925 ;
        RECT 121.845 106.915 122.635 107.165 ;
        RECT 122.840 106.745 123.010 107.455 ;
        RECT 123.180 106.945 123.535 107.165 ;
        RECT 121.505 106.575 123.195 106.745 ;
        RECT 120.010 105.975 120.470 106.265 ;
        RECT 121.165 106.235 122.665 106.405 ;
        RECT 121.165 106.095 121.335 106.235 ;
        RECT 120.775 105.925 121.335 106.095 ;
        RECT 119.250 105.295 119.500 105.755 ;
        RECT 119.670 105.465 120.540 105.805 ;
        RECT 120.775 105.465 120.945 105.925 ;
        RECT 121.780 105.895 122.855 106.065 ;
        RECT 121.115 105.295 121.485 105.755 ;
        RECT 121.780 105.555 121.950 105.895 ;
        RECT 122.120 105.295 122.450 105.725 ;
        RECT 122.685 105.555 122.855 105.895 ;
        RECT 123.025 105.795 123.195 106.575 ;
        RECT 123.365 106.355 123.535 106.945 ;
        RECT 123.705 106.545 124.055 107.165 ;
        RECT 123.365 105.965 123.830 106.355 ;
        RECT 124.225 106.095 124.395 107.455 ;
        RECT 124.565 106.265 125.025 107.315 ;
        RECT 124.000 105.925 124.395 106.095 ;
        RECT 124.000 105.795 124.170 105.925 ;
        RECT 123.025 105.465 123.705 105.795 ;
        RECT 123.920 105.465 124.170 105.795 ;
        RECT 124.340 105.295 124.590 105.755 ;
        RECT 124.760 105.480 125.085 106.265 ;
        RECT 125.255 105.465 125.425 107.585 ;
        RECT 125.595 107.465 125.925 107.845 ;
        RECT 126.095 107.295 126.350 107.585 ;
        RECT 125.600 107.125 126.350 107.295 ;
        RECT 125.600 106.135 125.830 107.125 ;
        RECT 126.525 107.095 127.735 107.845 ;
        RECT 126.000 106.305 126.350 106.955 ;
        RECT 126.525 106.385 127.045 106.925 ;
        RECT 127.215 106.555 127.735 107.095 ;
        RECT 125.600 105.965 126.350 106.135 ;
        RECT 125.595 105.295 125.925 105.795 ;
        RECT 126.095 105.465 126.350 105.965 ;
        RECT 126.525 105.295 127.735 106.385 ;
        RECT 14.660 105.125 127.820 105.295 ;
        RECT 14.745 104.035 15.955 105.125 ;
        RECT 14.745 103.325 15.265 103.865 ;
        RECT 15.435 103.495 15.955 104.035 ;
        RECT 16.125 104.035 18.715 105.125 ;
        RECT 18.890 104.690 24.235 105.125 ;
        RECT 16.125 103.515 17.335 104.035 ;
        RECT 17.505 103.345 18.715 103.865 ;
        RECT 20.480 103.440 20.830 104.690 ;
        RECT 24.405 103.960 24.695 105.125 ;
        RECT 24.865 104.035 26.075 105.125 ;
        RECT 14.745 102.575 15.955 103.325 ;
        RECT 16.125 102.575 18.715 103.345 ;
        RECT 22.310 103.120 22.650 103.950 ;
        RECT 24.865 103.495 25.385 104.035 ;
        RECT 26.285 103.985 26.515 105.125 ;
        RECT 26.685 103.975 27.015 104.955 ;
        RECT 27.185 103.985 27.395 105.125 ;
        RECT 27.625 104.050 27.895 104.955 ;
        RECT 28.065 104.365 28.395 105.125 ;
        RECT 28.575 104.195 28.745 104.955 ;
        RECT 29.315 104.285 29.485 105.125 ;
        RECT 25.555 103.325 26.075 103.865 ;
        RECT 26.265 103.565 26.595 103.815 ;
        RECT 18.890 102.575 24.235 103.120 ;
        RECT 24.405 102.575 24.695 103.300 ;
        RECT 24.865 102.575 26.075 103.325 ;
        RECT 26.285 102.575 26.515 103.395 ;
        RECT 26.765 103.375 27.015 103.975 ;
        RECT 26.685 102.745 27.015 103.375 ;
        RECT 27.185 102.575 27.395 103.395 ;
        RECT 27.625 103.250 27.795 104.050 ;
        RECT 28.080 104.025 28.745 104.195 ;
        RECT 29.695 104.115 29.945 104.955 ;
        RECT 30.155 104.285 30.325 105.125 ;
        RECT 30.495 104.115 30.785 104.955 ;
        RECT 28.080 103.880 28.250 104.025 ;
        RECT 27.965 103.550 28.250 103.880 ;
        RECT 29.060 103.945 30.785 104.115 ;
        RECT 30.995 104.065 31.165 105.125 ;
        RECT 31.460 104.745 31.790 105.125 ;
        RECT 31.970 104.575 32.140 104.865 ;
        RECT 32.310 104.665 32.560 105.125 ;
        RECT 31.340 104.405 32.140 104.575 ;
        RECT 32.730 104.615 33.600 104.955 ;
        RECT 28.080 103.295 28.250 103.550 ;
        RECT 28.485 103.475 28.815 103.845 ;
        RECT 29.060 103.395 29.470 103.945 ;
        RECT 31.340 103.785 31.510 104.405 ;
        RECT 32.730 104.235 32.900 104.615 ;
        RECT 33.835 104.495 34.005 104.955 ;
        RECT 34.175 104.665 34.545 105.125 ;
        RECT 34.840 104.525 35.010 104.865 ;
        RECT 35.180 104.695 35.510 105.125 ;
        RECT 35.745 104.525 35.915 104.865 ;
        RECT 31.680 104.065 32.900 104.235 ;
        RECT 33.070 104.155 33.530 104.445 ;
        RECT 33.835 104.325 34.395 104.495 ;
        RECT 34.840 104.355 35.915 104.525 ;
        RECT 36.085 104.625 36.765 104.955 ;
        RECT 36.980 104.625 37.230 104.955 ;
        RECT 37.400 104.665 37.650 105.125 ;
        RECT 34.225 104.185 34.395 104.325 ;
        RECT 33.070 104.145 34.035 104.155 ;
        RECT 32.730 103.975 32.900 104.065 ;
        RECT 33.360 103.985 34.035 104.145 ;
        RECT 31.340 103.775 31.685 103.785 ;
        RECT 29.655 103.565 31.685 103.775 ;
        RECT 27.625 102.745 27.885 103.250 ;
        RECT 28.080 103.125 28.745 103.295 ;
        RECT 29.060 103.225 30.825 103.395 ;
        RECT 28.065 102.575 28.395 102.955 ;
        RECT 28.575 102.745 28.745 103.125 ;
        RECT 29.315 102.575 29.485 103.045 ;
        RECT 29.655 102.745 29.985 103.225 ;
        RECT 30.155 102.575 30.325 103.045 ;
        RECT 30.495 102.745 30.825 103.225 ;
        RECT 30.995 102.575 31.165 103.385 ;
        RECT 31.360 103.310 31.685 103.565 ;
        RECT 31.365 102.955 31.685 103.310 ;
        RECT 31.855 103.525 32.395 103.895 ;
        RECT 32.730 103.805 33.135 103.975 ;
        RECT 31.855 103.125 32.095 103.525 ;
        RECT 32.575 103.355 32.795 103.635 ;
        RECT 32.265 103.185 32.795 103.355 ;
        RECT 32.265 102.955 32.435 103.185 ;
        RECT 32.965 103.025 33.135 103.805 ;
        RECT 33.305 103.195 33.655 103.815 ;
        RECT 33.825 103.195 34.035 103.985 ;
        RECT 34.225 104.015 35.725 104.185 ;
        RECT 34.225 103.325 34.395 104.015 ;
        RECT 36.085 103.845 36.255 104.625 ;
        RECT 37.060 104.495 37.230 104.625 ;
        RECT 34.565 103.675 36.255 103.845 ;
        RECT 36.425 104.065 36.890 104.455 ;
        RECT 37.060 104.325 37.455 104.495 ;
        RECT 34.565 103.495 34.735 103.675 ;
        RECT 31.365 102.785 32.435 102.955 ;
        RECT 32.605 102.575 32.795 103.015 ;
        RECT 32.965 102.745 33.915 103.025 ;
        RECT 34.225 102.935 34.485 103.325 ;
        RECT 34.905 103.255 35.695 103.505 ;
        RECT 34.135 102.765 34.485 102.935 ;
        RECT 34.695 102.575 35.025 103.035 ;
        RECT 35.900 102.965 36.070 103.675 ;
        RECT 36.425 103.475 36.595 104.065 ;
        RECT 36.240 103.255 36.595 103.475 ;
        RECT 36.765 103.255 37.115 103.875 ;
        RECT 37.285 102.965 37.455 104.325 ;
        RECT 37.820 104.155 38.145 104.940 ;
        RECT 37.625 103.105 38.085 104.155 ;
        RECT 35.900 102.795 36.755 102.965 ;
        RECT 36.960 102.795 37.455 102.965 ;
        RECT 37.625 102.575 37.955 102.935 ;
        RECT 38.315 102.835 38.485 104.955 ;
        RECT 38.655 104.625 38.985 105.125 ;
        RECT 39.155 104.455 39.410 104.955 ;
        RECT 38.660 104.285 39.410 104.455 ;
        RECT 39.590 104.455 39.845 104.955 ;
        RECT 40.015 104.625 40.345 105.125 ;
        RECT 39.590 104.285 40.340 104.455 ;
        RECT 38.660 103.295 38.890 104.285 ;
        RECT 39.060 103.465 39.410 104.115 ;
        RECT 39.590 103.465 39.940 104.115 ;
        RECT 40.110 103.295 40.340 104.285 ;
        RECT 38.660 103.125 39.410 103.295 ;
        RECT 38.655 102.575 38.985 102.955 ;
        RECT 39.155 102.835 39.410 103.125 ;
        RECT 39.590 103.125 40.340 103.295 ;
        RECT 39.590 102.835 39.845 103.125 ;
        RECT 40.015 102.575 40.345 102.955 ;
        RECT 40.515 102.835 40.685 104.955 ;
        RECT 40.855 104.155 41.180 104.940 ;
        RECT 41.350 104.665 41.600 105.125 ;
        RECT 41.770 104.625 42.020 104.955 ;
        RECT 42.235 104.625 42.915 104.955 ;
        RECT 41.770 104.495 41.940 104.625 ;
        RECT 41.545 104.325 41.940 104.495 ;
        RECT 40.915 103.105 41.375 104.155 ;
        RECT 41.545 102.965 41.715 104.325 ;
        RECT 42.110 104.065 42.575 104.455 ;
        RECT 41.885 103.255 42.235 103.875 ;
        RECT 42.405 103.475 42.575 104.065 ;
        RECT 42.745 103.845 42.915 104.625 ;
        RECT 43.085 104.525 43.255 104.865 ;
        RECT 43.490 104.695 43.820 105.125 ;
        RECT 43.990 104.525 44.160 104.865 ;
        RECT 44.455 104.665 44.825 105.125 ;
        RECT 43.085 104.355 44.160 104.525 ;
        RECT 44.995 104.495 45.165 104.955 ;
        RECT 45.400 104.615 46.270 104.955 ;
        RECT 46.440 104.665 46.690 105.125 ;
        RECT 44.605 104.325 45.165 104.495 ;
        RECT 44.605 104.185 44.775 104.325 ;
        RECT 43.275 104.015 44.775 104.185 ;
        RECT 45.470 104.155 45.930 104.445 ;
        RECT 42.745 103.675 44.435 103.845 ;
        RECT 42.405 103.255 42.760 103.475 ;
        RECT 42.930 102.965 43.100 103.675 ;
        RECT 43.305 103.255 44.095 103.505 ;
        RECT 44.265 103.495 44.435 103.675 ;
        RECT 44.605 103.325 44.775 104.015 ;
        RECT 41.045 102.575 41.375 102.935 ;
        RECT 41.545 102.795 42.040 102.965 ;
        RECT 42.245 102.795 43.100 102.965 ;
        RECT 43.975 102.575 44.305 103.035 ;
        RECT 44.515 102.935 44.775 103.325 ;
        RECT 44.965 104.145 45.930 104.155 ;
        RECT 46.100 104.235 46.270 104.615 ;
        RECT 46.860 104.575 47.030 104.865 ;
        RECT 47.210 104.745 47.540 105.125 ;
        RECT 46.860 104.405 47.660 104.575 ;
        RECT 44.965 103.985 45.640 104.145 ;
        RECT 46.100 104.065 47.320 104.235 ;
        RECT 44.965 103.195 45.175 103.985 ;
        RECT 46.100 103.975 46.270 104.065 ;
        RECT 45.345 103.195 45.695 103.815 ;
        RECT 45.865 103.805 46.270 103.975 ;
        RECT 45.865 103.025 46.035 103.805 ;
        RECT 46.205 103.355 46.425 103.635 ;
        RECT 46.605 103.525 47.145 103.895 ;
        RECT 47.490 103.785 47.660 104.405 ;
        RECT 47.835 104.065 48.005 105.125 ;
        RECT 48.215 104.115 48.505 104.955 ;
        RECT 48.675 104.285 48.845 105.125 ;
        RECT 49.055 104.115 49.305 104.955 ;
        RECT 49.515 104.285 49.685 105.125 ;
        RECT 48.215 103.945 49.940 104.115 ;
        RECT 50.165 103.960 50.455 105.125 ;
        RECT 50.625 104.035 51.835 105.125 ;
        RECT 52.005 104.035 55.515 105.125 ;
        RECT 46.205 103.185 46.735 103.355 ;
        RECT 44.515 102.765 44.865 102.935 ;
        RECT 45.085 102.745 46.035 103.025 ;
        RECT 46.205 102.575 46.395 103.015 ;
        RECT 46.565 102.955 46.735 103.185 ;
        RECT 46.905 103.125 47.145 103.525 ;
        RECT 47.315 103.775 47.660 103.785 ;
        RECT 47.315 103.565 49.345 103.775 ;
        RECT 47.315 103.310 47.640 103.565 ;
        RECT 49.530 103.395 49.940 103.945 ;
        RECT 50.625 103.495 51.145 104.035 ;
        RECT 47.315 102.955 47.635 103.310 ;
        RECT 46.565 102.785 47.635 102.955 ;
        RECT 47.835 102.575 48.005 103.385 ;
        RECT 48.175 103.225 49.940 103.395 ;
        RECT 51.315 103.325 51.835 103.865 ;
        RECT 52.005 103.515 53.695 104.035 ;
        RECT 55.745 103.985 55.955 105.125 ;
        RECT 56.125 103.975 56.455 104.955 ;
        RECT 56.625 103.985 56.855 105.125 ;
        RECT 57.065 104.035 58.275 105.125 ;
        RECT 58.755 104.285 58.925 105.125 ;
        RECT 59.135 104.115 59.385 104.955 ;
        RECT 59.595 104.285 59.765 105.125 ;
        RECT 59.935 104.115 60.225 104.955 ;
        RECT 53.865 103.345 55.515 103.865 ;
        RECT 48.175 102.745 48.505 103.225 ;
        RECT 48.675 102.575 48.845 103.045 ;
        RECT 49.015 102.745 49.345 103.225 ;
        RECT 49.515 102.575 49.685 103.045 ;
        RECT 50.165 102.575 50.455 103.300 ;
        RECT 50.625 102.575 51.835 103.325 ;
        RECT 52.005 102.575 55.515 103.345 ;
        RECT 55.745 102.575 55.955 103.395 ;
        RECT 56.125 103.375 56.375 103.975 ;
        RECT 56.545 103.565 56.875 103.815 ;
        RECT 57.065 103.495 57.585 104.035 ;
        RECT 58.500 103.945 60.225 104.115 ;
        RECT 60.435 104.065 60.605 105.125 ;
        RECT 60.900 104.745 61.230 105.125 ;
        RECT 61.410 104.575 61.580 104.865 ;
        RECT 61.750 104.665 62.000 105.125 ;
        RECT 60.780 104.405 61.580 104.575 ;
        RECT 62.170 104.615 63.040 104.955 ;
        RECT 56.125 102.745 56.455 103.375 ;
        RECT 56.625 102.575 56.855 103.395 ;
        RECT 57.755 103.325 58.275 103.865 ;
        RECT 57.065 102.575 58.275 103.325 ;
        RECT 58.500 103.395 58.910 103.945 ;
        RECT 60.780 103.785 60.950 104.405 ;
        RECT 62.170 104.235 62.340 104.615 ;
        RECT 63.275 104.495 63.445 104.955 ;
        RECT 63.615 104.665 63.985 105.125 ;
        RECT 64.280 104.525 64.450 104.865 ;
        RECT 64.620 104.695 64.950 105.125 ;
        RECT 65.185 104.525 65.355 104.865 ;
        RECT 61.120 104.065 62.340 104.235 ;
        RECT 62.510 104.155 62.970 104.445 ;
        RECT 63.275 104.325 63.835 104.495 ;
        RECT 64.280 104.355 65.355 104.525 ;
        RECT 65.525 104.625 66.205 104.955 ;
        RECT 66.420 104.625 66.670 104.955 ;
        RECT 66.840 104.665 67.090 105.125 ;
        RECT 63.665 104.185 63.835 104.325 ;
        RECT 62.510 104.145 63.475 104.155 ;
        RECT 62.170 103.975 62.340 104.065 ;
        RECT 62.800 103.985 63.475 104.145 ;
        RECT 60.780 103.775 61.125 103.785 ;
        RECT 59.095 103.565 61.125 103.775 ;
        RECT 58.500 103.225 60.265 103.395 ;
        RECT 58.755 102.575 58.925 103.045 ;
        RECT 59.095 102.745 59.425 103.225 ;
        RECT 59.595 102.575 59.765 103.045 ;
        RECT 59.935 102.745 60.265 103.225 ;
        RECT 60.435 102.575 60.605 103.385 ;
        RECT 60.800 103.310 61.125 103.565 ;
        RECT 60.805 102.955 61.125 103.310 ;
        RECT 61.295 103.525 61.835 103.895 ;
        RECT 62.170 103.805 62.575 103.975 ;
        RECT 61.295 103.125 61.535 103.525 ;
        RECT 62.015 103.355 62.235 103.635 ;
        RECT 61.705 103.185 62.235 103.355 ;
        RECT 61.705 102.955 61.875 103.185 ;
        RECT 62.405 103.025 62.575 103.805 ;
        RECT 62.745 103.195 63.095 103.815 ;
        RECT 63.265 103.195 63.475 103.985 ;
        RECT 63.665 104.015 65.165 104.185 ;
        RECT 63.665 103.325 63.835 104.015 ;
        RECT 65.525 103.845 65.695 104.625 ;
        RECT 66.500 104.495 66.670 104.625 ;
        RECT 64.005 103.675 65.695 103.845 ;
        RECT 65.865 104.065 66.330 104.455 ;
        RECT 66.500 104.325 66.895 104.495 ;
        RECT 64.005 103.495 64.175 103.675 ;
        RECT 60.805 102.785 61.875 102.955 ;
        RECT 62.045 102.575 62.235 103.015 ;
        RECT 62.405 102.745 63.355 103.025 ;
        RECT 63.665 102.935 63.925 103.325 ;
        RECT 64.345 103.255 65.135 103.505 ;
        RECT 63.575 102.765 63.925 102.935 ;
        RECT 64.135 102.575 64.465 103.035 ;
        RECT 65.340 102.965 65.510 103.675 ;
        RECT 65.865 103.475 66.035 104.065 ;
        RECT 65.680 103.255 66.035 103.475 ;
        RECT 66.205 103.255 66.555 103.875 ;
        RECT 66.725 102.965 66.895 104.325 ;
        RECT 67.260 104.155 67.585 104.940 ;
        RECT 67.065 103.105 67.525 104.155 ;
        RECT 65.340 102.795 66.195 102.965 ;
        RECT 66.400 102.795 66.895 102.965 ;
        RECT 67.065 102.575 67.395 102.935 ;
        RECT 67.755 102.835 67.925 104.955 ;
        RECT 68.095 104.625 68.425 105.125 ;
        RECT 68.595 104.455 68.850 104.955 ;
        RECT 68.100 104.285 68.850 104.455 ;
        RECT 68.100 103.295 68.330 104.285 ;
        RECT 68.500 103.465 68.850 104.115 ;
        RECT 69.025 104.035 70.235 105.125 ;
        RECT 70.410 104.690 75.755 105.125 ;
        RECT 69.025 103.495 69.545 104.035 ;
        RECT 69.715 103.325 70.235 103.865 ;
        RECT 72.000 103.440 72.350 104.690 ;
        RECT 75.925 103.960 76.215 105.125 ;
        RECT 76.695 104.285 76.865 105.125 ;
        RECT 77.075 104.115 77.325 104.955 ;
        RECT 77.535 104.285 77.705 105.125 ;
        RECT 77.875 104.115 78.165 104.955 ;
        RECT 68.100 103.125 68.850 103.295 ;
        RECT 68.095 102.575 68.425 102.955 ;
        RECT 68.595 102.835 68.850 103.125 ;
        RECT 69.025 102.575 70.235 103.325 ;
        RECT 73.830 103.120 74.170 103.950 ;
        RECT 76.440 103.945 78.165 104.115 ;
        RECT 78.375 104.065 78.545 105.125 ;
        RECT 78.840 104.745 79.170 105.125 ;
        RECT 79.350 104.575 79.520 104.865 ;
        RECT 79.690 104.665 79.940 105.125 ;
        RECT 78.720 104.405 79.520 104.575 ;
        RECT 80.110 104.615 80.980 104.955 ;
        RECT 76.440 103.395 76.850 103.945 ;
        RECT 78.720 103.785 78.890 104.405 ;
        RECT 80.110 104.235 80.280 104.615 ;
        RECT 81.215 104.495 81.385 104.955 ;
        RECT 81.555 104.665 81.925 105.125 ;
        RECT 82.220 104.525 82.390 104.865 ;
        RECT 82.560 104.695 82.890 105.125 ;
        RECT 83.125 104.525 83.295 104.865 ;
        RECT 79.060 104.065 80.280 104.235 ;
        RECT 80.450 104.155 80.910 104.445 ;
        RECT 81.215 104.325 81.775 104.495 ;
        RECT 82.220 104.355 83.295 104.525 ;
        RECT 83.465 104.625 84.145 104.955 ;
        RECT 84.360 104.625 84.610 104.955 ;
        RECT 84.780 104.665 85.030 105.125 ;
        RECT 81.605 104.185 81.775 104.325 ;
        RECT 80.450 104.145 81.415 104.155 ;
        RECT 80.110 103.975 80.280 104.065 ;
        RECT 80.740 103.985 81.415 104.145 ;
        RECT 78.720 103.775 79.065 103.785 ;
        RECT 77.035 103.565 79.065 103.775 ;
        RECT 70.410 102.575 75.755 103.120 ;
        RECT 75.925 102.575 76.215 103.300 ;
        RECT 76.440 103.225 78.205 103.395 ;
        RECT 76.695 102.575 76.865 103.045 ;
        RECT 77.035 102.745 77.365 103.225 ;
        RECT 77.535 102.575 77.705 103.045 ;
        RECT 77.875 102.745 78.205 103.225 ;
        RECT 78.375 102.575 78.545 103.385 ;
        RECT 78.740 103.310 79.065 103.565 ;
        RECT 78.745 102.955 79.065 103.310 ;
        RECT 79.235 103.525 79.775 103.895 ;
        RECT 80.110 103.805 80.515 103.975 ;
        RECT 79.235 103.125 79.475 103.525 ;
        RECT 79.955 103.355 80.175 103.635 ;
        RECT 79.645 103.185 80.175 103.355 ;
        RECT 79.645 102.955 79.815 103.185 ;
        RECT 80.345 103.025 80.515 103.805 ;
        RECT 80.685 103.195 81.035 103.815 ;
        RECT 81.205 103.195 81.415 103.985 ;
        RECT 81.605 104.015 83.105 104.185 ;
        RECT 81.605 103.325 81.775 104.015 ;
        RECT 83.465 103.845 83.635 104.625 ;
        RECT 84.440 104.495 84.610 104.625 ;
        RECT 81.945 103.675 83.635 103.845 ;
        RECT 83.805 104.065 84.270 104.455 ;
        RECT 84.440 104.325 84.835 104.495 ;
        RECT 81.945 103.495 82.115 103.675 ;
        RECT 78.745 102.785 79.815 102.955 ;
        RECT 79.985 102.575 80.175 103.015 ;
        RECT 80.345 102.745 81.295 103.025 ;
        RECT 81.605 102.935 81.865 103.325 ;
        RECT 82.285 103.255 83.075 103.505 ;
        RECT 81.515 102.765 81.865 102.935 ;
        RECT 82.075 102.575 82.405 103.035 ;
        RECT 83.280 102.965 83.450 103.675 ;
        RECT 83.805 103.475 83.975 104.065 ;
        RECT 83.620 103.255 83.975 103.475 ;
        RECT 84.145 103.255 84.495 103.875 ;
        RECT 84.665 102.965 84.835 104.325 ;
        RECT 85.200 104.155 85.525 104.940 ;
        RECT 85.005 103.105 85.465 104.155 ;
        RECT 83.280 102.795 84.135 102.965 ;
        RECT 84.340 102.795 84.835 102.965 ;
        RECT 85.005 102.575 85.335 102.935 ;
        RECT 85.695 102.835 85.865 104.955 ;
        RECT 86.035 104.625 86.365 105.125 ;
        RECT 86.535 104.455 86.790 104.955 ;
        RECT 86.040 104.285 86.790 104.455 ;
        RECT 87.275 104.285 87.445 105.125 ;
        RECT 86.040 103.295 86.270 104.285 ;
        RECT 87.655 104.115 87.905 104.955 ;
        RECT 88.115 104.285 88.285 105.125 ;
        RECT 88.455 104.115 88.745 104.955 ;
        RECT 86.440 103.465 86.790 104.115 ;
        RECT 87.020 103.945 88.745 104.115 ;
        RECT 88.955 104.065 89.125 105.125 ;
        RECT 89.420 104.745 89.750 105.125 ;
        RECT 89.930 104.575 90.100 104.865 ;
        RECT 90.270 104.665 90.520 105.125 ;
        RECT 89.300 104.405 90.100 104.575 ;
        RECT 90.690 104.615 91.560 104.955 ;
        RECT 87.020 103.395 87.430 103.945 ;
        RECT 89.300 103.785 89.470 104.405 ;
        RECT 90.690 104.235 90.860 104.615 ;
        RECT 91.795 104.495 91.965 104.955 ;
        RECT 92.135 104.665 92.505 105.125 ;
        RECT 92.800 104.525 92.970 104.865 ;
        RECT 93.140 104.695 93.470 105.125 ;
        RECT 93.705 104.525 93.875 104.865 ;
        RECT 89.640 104.065 90.860 104.235 ;
        RECT 91.030 104.155 91.490 104.445 ;
        RECT 91.795 104.325 92.355 104.495 ;
        RECT 92.800 104.355 93.875 104.525 ;
        RECT 94.045 104.625 94.725 104.955 ;
        RECT 94.940 104.625 95.190 104.955 ;
        RECT 95.360 104.665 95.610 105.125 ;
        RECT 92.185 104.185 92.355 104.325 ;
        RECT 91.030 104.145 91.995 104.155 ;
        RECT 90.690 103.975 90.860 104.065 ;
        RECT 91.320 103.985 91.995 104.145 ;
        RECT 89.300 103.775 89.645 103.785 ;
        RECT 87.615 103.565 89.645 103.775 ;
        RECT 86.040 103.125 86.790 103.295 ;
        RECT 87.020 103.225 88.785 103.395 ;
        RECT 86.035 102.575 86.365 102.955 ;
        RECT 86.535 102.835 86.790 103.125 ;
        RECT 87.275 102.575 87.445 103.045 ;
        RECT 87.615 102.745 87.945 103.225 ;
        RECT 88.115 102.575 88.285 103.045 ;
        RECT 88.455 102.745 88.785 103.225 ;
        RECT 88.955 102.575 89.125 103.385 ;
        RECT 89.320 103.310 89.645 103.565 ;
        RECT 89.325 102.955 89.645 103.310 ;
        RECT 89.815 103.525 90.355 103.895 ;
        RECT 90.690 103.805 91.095 103.975 ;
        RECT 89.815 103.125 90.055 103.525 ;
        RECT 90.535 103.355 90.755 103.635 ;
        RECT 90.225 103.185 90.755 103.355 ;
        RECT 90.225 102.955 90.395 103.185 ;
        RECT 90.925 103.025 91.095 103.805 ;
        RECT 91.265 103.195 91.615 103.815 ;
        RECT 91.785 103.195 91.995 103.985 ;
        RECT 92.185 104.015 93.685 104.185 ;
        RECT 92.185 103.325 92.355 104.015 ;
        RECT 94.045 103.845 94.215 104.625 ;
        RECT 95.020 104.495 95.190 104.625 ;
        RECT 92.525 103.675 94.215 103.845 ;
        RECT 94.385 104.065 94.850 104.455 ;
        RECT 95.020 104.325 95.415 104.495 ;
        RECT 92.525 103.495 92.695 103.675 ;
        RECT 89.325 102.785 90.395 102.955 ;
        RECT 90.565 102.575 90.755 103.015 ;
        RECT 90.925 102.745 91.875 103.025 ;
        RECT 92.185 102.935 92.445 103.325 ;
        RECT 92.865 103.255 93.655 103.505 ;
        RECT 92.095 102.765 92.445 102.935 ;
        RECT 92.655 102.575 92.985 103.035 ;
        RECT 93.860 102.965 94.030 103.675 ;
        RECT 94.385 103.475 94.555 104.065 ;
        RECT 94.200 103.255 94.555 103.475 ;
        RECT 94.725 103.255 95.075 103.875 ;
        RECT 95.245 102.965 95.415 104.325 ;
        RECT 95.780 104.155 96.105 104.940 ;
        RECT 95.585 103.105 96.045 104.155 ;
        RECT 93.860 102.795 94.715 102.965 ;
        RECT 94.920 102.795 95.415 102.965 ;
        RECT 95.585 102.575 95.915 102.935 ;
        RECT 96.275 102.835 96.445 104.955 ;
        RECT 96.615 104.625 96.945 105.125 ;
        RECT 97.115 104.455 97.370 104.955 ;
        RECT 96.620 104.285 97.370 104.455 ;
        RECT 96.620 103.295 96.850 104.285 ;
        RECT 97.020 103.465 97.370 104.115 ;
        RECT 98.525 103.985 98.735 105.125 ;
        RECT 98.905 103.975 99.235 104.955 ;
        RECT 99.405 103.985 99.635 105.125 ;
        RECT 99.845 104.035 101.515 105.125 ;
        RECT 96.620 103.125 97.370 103.295 ;
        RECT 96.615 102.575 96.945 102.955 ;
        RECT 97.115 102.835 97.370 103.125 ;
        RECT 98.525 102.575 98.735 103.395 ;
        RECT 98.905 103.375 99.155 103.975 ;
        RECT 99.325 103.565 99.655 103.815 ;
        RECT 99.845 103.515 100.595 104.035 ;
        RECT 101.685 103.960 101.975 105.125 ;
        RECT 102.145 104.035 103.355 105.125 ;
        RECT 103.530 104.455 103.785 104.955 ;
        RECT 103.955 104.625 104.285 105.125 ;
        RECT 103.530 104.285 104.280 104.455 ;
        RECT 98.905 102.745 99.235 103.375 ;
        RECT 99.405 102.575 99.635 103.395 ;
        RECT 100.765 103.345 101.515 103.865 ;
        RECT 102.145 103.495 102.665 104.035 ;
        RECT 99.845 102.575 101.515 103.345 ;
        RECT 102.835 103.325 103.355 103.865 ;
        RECT 103.530 103.465 103.880 104.115 ;
        RECT 101.685 102.575 101.975 103.300 ;
        RECT 102.145 102.575 103.355 103.325 ;
        RECT 104.050 103.295 104.280 104.285 ;
        RECT 103.530 103.125 104.280 103.295 ;
        RECT 103.530 102.835 103.785 103.125 ;
        RECT 103.955 102.575 104.285 102.955 ;
        RECT 104.455 102.835 104.625 104.955 ;
        RECT 104.795 104.155 105.120 104.940 ;
        RECT 105.290 104.665 105.540 105.125 ;
        RECT 105.710 104.625 105.960 104.955 ;
        RECT 106.175 104.625 106.855 104.955 ;
        RECT 105.710 104.495 105.880 104.625 ;
        RECT 105.485 104.325 105.880 104.495 ;
        RECT 104.855 103.105 105.315 104.155 ;
        RECT 105.485 102.965 105.655 104.325 ;
        RECT 106.050 104.065 106.515 104.455 ;
        RECT 105.825 103.255 106.175 103.875 ;
        RECT 106.345 103.475 106.515 104.065 ;
        RECT 106.685 103.845 106.855 104.625 ;
        RECT 107.025 104.525 107.195 104.865 ;
        RECT 107.430 104.695 107.760 105.125 ;
        RECT 107.930 104.525 108.100 104.865 ;
        RECT 108.395 104.665 108.765 105.125 ;
        RECT 107.025 104.355 108.100 104.525 ;
        RECT 108.935 104.495 109.105 104.955 ;
        RECT 109.340 104.615 110.210 104.955 ;
        RECT 110.380 104.665 110.630 105.125 ;
        RECT 108.545 104.325 109.105 104.495 ;
        RECT 108.545 104.185 108.715 104.325 ;
        RECT 107.215 104.015 108.715 104.185 ;
        RECT 109.410 104.155 109.870 104.445 ;
        RECT 106.685 103.675 108.375 103.845 ;
        RECT 106.345 103.255 106.700 103.475 ;
        RECT 106.870 102.965 107.040 103.675 ;
        RECT 107.245 103.255 108.035 103.505 ;
        RECT 108.205 103.495 108.375 103.675 ;
        RECT 108.545 103.325 108.715 104.015 ;
        RECT 104.985 102.575 105.315 102.935 ;
        RECT 105.485 102.795 105.980 102.965 ;
        RECT 106.185 102.795 107.040 102.965 ;
        RECT 107.915 102.575 108.245 103.035 ;
        RECT 108.455 102.935 108.715 103.325 ;
        RECT 108.905 104.145 109.870 104.155 ;
        RECT 110.040 104.235 110.210 104.615 ;
        RECT 110.800 104.575 110.970 104.865 ;
        RECT 111.150 104.745 111.480 105.125 ;
        RECT 110.800 104.405 111.600 104.575 ;
        RECT 108.905 103.985 109.580 104.145 ;
        RECT 110.040 104.065 111.260 104.235 ;
        RECT 108.905 103.195 109.115 103.985 ;
        RECT 110.040 103.975 110.210 104.065 ;
        RECT 109.285 103.195 109.635 103.815 ;
        RECT 109.805 103.805 110.210 103.975 ;
        RECT 109.805 103.025 109.975 103.805 ;
        RECT 110.145 103.355 110.365 103.635 ;
        RECT 110.545 103.525 111.085 103.895 ;
        RECT 111.430 103.785 111.600 104.405 ;
        RECT 111.775 104.065 111.945 105.125 ;
        RECT 112.155 104.115 112.445 104.955 ;
        RECT 112.615 104.285 112.785 105.125 ;
        RECT 112.995 104.115 113.245 104.955 ;
        RECT 113.455 104.285 113.625 105.125 ;
        RECT 114.415 104.285 114.585 105.125 ;
        RECT 114.795 104.115 115.045 104.955 ;
        RECT 115.255 104.285 115.425 105.125 ;
        RECT 115.595 104.115 115.885 104.955 ;
        RECT 112.155 103.945 113.880 104.115 ;
        RECT 110.145 103.185 110.675 103.355 ;
        RECT 108.455 102.765 108.805 102.935 ;
        RECT 109.025 102.745 109.975 103.025 ;
        RECT 110.145 102.575 110.335 103.015 ;
        RECT 110.505 102.955 110.675 103.185 ;
        RECT 110.845 103.125 111.085 103.525 ;
        RECT 111.255 103.775 111.600 103.785 ;
        RECT 111.255 103.565 113.285 103.775 ;
        RECT 111.255 103.310 111.580 103.565 ;
        RECT 113.470 103.395 113.880 103.945 ;
        RECT 111.255 102.955 111.575 103.310 ;
        RECT 110.505 102.785 111.575 102.955 ;
        RECT 111.775 102.575 111.945 103.385 ;
        RECT 112.115 103.225 113.880 103.395 ;
        RECT 114.160 103.945 115.885 104.115 ;
        RECT 116.095 104.065 116.265 105.125 ;
        RECT 116.560 104.745 116.890 105.125 ;
        RECT 117.070 104.575 117.240 104.865 ;
        RECT 117.410 104.665 117.660 105.125 ;
        RECT 116.440 104.405 117.240 104.575 ;
        RECT 117.830 104.615 118.700 104.955 ;
        RECT 114.160 103.395 114.570 103.945 ;
        RECT 116.440 103.785 116.610 104.405 ;
        RECT 117.830 104.235 118.000 104.615 ;
        RECT 118.935 104.495 119.105 104.955 ;
        RECT 119.275 104.665 119.645 105.125 ;
        RECT 119.940 104.525 120.110 104.865 ;
        RECT 120.280 104.695 120.610 105.125 ;
        RECT 120.845 104.525 121.015 104.865 ;
        RECT 116.780 104.065 118.000 104.235 ;
        RECT 118.170 104.155 118.630 104.445 ;
        RECT 118.935 104.325 119.495 104.495 ;
        RECT 119.940 104.355 121.015 104.525 ;
        RECT 121.185 104.625 121.865 104.955 ;
        RECT 122.080 104.625 122.330 104.955 ;
        RECT 122.500 104.665 122.750 105.125 ;
        RECT 119.325 104.185 119.495 104.325 ;
        RECT 118.170 104.145 119.135 104.155 ;
        RECT 117.830 103.975 118.000 104.065 ;
        RECT 118.460 103.985 119.135 104.145 ;
        RECT 116.440 103.775 116.785 103.785 ;
        RECT 114.755 103.565 116.785 103.775 ;
        RECT 114.160 103.225 115.925 103.395 ;
        RECT 112.115 102.745 112.445 103.225 ;
        RECT 112.615 102.575 112.785 103.045 ;
        RECT 112.955 102.745 113.285 103.225 ;
        RECT 113.455 102.575 113.625 103.045 ;
        RECT 114.415 102.575 114.585 103.045 ;
        RECT 114.755 102.745 115.085 103.225 ;
        RECT 115.255 102.575 115.425 103.045 ;
        RECT 115.595 102.745 115.925 103.225 ;
        RECT 116.095 102.575 116.265 103.385 ;
        RECT 116.460 103.310 116.785 103.565 ;
        RECT 116.465 102.955 116.785 103.310 ;
        RECT 116.955 103.525 117.495 103.895 ;
        RECT 117.830 103.805 118.235 103.975 ;
        RECT 116.955 103.125 117.195 103.525 ;
        RECT 117.675 103.355 117.895 103.635 ;
        RECT 117.365 103.185 117.895 103.355 ;
        RECT 117.365 102.955 117.535 103.185 ;
        RECT 118.065 103.025 118.235 103.805 ;
        RECT 118.405 103.195 118.755 103.815 ;
        RECT 118.925 103.195 119.135 103.985 ;
        RECT 119.325 104.015 120.825 104.185 ;
        RECT 119.325 103.325 119.495 104.015 ;
        RECT 121.185 103.845 121.355 104.625 ;
        RECT 122.160 104.495 122.330 104.625 ;
        RECT 119.665 103.675 121.355 103.845 ;
        RECT 121.525 104.065 121.990 104.455 ;
        RECT 122.160 104.325 122.555 104.495 ;
        RECT 119.665 103.495 119.835 103.675 ;
        RECT 116.465 102.785 117.535 102.955 ;
        RECT 117.705 102.575 117.895 103.015 ;
        RECT 118.065 102.745 119.015 103.025 ;
        RECT 119.325 102.935 119.585 103.325 ;
        RECT 120.005 103.255 120.795 103.505 ;
        RECT 119.235 102.765 119.585 102.935 ;
        RECT 119.795 102.575 120.125 103.035 ;
        RECT 121.000 102.965 121.170 103.675 ;
        RECT 121.525 103.475 121.695 104.065 ;
        RECT 121.340 103.255 121.695 103.475 ;
        RECT 121.865 103.255 122.215 103.875 ;
        RECT 122.385 102.965 122.555 104.325 ;
        RECT 122.920 104.155 123.245 104.940 ;
        RECT 122.725 103.105 123.185 104.155 ;
        RECT 121.000 102.795 121.855 102.965 ;
        RECT 122.060 102.795 122.555 102.965 ;
        RECT 122.725 102.575 123.055 102.935 ;
        RECT 123.415 102.835 123.585 104.955 ;
        RECT 123.755 104.625 124.085 105.125 ;
        RECT 124.255 104.455 124.510 104.955 ;
        RECT 123.760 104.285 124.510 104.455 ;
        RECT 123.760 103.295 123.990 104.285 ;
        RECT 124.160 103.465 124.510 104.115 ;
        RECT 125.145 104.050 125.415 104.955 ;
        RECT 125.585 104.365 125.915 105.125 ;
        RECT 126.095 104.195 126.275 104.955 ;
        RECT 123.760 103.125 124.510 103.295 ;
        RECT 123.755 102.575 124.085 102.955 ;
        RECT 124.255 102.835 124.510 103.125 ;
        RECT 125.145 103.250 125.325 104.050 ;
        RECT 125.600 104.025 126.275 104.195 ;
        RECT 126.525 104.035 127.735 105.125 ;
        RECT 125.600 103.880 125.770 104.025 ;
        RECT 125.495 103.550 125.770 103.880 ;
        RECT 125.600 103.295 125.770 103.550 ;
        RECT 125.995 103.475 126.335 103.845 ;
        RECT 126.525 103.495 127.045 104.035 ;
        RECT 127.215 103.325 127.735 103.865 ;
        RECT 125.145 102.745 125.405 103.250 ;
        RECT 125.600 103.125 126.265 103.295 ;
        RECT 125.585 102.575 125.915 102.955 ;
        RECT 126.095 102.745 126.265 103.125 ;
        RECT 126.525 102.575 127.735 103.325 ;
        RECT 14.660 102.405 127.820 102.575 ;
        RECT 14.745 101.655 15.955 102.405 ;
        RECT 14.745 101.115 15.265 101.655 ;
        RECT 16.125 101.635 18.715 102.405 ;
        RECT 18.890 101.860 24.235 102.405 ;
        RECT 15.435 100.945 15.955 101.485 ;
        RECT 14.745 99.855 15.955 100.945 ;
        RECT 16.125 100.945 17.335 101.465 ;
        RECT 17.505 101.115 18.715 101.635 ;
        RECT 16.125 99.855 18.715 100.945 ;
        RECT 20.480 100.290 20.830 101.540 ;
        RECT 22.310 101.030 22.650 101.860 ;
        RECT 24.405 101.680 24.695 102.405 ;
        RECT 24.865 101.655 26.075 102.405 ;
        RECT 26.250 101.860 31.595 102.405 ;
        RECT 31.770 101.860 37.115 102.405 ;
        RECT 18.890 99.855 24.235 100.290 ;
        RECT 24.405 99.855 24.695 101.020 ;
        RECT 24.865 100.945 25.385 101.485 ;
        RECT 25.555 101.115 26.075 101.655 ;
        RECT 24.865 99.855 26.075 100.945 ;
        RECT 27.840 100.290 28.190 101.540 ;
        RECT 29.670 101.030 30.010 101.860 ;
        RECT 33.360 100.290 33.710 101.540 ;
        RECT 35.190 101.030 35.530 101.860 ;
        RECT 37.285 101.680 37.575 102.405 ;
        RECT 37.745 101.655 38.955 102.405 ;
        RECT 39.130 101.860 44.475 102.405 ;
        RECT 44.650 101.860 49.995 102.405 ;
        RECT 26.250 99.855 31.595 100.290 ;
        RECT 31.770 99.855 37.115 100.290 ;
        RECT 37.285 99.855 37.575 101.020 ;
        RECT 37.745 100.945 38.265 101.485 ;
        RECT 38.435 101.115 38.955 101.655 ;
        RECT 37.745 99.855 38.955 100.945 ;
        RECT 40.720 100.290 41.070 101.540 ;
        RECT 42.550 101.030 42.890 101.860 ;
        RECT 46.240 100.290 46.590 101.540 ;
        RECT 48.070 101.030 48.410 101.860 ;
        RECT 50.165 101.680 50.455 102.405 ;
        RECT 50.630 101.860 55.975 102.405 ;
        RECT 56.150 101.860 61.495 102.405 ;
        RECT 39.130 99.855 44.475 100.290 ;
        RECT 44.650 99.855 49.995 100.290 ;
        RECT 50.165 99.855 50.455 101.020 ;
        RECT 52.220 100.290 52.570 101.540 ;
        RECT 54.050 101.030 54.390 101.860 ;
        RECT 57.740 100.290 58.090 101.540 ;
        RECT 59.570 101.030 59.910 101.860 ;
        RECT 61.705 101.585 61.935 102.405 ;
        RECT 62.105 101.605 62.435 102.235 ;
        RECT 61.685 101.165 62.015 101.415 ;
        RECT 62.185 101.005 62.435 101.605 ;
        RECT 62.605 101.585 62.815 102.405 ;
        RECT 63.045 101.680 63.335 102.405 ;
        RECT 64.465 101.585 64.695 102.405 ;
        RECT 64.865 101.605 65.195 102.235 ;
        RECT 64.445 101.165 64.775 101.415 ;
        RECT 50.630 99.855 55.975 100.290 ;
        RECT 56.150 99.855 61.495 100.290 ;
        RECT 61.705 99.855 61.935 100.995 ;
        RECT 62.105 100.025 62.435 101.005 ;
        RECT 62.605 99.855 62.815 100.995 ;
        RECT 63.045 99.855 63.335 101.020 ;
        RECT 64.945 101.005 65.195 101.605 ;
        RECT 65.365 101.585 65.575 102.405 ;
        RECT 66.725 101.635 70.235 102.405 ;
        RECT 70.410 101.860 75.755 102.405 ;
        RECT 64.465 99.855 64.695 100.995 ;
        RECT 64.865 100.025 65.195 101.005 ;
        RECT 65.365 99.855 65.575 100.995 ;
        RECT 66.725 100.945 68.415 101.465 ;
        RECT 68.585 101.115 70.235 101.635 ;
        RECT 66.725 99.855 70.235 100.945 ;
        RECT 72.000 100.290 72.350 101.540 ;
        RECT 73.830 101.030 74.170 101.860 ;
        RECT 75.925 101.680 76.215 102.405 ;
        RECT 76.385 101.655 77.595 102.405 ;
        RECT 77.770 101.860 83.115 102.405 ;
        RECT 83.290 101.860 88.635 102.405 ;
        RECT 70.410 99.855 75.755 100.290 ;
        RECT 75.925 99.855 76.215 101.020 ;
        RECT 76.385 100.945 76.905 101.485 ;
        RECT 77.075 101.115 77.595 101.655 ;
        RECT 76.385 99.855 77.595 100.945 ;
        RECT 79.360 100.290 79.710 101.540 ;
        RECT 81.190 101.030 81.530 101.860 ;
        RECT 84.880 100.290 85.230 101.540 ;
        RECT 86.710 101.030 87.050 101.860 ;
        RECT 88.805 101.680 89.095 102.405 ;
        RECT 89.265 101.655 90.475 102.405 ;
        RECT 90.650 101.860 95.995 102.405 ;
        RECT 96.170 101.860 101.515 102.405 ;
        RECT 77.770 99.855 83.115 100.290 ;
        RECT 83.290 99.855 88.635 100.290 ;
        RECT 88.805 99.855 89.095 101.020 ;
        RECT 89.265 100.945 89.785 101.485 ;
        RECT 89.955 101.115 90.475 101.655 ;
        RECT 89.265 99.855 90.475 100.945 ;
        RECT 92.240 100.290 92.590 101.540 ;
        RECT 94.070 101.030 94.410 101.860 ;
        RECT 97.760 100.290 98.110 101.540 ;
        RECT 99.590 101.030 99.930 101.860 ;
        RECT 101.685 101.680 101.975 102.405 ;
        RECT 102.145 101.655 103.355 102.405 ;
        RECT 103.530 101.860 108.875 102.405 ;
        RECT 109.050 101.860 114.395 102.405 ;
        RECT 90.650 99.855 95.995 100.290 ;
        RECT 96.170 99.855 101.515 100.290 ;
        RECT 101.685 99.855 101.975 101.020 ;
        RECT 102.145 100.945 102.665 101.485 ;
        RECT 102.835 101.115 103.355 101.655 ;
        RECT 102.145 99.855 103.355 100.945 ;
        RECT 105.120 100.290 105.470 101.540 ;
        RECT 106.950 101.030 107.290 101.860 ;
        RECT 110.640 100.290 110.990 101.540 ;
        RECT 112.470 101.030 112.810 101.860 ;
        RECT 114.565 101.680 114.855 102.405 ;
        RECT 115.485 101.635 118.995 102.405 ;
        RECT 103.530 99.855 108.875 100.290 ;
        RECT 109.050 99.855 114.395 100.290 ;
        RECT 114.565 99.855 114.855 101.020 ;
        RECT 115.485 100.945 117.175 101.465 ;
        RECT 117.345 101.115 118.995 101.635 ;
        RECT 119.205 101.585 119.435 102.405 ;
        RECT 119.605 101.605 119.935 102.235 ;
        RECT 119.185 101.165 119.515 101.415 ;
        RECT 119.685 101.005 119.935 101.605 ;
        RECT 120.105 101.585 120.315 102.405 ;
        RECT 121.010 101.860 126.355 102.405 ;
        RECT 115.485 99.855 118.995 100.945 ;
        RECT 119.205 99.855 119.435 100.995 ;
        RECT 119.605 100.025 119.935 101.005 ;
        RECT 120.105 99.855 120.315 100.995 ;
        RECT 122.600 100.290 122.950 101.540 ;
        RECT 124.430 101.030 124.770 101.860 ;
        RECT 126.525 101.655 127.735 102.405 ;
        RECT 126.525 100.945 127.045 101.485 ;
        RECT 127.215 101.115 127.735 101.655 ;
        RECT 121.010 99.855 126.355 100.290 ;
        RECT 126.525 99.855 127.735 100.945 ;
        RECT 14.660 99.685 127.820 99.855 ;
        RECT 19.165 66.070 30.165 66.940 ;
        RECT 19.165 54.930 20.835 66.070 ;
        RECT 21.465 65.555 26.465 65.725 ;
        RECT 21.235 55.300 21.405 65.340 ;
        RECT 26.525 55.300 26.695 65.340 ;
        RECT 27.095 54.930 27.265 66.070 ;
        RECT 27.895 65.555 28.895 65.725 ;
        RECT 27.665 55.300 27.835 65.340 ;
        RECT 28.955 55.300 29.125 65.340 ;
        RECT 29.525 54.930 30.165 66.070 ;
        RECT 19.165 52.860 30.165 54.930 ;
        RECT 19.165 49.370 21.005 52.860 ;
        RECT 22.765 52.780 30.165 52.860 ;
        RECT 21.635 52.350 22.135 52.520 ;
        RECT 21.405 50.095 21.575 52.135 ;
        RECT 22.195 50.095 22.365 52.135 ;
        RECT 21.635 49.710 22.135 49.880 ;
        RECT 22.765 49.370 25.085 52.780 ;
        RECT 25.715 52.270 26.215 52.440 ;
        RECT 19.165 48.650 25.085 49.370 ;
        RECT 19.135 48.040 23.045 48.260 ;
        RECT 19.135 45.640 20.855 48.040 ;
        RECT 21.485 47.530 21.985 47.700 ;
        RECT 21.255 46.320 21.425 47.360 ;
        RECT 22.045 46.320 22.215 47.360 ;
        RECT 21.485 45.980 21.985 46.150 ;
        RECT 22.615 45.640 23.045 48.040 ;
        RECT 24.025 46.290 25.085 48.650 ;
        RECT 25.485 47.015 25.655 52.055 ;
        RECT 26.275 47.015 26.445 52.055 ;
        RECT 25.715 46.630 26.215 46.800 ;
        RECT 26.845 46.290 27.015 52.780 ;
        RECT 27.645 52.270 28.145 52.440 ;
        RECT 27.415 47.015 27.585 52.055 ;
        RECT 28.205 47.015 28.375 52.055 ;
        RECT 27.645 46.630 28.145 46.800 ;
        RECT 28.775 46.290 30.165 52.780 ;
        RECT 30.365 66.080 41.365 66.950 ;
        RECT 30.365 54.940 32.035 66.080 ;
        RECT 32.665 65.565 37.665 65.735 ;
        RECT 32.435 55.310 32.605 65.350 ;
        RECT 37.725 55.310 37.895 65.350 ;
        RECT 38.295 54.940 38.465 66.080 ;
        RECT 39.095 65.565 40.095 65.735 ;
        RECT 38.865 55.310 39.035 65.350 ;
        RECT 40.155 55.310 40.325 65.350 ;
        RECT 40.725 54.940 41.365 66.080 ;
        RECT 30.365 52.870 41.365 54.940 ;
        RECT 30.365 49.380 32.205 52.870 ;
        RECT 33.965 52.790 41.365 52.870 ;
        RECT 32.835 52.360 33.335 52.530 ;
        RECT 32.605 50.105 32.775 52.145 ;
        RECT 33.395 50.105 33.565 52.145 ;
        RECT 32.835 49.720 33.335 49.890 ;
        RECT 33.965 49.380 36.285 52.790 ;
        RECT 36.915 52.280 37.415 52.450 ;
        RECT 30.365 48.660 36.285 49.380 ;
        RECT 24.025 45.800 30.165 46.290 ;
        RECT 30.335 48.050 34.245 48.270 ;
        RECT 19.135 45.370 23.045 45.640 ;
        RECT 30.335 45.650 32.055 48.050 ;
        RECT 32.685 47.540 33.185 47.710 ;
        RECT 32.455 46.330 32.625 47.370 ;
        RECT 33.245 46.330 33.415 47.370 ;
        RECT 32.685 45.990 33.185 46.160 ;
        RECT 33.815 45.650 34.245 48.050 ;
        RECT 35.225 46.300 36.285 48.660 ;
        RECT 36.685 47.025 36.855 52.065 ;
        RECT 37.475 47.025 37.645 52.065 ;
        RECT 36.915 46.640 37.415 46.810 ;
        RECT 38.045 46.300 38.215 52.790 ;
        RECT 38.845 52.280 39.345 52.450 ;
        RECT 38.615 47.025 38.785 52.065 ;
        RECT 39.405 47.025 39.575 52.065 ;
        RECT 38.845 46.640 39.345 46.810 ;
        RECT 39.975 46.300 41.365 52.790 ;
        RECT 41.585 66.050 52.585 66.920 ;
        RECT 41.585 54.910 43.255 66.050 ;
        RECT 43.885 65.535 48.885 65.705 ;
        RECT 43.655 55.280 43.825 65.320 ;
        RECT 48.945 55.280 49.115 65.320 ;
        RECT 49.515 54.910 49.685 66.050 ;
        RECT 50.315 65.535 51.315 65.705 ;
        RECT 50.085 55.280 50.255 65.320 ;
        RECT 51.375 55.280 51.545 65.320 ;
        RECT 51.945 54.910 52.585 66.050 ;
        RECT 41.585 52.840 52.585 54.910 ;
        RECT 41.585 49.350 43.425 52.840 ;
        RECT 45.185 52.760 52.585 52.840 ;
        RECT 44.055 52.330 44.555 52.500 ;
        RECT 43.825 50.075 43.995 52.115 ;
        RECT 44.615 50.075 44.785 52.115 ;
        RECT 44.055 49.690 44.555 49.860 ;
        RECT 45.185 49.350 47.505 52.760 ;
        RECT 48.135 52.250 48.635 52.420 ;
        RECT 41.585 48.630 47.505 49.350 ;
        RECT 35.225 45.810 41.365 46.300 ;
        RECT 41.555 48.020 45.465 48.240 ;
        RECT 30.335 45.380 34.245 45.650 ;
        RECT 41.555 45.620 43.275 48.020 ;
        RECT 43.905 47.510 44.405 47.680 ;
        RECT 43.675 46.300 43.845 47.340 ;
        RECT 44.465 46.300 44.635 47.340 ;
        RECT 43.905 45.960 44.405 46.130 ;
        RECT 45.035 45.620 45.465 48.020 ;
        RECT 46.445 46.270 47.505 48.630 ;
        RECT 47.905 46.995 48.075 52.035 ;
        RECT 48.695 46.995 48.865 52.035 ;
        RECT 48.135 46.610 48.635 46.780 ;
        RECT 49.265 46.270 49.435 52.760 ;
        RECT 50.065 52.250 50.565 52.420 ;
        RECT 49.835 46.995 50.005 52.035 ;
        RECT 50.625 46.995 50.795 52.035 ;
        RECT 50.065 46.610 50.565 46.780 ;
        RECT 51.195 46.270 52.585 52.760 ;
        RECT 52.835 66.030 63.835 66.900 ;
        RECT 52.835 54.890 54.505 66.030 ;
        RECT 55.135 65.515 60.135 65.685 ;
        RECT 54.905 55.260 55.075 65.300 ;
        RECT 60.195 55.260 60.365 65.300 ;
        RECT 60.765 54.890 60.935 66.030 ;
        RECT 61.565 65.515 62.565 65.685 ;
        RECT 61.335 55.260 61.505 65.300 ;
        RECT 62.625 55.260 62.795 65.300 ;
        RECT 63.195 54.890 63.835 66.030 ;
        RECT 52.835 52.820 63.835 54.890 ;
        RECT 52.835 49.330 54.675 52.820 ;
        RECT 56.435 52.740 63.835 52.820 ;
        RECT 55.305 52.310 55.805 52.480 ;
        RECT 55.075 50.055 55.245 52.095 ;
        RECT 55.865 50.055 56.035 52.095 ;
        RECT 55.305 49.670 55.805 49.840 ;
        RECT 56.435 49.330 58.755 52.740 ;
        RECT 59.385 52.230 59.885 52.400 ;
        RECT 52.835 48.610 58.755 49.330 ;
        RECT 46.445 45.780 52.585 46.270 ;
        RECT 52.805 48.000 56.715 48.220 ;
        RECT 41.555 45.350 45.465 45.620 ;
        RECT 52.805 45.600 54.525 48.000 ;
        RECT 55.155 47.490 55.655 47.660 ;
        RECT 54.925 46.280 55.095 47.320 ;
        RECT 55.715 46.280 55.885 47.320 ;
        RECT 55.155 45.940 55.655 46.110 ;
        RECT 56.285 45.600 56.715 48.000 ;
        RECT 57.695 46.250 58.755 48.610 ;
        RECT 59.155 46.975 59.325 52.015 ;
        RECT 59.945 46.975 60.115 52.015 ;
        RECT 59.385 46.590 59.885 46.760 ;
        RECT 60.515 46.250 60.685 52.740 ;
        RECT 61.315 52.230 61.815 52.400 ;
        RECT 61.085 46.975 61.255 52.015 ;
        RECT 61.875 46.975 62.045 52.015 ;
        RECT 61.315 46.590 61.815 46.760 ;
        RECT 62.445 46.250 63.835 52.740 ;
        RECT 64.055 66.020 75.055 66.890 ;
        RECT 64.055 54.880 65.725 66.020 ;
        RECT 66.355 65.505 71.355 65.675 ;
        RECT 66.125 55.250 66.295 65.290 ;
        RECT 71.415 55.250 71.585 65.290 ;
        RECT 71.985 54.880 72.155 66.020 ;
        RECT 72.785 65.505 73.785 65.675 ;
        RECT 72.555 55.250 72.725 65.290 ;
        RECT 73.845 55.250 74.015 65.290 ;
        RECT 74.415 54.880 75.055 66.020 ;
        RECT 64.055 52.810 75.055 54.880 ;
        RECT 64.055 49.320 65.895 52.810 ;
        RECT 67.655 52.730 75.055 52.810 ;
        RECT 66.525 52.300 67.025 52.470 ;
        RECT 66.295 50.045 66.465 52.085 ;
        RECT 67.085 50.045 67.255 52.085 ;
        RECT 66.525 49.660 67.025 49.830 ;
        RECT 67.655 49.320 69.975 52.730 ;
        RECT 70.605 52.220 71.105 52.390 ;
        RECT 64.055 48.600 69.975 49.320 ;
        RECT 57.695 45.760 63.835 46.250 ;
        RECT 64.025 47.990 67.935 48.210 ;
        RECT 52.805 45.330 56.715 45.600 ;
        RECT 64.025 45.590 65.745 47.990 ;
        RECT 66.375 47.480 66.875 47.650 ;
        RECT 66.145 46.270 66.315 47.310 ;
        RECT 66.935 46.270 67.105 47.310 ;
        RECT 66.375 45.930 66.875 46.100 ;
        RECT 67.505 45.590 67.935 47.990 ;
        RECT 68.915 46.240 69.975 48.600 ;
        RECT 70.375 46.965 70.545 52.005 ;
        RECT 71.165 46.965 71.335 52.005 ;
        RECT 70.605 46.580 71.105 46.750 ;
        RECT 71.735 46.240 71.905 52.730 ;
        RECT 72.535 52.220 73.035 52.390 ;
        RECT 72.305 46.965 72.475 52.005 ;
        RECT 73.095 46.965 73.265 52.005 ;
        RECT 72.535 46.580 73.035 46.750 ;
        RECT 73.665 46.240 75.055 52.730 ;
        RECT 75.295 66.010 86.295 66.880 ;
        RECT 75.295 54.870 76.965 66.010 ;
        RECT 77.595 65.495 82.595 65.665 ;
        RECT 77.365 55.240 77.535 65.280 ;
        RECT 82.655 55.240 82.825 65.280 ;
        RECT 83.225 54.870 83.395 66.010 ;
        RECT 84.025 65.495 85.025 65.665 ;
        RECT 83.795 55.240 83.965 65.280 ;
        RECT 85.085 55.240 85.255 65.280 ;
        RECT 85.655 54.870 86.295 66.010 ;
        RECT 75.295 52.800 86.295 54.870 ;
        RECT 75.295 49.310 77.135 52.800 ;
        RECT 78.895 52.720 86.295 52.800 ;
        RECT 77.765 52.290 78.265 52.460 ;
        RECT 77.535 50.035 77.705 52.075 ;
        RECT 78.325 50.035 78.495 52.075 ;
        RECT 77.765 49.650 78.265 49.820 ;
        RECT 78.895 49.310 81.215 52.720 ;
        RECT 81.845 52.210 82.345 52.380 ;
        RECT 75.295 48.590 81.215 49.310 ;
        RECT 68.915 45.750 75.055 46.240 ;
        RECT 75.265 47.980 79.175 48.200 ;
        RECT 64.025 45.320 67.935 45.590 ;
        RECT 75.265 45.580 76.985 47.980 ;
        RECT 77.615 47.470 78.115 47.640 ;
        RECT 77.385 46.260 77.555 47.300 ;
        RECT 78.175 46.260 78.345 47.300 ;
        RECT 77.615 45.920 78.115 46.090 ;
        RECT 78.745 45.580 79.175 47.980 ;
        RECT 80.155 46.230 81.215 48.590 ;
        RECT 81.615 46.955 81.785 51.995 ;
        RECT 82.405 46.955 82.575 51.995 ;
        RECT 81.845 46.570 82.345 46.740 ;
        RECT 82.975 46.230 83.145 52.720 ;
        RECT 83.775 52.210 84.275 52.380 ;
        RECT 83.545 46.955 83.715 51.995 ;
        RECT 84.335 46.955 84.505 51.995 ;
        RECT 83.775 46.570 84.275 46.740 ;
        RECT 84.905 46.230 86.295 52.720 ;
        RECT 86.545 66.020 97.545 66.890 ;
        RECT 131.125 66.880 140.025 66.890 ;
        RECT 86.545 54.880 88.215 66.020 ;
        RECT 88.845 65.505 93.845 65.675 ;
        RECT 88.615 55.250 88.785 65.290 ;
        RECT 93.905 55.250 94.075 65.290 ;
        RECT 94.475 54.880 94.645 66.020 ;
        RECT 95.275 65.505 96.275 65.675 ;
        RECT 95.045 55.250 95.215 65.290 ;
        RECT 96.335 55.250 96.505 65.290 ;
        RECT 96.905 54.880 97.545 66.020 ;
        RECT 86.545 52.810 97.545 54.880 ;
        RECT 86.545 49.320 88.385 52.810 ;
        RECT 90.145 52.730 97.545 52.810 ;
        RECT 89.015 52.300 89.515 52.470 ;
        RECT 88.785 50.045 88.955 52.085 ;
        RECT 89.575 50.045 89.745 52.085 ;
        RECT 89.015 49.660 89.515 49.830 ;
        RECT 90.145 49.320 92.465 52.730 ;
        RECT 93.095 52.220 93.595 52.390 ;
        RECT 86.545 48.600 92.465 49.320 ;
        RECT 80.155 45.740 86.295 46.230 ;
        RECT 86.515 47.990 90.425 48.210 ;
        RECT 75.265 45.310 79.175 45.580 ;
        RECT 86.515 45.590 88.235 47.990 ;
        RECT 88.865 47.480 89.365 47.650 ;
        RECT 88.635 46.270 88.805 47.310 ;
        RECT 89.425 46.270 89.595 47.310 ;
        RECT 88.865 45.930 89.365 46.100 ;
        RECT 89.995 45.590 90.425 47.990 ;
        RECT 91.405 46.240 92.465 48.600 ;
        RECT 92.865 46.965 93.035 52.005 ;
        RECT 93.655 46.965 93.825 52.005 ;
        RECT 93.095 46.580 93.595 46.750 ;
        RECT 94.225 46.240 94.395 52.730 ;
        RECT 95.025 52.220 95.525 52.390 ;
        RECT 94.795 46.965 94.965 52.005 ;
        RECT 95.585 46.965 95.755 52.005 ;
        RECT 95.025 46.580 95.525 46.750 ;
        RECT 96.155 46.240 97.545 52.730 ;
        RECT 97.825 66.010 108.825 66.880 ;
        RECT 97.825 54.870 99.495 66.010 ;
        RECT 100.125 65.495 105.125 65.665 ;
        RECT 99.895 55.240 100.065 65.280 ;
        RECT 105.185 55.240 105.355 65.280 ;
        RECT 105.755 54.870 105.925 66.010 ;
        RECT 106.555 65.495 107.555 65.665 ;
        RECT 106.325 55.240 106.495 65.280 ;
        RECT 107.615 55.240 107.785 65.280 ;
        RECT 108.185 54.870 108.825 66.010 ;
        RECT 97.825 52.800 108.825 54.870 ;
        RECT 97.825 49.310 99.665 52.800 ;
        RECT 101.425 52.720 108.825 52.800 ;
        RECT 100.295 52.290 100.795 52.460 ;
        RECT 100.065 50.035 100.235 52.075 ;
        RECT 100.855 50.035 101.025 52.075 ;
        RECT 100.295 49.650 100.795 49.820 ;
        RECT 101.425 49.310 103.745 52.720 ;
        RECT 104.375 52.210 104.875 52.380 ;
        RECT 97.825 48.590 103.745 49.310 ;
        RECT 91.405 45.750 97.545 46.240 ;
        RECT 97.795 47.980 101.705 48.200 ;
        RECT 86.515 45.320 90.425 45.590 ;
        RECT 97.795 45.580 99.515 47.980 ;
        RECT 100.145 47.470 100.645 47.640 ;
        RECT 99.915 46.260 100.085 47.300 ;
        RECT 100.705 46.260 100.875 47.300 ;
        RECT 100.145 45.920 100.645 46.090 ;
        RECT 101.275 45.580 101.705 47.980 ;
        RECT 102.685 46.230 103.745 48.590 ;
        RECT 104.145 46.955 104.315 51.995 ;
        RECT 104.935 46.955 105.105 51.995 ;
        RECT 104.375 46.570 104.875 46.740 ;
        RECT 105.505 46.230 105.675 52.720 ;
        RECT 106.305 52.210 106.805 52.380 ;
        RECT 106.075 46.955 106.245 51.995 ;
        RECT 106.865 46.955 107.035 51.995 ;
        RECT 106.305 46.570 106.805 46.740 ;
        RECT 107.435 46.230 108.825 52.720 ;
        RECT 109.095 66.010 120.095 66.880 ;
        RECT 109.095 54.870 110.765 66.010 ;
        RECT 111.395 65.495 116.395 65.665 ;
        RECT 111.165 55.240 111.335 65.280 ;
        RECT 116.455 55.240 116.625 65.280 ;
        RECT 117.025 54.870 117.195 66.010 ;
        RECT 117.825 65.495 118.825 65.665 ;
        RECT 117.595 55.240 117.765 65.280 ;
        RECT 118.885 55.240 119.055 65.280 ;
        RECT 119.455 54.870 120.095 66.010 ;
        RECT 109.095 52.800 120.095 54.870 ;
        RECT 109.095 49.310 110.935 52.800 ;
        RECT 112.695 52.720 120.095 52.800 ;
        RECT 111.565 52.290 112.065 52.460 ;
        RECT 111.335 50.035 111.505 52.075 ;
        RECT 112.125 50.035 112.295 52.075 ;
        RECT 111.565 49.650 112.065 49.820 ;
        RECT 112.695 49.310 115.015 52.720 ;
        RECT 115.645 52.210 116.145 52.380 ;
        RECT 109.095 48.590 115.015 49.310 ;
        RECT 102.685 45.740 108.825 46.230 ;
        RECT 109.065 47.980 112.975 48.200 ;
        RECT 97.795 45.310 101.705 45.580 ;
        RECT 109.065 45.580 110.785 47.980 ;
        RECT 111.415 47.470 111.915 47.640 ;
        RECT 111.185 46.260 111.355 47.300 ;
        RECT 111.975 46.260 112.145 47.300 ;
        RECT 111.415 45.920 111.915 46.090 ;
        RECT 112.545 45.580 112.975 47.980 ;
        RECT 113.955 46.230 115.015 48.590 ;
        RECT 115.415 46.955 115.585 51.995 ;
        RECT 116.205 46.955 116.375 51.995 ;
        RECT 115.645 46.570 116.145 46.740 ;
        RECT 116.775 46.230 116.945 52.720 ;
        RECT 117.575 52.210 118.075 52.380 ;
        RECT 117.345 46.955 117.515 51.995 ;
        RECT 118.135 46.955 118.305 51.995 ;
        RECT 117.575 46.570 118.075 46.740 ;
        RECT 118.705 46.230 120.095 52.720 ;
        RECT 120.345 66.010 140.025 66.880 ;
        RECT 120.345 54.870 122.015 66.010 ;
        RECT 122.645 65.495 127.645 65.665 ;
        RECT 122.415 55.240 122.585 65.280 ;
        RECT 127.705 55.240 127.875 65.280 ;
        RECT 128.275 54.870 128.445 66.010 ;
        RECT 130.705 65.980 140.025 66.010 ;
        RECT 129.075 65.495 130.075 65.665 ;
        RECT 128.845 55.240 129.015 65.280 ;
        RECT 130.135 55.240 130.305 65.280 ;
        RECT 130.705 54.870 132.765 65.980 ;
        RECT 133.395 65.465 138.395 65.635 ;
        RECT 133.165 55.210 133.335 65.250 ;
        RECT 138.455 55.210 138.625 65.250 ;
        RECT 120.345 54.840 132.765 54.870 ;
        RECT 139.025 54.840 140.025 65.980 ;
        RECT 120.345 54.720 140.025 54.840 ;
        RECT 120.345 53.550 140.035 54.720 ;
        RECT 120.345 52.800 131.345 53.550 ;
        RECT 120.345 49.310 122.185 52.800 ;
        RECT 123.945 52.720 131.345 52.800 ;
        RECT 122.815 52.290 123.315 52.460 ;
        RECT 122.585 50.035 122.755 52.075 ;
        RECT 123.375 50.035 123.545 52.075 ;
        RECT 122.815 49.650 123.315 49.820 ;
        RECT 123.945 49.310 126.265 52.720 ;
        RECT 126.895 52.210 127.395 52.380 ;
        RECT 120.345 48.590 126.265 49.310 ;
        RECT 113.955 45.740 120.095 46.230 ;
        RECT 120.315 47.980 124.225 48.200 ;
        RECT 109.065 45.310 112.975 45.580 ;
        RECT 120.315 45.580 122.035 47.980 ;
        RECT 122.665 47.470 123.165 47.640 ;
        RECT 122.435 46.260 122.605 47.300 ;
        RECT 123.225 46.260 123.395 47.300 ;
        RECT 122.665 45.920 123.165 46.090 ;
        RECT 123.795 45.580 124.225 47.980 ;
        RECT 125.205 46.230 126.265 48.590 ;
        RECT 126.665 46.955 126.835 51.995 ;
        RECT 127.455 46.955 127.625 51.995 ;
        RECT 126.895 46.570 127.395 46.740 ;
        RECT 128.025 46.230 128.195 52.720 ;
        RECT 128.825 52.210 129.325 52.380 ;
        RECT 128.595 46.955 128.765 51.995 ;
        RECT 129.385 46.955 129.555 51.995 ;
        RECT 128.825 46.570 129.325 46.740 ;
        RECT 129.955 46.230 131.345 52.720 ;
        RECT 125.205 45.740 131.345 46.230 ;
        RECT 120.315 45.310 124.225 45.580 ;
        RECT 25.695 39.770 29.605 40.040 ;
        RECT 18.575 39.120 24.715 39.610 ;
        RECT 18.575 32.630 19.965 39.120 ;
        RECT 20.595 38.610 21.095 38.780 ;
        RECT 20.365 33.355 20.535 38.395 ;
        RECT 21.155 33.355 21.325 38.395 ;
        RECT 20.595 32.970 21.095 33.140 ;
        RECT 21.725 32.630 21.895 39.120 ;
        RECT 22.525 38.610 23.025 38.780 ;
        RECT 22.295 33.355 22.465 38.395 ;
        RECT 23.085 33.355 23.255 38.395 ;
        RECT 23.655 36.760 24.715 39.120 ;
        RECT 25.695 37.370 26.125 39.770 ;
        RECT 26.755 39.260 27.255 39.430 ;
        RECT 26.525 38.050 26.695 39.090 ;
        RECT 27.315 38.050 27.485 39.090 ;
        RECT 26.755 37.710 27.255 37.880 ;
        RECT 27.885 37.370 29.605 39.770 ;
        RECT 36.975 39.770 40.885 40.040 ;
        RECT 25.695 37.150 29.605 37.370 ;
        RECT 29.855 39.120 35.995 39.610 ;
        RECT 23.655 36.040 29.575 36.760 ;
        RECT 22.525 32.970 23.025 33.140 ;
        RECT 23.655 32.630 25.975 36.040 ;
        RECT 26.605 35.530 27.105 35.700 ;
        RECT 26.375 33.275 26.545 35.315 ;
        RECT 27.165 33.275 27.335 35.315 ;
        RECT 26.605 32.890 27.105 33.060 ;
        RECT 18.575 32.550 25.975 32.630 ;
        RECT 27.735 32.550 29.575 36.040 ;
        RECT 18.575 30.480 29.575 32.550 ;
        RECT 18.575 19.340 19.215 30.480 ;
        RECT 19.615 20.070 19.785 30.110 ;
        RECT 20.905 20.070 21.075 30.110 ;
        RECT 19.845 19.685 20.845 19.855 ;
        RECT 21.475 19.340 21.645 30.480 ;
        RECT 22.045 20.070 22.215 30.110 ;
        RECT 27.335 20.070 27.505 30.110 ;
        RECT 22.275 19.685 27.275 19.855 ;
        RECT 27.905 19.340 29.575 30.480 ;
        RECT 18.575 18.470 29.575 19.340 ;
        RECT 29.855 32.630 31.245 39.120 ;
        RECT 31.875 38.610 32.375 38.780 ;
        RECT 31.645 33.355 31.815 38.395 ;
        RECT 32.435 33.355 32.605 38.395 ;
        RECT 31.875 32.970 32.375 33.140 ;
        RECT 33.005 32.630 33.175 39.120 ;
        RECT 33.805 38.610 34.305 38.780 ;
        RECT 33.575 33.355 33.745 38.395 ;
        RECT 34.365 33.355 34.535 38.395 ;
        RECT 34.935 36.760 35.995 39.120 ;
        RECT 36.975 37.370 37.405 39.770 ;
        RECT 38.035 39.260 38.535 39.430 ;
        RECT 37.805 38.050 37.975 39.090 ;
        RECT 38.595 38.050 38.765 39.090 ;
        RECT 38.035 37.710 38.535 37.880 ;
        RECT 39.165 37.370 40.885 39.770 ;
        RECT 48.265 39.750 52.175 40.020 ;
        RECT 36.975 37.150 40.885 37.370 ;
        RECT 41.145 39.100 47.285 39.590 ;
        RECT 34.935 36.040 40.855 36.760 ;
        RECT 33.805 32.970 34.305 33.140 ;
        RECT 34.935 32.630 37.255 36.040 ;
        RECT 37.885 35.530 38.385 35.700 ;
        RECT 37.655 33.275 37.825 35.315 ;
        RECT 38.445 33.275 38.615 35.315 ;
        RECT 37.885 32.890 38.385 33.060 ;
        RECT 29.855 32.550 37.255 32.630 ;
        RECT 39.015 32.550 40.855 36.040 ;
        RECT 29.855 30.480 40.855 32.550 ;
        RECT 29.855 19.340 30.495 30.480 ;
        RECT 30.895 20.070 31.065 30.110 ;
        RECT 32.185 20.070 32.355 30.110 ;
        RECT 31.125 19.685 32.125 19.855 ;
        RECT 32.755 19.340 32.925 30.480 ;
        RECT 33.325 20.070 33.495 30.110 ;
        RECT 38.615 20.070 38.785 30.110 ;
        RECT 33.555 19.685 38.555 19.855 ;
        RECT 39.185 19.340 40.855 30.480 ;
        RECT 29.855 18.470 40.855 19.340 ;
        RECT 41.145 32.610 42.535 39.100 ;
        RECT 43.165 38.590 43.665 38.760 ;
        RECT 42.935 33.335 43.105 38.375 ;
        RECT 43.725 33.335 43.895 38.375 ;
        RECT 43.165 32.950 43.665 33.120 ;
        RECT 44.295 32.610 44.465 39.100 ;
        RECT 45.095 38.590 45.595 38.760 ;
        RECT 44.865 33.335 45.035 38.375 ;
        RECT 45.655 33.335 45.825 38.375 ;
        RECT 46.225 36.740 47.285 39.100 ;
        RECT 48.265 37.350 48.695 39.750 ;
        RECT 49.325 39.240 49.825 39.410 ;
        RECT 49.095 38.030 49.265 39.070 ;
        RECT 49.885 38.030 50.055 39.070 ;
        RECT 49.325 37.690 49.825 37.860 ;
        RECT 50.455 37.350 52.175 39.750 ;
        RECT 59.485 39.750 63.395 40.020 ;
        RECT 48.265 37.130 52.175 37.350 ;
        RECT 52.365 39.100 58.505 39.590 ;
        RECT 46.225 36.020 52.145 36.740 ;
        RECT 45.095 32.950 45.595 33.120 ;
        RECT 46.225 32.610 48.545 36.020 ;
        RECT 49.175 35.510 49.675 35.680 ;
        RECT 48.945 33.255 49.115 35.295 ;
        RECT 49.735 33.255 49.905 35.295 ;
        RECT 49.175 32.870 49.675 33.040 ;
        RECT 41.145 32.530 48.545 32.610 ;
        RECT 50.305 32.530 52.145 36.020 ;
        RECT 41.145 30.460 52.145 32.530 ;
        RECT 41.145 19.320 41.785 30.460 ;
        RECT 42.185 20.050 42.355 30.090 ;
        RECT 43.475 20.050 43.645 30.090 ;
        RECT 42.415 19.665 43.415 19.835 ;
        RECT 44.045 19.320 44.215 30.460 ;
        RECT 44.615 20.050 44.785 30.090 ;
        RECT 49.905 20.050 50.075 30.090 ;
        RECT 44.845 19.665 49.845 19.835 ;
        RECT 50.475 19.320 52.145 30.460 ;
        RECT 41.145 18.450 52.145 19.320 ;
        RECT 52.365 32.610 53.755 39.100 ;
        RECT 54.385 38.590 54.885 38.760 ;
        RECT 54.155 33.335 54.325 38.375 ;
        RECT 54.945 33.335 55.115 38.375 ;
        RECT 54.385 32.950 54.885 33.120 ;
        RECT 55.515 32.610 55.685 39.100 ;
        RECT 56.315 38.590 56.815 38.760 ;
        RECT 56.085 33.335 56.255 38.375 ;
        RECT 56.875 33.335 57.045 38.375 ;
        RECT 57.445 36.740 58.505 39.100 ;
        RECT 59.485 37.350 59.915 39.750 ;
        RECT 60.545 39.240 61.045 39.410 ;
        RECT 60.315 38.030 60.485 39.070 ;
        RECT 61.105 38.030 61.275 39.070 ;
        RECT 60.545 37.690 61.045 37.860 ;
        RECT 61.675 37.350 63.395 39.750 ;
        RECT 70.685 39.750 74.595 40.020 ;
        RECT 59.485 37.130 63.395 37.350 ;
        RECT 63.565 39.100 69.705 39.590 ;
        RECT 57.445 36.020 63.365 36.740 ;
        RECT 56.315 32.950 56.815 33.120 ;
        RECT 57.445 32.610 59.765 36.020 ;
        RECT 60.395 35.510 60.895 35.680 ;
        RECT 60.165 33.255 60.335 35.295 ;
        RECT 60.955 33.255 61.125 35.295 ;
        RECT 60.395 32.870 60.895 33.040 ;
        RECT 52.365 32.530 59.765 32.610 ;
        RECT 61.525 32.530 63.365 36.020 ;
        RECT 52.365 30.460 63.365 32.530 ;
        RECT 52.365 19.320 53.005 30.460 ;
        RECT 53.405 20.050 53.575 30.090 ;
        RECT 54.695 20.050 54.865 30.090 ;
        RECT 53.635 19.665 54.635 19.835 ;
        RECT 55.265 19.320 55.435 30.460 ;
        RECT 55.835 20.050 56.005 30.090 ;
        RECT 61.125 20.050 61.295 30.090 ;
        RECT 56.065 19.665 61.065 19.835 ;
        RECT 61.695 19.320 63.365 30.460 ;
        RECT 52.365 18.450 63.365 19.320 ;
        RECT 63.565 32.610 64.955 39.100 ;
        RECT 65.585 38.590 66.085 38.760 ;
        RECT 65.355 33.335 65.525 38.375 ;
        RECT 66.145 33.335 66.315 38.375 ;
        RECT 65.585 32.950 66.085 33.120 ;
        RECT 66.715 32.610 66.885 39.100 ;
        RECT 67.515 38.590 68.015 38.760 ;
        RECT 67.285 33.335 67.455 38.375 ;
        RECT 68.075 33.335 68.245 38.375 ;
        RECT 68.645 36.740 69.705 39.100 ;
        RECT 70.685 37.350 71.115 39.750 ;
        RECT 71.745 39.240 72.245 39.410 ;
        RECT 71.515 38.030 71.685 39.070 ;
        RECT 72.305 38.030 72.475 39.070 ;
        RECT 71.745 37.690 72.245 37.860 ;
        RECT 72.875 37.350 74.595 39.750 ;
        RECT 81.975 39.740 85.885 40.010 ;
        RECT 70.685 37.130 74.595 37.350 ;
        RECT 74.855 39.090 80.995 39.580 ;
        RECT 68.645 36.020 74.565 36.740 ;
        RECT 67.515 32.950 68.015 33.120 ;
        RECT 68.645 32.610 70.965 36.020 ;
        RECT 71.595 35.510 72.095 35.680 ;
        RECT 71.365 33.255 71.535 35.295 ;
        RECT 72.155 33.255 72.325 35.295 ;
        RECT 71.595 32.870 72.095 33.040 ;
        RECT 63.565 32.530 70.965 32.610 ;
        RECT 72.725 32.530 74.565 36.020 ;
        RECT 63.565 30.460 74.565 32.530 ;
        RECT 63.565 19.320 64.205 30.460 ;
        RECT 64.605 20.050 64.775 30.090 ;
        RECT 65.895 20.050 66.065 30.090 ;
        RECT 64.835 19.665 65.835 19.835 ;
        RECT 66.465 19.320 66.635 30.460 ;
        RECT 67.035 20.050 67.205 30.090 ;
        RECT 72.325 20.050 72.495 30.090 ;
        RECT 67.265 19.665 72.265 19.835 ;
        RECT 72.895 19.320 74.565 30.460 ;
        RECT 63.565 18.450 74.565 19.320 ;
        RECT 74.855 32.600 76.245 39.090 ;
        RECT 76.875 38.580 77.375 38.750 ;
        RECT 76.645 33.325 76.815 38.365 ;
        RECT 77.435 33.325 77.605 38.365 ;
        RECT 76.875 32.940 77.375 33.110 ;
        RECT 78.005 32.600 78.175 39.090 ;
        RECT 78.805 38.580 79.305 38.750 ;
        RECT 78.575 33.325 78.745 38.365 ;
        RECT 79.365 33.325 79.535 38.365 ;
        RECT 79.935 36.730 80.995 39.090 ;
        RECT 81.975 37.340 82.405 39.740 ;
        RECT 83.035 39.230 83.535 39.400 ;
        RECT 82.805 38.020 82.975 39.060 ;
        RECT 83.595 38.020 83.765 39.060 ;
        RECT 83.035 37.680 83.535 37.850 ;
        RECT 84.165 37.340 85.885 39.740 ;
        RECT 93.215 39.760 97.125 40.030 ;
        RECT 81.975 37.120 85.885 37.340 ;
        RECT 86.095 39.110 92.235 39.600 ;
        RECT 79.935 36.010 85.855 36.730 ;
        RECT 78.805 32.940 79.305 33.110 ;
        RECT 79.935 32.600 82.255 36.010 ;
        RECT 82.885 35.500 83.385 35.670 ;
        RECT 82.655 33.245 82.825 35.285 ;
        RECT 83.445 33.245 83.615 35.285 ;
        RECT 82.885 32.860 83.385 33.030 ;
        RECT 74.855 32.520 82.255 32.600 ;
        RECT 84.015 32.520 85.855 36.010 ;
        RECT 74.855 30.450 85.855 32.520 ;
        RECT 74.855 19.310 75.495 30.450 ;
        RECT 75.895 20.040 76.065 30.080 ;
        RECT 77.185 20.040 77.355 30.080 ;
        RECT 76.125 19.655 77.125 19.825 ;
        RECT 77.755 19.310 77.925 30.450 ;
        RECT 78.325 20.040 78.495 30.080 ;
        RECT 83.615 20.040 83.785 30.080 ;
        RECT 78.555 19.655 83.555 19.825 ;
        RECT 84.185 19.310 85.855 30.450 ;
        RECT 74.855 18.440 85.855 19.310 ;
        RECT 86.095 32.620 87.485 39.110 ;
        RECT 88.115 38.600 88.615 38.770 ;
        RECT 87.885 33.345 88.055 38.385 ;
        RECT 88.675 33.345 88.845 38.385 ;
        RECT 88.115 32.960 88.615 33.130 ;
        RECT 89.245 32.620 89.415 39.110 ;
        RECT 90.045 38.600 90.545 38.770 ;
        RECT 89.815 33.345 89.985 38.385 ;
        RECT 90.605 33.345 90.775 38.385 ;
        RECT 91.175 36.750 92.235 39.110 ;
        RECT 93.215 37.360 93.645 39.760 ;
        RECT 94.275 39.250 94.775 39.420 ;
        RECT 94.045 38.040 94.215 39.080 ;
        RECT 94.835 38.040 95.005 39.080 ;
        RECT 94.275 37.700 94.775 37.870 ;
        RECT 95.405 37.360 97.125 39.760 ;
        RECT 104.425 39.780 108.335 40.050 ;
        RECT 93.215 37.140 97.125 37.360 ;
        RECT 97.305 39.130 103.445 39.620 ;
        RECT 91.175 36.030 97.095 36.750 ;
        RECT 90.045 32.960 90.545 33.130 ;
        RECT 91.175 32.620 93.495 36.030 ;
        RECT 94.125 35.520 94.625 35.690 ;
        RECT 93.895 33.265 94.065 35.305 ;
        RECT 94.685 33.265 94.855 35.305 ;
        RECT 94.125 32.880 94.625 33.050 ;
        RECT 86.095 32.540 93.495 32.620 ;
        RECT 95.255 32.540 97.095 36.030 ;
        RECT 86.095 30.470 97.095 32.540 ;
        RECT 86.095 19.330 86.735 30.470 ;
        RECT 87.135 20.060 87.305 30.100 ;
        RECT 88.425 20.060 88.595 30.100 ;
        RECT 87.365 19.675 88.365 19.845 ;
        RECT 88.995 19.330 89.165 30.470 ;
        RECT 89.565 20.060 89.735 30.100 ;
        RECT 94.855 20.060 95.025 30.100 ;
        RECT 89.795 19.675 94.795 19.845 ;
        RECT 95.425 19.330 97.095 30.470 ;
        RECT 86.095 18.460 97.095 19.330 ;
        RECT 97.305 32.640 98.695 39.130 ;
        RECT 99.325 38.620 99.825 38.790 ;
        RECT 99.095 33.365 99.265 38.405 ;
        RECT 99.885 33.365 100.055 38.405 ;
        RECT 99.325 32.980 99.825 33.150 ;
        RECT 100.455 32.640 100.625 39.130 ;
        RECT 101.255 38.620 101.755 38.790 ;
        RECT 101.025 33.365 101.195 38.405 ;
        RECT 101.815 33.365 101.985 38.405 ;
        RECT 102.385 36.770 103.445 39.130 ;
        RECT 104.425 37.380 104.855 39.780 ;
        RECT 105.485 39.270 105.985 39.440 ;
        RECT 105.255 38.060 105.425 39.100 ;
        RECT 106.045 38.060 106.215 39.100 ;
        RECT 105.485 37.720 105.985 37.890 ;
        RECT 106.615 37.380 108.335 39.780 ;
        RECT 115.625 39.820 119.535 40.090 ;
        RECT 104.425 37.160 108.335 37.380 ;
        RECT 108.505 39.170 114.645 39.660 ;
        RECT 102.385 36.050 108.305 36.770 ;
        RECT 101.255 32.980 101.755 33.150 ;
        RECT 102.385 32.640 104.705 36.050 ;
        RECT 105.335 35.540 105.835 35.710 ;
        RECT 105.105 33.285 105.275 35.325 ;
        RECT 105.895 33.285 106.065 35.325 ;
        RECT 105.335 32.900 105.835 33.070 ;
        RECT 97.305 32.560 104.705 32.640 ;
        RECT 106.465 32.560 108.305 36.050 ;
        RECT 97.305 30.490 108.305 32.560 ;
        RECT 97.305 19.350 97.945 30.490 ;
        RECT 98.345 20.080 98.515 30.120 ;
        RECT 99.635 20.080 99.805 30.120 ;
        RECT 98.575 19.695 99.575 19.865 ;
        RECT 100.205 19.350 100.375 30.490 ;
        RECT 100.775 20.080 100.945 30.120 ;
        RECT 106.065 20.080 106.235 30.120 ;
        RECT 101.005 19.695 106.005 19.865 ;
        RECT 106.635 19.350 108.305 30.490 ;
        RECT 97.305 18.480 108.305 19.350 ;
        RECT 108.505 32.680 109.895 39.170 ;
        RECT 110.525 38.660 111.025 38.830 ;
        RECT 110.295 33.405 110.465 38.445 ;
        RECT 111.085 33.405 111.255 38.445 ;
        RECT 110.525 33.020 111.025 33.190 ;
        RECT 111.655 32.680 111.825 39.170 ;
        RECT 112.455 38.660 112.955 38.830 ;
        RECT 112.225 33.405 112.395 38.445 ;
        RECT 113.015 33.405 113.185 38.445 ;
        RECT 113.585 36.810 114.645 39.170 ;
        RECT 115.625 37.420 116.055 39.820 ;
        RECT 116.685 39.310 117.185 39.480 ;
        RECT 116.455 38.100 116.625 39.140 ;
        RECT 117.245 38.100 117.415 39.140 ;
        RECT 116.685 37.760 117.185 37.930 ;
        RECT 117.815 37.420 119.535 39.820 ;
        RECT 126.835 39.840 130.745 40.110 ;
        RECT 115.625 37.200 119.535 37.420 ;
        RECT 119.715 39.190 125.855 39.680 ;
        RECT 113.585 36.090 119.505 36.810 ;
        RECT 112.455 33.020 112.955 33.190 ;
        RECT 113.585 32.680 115.905 36.090 ;
        RECT 116.535 35.580 117.035 35.750 ;
        RECT 116.305 33.325 116.475 35.365 ;
        RECT 117.095 33.325 117.265 35.365 ;
        RECT 116.535 32.940 117.035 33.110 ;
        RECT 108.505 32.600 115.905 32.680 ;
        RECT 117.665 32.600 119.505 36.090 ;
        RECT 108.505 30.530 119.505 32.600 ;
        RECT 108.505 19.390 109.145 30.530 ;
        RECT 109.545 20.120 109.715 30.160 ;
        RECT 110.835 20.120 111.005 30.160 ;
        RECT 109.775 19.735 110.775 19.905 ;
        RECT 111.405 19.390 111.575 30.530 ;
        RECT 111.975 20.120 112.145 30.160 ;
        RECT 117.265 20.120 117.435 30.160 ;
        RECT 112.205 19.735 117.205 19.905 ;
        RECT 117.835 19.390 119.505 30.530 ;
        RECT 108.505 18.520 119.505 19.390 ;
        RECT 119.715 32.700 121.105 39.190 ;
        RECT 121.735 38.680 122.235 38.850 ;
        RECT 121.505 33.425 121.675 38.465 ;
        RECT 122.295 33.425 122.465 38.465 ;
        RECT 121.735 33.040 122.235 33.210 ;
        RECT 122.865 32.700 123.035 39.190 ;
        RECT 123.665 38.680 124.165 38.850 ;
        RECT 123.435 33.425 123.605 38.465 ;
        RECT 124.225 33.425 124.395 38.465 ;
        RECT 124.795 36.830 125.855 39.190 ;
        RECT 126.835 37.440 127.265 39.840 ;
        RECT 127.895 39.330 128.395 39.500 ;
        RECT 127.665 38.120 127.835 39.160 ;
        RECT 128.455 38.120 128.625 39.160 ;
        RECT 127.895 37.780 128.395 37.950 ;
        RECT 129.025 37.440 130.745 39.840 ;
        RECT 126.835 37.220 130.745 37.440 ;
        RECT 124.795 36.110 130.715 36.830 ;
        RECT 123.665 33.040 124.165 33.210 ;
        RECT 124.795 32.700 127.115 36.110 ;
        RECT 127.745 35.600 128.245 35.770 ;
        RECT 127.515 33.345 127.685 35.385 ;
        RECT 128.305 33.345 128.475 35.385 ;
        RECT 127.745 32.960 128.245 33.130 ;
        RECT 119.715 32.620 127.115 32.700 ;
        RECT 128.875 32.620 130.715 36.110 ;
        RECT 119.715 31.140 130.715 32.620 ;
        RECT 119.715 30.550 139.465 31.140 ;
        RECT 119.715 19.410 120.355 30.550 ;
        RECT 120.755 20.140 120.925 30.180 ;
        RECT 122.045 20.140 122.215 30.180 ;
        RECT 120.985 19.755 121.985 19.925 ;
        RECT 122.615 19.410 122.785 30.550 ;
        RECT 129.045 30.520 139.465 30.550 ;
        RECT 123.185 20.140 123.355 30.180 ;
        RECT 128.475 20.140 128.645 30.180 ;
        RECT 123.415 19.755 128.415 19.925 ;
        RECT 129.045 19.410 132.075 30.520 ;
        RECT 132.475 20.110 132.645 30.150 ;
        RECT 137.765 20.110 137.935 30.150 ;
        RECT 132.705 19.725 137.705 19.895 ;
        RECT 119.715 19.380 132.075 19.410 ;
        RECT 138.335 19.380 139.465 30.520 ;
        RECT 119.715 18.540 139.465 19.380 ;
        RECT 131.925 18.520 139.465 18.540 ;
      LAYER met1 ;
        RECT 135.340 223.880 136.790 225.180 ;
        RECT 14.660 211.050 127.820 211.530 ;
        RECT 14.660 208.330 127.820 208.810 ;
        RECT 14.660 205.610 127.820 206.090 ;
        RECT 64.885 205.070 65.175 205.115 ;
        RECT 67.285 205.070 67.575 205.115 ;
        RECT 70.525 205.070 71.175 205.115 ;
        RECT 64.885 204.930 71.175 205.070 ;
        RECT 64.885 204.885 65.175 204.930 ;
        RECT 67.285 204.885 67.875 204.930 ;
        RECT 70.525 204.885 71.175 204.930 ;
        RECT 62.585 204.730 62.875 204.775 ;
        RECT 63.950 204.730 64.270 204.790 ;
        RECT 64.425 204.730 64.715 204.775 ;
        RECT 62.585 204.590 64.715 204.730 ;
        RECT 62.585 204.545 62.875 204.590 ;
        RECT 63.950 204.530 64.270 204.590 ;
        RECT 64.425 204.545 64.715 204.590 ;
        RECT 67.585 204.570 67.875 204.885 ;
        RECT 68.665 204.730 68.955 204.775 ;
        RECT 72.245 204.730 72.535 204.775 ;
        RECT 74.080 204.730 74.370 204.775 ;
        RECT 68.665 204.590 74.370 204.730 ;
        RECT 68.665 204.545 68.955 204.590 ;
        RECT 72.245 204.545 72.535 204.590 ;
        RECT 74.080 204.545 74.370 204.590 ;
        RECT 73.150 204.190 73.470 204.450 ;
        RECT 74.530 204.190 74.850 204.450 ;
        RECT 68.665 204.050 68.955 204.095 ;
        RECT 71.785 204.050 72.075 204.095 ;
        RECT 73.675 204.050 73.965 204.095 ;
        RECT 68.665 203.910 73.965 204.050 ;
        RECT 68.665 203.865 68.955 203.910 ;
        RECT 71.785 203.865 72.075 203.910 ;
        RECT 73.675 203.865 73.965 203.910 ;
        RECT 61.190 203.710 61.510 203.770 ;
        RECT 62.125 203.710 62.415 203.755 ;
        RECT 61.190 203.570 62.415 203.710 ;
        RECT 61.190 203.510 61.510 203.570 ;
        RECT 62.125 203.525 62.415 203.570 ;
        RECT 65.805 203.710 66.095 203.755 ;
        RECT 67.170 203.710 67.490 203.770 ;
        RECT 65.805 203.570 67.490 203.710 ;
        RECT 65.805 203.525 66.095 203.570 ;
        RECT 67.170 203.510 67.490 203.570 ;
        RECT 14.660 202.890 127.820 203.370 ;
        RECT 73.150 202.490 73.470 202.750 ;
        RECT 62.685 202.350 62.975 202.395 ;
        RECT 65.805 202.350 66.095 202.395 ;
        RECT 67.695 202.350 67.985 202.395 ;
        RECT 62.685 202.210 67.985 202.350 ;
        RECT 62.685 202.165 62.975 202.210 ;
        RECT 65.805 202.165 66.095 202.210 ;
        RECT 67.695 202.165 67.985 202.210 ;
        RECT 106.845 202.350 107.135 202.395 ;
        RECT 109.965 202.350 110.255 202.395 ;
        RECT 111.855 202.350 112.145 202.395 ;
        RECT 106.845 202.210 112.145 202.350 ;
        RECT 106.845 202.165 107.135 202.210 ;
        RECT 109.965 202.165 110.255 202.210 ;
        RECT 111.855 202.165 112.145 202.210 ;
        RECT 61.190 201.810 61.510 202.070 ;
        RECT 103.050 202.010 103.370 202.070 ;
        RECT 103.985 202.010 104.275 202.055 ;
        RECT 103.050 201.870 104.275 202.010 ;
        RECT 103.050 201.810 103.370 201.870 ;
        RECT 103.985 201.825 104.275 201.870 ;
        RECT 61.280 201.670 61.420 201.810 ;
        RECT 61.605 201.670 61.895 201.690 ;
        RECT 61.280 201.530 61.895 201.670 ;
        RECT 61.605 201.375 61.895 201.530 ;
        RECT 62.685 201.670 62.975 201.715 ;
        RECT 66.265 201.670 66.555 201.715 ;
        RECT 68.100 201.670 68.390 201.715 ;
        RECT 62.685 201.530 68.390 201.670 ;
        RECT 62.685 201.485 62.975 201.530 ;
        RECT 66.265 201.485 66.555 201.530 ;
        RECT 68.100 201.485 68.390 201.530 ;
        RECT 68.550 201.470 68.870 201.730 ;
        RECT 69.930 201.670 70.250 201.730 ;
        RECT 72.245 201.670 72.535 201.715 ;
        RECT 69.930 201.530 72.535 201.670 ;
        RECT 69.930 201.470 70.250 201.530 ;
        RECT 72.245 201.485 72.535 201.530 ;
        RECT 74.070 201.670 74.390 201.730 ;
        RECT 74.545 201.670 74.835 201.715 ;
        RECT 74.070 201.530 74.835 201.670 ;
        RECT 74.070 201.470 74.390 201.530 ;
        RECT 74.545 201.485 74.835 201.530 ;
        RECT 75.005 201.670 75.295 201.715 ;
        RECT 75.910 201.670 76.230 201.730 ;
        RECT 75.005 201.530 76.230 201.670 ;
        RECT 75.005 201.485 75.295 201.530 ;
        RECT 75.910 201.470 76.230 201.530 ;
        RECT 99.370 201.670 99.690 201.730 ;
        RECT 100.305 201.670 100.595 201.715 ;
        RECT 99.370 201.530 100.595 201.670 ;
        RECT 99.370 201.470 99.690 201.530 ;
        RECT 100.305 201.485 100.595 201.530 ;
        RECT 100.750 201.470 101.070 201.730 ;
        RECT 58.445 201.145 58.735 201.375 ;
        RECT 61.305 201.330 61.895 201.375 ;
        RECT 64.545 201.330 65.195 201.375 ;
        RECT 61.305 201.190 65.195 201.330 ;
        RECT 61.305 201.145 61.595 201.190 ;
        RECT 64.545 201.145 65.195 201.190 ;
        RECT 67.185 201.330 67.475 201.375 ;
        RECT 67.630 201.330 67.950 201.390 ;
        RECT 105.765 201.375 106.055 201.690 ;
        RECT 106.845 201.670 107.135 201.715 ;
        RECT 110.425 201.670 110.715 201.715 ;
        RECT 112.260 201.670 112.550 201.715 ;
        RECT 106.845 201.530 112.550 201.670 ;
        RECT 106.845 201.485 107.135 201.530 ;
        RECT 110.425 201.485 110.715 201.530 ;
        RECT 112.260 201.485 112.550 201.530 ;
        RECT 112.710 201.470 113.030 201.730 ;
        RECT 109.030 201.375 109.350 201.390 ;
        RECT 67.185 201.190 67.950 201.330 ;
        RECT 67.185 201.145 67.475 201.190 ;
        RECT 58.520 200.990 58.660 201.145 ;
        RECT 67.630 201.130 67.950 201.190 ;
        RECT 105.465 201.330 106.055 201.375 ;
        RECT 108.705 201.330 109.355 201.375 ;
        RECT 105.465 201.190 109.355 201.330 ;
        RECT 105.465 201.145 105.755 201.190 ;
        RECT 108.705 201.145 109.355 201.190 ;
        RECT 109.030 201.130 109.350 201.145 ;
        RECT 111.330 201.130 111.650 201.390 ;
        RECT 69.470 200.990 69.790 201.050 ;
        RECT 58.520 200.850 69.790 200.990 ;
        RECT 69.470 200.790 69.790 200.850 ;
        RECT 14.660 200.170 127.820 200.650 ;
        RECT 67.630 199.770 67.950 200.030 ;
        RECT 69.930 199.770 70.250 200.030 ;
        RECT 74.990 199.970 75.310 200.030 ;
        RECT 99.370 199.970 99.690 200.030 ;
        RECT 109.030 199.970 109.350 200.030 ;
        RECT 109.505 199.970 109.795 200.015 ;
        RECT 74.990 199.830 105.580 199.970 ;
        RECT 74.990 199.770 75.310 199.830 ;
        RECT 70.390 199.675 70.710 199.690 ;
        RECT 70.390 199.445 70.995 199.675 ;
        RECT 71.785 199.630 72.075 199.675 ;
        RECT 73.150 199.630 73.470 199.690 ;
        RECT 71.785 199.490 73.470 199.630 ;
        RECT 71.785 199.445 72.075 199.490 ;
        RECT 70.390 199.430 70.710 199.445 ;
        RECT 73.150 199.430 73.470 199.490 ;
        RECT 73.725 199.630 74.015 199.675 ;
        RECT 75.910 199.630 76.230 199.690 ;
        RECT 76.965 199.630 77.615 199.675 ;
        RECT 73.725 199.490 77.615 199.630 ;
        RECT 73.725 199.445 74.315 199.490 ;
        RECT 66.710 199.090 67.030 199.350 ;
        RECT 74.025 199.130 74.315 199.445 ;
        RECT 75.910 199.430 76.230 199.490 ;
        RECT 76.965 199.445 77.615 199.490 ;
        RECT 79.590 199.430 79.910 199.690 ;
        RECT 75.105 199.290 75.395 199.335 ;
        RECT 78.685 199.290 78.975 199.335 ;
        RECT 80.520 199.290 80.810 199.335 ;
        RECT 75.105 199.150 80.810 199.290 ;
        RECT 87.040 199.290 87.180 199.830 ;
        RECT 99.370 199.770 99.690 199.830 ;
        RECT 87.885 199.630 88.175 199.675 ;
        RECT 90.745 199.630 91.035 199.675 ;
        RECT 93.985 199.630 94.635 199.675 ;
        RECT 87.885 199.490 94.635 199.630 ;
        RECT 87.885 199.445 88.175 199.490 ;
        RECT 90.745 199.445 91.335 199.490 ;
        RECT 93.985 199.445 94.635 199.490 ;
        RECT 87.425 199.290 87.715 199.335 ;
        RECT 87.040 199.150 87.715 199.290 ;
        RECT 75.105 199.105 75.395 199.150 ;
        RECT 78.685 199.105 78.975 199.150 ;
        RECT 80.520 199.105 80.810 199.150 ;
        RECT 87.425 199.105 87.715 199.150 ;
        RECT 91.045 199.130 91.335 199.445 ;
        RECT 96.610 199.430 96.930 199.690 ;
        RECT 99.945 199.630 100.235 199.675 ;
        RECT 100.750 199.630 101.070 199.690 ;
        RECT 103.185 199.630 103.835 199.675 ;
        RECT 99.945 199.490 103.835 199.630 ;
        RECT 105.440 199.630 105.580 199.830 ;
        RECT 109.030 199.830 109.795 199.970 ;
        RECT 109.030 199.770 109.350 199.830 ;
        RECT 109.505 199.785 109.795 199.830 ;
        RECT 105.440 199.490 109.260 199.630 ;
        RECT 99.945 199.445 100.535 199.490 ;
        RECT 92.125 199.290 92.415 199.335 ;
        RECT 95.705 199.290 95.995 199.335 ;
        RECT 97.540 199.290 97.830 199.335 ;
        RECT 92.125 199.150 97.830 199.290 ;
        RECT 92.125 199.105 92.415 199.150 ;
        RECT 95.705 199.105 95.995 199.150 ;
        RECT 97.540 199.105 97.830 199.150 ;
        RECT 100.245 199.130 100.535 199.445 ;
        RECT 100.750 199.430 101.070 199.490 ;
        RECT 103.185 199.445 103.835 199.490 ;
        RECT 101.325 199.290 101.615 199.335 ;
        RECT 104.905 199.290 105.195 199.335 ;
        RECT 106.740 199.290 107.030 199.335 ;
        RECT 101.325 199.150 107.030 199.290 ;
        RECT 101.325 199.105 101.615 199.150 ;
        RECT 104.905 199.105 105.195 199.150 ;
        RECT 106.740 199.105 107.030 199.150 ;
        RECT 108.570 199.090 108.890 199.350 ;
        RECT 109.120 199.335 109.260 199.490 ;
        RECT 109.045 199.105 109.335 199.335 ;
        RECT 69.930 198.950 70.250 199.010 ;
        RECT 72.245 198.950 72.535 198.995 ;
        RECT 69.930 198.810 72.535 198.950 ;
        RECT 69.930 198.750 70.250 198.810 ;
        RECT 72.245 198.765 72.535 198.810 ;
        RECT 74.530 198.950 74.850 199.010 ;
        RECT 75.910 198.950 76.230 199.010 ;
        RECT 80.985 198.950 81.275 198.995 ;
        RECT 98.005 198.950 98.295 198.995 ;
        RECT 74.530 198.810 98.295 198.950 ;
        RECT 74.530 198.750 74.850 198.810 ;
        RECT 75.910 198.750 76.230 198.810 ;
        RECT 80.985 198.765 81.275 198.810 ;
        RECT 98.005 198.765 98.295 198.810 ;
        RECT 105.825 198.950 106.115 198.995 ;
        RECT 107.205 198.950 107.495 198.995 ;
        RECT 112.250 198.950 112.570 199.010 ;
        RECT 105.825 198.810 106.960 198.950 ;
        RECT 105.825 198.765 106.115 198.810 ;
        RECT 75.105 198.610 75.395 198.655 ;
        RECT 78.225 198.610 78.515 198.655 ;
        RECT 80.115 198.610 80.405 198.655 ;
        RECT 75.105 198.470 80.405 198.610 ;
        RECT 75.105 198.425 75.395 198.470 ;
        RECT 78.225 198.425 78.515 198.470 ;
        RECT 80.115 198.425 80.405 198.470 ;
        RECT 92.125 198.610 92.415 198.655 ;
        RECT 95.245 198.610 95.535 198.655 ;
        RECT 97.135 198.610 97.425 198.655 ;
        RECT 92.125 198.470 97.425 198.610 ;
        RECT 92.125 198.425 92.415 198.470 ;
        RECT 95.245 198.425 95.535 198.470 ;
        RECT 97.135 198.425 97.425 198.470 ;
        RECT 101.325 198.610 101.615 198.655 ;
        RECT 104.445 198.610 104.735 198.655 ;
        RECT 106.335 198.610 106.625 198.655 ;
        RECT 101.325 198.470 106.625 198.610 ;
        RECT 106.820 198.610 106.960 198.810 ;
        RECT 107.205 198.810 112.570 198.950 ;
        RECT 107.205 198.765 107.495 198.810 ;
        RECT 112.250 198.750 112.570 198.810 ;
        RECT 107.665 198.610 107.955 198.655 ;
        RECT 106.820 198.470 107.955 198.610 ;
        RECT 101.325 198.425 101.615 198.470 ;
        RECT 104.445 198.425 104.735 198.470 ;
        RECT 106.335 198.425 106.625 198.470 ;
        RECT 107.665 198.425 107.955 198.470 ;
        RECT 70.865 198.270 71.155 198.315 ;
        RECT 73.610 198.270 73.930 198.330 ;
        RECT 70.865 198.130 73.930 198.270 ;
        RECT 70.865 198.085 71.155 198.130 ;
        RECT 73.610 198.070 73.930 198.130 ;
        RECT 89.265 198.270 89.555 198.315 ;
        RECT 91.090 198.270 91.410 198.330 ;
        RECT 89.265 198.130 91.410 198.270 ;
        RECT 89.265 198.085 89.555 198.130 ;
        RECT 91.090 198.070 91.410 198.130 ;
        RECT 98.465 198.270 98.755 198.315 ;
        RECT 98.910 198.270 99.230 198.330 ;
        RECT 98.465 198.130 99.230 198.270 ;
        RECT 98.465 198.085 98.755 198.130 ;
        RECT 98.910 198.070 99.230 198.130 ;
        RECT 14.660 197.450 127.820 197.930 ;
        RECT 65.790 197.050 66.110 197.310 ;
        RECT 66.710 197.050 67.030 197.310 ;
        RECT 70.850 197.250 71.170 197.310 ;
        RECT 72.705 197.250 72.995 197.295 ;
        RECT 79.145 197.250 79.435 197.295 ;
        RECT 79.590 197.250 79.910 197.310 ;
        RECT 68.180 197.110 77.980 197.250 ;
        RECT 68.180 196.615 68.320 197.110 ;
        RECT 70.850 197.050 71.170 197.110 ;
        RECT 72.705 197.065 72.995 197.110 ;
        RECT 69.010 196.910 69.330 196.970 ;
        RECT 68.640 196.770 69.330 196.910 ;
        RECT 68.640 196.615 68.780 196.770 ;
        RECT 69.010 196.710 69.330 196.770 ;
        RECT 68.105 196.385 68.395 196.615 ;
        RECT 68.565 196.385 68.855 196.615 ;
        RECT 69.470 196.570 69.790 196.630 ;
        RECT 72.230 196.570 72.550 196.630 ;
        RECT 69.470 196.430 73.380 196.570 ;
        RECT 69.470 196.370 69.790 196.430 ;
        RECT 72.230 196.370 72.550 196.430 ;
        RECT 62.585 196.230 62.875 196.275 ;
        RECT 63.950 196.230 64.270 196.290 ;
        RECT 62.585 196.090 64.270 196.230 ;
        RECT 62.585 196.045 62.875 196.090 ;
        RECT 63.950 196.030 64.270 196.090 ;
        RECT 69.030 196.200 69.320 196.275 ;
        RECT 69.030 196.060 69.700 196.200 ;
        RECT 69.030 196.045 69.320 196.060 ;
        RECT 64.885 195.890 65.175 195.935 ;
        RECT 69.560 195.890 69.700 196.060 ;
        RECT 71.770 196.030 72.090 196.290 ;
        RECT 73.240 196.275 73.380 196.430 ;
        RECT 73.610 196.370 73.930 196.630 ;
        RECT 74.990 196.570 75.310 196.630 ;
        RECT 77.305 196.570 77.595 196.615 ;
        RECT 74.990 196.430 77.595 196.570 ;
        RECT 74.990 196.370 75.310 196.430 ;
        RECT 77.305 196.385 77.595 196.430 ;
        RECT 77.840 196.275 77.980 197.110 ;
        RECT 79.145 197.110 79.910 197.250 ;
        RECT 79.145 197.065 79.435 197.110 ;
        RECT 79.590 197.050 79.910 197.110 ;
        RECT 95.245 197.250 95.535 197.295 ;
        RECT 96.610 197.250 96.930 197.310 ;
        RECT 95.245 197.110 96.930 197.250 ;
        RECT 95.245 197.065 95.535 197.110 ;
        RECT 96.610 197.050 96.930 197.110 ;
        RECT 101.225 197.250 101.515 197.295 ;
        RECT 108.570 197.250 108.890 197.310 ;
        RECT 101.225 197.110 108.890 197.250 ;
        RECT 101.225 197.065 101.515 197.110 ;
        RECT 108.570 197.050 108.890 197.110 ;
        RECT 110.425 197.250 110.715 197.295 ;
        RECT 111.330 197.250 111.650 197.310 ;
        RECT 110.425 197.110 111.650 197.250 ;
        RECT 110.425 197.065 110.715 197.110 ;
        RECT 111.330 197.050 111.650 197.110 ;
        RECT 91.180 196.770 98.680 196.910 ;
        RECT 91.180 196.615 91.320 196.770 ;
        RECT 91.105 196.385 91.395 196.615 ;
        RECT 91.550 196.570 91.870 196.630 ;
        RECT 98.540 196.615 98.680 196.770 ;
        RECT 108.125 196.725 108.415 196.955 ;
        RECT 98.465 196.570 98.755 196.615 ;
        RECT 105.350 196.570 105.670 196.630 ;
        RECT 91.550 196.430 96.840 196.570 ;
        RECT 91.550 196.370 91.870 196.430 ;
        RECT 73.165 196.045 73.455 196.275 ;
        RECT 74.545 196.230 74.835 196.275 ;
        RECT 73.700 196.090 74.835 196.230 ;
        RECT 73.700 195.950 73.840 196.090 ;
        RECT 74.545 196.045 74.835 196.090 ;
        RECT 77.765 196.045 78.055 196.275 ;
        RECT 94.325 196.230 94.615 196.275 ;
        RECT 93.940 196.090 94.615 196.230 ;
        RECT 96.700 196.230 96.840 196.430 ;
        RECT 98.465 196.430 105.670 196.570 ;
        RECT 98.465 196.385 98.755 196.430 ;
        RECT 105.350 196.370 105.670 196.430 ;
        RECT 99.385 196.230 99.675 196.275 ;
        RECT 105.810 196.230 106.130 196.290 ;
        RECT 96.700 196.090 106.130 196.230 ;
        RECT 108.200 196.230 108.340 196.725 ;
        RECT 109.505 196.230 109.795 196.275 ;
        RECT 108.200 196.090 109.795 196.230 ;
        RECT 73.610 195.890 73.930 195.950 ;
        RECT 75.465 195.890 75.755 195.935 ;
        RECT 64.885 195.750 68.320 195.890 ;
        RECT 69.560 195.750 73.930 195.890 ;
        RECT 64.885 195.705 65.175 195.750 ;
        RECT 61.650 195.550 61.970 195.610 ;
        RECT 62.125 195.550 62.415 195.595 ;
        RECT 61.650 195.410 62.415 195.550 ;
        RECT 61.650 195.350 61.970 195.410 ;
        RECT 62.125 195.365 62.415 195.410 ;
        RECT 65.935 195.550 66.225 195.595 ;
        RECT 67.185 195.550 67.475 195.595 ;
        RECT 65.935 195.410 67.475 195.550 ;
        RECT 68.180 195.550 68.320 195.750 ;
        RECT 73.610 195.690 73.930 195.750 ;
        RECT 74.620 195.750 75.755 195.890 ;
        RECT 74.620 195.610 74.760 195.750 ;
        RECT 75.465 195.705 75.755 195.750 ;
        RECT 70.390 195.550 70.710 195.610 ;
        RECT 68.180 195.410 70.710 195.550 ;
        RECT 65.935 195.365 66.225 195.410 ;
        RECT 67.185 195.365 67.475 195.410 ;
        RECT 70.390 195.350 70.710 195.410 ;
        RECT 74.530 195.350 74.850 195.610 ;
        RECT 86.030 195.550 86.350 195.610 ;
        RECT 93.940 195.595 94.080 196.090 ;
        RECT 94.325 196.045 94.615 196.090 ;
        RECT 99.385 196.045 99.675 196.090 ;
        RECT 105.810 196.030 106.130 196.090 ;
        RECT 109.505 196.045 109.795 196.090 ;
        RECT 98.910 195.890 99.230 195.950 ;
        RECT 104.890 195.890 105.210 195.950 ;
        RECT 106.285 195.890 106.575 195.935 ;
        RECT 98.910 195.750 106.575 195.890 ;
        RECT 98.910 195.690 99.230 195.750 ;
        RECT 104.890 195.690 105.210 195.750 ;
        RECT 106.285 195.705 106.575 195.750 ;
        RECT 92.025 195.550 92.315 195.595 ;
        RECT 86.030 195.410 92.315 195.550 ;
        RECT 86.030 195.350 86.350 195.410 ;
        RECT 92.025 195.365 92.315 195.410 ;
        RECT 93.865 195.365 94.155 195.595 ;
        RECT 105.810 195.350 106.130 195.610 ;
        RECT 14.660 194.730 127.820 195.210 ;
        RECT 71.770 194.330 72.090 194.590 ;
        RECT 73.150 194.530 73.470 194.590 ;
        RECT 74.990 194.530 75.310 194.590 ;
        RECT 73.150 194.390 75.310 194.530 ;
        RECT 73.150 194.330 73.470 194.390 ;
        RECT 74.990 194.330 75.310 194.390 ;
        RECT 88.345 194.345 88.635 194.575 ;
        RECT 108.585 194.345 108.875 194.575 ;
        RECT 55.210 194.190 55.530 194.250 ;
        RECT 52.080 194.050 55.530 194.190 ;
        RECT 52.080 193.895 52.220 194.050 ;
        RECT 55.210 193.990 55.530 194.050 ;
        RECT 57.045 194.190 57.695 194.235 ;
        RECT 60.645 194.190 60.935 194.235 ;
        RECT 61.650 194.190 61.970 194.250 ;
        RECT 57.045 194.050 61.970 194.190 ;
        RECT 57.045 194.005 57.695 194.050 ;
        RECT 60.345 194.005 60.935 194.050 ;
        RECT 49.705 193.850 49.995 193.895 ;
        RECT 52.005 193.850 52.295 193.895 ;
        RECT 49.705 193.710 52.295 193.850 ;
        RECT 49.705 193.665 49.995 193.710 ;
        RECT 52.005 193.665 52.295 193.710 ;
        RECT 53.850 193.850 54.140 193.895 ;
        RECT 55.685 193.850 55.975 193.895 ;
        RECT 59.265 193.850 59.555 193.895 ;
        RECT 53.850 193.710 59.555 193.850 ;
        RECT 53.850 193.665 54.140 193.710 ;
        RECT 55.685 193.665 55.975 193.710 ;
        RECT 59.265 193.665 59.555 193.710 ;
        RECT 60.345 193.690 60.635 194.005 ;
        RECT 61.650 193.990 61.970 194.050 ;
        RECT 67.645 193.665 67.935 193.895 ;
        RECT 69.010 193.850 69.330 193.910 ;
        RECT 74.530 193.850 74.850 193.910 ;
        RECT 69.010 193.710 74.850 193.850 ;
        RECT 53.385 193.510 53.675 193.555 ;
        RECT 56.590 193.510 56.910 193.570 ;
        RECT 53.385 193.370 56.910 193.510 ;
        RECT 53.385 193.325 53.675 193.370 ;
        RECT 56.590 193.310 56.910 193.370 ;
        RECT 65.790 193.510 66.110 193.570 ;
        RECT 67.185 193.510 67.475 193.555 ;
        RECT 65.790 193.370 67.475 193.510 ;
        RECT 65.790 193.310 66.110 193.370 ;
        RECT 67.185 193.325 67.475 193.370 ;
        RECT 54.255 193.170 54.545 193.215 ;
        RECT 56.145 193.170 56.435 193.215 ;
        RECT 59.265 193.170 59.555 193.215 ;
        RECT 54.255 193.030 59.555 193.170 ;
        RECT 54.255 192.985 54.545 193.030 ;
        RECT 56.145 192.985 56.435 193.030 ;
        RECT 59.265 192.985 59.555 193.030 ;
        RECT 62.125 193.170 62.415 193.215 ;
        RECT 67.720 193.170 67.860 193.665 ;
        RECT 69.010 193.650 69.330 193.710 ;
        RECT 74.530 193.650 74.850 193.710 ;
        RECT 75.465 193.665 75.755 193.895 ;
        RECT 84.190 193.850 84.510 193.910 ;
        RECT 86.505 193.850 86.795 193.895 ;
        RECT 84.190 193.710 86.795 193.850 ;
        RECT 88.420 193.850 88.560 194.345 ;
        RECT 103.050 194.190 103.370 194.250 ;
        RECT 105.810 194.190 106.130 194.250 ;
        RECT 106.745 194.190 107.035 194.235 ;
        RECT 103.050 194.050 107.035 194.190 ;
        RECT 103.050 193.990 103.370 194.050 ;
        RECT 105.810 193.990 106.130 194.050 ;
        RECT 106.745 194.005 107.035 194.050 ;
        RECT 89.725 193.850 90.015 193.895 ;
        RECT 88.420 193.710 90.015 193.850 ;
        RECT 70.390 193.510 70.710 193.570 ;
        RECT 73.610 193.510 73.930 193.570 ;
        RECT 75.540 193.510 75.680 193.665 ;
        RECT 84.190 193.650 84.510 193.710 ;
        RECT 86.505 193.665 86.795 193.710 ;
        RECT 89.725 193.665 90.015 193.710 ;
        RECT 99.370 193.850 99.690 193.910 ;
        RECT 102.590 193.850 102.910 193.910 ;
        RECT 103.525 193.850 103.815 193.895 ;
        RECT 99.370 193.710 103.815 193.850 ;
        RECT 108.660 193.850 108.800 194.345 ;
        RECT 109.045 193.850 109.335 193.895 ;
        RECT 108.660 193.710 109.335 193.850 ;
        RECT 99.370 193.650 99.690 193.710 ;
        RECT 102.590 193.650 102.910 193.710 ;
        RECT 103.525 193.665 103.815 193.710 ;
        RECT 109.045 193.665 109.335 193.710 ;
        RECT 70.390 193.370 75.680 193.510 ;
        RECT 70.390 193.310 70.710 193.370 ;
        RECT 73.610 193.310 73.930 193.370 ;
        RECT 85.110 193.310 85.430 193.570 ;
        RECT 86.030 193.310 86.350 193.570 ;
        RECT 105.350 193.510 105.670 193.570 ;
        RECT 105.825 193.510 106.115 193.555 ;
        RECT 105.350 193.370 106.115 193.510 ;
        RECT 105.350 193.310 105.670 193.370 ;
        RECT 105.825 193.325 106.115 193.370 ;
        RECT 106.285 193.325 106.575 193.555 ;
        RECT 103.510 193.170 103.830 193.230 ;
        RECT 106.360 193.170 106.500 193.325 ;
        RECT 62.125 193.030 69.700 193.170 ;
        RECT 62.125 192.985 62.415 193.030 ;
        RECT 69.560 192.890 69.700 193.030 ;
        RECT 103.510 193.030 106.500 193.170 ;
        RECT 103.510 192.970 103.830 193.030 ;
        RECT 46.010 192.830 46.330 192.890 ;
        RECT 49.245 192.830 49.535 192.875 ;
        RECT 46.010 192.690 49.535 192.830 ;
        RECT 46.010 192.630 46.330 192.690 ;
        RECT 49.245 192.645 49.535 192.690 ;
        RECT 52.465 192.830 52.755 192.875 ;
        RECT 52.910 192.830 53.230 192.890 ;
        RECT 52.465 192.690 53.230 192.830 ;
        RECT 52.465 192.645 52.755 192.690 ;
        RECT 52.910 192.630 53.230 192.690 ;
        RECT 54.705 192.830 54.995 192.875 ;
        RECT 66.265 192.830 66.555 192.875 ;
        RECT 54.705 192.690 66.555 192.830 ;
        RECT 54.705 192.645 54.995 192.690 ;
        RECT 66.265 192.645 66.555 192.690 ;
        RECT 69.470 192.630 69.790 192.890 ;
        RECT 90.630 192.630 90.950 192.890 ;
        RECT 103.970 192.630 104.290 192.890 ;
        RECT 109.965 192.830 110.255 192.875 ;
        RECT 110.870 192.830 111.190 192.890 ;
        RECT 109.965 192.690 111.190 192.830 ;
        RECT 109.965 192.645 110.255 192.690 ;
        RECT 110.870 192.630 111.190 192.690 ;
        RECT 14.660 192.010 127.820 192.490 ;
        RECT 65.790 191.810 66.110 191.870 ;
        RECT 69.485 191.810 69.775 191.855 ;
        RECT 65.790 191.670 69.775 191.810 ;
        RECT 65.790 191.610 66.110 191.670 ;
        RECT 69.485 191.625 69.775 191.670 ;
        RECT 44.600 191.470 44.890 191.515 ;
        RECT 47.380 191.470 47.670 191.515 ;
        RECT 49.240 191.470 49.530 191.515 ;
        RECT 44.600 191.330 49.530 191.470 ;
        RECT 44.600 191.285 44.890 191.330 ;
        RECT 47.380 191.285 47.670 191.330 ;
        RECT 49.240 191.285 49.530 191.330 ;
        RECT 54.720 191.470 55.010 191.515 ;
        RECT 57.500 191.470 57.790 191.515 ;
        RECT 59.360 191.470 59.650 191.515 ;
        RECT 54.720 191.330 59.650 191.470 ;
        RECT 54.720 191.285 55.010 191.330 ;
        RECT 57.500 191.285 57.790 191.330 ;
        RECT 59.360 191.285 59.650 191.330 ;
        RECT 88.300 191.470 88.590 191.515 ;
        RECT 91.080 191.470 91.370 191.515 ;
        RECT 92.940 191.470 93.230 191.515 ;
        RECT 88.300 191.330 93.230 191.470 ;
        RECT 88.300 191.285 88.590 191.330 ;
        RECT 91.080 191.285 91.370 191.330 ;
        RECT 92.940 191.285 93.230 191.330 ;
        RECT 106.385 191.470 106.675 191.515 ;
        RECT 109.505 191.470 109.795 191.515 ;
        RECT 111.395 191.470 111.685 191.515 ;
        RECT 106.385 191.330 111.685 191.470 ;
        RECT 106.385 191.285 106.675 191.330 ;
        RECT 109.505 191.285 109.795 191.330 ;
        RECT 111.395 191.285 111.685 191.330 ;
        RECT 40.735 191.130 41.025 191.175 ;
        RECT 42.790 191.130 43.110 191.190 ;
        RECT 40.735 190.990 43.110 191.130 ;
        RECT 40.735 190.945 41.025 190.990 ;
        RECT 42.790 190.930 43.110 190.990 ;
        RECT 49.705 191.130 49.995 191.175 ;
        RECT 56.590 191.130 56.910 191.190 ;
        RECT 49.705 190.990 57.740 191.130 ;
        RECT 49.705 190.945 49.995 190.990 ;
        RECT 56.590 190.930 56.910 190.990 ;
        RECT 44.600 190.790 44.890 190.835 ;
        RECT 47.865 190.790 48.155 190.835 ;
        RECT 49.230 190.790 49.550 190.850 ;
        RECT 44.600 190.650 47.135 190.790 ;
        RECT 44.600 190.605 44.890 190.650 ;
        RECT 46.010 190.495 46.330 190.510 ;
        RECT 42.740 190.450 43.030 190.495 ;
        RECT 46.000 190.450 46.330 190.495 ;
        RECT 42.740 190.310 46.330 190.450 ;
        RECT 42.740 190.265 43.030 190.310 ;
        RECT 46.000 190.265 46.330 190.310 ;
        RECT 46.920 190.495 47.135 190.650 ;
        RECT 47.865 190.650 49.550 190.790 ;
        RECT 47.865 190.605 48.155 190.650 ;
        RECT 49.230 190.590 49.550 190.650 ;
        RECT 54.720 190.790 55.010 190.835 ;
        RECT 57.600 190.790 57.740 190.990 ;
        RECT 57.970 190.930 58.290 191.190 ;
        RECT 82.810 191.130 83.130 191.190 ;
        RECT 84.435 191.130 84.725 191.175 ;
        RECT 86.030 191.130 86.350 191.190 ;
        RECT 82.810 190.990 86.350 191.130 ;
        RECT 82.810 190.930 83.130 190.990 ;
        RECT 84.435 190.945 84.725 190.990 ;
        RECT 86.030 190.930 86.350 190.990 ;
        RECT 90.630 191.130 90.950 191.190 ;
        RECT 91.565 191.130 91.855 191.175 ;
        RECT 90.630 190.990 91.855 191.130 ;
        RECT 90.630 190.930 90.950 190.990 ;
        RECT 91.565 190.945 91.855 190.990 ;
        RECT 110.870 190.930 111.190 191.190 ;
        RECT 59.825 190.790 60.115 190.835 ;
        RECT 68.550 190.790 68.870 190.850 ;
        RECT 54.720 190.650 57.255 190.790 ;
        RECT 57.600 190.650 68.870 190.790 ;
        RECT 54.720 190.605 55.010 190.650 ;
        RECT 52.910 190.495 53.230 190.510 ;
        RECT 57.040 190.495 57.255 190.650 ;
        RECT 59.825 190.605 60.115 190.650 ;
        RECT 68.550 190.590 68.870 190.650 ;
        RECT 69.025 190.790 69.315 190.835 ;
        RECT 70.390 190.790 70.710 190.850 ;
        RECT 69.025 190.650 70.710 190.790 ;
        RECT 69.025 190.605 69.315 190.650 ;
        RECT 70.390 190.590 70.710 190.650 ;
        RECT 70.865 190.790 71.155 190.835 ;
        RECT 72.230 190.790 72.550 190.850 ;
        RECT 70.865 190.650 72.550 190.790 ;
        RECT 70.865 190.605 71.155 190.650 ;
        RECT 46.920 190.450 47.210 190.495 ;
        RECT 48.780 190.450 49.070 190.495 ;
        RECT 46.920 190.310 49.070 190.450 ;
        RECT 46.920 190.265 47.210 190.310 ;
        RECT 48.780 190.265 49.070 190.310 ;
        RECT 52.860 190.450 53.230 190.495 ;
        RECT 56.120 190.450 56.410 190.495 ;
        RECT 52.860 190.310 56.410 190.450 ;
        RECT 52.860 190.265 53.230 190.310 ;
        RECT 56.120 190.265 56.410 190.310 ;
        RECT 57.040 190.450 57.330 190.495 ;
        RECT 58.900 190.450 59.190 190.495 ;
        RECT 57.040 190.310 59.190 190.450 ;
        RECT 57.040 190.265 57.330 190.310 ;
        RECT 58.900 190.265 59.190 190.310 ;
        RECT 64.870 190.450 65.190 190.510 ;
        RECT 70.940 190.450 71.080 190.605 ;
        RECT 72.230 190.590 72.550 190.650 ;
        RECT 81.445 190.790 81.735 190.835 ;
        RECT 83.270 190.790 83.590 190.850 ;
        RECT 83.745 190.790 84.035 190.835 ;
        RECT 81.445 190.650 84.035 190.790 ;
        RECT 81.445 190.605 81.735 190.650 ;
        RECT 83.270 190.590 83.590 190.650 ;
        RECT 83.745 190.605 84.035 190.650 ;
        RECT 88.300 190.790 88.590 190.835 ;
        RECT 88.300 190.650 90.835 190.790 ;
        RECT 88.300 190.605 88.590 190.650 ;
        RECT 90.620 190.495 90.835 190.650 ;
        RECT 93.390 190.590 93.710 190.850 ;
        RECT 64.870 190.310 71.080 190.450 ;
        RECT 81.905 190.450 82.195 190.495 ;
        RECT 86.440 190.450 86.730 190.495 ;
        RECT 89.700 190.450 89.990 190.495 ;
        RECT 81.905 190.310 89.990 190.450 ;
        RECT 46.010 190.250 46.330 190.265 ;
        RECT 52.910 190.250 53.230 190.265 ;
        RECT 64.870 190.250 65.190 190.310 ;
        RECT 81.905 190.265 82.195 190.310 ;
        RECT 86.440 190.265 86.730 190.310 ;
        RECT 89.700 190.265 89.990 190.310 ;
        RECT 90.620 190.450 90.910 190.495 ;
        RECT 92.480 190.450 92.770 190.495 ;
        RECT 90.620 190.310 92.770 190.450 ;
        RECT 90.620 190.265 90.910 190.310 ;
        RECT 92.480 190.265 92.770 190.310 ;
        RECT 103.970 190.450 104.290 190.510 ;
        RECT 105.305 190.495 105.595 190.810 ;
        RECT 106.385 190.790 106.675 190.835 ;
        RECT 109.965 190.790 110.255 190.835 ;
        RECT 111.800 190.790 112.090 190.835 ;
        RECT 106.385 190.650 112.090 190.790 ;
        RECT 106.385 190.605 106.675 190.650 ;
        RECT 109.965 190.605 110.255 190.650 ;
        RECT 111.800 190.605 112.090 190.650 ;
        RECT 112.250 190.590 112.570 190.850 ;
        RECT 113.630 190.790 113.950 190.850 ;
        RECT 118.705 190.790 118.995 190.835 ;
        RECT 113.630 190.650 118.995 190.790 ;
        RECT 113.630 190.590 113.950 190.650 ;
        RECT 118.705 190.605 118.995 190.650 ;
        RECT 105.005 190.450 105.595 190.495 ;
        RECT 108.245 190.450 108.895 190.495 ;
        RECT 103.970 190.310 108.895 190.450 ;
        RECT 103.970 190.250 104.290 190.310 ;
        RECT 105.005 190.265 105.295 190.310 ;
        RECT 108.245 190.265 108.895 190.310 ;
        RECT 51.070 190.155 51.390 190.170 ;
        RECT 50.855 189.925 51.390 190.155 ;
        RECT 51.070 189.910 51.390 189.925 ;
        RECT 69.010 190.110 69.330 190.170 ;
        RECT 69.945 190.110 70.235 190.155 ;
        RECT 69.010 189.970 70.235 190.110 ;
        RECT 69.010 189.910 69.330 189.970 ;
        RECT 69.945 189.925 70.235 189.970 ;
        RECT 70.405 190.110 70.695 190.155 ;
        RECT 70.850 190.110 71.170 190.170 ;
        RECT 70.405 189.970 71.170 190.110 ;
        RECT 70.405 189.925 70.695 189.970 ;
        RECT 70.850 189.910 71.170 189.970 ;
        RECT 83.285 190.110 83.575 190.155 ;
        RECT 83.730 190.110 84.050 190.170 ;
        RECT 83.285 189.970 84.050 190.110 ;
        RECT 83.285 189.925 83.575 189.970 ;
        RECT 83.730 189.910 84.050 189.970 ;
        RECT 103.510 189.910 103.830 190.170 ;
        RECT 118.245 190.110 118.535 190.155 ;
        RECT 118.690 190.110 119.010 190.170 ;
        RECT 118.245 189.970 119.010 190.110 ;
        RECT 118.245 189.925 118.535 189.970 ;
        RECT 118.690 189.910 119.010 189.970 ;
        RECT 14.660 189.290 127.820 189.770 ;
        RECT 54.765 188.905 55.055 189.135 ;
        RECT 54.840 188.750 54.980 188.905 ;
        RECT 57.970 188.890 58.290 189.150 ;
        RECT 63.950 189.090 64.270 189.150 ;
        RECT 74.070 189.090 74.390 189.150 ;
        RECT 76.370 189.090 76.690 189.150 ;
        RECT 63.950 188.950 76.690 189.090 ;
        RECT 63.950 188.890 64.270 188.950 ;
        RECT 54.840 188.610 57.280 188.750 ;
        RECT 42.790 188.410 43.110 188.470 ;
        RECT 48.325 188.410 48.615 188.455 ;
        RECT 42.790 188.270 48.615 188.410 ;
        RECT 42.790 188.210 43.110 188.270 ;
        RECT 48.325 188.225 48.615 188.270 ;
        RECT 48.785 188.410 49.075 188.455 ;
        RECT 51.070 188.410 51.390 188.470 ;
        RECT 52.465 188.410 52.755 188.455 ;
        RECT 48.785 188.270 52.755 188.410 ;
        RECT 48.785 188.225 49.075 188.270 ;
        RECT 51.070 188.210 51.390 188.270 ;
        RECT 52.465 188.225 52.755 188.270 ;
        RECT 52.925 188.410 53.215 188.455 ;
        RECT 53.370 188.410 53.690 188.470 ;
        RECT 52.925 188.270 53.690 188.410 ;
        RECT 52.925 188.225 53.215 188.270 ;
        RECT 53.370 188.210 53.690 188.270 ;
        RECT 55.670 188.210 55.990 188.470 ;
        RECT 57.140 188.455 57.280 188.610 ;
        RECT 65.420 188.455 65.560 188.950 ;
        RECT 74.070 188.890 74.390 188.950 ;
        RECT 76.370 188.890 76.690 188.950 ;
        RECT 89.265 188.905 89.555 189.135 ;
        RECT 67.170 188.550 67.490 188.810 ;
        RECT 81.380 188.750 81.670 188.795 ;
        RECT 83.730 188.750 84.050 188.810 ;
        RECT 84.640 188.750 84.930 188.795 ;
        RECT 81.380 188.610 84.930 188.750 ;
        RECT 81.380 188.565 81.670 188.610 ;
        RECT 83.730 188.550 84.050 188.610 ;
        RECT 84.640 188.565 84.930 188.610 ;
        RECT 85.560 188.750 85.850 188.795 ;
        RECT 87.420 188.750 87.710 188.795 ;
        RECT 85.560 188.610 87.710 188.750 ;
        RECT 85.560 188.565 85.850 188.610 ;
        RECT 87.420 188.565 87.710 188.610 ;
        RECT 57.065 188.225 57.355 188.455 ;
        RECT 65.345 188.225 65.635 188.455 ;
        RECT 67.630 188.410 67.950 188.470 ;
        RECT 69.930 188.410 70.250 188.470 ;
        RECT 70.865 188.410 71.155 188.455 ;
        RECT 67.630 188.270 71.155 188.410 ;
        RECT 67.630 188.210 67.950 188.270 ;
        RECT 69.930 188.210 70.250 188.270 ;
        RECT 70.865 188.225 71.155 188.270 ;
        RECT 73.165 188.410 73.455 188.455 ;
        RECT 74.530 188.410 74.850 188.470 ;
        RECT 73.165 188.270 74.850 188.410 ;
        RECT 73.165 188.225 73.455 188.270 ;
        RECT 41.870 188.070 42.190 188.130 ;
        RECT 47.405 188.070 47.695 188.115 ;
        RECT 51.545 188.070 51.835 188.115 ;
        RECT 41.870 187.930 51.835 188.070 ;
        RECT 41.870 187.870 42.190 187.930 ;
        RECT 47.405 187.885 47.695 187.930 ;
        RECT 51.545 187.885 51.835 187.930 ;
        RECT 56.130 187.870 56.450 188.130 ;
        RECT 65.790 187.870 66.110 188.130 ;
        RECT 69.010 188.070 69.330 188.130 ;
        RECT 73.240 188.070 73.380 188.225 ;
        RECT 74.530 188.210 74.850 188.270 ;
        RECT 83.240 188.410 83.530 188.455 ;
        RECT 85.560 188.410 85.775 188.565 ;
        RECT 83.240 188.270 85.775 188.410 ;
        RECT 86.505 188.410 86.795 188.455 ;
        RECT 89.340 188.410 89.480 188.905 ;
        RECT 104.430 188.795 104.750 188.810 ;
        RECT 100.865 188.750 101.155 188.795 ;
        RECT 104.105 188.750 104.755 188.795 ;
        RECT 100.865 188.610 104.755 188.750 ;
        RECT 100.865 188.565 101.455 188.610 ;
        RECT 104.105 188.565 104.755 188.610 ;
        RECT 116.505 188.750 116.795 188.795 ;
        RECT 118.690 188.750 119.010 188.810 ;
        RECT 119.745 188.750 120.395 188.795 ;
        RECT 116.505 188.610 120.395 188.750 ;
        RECT 116.505 188.565 117.095 188.610 ;
        RECT 86.505 188.270 89.480 188.410 ;
        RECT 83.240 188.225 83.530 188.270 ;
        RECT 86.505 188.225 86.795 188.270 ;
        RECT 90.170 188.210 90.490 188.470 ;
        RECT 101.165 188.250 101.455 188.565 ;
        RECT 104.430 188.550 104.750 188.565 ;
        RECT 102.245 188.410 102.535 188.455 ;
        RECT 105.825 188.410 106.115 188.455 ;
        RECT 107.660 188.410 107.950 188.455 ;
        RECT 102.245 188.270 107.950 188.410 ;
        RECT 102.245 188.225 102.535 188.270 ;
        RECT 105.825 188.225 106.115 188.270 ;
        RECT 107.660 188.225 107.950 188.270 ;
        RECT 116.805 188.250 117.095 188.565 ;
        RECT 118.690 188.550 119.010 188.610 ;
        RECT 119.745 188.565 120.395 188.610 ;
        RECT 117.885 188.410 118.175 188.455 ;
        RECT 121.465 188.410 121.755 188.455 ;
        RECT 123.300 188.410 123.590 188.455 ;
        RECT 117.885 188.270 123.590 188.410 ;
        RECT 117.885 188.225 118.175 188.270 ;
        RECT 121.465 188.225 121.755 188.270 ;
        RECT 123.300 188.225 123.590 188.270 ;
        RECT 69.010 187.930 73.380 188.070 ;
        RECT 79.375 188.070 79.665 188.115 ;
        RECT 84.190 188.070 84.510 188.130 ;
        RECT 79.375 187.930 84.510 188.070 ;
        RECT 69.010 187.870 69.330 187.930 ;
        RECT 79.375 187.885 79.665 187.930 ;
        RECT 84.190 187.870 84.510 187.930 ;
        RECT 88.345 188.070 88.635 188.115 ;
        RECT 93.390 188.070 93.710 188.130 ;
        RECT 88.345 187.930 93.710 188.070 ;
        RECT 88.345 187.885 88.635 187.930 ;
        RECT 68.105 187.730 68.395 187.775 ;
        RECT 70.390 187.730 70.710 187.790 ;
        RECT 68.105 187.590 70.710 187.730 ;
        RECT 68.105 187.545 68.395 187.590 ;
        RECT 70.390 187.530 70.710 187.590 ;
        RECT 83.240 187.730 83.530 187.775 ;
        RECT 86.020 187.730 86.310 187.775 ;
        RECT 87.880 187.730 88.170 187.775 ;
        RECT 83.240 187.590 88.170 187.730 ;
        RECT 83.240 187.545 83.530 187.590 ;
        RECT 86.020 187.545 86.310 187.590 ;
        RECT 87.880 187.545 88.170 187.590 ;
        RECT 50.625 187.390 50.915 187.435 ;
        RECT 51.530 187.390 51.850 187.450 ;
        RECT 50.625 187.250 51.850 187.390 ;
        RECT 50.625 187.205 50.915 187.250 ;
        RECT 51.530 187.190 51.850 187.250 ;
        RECT 69.945 187.390 70.235 187.435 ;
        RECT 70.850 187.390 71.170 187.450 ;
        RECT 69.945 187.250 71.170 187.390 ;
        RECT 69.945 187.205 70.235 187.250 ;
        RECT 70.850 187.190 71.170 187.250 ;
        RECT 73.625 187.390 73.915 187.435 ;
        RECT 74.070 187.390 74.390 187.450 ;
        RECT 73.625 187.250 74.390 187.390 ;
        RECT 73.625 187.205 73.915 187.250 ;
        RECT 74.070 187.190 74.390 187.250 ;
        RECT 75.910 187.390 76.230 187.450 ;
        RECT 87.410 187.390 87.730 187.450 ;
        RECT 88.420 187.390 88.560 187.885 ;
        RECT 93.390 187.870 93.710 187.930 ;
        RECT 108.125 188.070 108.415 188.115 ;
        RECT 112.250 188.070 112.570 188.130 ;
        RECT 123.765 188.070 124.055 188.115 ;
        RECT 125.590 188.070 125.910 188.130 ;
        RECT 108.125 187.930 125.910 188.070 ;
        RECT 108.125 187.885 108.415 187.930 ;
        RECT 112.250 187.870 112.570 187.930 ;
        RECT 123.765 187.885 124.055 187.930 ;
        RECT 125.590 187.870 125.910 187.930 ;
        RECT 102.245 187.730 102.535 187.775 ;
        RECT 105.365 187.730 105.655 187.775 ;
        RECT 107.255 187.730 107.545 187.775 ;
        RECT 102.245 187.590 107.545 187.730 ;
        RECT 102.245 187.545 102.535 187.590 ;
        RECT 105.365 187.545 105.655 187.590 ;
        RECT 107.255 187.545 107.545 187.590 ;
        RECT 117.885 187.730 118.175 187.775 ;
        RECT 121.005 187.730 121.295 187.775 ;
        RECT 122.895 187.730 123.185 187.775 ;
        RECT 117.885 187.590 123.185 187.730 ;
        RECT 117.885 187.545 118.175 187.590 ;
        RECT 121.005 187.545 121.295 187.590 ;
        RECT 122.895 187.545 123.185 187.590 ;
        RECT 75.910 187.250 88.560 187.390 ;
        RECT 75.910 187.190 76.230 187.250 ;
        RECT 87.410 187.190 87.730 187.250 ;
        RECT 99.370 187.190 99.690 187.450 ;
        RECT 106.840 187.390 107.130 187.435 ;
        RECT 108.110 187.390 108.430 187.450 ;
        RECT 106.840 187.250 108.430 187.390 ;
        RECT 106.840 187.205 107.130 187.250 ;
        RECT 108.110 187.190 108.430 187.250 ;
        RECT 115.025 187.390 115.315 187.435 ;
        RECT 117.310 187.390 117.630 187.450 ;
        RECT 115.025 187.250 117.630 187.390 ;
        RECT 115.025 187.205 115.315 187.250 ;
        RECT 117.310 187.190 117.630 187.250 ;
        RECT 122.480 187.390 122.770 187.435 ;
        RECT 124.210 187.390 124.530 187.450 ;
        RECT 122.480 187.250 124.530 187.390 ;
        RECT 122.480 187.205 122.770 187.250 ;
        RECT 124.210 187.190 124.530 187.250 ;
        RECT 14.660 186.570 127.820 187.050 ;
        RECT 49.230 186.370 49.550 186.430 ;
        RECT 50.625 186.370 50.915 186.415 ;
        RECT 49.230 186.230 50.915 186.370 ;
        RECT 49.230 186.170 49.550 186.230 ;
        RECT 50.625 186.185 50.915 186.230 ;
        RECT 86.505 186.370 86.795 186.415 ;
        RECT 90.170 186.370 90.490 186.430 ;
        RECT 86.505 186.230 90.490 186.370 ;
        RECT 86.505 186.185 86.795 186.230 ;
        RECT 90.170 186.170 90.490 186.230 ;
        RECT 108.110 186.170 108.430 186.430 ;
        RECT 124.210 186.170 124.530 186.430 ;
        RECT 56.560 186.030 56.850 186.075 ;
        RECT 59.340 186.030 59.630 186.075 ;
        RECT 61.200 186.030 61.490 186.075 ;
        RECT 56.560 185.890 61.490 186.030 ;
        RECT 56.560 185.845 56.850 185.890 ;
        RECT 59.340 185.845 59.630 185.890 ;
        RECT 61.200 185.845 61.490 185.890 ;
        RECT 66.250 185.830 66.570 186.090 ;
        RECT 69.585 186.030 69.875 186.075 ;
        RECT 72.705 186.030 72.995 186.075 ;
        RECT 74.595 186.030 74.885 186.075 ;
        RECT 69.585 185.890 74.885 186.030 ;
        RECT 69.585 185.845 69.875 185.890 ;
        RECT 72.705 185.845 72.995 185.890 ;
        RECT 74.595 185.845 74.885 185.890 ;
        RECT 104.430 186.030 104.750 186.090 ;
        RECT 107.205 186.030 107.495 186.075 ;
        RECT 104.430 185.890 107.495 186.030 ;
        RECT 104.430 185.830 104.750 185.890 ;
        RECT 107.205 185.845 107.495 185.890 ;
        RECT 115.025 186.030 115.315 186.075 ;
        RECT 116.850 186.030 117.170 186.090 ;
        RECT 115.025 185.890 117.170 186.030 ;
        RECT 115.025 185.845 115.315 185.890 ;
        RECT 116.850 185.830 117.170 185.890 ;
        RECT 117.885 186.030 118.175 186.075 ;
        RECT 121.005 186.030 121.295 186.075 ;
        RECT 122.895 186.030 123.185 186.075 ;
        RECT 117.885 185.890 123.185 186.030 ;
        RECT 117.885 185.845 118.175 185.890 ;
        RECT 121.005 185.845 121.295 185.890 ;
        RECT 122.895 185.845 123.185 185.890 ;
        RECT 31.290 185.690 31.610 185.750 ;
        RECT 37.745 185.690 38.035 185.735 ;
        RECT 31.290 185.550 38.035 185.690 ;
        RECT 31.290 185.490 31.610 185.550 ;
        RECT 37.745 185.505 38.035 185.550 ;
        RECT 38.665 185.690 38.955 185.735 ;
        RECT 41.870 185.690 42.190 185.750 ;
        RECT 38.665 185.550 42.190 185.690 ;
        RECT 38.665 185.505 38.955 185.550 ;
        RECT 41.870 185.490 42.190 185.550 ;
        RECT 42.330 185.690 42.650 185.750 ;
        RECT 42.805 185.690 43.095 185.735 ;
        RECT 42.330 185.550 43.095 185.690 ;
        RECT 42.330 185.490 42.650 185.550 ;
        RECT 42.805 185.505 43.095 185.550 ;
        RECT 63.045 185.690 63.335 185.735 ;
        RECT 64.870 185.690 65.190 185.750 ;
        RECT 63.045 185.550 65.190 185.690 ;
        RECT 63.045 185.505 63.335 185.550 ;
        RECT 64.870 185.490 65.190 185.550 ;
        RECT 65.470 185.690 65.760 185.735 ;
        RECT 67.170 185.690 67.490 185.750 ;
        RECT 65.470 185.550 67.490 185.690 ;
        RECT 65.470 185.505 65.760 185.550 ;
        RECT 67.170 185.490 67.490 185.550 ;
        RECT 74.070 185.490 74.390 185.750 ;
        RECT 75.465 185.690 75.755 185.735 ;
        RECT 75.910 185.690 76.230 185.750 ;
        RECT 75.465 185.550 76.230 185.690 ;
        RECT 75.465 185.505 75.755 185.550 ;
        RECT 75.910 185.490 76.230 185.550 ;
        RECT 83.745 185.690 84.035 185.735 ;
        RECT 85.110 185.690 85.430 185.750 ;
        RECT 98.005 185.690 98.295 185.735 ;
        RECT 103.065 185.690 103.355 185.735 ;
        RECT 105.350 185.690 105.670 185.750 ;
        RECT 125.590 185.690 125.910 185.750 ;
        RECT 83.745 185.550 105.670 185.690 ;
        RECT 83.745 185.505 84.035 185.550 ;
        RECT 85.110 185.490 85.430 185.550 ;
        RECT 98.005 185.505 98.295 185.550 ;
        RECT 103.065 185.505 103.355 185.550 ;
        RECT 105.350 185.490 105.670 185.550 ;
        RECT 124.300 185.550 125.910 185.690 ;
        RECT 124.300 185.410 124.440 185.550 ;
        RECT 125.590 185.490 125.910 185.550 ;
        RECT 33.145 185.350 33.435 185.395 ;
        RECT 34.050 185.350 34.370 185.410 ;
        RECT 33.145 185.210 34.370 185.350 ;
        RECT 33.145 185.165 33.435 185.210 ;
        RECT 34.050 185.150 34.370 185.210 ;
        RECT 43.265 185.165 43.555 185.395 ;
        RECT 37.285 185.010 37.575 185.055 ;
        RECT 42.330 185.010 42.650 185.070 ;
        RECT 37.285 184.870 42.650 185.010 ;
        RECT 37.285 184.825 37.575 184.870 ;
        RECT 42.330 184.810 42.650 184.870 ;
        RECT 42.790 185.010 43.110 185.070 ;
        RECT 43.340 185.010 43.480 185.165 ;
        RECT 51.530 185.150 51.850 185.410 ;
        RECT 56.560 185.350 56.850 185.395 ;
        RECT 56.560 185.210 59.095 185.350 ;
        RECT 56.560 185.165 56.850 185.210 ;
        RECT 42.790 184.870 43.480 185.010 ;
        RECT 54.700 185.010 54.990 185.055 ;
        RECT 56.130 185.010 56.450 185.070 ;
        RECT 58.880 185.055 59.095 185.210 ;
        RECT 59.810 185.150 60.130 185.410 ;
        RECT 61.665 185.165 61.955 185.395 ;
        RECT 64.425 185.350 64.715 185.395 ;
        RECT 67.630 185.350 67.950 185.410 ;
        RECT 64.425 185.210 67.950 185.350 ;
        RECT 64.425 185.165 64.715 185.210 ;
        RECT 57.960 185.010 58.250 185.055 ;
        RECT 54.700 184.870 58.250 185.010 ;
        RECT 42.790 184.810 43.110 184.870 ;
        RECT 54.700 184.825 54.990 184.870 ;
        RECT 56.130 184.810 56.450 184.870 ;
        RECT 57.960 184.825 58.250 184.870 ;
        RECT 58.880 185.010 59.170 185.055 ;
        RECT 60.740 185.010 61.030 185.055 ;
        RECT 58.880 184.870 61.030 185.010 ;
        RECT 58.880 184.825 59.170 184.870 ;
        RECT 60.740 184.825 61.030 184.870 ;
        RECT 32.670 184.470 32.990 184.730 ;
        RECT 35.445 184.670 35.735 184.715 ;
        RECT 36.350 184.670 36.670 184.730 ;
        RECT 35.445 184.530 36.670 184.670 ;
        RECT 35.445 184.485 35.735 184.530 ;
        RECT 36.350 184.470 36.670 184.530 ;
        RECT 43.250 184.670 43.570 184.730 ;
        RECT 45.105 184.670 45.395 184.715 ;
        RECT 43.250 184.530 45.395 184.670 ;
        RECT 43.250 184.470 43.570 184.530 ;
        RECT 45.105 184.485 45.395 184.530 ;
        RECT 52.695 184.670 52.985 184.715 ;
        RECT 53.370 184.670 53.690 184.730 ;
        RECT 52.695 184.530 53.690 184.670 ;
        RECT 52.695 184.485 52.985 184.530 ;
        RECT 53.370 184.470 53.690 184.530 ;
        RECT 56.590 184.670 56.910 184.730 ;
        RECT 61.740 184.670 61.880 185.165 ;
        RECT 67.630 185.150 67.950 185.210 ;
        RECT 65.790 185.010 66.110 185.070 ;
        RECT 68.505 185.055 68.795 185.370 ;
        RECT 69.585 185.350 69.875 185.395 ;
        RECT 73.165 185.350 73.455 185.395 ;
        RECT 75.000 185.350 75.290 185.395 ;
        RECT 69.585 185.210 75.290 185.350 ;
        RECT 69.585 185.165 69.875 185.210 ;
        RECT 73.165 185.165 73.455 185.210 ;
        RECT 75.000 185.165 75.290 185.210 ;
        RECT 82.365 185.350 82.655 185.395 ;
        RECT 83.270 185.350 83.590 185.410 ;
        RECT 82.365 185.210 83.590 185.350 ;
        RECT 82.365 185.165 82.655 185.210 ;
        RECT 83.270 185.150 83.590 185.210 ;
        RECT 99.370 185.350 99.690 185.410 ;
        RECT 102.130 185.350 102.450 185.410 ;
        RECT 103.985 185.350 104.275 185.395 ;
        RECT 107.665 185.350 107.955 185.395 ;
        RECT 99.370 185.210 104.275 185.350 ;
        RECT 99.370 185.150 99.690 185.210 ;
        RECT 102.130 185.150 102.450 185.210 ;
        RECT 103.985 185.165 104.275 185.210 ;
        RECT 104.520 185.210 107.955 185.350 ;
        RECT 68.205 185.010 68.795 185.055 ;
        RECT 71.445 185.010 72.095 185.055 ;
        RECT 65.790 184.870 72.095 185.010 ;
        RECT 65.790 184.810 66.110 184.870 ;
        RECT 68.205 184.825 68.495 184.870 ;
        RECT 71.445 184.825 72.095 184.870 ;
        RECT 80.050 185.010 80.370 185.070 ;
        RECT 84.665 185.010 84.955 185.055 ;
        RECT 80.050 184.870 84.955 185.010 ;
        RECT 80.050 184.810 80.370 184.870 ;
        RECT 84.665 184.825 84.955 184.870 ;
        RECT 102.590 185.010 102.910 185.070 ;
        RECT 104.520 185.010 104.660 185.210 ;
        RECT 107.665 185.165 107.955 185.210 ;
        RECT 109.045 185.165 109.335 185.395 ;
        RECT 109.120 185.010 109.260 185.165 ;
        RECT 113.630 185.150 113.950 185.410 ;
        RECT 116.805 185.055 117.095 185.370 ;
        RECT 117.885 185.350 118.175 185.395 ;
        RECT 121.465 185.350 121.755 185.395 ;
        RECT 123.300 185.350 123.590 185.395 ;
        RECT 117.885 185.210 123.590 185.350 ;
        RECT 117.885 185.165 118.175 185.210 ;
        RECT 121.465 185.165 121.755 185.210 ;
        RECT 123.300 185.165 123.590 185.210 ;
        RECT 123.765 185.350 124.055 185.395 ;
        RECT 124.210 185.350 124.530 185.410 ;
        RECT 123.765 185.210 124.530 185.350 ;
        RECT 123.765 185.165 124.055 185.210 ;
        RECT 124.210 185.150 124.530 185.210 ;
        RECT 125.145 185.165 125.435 185.395 ;
        RECT 102.590 184.870 104.660 185.010 ;
        RECT 106.360 184.870 109.260 185.010 ;
        RECT 114.105 185.010 114.395 185.055 ;
        RECT 116.505 185.010 117.095 185.055 ;
        RECT 119.745 185.010 120.395 185.055 ;
        RECT 114.105 184.870 120.395 185.010 ;
        RECT 102.590 184.810 102.910 184.870 ;
        RECT 56.590 184.530 61.880 184.670 ;
        RECT 64.885 184.670 65.175 184.715 ;
        RECT 66.710 184.670 67.030 184.730 ;
        RECT 64.885 184.530 67.030 184.670 ;
        RECT 56.590 184.470 56.910 184.530 ;
        RECT 64.885 184.485 65.175 184.530 ;
        RECT 66.710 184.470 67.030 184.530 ;
        RECT 81.905 184.670 82.195 184.715 ;
        RECT 82.350 184.670 82.670 184.730 ;
        RECT 81.905 184.530 82.670 184.670 ;
        RECT 81.905 184.485 82.195 184.530 ;
        RECT 82.350 184.470 82.670 184.530 ;
        RECT 84.190 184.470 84.510 184.730 ;
        RECT 98.925 184.670 99.215 184.715 ;
        RECT 99.830 184.670 100.150 184.730 ;
        RECT 98.925 184.530 100.150 184.670 ;
        RECT 98.925 184.485 99.215 184.530 ;
        RECT 99.830 184.470 100.150 184.530 ;
        RECT 101.225 184.670 101.515 184.715 ;
        RECT 103.510 184.670 103.830 184.730 ;
        RECT 101.225 184.530 103.830 184.670 ;
        RECT 101.225 184.485 101.515 184.530 ;
        RECT 103.510 184.470 103.830 184.530 ;
        RECT 103.970 184.670 104.290 184.730 ;
        RECT 106.360 184.715 106.500 184.870 ;
        RECT 114.105 184.825 114.395 184.870 ;
        RECT 116.505 184.825 116.795 184.870 ;
        RECT 119.745 184.825 120.395 184.870 ;
        RECT 122.370 184.810 122.690 185.070 ;
        RECT 104.445 184.670 104.735 184.715 ;
        RECT 103.970 184.530 104.735 184.670 ;
        RECT 103.970 184.470 104.290 184.530 ;
        RECT 104.445 184.485 104.735 184.530 ;
        RECT 106.285 184.485 106.575 184.715 ;
        RECT 118.690 184.670 119.010 184.730 ;
        RECT 125.220 184.670 125.360 185.165 ;
        RECT 118.690 184.530 125.360 184.670 ;
        RECT 118.690 184.470 119.010 184.530 ;
        RECT 14.660 183.850 127.820 184.330 ;
        RECT 28.085 183.650 28.375 183.695 ;
        RECT 31.290 183.650 31.610 183.710 ;
        RECT 28.085 183.510 31.610 183.650 ;
        RECT 28.085 183.465 28.375 183.510 ;
        RECT 31.290 183.450 31.610 183.510 ;
        RECT 58.905 183.650 59.195 183.695 ;
        RECT 59.810 183.650 60.130 183.710 ;
        RECT 58.905 183.510 60.130 183.650 ;
        RECT 58.905 183.465 59.195 183.510 ;
        RECT 59.810 183.450 60.130 183.510 ;
        RECT 66.265 183.465 66.555 183.695 ;
        RECT 67.170 183.650 67.490 183.710 ;
        RECT 68.565 183.650 68.855 183.695 ;
        RECT 100.290 183.650 100.610 183.710 ;
        RECT 102.605 183.650 102.895 183.695 ;
        RECT 67.170 183.510 68.855 183.650 ;
        RECT 32.670 183.355 32.990 183.370 ;
        RECT 29.565 183.310 29.855 183.355 ;
        RECT 32.670 183.310 33.455 183.355 ;
        RECT 29.565 183.170 33.455 183.310 ;
        RECT 29.565 183.125 30.155 183.170 ;
        RECT 29.865 182.810 30.155 183.125 ;
        RECT 32.670 183.125 33.455 183.170 ;
        RECT 32.670 183.110 32.990 183.125 ;
        RECT 35.430 183.110 35.750 183.370 ;
        RECT 35.890 183.310 36.210 183.370 ;
        RECT 39.225 183.310 39.515 183.355 ;
        RECT 42.465 183.310 43.115 183.355 ;
        RECT 35.890 183.170 43.115 183.310 ;
        RECT 66.340 183.310 66.480 183.465 ;
        RECT 67.170 183.450 67.490 183.510 ;
        RECT 68.565 183.465 68.855 183.510 ;
        RECT 92.100 183.510 100.610 183.650 ;
        RECT 69.010 183.310 69.330 183.370 ;
        RECT 66.340 183.170 69.330 183.310 ;
        RECT 35.890 183.110 36.210 183.170 ;
        RECT 39.225 183.125 39.815 183.170 ;
        RECT 42.465 183.125 43.115 183.170 ;
        RECT 30.945 182.970 31.235 183.015 ;
        RECT 34.525 182.970 34.815 183.015 ;
        RECT 36.360 182.970 36.650 183.015 ;
        RECT 30.945 182.830 36.650 182.970 ;
        RECT 30.945 182.785 31.235 182.830 ;
        RECT 34.525 182.785 34.815 182.830 ;
        RECT 36.360 182.785 36.650 182.830 ;
        RECT 39.525 182.810 39.815 183.125 ;
        RECT 69.010 183.110 69.330 183.170 ;
        RECT 70.865 183.310 71.155 183.355 ;
        RECT 72.230 183.310 72.550 183.370 ;
        RECT 70.865 183.170 72.550 183.310 ;
        RECT 70.865 183.125 71.155 183.170 ;
        RECT 72.230 183.110 72.550 183.170 ;
        RECT 76.370 183.110 76.690 183.370 ;
        RECT 80.165 183.310 80.455 183.355 ;
        RECT 82.350 183.310 82.670 183.370 ;
        RECT 83.405 183.310 84.055 183.355 ;
        RECT 80.165 183.170 84.055 183.310 ;
        RECT 80.165 183.125 80.755 183.170 ;
        RECT 40.605 182.970 40.895 183.015 ;
        RECT 44.185 182.970 44.475 183.015 ;
        RECT 46.020 182.970 46.310 183.015 ;
        RECT 40.605 182.830 46.310 182.970 ;
        RECT 40.605 182.785 40.895 182.830 ;
        RECT 44.185 182.785 44.475 182.830 ;
        RECT 46.020 182.785 46.310 182.830 ;
        RECT 57.970 182.770 58.290 183.030 ;
        RECT 65.345 182.970 65.635 183.015 ;
        RECT 66.710 182.970 67.030 183.030 ;
        RECT 68.105 182.970 68.395 183.015 ;
        RECT 65.345 182.830 68.395 182.970 ;
        RECT 65.345 182.785 65.635 182.830 ;
        RECT 66.710 182.770 67.030 182.830 ;
        RECT 68.105 182.785 68.395 182.830 ;
        RECT 74.990 182.770 75.310 183.030 ;
        RECT 80.465 182.810 80.755 183.125 ;
        RECT 82.350 183.110 82.670 183.170 ;
        RECT 83.405 183.125 84.055 183.170 ;
        RECT 86.045 183.310 86.335 183.355 ;
        RECT 86.490 183.310 86.810 183.370 ;
        RECT 86.045 183.170 86.810 183.310 ;
        RECT 86.045 183.125 86.335 183.170 ;
        RECT 86.490 183.110 86.810 183.170 ;
        RECT 81.545 182.970 81.835 183.015 ;
        RECT 85.125 182.970 85.415 183.015 ;
        RECT 86.960 182.970 87.250 183.015 ;
        RECT 81.545 182.830 87.250 182.970 ;
        RECT 81.545 182.785 81.835 182.830 ;
        RECT 85.125 182.785 85.415 182.830 ;
        RECT 86.960 182.785 87.250 182.830 ;
        RECT 87.410 182.770 87.730 183.030 ;
        RECT 90.630 182.770 90.950 183.030 ;
        RECT 92.100 183.015 92.240 183.510 ;
        RECT 100.290 183.450 100.610 183.510 ;
        RECT 100.840 183.510 102.895 183.650 ;
        RECT 100.840 183.355 100.980 183.510 ;
        RECT 102.605 183.465 102.895 183.510 ;
        RECT 118.690 183.450 119.010 183.710 ;
        RECT 120.545 183.650 120.835 183.695 ;
        RECT 122.370 183.650 122.690 183.710 ;
        RECT 120.545 183.510 122.690 183.650 ;
        RECT 120.545 183.465 120.835 183.510 ;
        RECT 122.370 183.450 122.690 183.510 ;
        RECT 92.485 183.310 92.775 183.355 ;
        RECT 94.885 183.310 95.175 183.355 ;
        RECT 98.125 183.310 98.775 183.355 ;
        RECT 92.485 183.170 98.775 183.310 ;
        RECT 92.485 183.125 92.775 183.170 ;
        RECT 94.885 183.125 95.475 183.170 ;
        RECT 98.125 183.125 98.775 183.170 ;
        RECT 100.765 183.125 101.055 183.355 ;
        RECT 101.210 183.310 101.530 183.370 ;
        RECT 110.885 183.310 111.175 183.355 ;
        RECT 101.210 183.170 111.175 183.310 ;
        RECT 92.025 182.785 92.315 183.015 ;
        RECT 95.185 182.810 95.475 183.125 ;
        RECT 101.210 183.110 101.530 183.170 ;
        RECT 110.885 183.125 111.175 183.170 ;
        RECT 96.265 182.970 96.555 183.015 ;
        RECT 99.845 182.970 100.135 183.015 ;
        RECT 101.680 182.970 101.970 183.015 ;
        RECT 96.265 182.830 101.970 182.970 ;
        RECT 96.265 182.785 96.555 182.830 ;
        RECT 99.845 182.785 100.135 182.830 ;
        RECT 101.680 182.785 101.970 182.830 ;
        RECT 103.510 182.770 103.830 183.030 ;
        RECT 107.665 182.785 107.955 183.015 ;
        RECT 109.030 182.970 109.350 183.030 ;
        RECT 110.425 182.970 110.715 183.015 ;
        RECT 109.030 182.830 110.715 182.970 ;
        RECT 30.370 182.630 30.690 182.690 ;
        RECT 36.825 182.630 37.115 182.675 ;
        RECT 30.370 182.490 37.115 182.630 ;
        RECT 30.370 182.430 30.690 182.490 ;
        RECT 36.825 182.445 37.115 182.490 ;
        RECT 45.090 182.430 45.410 182.690 ;
        RECT 46.485 182.630 46.775 182.675 ;
        RECT 56.590 182.630 56.910 182.690 ;
        RECT 46.485 182.490 56.910 182.630 ;
        RECT 46.485 182.445 46.775 182.490 ;
        RECT 56.590 182.430 56.910 182.490 ;
        RECT 100.750 182.630 101.070 182.690 ;
        RECT 102.145 182.630 102.435 182.675 ;
        RECT 100.750 182.490 102.435 182.630 ;
        RECT 100.750 182.430 101.070 182.490 ;
        RECT 102.145 182.445 102.435 182.490 ;
        RECT 30.945 182.290 31.235 182.335 ;
        RECT 34.065 182.290 34.355 182.335 ;
        RECT 35.955 182.290 36.245 182.335 ;
        RECT 30.945 182.150 36.245 182.290 ;
        RECT 30.945 182.105 31.235 182.150 ;
        RECT 34.065 182.105 34.355 182.150 ;
        RECT 35.955 182.105 36.245 182.150 ;
        RECT 40.605 182.290 40.895 182.335 ;
        RECT 43.725 182.290 44.015 182.335 ;
        RECT 45.615 182.290 45.905 182.335 ;
        RECT 40.605 182.150 45.905 182.290 ;
        RECT 40.605 182.105 40.895 182.150 ;
        RECT 43.725 182.105 44.015 182.150 ;
        RECT 45.615 182.105 45.905 182.150 ;
        RECT 70.850 182.090 71.170 182.350 ;
        RECT 81.545 182.290 81.835 182.335 ;
        RECT 84.665 182.290 84.955 182.335 ;
        RECT 86.555 182.290 86.845 182.335 ;
        RECT 81.545 182.150 86.845 182.290 ;
        RECT 81.545 182.105 81.835 182.150 ;
        RECT 84.665 182.105 84.955 182.150 ;
        RECT 86.555 182.105 86.845 182.150 ;
        RECT 96.265 182.290 96.555 182.335 ;
        RECT 99.385 182.290 99.675 182.335 ;
        RECT 101.275 182.290 101.565 182.335 ;
        RECT 96.265 182.150 101.565 182.290 ;
        RECT 96.265 182.105 96.555 182.150 ;
        RECT 99.385 182.105 99.675 182.150 ;
        RECT 101.275 182.105 101.565 182.150 ;
        RECT 107.740 182.290 107.880 182.785 ;
        RECT 109.030 182.770 109.350 182.830 ;
        RECT 110.425 182.785 110.715 182.830 ;
        RECT 116.850 182.770 117.170 183.030 ;
        RECT 119.610 182.770 119.930 183.030 ;
        RECT 109.965 182.630 110.255 182.675 ;
        RECT 115.945 182.630 116.235 182.675 ;
        RECT 109.965 182.490 116.235 182.630 ;
        RECT 109.965 182.445 110.255 182.490 ;
        RECT 115.945 182.445 116.235 182.490 ;
        RECT 116.405 182.630 116.695 182.675 ;
        RECT 117.310 182.630 117.630 182.690 ;
        RECT 116.405 182.490 117.630 182.630 ;
        RECT 116.405 182.445 116.695 182.490 ;
        RECT 113.630 182.290 113.950 182.350 ;
        RECT 107.740 182.150 113.950 182.290 ;
        RECT 116.020 182.290 116.160 182.445 ;
        RECT 117.310 182.430 117.630 182.490 ;
        RECT 118.230 182.290 118.550 182.350 ;
        RECT 116.020 182.150 118.550 182.290 ;
        RECT 37.745 181.950 38.035 181.995 ;
        RECT 42.330 181.950 42.650 182.010 ;
        RECT 37.745 181.810 42.650 181.950 ;
        RECT 37.745 181.765 38.035 181.810 ;
        RECT 42.330 181.750 42.650 181.810 ;
        RECT 66.250 181.950 66.570 182.010 ;
        RECT 67.185 181.950 67.475 181.995 ;
        RECT 66.250 181.810 67.475 181.950 ;
        RECT 66.250 181.750 66.570 181.810 ;
        RECT 67.185 181.765 67.475 181.810 ;
        RECT 78.685 181.950 78.975 181.995 ;
        RECT 80.050 181.950 80.370 182.010 ;
        RECT 78.685 181.810 80.370 181.950 ;
        RECT 78.685 181.765 78.975 181.810 ;
        RECT 80.050 181.750 80.370 181.810 ;
        RECT 91.090 181.950 91.410 182.010 ;
        RECT 91.565 181.950 91.855 181.995 ;
        RECT 91.090 181.810 91.855 181.950 ;
        RECT 91.090 181.750 91.410 181.810 ;
        RECT 91.565 181.765 91.855 181.810 ;
        RECT 93.405 181.950 93.695 181.995 ;
        RECT 99.830 181.950 100.150 182.010 ;
        RECT 93.405 181.810 100.150 181.950 ;
        RECT 93.405 181.765 93.695 181.810 ;
        RECT 99.830 181.750 100.150 181.810 ;
        RECT 100.290 181.950 100.610 182.010 ;
        RECT 107.740 181.950 107.880 182.150 ;
        RECT 113.630 182.090 113.950 182.150 ;
        RECT 118.230 182.090 118.550 182.150 ;
        RECT 100.290 181.810 107.880 181.950 ;
        RECT 100.290 181.750 100.610 181.810 ;
        RECT 108.110 181.750 108.430 182.010 ;
        RECT 112.725 181.950 113.015 181.995 ;
        RECT 113.170 181.950 113.490 182.010 ;
        RECT 112.725 181.810 113.490 181.950 ;
        RECT 112.725 181.765 113.015 181.810 ;
        RECT 113.170 181.750 113.490 181.810 ;
        RECT 14.660 181.130 127.820 181.610 ;
        RECT 35.890 180.930 36.210 180.990 ;
        RECT 36.365 180.930 36.655 180.975 ;
        RECT 35.890 180.790 36.655 180.930 ;
        RECT 35.890 180.730 36.210 180.790 ;
        RECT 36.365 180.745 36.655 180.790 ;
        RECT 44.185 180.930 44.475 180.975 ;
        RECT 45.090 180.930 45.410 180.990 ;
        RECT 44.185 180.790 45.410 180.930 ;
        RECT 44.185 180.745 44.475 180.790 ;
        RECT 45.090 180.730 45.410 180.790 ;
        RECT 57.525 180.930 57.815 180.975 ;
        RECT 57.970 180.930 58.290 180.990 ;
        RECT 57.525 180.790 58.290 180.930 ;
        RECT 57.525 180.745 57.815 180.790 ;
        RECT 57.970 180.730 58.290 180.790 ;
        RECT 119.610 180.930 119.930 180.990 ;
        RECT 121.465 180.930 121.755 180.975 ;
        RECT 119.610 180.790 121.755 180.930 ;
        RECT 119.610 180.730 119.930 180.790 ;
        RECT 121.465 180.745 121.755 180.790 ;
        RECT 25.735 180.590 26.025 180.635 ;
        RECT 27.625 180.590 27.915 180.635 ;
        RECT 30.745 180.590 31.035 180.635 ;
        RECT 25.735 180.450 31.035 180.590 ;
        RECT 25.735 180.405 26.025 180.450 ;
        RECT 27.625 180.405 27.915 180.450 ;
        RECT 30.745 180.405 31.035 180.450 ;
        RECT 35.430 180.590 35.750 180.650 ;
        RECT 37.285 180.590 37.575 180.635 ;
        RECT 55.670 180.590 55.990 180.650 ;
        RECT 35.430 180.450 37.575 180.590 ;
        RECT 35.430 180.390 35.750 180.450 ;
        RECT 37.285 180.405 37.575 180.450 ;
        RECT 52.540 180.450 55.990 180.590 ;
        RECT 23.485 180.250 23.775 180.295 ;
        RECT 23.485 180.110 31.980 180.250 ;
        RECT 23.485 180.065 23.775 180.110 ;
        RECT 23.010 179.710 23.330 179.970 ;
        RECT 24.865 179.725 25.155 179.955 ;
        RECT 25.330 179.910 25.620 179.955 ;
        RECT 27.165 179.910 27.455 179.955 ;
        RECT 30.745 179.910 31.035 179.955 ;
        RECT 31.840 179.930 31.980 180.110 ;
        RECT 25.330 179.770 31.035 179.910 ;
        RECT 25.330 179.725 25.620 179.770 ;
        RECT 27.165 179.725 27.455 179.770 ;
        RECT 30.745 179.725 31.035 179.770 ;
        RECT 24.940 179.230 25.080 179.725 ;
        RECT 26.230 179.370 26.550 179.630 ;
        RECT 31.825 179.615 32.115 179.930 ;
        RECT 34.050 179.910 34.370 179.970 ;
        RECT 35.890 179.910 36.210 179.970 ;
        RECT 34.050 179.770 36.210 179.910 ;
        RECT 34.050 179.710 34.370 179.770 ;
        RECT 35.890 179.710 36.210 179.770 ;
        RECT 36.350 179.910 36.670 179.970 ;
        RECT 38.205 179.910 38.495 179.955 ;
        RECT 36.350 179.770 38.495 179.910 ;
        RECT 36.350 179.710 36.670 179.770 ;
        RECT 38.205 179.725 38.495 179.770 ;
        RECT 43.250 179.710 43.570 179.970 ;
        RECT 52.540 179.955 52.680 180.450 ;
        RECT 55.670 180.390 55.990 180.450 ;
        RECT 87.065 180.590 87.355 180.635 ;
        RECT 90.185 180.590 90.475 180.635 ;
        RECT 92.075 180.590 92.365 180.635 ;
        RECT 87.065 180.450 92.365 180.590 ;
        RECT 87.065 180.405 87.355 180.450 ;
        RECT 90.185 180.405 90.475 180.450 ;
        RECT 92.075 180.405 92.365 180.450 ;
        RECT 111.445 180.590 111.735 180.635 ;
        RECT 114.565 180.590 114.855 180.635 ;
        RECT 116.455 180.590 116.745 180.635 ;
        RECT 111.445 180.450 116.745 180.590 ;
        RECT 111.445 180.405 111.735 180.450 ;
        RECT 114.565 180.405 114.855 180.450 ;
        RECT 116.455 180.405 116.745 180.450 ;
        RECT 54.750 180.050 55.070 180.310 ;
        RECT 80.510 180.250 80.830 180.310 ;
        RECT 85.110 180.250 85.430 180.310 ;
        RECT 80.510 180.110 85.430 180.250 ;
        RECT 80.510 180.050 80.830 180.110 ;
        RECT 85.110 180.050 85.430 180.110 ;
        RECT 91.090 180.250 91.410 180.310 ;
        RECT 91.565 180.250 91.855 180.295 ;
        RECT 91.090 180.110 91.855 180.250 ;
        RECT 91.090 180.050 91.410 180.110 ;
        RECT 91.565 180.065 91.855 180.110 ;
        RECT 109.030 180.250 109.350 180.310 ;
        RECT 109.030 180.110 118.000 180.250 ;
        RECT 109.030 180.050 109.350 180.110 ;
        RECT 49.705 179.910 49.995 179.955 ;
        RECT 52.465 179.910 52.755 179.955 ;
        RECT 49.705 179.770 52.755 179.910 ;
        RECT 49.705 179.725 49.995 179.770 ;
        RECT 52.465 179.725 52.755 179.770 ;
        RECT 53.370 179.910 53.690 179.970 ;
        RECT 55.225 179.910 55.515 179.955 ;
        RECT 53.370 179.770 55.515 179.910 ;
        RECT 53.370 179.710 53.690 179.770 ;
        RECT 55.225 179.725 55.515 179.770 ;
        RECT 57.970 179.710 58.290 179.970 ;
        RECT 63.950 179.910 64.270 179.970 ;
        RECT 74.990 179.910 75.310 179.970 ;
        RECT 77.305 179.910 77.595 179.955 ;
        RECT 63.950 179.770 77.595 179.910 ;
        RECT 63.950 179.710 64.270 179.770 ;
        RECT 74.990 179.710 75.310 179.770 ;
        RECT 77.305 179.725 77.595 179.770 ;
        RECT 78.685 179.910 78.975 179.955 ;
        RECT 83.270 179.910 83.590 179.970 ;
        RECT 78.685 179.770 83.590 179.910 ;
        RECT 78.685 179.725 78.975 179.770 ;
        RECT 83.270 179.710 83.590 179.770 ;
        RECT 28.525 179.570 29.175 179.615 ;
        RECT 31.825 179.570 32.415 179.615 ;
        RECT 28.525 179.430 32.415 179.570 ;
        RECT 28.525 179.385 29.175 179.430 ;
        RECT 32.125 179.385 32.415 179.430 ;
        RECT 54.290 179.570 54.610 179.630 ;
        RECT 55.685 179.570 55.975 179.615 ;
        RECT 54.290 179.430 55.975 179.570 ;
        RECT 54.290 179.370 54.610 179.430 ;
        RECT 55.685 179.385 55.975 179.430 ;
        RECT 72.230 179.570 72.550 179.630 ;
        RECT 85.985 179.615 86.275 179.930 ;
        RECT 87.065 179.910 87.355 179.955 ;
        RECT 90.645 179.910 90.935 179.955 ;
        RECT 92.480 179.910 92.770 179.955 ;
        RECT 87.065 179.770 92.770 179.910 ;
        RECT 87.065 179.725 87.355 179.770 ;
        RECT 90.645 179.725 90.935 179.770 ;
        RECT 92.480 179.725 92.770 179.770 ;
        RECT 92.945 179.910 93.235 179.955 ;
        RECT 100.750 179.910 101.070 179.970 ;
        RECT 92.945 179.770 101.070 179.910 ;
        RECT 92.945 179.725 93.235 179.770 ;
        RECT 81.905 179.570 82.195 179.615 ;
        RECT 85.685 179.570 86.275 179.615 ;
        RECT 87.870 179.570 88.190 179.630 ;
        RECT 88.925 179.570 89.575 179.615 ;
        RECT 93.020 179.570 93.160 179.725 ;
        RECT 100.750 179.710 101.070 179.770 ;
        RECT 72.230 179.430 84.420 179.570 ;
        RECT 72.230 179.370 72.550 179.430 ;
        RECT 81.905 179.385 82.195 179.430 ;
        RECT 84.280 179.290 84.420 179.430 ;
        RECT 85.685 179.430 89.575 179.570 ;
        RECT 85.685 179.385 85.975 179.430 ;
        RECT 87.870 179.370 88.190 179.430 ;
        RECT 88.925 179.385 89.575 179.430 ;
        RECT 92.560 179.430 93.160 179.570 ;
        RECT 108.110 179.570 108.430 179.630 ;
        RECT 110.365 179.615 110.655 179.930 ;
        RECT 111.445 179.910 111.735 179.955 ;
        RECT 115.025 179.910 115.315 179.955 ;
        RECT 116.860 179.910 117.150 179.955 ;
        RECT 111.445 179.770 117.150 179.910 ;
        RECT 111.445 179.725 111.735 179.770 ;
        RECT 115.025 179.725 115.315 179.770 ;
        RECT 116.860 179.725 117.150 179.770 ;
        RECT 117.325 179.725 117.615 179.955 ;
        RECT 117.860 179.910 118.000 180.110 ;
        RECT 118.230 180.050 118.550 180.310 ;
        RECT 119.625 179.910 119.915 179.955 ;
        RECT 117.860 179.770 119.915 179.910 ;
        RECT 119.625 179.725 119.915 179.770 ;
        RECT 110.065 179.570 110.655 179.615 ;
        RECT 113.305 179.570 113.955 179.615 ;
        RECT 108.110 179.430 113.955 179.570 ;
        RECT 30.370 179.230 30.690 179.290 ;
        RECT 24.940 179.090 30.690 179.230 ;
        RECT 30.370 179.030 30.690 179.090 ;
        RECT 30.830 179.230 31.150 179.290 ;
        RECT 33.605 179.230 33.895 179.275 ;
        RECT 30.830 179.090 33.895 179.230 ;
        RECT 30.830 179.030 31.150 179.090 ;
        RECT 33.605 179.045 33.895 179.090 ;
        RECT 49.230 179.030 49.550 179.290 ;
        RECT 52.925 179.230 53.215 179.275 ;
        RECT 55.210 179.230 55.530 179.290 ;
        RECT 52.925 179.090 55.530 179.230 ;
        RECT 52.925 179.045 53.215 179.090 ;
        RECT 55.210 179.030 55.530 179.090 ;
        RECT 58.905 179.230 59.195 179.275 ;
        RECT 60.270 179.230 60.590 179.290 ;
        RECT 58.905 179.090 60.590 179.230 ;
        RECT 58.905 179.045 59.195 179.090 ;
        RECT 60.270 179.030 60.590 179.090 ;
        RECT 80.050 179.230 80.370 179.290 ;
        RECT 81.445 179.230 81.735 179.275 ;
        RECT 80.050 179.090 81.735 179.230 ;
        RECT 80.050 179.030 80.370 179.090 ;
        RECT 81.445 179.045 81.735 179.090 ;
        RECT 83.730 179.030 84.050 179.290 ;
        RECT 84.190 179.030 84.510 179.290 ;
        RECT 87.410 179.230 87.730 179.290 ;
        RECT 91.090 179.230 91.410 179.290 ;
        RECT 92.560 179.230 92.700 179.430 ;
        RECT 108.110 179.370 108.430 179.430 ;
        RECT 110.065 179.385 110.355 179.430 ;
        RECT 113.305 179.385 113.955 179.430 ;
        RECT 115.930 179.370 116.250 179.630 ;
        RECT 117.400 179.570 117.540 179.725 ;
        RECT 124.210 179.570 124.530 179.630 ;
        RECT 117.400 179.430 124.530 179.570 ;
        RECT 124.210 179.370 124.530 179.430 ;
        RECT 87.410 179.090 92.700 179.230 ;
        RECT 108.585 179.230 108.875 179.275 ;
        RECT 109.030 179.230 109.350 179.290 ;
        RECT 108.585 179.090 109.350 179.230 ;
        RECT 87.410 179.030 87.730 179.090 ;
        RECT 91.090 179.030 91.410 179.090 ;
        RECT 108.585 179.045 108.875 179.090 ;
        RECT 109.030 179.030 109.350 179.090 ;
        RECT 114.550 179.230 114.870 179.290 ;
        RECT 116.850 179.230 117.170 179.290 ;
        RECT 119.165 179.230 119.455 179.275 ;
        RECT 114.550 179.090 119.455 179.230 ;
        RECT 114.550 179.030 114.870 179.090 ;
        RECT 116.850 179.030 117.170 179.090 ;
        RECT 119.165 179.045 119.455 179.090 ;
        RECT 14.660 178.410 127.820 178.890 ;
        RECT 26.230 178.210 26.550 178.270 ;
        RECT 28.085 178.210 28.375 178.255 ;
        RECT 26.230 178.070 28.375 178.210 ;
        RECT 26.230 178.010 26.550 178.070 ;
        RECT 28.085 178.025 28.375 178.070 ;
        RECT 29.465 178.025 29.755 178.255 ;
        RECT 29.005 177.530 29.295 177.575 ;
        RECT 29.540 177.530 29.680 178.025 ;
        RECT 49.230 178.010 49.550 178.270 ;
        RECT 70.850 178.210 71.170 178.270 ;
        RECT 73.150 178.210 73.470 178.270 ;
        RECT 70.850 178.070 73.470 178.210 ;
        RECT 70.850 178.010 71.170 178.070 ;
        RECT 73.150 178.010 73.470 178.070 ;
        RECT 84.190 178.210 84.510 178.270 ;
        RECT 89.265 178.210 89.555 178.255 ;
        RECT 90.630 178.210 90.950 178.270 ;
        RECT 84.190 178.070 88.100 178.210 ;
        RECT 84.190 178.010 84.510 178.070 ;
        RECT 45.500 177.870 45.790 177.915 ;
        RECT 48.760 177.870 49.050 177.915 ;
        RECT 49.320 177.870 49.460 178.010 ;
        RECT 55.210 177.915 55.530 177.930 ;
        RECT 45.500 177.730 49.460 177.870 ;
        RECT 49.680 177.870 49.970 177.915 ;
        RECT 51.540 177.870 51.830 177.915 ;
        RECT 49.680 177.730 51.830 177.870 ;
        RECT 45.500 177.685 45.790 177.730 ;
        RECT 48.760 177.685 49.050 177.730 ;
        RECT 49.680 177.685 49.970 177.730 ;
        RECT 51.540 177.685 51.830 177.730 ;
        RECT 55.160 177.870 55.530 177.915 ;
        RECT 58.420 177.870 58.710 177.915 ;
        RECT 55.160 177.730 58.710 177.870 ;
        RECT 55.160 177.685 55.530 177.730 ;
        RECT 58.420 177.685 58.710 177.730 ;
        RECT 59.340 177.870 59.630 177.915 ;
        RECT 61.200 177.870 61.490 177.915 ;
        RECT 59.340 177.730 61.490 177.870 ;
        RECT 59.340 177.685 59.630 177.730 ;
        RECT 61.200 177.685 61.490 177.730 ;
        RECT 29.005 177.390 29.680 177.530 ;
        RECT 29.005 177.345 29.295 177.390 ;
        RECT 31.290 177.330 31.610 177.590 ;
        RECT 47.360 177.530 47.650 177.575 ;
        RECT 49.680 177.530 49.895 177.685 ;
        RECT 55.210 177.670 55.530 177.685 ;
        RECT 47.360 177.390 49.895 177.530 ;
        RECT 57.020 177.530 57.310 177.575 ;
        RECT 59.340 177.530 59.555 177.685 ;
        RECT 87.410 177.670 87.730 177.930 ;
        RECT 87.960 177.870 88.100 178.070 ;
        RECT 89.265 178.070 90.950 178.210 ;
        RECT 89.265 178.025 89.555 178.070 ;
        RECT 90.630 178.010 90.950 178.070 ;
        RECT 114.105 178.210 114.395 178.255 ;
        RECT 115.930 178.210 116.250 178.270 ;
        RECT 114.105 178.070 116.250 178.210 ;
        RECT 114.105 178.025 114.395 178.070 ;
        RECT 115.930 178.010 116.250 178.070 ;
        RECT 91.565 177.870 91.855 177.915 ;
        RECT 87.960 177.730 91.855 177.870 ;
        RECT 91.565 177.685 91.855 177.730 ;
        RECT 57.020 177.390 59.555 177.530 ;
        RECT 47.360 177.345 47.650 177.390 ;
        RECT 57.020 177.345 57.310 177.390 ;
        RECT 60.270 177.330 60.590 177.590 ;
        RECT 69.930 177.530 70.250 177.590 ;
        RECT 71.785 177.530 72.075 177.575 ;
        RECT 69.930 177.390 72.075 177.530 ;
        RECT 69.930 177.330 70.250 177.390 ;
        RECT 71.785 177.345 72.075 177.390 ;
        RECT 72.705 177.530 72.995 177.575 ;
        RECT 73.610 177.530 73.930 177.590 ;
        RECT 72.705 177.390 73.930 177.530 ;
        RECT 72.705 177.345 72.995 177.390 ;
        RECT 73.610 177.330 73.930 177.390 ;
        RECT 79.590 177.330 79.910 177.590 ;
        RECT 91.105 177.530 91.395 177.575 ;
        RECT 99.830 177.530 100.150 177.590 ;
        RECT 91.105 177.390 100.150 177.530 ;
        RECT 91.105 177.345 91.395 177.390 ;
        RECT 99.830 177.330 100.150 177.390 ;
        RECT 100.290 177.330 100.610 177.590 ;
        RECT 101.670 177.330 101.990 177.590 ;
        RECT 113.170 177.330 113.490 177.590 ;
        RECT 115.930 177.530 116.250 177.590 ;
        RECT 118.230 177.530 118.550 177.590 ;
        RECT 115.930 177.390 118.550 177.530 ;
        RECT 115.930 177.330 116.250 177.390 ;
        RECT 118.230 177.330 118.550 177.390 ;
        RECT 30.830 177.190 31.150 177.250 ;
        RECT 31.765 177.190 32.055 177.235 ;
        RECT 30.830 177.050 32.055 177.190 ;
        RECT 30.830 176.990 31.150 177.050 ;
        RECT 31.765 177.005 32.055 177.050 ;
        RECT 32.685 177.190 32.975 177.235 ;
        RECT 41.870 177.190 42.190 177.250 ;
        RECT 32.685 177.050 42.190 177.190 ;
        RECT 32.685 177.005 32.975 177.050 ;
        RECT 29.910 176.850 30.230 176.910 ;
        RECT 32.760 176.850 32.900 177.005 ;
        RECT 41.870 176.990 42.190 177.050 ;
        RECT 50.610 176.990 50.930 177.250 ;
        RECT 52.465 177.190 52.755 177.235 ;
        RECT 56.590 177.190 56.910 177.250 ;
        RECT 62.125 177.190 62.415 177.235 ;
        RECT 52.465 177.050 62.415 177.190 ;
        RECT 52.465 177.005 52.755 177.050 ;
        RECT 56.590 176.990 56.910 177.050 ;
        RECT 62.125 177.005 62.415 177.050 ;
        RECT 72.245 177.190 72.535 177.235 ;
        RECT 72.245 177.050 72.920 177.190 ;
        RECT 72.245 177.005 72.535 177.050 ;
        RECT 72.780 176.910 72.920 177.050 ;
        RECT 73.150 176.990 73.470 177.250 ;
        RECT 85.110 177.190 85.430 177.250 ;
        RECT 92.025 177.190 92.315 177.235 ;
        RECT 85.110 177.050 92.315 177.190 ;
        RECT 85.110 176.990 85.430 177.050 ;
        RECT 92.025 177.005 92.315 177.050 ;
        RECT 110.425 177.190 110.715 177.235 ;
        RECT 111.790 177.190 112.110 177.250 ;
        RECT 110.425 177.050 112.110 177.190 ;
        RECT 110.425 177.005 110.715 177.050 ;
        RECT 111.790 176.990 112.110 177.050 ;
        RECT 29.910 176.710 32.900 176.850 ;
        RECT 47.360 176.850 47.650 176.895 ;
        RECT 50.140 176.850 50.430 176.895 ;
        RECT 52.000 176.850 52.290 176.895 ;
        RECT 47.360 176.710 52.290 176.850 ;
        RECT 29.910 176.650 30.230 176.710 ;
        RECT 47.360 176.665 47.650 176.710 ;
        RECT 50.140 176.665 50.430 176.710 ;
        RECT 52.000 176.665 52.290 176.710 ;
        RECT 57.020 176.850 57.310 176.895 ;
        RECT 59.800 176.850 60.090 176.895 ;
        RECT 61.660 176.850 61.950 176.895 ;
        RECT 57.020 176.710 61.950 176.850 ;
        RECT 57.020 176.665 57.310 176.710 ;
        RECT 59.800 176.665 60.090 176.710 ;
        RECT 61.660 176.665 61.950 176.710 ;
        RECT 72.690 176.650 73.010 176.910 ;
        RECT 43.495 176.510 43.785 176.555 ;
        RECT 46.930 176.510 47.250 176.570 ;
        RECT 43.495 176.370 47.250 176.510 ;
        RECT 43.495 176.325 43.785 176.370 ;
        RECT 46.930 176.310 47.250 176.370 ;
        RECT 53.155 176.510 53.445 176.555 ;
        RECT 54.290 176.510 54.610 176.570 ;
        RECT 53.155 176.370 54.610 176.510 ;
        RECT 53.155 176.325 53.445 176.370 ;
        RECT 54.290 176.310 54.610 176.370 ;
        RECT 70.865 176.510 71.155 176.555 ;
        RECT 71.310 176.510 71.630 176.570 ;
        RECT 70.865 176.370 71.630 176.510 ;
        RECT 70.865 176.325 71.155 176.370 ;
        RECT 71.310 176.310 71.630 176.370 ;
        RECT 99.370 176.510 99.690 176.570 ;
        RECT 99.845 176.510 100.135 176.555 ;
        RECT 99.370 176.370 100.135 176.510 ;
        RECT 99.370 176.310 99.690 176.370 ;
        RECT 99.845 176.325 100.135 176.370 ;
        RECT 14.660 175.690 127.820 176.170 ;
        RECT 29.910 175.290 30.230 175.550 ;
        RECT 35.445 175.490 35.735 175.535 ;
        RECT 40.030 175.490 40.350 175.550 ;
        RECT 50.610 175.490 50.930 175.550 ;
        RECT 51.545 175.490 51.835 175.535 ;
        RECT 35.445 175.350 44.860 175.490 ;
        RECT 35.445 175.305 35.735 175.350 ;
        RECT 40.030 175.290 40.350 175.350 ;
        RECT 30.000 175.150 30.140 175.290 ;
        RECT 29.540 175.010 30.140 175.150 ;
        RECT 38.305 175.150 38.595 175.195 ;
        RECT 41.425 175.150 41.715 175.195 ;
        RECT 43.315 175.150 43.605 175.195 ;
        RECT 38.305 175.010 43.605 175.150 ;
        RECT 29.540 174.855 29.680 175.010 ;
        RECT 38.305 174.965 38.595 175.010 ;
        RECT 41.425 174.965 41.715 175.010 ;
        RECT 43.315 174.965 43.605 175.010 ;
        RECT 29.465 174.625 29.755 174.855 ;
        RECT 29.910 174.810 30.230 174.870 ;
        RECT 35.890 174.810 36.210 174.870 ;
        RECT 29.910 174.670 36.210 174.810 ;
        RECT 29.910 174.610 30.230 174.670 ;
        RECT 30.385 174.470 30.675 174.515 ;
        RECT 30.830 174.470 31.150 174.530 ;
        RECT 34.140 174.515 34.280 174.670 ;
        RECT 35.890 174.610 36.210 174.670 ;
        RECT 36.810 174.810 37.130 174.870 ;
        RECT 42.805 174.810 43.095 174.855 ;
        RECT 36.810 174.670 43.095 174.810 ;
        RECT 36.810 174.610 37.130 174.670 ;
        RECT 42.805 174.625 43.095 174.670 ;
        RECT 30.385 174.330 31.150 174.470 ;
        RECT 30.385 174.285 30.675 174.330 ;
        RECT 30.830 174.270 31.150 174.330 ;
        RECT 34.065 174.285 34.355 174.515 ;
        RECT 29.925 174.130 30.215 174.175 ;
        RECT 32.670 174.130 32.990 174.190 ;
        RECT 37.225 174.175 37.515 174.490 ;
        RECT 38.305 174.470 38.595 174.515 ;
        RECT 41.885 174.470 42.175 174.515 ;
        RECT 43.720 174.470 44.010 174.515 ;
        RECT 38.305 174.330 44.010 174.470 ;
        RECT 38.305 174.285 38.595 174.330 ;
        RECT 41.885 174.285 42.175 174.330 ;
        RECT 43.720 174.285 44.010 174.330 ;
        RECT 44.170 174.270 44.490 174.530 ;
        RECT 44.720 174.470 44.860 175.350 ;
        RECT 47.020 175.350 49.920 175.490 ;
        RECT 47.020 175.150 47.160 175.350 ;
        RECT 46.560 175.010 47.160 175.150 ;
        RECT 46.560 174.870 46.700 175.010 ;
        RECT 49.245 174.965 49.535 175.195 ;
        RECT 49.780 175.150 49.920 175.350 ;
        RECT 50.610 175.350 51.835 175.490 ;
        RECT 50.610 175.290 50.930 175.350 ;
        RECT 51.545 175.305 51.835 175.350 ;
        RECT 57.065 175.490 57.355 175.535 ;
        RECT 57.970 175.490 58.290 175.550 ;
        RECT 57.065 175.350 58.290 175.490 ;
        RECT 57.065 175.305 57.355 175.350 ;
        RECT 57.970 175.290 58.290 175.350 ;
        RECT 69.010 175.490 69.330 175.550 ;
        RECT 74.530 175.490 74.850 175.550 ;
        RECT 79.145 175.490 79.435 175.535 ;
        RECT 69.010 175.350 71.080 175.490 ;
        RECT 69.010 175.290 69.330 175.350 ;
        RECT 49.780 175.010 54.520 175.150 ;
        RECT 46.470 174.610 46.790 174.870 ;
        RECT 46.930 174.810 47.250 174.870 ;
        RECT 46.930 174.670 48.540 174.810 ;
        RECT 46.930 174.610 47.250 174.670 ;
        RECT 47.405 174.470 47.695 174.515 ;
        RECT 44.720 174.330 47.695 174.470 ;
        RECT 47.405 174.285 47.695 174.330 ;
        RECT 29.925 173.990 32.990 174.130 ;
        RECT 29.925 173.945 30.215 173.990 ;
        RECT 32.670 173.930 32.990 173.990 ;
        RECT 34.525 174.130 34.815 174.175 ;
        RECT 36.925 174.130 37.515 174.175 ;
        RECT 40.165 174.130 40.815 174.175 ;
        RECT 34.525 173.990 40.815 174.130 ;
        RECT 48.400 174.130 48.540 174.670 ;
        RECT 49.320 174.470 49.460 174.965 ;
        RECT 54.380 174.855 54.520 175.010 ;
        RECT 54.305 174.810 54.595 174.855 ;
        RECT 54.750 174.810 55.070 174.870 ;
        RECT 69.100 174.855 69.240 175.290 ;
        RECT 70.390 175.150 70.710 175.210 ;
        RECT 70.940 175.195 71.080 175.350 ;
        RECT 74.530 175.350 79.435 175.490 ;
        RECT 74.530 175.290 74.850 175.350 ;
        RECT 79.145 175.305 79.435 175.350 ;
        RECT 80.510 175.290 80.830 175.550 ;
        RECT 86.490 175.290 86.810 175.550 ;
        RECT 87.425 175.490 87.715 175.535 ;
        RECT 87.870 175.490 88.190 175.550 ;
        RECT 100.290 175.490 100.610 175.550 ;
        RECT 87.425 175.350 88.190 175.490 ;
        RECT 87.425 175.305 87.715 175.350 ;
        RECT 87.870 175.290 88.190 175.350 ;
        RECT 90.260 175.350 100.610 175.490 ;
        RECT 69.560 175.010 70.710 175.150 ;
        RECT 69.560 174.855 69.700 175.010 ;
        RECT 70.390 174.950 70.710 175.010 ;
        RECT 70.865 175.150 71.155 175.195 ;
        RECT 74.070 175.150 74.390 175.210 ;
        RECT 70.865 175.010 77.980 175.150 ;
        RECT 70.865 174.965 71.155 175.010 ;
        RECT 74.070 174.950 74.390 175.010 ;
        RECT 54.305 174.670 55.070 174.810 ;
        RECT 54.305 174.625 54.595 174.670 ;
        RECT 54.750 174.610 55.070 174.670 ;
        RECT 69.025 174.625 69.315 174.855 ;
        RECT 69.485 174.625 69.775 174.855 ;
        RECT 71.770 174.810 72.090 174.870 ;
        RECT 73.610 174.810 73.930 174.870 ;
        RECT 77.840 174.855 77.980 175.010 ;
        RECT 77.305 174.810 77.595 174.855 ;
        RECT 70.020 174.670 72.090 174.810 ;
        RECT 50.625 174.470 50.915 174.515 ;
        RECT 49.320 174.330 50.915 174.470 ;
        RECT 50.625 174.285 50.915 174.330 ;
        RECT 68.105 174.285 68.395 174.515 ;
        RECT 68.565 174.470 68.855 174.515 ;
        RECT 70.020 174.470 70.160 174.670 ;
        RECT 71.770 174.610 72.090 174.670 ;
        RECT 72.320 174.670 77.595 174.810 ;
        RECT 68.565 174.330 70.160 174.470 ;
        RECT 70.390 174.470 70.710 174.530 ;
        RECT 72.320 174.470 72.460 174.670 ;
        RECT 73.610 174.610 73.930 174.670 ;
        RECT 77.305 174.625 77.595 174.670 ;
        RECT 77.765 174.625 78.055 174.855 ;
        RECT 83.270 174.810 83.590 174.870 ;
        RECT 83.270 174.670 88.100 174.810 ;
        RECT 83.270 174.610 83.590 174.670 ;
        RECT 76.845 174.470 77.135 174.515 ;
        RECT 78.225 174.470 78.515 174.515 ;
        RECT 70.390 174.330 72.460 174.470 ;
        RECT 72.780 174.330 77.135 174.470 ;
        RECT 68.565 174.285 68.855 174.330 ;
        RECT 49.690 174.130 50.010 174.190 ;
        RECT 55.225 174.130 55.515 174.175 ;
        RECT 48.400 173.990 55.515 174.130 ;
        RECT 34.525 173.945 34.815 173.990 ;
        RECT 36.925 173.945 37.215 173.990 ;
        RECT 40.165 173.945 40.815 173.990 ;
        RECT 49.690 173.930 50.010 173.990 ;
        RECT 55.225 173.945 55.515 173.990 ;
        RECT 67.170 173.930 67.490 174.190 ;
        RECT 68.180 174.130 68.320 174.285 ;
        RECT 70.390 174.270 70.710 174.330 ;
        RECT 72.780 174.190 72.920 174.330 ;
        RECT 76.845 174.285 77.135 174.330 ;
        RECT 77.380 174.330 78.515 174.470 ;
        RECT 70.865 174.130 71.155 174.175 ;
        RECT 72.690 174.130 73.010 174.190 ;
        RECT 68.180 173.990 73.010 174.130 ;
        RECT 70.865 173.945 71.155 173.990 ;
        RECT 72.690 173.930 73.010 173.990 ;
        RECT 74.545 174.130 74.835 174.175 ;
        RECT 75.910 174.130 76.230 174.190 ;
        RECT 74.545 173.990 76.230 174.130 ;
        RECT 74.545 173.945 74.835 173.990 ;
        RECT 75.910 173.930 76.230 173.990 ;
        RECT 32.225 173.790 32.515 173.835 ;
        RECT 33.590 173.790 33.910 173.850 ;
        RECT 32.225 173.650 33.910 173.790 ;
        RECT 32.225 173.605 32.515 173.650 ;
        RECT 33.590 173.590 33.910 173.650 ;
        RECT 54.290 173.790 54.610 173.850 ;
        RECT 54.765 173.790 55.055 173.835 ;
        RECT 54.290 173.650 55.055 173.790 ;
        RECT 54.290 173.590 54.610 173.650 ;
        RECT 54.765 173.605 55.055 173.650 ;
        RECT 71.770 173.790 72.090 173.850 ;
        RECT 73.150 173.790 73.470 173.850 ;
        RECT 77.380 173.790 77.520 174.330 ;
        RECT 78.225 174.285 78.515 174.330 ;
        RECT 83.730 174.470 84.050 174.530 ;
        RECT 87.960 174.515 88.100 174.670 ;
        RECT 85.585 174.470 85.875 174.515 ;
        RECT 83.730 174.330 85.875 174.470 ;
        RECT 83.730 174.270 84.050 174.330 ;
        RECT 85.585 174.285 85.875 174.330 ;
        RECT 87.885 174.470 88.175 174.515 ;
        RECT 90.260 174.470 90.400 175.350 ;
        RECT 100.290 175.290 100.610 175.350 ;
        RECT 101.210 175.290 101.530 175.550 ;
        RECT 93.355 175.150 93.645 175.195 ;
        RECT 95.245 175.150 95.535 175.195 ;
        RECT 98.365 175.150 98.655 175.195 ;
        RECT 93.355 175.010 98.655 175.150 ;
        RECT 93.355 174.965 93.645 175.010 ;
        RECT 95.245 174.965 95.535 175.010 ;
        RECT 98.365 174.965 98.655 175.010 ;
        RECT 113.630 175.150 113.950 175.210 ;
        RECT 119.165 175.150 119.455 175.195 ;
        RECT 113.630 175.010 118.000 175.150 ;
        RECT 113.630 174.950 113.950 175.010 ;
        RECT 115.930 174.610 116.250 174.870 ;
        RECT 87.885 174.330 90.400 174.470 ;
        RECT 91.090 174.470 91.410 174.530 ;
        RECT 92.485 174.470 92.775 174.515 ;
        RECT 91.090 174.330 92.775 174.470 ;
        RECT 87.885 174.285 88.175 174.330 ;
        RECT 91.090 174.270 91.410 174.330 ;
        RECT 92.485 174.285 92.775 174.330 ;
        RECT 92.950 174.470 93.240 174.515 ;
        RECT 94.785 174.470 95.075 174.515 ;
        RECT 98.365 174.470 98.655 174.515 ;
        RECT 92.950 174.330 98.655 174.470 ;
        RECT 92.950 174.285 93.240 174.330 ;
        RECT 94.785 174.285 95.075 174.330 ;
        RECT 98.365 174.285 98.655 174.330 ;
        RECT 99.370 174.490 99.690 174.530 ;
        RECT 99.370 174.270 99.735 174.490 ;
        RECT 111.790 174.270 112.110 174.530 ;
        RECT 117.310 174.270 117.630 174.530 ;
        RECT 117.860 174.470 118.000 175.010 ;
        RECT 119.165 175.010 122.140 175.150 ;
        RECT 119.165 174.965 119.455 175.010 ;
        RECT 118.690 174.810 119.010 174.870 ;
        RECT 120.085 174.810 120.375 174.855 ;
        RECT 118.690 174.670 120.375 174.810 ;
        RECT 118.690 174.610 119.010 174.670 ;
        RECT 120.085 174.625 120.375 174.670 ;
        RECT 122.000 174.515 122.140 175.010 ;
        RECT 135.635 174.550 136.775 223.880 ;
        RECT 138.130 223.810 139.580 225.110 ;
        RECT 143.180 223.840 144.630 225.140 ;
        RECT 119.625 174.470 119.915 174.515 ;
        RECT 117.860 174.330 119.915 174.470 ;
        RECT 119.625 174.285 119.915 174.330 ;
        RECT 121.925 174.285 122.215 174.515 ;
        RECT 77.750 174.130 78.070 174.190 ;
        RECT 80.065 174.130 80.355 174.175 ;
        RECT 77.750 173.990 80.355 174.130 ;
        RECT 77.750 173.930 78.070 173.990 ;
        RECT 80.065 173.945 80.355 173.990 ;
        RECT 93.865 174.130 94.155 174.175 ;
        RECT 94.310 174.130 94.630 174.190 ;
        RECT 99.445 174.175 99.735 174.270 ;
        RECT 93.865 173.990 94.630 174.130 ;
        RECT 93.865 173.945 94.155 173.990 ;
        RECT 94.310 173.930 94.630 173.990 ;
        RECT 96.145 174.130 96.795 174.175 ;
        RECT 99.445 174.130 100.035 174.175 ;
        RECT 96.145 173.990 100.035 174.130 ;
        RECT 111.880 174.130 112.020 174.270 ;
        RECT 124.210 174.130 124.530 174.190 ;
        RECT 111.880 173.990 124.530 174.130 ;
        RECT 96.145 173.945 96.795 173.990 ;
        RECT 99.745 173.945 100.035 173.990 ;
        RECT 124.210 173.930 124.530 173.990 ;
        RECT 71.770 173.650 77.520 173.790 ;
        RECT 71.770 173.590 72.090 173.650 ;
        RECT 73.150 173.590 73.470 173.650 ;
        RECT 116.850 173.590 117.170 173.850 ;
        RECT 122.830 173.590 123.150 173.850 ;
        RECT 14.660 172.970 127.820 173.450 ;
        RECT 135.580 173.430 136.830 174.550 ;
        RECT 135.635 173.420 136.775 173.430 ;
        RECT 32.685 172.770 32.975 172.815 ;
        RECT 30.920 172.630 32.975 172.770 ;
        RECT 30.920 172.475 31.060 172.630 ;
        RECT 32.685 172.585 32.975 172.630 ;
        RECT 36.810 172.570 37.130 172.830 ;
        RECT 37.745 172.585 38.035 172.815 ;
        RECT 22.565 172.430 22.855 172.475 ;
        RECT 24.965 172.430 25.255 172.475 ;
        RECT 28.205 172.430 28.855 172.475 ;
        RECT 22.565 172.290 28.855 172.430 ;
        RECT 22.565 172.245 22.855 172.290 ;
        RECT 24.965 172.245 25.555 172.290 ;
        RECT 28.205 172.245 28.855 172.290 ;
        RECT 30.845 172.245 31.135 172.475 ;
        RECT 22.105 172.090 22.395 172.135 ;
        RECT 22.105 171.950 22.780 172.090 ;
        RECT 22.105 171.905 22.395 171.950 ;
        RECT 22.640 171.810 22.780 171.950 ;
        RECT 25.265 171.930 25.555 172.245 ;
        RECT 26.345 172.090 26.635 172.135 ;
        RECT 29.925 172.090 30.215 172.135 ;
        RECT 31.760 172.090 32.050 172.135 ;
        RECT 26.345 171.950 32.050 172.090 ;
        RECT 26.345 171.905 26.635 171.950 ;
        RECT 29.925 171.905 30.215 171.950 ;
        RECT 31.760 171.905 32.050 171.950 ;
        RECT 33.590 171.890 33.910 172.150 ;
        RECT 35.905 172.090 36.195 172.135 ;
        RECT 37.820 172.090 37.960 172.585 ;
        RECT 40.030 172.570 40.350 172.830 ;
        RECT 44.170 172.570 44.490 172.830 ;
        RECT 54.750 172.770 55.070 172.830 ;
        RECT 57.525 172.770 57.815 172.815 ;
        RECT 54.750 172.630 57.815 172.770 ;
        RECT 54.750 172.570 55.070 172.630 ;
        RECT 57.525 172.585 57.815 172.630 ;
        RECT 64.870 172.770 65.190 172.830 ;
        RECT 97.990 172.770 98.310 172.830 ;
        RECT 64.870 172.630 77.980 172.770 ;
        RECT 64.870 172.570 65.190 172.630 ;
        RECT 44.260 172.430 44.400 172.570 ;
        RECT 53.385 172.430 53.675 172.475 ;
        RECT 56.590 172.430 56.910 172.490 ;
        RECT 76.370 172.430 76.690 172.490 ;
        RECT 44.260 172.290 56.910 172.430 ;
        RECT 53.385 172.245 53.675 172.290 ;
        RECT 56.590 172.230 56.910 172.290 ;
        RECT 57.140 172.290 76.690 172.430 ;
        RECT 77.840 172.430 77.980 172.630 ;
        RECT 81.060 172.630 98.310 172.770 ;
        RECT 81.060 172.430 81.200 172.630 ;
        RECT 97.990 172.570 98.310 172.630 ;
        RECT 98.465 172.770 98.755 172.815 ;
        RECT 101.210 172.770 101.530 172.830 ;
        RECT 98.465 172.630 101.530 172.770 ;
        RECT 98.465 172.585 98.755 172.630 ;
        RECT 101.210 172.570 101.530 172.630 ;
        RECT 102.145 172.585 102.435 172.815 ;
        RECT 102.590 172.770 102.910 172.830 ;
        RECT 119.610 172.770 119.930 172.830 ;
        RECT 102.590 172.630 119.930 172.770 ;
        RECT 84.650 172.475 84.970 172.490 ;
        RECT 77.840 172.290 81.200 172.430 ;
        RECT 81.380 172.430 81.670 172.475 ;
        RECT 84.640 172.430 84.970 172.475 ;
        RECT 81.380 172.290 84.970 172.430 ;
        RECT 35.905 171.950 37.960 172.090 ;
        RECT 39.585 172.090 39.875 172.135 ;
        RECT 43.710 172.090 44.030 172.150 ;
        RECT 39.585 171.950 44.030 172.090 ;
        RECT 35.905 171.905 36.195 171.950 ;
        RECT 39.585 171.905 39.875 171.950 ;
        RECT 22.550 171.550 22.870 171.810 ;
        RECT 30.370 171.750 30.690 171.810 ;
        RECT 32.225 171.750 32.515 171.795 ;
        RECT 30.370 171.610 32.515 171.750 ;
        RECT 30.370 171.550 30.690 171.610 ;
        RECT 32.225 171.565 32.515 171.610 ;
        RECT 32.670 171.750 32.990 171.810 ;
        RECT 39.660 171.750 39.800 171.905 ;
        RECT 43.710 171.890 44.030 171.950 ;
        RECT 50.610 171.890 50.930 172.150 ;
        RECT 32.670 171.610 39.800 171.750 ;
        RECT 40.965 171.750 41.255 171.795 ;
        RECT 41.870 171.750 42.190 171.810 ;
        RECT 46.470 171.750 46.790 171.810 ;
        RECT 40.965 171.610 46.790 171.750 ;
        RECT 32.670 171.550 32.990 171.610 ;
        RECT 40.965 171.565 41.255 171.610 ;
        RECT 41.870 171.550 42.190 171.610 ;
        RECT 46.470 171.550 46.790 171.610 ;
        RECT 26.345 171.410 26.635 171.455 ;
        RECT 29.465 171.410 29.755 171.455 ;
        RECT 31.355 171.410 31.645 171.455 ;
        RECT 26.345 171.270 31.645 171.410 ;
        RECT 26.345 171.225 26.635 171.270 ;
        RECT 29.465 171.225 29.755 171.270 ;
        RECT 31.355 171.225 31.645 171.270 ;
        RECT 23.485 171.070 23.775 171.115 ;
        RECT 32.760 171.070 32.900 171.550 ;
        RECT 36.350 171.410 36.670 171.470 ;
        RECT 57.140 171.410 57.280 172.290 ;
        RECT 76.370 172.230 76.690 172.290 ;
        RECT 81.380 172.245 81.670 172.290 ;
        RECT 84.640 172.245 84.970 172.290 ;
        RECT 84.650 172.230 84.970 172.245 ;
        RECT 85.560 172.430 85.850 172.475 ;
        RECT 87.420 172.430 87.710 172.475 ;
        RECT 85.560 172.290 87.710 172.430 ;
        RECT 85.560 172.245 85.850 172.290 ;
        RECT 87.420 172.245 87.710 172.290 ;
        RECT 94.310 172.430 94.630 172.490 ;
        RECT 102.220 172.430 102.360 172.585 ;
        RECT 102.590 172.570 102.910 172.630 ;
        RECT 119.610 172.570 119.930 172.630 ;
        RECT 117.310 172.430 117.630 172.490 ;
        RECT 94.310 172.290 102.360 172.430 ;
        RECT 111.420 172.290 117.630 172.430 ;
        RECT 58.905 171.905 59.195 172.135 ;
        RECT 65.805 172.090 66.095 172.135 ;
        RECT 66.265 172.090 66.555 172.135 ;
        RECT 67.170 172.090 67.490 172.150 ;
        RECT 68.550 172.090 68.870 172.150 ;
        RECT 65.805 171.950 68.870 172.090 ;
        RECT 65.805 171.905 66.095 171.950 ;
        RECT 66.265 171.905 66.555 171.950 ;
        RECT 58.980 171.750 59.120 171.905 ;
        RECT 67.170 171.890 67.490 171.950 ;
        RECT 68.550 171.890 68.870 171.950 ;
        RECT 69.930 172.090 70.250 172.150 ;
        RECT 70.405 172.090 70.695 172.135 ;
        RECT 69.930 171.950 70.695 172.090 ;
        RECT 69.930 171.890 70.250 171.950 ;
        RECT 70.405 171.905 70.695 171.950 ;
        RECT 72.690 171.890 73.010 172.150 ;
        RECT 73.150 171.890 73.470 172.150 ;
        RECT 73.610 171.890 73.930 172.150 ;
        RECT 74.070 171.890 74.390 172.150 ;
        RECT 76.845 171.905 77.135 172.135 ;
        RECT 83.240 172.090 83.530 172.135 ;
        RECT 85.560 172.090 85.775 172.245 ;
        RECT 94.310 172.230 94.630 172.290 ;
        RECT 83.240 171.950 85.775 172.090 ;
        RECT 88.345 172.090 88.635 172.135 ;
        RECT 91.090 172.090 91.410 172.150 ;
        RECT 93.850 172.090 94.170 172.150 ;
        RECT 88.345 171.950 94.170 172.090 ;
        RECT 83.240 171.905 83.530 171.950 ;
        RECT 88.345 171.905 88.635 171.950 ;
        RECT 69.470 171.750 69.790 171.810 ;
        RECT 76.920 171.750 77.060 171.905 ;
        RECT 91.090 171.890 91.410 171.950 ;
        RECT 93.850 171.890 94.170 171.950 ;
        RECT 98.925 171.905 99.215 172.135 ;
        RECT 103.065 172.090 103.355 172.135 ;
        RECT 100.840 171.950 103.355 172.090 ;
        RECT 58.980 171.610 77.060 171.750 ;
        RECT 78.225 171.750 78.515 171.795 ;
        RECT 85.110 171.750 85.430 171.810 ;
        RECT 78.225 171.610 85.430 171.750 ;
        RECT 69.470 171.550 69.790 171.610 ;
        RECT 78.225 171.565 78.515 171.610 ;
        RECT 85.110 171.550 85.430 171.610 ;
        RECT 86.505 171.750 86.795 171.795 ;
        RECT 89.250 171.750 89.570 171.810 ;
        RECT 86.505 171.610 89.570 171.750 ;
        RECT 86.505 171.565 86.795 171.610 ;
        RECT 89.250 171.550 89.570 171.610 ;
        RECT 97.530 171.550 97.850 171.810 ;
        RECT 36.350 171.270 57.280 171.410 ;
        RECT 83.240 171.410 83.530 171.455 ;
        RECT 86.020 171.410 86.310 171.455 ;
        RECT 87.880 171.410 88.170 171.455 ;
        RECT 83.240 171.270 88.170 171.410 ;
        RECT 36.350 171.210 36.670 171.270 ;
        RECT 83.240 171.225 83.530 171.270 ;
        RECT 86.020 171.225 86.310 171.270 ;
        RECT 87.880 171.225 88.170 171.270 ;
        RECT 23.485 170.930 32.900 171.070 ;
        RECT 23.485 170.885 23.775 170.930 ;
        RECT 67.170 170.870 67.490 171.130 ;
        RECT 70.390 171.070 70.710 171.130 ;
        RECT 70.865 171.070 71.155 171.115 ;
        RECT 70.390 170.930 71.155 171.070 ;
        RECT 70.390 170.870 70.710 170.930 ;
        RECT 70.865 170.885 71.155 170.930 ;
        RECT 71.770 170.870 72.090 171.130 ;
        RECT 79.130 171.115 79.450 171.130 ;
        RECT 79.130 171.070 79.665 171.115 ;
        RECT 84.190 171.070 84.510 171.130 ;
        RECT 99.000 171.070 99.140 171.905 ;
        RECT 100.840 171.455 100.980 171.950 ;
        RECT 103.065 171.905 103.355 171.950 ;
        RECT 105.810 172.090 106.130 172.150 ;
        RECT 111.420 172.135 111.560 172.290 ;
        RECT 117.310 172.230 117.630 172.290 ;
        RECT 118.345 172.430 118.635 172.475 ;
        RECT 121.585 172.430 122.235 172.475 ;
        RECT 118.345 172.290 122.235 172.430 ;
        RECT 118.345 172.245 118.935 172.290 ;
        RECT 121.585 172.245 122.235 172.290 ;
        RECT 122.830 172.430 123.150 172.490 ;
        RECT 124.225 172.430 124.515 172.475 ;
        RECT 122.830 172.290 124.515 172.430 ;
        RECT 118.645 172.150 118.935 172.245 ;
        RECT 122.830 172.230 123.150 172.290 ;
        RECT 124.225 172.245 124.515 172.290 ;
        RECT 134.290 172.170 136.690 172.190 ;
        RECT 110.425 172.090 110.715 172.135 ;
        RECT 105.810 171.950 110.715 172.090 ;
        RECT 105.810 171.890 106.130 171.950 ;
        RECT 110.425 171.905 110.715 171.950 ;
        RECT 110.885 171.905 111.175 172.135 ;
        RECT 111.345 171.905 111.635 172.135 ;
        RECT 109.950 171.750 110.270 171.810 ;
        RECT 110.960 171.750 111.100 171.905 ;
        RECT 112.250 171.890 112.570 172.150 ;
        RECT 114.090 172.090 114.410 172.150 ;
        RECT 115.485 172.090 115.775 172.135 ;
        RECT 114.090 171.950 115.775 172.090 ;
        RECT 114.090 171.890 114.410 171.950 ;
        RECT 115.485 171.905 115.775 171.950 ;
        RECT 118.645 171.930 119.010 172.150 ;
        RECT 118.690 171.890 119.010 171.930 ;
        RECT 119.725 172.090 120.015 172.135 ;
        RECT 123.305 172.090 123.595 172.135 ;
        RECT 125.140 172.090 125.430 172.135 ;
        RECT 119.725 171.950 125.430 172.090 ;
        RECT 119.725 171.905 120.015 171.950 ;
        RECT 123.305 171.905 123.595 171.950 ;
        RECT 125.140 171.905 125.430 171.950 ;
        RECT 133.920 171.930 136.690 172.170 ;
        RECT 138.330 171.930 139.470 223.810 ;
        RECT 109.950 171.610 111.100 171.750 ;
        RECT 124.210 171.750 124.530 171.810 ;
        RECT 125.605 171.750 125.895 171.795 ;
        RECT 124.210 171.610 125.895 171.750 ;
        RECT 109.950 171.550 110.270 171.610 ;
        RECT 124.210 171.550 124.530 171.610 ;
        RECT 125.605 171.565 125.895 171.610 ;
        RECT 100.765 171.225 101.055 171.455 ;
        RECT 110.410 171.410 110.730 171.470 ;
        RECT 116.850 171.410 117.170 171.470 ;
        RECT 110.410 171.270 117.170 171.410 ;
        RECT 110.410 171.210 110.730 171.270 ;
        RECT 116.850 171.210 117.170 171.270 ;
        RECT 119.725 171.410 120.015 171.455 ;
        RECT 122.845 171.410 123.135 171.455 ;
        RECT 124.735 171.410 125.025 171.455 ;
        RECT 119.725 171.270 125.025 171.410 ;
        RECT 119.725 171.225 120.015 171.270 ;
        RECT 122.845 171.225 123.135 171.270 ;
        RECT 124.735 171.225 125.025 171.270 ;
        RECT 79.130 170.930 99.140 171.070 ;
        RECT 109.045 171.070 109.335 171.115 ;
        RECT 109.490 171.070 109.810 171.130 ;
        RECT 109.045 170.930 109.810 171.070 ;
        RECT 79.130 170.885 79.665 170.930 ;
        RECT 79.130 170.870 79.450 170.885 ;
        RECT 84.190 170.870 84.510 170.930 ;
        RECT 109.045 170.885 109.335 170.930 ;
        RECT 109.490 170.870 109.810 170.930 ;
        RECT 116.390 170.870 116.710 171.130 ;
        RECT 133.920 170.790 139.470 171.930 ;
        RECT 14.660 170.250 127.820 170.730 ;
        RECT 133.920 170.600 136.690 170.790 ;
        RECT 133.920 170.590 134.760 170.600 ;
        RECT 41.870 170.050 42.190 170.110 ;
        RECT 57.050 170.050 57.370 170.110 ;
        RECT 41.870 169.910 57.370 170.050 ;
        RECT 41.870 169.850 42.190 169.910 ;
        RECT 57.050 169.850 57.370 169.910 ;
        RECT 63.045 170.050 63.335 170.095 ;
        RECT 63.950 170.050 64.270 170.110 ;
        RECT 63.045 169.910 64.270 170.050 ;
        RECT 63.045 169.865 63.335 169.910 ;
        RECT 63.950 169.850 64.270 169.910 ;
        RECT 69.470 169.850 69.790 170.110 ;
        RECT 75.005 170.050 75.295 170.095 ;
        RECT 76.370 170.050 76.690 170.110 ;
        RECT 75.005 169.910 76.690 170.050 ;
        RECT 75.005 169.865 75.295 169.910 ;
        RECT 76.370 169.850 76.690 169.910 ;
        RECT 84.650 170.050 84.970 170.110 ;
        RECT 88.345 170.050 88.635 170.095 ;
        RECT 84.650 169.910 88.635 170.050 ;
        RECT 84.650 169.850 84.970 169.910 ;
        RECT 88.345 169.865 88.635 169.910 ;
        RECT 89.250 169.850 89.570 170.110 ;
        RECT 102.590 170.050 102.910 170.110 ;
        RECT 97.160 169.910 102.910 170.050 ;
        RECT 42.790 169.710 43.110 169.770 ;
        RECT 55.210 169.710 55.530 169.770 ;
        RECT 74.070 169.710 74.390 169.770 ;
        RECT 85.110 169.710 85.430 169.770 ;
        RECT 86.950 169.710 87.270 169.770 ;
        RECT 42.790 169.570 49.000 169.710 ;
        RECT 42.790 169.510 43.110 169.570 ;
        RECT 29.910 169.370 30.230 169.430 ;
        RECT 40.045 169.370 40.335 169.415 ;
        RECT 29.910 169.230 40.335 169.370 ;
        RECT 29.910 169.170 30.230 169.230 ;
        RECT 40.045 169.185 40.335 169.230 ;
        RECT 22.550 168.830 22.870 169.090 ;
        RECT 41.425 169.030 41.715 169.075 ;
        RECT 41.870 169.030 42.190 169.090 ;
        RECT 41.425 168.890 42.190 169.030 ;
        RECT 41.425 168.845 41.715 168.890 ;
        RECT 41.870 168.830 42.190 168.890 ;
        RECT 42.805 169.030 43.095 169.075 ;
        RECT 42.805 168.890 43.480 169.030 ;
        RECT 42.805 168.845 43.095 168.890 ;
        RECT 22.090 168.150 22.410 168.410 ;
        RECT 43.340 168.350 43.480 168.890 ;
        RECT 43.710 168.830 44.030 169.090 ;
        RECT 44.185 168.845 44.475 169.075 ;
        RECT 44.645 169.030 44.935 169.075 ;
        RECT 45.550 169.030 45.870 169.090 ;
        RECT 48.860 169.075 49.000 169.570 ;
        RECT 49.780 169.570 55.530 169.710 ;
        RECT 49.780 169.075 49.920 169.570 ;
        RECT 55.210 169.510 55.530 169.570 ;
        RECT 70.020 169.570 74.390 169.710 ;
        RECT 64.870 169.370 65.190 169.430 ;
        RECT 70.020 169.415 70.160 169.570 ;
        RECT 74.070 169.510 74.390 169.570 ;
        RECT 84.740 169.570 87.270 169.710 ;
        RECT 69.025 169.370 69.315 169.415 ;
        RECT 53.460 169.230 65.190 169.370 ;
        RECT 44.645 168.890 45.870 169.030 ;
        RECT 44.645 168.845 44.935 168.890 ;
        RECT 44.260 168.690 44.400 168.845 ;
        RECT 45.550 168.830 45.870 168.890 ;
        RECT 47.865 168.845 48.155 169.075 ;
        RECT 48.325 168.845 48.615 169.075 ;
        RECT 48.785 168.845 49.075 169.075 ;
        RECT 49.705 168.845 49.995 169.075 ;
        RECT 52.450 169.030 52.770 169.090 ;
        RECT 53.460 169.075 53.600 169.230 ;
        RECT 64.870 169.170 65.190 169.230 ;
        RECT 65.880 169.230 69.315 169.370 ;
        RECT 65.880 169.090 66.020 169.230 ;
        RECT 69.025 169.185 69.315 169.230 ;
        RECT 69.945 169.185 70.235 169.415 ;
        RECT 70.390 169.370 70.710 169.430 ;
        RECT 84.740 169.415 84.880 169.570 ;
        RECT 85.110 169.510 85.430 169.570 ;
        RECT 86.950 169.510 87.270 169.570 ;
        RECT 87.425 169.525 87.715 169.755 ;
        RECT 70.390 169.230 75.680 169.370 ;
        RECT 70.390 169.170 70.710 169.230 ;
        RECT 75.540 169.090 75.680 169.230 ;
        RECT 84.665 169.185 84.955 169.415 ;
        RECT 87.500 169.370 87.640 169.525 ;
        RECT 87.500 169.230 90.400 169.370 ;
        RECT 53.385 169.030 53.675 169.075 ;
        RECT 52.450 168.890 53.675 169.030 ;
        RECT 45.090 168.690 45.410 168.750 ;
        RECT 44.260 168.550 45.410 168.690 ;
        RECT 45.090 168.490 45.410 168.550 ;
        RECT 44.170 168.350 44.490 168.410 ;
        RECT 43.340 168.210 44.490 168.350 ;
        RECT 44.170 168.150 44.490 168.210 ;
        RECT 46.010 168.150 46.330 168.410 ;
        RECT 46.470 168.150 46.790 168.410 ;
        RECT 47.940 168.350 48.080 168.845 ;
        RECT 48.400 168.690 48.540 168.845 ;
        RECT 52.450 168.830 52.770 168.890 ;
        RECT 53.385 168.845 53.675 168.890 ;
        RECT 53.830 168.830 54.150 169.090 ;
        RECT 54.290 168.830 54.610 169.090 ;
        RECT 55.210 168.830 55.530 169.090 ;
        RECT 65.790 168.830 66.110 169.090 ;
        RECT 68.550 168.830 68.870 169.090 ;
        RECT 71.770 168.830 72.090 169.090 ;
        RECT 73.165 168.845 73.455 169.075 ;
        RECT 53.920 168.690 54.060 168.830 ;
        RECT 48.400 168.550 54.060 168.690 ;
        RECT 57.050 168.690 57.370 168.750 ;
        RECT 63.505 168.690 63.795 168.735 ;
        RECT 73.240 168.690 73.380 168.845 ;
        RECT 74.070 168.830 74.390 169.090 ;
        RECT 75.450 168.830 75.770 169.090 ;
        RECT 84.190 169.030 84.510 169.090 ;
        RECT 85.125 169.030 85.415 169.075 ;
        RECT 84.190 168.890 85.415 169.030 ;
        RECT 84.190 168.830 84.510 168.890 ;
        RECT 85.125 168.845 85.415 168.890 ;
        RECT 87.410 169.030 87.730 169.090 ;
        RECT 90.260 169.075 90.400 169.230 ;
        RECT 88.805 169.030 89.095 169.075 ;
        RECT 87.410 168.890 89.095 169.030 ;
        RECT 87.410 168.830 87.730 168.890 ;
        RECT 88.805 168.845 89.095 168.890 ;
        RECT 90.185 168.845 90.475 169.075 ;
        RECT 74.530 168.690 74.850 168.750 ;
        RECT 97.160 168.690 97.300 169.910 ;
        RECT 102.590 169.850 102.910 169.910 ;
        RECT 114.090 169.850 114.410 170.110 ;
        RECT 115.930 169.710 116.250 169.770 ;
        RECT 101.300 169.570 116.250 169.710 ;
        RECT 97.530 169.370 97.850 169.430 ;
        RECT 98.005 169.370 98.295 169.415 ;
        RECT 101.300 169.370 101.440 169.570 ;
        RECT 97.530 169.230 101.440 169.370 ;
        RECT 101.670 169.370 101.990 169.430 ;
        RECT 111.420 169.415 111.560 169.570 ;
        RECT 115.930 169.510 116.250 169.570 ;
        RECT 118.660 169.710 118.950 169.755 ;
        RECT 121.440 169.710 121.730 169.755 ;
        RECT 123.300 169.710 123.590 169.755 ;
        RECT 118.660 169.570 123.590 169.710 ;
        RECT 118.660 169.525 118.950 169.570 ;
        RECT 121.440 169.525 121.730 169.570 ;
        RECT 123.300 169.525 123.590 169.570 ;
        RECT 101.670 169.230 107.420 169.370 ;
        RECT 97.530 169.170 97.850 169.230 ;
        RECT 98.005 169.185 98.295 169.230 ;
        RECT 57.050 168.550 71.310 168.690 ;
        RECT 73.240 168.550 74.850 168.690 ;
        RECT 57.050 168.490 57.370 168.550 ;
        RECT 63.505 168.505 63.795 168.550 ;
        RECT 49.230 168.350 49.550 168.410 ;
        RECT 47.940 168.210 49.550 168.350 ;
        RECT 49.230 168.150 49.550 168.210 ;
        RECT 51.990 168.150 52.310 168.410 ;
        RECT 66.710 168.150 67.030 168.410 ;
        RECT 71.170 168.350 71.310 168.550 ;
        RECT 74.530 168.490 74.850 168.550 ;
        RECT 84.740 168.550 97.300 168.690 ;
        RECT 84.740 168.350 84.880 168.550 ;
        RECT 71.170 168.210 84.880 168.350 ;
        RECT 85.110 168.350 85.430 168.410 ;
        RECT 85.585 168.350 85.875 168.395 ;
        RECT 85.110 168.210 85.875 168.350 ;
        RECT 85.110 168.150 85.430 168.210 ;
        RECT 85.585 168.165 85.875 168.210 ;
        RECT 86.950 168.350 87.270 168.410 ;
        RECT 91.090 168.350 91.410 168.410 ;
        RECT 98.080 168.350 98.220 169.185 ;
        RECT 101.670 169.170 101.990 169.230 ;
        RECT 103.065 169.030 103.355 169.075 ;
        RECT 101.300 168.890 103.355 169.030 ;
        RECT 86.950 168.210 98.220 168.350 ;
        RECT 98.450 168.350 98.770 168.410 ;
        RECT 98.925 168.350 99.215 168.395 ;
        RECT 98.450 168.210 99.215 168.350 ;
        RECT 86.950 168.150 87.270 168.210 ;
        RECT 91.090 168.150 91.410 168.210 ;
        RECT 98.450 168.150 98.770 168.210 ;
        RECT 98.925 168.165 99.215 168.210 ;
        RECT 99.385 168.350 99.675 168.395 ;
        RECT 100.290 168.350 100.610 168.410 ;
        RECT 101.300 168.395 101.440 168.890 ;
        RECT 103.065 168.845 103.355 168.890 ;
        RECT 105.810 169.030 106.130 169.090 ;
        RECT 106.285 169.030 106.575 169.075 ;
        RECT 105.810 168.890 106.575 169.030 ;
        RECT 105.810 168.830 106.130 168.890 ;
        RECT 106.285 168.845 106.575 168.890 ;
        RECT 106.730 168.830 107.050 169.090 ;
        RECT 107.280 169.075 107.420 169.230 ;
        RECT 111.345 169.185 111.635 169.415 ;
        RECT 116.390 169.370 116.710 169.430 ;
        RECT 121.925 169.370 122.215 169.415 ;
        RECT 116.390 169.230 122.215 169.370 ;
        RECT 116.390 169.170 116.710 169.230 ;
        RECT 121.925 169.185 122.215 169.230 ;
        RECT 107.205 168.845 107.495 169.075 ;
        RECT 108.125 169.030 108.415 169.075 ;
        RECT 110.870 169.030 111.190 169.090 ;
        RECT 112.250 169.030 112.570 169.090 ;
        RECT 108.125 168.890 112.570 169.030 ;
        RECT 108.125 168.845 108.415 168.890 ;
        RECT 110.870 168.830 111.190 168.890 ;
        RECT 112.250 168.830 112.570 168.890 ;
        RECT 118.660 169.030 118.950 169.075 ;
        RECT 123.765 169.030 124.055 169.075 ;
        RECT 124.210 169.030 124.530 169.090 ;
        RECT 118.660 168.890 121.195 169.030 ;
        RECT 118.660 168.845 118.950 168.890 ;
        RECT 101.670 168.690 101.990 168.750 ;
        RECT 116.850 168.735 117.170 168.750 ;
        RECT 120.980 168.735 121.195 168.890 ;
        RECT 123.765 168.890 124.530 169.030 ;
        RECT 123.765 168.845 124.055 168.890 ;
        RECT 124.210 168.830 124.530 168.890 ;
        RECT 125.145 169.030 125.435 169.075 ;
        RECT 130.190 169.030 130.510 169.090 ;
        RECT 125.145 168.890 130.510 169.030 ;
        RECT 125.145 168.845 125.435 168.890 ;
        RECT 130.190 168.830 130.510 168.890 ;
        RECT 111.805 168.690 112.095 168.735 ;
        RECT 114.795 168.690 115.085 168.735 ;
        RECT 101.670 168.550 115.085 168.690 ;
        RECT 101.670 168.490 101.990 168.550 ;
        RECT 111.805 168.505 112.095 168.550 ;
        RECT 114.795 168.505 115.085 168.550 ;
        RECT 116.800 168.690 117.170 168.735 ;
        RECT 120.060 168.690 120.350 168.735 ;
        RECT 116.800 168.550 120.350 168.690 ;
        RECT 116.800 168.505 117.170 168.550 ;
        RECT 120.060 168.505 120.350 168.550 ;
        RECT 120.980 168.690 121.270 168.735 ;
        RECT 122.840 168.690 123.130 168.735 ;
        RECT 120.980 168.550 123.130 168.690 ;
        RECT 120.980 168.505 121.270 168.550 ;
        RECT 122.840 168.505 123.130 168.550 ;
        RECT 116.850 168.490 117.170 168.505 ;
        RECT 99.385 168.210 100.610 168.350 ;
        RECT 99.385 168.165 99.675 168.210 ;
        RECT 100.290 168.150 100.610 168.210 ;
        RECT 101.225 168.165 101.515 168.395 ;
        RECT 103.970 168.150 104.290 168.410 ;
        RECT 104.905 168.350 105.195 168.395 ;
        RECT 105.350 168.350 105.670 168.410 ;
        RECT 104.905 168.210 105.670 168.350 ;
        RECT 104.905 168.165 105.195 168.210 ;
        RECT 105.350 168.150 105.670 168.210 ;
        RECT 110.410 168.350 110.730 168.410 ;
        RECT 112.265 168.350 112.555 168.395 ;
        RECT 110.410 168.210 112.555 168.350 ;
        RECT 110.410 168.150 110.730 168.210 ;
        RECT 112.265 168.165 112.555 168.210 ;
        RECT 119.610 168.350 119.930 168.410 ;
        RECT 124.685 168.350 124.975 168.395 ;
        RECT 119.610 168.210 124.975 168.350 ;
        RECT 119.610 168.150 119.930 168.210 ;
        RECT 124.685 168.165 124.975 168.210 ;
        RECT 14.660 167.530 127.820 168.010 ;
        RECT 52.910 167.330 53.230 167.390 ;
        RECT 66.710 167.330 67.030 167.390 ;
        RECT 80.510 167.330 80.830 167.390 ;
        RECT 87.410 167.330 87.730 167.390 ;
        RECT 97.990 167.330 98.310 167.390 ;
        RECT 105.810 167.330 106.130 167.390 ;
        RECT 108.570 167.330 108.890 167.390 ;
        RECT 52.910 167.190 80.830 167.330 ;
        RECT 52.910 167.130 53.230 167.190 ;
        RECT 66.710 167.130 67.030 167.190 ;
        RECT 19.445 166.990 19.735 167.035 ;
        RECT 22.090 166.990 22.410 167.050 ;
        RECT 22.685 166.990 23.335 167.035 ;
        RECT 19.445 166.850 23.335 166.990 ;
        RECT 19.445 166.805 20.035 166.850 ;
        RECT 19.745 166.490 20.035 166.805 ;
        RECT 22.090 166.790 22.410 166.850 ;
        RECT 22.685 166.805 23.335 166.850 ;
        RECT 36.350 166.790 36.670 167.050 ;
        RECT 44.170 166.990 44.490 167.050 ;
        RECT 55.210 166.990 55.530 167.050 ;
        RECT 59.350 166.990 59.670 167.050 ;
        RECT 43.800 166.850 47.620 166.990 ;
        RECT 20.825 166.650 21.115 166.695 ;
        RECT 24.405 166.650 24.695 166.695 ;
        RECT 26.240 166.650 26.530 166.695 ;
        RECT 20.825 166.510 26.530 166.650 ;
        RECT 20.825 166.465 21.115 166.510 ;
        RECT 24.405 166.465 24.695 166.510 ;
        RECT 26.240 166.465 26.530 166.510 ;
        RECT 26.705 166.650 26.995 166.695 ;
        RECT 28.530 166.650 28.850 166.710 ;
        RECT 30.370 166.650 30.690 166.710 ;
        RECT 26.705 166.510 30.690 166.650 ;
        RECT 26.705 166.465 26.995 166.510 ;
        RECT 28.530 166.450 28.850 166.510 ;
        RECT 30.370 166.450 30.690 166.510 ;
        RECT 37.730 166.450 38.050 166.710 ;
        RECT 40.045 166.465 40.335 166.695 ;
        RECT 40.490 166.650 40.810 166.710 ;
        RECT 40.965 166.650 41.255 166.695 ;
        RECT 40.490 166.510 41.255 166.650 ;
        RECT 25.310 166.110 25.630 166.370 ;
        RECT 40.120 166.310 40.260 166.465 ;
        RECT 40.490 166.450 40.810 166.510 ;
        RECT 40.965 166.465 41.255 166.510 ;
        RECT 41.410 166.450 41.730 166.710 ;
        RECT 43.800 166.695 43.940 166.850 ;
        RECT 44.170 166.790 44.490 166.850 ;
        RECT 41.885 166.650 42.175 166.695 ;
        RECT 41.885 166.510 42.560 166.650 ;
        RECT 41.885 166.465 42.175 166.510 ;
        RECT 40.120 166.170 41.180 166.310 ;
        RECT 41.040 166.030 41.180 166.170 ;
        RECT 20.825 165.970 21.115 166.015 ;
        RECT 23.945 165.970 24.235 166.015 ;
        RECT 25.835 165.970 26.125 166.015 ;
        RECT 20.825 165.830 26.125 165.970 ;
        RECT 20.825 165.785 21.115 165.830 ;
        RECT 23.945 165.785 24.235 165.830 ;
        RECT 25.835 165.785 26.125 165.830 ;
        RECT 30.830 165.970 31.150 166.030 ;
        RECT 30.830 165.830 40.720 165.970 ;
        RECT 30.830 165.770 31.150 165.830 ;
        RECT 17.950 165.430 18.270 165.690 ;
        RECT 21.630 165.630 21.950 165.690 ;
        RECT 35.890 165.630 36.210 165.690 ;
        RECT 21.630 165.490 36.210 165.630 ;
        RECT 21.630 165.430 21.950 165.490 ;
        RECT 35.890 165.430 36.210 165.490 ;
        RECT 38.650 165.430 38.970 165.690 ;
        RECT 40.580 165.630 40.720 165.830 ;
        RECT 40.950 165.770 41.270 166.030 ;
        RECT 42.420 165.970 42.560 166.510 ;
        RECT 43.725 166.465 44.015 166.695 ;
        RECT 44.645 166.465 44.935 166.695 ;
        RECT 43.250 166.310 43.570 166.370 ;
        RECT 44.720 166.310 44.860 166.465 ;
        RECT 45.090 166.450 45.410 166.710 ;
        RECT 45.550 166.650 45.870 166.710 ;
        RECT 46.930 166.650 47.250 166.710 ;
        RECT 47.480 166.695 47.620 166.850 ;
        RECT 48.860 166.850 53.140 166.990 ;
        RECT 48.860 166.695 49.000 166.850 ;
        RECT 45.550 166.510 47.250 166.650 ;
        RECT 45.550 166.450 45.870 166.510 ;
        RECT 46.930 166.450 47.250 166.510 ;
        RECT 47.405 166.465 47.695 166.695 ;
        RECT 48.325 166.465 48.615 166.695 ;
        RECT 48.785 166.465 49.075 166.695 ;
        RECT 49.230 166.650 49.550 166.710 ;
        RECT 52.450 166.650 52.770 166.710 ;
        RECT 53.000 166.695 53.140 166.850 ;
        RECT 54.380 166.850 59.670 166.990 ;
        RECT 49.230 166.510 52.770 166.650 ;
        RECT 43.250 166.170 44.860 166.310 ;
        RECT 43.250 166.110 43.570 166.170 ;
        RECT 45.640 165.970 45.780 166.450 ;
        RECT 42.420 165.830 45.780 165.970 ;
        RECT 47.480 165.970 47.620 166.465 ;
        RECT 48.400 166.310 48.540 166.465 ;
        RECT 49.230 166.450 49.550 166.510 ;
        RECT 52.450 166.450 52.770 166.510 ;
        RECT 52.925 166.465 53.215 166.695 ;
        RECT 49.690 166.310 50.010 166.370 ;
        RECT 48.400 166.170 50.010 166.310 ;
        RECT 49.690 166.110 50.010 166.170 ;
        RECT 50.625 166.310 50.915 166.355 ;
        RECT 51.530 166.310 51.850 166.370 ;
        RECT 50.625 166.170 51.850 166.310 ;
        RECT 53.000 166.310 53.140 166.465 ;
        RECT 53.370 166.450 53.690 166.710 ;
        RECT 54.380 166.695 54.520 166.850 ;
        RECT 55.210 166.790 55.530 166.850 ;
        RECT 59.350 166.790 59.670 166.850 ;
        RECT 54.305 166.465 54.595 166.695 ;
        RECT 55.670 166.450 55.990 166.710 ;
        RECT 57.050 166.450 57.370 166.710 ;
        RECT 58.430 166.650 58.750 166.710 ;
        RECT 61.665 166.650 61.955 166.695 ;
        RECT 63.950 166.650 64.270 166.710 ;
        RECT 58.430 166.510 64.270 166.650 ;
        RECT 58.430 166.450 58.750 166.510 ;
        RECT 61.665 166.465 61.955 166.510 ;
        RECT 63.950 166.450 64.270 166.510 ;
        RECT 65.790 166.450 66.110 166.710 ;
        RECT 75.450 166.450 75.770 166.710 ;
        RECT 76.385 166.465 76.675 166.695 ;
        RECT 53.830 166.310 54.150 166.370 ;
        RECT 67.170 166.310 67.490 166.370 ;
        RECT 76.460 166.310 76.600 166.465 ;
        RECT 77.290 166.450 77.610 166.710 ;
        RECT 77.840 166.695 77.980 167.190 ;
        RECT 80.510 167.130 80.830 167.190 ;
        RECT 81.060 167.190 82.120 167.330 ;
        RECT 77.765 166.465 78.055 166.695 ;
        RECT 78.325 166.650 78.615 166.695 ;
        RECT 79.590 166.650 79.910 166.710 ;
        RECT 81.060 166.695 81.200 167.190 ;
        RECT 81.980 166.990 82.120 167.190 ;
        RECT 87.410 167.190 93.160 167.330 ;
        RECT 87.410 167.130 87.730 167.190 ;
        RECT 93.020 166.990 93.160 167.190 ;
        RECT 97.990 167.190 108.890 167.330 ;
        RECT 97.990 167.130 98.310 167.190 ;
        RECT 105.810 167.130 106.130 167.190 ;
        RECT 108.570 167.130 108.890 167.190 ;
        RECT 95.705 166.990 95.995 167.035 ;
        RECT 98.860 166.990 99.150 167.035 ;
        RECT 102.120 166.990 102.410 167.035 ;
        RECT 81.980 166.850 92.700 166.990 ;
        RECT 93.020 166.850 95.460 166.990 ;
        RECT 78.300 166.640 78.615 166.650 ;
        RECT 79.220 166.640 79.910 166.650 ;
        RECT 78.300 166.510 79.910 166.640 ;
        RECT 78.300 166.500 79.360 166.510 ;
        RECT 78.325 166.465 78.615 166.500 ;
        RECT 79.590 166.450 79.910 166.510 ;
        RECT 80.065 166.465 80.355 166.695 ;
        RECT 80.985 166.465 81.275 166.695 ;
        RECT 80.140 166.310 80.280 166.465 ;
        RECT 81.430 166.450 81.750 166.710 ;
        RECT 81.890 166.450 82.210 166.710 ;
        RECT 86.030 166.450 86.350 166.710 ;
        RECT 53.000 166.170 67.490 166.310 ;
        RECT 50.625 166.125 50.915 166.170 ;
        RECT 51.530 166.110 51.850 166.170 ;
        RECT 53.830 166.110 54.150 166.170 ;
        RECT 67.170 166.110 67.490 166.170 ;
        RECT 74.620 166.170 80.280 166.310 ;
        RECT 85.110 166.310 85.430 166.370 ;
        RECT 86.505 166.310 86.795 166.355 ;
        RECT 85.110 166.170 86.795 166.310 ;
        RECT 74.620 166.015 74.760 166.170 ;
        RECT 78.760 166.030 78.900 166.170 ;
        RECT 85.110 166.110 85.430 166.170 ;
        RECT 86.505 166.125 86.795 166.170 ;
        RECT 86.950 166.110 87.270 166.370 ;
        RECT 92.560 166.310 92.700 166.850 ;
        RECT 92.945 166.650 93.235 166.695 ;
        RECT 94.310 166.650 94.630 166.710 ;
        RECT 95.320 166.695 95.460 166.850 ;
        RECT 95.705 166.850 102.410 166.990 ;
        RECT 95.705 166.805 95.995 166.850 ;
        RECT 98.860 166.805 99.150 166.850 ;
        RECT 102.120 166.805 102.410 166.850 ;
        RECT 103.040 166.990 103.330 167.035 ;
        RECT 104.900 166.990 105.190 167.035 ;
        RECT 116.405 166.990 116.695 167.035 ;
        RECT 116.850 166.990 117.170 167.050 ;
        RECT 103.040 166.850 105.190 166.990 ;
        RECT 103.040 166.805 103.330 166.850 ;
        RECT 104.900 166.805 105.190 166.850 ;
        RECT 105.440 166.850 116.160 166.990 ;
        RECT 92.945 166.510 94.630 166.650 ;
        RECT 92.945 166.465 93.235 166.510 ;
        RECT 94.310 166.450 94.630 166.510 ;
        RECT 95.245 166.650 95.535 166.695 ;
        RECT 100.720 166.650 101.010 166.695 ;
        RECT 103.040 166.650 103.255 166.805 ;
        RECT 95.245 166.510 100.520 166.650 ;
        RECT 95.245 166.465 95.535 166.510 ;
        RECT 94.770 166.310 95.090 166.370 ;
        RECT 96.855 166.310 97.145 166.355 ;
        RECT 98.450 166.310 98.770 166.370 ;
        RECT 92.560 166.170 98.770 166.310 ;
        RECT 100.380 166.310 100.520 166.510 ;
        RECT 100.720 166.510 103.255 166.650 ;
        RECT 100.720 166.465 101.010 166.510 ;
        RECT 103.970 166.450 104.290 166.710 ;
        RECT 105.440 166.310 105.580 166.850 ;
        RECT 108.570 166.650 108.890 166.710 ;
        RECT 109.505 166.650 109.795 166.695 ;
        RECT 108.570 166.510 109.795 166.650 ;
        RECT 108.570 166.450 108.890 166.510 ;
        RECT 109.505 166.465 109.795 166.510 ;
        RECT 109.950 166.450 110.270 166.710 ;
        RECT 110.410 166.450 110.730 166.710 ;
        RECT 111.330 166.450 111.650 166.710 ;
        RECT 116.020 166.695 116.160 166.850 ;
        RECT 116.405 166.850 117.170 166.990 ;
        RECT 116.405 166.805 116.695 166.850 ;
        RECT 116.850 166.790 117.170 166.850 ;
        RECT 115.945 166.650 116.235 166.695 ;
        RECT 118.245 166.650 118.535 166.695 ;
        RECT 118.690 166.650 119.010 166.710 ;
        RECT 115.945 166.510 119.010 166.650 ;
        RECT 115.945 166.465 116.235 166.510 ;
        RECT 118.245 166.465 118.535 166.510 ;
        RECT 118.690 166.450 119.010 166.510 ;
        RECT 119.610 166.450 119.930 166.710 ;
        RECT 100.380 166.170 105.580 166.310 ;
        RECT 105.825 166.310 106.115 166.355 ;
        RECT 124.210 166.310 124.530 166.370 ;
        RECT 105.825 166.170 124.530 166.310 ;
        RECT 94.770 166.110 95.090 166.170 ;
        RECT 96.855 166.125 97.145 166.170 ;
        RECT 98.450 166.110 98.770 166.170 ;
        RECT 105.825 166.125 106.115 166.170 ;
        RECT 124.210 166.110 124.530 166.170 ;
        RECT 74.545 165.970 74.835 166.015 ;
        RECT 47.480 165.830 74.835 165.970 ;
        RECT 74.545 165.785 74.835 165.830 ;
        RECT 78.670 165.770 78.990 166.030 ;
        RECT 100.720 165.970 101.010 166.015 ;
        RECT 103.500 165.970 103.790 166.015 ;
        RECT 105.360 165.970 105.650 166.015 ;
        RECT 100.720 165.830 105.650 165.970 ;
        RECT 100.720 165.785 101.010 165.830 ;
        RECT 103.500 165.785 103.790 165.830 ;
        RECT 105.360 165.785 105.650 165.830 ;
        RECT 42.790 165.630 43.110 165.690 ;
        RECT 40.580 165.490 43.110 165.630 ;
        RECT 42.790 165.430 43.110 165.490 ;
        RECT 43.250 165.430 43.570 165.690 ;
        RECT 46.010 165.630 46.330 165.690 ;
        RECT 46.945 165.630 47.235 165.675 ;
        RECT 46.010 165.490 47.235 165.630 ;
        RECT 46.010 165.430 46.330 165.490 ;
        RECT 46.945 165.445 47.235 165.490 ;
        RECT 50.610 165.630 50.930 165.690 ;
        RECT 51.085 165.630 51.375 165.675 ;
        RECT 50.610 165.490 51.375 165.630 ;
        RECT 50.610 165.430 50.930 165.490 ;
        RECT 51.085 165.445 51.375 165.490 ;
        RECT 61.190 165.630 61.510 165.690 ;
        RECT 62.125 165.630 62.415 165.675 ;
        RECT 61.190 165.490 62.415 165.630 ;
        RECT 61.190 165.430 61.510 165.490 ;
        RECT 62.125 165.445 62.415 165.490 ;
        RECT 66.725 165.630 67.015 165.675 ;
        RECT 67.170 165.630 67.490 165.690 ;
        RECT 66.725 165.490 67.490 165.630 ;
        RECT 66.725 165.445 67.015 165.490 ;
        RECT 67.170 165.430 67.490 165.490 ;
        RECT 79.605 165.630 79.895 165.675 ;
        RECT 80.050 165.630 80.370 165.690 ;
        RECT 79.605 165.490 80.370 165.630 ;
        RECT 79.605 165.445 79.895 165.490 ;
        RECT 80.050 165.430 80.370 165.490 ;
        RECT 83.270 165.430 83.590 165.690 ;
        RECT 84.190 165.430 84.510 165.690 ;
        RECT 93.865 165.630 94.155 165.675 ;
        RECT 96.610 165.630 96.930 165.690 ;
        RECT 93.865 165.490 96.930 165.630 ;
        RECT 93.865 165.445 94.155 165.490 ;
        RECT 96.610 165.430 96.930 165.490 ;
        RECT 108.125 165.630 108.415 165.675 ;
        RECT 110.410 165.630 110.730 165.690 ;
        RECT 108.125 165.490 110.730 165.630 ;
        RECT 108.125 165.445 108.415 165.490 ;
        RECT 110.410 165.430 110.730 165.490 ;
        RECT 135.580 165.470 136.830 166.590 ;
        RECT 14.660 164.810 127.820 165.290 ;
        RECT 17.950 164.610 18.270 164.670 ;
        RECT 25.310 164.610 25.630 164.670 ;
        RECT 25.785 164.610 26.075 164.655 ;
        RECT 39.570 164.610 39.890 164.670 ;
        RECT 17.950 164.470 23.010 164.610 ;
        RECT 17.950 164.410 18.270 164.470 ;
        RECT 21.170 163.730 21.490 163.990 ;
        RECT 21.720 163.975 21.860 164.470 ;
        RECT 22.870 164.270 23.010 164.470 ;
        RECT 25.310 164.470 26.075 164.610 ;
        RECT 25.310 164.410 25.630 164.470 ;
        RECT 25.785 164.425 26.075 164.470 ;
        RECT 33.680 164.470 39.890 164.610 ;
        RECT 33.680 164.270 33.820 164.470 ;
        RECT 39.570 164.410 39.890 164.470 ;
        RECT 42.330 164.610 42.650 164.670 ;
        RECT 45.550 164.610 45.870 164.670 ;
        RECT 42.330 164.470 45.870 164.610 ;
        RECT 42.330 164.410 42.650 164.470 ;
        RECT 45.550 164.410 45.870 164.470 ;
        RECT 67.170 164.610 67.490 164.670 ;
        RECT 74.990 164.610 75.310 164.670 ;
        RECT 83.270 164.610 83.590 164.670 ;
        RECT 92.945 164.610 93.235 164.655 ;
        RECT 94.310 164.610 94.630 164.670 ;
        RECT 67.170 164.470 71.310 164.610 ;
        RECT 67.170 164.410 67.490 164.470 ;
        RECT 22.870 164.130 33.820 164.270 ;
        RECT 34.165 164.270 34.455 164.315 ;
        RECT 37.285 164.270 37.575 164.315 ;
        RECT 39.175 164.270 39.465 164.315 ;
        RECT 34.165 164.130 39.465 164.270 ;
        RECT 34.165 164.085 34.455 164.130 ;
        RECT 37.285 164.085 37.575 164.130 ;
        RECT 39.175 164.085 39.465 164.130 ;
        RECT 41.410 164.270 41.730 164.330 ;
        RECT 45.090 164.270 45.410 164.330 ;
        RECT 41.410 164.130 45.410 164.270 ;
        RECT 41.410 164.070 41.730 164.130 ;
        RECT 21.645 163.745 21.935 163.975 ;
        RECT 31.305 163.930 31.595 163.975 ;
        RECT 36.350 163.930 36.670 163.990 ;
        RECT 22.870 163.790 28.760 163.930 ;
        RECT 22.870 163.310 23.010 163.790 ;
        RECT 28.620 163.635 28.760 163.790 ;
        RECT 31.305 163.790 36.670 163.930 ;
        RECT 31.305 163.745 31.595 163.790 ;
        RECT 36.350 163.730 36.670 163.790 ;
        RECT 38.650 163.730 38.970 163.990 ;
        RECT 40.580 163.790 42.100 163.930 ;
        RECT 24.865 163.590 25.155 163.635 ;
        RECT 22.550 163.110 23.010 163.310 ;
        RECT 24.020 163.450 25.155 163.590 ;
        RECT 22.550 163.050 22.870 163.110 ;
        RECT 21.630 162.910 21.950 162.970 ;
        RECT 24.020 162.955 24.160 163.450 ;
        RECT 24.865 163.405 25.155 163.450 ;
        RECT 28.545 163.590 28.835 163.635 ;
        RECT 29.910 163.590 30.230 163.650 ;
        RECT 28.545 163.450 30.230 163.590 ;
        RECT 28.545 163.405 28.835 163.450 ;
        RECT 29.910 163.390 30.230 163.450 ;
        RECT 33.085 163.295 33.375 163.610 ;
        RECT 34.165 163.590 34.455 163.635 ;
        RECT 37.745 163.590 38.035 163.635 ;
        RECT 39.580 163.590 39.870 163.635 ;
        RECT 34.165 163.450 39.870 163.590 ;
        RECT 34.165 163.405 34.455 163.450 ;
        RECT 37.745 163.405 38.035 163.450 ;
        RECT 39.580 163.405 39.870 163.450 ;
        RECT 40.030 163.390 40.350 163.650 ;
        RECT 29.005 163.250 29.295 163.295 ;
        RECT 32.785 163.250 33.375 163.295 ;
        RECT 36.025 163.250 36.675 163.295 ;
        RECT 29.005 163.110 36.675 163.250 ;
        RECT 29.005 163.065 29.295 163.110 ;
        RECT 32.785 163.065 33.075 163.110 ;
        RECT 36.025 163.065 36.675 163.110 ;
        RECT 22.105 162.910 22.395 162.955 ;
        RECT 21.630 162.770 22.395 162.910 ;
        RECT 21.630 162.710 21.950 162.770 ;
        RECT 22.105 162.725 22.395 162.770 ;
        RECT 23.945 162.725 24.235 162.955 ;
        RECT 30.370 162.710 30.690 162.970 ;
        RECT 31.290 162.910 31.610 162.970 ;
        RECT 40.580 162.910 40.720 163.790 ;
        RECT 40.950 163.390 41.270 163.650 ;
        RECT 41.960 163.635 42.100 163.790 ;
        RECT 42.420 163.635 42.560 164.130 ;
        RECT 45.090 164.070 45.410 164.130 ;
        RECT 63.920 164.270 64.210 164.315 ;
        RECT 66.700 164.270 66.990 164.315 ;
        RECT 68.560 164.270 68.850 164.315 ;
        RECT 63.920 164.130 68.850 164.270 ;
        RECT 71.170 164.270 71.310 164.470 ;
        RECT 74.990 164.470 83.590 164.610 ;
        RECT 74.990 164.410 75.310 164.470 ;
        RECT 83.270 164.410 83.590 164.470 ;
        RECT 87.040 164.470 92.700 164.610 ;
        RECT 87.040 164.270 87.180 164.470 ;
        RECT 71.170 164.130 87.180 164.270 ;
        RECT 87.380 164.270 87.670 164.315 ;
        RECT 90.160 164.270 90.450 164.315 ;
        RECT 92.020 164.270 92.310 164.315 ;
        RECT 87.380 164.130 92.310 164.270 ;
        RECT 92.560 164.270 92.700 164.470 ;
        RECT 92.945 164.470 94.630 164.610 ;
        RECT 92.945 164.425 93.235 164.470 ;
        RECT 94.310 164.410 94.630 164.470 ;
        RECT 108.570 164.610 108.890 164.670 ;
        RECT 112.250 164.610 112.570 164.670 ;
        RECT 108.570 164.470 112.570 164.610 ;
        RECT 108.570 164.410 108.890 164.470 ;
        RECT 112.250 164.410 112.570 164.470 ;
        RECT 111.330 164.270 111.650 164.330 ;
        RECT 92.560 164.130 100.060 164.270 ;
        RECT 63.920 164.085 64.210 164.130 ;
        RECT 66.700 164.085 66.990 164.130 ;
        RECT 68.560 164.085 68.850 164.130 ;
        RECT 87.380 164.085 87.670 164.130 ;
        RECT 90.160 164.085 90.450 164.130 ;
        RECT 92.020 164.085 92.310 164.130 ;
        RECT 56.590 163.930 56.910 163.990 ;
        RECT 42.880 163.790 46.700 163.930 ;
        RECT 42.880 163.635 43.020 163.790 ;
        RECT 41.885 163.405 42.175 163.635 ;
        RECT 42.345 163.405 42.635 163.635 ;
        RECT 42.805 163.405 43.095 163.635 ;
        RECT 44.170 163.590 44.490 163.650 ;
        RECT 44.645 163.590 44.935 163.635 ;
        RECT 44.170 163.450 44.935 163.590 ;
        RECT 44.170 163.390 44.490 163.450 ;
        RECT 44.645 163.405 44.935 163.450 ;
        RECT 45.550 163.390 45.870 163.650 ;
        RECT 46.560 163.635 46.700 163.790 ;
        RECT 56.590 163.790 66.940 163.930 ;
        RECT 56.590 163.730 56.910 163.790 ;
        RECT 46.025 163.405 46.315 163.635 ;
        RECT 46.485 163.590 46.775 163.635 ;
        RECT 46.930 163.590 47.250 163.650 ;
        RECT 50.150 163.590 50.470 163.650 ;
        RECT 46.485 163.450 50.470 163.590 ;
        RECT 46.485 163.405 46.775 163.450 ;
        RECT 41.040 163.250 41.180 163.390 ;
        RECT 44.260 163.250 44.400 163.390 ;
        RECT 41.040 163.110 44.400 163.250 ;
        RECT 45.090 163.250 45.410 163.310 ;
        RECT 46.100 163.250 46.240 163.405 ;
        RECT 46.930 163.390 47.250 163.450 ;
        RECT 50.150 163.390 50.470 163.450 ;
        RECT 63.920 163.590 64.210 163.635 ;
        RECT 66.800 163.590 66.940 163.790 ;
        RECT 67.170 163.730 67.490 163.990 ;
        RECT 83.515 163.930 83.805 163.975 ;
        RECT 85.110 163.930 85.430 163.990 ;
        RECT 81.520 163.790 85.430 163.930 ;
        RECT 67.630 163.590 67.950 163.650 ;
        RECT 69.025 163.590 69.315 163.635 ;
        RECT 63.920 163.450 66.455 163.590 ;
        RECT 66.800 163.450 69.315 163.590 ;
        RECT 63.920 163.405 64.210 163.450 ;
        RECT 52.910 163.250 53.230 163.310 ;
        RECT 45.090 163.110 53.230 163.250 ;
        RECT 45.090 163.050 45.410 163.110 ;
        RECT 52.910 163.050 53.230 163.110 ;
        RECT 59.350 163.250 59.670 163.310 ;
        RECT 61.190 163.250 61.510 163.310 ;
        RECT 66.240 163.295 66.455 163.450 ;
        RECT 67.630 163.390 67.950 163.450 ;
        RECT 69.025 163.405 69.315 163.450 ;
        RECT 75.450 163.390 75.770 163.650 ;
        RECT 78.670 163.590 78.990 163.650 ;
        RECT 79.590 163.590 79.910 163.650 ;
        RECT 78.670 163.450 80.280 163.590 ;
        RECT 78.670 163.390 78.990 163.450 ;
        RECT 79.590 163.390 79.910 163.450 ;
        RECT 62.060 163.250 62.350 163.295 ;
        RECT 65.320 163.250 65.610 163.295 ;
        RECT 59.350 163.110 60.960 163.250 ;
        RECT 59.350 163.050 59.670 163.110 ;
        RECT 31.290 162.770 40.720 162.910 ;
        RECT 31.290 162.710 31.610 162.770 ;
        RECT 44.170 162.710 44.490 162.970 ;
        RECT 47.865 162.910 48.155 162.955 ;
        RECT 52.450 162.910 52.770 162.970 ;
        RECT 60.270 162.955 60.590 162.970 ;
        RECT 47.865 162.770 52.770 162.910 ;
        RECT 47.865 162.725 48.155 162.770 ;
        RECT 52.450 162.710 52.770 162.770 ;
        RECT 60.055 162.725 60.590 162.955 ;
        RECT 60.820 162.910 60.960 163.110 ;
        RECT 61.190 163.110 65.610 163.250 ;
        RECT 61.190 163.050 61.510 163.110 ;
        RECT 62.060 163.065 62.350 163.110 ;
        RECT 65.320 163.065 65.610 163.110 ;
        RECT 66.240 163.250 66.530 163.295 ;
        RECT 68.100 163.250 68.390 163.295 ;
        RECT 80.140 163.250 80.280 163.450 ;
        RECT 80.510 163.390 80.830 163.650 ;
        RECT 80.970 163.390 81.290 163.650 ;
        RECT 81.520 163.635 81.660 163.790 ;
        RECT 83.515 163.745 83.805 163.790 ;
        RECT 85.110 163.730 85.430 163.790 ;
        RECT 85.570 163.930 85.890 163.990 ;
        RECT 90.645 163.930 90.935 163.975 ;
        RECT 85.570 163.790 90.935 163.930 ;
        RECT 85.570 163.730 85.890 163.790 ;
        RECT 90.645 163.745 90.935 163.790 ;
        RECT 92.485 163.930 92.775 163.975 ;
        RECT 93.850 163.930 94.170 163.990 ;
        RECT 95.705 163.930 95.995 163.975 ;
        RECT 92.485 163.790 94.170 163.930 ;
        RECT 92.485 163.745 92.775 163.790 ;
        RECT 93.850 163.730 94.170 163.790 ;
        RECT 94.400 163.790 95.995 163.930 ;
        RECT 81.445 163.405 81.735 163.635 ;
        RECT 82.365 163.405 82.655 163.635 ;
        RECT 87.380 163.590 87.670 163.635 ;
        RECT 91.090 163.590 91.410 163.650 ;
        RECT 94.400 163.590 94.540 163.790 ;
        RECT 95.705 163.745 95.995 163.790 ;
        RECT 87.380 163.450 89.915 163.590 ;
        RECT 87.380 163.405 87.670 163.450 ;
        RECT 82.440 163.250 82.580 163.405 ;
        RECT 66.240 163.110 68.390 163.250 ;
        RECT 66.240 163.065 66.530 163.110 ;
        RECT 68.100 163.065 68.390 163.110 ;
        RECT 74.620 163.110 79.820 163.250 ;
        RECT 80.140 163.110 82.580 163.250 ;
        RECT 85.520 163.250 85.810 163.295 ;
        RECT 86.490 163.250 86.810 163.310 ;
        RECT 89.700 163.295 89.915 163.450 ;
        RECT 91.090 163.450 94.540 163.590 ;
        RECT 91.090 163.390 91.410 163.450 ;
        RECT 94.770 163.390 95.090 163.650 ;
        RECT 97.990 163.590 98.310 163.650 ;
        RECT 99.920 163.635 100.060 164.130 ;
        RECT 101.300 164.130 111.650 164.270 ;
        RECT 101.300 163.650 101.440 164.130 ;
        RECT 111.330 164.070 111.650 164.130 ;
        RECT 109.030 163.930 109.350 163.990 ;
        RECT 111.420 163.930 111.560 164.070 ;
        RECT 109.030 163.790 110.640 163.930 ;
        RECT 109.030 163.730 109.350 163.790 ;
        RECT 99.385 163.590 99.675 163.635 ;
        RECT 97.990 163.450 99.675 163.590 ;
        RECT 97.990 163.390 98.310 163.450 ;
        RECT 99.385 163.405 99.675 163.450 ;
        RECT 99.845 163.405 100.135 163.635 ;
        RECT 88.780 163.250 89.070 163.295 ;
        RECT 85.520 163.110 89.070 163.250 ;
        RECT 74.620 162.955 74.760 163.110 ;
        RECT 74.545 162.910 74.835 162.955 ;
        RECT 60.820 162.770 74.835 162.910 ;
        RECT 74.545 162.725 74.835 162.770 ;
        RECT 76.370 162.910 76.690 162.970 ;
        RECT 79.145 162.910 79.435 162.955 ;
        RECT 76.370 162.770 79.435 162.910 ;
        RECT 79.680 162.910 79.820 163.110 ;
        RECT 85.520 163.065 85.810 163.110 ;
        RECT 86.490 163.050 86.810 163.110 ;
        RECT 88.780 163.065 89.070 163.110 ;
        RECT 89.700 163.250 89.990 163.295 ;
        RECT 91.560 163.250 91.850 163.295 ;
        RECT 89.700 163.110 91.850 163.250 ;
        RECT 99.920 163.250 100.060 163.405 ;
        RECT 100.290 163.390 100.610 163.650 ;
        RECT 101.210 163.390 101.530 163.650 ;
        RECT 108.570 163.590 108.890 163.650 ;
        RECT 109.505 163.590 109.795 163.635 ;
        RECT 108.570 163.450 109.795 163.590 ;
        RECT 108.570 163.390 108.890 163.450 ;
        RECT 109.505 163.405 109.795 163.450 ;
        RECT 109.950 163.390 110.270 163.650 ;
        RECT 110.500 163.635 110.640 163.790 ;
        RECT 111.420 163.790 115.240 163.930 ;
        RECT 111.420 163.635 111.560 163.790 ;
        RECT 110.425 163.405 110.715 163.635 ;
        RECT 111.345 163.405 111.635 163.635 ;
        RECT 112.250 163.590 112.570 163.650 ;
        RECT 113.185 163.590 113.475 163.635 ;
        RECT 112.250 163.450 113.475 163.590 ;
        RECT 112.250 163.390 112.570 163.450 ;
        RECT 113.185 163.405 113.475 163.450 ;
        RECT 113.645 163.405 113.935 163.635 ;
        RECT 114.105 163.590 114.395 163.635 ;
        RECT 114.550 163.590 114.870 163.650 ;
        RECT 115.100 163.635 115.240 163.790 ;
        RECT 114.105 163.450 114.870 163.590 ;
        RECT 114.105 163.405 114.395 163.450 ;
        RECT 106.270 163.250 106.590 163.310 ;
        RECT 110.040 163.250 110.180 163.390 ;
        RECT 113.720 163.250 113.860 163.405 ;
        RECT 114.550 163.390 114.870 163.450 ;
        RECT 115.025 163.405 115.315 163.635 ;
        RECT 99.920 163.110 113.860 163.250 ;
        RECT 89.700 163.065 89.990 163.110 ;
        RECT 91.560 163.065 91.850 163.110 ;
        RECT 106.270 163.050 106.590 163.110 ;
        RECT 83.730 162.910 84.050 162.970 ;
        RECT 79.680 162.770 84.050 162.910 ;
        RECT 60.270 162.710 60.590 162.725 ;
        RECT 76.370 162.710 76.690 162.770 ;
        RECT 79.145 162.725 79.435 162.770 ;
        RECT 83.730 162.710 84.050 162.770 ;
        RECT 86.030 162.910 86.350 162.970 ;
        RECT 95.245 162.910 95.535 162.955 ;
        RECT 86.030 162.770 95.535 162.910 ;
        RECT 86.030 162.710 86.350 162.770 ;
        RECT 95.245 162.725 95.535 162.770 ;
        RECT 96.150 162.910 96.470 162.970 ;
        RECT 98.005 162.910 98.295 162.955 ;
        RECT 96.150 162.770 98.295 162.910 ;
        RECT 96.150 162.710 96.470 162.770 ;
        RECT 98.005 162.725 98.295 162.770 ;
        RECT 108.125 162.910 108.415 162.955 ;
        RECT 109.030 162.910 109.350 162.970 ;
        RECT 108.125 162.770 109.350 162.910 ;
        RECT 108.125 162.725 108.415 162.770 ;
        RECT 109.030 162.710 109.350 162.770 ;
        RECT 110.870 162.910 111.190 162.970 ;
        RECT 111.805 162.910 112.095 162.955 ;
        RECT 110.870 162.770 112.095 162.910 ;
        RECT 110.870 162.710 111.190 162.770 ;
        RECT 111.805 162.725 112.095 162.770 ;
        RECT 14.660 162.090 127.820 162.570 ;
        RECT 28.530 161.890 28.850 161.950 ;
        RECT 28.530 161.750 36.120 161.890 ;
        RECT 28.530 161.690 28.850 161.750 ;
        RECT 17.950 161.550 18.270 161.610 ;
        RECT 18.525 161.550 18.815 161.595 ;
        RECT 21.765 161.550 22.415 161.595 ;
        RECT 17.950 161.410 22.415 161.550 ;
        RECT 17.950 161.350 18.270 161.410 ;
        RECT 18.525 161.365 19.115 161.410 ;
        RECT 21.765 161.365 22.415 161.410 ;
        RECT 18.825 161.050 19.115 161.365 ;
        RECT 19.905 161.210 20.195 161.255 ;
        RECT 23.485 161.210 23.775 161.255 ;
        RECT 25.320 161.210 25.610 161.255 ;
        RECT 19.905 161.070 25.610 161.210 ;
        RECT 19.905 161.025 20.195 161.070 ;
        RECT 23.485 161.025 23.775 161.070 ;
        RECT 25.320 161.025 25.610 161.070 ;
        RECT 25.785 161.210 26.075 161.255 ;
        RECT 26.690 161.210 27.010 161.270 ;
        RECT 28.620 161.210 28.760 161.690 ;
        RECT 34.970 161.350 35.290 161.610 ;
        RECT 35.980 161.255 36.120 161.750 ;
        RECT 37.730 161.690 38.050 161.950 ;
        RECT 39.570 161.690 39.890 161.950 ;
        RECT 40.045 161.705 40.335 161.935 ;
        RECT 51.070 161.890 51.390 161.950 ;
        RECT 50.700 161.750 51.390 161.890 ;
        RECT 36.350 161.550 36.670 161.610 ;
        RECT 40.120 161.550 40.260 161.705 ;
        RECT 36.350 161.410 40.260 161.550 ;
        RECT 36.350 161.350 36.670 161.410 ;
        RECT 25.785 161.070 28.760 161.210 ;
        RECT 35.905 161.210 36.195 161.255 ;
        RECT 40.030 161.210 40.350 161.270 ;
        RECT 35.905 161.070 40.350 161.210 ;
        RECT 25.785 161.025 26.075 161.070 ;
        RECT 26.690 161.010 27.010 161.070 ;
        RECT 35.905 161.025 36.195 161.070 ;
        RECT 40.030 161.010 40.350 161.070 ;
        RECT 49.690 161.010 50.010 161.270 ;
        RECT 50.700 161.255 50.840 161.750 ;
        RECT 51.070 161.690 51.390 161.750 ;
        RECT 62.585 161.705 62.875 161.935 ;
        RECT 64.885 161.890 65.175 161.935 ;
        RECT 66.710 161.890 67.030 161.950 ;
        RECT 64.885 161.750 67.030 161.890 ;
        RECT 64.885 161.705 65.175 161.750 ;
        RECT 50.165 161.025 50.455 161.255 ;
        RECT 50.625 161.025 50.915 161.255 ;
        RECT 51.545 161.210 51.835 161.255 ;
        RECT 53.830 161.210 54.150 161.270 ;
        RECT 51.545 161.070 54.150 161.210 ;
        RECT 51.545 161.025 51.835 161.070 ;
        RECT 24.390 160.670 24.710 160.930 ;
        RECT 40.505 160.685 40.795 160.915 ;
        RECT 50.240 160.870 50.380 161.025 ;
        RECT 53.830 161.010 54.150 161.070 ;
        RECT 58.430 161.010 58.750 161.270 ;
        RECT 60.730 161.010 61.050 161.270 ;
        RECT 62.660 161.210 62.800 161.705 ;
        RECT 66.710 161.690 67.030 161.750 ;
        RECT 74.530 161.690 74.850 161.950 ;
        RECT 80.970 161.890 81.290 161.950 ;
        RECT 80.970 161.750 81.660 161.890 ;
        RECT 80.970 161.690 81.290 161.750 ;
        RECT 67.185 161.550 67.475 161.595 ;
        RECT 74.070 161.550 74.390 161.610 ;
        RECT 64.960 161.410 67.475 161.550 ;
        RECT 64.960 161.270 65.100 161.410 ;
        RECT 67.185 161.365 67.475 161.410 ;
        RECT 67.720 161.410 74.390 161.550 ;
        RECT 63.965 161.210 64.255 161.255 ;
        RECT 62.660 161.070 64.255 161.210 ;
        RECT 63.965 161.025 64.255 161.070 ;
        RECT 64.870 161.010 65.190 161.270 ;
        RECT 65.330 161.210 65.650 161.270 ;
        RECT 66.265 161.210 66.555 161.255 ;
        RECT 65.330 161.070 66.555 161.210 ;
        RECT 65.330 161.010 65.650 161.070 ;
        RECT 66.265 161.025 66.555 161.070 ;
        RECT 66.725 161.210 67.015 161.255 ;
        RECT 67.720 161.210 67.860 161.410 ;
        RECT 74.070 161.350 74.390 161.410 ;
        RECT 66.725 161.070 67.860 161.210 ;
        RECT 66.725 161.025 67.015 161.070 ;
        RECT 68.090 161.010 68.410 161.270 ;
        RECT 74.620 161.255 74.760 161.690 ;
        RECT 74.545 161.210 74.835 161.255 ;
        RECT 74.160 161.070 74.835 161.210 ;
        RECT 74.160 160.930 74.300 161.070 ;
        RECT 74.545 161.025 74.835 161.070 ;
        RECT 79.590 161.210 79.910 161.270 ;
        RECT 81.520 161.255 81.660 161.750 ;
        RECT 85.570 161.690 85.890 161.950 ;
        RECT 86.490 161.690 86.810 161.950 ;
        RECT 101.210 161.890 101.530 161.950 ;
        RECT 104.890 161.890 105.210 161.950 ;
        RECT 87.500 161.750 101.530 161.890 ;
        RECT 83.730 161.550 84.050 161.610 ;
        RECT 87.500 161.550 87.640 161.750 ;
        RECT 101.210 161.690 101.530 161.750 ;
        RECT 103.600 161.750 105.210 161.890 ;
        RECT 83.730 161.410 87.640 161.550 ;
        RECT 87.885 161.550 88.175 161.595 ;
        RECT 91.500 161.550 91.790 161.595 ;
        RECT 94.760 161.550 95.050 161.595 ;
        RECT 87.885 161.410 95.050 161.550 ;
        RECT 83.730 161.350 84.050 161.410 ;
        RECT 87.885 161.365 88.175 161.410 ;
        RECT 91.500 161.365 91.790 161.410 ;
        RECT 94.760 161.365 95.050 161.410 ;
        RECT 95.680 161.550 95.970 161.595 ;
        RECT 97.540 161.550 97.830 161.595 ;
        RECT 95.680 161.410 97.830 161.550 ;
        RECT 95.680 161.365 95.970 161.410 ;
        RECT 97.540 161.365 97.830 161.410 ;
        RECT 80.065 161.210 80.355 161.255 ;
        RECT 79.590 161.070 80.355 161.210 ;
        RECT 79.590 161.010 79.910 161.070 ;
        RECT 80.065 161.025 80.355 161.070 ;
        RECT 80.985 161.025 81.275 161.255 ;
        RECT 81.445 161.025 81.735 161.255 ;
        RECT 52.910 160.870 53.230 160.930 ;
        RECT 50.240 160.730 53.230 160.870 ;
        RECT 19.905 160.530 20.195 160.575 ;
        RECT 23.025 160.530 23.315 160.575 ;
        RECT 24.915 160.530 25.205 160.575 ;
        RECT 19.905 160.390 25.205 160.530 ;
        RECT 19.905 160.345 20.195 160.390 ;
        RECT 23.025 160.345 23.315 160.390 ;
        RECT 24.915 160.345 25.205 160.390 ;
        RECT 35.890 160.530 36.210 160.590 ;
        RECT 40.580 160.530 40.720 160.685 ;
        RECT 52.910 160.670 53.230 160.730 ;
        RECT 59.825 160.685 60.115 160.915 ;
        RECT 35.890 160.390 40.720 160.530 ;
        RECT 35.890 160.330 36.210 160.390 ;
        RECT 17.045 160.190 17.335 160.235 ;
        RECT 21.630 160.190 21.950 160.250 ;
        RECT 17.045 160.050 21.950 160.190 ;
        RECT 17.045 160.005 17.335 160.050 ;
        RECT 21.630 159.990 21.950 160.050 ;
        RECT 44.630 160.190 44.950 160.250 ;
        RECT 48.325 160.190 48.615 160.235 ;
        RECT 44.630 160.050 48.615 160.190 ;
        RECT 44.630 159.990 44.950 160.050 ;
        RECT 48.325 160.005 48.615 160.050 ;
        RECT 57.970 159.990 58.290 160.250 ;
        RECT 59.900 160.190 60.040 160.685 ;
        RECT 60.270 160.670 60.590 160.930 ;
        RECT 74.070 160.670 74.390 160.930 ;
        RECT 61.190 160.530 61.510 160.590 ;
        RECT 81.060 160.530 81.200 161.025 ;
        RECT 81.890 161.010 82.210 161.270 ;
        RECT 84.190 161.210 84.510 161.270 ;
        RECT 84.665 161.210 84.955 161.255 ;
        RECT 84.190 161.070 84.955 161.210 ;
        RECT 84.190 161.010 84.510 161.070 ;
        RECT 84.665 161.025 84.955 161.070 ;
        RECT 86.965 161.210 87.255 161.255 ;
        RECT 87.410 161.210 87.730 161.270 ;
        RECT 86.965 161.070 87.730 161.210 ;
        RECT 86.965 161.025 87.255 161.070 ;
        RECT 87.410 161.010 87.730 161.070 ;
        RECT 93.360 161.210 93.650 161.255 ;
        RECT 95.680 161.210 95.895 161.365 ;
        RECT 93.360 161.070 95.895 161.210 ;
        RECT 93.360 161.025 93.650 161.070 ;
        RECT 96.610 161.010 96.930 161.270 ;
        RECT 101.670 161.210 101.990 161.270 ;
        RECT 103.600 161.255 103.740 161.750 ;
        RECT 104.890 161.690 105.210 161.750 ;
        RECT 102.605 161.210 102.895 161.255 ;
        RECT 101.670 161.070 102.895 161.210 ;
        RECT 101.670 161.010 101.990 161.070 ;
        RECT 102.605 161.025 102.895 161.070 ;
        RECT 103.525 161.025 103.815 161.255 ;
        RECT 103.970 161.010 104.290 161.270 ;
        RECT 104.445 161.210 104.735 161.255 ;
        RECT 104.890 161.210 105.210 161.270 ;
        RECT 104.445 161.070 105.210 161.210 ;
        RECT 104.445 161.025 104.735 161.070 ;
        RECT 104.890 161.010 105.210 161.070 ;
        RECT 115.470 161.210 115.790 161.270 ;
        RECT 118.690 161.210 119.010 161.270 ;
        RECT 115.470 161.070 119.010 161.210 ;
        RECT 115.470 161.010 115.790 161.070 ;
        RECT 118.690 161.010 119.010 161.070 ;
        RECT 83.270 160.670 83.590 160.930 ;
        RECT 93.850 160.870 94.170 160.930 ;
        RECT 97.070 160.870 97.390 160.930 ;
        RECT 98.465 160.870 98.755 160.915 ;
        RECT 93.850 160.730 98.755 160.870 ;
        RECT 93.850 160.670 94.170 160.730 ;
        RECT 97.070 160.670 97.390 160.730 ;
        RECT 98.465 160.685 98.755 160.730 ;
        RECT 86.030 160.530 86.350 160.590 ;
        RECT 89.495 160.530 89.785 160.575 ;
        RECT 61.190 160.390 73.840 160.530 ;
        RECT 81.060 160.390 89.785 160.530 ;
        RECT 61.190 160.330 61.510 160.390 ;
        RECT 64.870 160.190 65.190 160.250 ;
        RECT 59.900 160.050 65.190 160.190 ;
        RECT 64.870 159.990 65.190 160.050 ;
        RECT 65.345 160.190 65.635 160.235 ;
        RECT 65.790 160.190 66.110 160.250 ;
        RECT 73.700 160.235 73.840 160.390 ;
        RECT 86.030 160.330 86.350 160.390 ;
        RECT 89.495 160.345 89.785 160.390 ;
        RECT 93.360 160.530 93.650 160.575 ;
        RECT 96.140 160.530 96.430 160.575 ;
        RECT 98.000 160.530 98.290 160.575 ;
        RECT 93.360 160.390 98.290 160.530 ;
        RECT 93.360 160.345 93.650 160.390 ;
        RECT 96.140 160.345 96.430 160.390 ;
        RECT 98.000 160.345 98.290 160.390 ;
        RECT 65.345 160.050 66.110 160.190 ;
        RECT 65.345 160.005 65.635 160.050 ;
        RECT 65.790 159.990 66.110 160.050 ;
        RECT 73.625 160.190 73.915 160.235 ;
        RECT 99.370 160.190 99.690 160.250 ;
        RECT 73.625 160.050 99.690 160.190 ;
        RECT 73.625 160.005 73.915 160.050 ;
        RECT 99.370 159.990 99.690 160.050 ;
        RECT 105.810 159.990 106.130 160.250 ;
        RECT 119.150 159.990 119.470 160.250 ;
        RECT 14.660 159.370 127.820 159.850 ;
        RECT 17.950 158.970 18.270 159.230 ;
        RECT 24.390 159.170 24.710 159.230 ;
        RECT 24.865 159.170 25.155 159.215 ;
        RECT 24.390 159.030 25.155 159.170 ;
        RECT 24.390 158.970 24.710 159.030 ;
        RECT 24.865 158.985 25.155 159.030 ;
        RECT 39.570 159.170 39.890 159.230 ;
        RECT 57.510 159.170 57.830 159.230 ;
        RECT 58.675 159.170 58.965 159.215 ;
        RECT 68.090 159.170 68.410 159.230 ;
        RECT 39.570 159.030 49.000 159.170 ;
        RECT 39.570 158.970 39.890 159.030 ;
        RECT 23.945 158.645 24.235 158.875 ;
        RECT 34.480 158.830 34.770 158.875 ;
        RECT 37.260 158.830 37.550 158.875 ;
        RECT 39.120 158.830 39.410 158.875 ;
        RECT 34.480 158.690 39.410 158.830 ;
        RECT 34.480 158.645 34.770 158.690 ;
        RECT 37.260 158.645 37.550 158.690 ;
        RECT 39.120 158.645 39.410 158.690 ;
        RECT 21.170 158.290 21.490 158.550 ;
        RECT 18.425 158.150 18.715 158.195 ;
        RECT 18.885 158.150 19.175 158.195 ;
        RECT 22.550 158.150 22.870 158.210 ;
        RECT 18.425 158.010 22.870 158.150 ;
        RECT 24.020 158.150 24.160 158.645 ;
        RECT 30.615 158.490 30.905 158.535 ;
        RECT 34.050 158.490 34.370 158.550 ;
        RECT 30.615 158.350 34.370 158.490 ;
        RECT 30.615 158.305 30.905 158.350 ;
        RECT 34.050 158.290 34.370 158.350 ;
        RECT 39.585 158.490 39.875 158.535 ;
        RECT 40.030 158.490 40.350 158.550 ;
        RECT 39.585 158.350 40.350 158.490 ;
        RECT 39.585 158.305 39.875 158.350 ;
        RECT 40.030 158.290 40.350 158.350 ;
        RECT 25.785 158.150 26.075 158.195 ;
        RECT 24.020 158.010 26.075 158.150 ;
        RECT 18.425 157.965 18.715 158.010 ;
        RECT 18.885 157.965 19.175 158.010 ;
        RECT 22.550 157.950 22.870 158.010 ;
        RECT 25.785 157.965 26.075 158.010 ;
        RECT 34.480 158.150 34.770 158.195 ;
        RECT 37.745 158.150 38.035 158.195 ;
        RECT 34.480 158.010 37.015 158.150 ;
        RECT 34.480 157.965 34.770 158.010 ;
        RECT 30.370 157.810 30.690 157.870 ;
        RECT 36.800 157.855 37.015 158.010 ;
        RECT 37.745 158.010 40.260 158.150 ;
        RECT 37.745 157.965 38.035 158.010 ;
        RECT 32.620 157.810 32.910 157.855 ;
        RECT 35.880 157.810 36.170 157.855 ;
        RECT 30.370 157.670 36.170 157.810 ;
        RECT 30.370 157.610 30.690 157.670 ;
        RECT 32.620 157.625 32.910 157.670 ;
        RECT 35.880 157.625 36.170 157.670 ;
        RECT 36.800 157.810 37.090 157.855 ;
        RECT 38.660 157.810 38.950 157.855 ;
        RECT 36.800 157.670 38.950 157.810 ;
        RECT 36.800 157.625 37.090 157.670 ;
        RECT 38.660 157.625 38.950 157.670 ;
        RECT 19.345 157.470 19.635 157.515 ;
        RECT 19.790 157.470 20.110 157.530 ;
        RECT 19.345 157.330 20.110 157.470 ;
        RECT 19.345 157.285 19.635 157.330 ;
        RECT 19.790 157.270 20.110 157.330 ;
        RECT 21.630 157.270 21.950 157.530 ;
        RECT 22.105 157.470 22.395 157.515 ;
        RECT 22.550 157.470 22.870 157.530 ;
        RECT 40.120 157.515 40.260 158.010 ;
        RECT 40.950 157.950 41.270 158.210 ;
        RECT 48.860 158.195 49.000 159.030 ;
        RECT 57.510 159.030 68.410 159.170 ;
        RECT 57.510 158.970 57.830 159.030 ;
        RECT 58.675 158.985 58.965 159.030 ;
        RECT 68.090 158.970 68.410 159.030 ;
        RECT 70.850 159.170 71.170 159.230 ;
        RECT 71.325 159.170 71.615 159.215 ;
        RECT 70.850 159.030 71.615 159.170 ;
        RECT 70.850 158.970 71.170 159.030 ;
        RECT 71.325 158.985 71.615 159.030 ;
        RECT 99.370 159.170 99.690 159.230 ;
        RECT 104.430 159.170 104.750 159.230 ;
        RECT 99.370 159.030 104.750 159.170 ;
        RECT 99.370 158.970 99.690 159.030 ;
        RECT 104.430 158.970 104.750 159.030 ;
        RECT 109.950 158.970 110.270 159.230 ;
        RECT 61.190 158.830 61.510 158.890 ;
        RECT 49.320 158.690 61.510 158.830 ;
        RECT 47.865 157.965 48.155 158.195 ;
        RECT 48.325 157.965 48.615 158.195 ;
        RECT 48.785 157.965 49.075 158.195 ;
        RECT 22.105 157.330 22.870 157.470 ;
        RECT 22.105 157.285 22.395 157.330 ;
        RECT 22.550 157.270 22.870 157.330 ;
        RECT 40.045 157.285 40.335 157.515 ;
        RECT 45.550 157.470 45.870 157.530 ;
        RECT 46.485 157.470 46.775 157.515 ;
        RECT 45.550 157.330 46.775 157.470 ;
        RECT 47.940 157.470 48.080 157.965 ;
        RECT 48.400 157.810 48.540 157.965 ;
        RECT 49.320 157.810 49.460 158.690 ;
        RECT 61.190 158.630 61.510 158.690 ;
        RECT 62.540 158.830 62.830 158.875 ;
        RECT 65.320 158.830 65.610 158.875 ;
        RECT 67.180 158.830 67.470 158.875 ;
        RECT 62.540 158.690 67.470 158.830 ;
        RECT 62.540 158.645 62.830 158.690 ;
        RECT 65.320 158.645 65.610 158.690 ;
        RECT 67.180 158.645 67.470 158.690 ;
        RECT 73.625 158.830 73.915 158.875 ;
        RECT 107.665 158.830 107.955 158.875 ;
        RECT 118.345 158.830 118.635 158.875 ;
        RECT 121.465 158.830 121.755 158.875 ;
        RECT 123.355 158.830 123.645 158.875 ;
        RECT 73.625 158.690 77.060 158.830 ;
        RECT 73.625 158.645 73.915 158.690 ;
        RECT 65.790 158.290 66.110 158.550 ;
        RECT 67.630 158.290 67.950 158.550 ;
        RECT 74.070 158.490 74.390 158.550 ;
        RECT 72.320 158.350 74.390 158.490 ;
        RECT 49.690 157.950 50.010 158.210 ;
        RECT 58.890 158.150 59.210 158.210 ;
        RECT 61.650 158.150 61.970 158.210 ;
        RECT 72.320 158.195 72.460 158.350 ;
        RECT 74.070 158.290 74.390 158.350 ;
        RECT 58.890 158.010 61.970 158.150 ;
        RECT 58.890 157.950 59.210 158.010 ;
        RECT 61.650 157.950 61.970 158.010 ;
        RECT 62.540 158.150 62.830 158.195 ;
        RECT 70.405 158.150 70.695 158.195 ;
        RECT 62.540 158.010 65.075 158.150 ;
        RECT 62.540 157.965 62.830 158.010 ;
        RECT 50.610 157.810 50.930 157.870 ;
        RECT 48.400 157.670 50.930 157.810 ;
        RECT 50.610 157.610 50.930 157.670 ;
        RECT 57.970 157.810 58.290 157.870 ;
        RECT 64.860 157.855 65.075 158.010 ;
        RECT 70.405 158.010 71.310 158.150 ;
        RECT 70.405 157.965 70.695 158.010 ;
        RECT 60.680 157.810 60.970 157.855 ;
        RECT 63.940 157.810 64.230 157.855 ;
        RECT 57.970 157.670 64.230 157.810 ;
        RECT 57.970 157.610 58.290 157.670 ;
        RECT 60.680 157.625 60.970 157.670 ;
        RECT 63.940 157.625 64.230 157.670 ;
        RECT 64.860 157.810 65.150 157.855 ;
        RECT 66.720 157.810 67.010 157.855 ;
        RECT 64.860 157.670 67.010 157.810 ;
        RECT 71.170 157.810 71.310 158.010 ;
        RECT 72.245 157.965 72.535 158.195 ;
        RECT 72.705 157.965 72.995 158.195 ;
        RECT 75.450 158.150 75.770 158.210 ;
        RECT 76.385 158.150 76.675 158.195 ;
        RECT 75.450 158.010 76.675 158.150 ;
        RECT 71.770 157.810 72.090 157.870 ;
        RECT 72.780 157.810 72.920 157.965 ;
        RECT 75.450 157.950 75.770 158.010 ;
        RECT 76.385 157.965 76.675 158.010 ;
        RECT 71.170 157.670 72.920 157.810 ;
        RECT 76.920 157.810 77.060 158.690 ;
        RECT 107.665 158.690 113.860 158.830 ;
        RECT 107.665 158.645 107.955 158.690 ;
        RECT 105.810 158.490 106.130 158.550 ;
        RECT 109.505 158.490 109.795 158.535 ;
        RECT 113.170 158.490 113.490 158.550 ;
        RECT 105.810 158.350 109.795 158.490 ;
        RECT 105.810 158.290 106.130 158.350 ;
        RECT 109.505 158.305 109.795 158.350 ;
        RECT 111.880 158.350 113.490 158.490 ;
        RECT 113.720 158.490 113.860 158.690 ;
        RECT 118.345 158.690 123.645 158.830 ;
        RECT 118.345 158.645 118.635 158.690 ;
        RECT 121.465 158.645 121.755 158.690 ;
        RECT 123.355 158.645 123.645 158.690 ;
        RECT 120.070 158.490 120.390 158.550 ;
        RECT 113.720 158.350 120.390 158.490 ;
        RECT 101.670 158.150 101.990 158.210 ;
        RECT 103.065 158.150 103.355 158.195 ;
        RECT 84.970 158.010 103.355 158.150 ;
        RECT 80.510 157.810 80.830 157.870 ;
        RECT 76.920 157.670 80.830 157.810 ;
        RECT 64.860 157.625 65.150 157.670 ;
        RECT 66.720 157.625 67.010 157.670 ;
        RECT 71.770 157.610 72.090 157.670 ;
        RECT 80.510 157.610 80.830 157.670 ;
        RECT 49.230 157.470 49.550 157.530 ;
        RECT 51.070 157.470 51.390 157.530 ;
        RECT 69.470 157.470 69.790 157.530 ;
        RECT 47.940 157.330 69.790 157.470 ;
        RECT 45.550 157.270 45.870 157.330 ;
        RECT 46.485 157.285 46.775 157.330 ;
        RECT 49.230 157.270 49.550 157.330 ;
        RECT 51.070 157.270 51.390 157.330 ;
        RECT 69.470 157.270 69.790 157.330 ;
        RECT 72.690 157.470 73.010 157.530 ;
        RECT 74.990 157.470 75.310 157.530 ;
        RECT 72.690 157.330 75.310 157.470 ;
        RECT 72.690 157.270 73.010 157.330 ;
        RECT 74.990 157.270 75.310 157.330 ;
        RECT 77.290 157.470 77.610 157.530 ;
        RECT 84.970 157.470 85.110 158.010 ;
        RECT 101.670 157.950 101.990 158.010 ;
        RECT 103.065 157.965 103.355 158.010 ;
        RECT 103.970 157.950 104.290 158.210 ;
        RECT 104.430 157.950 104.750 158.210 ;
        RECT 104.890 157.950 105.210 158.210 ;
        RECT 108.585 158.150 108.875 158.195 ;
        RECT 109.030 158.150 109.350 158.210 ;
        RECT 111.880 158.195 112.020 158.350 ;
        RECT 113.170 158.290 113.490 158.350 ;
        RECT 120.070 158.290 120.390 158.350 ;
        RECT 108.585 158.010 109.350 158.150 ;
        RECT 108.585 157.965 108.875 158.010 ;
        RECT 109.030 157.950 109.350 158.010 ;
        RECT 111.805 157.965 112.095 158.195 ;
        RECT 112.250 157.950 112.570 158.210 ;
        RECT 112.750 158.150 113.040 158.195 ;
        RECT 112.750 158.010 113.400 158.150 ;
        RECT 112.750 157.965 113.040 158.010 ;
        RECT 103.510 157.810 103.830 157.870 ;
        RECT 104.980 157.810 105.120 157.950 ;
        RECT 103.510 157.670 105.120 157.810 ;
        RECT 109.965 157.810 110.255 157.855 ;
        RECT 110.425 157.810 110.715 157.855 ;
        RECT 109.965 157.670 110.715 157.810 ;
        RECT 103.510 157.610 103.830 157.670 ;
        RECT 109.965 157.625 110.255 157.670 ;
        RECT 110.425 157.625 110.715 157.670 ;
        RECT 113.260 157.810 113.400 158.010 ;
        RECT 113.630 157.950 113.950 158.210 ;
        RECT 117.265 157.855 117.555 158.170 ;
        RECT 118.345 158.150 118.635 158.195 ;
        RECT 121.925 158.150 122.215 158.195 ;
        RECT 123.760 158.150 124.050 158.195 ;
        RECT 118.345 158.010 124.050 158.150 ;
        RECT 118.345 157.965 118.635 158.010 ;
        RECT 121.925 157.965 122.215 158.010 ;
        RECT 123.760 157.965 124.050 158.010 ;
        RECT 124.210 158.150 124.530 158.210 ;
        RECT 126.050 158.150 126.370 158.210 ;
        RECT 124.210 158.010 126.370 158.150 ;
        RECT 124.210 157.950 124.530 158.010 ;
        RECT 126.050 157.950 126.370 158.010 ;
        RECT 116.965 157.810 117.555 157.855 ;
        RECT 119.150 157.810 119.470 157.870 ;
        RECT 120.205 157.810 120.855 157.855 ;
        RECT 113.260 157.670 115.700 157.810 ;
        RECT 77.290 157.330 85.110 157.470 ;
        RECT 105.810 157.470 106.130 157.530 ;
        RECT 106.285 157.470 106.575 157.515 ;
        RECT 105.810 157.330 106.575 157.470 ;
        RECT 77.290 157.270 77.610 157.330 ;
        RECT 105.810 157.270 106.130 157.330 ;
        RECT 106.285 157.285 106.575 157.330 ;
        RECT 111.790 157.470 112.110 157.530 ;
        RECT 113.260 157.470 113.400 157.670 ;
        RECT 115.560 157.515 115.700 157.670 ;
        RECT 116.965 157.670 120.855 157.810 ;
        RECT 116.965 157.625 117.255 157.670 ;
        RECT 119.150 157.610 119.470 157.670 ;
        RECT 120.205 157.625 120.855 157.670 ;
        RECT 121.450 157.810 121.770 157.870 ;
        RECT 122.845 157.810 123.135 157.855 ;
        RECT 121.450 157.670 123.135 157.810 ;
        RECT 121.450 157.610 121.770 157.670 ;
        RECT 122.845 157.625 123.135 157.670 ;
        RECT 111.790 157.330 113.400 157.470 ;
        RECT 115.485 157.470 115.775 157.515 ;
        RECT 118.230 157.470 118.550 157.530 ;
        RECT 115.485 157.330 118.550 157.470 ;
        RECT 111.790 157.270 112.110 157.330 ;
        RECT 115.485 157.285 115.775 157.330 ;
        RECT 118.230 157.270 118.550 157.330 ;
        RECT 14.660 156.650 127.820 157.130 ;
        RECT 27.165 156.450 27.455 156.495 ;
        RECT 25.400 156.310 27.455 156.450 ;
        RECT 25.400 156.155 25.540 156.310 ;
        RECT 27.165 156.265 27.455 156.310 ;
        RECT 36.825 156.450 37.115 156.495 ;
        RECT 40.950 156.450 41.270 156.510 ;
        RECT 42.805 156.450 43.095 156.495 ;
        RECT 57.970 156.450 58.290 156.510 ;
        RECT 36.825 156.310 41.270 156.450 ;
        RECT 36.825 156.265 37.115 156.310 ;
        RECT 40.950 156.250 41.270 156.310 ;
        RECT 41.960 156.310 43.095 156.450 ;
        RECT 19.445 156.110 19.735 156.155 ;
        RECT 22.685 156.110 23.335 156.155 ;
        RECT 19.445 155.970 23.335 156.110 ;
        RECT 19.445 155.925 20.035 155.970 ;
        RECT 22.685 155.925 23.335 155.970 ;
        RECT 25.325 155.925 25.615 156.155 ;
        RECT 19.745 155.830 20.035 155.925 ;
        RECT 34.970 155.910 35.290 156.170 ;
        RECT 19.745 155.610 20.110 155.830 ;
        RECT 19.790 155.570 20.110 155.610 ;
        RECT 20.825 155.770 21.115 155.815 ;
        RECT 24.405 155.770 24.695 155.815 ;
        RECT 26.240 155.770 26.530 155.815 ;
        RECT 20.825 155.630 26.530 155.770 ;
        RECT 20.825 155.585 21.115 155.630 ;
        RECT 24.405 155.585 24.695 155.630 ;
        RECT 26.240 155.585 26.530 155.630 ;
        RECT 28.070 155.570 28.390 155.830 ;
        RECT 28.990 155.770 29.310 155.830 ;
        RECT 41.960 155.770 42.100 156.310 ;
        RECT 42.805 156.265 43.095 156.310 ;
        RECT 43.340 156.310 48.080 156.450 ;
        RECT 28.990 155.630 42.100 155.770 ;
        RECT 28.990 155.570 29.310 155.630 ;
        RECT 17.965 155.430 18.255 155.475 ;
        RECT 22.550 155.430 22.870 155.490 ;
        RECT 17.965 155.290 22.870 155.430 ;
        RECT 17.965 155.245 18.255 155.290 ;
        RECT 22.550 155.230 22.870 155.290 ;
        RECT 26.690 155.230 27.010 155.490 ;
        RECT 34.065 155.245 34.355 155.475 ;
        RECT 20.825 155.090 21.115 155.135 ;
        RECT 23.945 155.090 24.235 155.135 ;
        RECT 25.835 155.090 26.125 155.135 ;
        RECT 20.825 154.950 26.125 155.090 ;
        RECT 34.140 155.090 34.280 155.245 ;
        RECT 34.510 155.230 34.830 155.490 ;
        RECT 34.970 155.430 35.290 155.490 ;
        RECT 36.350 155.430 36.670 155.490 ;
        RECT 43.340 155.430 43.480 156.310 ;
        RECT 45.105 156.110 45.395 156.155 ;
        RECT 45.565 156.110 45.855 156.155 ;
        RECT 45.105 155.970 45.855 156.110 ;
        RECT 45.105 155.925 45.395 155.970 ;
        RECT 45.565 155.925 45.855 155.970 ;
        RECT 43.710 155.570 44.030 155.830 ;
        RECT 46.930 155.570 47.250 155.830 ;
        RECT 47.390 155.570 47.710 155.830 ;
        RECT 47.940 155.815 48.080 156.310 ;
        RECT 48.400 156.310 58.290 156.450 ;
        RECT 47.865 155.585 48.155 155.815 ;
        RECT 48.400 155.770 48.540 156.310 ;
        RECT 57.970 156.250 58.290 156.310 ;
        RECT 69.470 156.450 69.790 156.510 ;
        RECT 103.510 156.450 103.830 156.510 ;
        RECT 69.470 156.310 107.420 156.450 ;
        RECT 69.470 156.250 69.790 156.310 ;
        RECT 49.690 156.110 50.010 156.170 ;
        RECT 49.320 155.970 50.010 156.110 ;
        RECT 49.320 155.815 49.460 155.970 ;
        RECT 49.690 155.910 50.010 155.970 ;
        RECT 65.345 156.110 65.635 156.155 ;
        RECT 68.500 156.110 68.790 156.155 ;
        RECT 71.760 156.110 72.050 156.155 ;
        RECT 65.345 155.970 72.050 156.110 ;
        RECT 65.345 155.925 65.635 155.970 ;
        RECT 68.500 155.925 68.790 155.970 ;
        RECT 71.760 155.925 72.050 155.970 ;
        RECT 72.680 156.110 72.970 156.155 ;
        RECT 74.540 156.110 74.830 156.155 ;
        RECT 72.680 155.970 74.830 156.110 ;
        RECT 72.680 155.925 72.970 155.970 ;
        RECT 74.540 155.925 74.830 155.970 ;
        RECT 48.785 155.770 49.075 155.815 ;
        RECT 48.400 155.630 49.075 155.770 ;
        RECT 48.785 155.585 49.075 155.630 ;
        RECT 49.245 155.585 49.535 155.815 ;
        RECT 50.165 155.585 50.455 155.815 ;
        RECT 34.970 155.290 43.480 155.430 ;
        RECT 34.970 155.230 35.290 155.290 ;
        RECT 36.350 155.230 36.670 155.290 ;
        RECT 44.630 155.230 44.950 155.490 ;
        RECT 50.240 155.430 50.380 155.585 ;
        RECT 50.610 155.570 50.930 155.830 ;
        RECT 51.070 155.570 51.390 155.830 ;
        RECT 59.350 155.570 59.670 155.830 ;
        RECT 60.270 155.570 60.590 155.830 ;
        RECT 60.745 155.585 61.035 155.815 ;
        RECT 45.180 155.290 50.380 155.430 ;
        RECT 35.890 155.090 36.210 155.150 ;
        RECT 45.180 155.090 45.320 155.290 ;
        RECT 53.370 155.090 53.690 155.150 ;
        RECT 34.140 154.950 36.210 155.090 ;
        RECT 20.825 154.905 21.115 154.950 ;
        RECT 23.945 154.905 24.235 154.950 ;
        RECT 25.835 154.905 26.125 154.950 ;
        RECT 35.890 154.890 36.210 154.950 ;
        RECT 36.440 154.950 45.320 155.090 ;
        RECT 49.320 154.950 53.690 155.090 ;
        RECT 21.630 154.750 21.950 154.810 ;
        RECT 36.440 154.750 36.580 154.950 ;
        RECT 21.630 154.610 36.580 154.750 ;
        RECT 21.630 154.550 21.950 154.610 ;
        RECT 44.630 154.550 44.950 154.810 ;
        RECT 47.390 154.750 47.710 154.810 ;
        RECT 49.320 154.750 49.460 154.950 ;
        RECT 53.370 154.890 53.690 154.950 ;
        RECT 60.270 155.090 60.590 155.150 ;
        RECT 60.820 155.090 60.960 155.585 ;
        RECT 61.190 155.570 61.510 155.830 ;
        RECT 61.650 155.770 61.970 155.830 ;
        RECT 64.885 155.770 65.175 155.815 ;
        RECT 61.650 155.630 65.175 155.770 ;
        RECT 61.650 155.570 61.970 155.630 ;
        RECT 64.885 155.585 65.175 155.630 ;
        RECT 70.360 155.770 70.650 155.815 ;
        RECT 72.680 155.770 72.895 155.925 ;
        RECT 75.450 155.910 75.770 156.170 ;
        RECT 70.360 155.630 72.895 155.770 ;
        RECT 75.540 155.770 75.680 155.910 ;
        RECT 77.290 155.770 77.610 155.830 ;
        RECT 75.540 155.630 77.610 155.770 ;
        RECT 70.360 155.585 70.650 155.630 ;
        RECT 77.290 155.570 77.610 155.630 ;
        RECT 93.850 155.570 94.170 155.830 ;
        RECT 98.540 155.770 98.680 156.310 ;
        RECT 103.510 156.250 103.830 156.310 ;
        RECT 104.430 156.110 104.750 156.170 ;
        RECT 99.460 155.970 106.960 156.110 ;
        RECT 99.460 155.815 99.600 155.970 ;
        RECT 98.925 155.770 99.215 155.815 ;
        RECT 98.540 155.630 99.215 155.770 ;
        RECT 98.925 155.585 99.215 155.630 ;
        RECT 99.385 155.585 99.675 155.815 ;
        RECT 99.830 155.570 100.150 155.830 ;
        RECT 100.765 155.770 101.055 155.815 ;
        RECT 101.670 155.770 101.990 155.830 ;
        RECT 100.765 155.630 101.990 155.770 ;
        RECT 100.765 155.585 101.055 155.630 ;
        RECT 101.670 155.570 101.990 155.630 ;
        RECT 102.130 155.770 102.450 155.830 ;
        RECT 103.140 155.815 103.280 155.970 ;
        RECT 104.430 155.910 104.750 155.970 ;
        RECT 102.605 155.770 102.895 155.815 ;
        RECT 102.130 155.630 102.895 155.770 ;
        RECT 102.130 155.570 102.450 155.630 ;
        RECT 102.605 155.585 102.895 155.630 ;
        RECT 103.065 155.585 103.355 155.815 ;
        RECT 103.510 155.570 103.830 155.830 ;
        RECT 105.365 155.585 105.655 155.815 ;
        RECT 62.570 155.430 62.890 155.490 ;
        RECT 65.330 155.430 65.650 155.490 ;
        RECT 62.570 155.290 65.650 155.430 ;
        RECT 62.570 155.230 62.890 155.290 ;
        RECT 65.330 155.230 65.650 155.290 ;
        RECT 73.610 155.230 73.930 155.490 ;
        RECT 75.465 155.430 75.755 155.475 ;
        RECT 97.070 155.430 97.390 155.490 ;
        RECT 75.465 155.290 97.390 155.430 ;
        RECT 101.760 155.430 101.900 155.570 ;
        RECT 105.440 155.430 105.580 155.585 ;
        RECT 106.270 155.570 106.590 155.830 ;
        RECT 106.820 155.815 106.960 155.970 ;
        RECT 107.280 155.815 107.420 156.310 ;
        RECT 111.790 156.250 112.110 156.510 ;
        RECT 115.945 156.110 116.235 156.155 ;
        RECT 119.100 156.110 119.390 156.155 ;
        RECT 122.360 156.110 122.650 156.155 ;
        RECT 115.945 155.970 122.650 156.110 ;
        RECT 115.945 155.925 116.235 155.970 ;
        RECT 119.100 155.925 119.390 155.970 ;
        RECT 122.360 155.925 122.650 155.970 ;
        RECT 123.280 156.110 123.570 156.155 ;
        RECT 125.140 156.110 125.430 156.155 ;
        RECT 123.280 155.970 125.430 156.110 ;
        RECT 123.280 155.925 123.570 155.970 ;
        RECT 125.140 155.925 125.430 155.970 ;
        RECT 106.745 155.585 107.035 155.815 ;
        RECT 107.205 155.585 107.495 155.815 ;
        RECT 108.570 155.770 108.890 155.830 ;
        RECT 112.265 155.770 112.555 155.815 ;
        RECT 108.570 155.630 112.555 155.770 ;
        RECT 108.570 155.570 108.890 155.630 ;
        RECT 112.265 155.585 112.555 155.630 ;
        RECT 115.470 155.570 115.790 155.830 ;
        RECT 120.960 155.770 121.250 155.815 ;
        RECT 123.280 155.770 123.495 155.925 ;
        RECT 120.960 155.630 123.495 155.770 ;
        RECT 120.960 155.585 121.250 155.630 ;
        RECT 126.050 155.570 126.370 155.830 ;
        RECT 101.760 155.290 105.580 155.430 ;
        RECT 111.345 155.430 111.635 155.475 ;
        RECT 112.710 155.430 113.030 155.490 ;
        RECT 111.345 155.290 113.030 155.430 ;
        RECT 75.465 155.245 75.755 155.290 ;
        RECT 97.070 155.230 97.390 155.290 ;
        RECT 111.345 155.245 111.635 155.290 ;
        RECT 112.710 155.230 113.030 155.290 ;
        RECT 124.210 155.230 124.530 155.490 ;
        RECT 60.270 154.950 60.960 155.090 ;
        RECT 61.190 155.090 61.510 155.150 ;
        RECT 66.495 155.090 66.785 155.135 ;
        RECT 61.190 154.950 66.785 155.090 ;
        RECT 60.270 154.890 60.590 154.950 ;
        RECT 61.190 154.890 61.510 154.950 ;
        RECT 66.495 154.905 66.785 154.950 ;
        RECT 70.360 155.090 70.650 155.135 ;
        RECT 73.140 155.090 73.430 155.135 ;
        RECT 75.000 155.090 75.290 155.135 ;
        RECT 70.360 154.950 75.290 155.090 ;
        RECT 70.360 154.905 70.650 154.950 ;
        RECT 73.140 154.905 73.430 154.950 ;
        RECT 75.000 154.905 75.290 154.950 ;
        RECT 104.430 155.090 104.750 155.150 ;
        RECT 108.585 155.090 108.875 155.135 ;
        RECT 104.430 154.950 108.875 155.090 ;
        RECT 104.430 154.890 104.750 154.950 ;
        RECT 108.585 154.905 108.875 154.950 ;
        RECT 117.095 155.090 117.385 155.135 ;
        RECT 117.770 155.090 118.090 155.150 ;
        RECT 117.095 154.950 118.090 155.090 ;
        RECT 117.095 154.905 117.385 154.950 ;
        RECT 117.770 154.890 118.090 154.950 ;
        RECT 120.960 155.090 121.250 155.135 ;
        RECT 123.740 155.090 124.030 155.135 ;
        RECT 125.600 155.090 125.890 155.135 ;
        RECT 120.960 154.950 125.890 155.090 ;
        RECT 120.960 154.905 121.250 154.950 ;
        RECT 123.740 154.905 124.030 154.950 ;
        RECT 125.600 154.905 125.890 154.950 ;
        RECT 47.390 154.610 49.460 154.750 ;
        RECT 51.070 154.750 51.390 154.810 ;
        RECT 52.465 154.750 52.755 154.795 ;
        RECT 51.070 154.610 52.755 154.750 ;
        RECT 47.390 154.550 47.710 154.610 ;
        RECT 51.070 154.550 51.390 154.610 ;
        RECT 52.465 154.565 52.755 154.610 ;
        RECT 63.950 154.750 64.270 154.810 ;
        RECT 76.385 154.750 76.675 154.795 ;
        RECT 81.430 154.750 81.750 154.810 ;
        RECT 63.950 154.610 81.750 154.750 ;
        RECT 63.950 154.550 64.270 154.610 ;
        RECT 76.385 154.565 76.675 154.610 ;
        RECT 81.430 154.550 81.750 154.610 ;
        RECT 94.785 154.750 95.075 154.795 ;
        RECT 95.690 154.750 96.010 154.810 ;
        RECT 94.785 154.610 96.010 154.750 ;
        RECT 94.785 154.565 95.075 154.610 ;
        RECT 95.690 154.550 96.010 154.610 ;
        RECT 97.530 154.550 97.850 154.810 ;
        RECT 104.890 154.550 105.210 154.810 ;
        RECT 114.105 154.750 114.395 154.795 ;
        RECT 118.690 154.750 119.010 154.810 ;
        RECT 114.105 154.610 119.010 154.750 ;
        RECT 114.105 154.565 114.395 154.610 ;
        RECT 118.690 154.550 119.010 154.610 ;
        RECT 14.660 153.930 127.820 154.410 ;
        RECT 23.945 153.730 24.235 153.775 ;
        RECT 28.070 153.730 28.390 153.790 ;
        RECT 23.945 153.590 28.390 153.730 ;
        RECT 23.945 153.545 24.235 153.590 ;
        RECT 28.070 153.530 28.390 153.590 ;
        RECT 39.125 153.545 39.415 153.775 ;
        RECT 39.200 153.110 39.340 153.545 ;
        RECT 45.090 153.530 45.410 153.790 ;
        RECT 50.150 153.730 50.470 153.790 ;
        RECT 48.860 153.590 50.470 153.730 ;
        RECT 43.725 153.205 44.015 153.435 ;
        RECT 48.860 153.390 49.000 153.590 ;
        RECT 50.150 153.530 50.470 153.590 ;
        RECT 50.625 153.730 50.915 153.775 ;
        RECT 53.370 153.730 53.690 153.790 ;
        RECT 73.150 153.730 73.470 153.790 ;
        RECT 75.005 153.730 75.295 153.775 ;
        RECT 50.625 153.590 53.140 153.730 ;
        RECT 50.625 153.545 50.915 153.590 ;
        RECT 45.180 153.250 49.000 153.390 ;
        RECT 21.170 152.850 21.490 153.110 ;
        RECT 36.350 152.850 36.670 153.110 ;
        RECT 39.110 152.850 39.430 153.110 ;
        RECT 39.570 153.050 39.890 153.110 ;
        RECT 43.800 153.050 43.940 153.205 ;
        RECT 45.180 153.050 45.320 153.250 ;
        RECT 49.690 153.190 50.010 153.450 ;
        RECT 53.000 153.390 53.140 153.590 ;
        RECT 53.370 153.590 71.080 153.730 ;
        RECT 53.370 153.530 53.690 153.590 ;
        RECT 70.940 153.450 71.080 153.590 ;
        RECT 73.150 153.590 75.295 153.730 ;
        RECT 73.150 153.530 73.470 153.590 ;
        RECT 75.005 153.545 75.295 153.590 ;
        RECT 75.910 153.730 76.230 153.790 ;
        RECT 76.845 153.730 77.135 153.775 ;
        RECT 117.770 153.730 118.090 153.790 ;
        RECT 75.910 153.590 77.135 153.730 ;
        RECT 75.910 153.530 76.230 153.590 ;
        RECT 76.845 153.545 77.135 153.590 ;
        RECT 112.340 153.590 118.090 153.730 ;
        RECT 54.290 153.390 54.610 153.450 ;
        RECT 70.850 153.390 71.170 153.450 ;
        RECT 79.130 153.390 79.450 153.450 ;
        RECT 53.000 153.250 54.610 153.390 ;
        RECT 54.290 153.190 54.610 153.250 ;
        RECT 66.800 153.250 70.620 153.390 ;
        RECT 66.800 153.110 66.940 153.250 ;
        RECT 39.570 152.910 43.940 153.050 ;
        RECT 44.720 152.910 45.320 153.050 ;
        RECT 39.570 152.850 39.890 152.910 ;
        RECT 36.810 152.510 37.130 152.770 ;
        RECT 44.720 152.755 44.860 152.910 ;
        RECT 45.550 152.850 45.870 153.110 ;
        RECT 58.445 153.050 58.735 153.095 ;
        RECT 46.100 152.910 58.735 153.050 ;
        RECT 46.100 152.755 46.240 152.910 ;
        RECT 58.445 152.865 58.735 152.910 ;
        RECT 64.870 153.050 65.190 153.110 ;
        RECT 66.265 153.050 66.555 153.095 ;
        RECT 66.710 153.050 67.030 153.110 ;
        RECT 64.870 152.910 67.030 153.050 ;
        RECT 64.870 152.850 65.190 152.910 ;
        RECT 66.265 152.865 66.555 152.910 ;
        RECT 66.710 152.850 67.030 152.910 ;
        RECT 67.630 153.050 67.950 153.110 ;
        RECT 70.480 153.050 70.620 153.250 ;
        RECT 70.850 153.250 79.450 153.390 ;
        RECT 70.850 153.190 71.170 153.250 ;
        RECT 79.130 153.190 79.450 153.250 ;
        RECT 91.205 153.390 91.495 153.435 ;
        RECT 94.325 153.390 94.615 153.435 ;
        RECT 96.215 153.390 96.505 153.435 ;
        RECT 91.205 153.250 96.505 153.390 ;
        RECT 91.205 153.205 91.495 153.250 ;
        RECT 94.325 153.205 94.615 153.250 ;
        RECT 96.215 153.205 96.505 153.250 ;
        RECT 103.510 153.190 103.830 153.450 ;
        RECT 112.340 153.390 112.480 153.590 ;
        RECT 117.770 153.530 118.090 153.590 ;
        RECT 121.450 153.530 121.770 153.790 ;
        RECT 122.845 153.730 123.135 153.775 ;
        RECT 124.210 153.730 124.530 153.790 ;
        RECT 122.845 153.590 124.530 153.730 ;
        RECT 122.845 153.545 123.135 153.590 ;
        RECT 124.210 153.530 124.530 153.590 ;
        RECT 111.880 153.250 112.480 153.390 ;
        RECT 112.710 153.390 113.030 153.450 ;
        RECT 112.710 153.250 117.080 153.390 ;
        RECT 71.325 153.050 71.615 153.095 ;
        RECT 67.630 152.910 70.160 153.050 ;
        RECT 70.480 152.910 71.615 153.050 ;
        RECT 67.630 152.850 67.950 152.910 ;
        RECT 44.645 152.525 44.935 152.755 ;
        RECT 46.025 152.525 46.315 152.755 ;
        RECT 46.485 152.710 46.775 152.755 ;
        RECT 46.930 152.710 47.250 152.770 ;
        RECT 46.485 152.570 47.250 152.710 ;
        RECT 46.485 152.525 46.775 152.570 ;
        RECT 46.930 152.510 47.250 152.570 ;
        RECT 47.405 152.525 47.695 152.755 ;
        RECT 47.865 152.525 48.155 152.755 ;
        RECT 48.325 152.710 48.615 152.755 ;
        RECT 49.230 152.710 49.550 152.770 ;
        RECT 52.005 152.710 52.295 152.755 ;
        RECT 48.325 152.570 52.295 152.710 ;
        RECT 48.325 152.525 48.615 152.570 ;
        RECT 21.645 152.370 21.935 152.415 ;
        RECT 22.550 152.370 22.870 152.430 ;
        RECT 47.480 152.370 47.620 152.525 ;
        RECT 21.645 152.230 47.620 152.370 ;
        RECT 47.940 152.370 48.080 152.525 ;
        RECT 49.230 152.510 49.550 152.570 ;
        RECT 52.005 152.525 52.295 152.570 ;
        RECT 52.465 152.525 52.755 152.755 ;
        RECT 52.925 152.525 53.215 152.755 ;
        RECT 50.150 152.370 50.470 152.430 ;
        RECT 52.540 152.370 52.680 152.525 ;
        RECT 47.940 152.230 52.680 152.370 ;
        RECT 21.645 152.185 21.935 152.230 ;
        RECT 22.550 152.170 22.870 152.230 ;
        RECT 50.150 152.170 50.470 152.230 ;
        RECT 22.090 151.830 22.410 152.090 ;
        RECT 34.510 152.030 34.830 152.090 ;
        RECT 37.285 152.030 37.575 152.075 ;
        RECT 49.230 152.030 49.550 152.090 ;
        RECT 34.510 151.890 49.550 152.030 ;
        RECT 53.000 152.030 53.140 152.525 ;
        RECT 53.830 152.510 54.150 152.770 ;
        RECT 59.810 152.510 60.130 152.770 ;
        RECT 60.270 152.510 60.590 152.770 ;
        RECT 60.730 152.510 61.050 152.770 ;
        RECT 61.650 152.710 61.970 152.770 ;
        RECT 63.950 152.710 64.270 152.770 ;
        RECT 69.485 152.710 69.775 152.755 ;
        RECT 61.650 152.570 64.270 152.710 ;
        RECT 61.650 152.510 61.970 152.570 ;
        RECT 63.950 152.510 64.270 152.570 ;
        RECT 69.100 152.570 69.775 152.710 ;
        RECT 70.020 152.710 70.160 152.910 ;
        RECT 71.325 152.865 71.615 152.910 ;
        RECT 72.320 152.910 76.600 153.050 ;
        RECT 70.850 152.710 71.170 152.770 ;
        RECT 72.320 152.710 72.460 152.910 ;
        RECT 70.020 152.570 72.460 152.710 ;
        RECT 74.085 152.710 74.375 152.755 ;
        RECT 75.450 152.710 75.770 152.770 ;
        RECT 76.460 152.755 76.600 152.910 ;
        RECT 77.750 152.850 78.070 153.110 ;
        RECT 95.690 152.850 96.010 153.110 ;
        RECT 97.070 152.850 97.390 153.110 ;
        RECT 103.600 153.050 103.740 153.190 ;
        RECT 103.600 152.910 104.660 153.050 ;
        RECT 74.085 152.570 75.770 152.710 ;
        RECT 60.820 152.370 60.960 152.510 ;
        RECT 66.725 152.370 67.015 152.415 ;
        RECT 60.820 152.230 67.015 152.370 ;
        RECT 66.725 152.185 67.015 152.230 ;
        RECT 53.830 152.030 54.150 152.090 ;
        RECT 53.000 151.890 54.150 152.030 ;
        RECT 34.510 151.830 34.830 151.890 ;
        RECT 37.285 151.845 37.575 151.890 ;
        RECT 49.230 151.830 49.550 151.890 ;
        RECT 53.830 151.830 54.150 151.890 ;
        RECT 66.250 152.030 66.570 152.090 ;
        RECT 69.100 152.075 69.240 152.570 ;
        RECT 69.485 152.525 69.775 152.570 ;
        RECT 70.850 152.510 71.170 152.570 ;
        RECT 74.085 152.525 74.375 152.570 ;
        RECT 75.450 152.510 75.770 152.570 ;
        RECT 76.385 152.525 76.675 152.755 ;
        RECT 77.290 152.710 77.610 152.770 ;
        RECT 78.225 152.710 78.515 152.755 ;
        RECT 77.290 152.570 78.515 152.710 ;
        RECT 77.290 152.510 77.610 152.570 ;
        RECT 78.225 152.525 78.515 152.570 ;
        RECT 86.950 152.510 87.270 152.770 ;
        RECT 72.705 152.370 72.995 152.415 ;
        RECT 78.685 152.370 78.975 152.415 ;
        RECT 82.365 152.370 82.655 152.415 ;
        RECT 72.705 152.230 82.655 152.370 ;
        RECT 72.705 152.185 72.995 152.230 ;
        RECT 78.685 152.185 78.975 152.230 ;
        RECT 82.365 152.185 82.655 152.230 ;
        RECT 84.205 152.370 84.495 152.415 ;
        RECT 86.490 152.370 86.810 152.430 ;
        RECT 90.125 152.415 90.415 152.730 ;
        RECT 91.205 152.710 91.495 152.755 ;
        RECT 94.785 152.710 95.075 152.755 ;
        RECT 96.620 152.710 96.910 152.755 ;
        RECT 91.205 152.570 96.910 152.710 ;
        RECT 91.205 152.525 91.495 152.570 ;
        RECT 94.785 152.525 95.075 152.570 ;
        RECT 96.620 152.525 96.910 152.570 ;
        RECT 101.670 152.710 101.990 152.770 ;
        RECT 102.605 152.710 102.895 152.755 ;
        RECT 101.670 152.570 102.895 152.710 ;
        RECT 101.670 152.510 101.990 152.570 ;
        RECT 102.605 152.525 102.895 152.570 ;
        RECT 103.050 152.710 103.370 152.770 ;
        RECT 103.525 152.710 103.815 152.755 ;
        RECT 103.050 152.570 103.815 152.710 ;
        RECT 103.050 152.510 103.370 152.570 ;
        RECT 103.525 152.525 103.815 152.570 ;
        RECT 103.970 152.510 104.290 152.770 ;
        RECT 104.520 152.755 104.660 152.910 ;
        RECT 104.980 152.910 108.340 153.050 ;
        RECT 104.445 152.525 104.735 152.755 ;
        RECT 84.205 152.230 86.810 152.370 ;
        RECT 84.205 152.185 84.495 152.230 ;
        RECT 86.490 152.170 86.810 152.230 ;
        RECT 87.425 152.370 87.715 152.415 ;
        RECT 89.825 152.370 90.415 152.415 ;
        RECT 93.065 152.370 93.715 152.415 ;
        RECT 87.425 152.230 93.715 152.370 ;
        RECT 87.425 152.185 87.715 152.230 ;
        RECT 89.825 152.185 90.115 152.230 ;
        RECT 93.065 152.185 93.715 152.230 ;
        RECT 99.830 152.370 100.150 152.430 ;
        RECT 104.980 152.370 105.120 152.910 ;
        RECT 107.650 152.510 107.970 152.770 ;
        RECT 108.200 152.755 108.340 152.910 ;
        RECT 108.125 152.525 108.415 152.755 ;
        RECT 108.570 152.510 108.890 152.770 ;
        RECT 109.505 152.710 109.795 152.755 ;
        RECT 110.885 152.710 111.175 152.755 ;
        RECT 111.330 152.710 111.650 152.770 ;
        RECT 111.880 152.755 112.020 153.250 ;
        RECT 112.710 153.190 113.030 153.250 ;
        RECT 116.940 153.095 117.080 153.250 ;
        RECT 116.865 152.865 117.155 153.095 ;
        RECT 109.505 152.570 111.650 152.710 ;
        RECT 109.505 152.525 109.795 152.570 ;
        RECT 110.885 152.525 111.175 152.570 ;
        RECT 111.330 152.510 111.650 152.570 ;
        RECT 111.805 152.525 112.095 152.755 ;
        RECT 112.250 152.510 112.570 152.770 ;
        RECT 112.725 152.525 113.015 152.755 ;
        RECT 99.830 152.230 105.120 152.370 ;
        RECT 99.830 152.170 100.150 152.230 ;
        RECT 105.810 152.170 106.130 152.430 ;
        RECT 107.740 152.370 107.880 152.510 ;
        RECT 112.800 152.370 112.940 152.525 ;
        RECT 118.230 152.510 118.550 152.770 ;
        RECT 118.690 152.710 119.010 152.770 ;
        RECT 120.545 152.710 120.835 152.755 ;
        RECT 118.690 152.570 120.835 152.710 ;
        RECT 118.690 152.510 119.010 152.570 ;
        RECT 120.545 152.525 120.835 152.570 ;
        RECT 121.925 152.525 122.215 152.755 ;
        RECT 113.170 152.370 113.490 152.430 ;
        RECT 122.000 152.370 122.140 152.525 ;
        RECT 107.740 152.230 113.490 152.370 ;
        RECT 113.170 152.170 113.490 152.230 ;
        RECT 120.160 152.230 122.140 152.370 ;
        RECT 67.185 152.030 67.475 152.075 ;
        RECT 66.250 151.890 67.475 152.030 ;
        RECT 66.250 151.830 66.570 151.890 ;
        RECT 67.185 151.845 67.475 151.890 ;
        RECT 69.025 151.845 69.315 152.075 ;
        RECT 70.405 152.030 70.695 152.075 ;
        RECT 73.610 152.030 73.930 152.090 ;
        RECT 70.405 151.890 73.930 152.030 ;
        RECT 70.405 151.845 70.695 151.890 ;
        RECT 73.610 151.830 73.930 151.890 ;
        RECT 74.990 152.030 75.310 152.090 ;
        RECT 77.750 152.030 78.070 152.090 ;
        RECT 74.990 151.890 78.070 152.030 ;
        RECT 74.990 151.830 75.310 151.890 ;
        RECT 77.750 151.830 78.070 151.890 ;
        RECT 88.330 151.830 88.650 152.090 ;
        RECT 103.970 152.030 104.290 152.090 ;
        RECT 106.285 152.030 106.575 152.075 ;
        RECT 103.970 151.890 106.575 152.030 ;
        RECT 103.970 151.830 104.290 151.890 ;
        RECT 106.285 151.845 106.575 151.890 ;
        RECT 114.090 151.830 114.410 152.090 ;
        RECT 117.785 152.030 118.075 152.075 ;
        RECT 118.230 152.030 118.550 152.090 ;
        RECT 120.160 152.075 120.300 152.230 ;
        RECT 117.785 151.890 118.550 152.030 ;
        RECT 117.785 151.845 118.075 151.890 ;
        RECT 118.230 151.830 118.550 151.890 ;
        RECT 120.085 151.845 120.375 152.075 ;
        RECT 14.660 151.210 127.820 151.690 ;
        RECT 24.390 151.010 24.710 151.070 ;
        RECT 46.485 151.010 46.775 151.055 ;
        RECT 49.245 151.010 49.535 151.055 ;
        RECT 54.765 151.010 55.055 151.055 ;
        RECT 24.390 150.870 46.775 151.010 ;
        RECT 24.390 150.810 24.710 150.870 ;
        RECT 46.485 150.825 46.775 150.870 ;
        RECT 47.020 150.870 49.535 151.010 ;
        RECT 18.065 150.670 18.355 150.715 ;
        RECT 18.870 150.670 19.190 150.730 ;
        RECT 21.305 150.670 21.955 150.715 ;
        RECT 18.065 150.530 21.955 150.670 ;
        RECT 18.065 150.485 18.655 150.530 ;
        RECT 18.365 150.170 18.655 150.485 ;
        RECT 18.870 150.470 19.190 150.530 ;
        RECT 21.305 150.485 21.955 150.530 ;
        RECT 31.745 150.670 32.395 150.715 ;
        RECT 34.510 150.670 34.830 150.730 ;
        RECT 35.345 150.670 35.635 150.715 ;
        RECT 31.745 150.530 35.635 150.670 ;
        RECT 31.745 150.485 32.395 150.530 ;
        RECT 34.510 150.470 34.830 150.530 ;
        RECT 35.045 150.485 35.635 150.530 ;
        RECT 43.710 150.670 44.030 150.730 ;
        RECT 47.020 150.670 47.160 150.870 ;
        RECT 49.245 150.825 49.535 150.870 ;
        RECT 51.160 150.870 55.055 151.010 ;
        RECT 43.710 150.530 47.160 150.670 ;
        RECT 48.785 150.670 49.075 150.715 ;
        RECT 51.160 150.670 51.300 150.870 ;
        RECT 54.765 150.825 55.055 150.870 ;
        RECT 56.130 151.010 56.450 151.070 ;
        RECT 59.810 151.010 60.130 151.070 ;
        RECT 73.165 151.010 73.455 151.055 ;
        RECT 92.945 151.010 93.235 151.055 ;
        RECT 93.850 151.010 94.170 151.070 ;
        RECT 109.030 151.010 109.350 151.070 ;
        RECT 56.130 150.870 85.110 151.010 ;
        RECT 56.130 150.810 56.450 150.870 ;
        RECT 59.810 150.810 60.130 150.870 ;
        RECT 73.165 150.825 73.455 150.870 ;
        RECT 48.785 150.530 51.300 150.670 ;
        RECT 51.545 150.670 51.835 150.715 ;
        RECT 58.445 150.670 58.735 150.715 ;
        RECT 74.530 150.670 74.850 150.730 ;
        RECT 79.130 150.670 79.450 150.730 ;
        RECT 51.545 150.530 58.735 150.670 ;
        RECT 19.445 150.330 19.735 150.375 ;
        RECT 23.025 150.330 23.315 150.375 ;
        RECT 24.860 150.330 25.150 150.375 ;
        RECT 19.445 150.190 25.150 150.330 ;
        RECT 19.445 150.145 19.735 150.190 ;
        RECT 23.025 150.145 23.315 150.190 ;
        RECT 24.860 150.145 25.150 150.190 ;
        RECT 28.550 150.330 28.840 150.375 ;
        RECT 30.385 150.330 30.675 150.375 ;
        RECT 33.965 150.330 34.255 150.375 ;
        RECT 28.550 150.190 34.255 150.330 ;
        RECT 28.550 150.145 28.840 150.190 ;
        RECT 30.385 150.145 30.675 150.190 ;
        RECT 33.965 150.145 34.255 150.190 ;
        RECT 35.045 150.170 35.335 150.485 ;
        RECT 43.710 150.470 44.030 150.530 ;
        RECT 48.785 150.485 49.075 150.530 ;
        RECT 51.545 150.485 51.835 150.530 ;
        RECT 58.445 150.485 58.735 150.530 ;
        RECT 59.440 150.530 61.880 150.670 ;
        RECT 39.110 150.330 39.430 150.390 ;
        RECT 39.585 150.330 39.875 150.375 ;
        RECT 39.110 150.190 39.875 150.330 ;
        RECT 39.110 150.130 39.430 150.190 ;
        RECT 39.585 150.145 39.875 150.190 ;
        RECT 46.470 150.330 46.790 150.390 ;
        RECT 47.405 150.330 47.695 150.375 ;
        RECT 46.470 150.190 47.695 150.330 ;
        RECT 46.470 150.130 46.790 150.190 ;
        RECT 47.405 150.145 47.695 150.190 ;
        RECT 50.165 150.330 50.455 150.375 ;
        RECT 51.990 150.330 52.310 150.390 ;
        RECT 50.165 150.190 52.310 150.330 ;
        RECT 50.165 150.145 50.455 150.190 ;
        RECT 51.990 150.130 52.310 150.190 ;
        RECT 56.130 150.130 56.450 150.390 ;
        RECT 56.605 150.145 56.895 150.375 ;
        RECT 57.065 150.330 57.355 150.375 ;
        RECT 57.510 150.330 57.830 150.390 ;
        RECT 57.065 150.190 57.830 150.330 ;
        RECT 57.065 150.145 57.355 150.190 ;
        RECT 20.710 149.990 21.030 150.050 ;
        RECT 23.945 149.990 24.235 150.035 ;
        RECT 20.710 149.850 24.235 149.990 ;
        RECT 20.710 149.790 21.030 149.850 ;
        RECT 23.945 149.805 24.235 149.850 ;
        RECT 25.325 149.990 25.615 150.035 ;
        RECT 26.690 149.990 27.010 150.050 ;
        RECT 28.070 149.990 28.390 150.050 ;
        RECT 25.325 149.850 28.390 149.990 ;
        RECT 25.325 149.805 25.615 149.850 ;
        RECT 26.690 149.790 27.010 149.850 ;
        RECT 28.070 149.790 28.390 149.850 ;
        RECT 29.465 149.990 29.755 150.035 ;
        RECT 29.465 149.850 38.880 149.990 ;
        RECT 29.465 149.805 29.755 149.850 ;
        RECT 38.740 149.695 38.880 149.850 ;
        RECT 48.325 149.805 48.615 150.035 ;
        RECT 19.445 149.650 19.735 149.695 ;
        RECT 22.565 149.650 22.855 149.695 ;
        RECT 24.455 149.650 24.745 149.695 ;
        RECT 19.445 149.510 24.745 149.650 ;
        RECT 19.445 149.465 19.735 149.510 ;
        RECT 22.565 149.465 22.855 149.510 ;
        RECT 24.455 149.465 24.745 149.510 ;
        RECT 28.955 149.650 29.245 149.695 ;
        RECT 30.845 149.650 31.135 149.695 ;
        RECT 33.965 149.650 34.255 149.695 ;
        RECT 28.955 149.510 34.255 149.650 ;
        RECT 28.955 149.465 29.245 149.510 ;
        RECT 30.845 149.465 31.135 149.510 ;
        RECT 33.965 149.465 34.255 149.510 ;
        RECT 38.665 149.465 38.955 149.695 ;
        RECT 48.400 149.650 48.540 149.805 ;
        RECT 51.070 149.790 51.390 150.050 ;
        RECT 56.680 149.990 56.820 150.145 ;
        RECT 57.510 150.130 57.830 150.190 ;
        RECT 57.970 150.330 58.290 150.390 ;
        RECT 59.440 150.330 59.580 150.530 ;
        RECT 61.740 150.390 61.880 150.530 ;
        RECT 74.530 150.530 77.980 150.670 ;
        RECT 74.530 150.470 74.850 150.530 ;
        RECT 57.970 150.190 59.580 150.330 ;
        RECT 57.970 150.130 58.290 150.190 ;
        RECT 59.810 150.130 60.130 150.390 ;
        RECT 60.270 150.130 60.590 150.390 ;
        RECT 60.745 150.145 61.035 150.375 ;
        RECT 60.360 149.990 60.500 150.130 ;
        RECT 56.680 149.850 60.500 149.990 ;
        RECT 60.820 149.990 60.960 150.145 ;
        RECT 61.650 150.130 61.970 150.390 ;
        RECT 72.230 150.130 72.550 150.390 ;
        RECT 74.085 150.145 74.375 150.375 ;
        RECT 66.250 149.990 66.570 150.050 ;
        RECT 60.820 149.850 66.570 149.990 ;
        RECT 54.290 149.650 54.610 149.710 ;
        RECT 48.400 149.510 54.610 149.650 ;
        RECT 60.360 149.650 60.500 149.850 ;
        RECT 66.250 149.790 66.570 149.850 ;
        RECT 70.850 149.990 71.170 150.050 ;
        RECT 74.160 149.990 74.300 150.145 ;
        RECT 75.910 150.130 76.230 150.390 ;
        RECT 76.845 150.330 77.135 150.375 ;
        RECT 77.290 150.330 77.610 150.390 ;
        RECT 77.840 150.375 77.980 150.530 ;
        RECT 78.300 150.530 82.580 150.670 ;
        RECT 78.300 150.375 78.440 150.530 ;
        RECT 79.130 150.470 79.450 150.530 ;
        RECT 76.845 150.190 77.610 150.330 ;
        RECT 76.845 150.145 77.135 150.190 ;
        RECT 77.290 150.130 77.610 150.190 ;
        RECT 77.765 150.145 78.055 150.375 ;
        RECT 78.225 150.145 78.515 150.375 ;
        RECT 78.685 150.330 78.975 150.375 ;
        RECT 80.510 150.330 80.830 150.390 ;
        RECT 82.440 150.375 82.580 150.530 ;
        RECT 81.905 150.330 82.195 150.375 ;
        RECT 78.685 150.190 82.195 150.330 ;
        RECT 78.685 150.145 78.975 150.190 ;
        RECT 80.510 150.130 80.830 150.190 ;
        RECT 81.905 150.145 82.195 150.190 ;
        RECT 82.365 150.145 82.655 150.375 ;
        RECT 82.825 150.330 83.115 150.375 ;
        RECT 83.270 150.330 83.590 150.390 ;
        RECT 82.825 150.190 83.590 150.330 ;
        RECT 82.825 150.145 83.115 150.190 ;
        RECT 83.270 150.130 83.590 150.190 ;
        RECT 83.730 150.130 84.050 150.390 ;
        RECT 84.970 150.330 85.110 150.870 ;
        RECT 92.945 150.870 94.170 151.010 ;
        RECT 92.945 150.825 93.235 150.870 ;
        RECT 93.850 150.810 94.170 150.870 ;
        RECT 99.920 150.870 109.350 151.010 ;
        RECT 88.330 150.670 88.650 150.730 ;
        RECT 90.645 150.670 90.935 150.715 ;
        RECT 99.920 150.670 100.060 150.870 ;
        RECT 109.030 150.810 109.350 150.870 ;
        RECT 111.805 151.010 112.095 151.055 ;
        RECT 114.550 151.010 114.870 151.070 ;
        RECT 111.805 150.870 114.870 151.010 ;
        RECT 111.805 150.825 112.095 150.870 ;
        RECT 114.550 150.810 114.870 150.870 ;
        RECT 88.330 150.530 100.060 150.670 ;
        RECT 88.330 150.470 88.650 150.530 ;
        RECT 90.645 150.485 90.935 150.530 ;
        RECT 103.970 150.470 104.290 150.730 ;
        RECT 109.505 150.670 109.795 150.715 ;
        RECT 114.090 150.670 114.410 150.730 ;
        RECT 109.505 150.530 114.410 150.670 ;
        RECT 109.505 150.485 109.795 150.530 ;
        RECT 114.090 150.470 114.410 150.530 ;
        RECT 84.970 150.190 90.860 150.330 ;
        RECT 70.850 149.850 74.300 149.990 ;
        RECT 86.490 149.990 86.810 150.050 ;
        RECT 89.725 149.990 90.015 150.035 ;
        RECT 86.490 149.850 90.015 149.990 ;
        RECT 90.720 149.990 90.860 150.190 ;
        RECT 91.090 150.130 91.410 150.390 ;
        RECT 105.350 150.130 105.670 150.390 ;
        RECT 105.810 150.330 106.130 150.390 ;
        RECT 110.425 150.330 110.715 150.375 ;
        RECT 105.810 150.190 110.715 150.330 ;
        RECT 105.810 150.130 106.130 150.190 ;
        RECT 110.425 150.145 110.715 150.190 ;
        RECT 110.870 150.130 111.190 150.390 ;
        RECT 99.370 149.990 99.690 150.050 ;
        RECT 90.720 149.850 99.690 149.990 ;
        RECT 70.850 149.790 71.170 149.850 ;
        RECT 86.490 149.790 86.810 149.850 ;
        RECT 89.725 149.805 90.015 149.850 ;
        RECT 99.370 149.790 99.690 149.850 ;
        RECT 104.430 149.790 104.750 150.050 ;
        RECT 111.330 149.990 111.650 150.050 ;
        RECT 113.630 149.990 113.950 150.050 ;
        RECT 105.900 149.850 113.950 149.990 ;
        RECT 78.670 149.650 78.990 149.710 ;
        RECT 80.525 149.650 80.815 149.695 ;
        RECT 60.360 149.510 75.220 149.650 ;
        RECT 54.290 149.450 54.610 149.510 ;
        RECT 16.585 149.310 16.875 149.355 ;
        RECT 22.090 149.310 22.410 149.370 ;
        RECT 16.585 149.170 22.410 149.310 ;
        RECT 16.585 149.125 16.875 149.170 ;
        RECT 22.090 149.110 22.410 149.170 ;
        RECT 36.810 149.110 37.130 149.370 ;
        RECT 48.785 149.310 49.075 149.355 ;
        RECT 49.230 149.310 49.550 149.370 ;
        RECT 48.785 149.170 49.550 149.310 ;
        RECT 48.785 149.125 49.075 149.170 ;
        RECT 49.230 149.110 49.550 149.170 ;
        RECT 50.610 149.110 50.930 149.370 ;
        RECT 64.870 149.110 65.190 149.370 ;
        RECT 75.080 149.355 75.220 149.510 ;
        RECT 78.670 149.510 80.815 149.650 ;
        RECT 78.670 149.450 78.990 149.510 ;
        RECT 80.525 149.465 80.815 149.510 ;
        RECT 80.970 149.450 81.290 149.710 ;
        RECT 81.430 149.650 81.750 149.710 ;
        RECT 101.210 149.650 101.530 149.710 ;
        RECT 105.900 149.650 106.040 149.850 ;
        RECT 111.330 149.790 111.650 149.850 ;
        RECT 113.630 149.790 113.950 149.850 ;
        RECT 81.430 149.510 106.040 149.650 ;
        RECT 106.285 149.650 106.575 149.695 ;
        RECT 120.990 149.650 121.310 149.710 ;
        RECT 106.285 149.510 121.310 149.650 ;
        RECT 81.430 149.450 81.750 149.510 ;
        RECT 101.210 149.450 101.530 149.510 ;
        RECT 106.285 149.465 106.575 149.510 ;
        RECT 120.990 149.450 121.310 149.510 ;
        RECT 75.005 149.310 75.295 149.355 ;
        RECT 76.830 149.310 77.150 149.370 ;
        RECT 75.005 149.170 77.150 149.310 ;
        RECT 75.005 149.125 75.295 149.170 ;
        RECT 76.830 149.110 77.150 149.170 ;
        RECT 80.065 149.310 80.355 149.355 ;
        RECT 81.060 149.310 81.200 149.450 ;
        RECT 80.065 149.170 81.200 149.310 ;
        RECT 82.350 149.310 82.670 149.370 ;
        RECT 99.830 149.310 100.150 149.370 ;
        RECT 82.350 149.170 100.150 149.310 ;
        RECT 80.065 149.125 80.355 149.170 ;
        RECT 82.350 149.110 82.670 149.170 ;
        RECT 99.830 149.110 100.150 149.170 ;
        RECT 103.970 149.110 104.290 149.370 ;
        RECT 110.885 149.310 111.175 149.355 ;
        RECT 111.790 149.310 112.110 149.370 ;
        RECT 110.885 149.170 112.110 149.310 ;
        RECT 110.885 149.125 111.175 149.170 ;
        RECT 111.790 149.110 112.110 149.170 ;
        RECT 14.660 148.490 127.820 148.970 ;
        RECT 18.870 148.290 19.190 148.350 ;
        RECT 19.345 148.290 19.635 148.335 ;
        RECT 18.870 148.150 19.635 148.290 ;
        RECT 18.870 148.090 19.190 148.150 ;
        RECT 19.345 148.105 19.635 148.150 ;
        RECT 33.145 148.290 33.435 148.335 ;
        RECT 34.510 148.290 34.830 148.350 ;
        RECT 33.145 148.150 34.830 148.290 ;
        RECT 33.145 148.105 33.435 148.150 ;
        RECT 34.510 148.090 34.830 148.150 ;
        RECT 77.305 148.290 77.595 148.335 ;
        RECT 85.570 148.290 85.890 148.350 ;
        RECT 77.305 148.150 85.890 148.290 ;
        RECT 77.305 148.105 77.595 148.150 ;
        RECT 85.570 148.090 85.890 148.150 ;
        RECT 97.545 148.290 97.835 148.335 ;
        RECT 97.990 148.290 98.310 148.350 ;
        RECT 97.545 148.150 98.310 148.290 ;
        RECT 97.545 148.105 97.835 148.150 ;
        RECT 97.990 148.090 98.310 148.150 ;
        RECT 109.030 148.090 109.350 148.350 ;
        RECT 49.690 147.950 50.010 148.010 ;
        RECT 73.150 147.950 73.470 148.010 ;
        RECT 83.730 147.950 84.050 148.010 ;
        RECT 49.690 147.810 77.520 147.950 ;
        RECT 49.690 147.750 50.010 147.810 ;
        RECT 73.150 147.750 73.470 147.810 ;
        RECT 77.380 147.670 77.520 147.810 ;
        RECT 78.760 147.810 84.050 147.950 ;
        RECT 21.170 147.410 21.490 147.670 ;
        RECT 75.450 147.610 75.770 147.670 ;
        RECT 77.290 147.610 77.610 147.670 ;
        RECT 78.760 147.610 78.900 147.810 ;
        RECT 83.730 147.750 84.050 147.810 ;
        RECT 112.710 147.950 113.030 148.010 ;
        RECT 112.710 147.810 117.080 147.950 ;
        RECT 112.710 147.750 113.030 147.810 ;
        RECT 75.450 147.470 76.600 147.610 ;
        RECT 75.450 147.410 75.770 147.470 ;
        RECT 19.805 147.270 20.095 147.315 ;
        RECT 20.250 147.270 20.570 147.330 ;
        RECT 19.805 147.130 20.570 147.270 ;
        RECT 19.805 147.085 20.095 147.130 ;
        RECT 20.250 147.070 20.570 147.130 ;
        RECT 32.685 147.085 32.975 147.315 ;
        RECT 22.105 146.930 22.395 146.975 ;
        RECT 27.610 146.930 27.930 146.990 ;
        RECT 22.105 146.790 27.930 146.930 ;
        RECT 22.105 146.745 22.395 146.790 ;
        RECT 27.610 146.730 27.930 146.790 ;
        RECT 30.830 146.930 31.150 146.990 ;
        RECT 32.760 146.930 32.900 147.085 ;
        RECT 34.050 147.070 34.370 147.330 ;
        RECT 41.870 147.070 42.190 147.330 ;
        RECT 55.670 147.270 55.990 147.330 ;
        RECT 61.205 147.270 61.495 147.315 ;
        RECT 63.030 147.270 63.350 147.330 ;
        RECT 55.670 147.130 63.350 147.270 ;
        RECT 55.670 147.070 55.990 147.130 ;
        RECT 61.205 147.085 61.495 147.130 ;
        RECT 63.030 147.070 63.350 147.130 ;
        RECT 63.490 147.270 63.810 147.330 ;
        RECT 65.805 147.270 66.095 147.315 ;
        RECT 63.490 147.130 66.095 147.270 ;
        RECT 63.490 147.070 63.810 147.130 ;
        RECT 65.805 147.085 66.095 147.130 ;
        RECT 70.850 147.270 71.170 147.330 ;
        RECT 71.325 147.270 71.615 147.315 ;
        RECT 70.850 147.130 71.615 147.270 ;
        RECT 70.850 147.070 71.170 147.130 ;
        RECT 71.325 147.085 71.615 147.130 ;
        RECT 73.625 147.270 73.915 147.315 ;
        RECT 75.910 147.270 76.230 147.330 ;
        RECT 76.460 147.315 76.600 147.470 ;
        RECT 77.290 147.470 78.900 147.610 ;
        RECT 77.290 147.410 77.610 147.470 ;
        RECT 78.760 147.315 78.900 147.470 ;
        RECT 79.130 147.610 79.450 147.670 ;
        RECT 97.085 147.610 97.375 147.655 ;
        RECT 97.530 147.610 97.850 147.670 ;
        RECT 79.130 147.470 80.280 147.610 ;
        RECT 79.130 147.410 79.450 147.470 ;
        RECT 73.625 147.130 76.230 147.270 ;
        RECT 73.625 147.085 73.915 147.130 ;
        RECT 75.910 147.070 76.230 147.130 ;
        RECT 76.385 147.085 76.675 147.315 ;
        RECT 78.685 147.085 78.975 147.315 ;
        RECT 79.590 147.070 79.910 147.330 ;
        RECT 80.140 147.315 80.280 147.470 ;
        RECT 97.085 147.470 97.850 147.610 ;
        RECT 97.085 147.425 97.375 147.470 ;
        RECT 97.530 147.410 97.850 147.470 ;
        RECT 106.270 147.610 106.590 147.670 ;
        RECT 108.125 147.610 108.415 147.655 ;
        RECT 113.170 147.610 113.490 147.670 ;
        RECT 116.940 147.655 117.080 147.810 ;
        RECT 120.085 147.765 120.375 147.995 ;
        RECT 106.270 147.470 108.415 147.610 ;
        RECT 106.270 147.410 106.590 147.470 ;
        RECT 108.125 147.425 108.415 147.470 ;
        RECT 111.880 147.470 113.490 147.610 ;
        RECT 80.065 147.085 80.355 147.315 ;
        RECT 80.510 147.270 80.830 147.330 ;
        RECT 81.890 147.270 82.210 147.330 ;
        RECT 80.510 147.130 82.210 147.270 ;
        RECT 80.510 147.070 80.830 147.130 ;
        RECT 81.890 147.070 82.210 147.130 ;
        RECT 83.270 147.270 83.590 147.330 ;
        RECT 83.745 147.270 84.035 147.315 ;
        RECT 83.270 147.130 84.035 147.270 ;
        RECT 83.270 147.070 83.590 147.130 ;
        RECT 83.745 147.085 84.035 147.130 ;
        RECT 84.190 147.070 84.510 147.330 ;
        RECT 84.665 147.085 84.955 147.315 ;
        RECT 40.490 146.930 40.810 146.990 ;
        RECT 43.265 146.930 43.555 146.975 ;
        RECT 30.830 146.790 43.555 146.930 ;
        RECT 30.830 146.730 31.150 146.790 ;
        RECT 40.490 146.730 40.810 146.790 ;
        RECT 43.265 146.745 43.555 146.790 ;
        RECT 59.350 146.930 59.670 146.990 ;
        RECT 84.280 146.930 84.420 147.070 ;
        RECT 59.350 146.790 84.420 146.930 ;
        RECT 84.740 146.930 84.880 147.085 ;
        RECT 85.570 147.070 85.890 147.330 ;
        RECT 93.405 147.270 93.695 147.315 ;
        RECT 94.310 147.270 94.630 147.330 ;
        RECT 93.405 147.130 94.630 147.270 ;
        RECT 93.405 147.085 93.695 147.130 ;
        RECT 94.310 147.070 94.630 147.130 ;
        RECT 96.150 147.070 96.470 147.330 ;
        RECT 99.370 147.315 99.690 147.330 ;
        RECT 99.285 147.085 99.690 147.315 ;
        RECT 99.370 147.070 99.690 147.085 ;
        RECT 99.830 147.070 100.150 147.330 ;
        RECT 100.290 147.070 100.610 147.330 ;
        RECT 101.210 147.070 101.530 147.330 ;
        RECT 109.045 147.270 109.335 147.315 ;
        RECT 109.490 147.270 109.810 147.330 ;
        RECT 111.880 147.315 112.020 147.470 ;
        RECT 113.170 147.410 113.490 147.470 ;
        RECT 116.865 147.425 117.155 147.655 ;
        RECT 109.045 147.130 109.810 147.270 ;
        RECT 109.045 147.085 109.335 147.130 ;
        RECT 109.490 147.070 109.810 147.130 ;
        RECT 111.805 147.085 112.095 147.315 ;
        RECT 112.250 147.070 112.570 147.330 ;
        RECT 112.725 147.085 113.015 147.315 ;
        RECT 86.030 146.930 86.350 146.990 ;
        RECT 84.740 146.790 86.350 146.930 ;
        RECT 59.350 146.730 59.670 146.790 ;
        RECT 21.630 146.390 21.950 146.650 ;
        RECT 23.945 146.590 24.235 146.635 ;
        RECT 25.310 146.590 25.630 146.650 ;
        RECT 23.945 146.450 25.630 146.590 ;
        RECT 23.945 146.405 24.235 146.450 ;
        RECT 25.310 146.390 25.630 146.450 ;
        RECT 34.970 146.390 35.290 146.650 ;
        RECT 56.130 146.590 56.450 146.650 ;
        RECT 60.745 146.590 61.035 146.635 ;
        RECT 56.130 146.450 61.035 146.590 ;
        RECT 56.130 146.390 56.450 146.450 ;
        RECT 60.745 146.405 61.035 146.450 ;
        RECT 61.190 146.590 61.510 146.650 ;
        RECT 64.885 146.590 65.175 146.635 ;
        RECT 61.190 146.450 65.175 146.590 ;
        RECT 61.190 146.390 61.510 146.450 ;
        RECT 64.885 146.405 65.175 146.450 ;
        RECT 71.770 146.590 72.090 146.650 ;
        RECT 74.620 146.635 74.760 146.790 ;
        RECT 86.030 146.730 86.350 146.790 ;
        RECT 97.545 146.930 97.835 146.975 ;
        RECT 98.005 146.930 98.295 146.975 ;
        RECT 97.545 146.790 98.295 146.930 ;
        RECT 99.920 146.930 100.060 147.070 ;
        RECT 106.270 146.930 106.590 146.990 ;
        RECT 99.920 146.790 106.590 146.930 ;
        RECT 97.545 146.745 97.835 146.790 ;
        RECT 98.005 146.745 98.295 146.790 ;
        RECT 106.270 146.730 106.590 146.790 ;
        RECT 107.665 146.930 107.955 146.975 ;
        RECT 110.425 146.930 110.715 146.975 ;
        RECT 107.665 146.790 110.715 146.930 ;
        RECT 107.665 146.745 107.955 146.790 ;
        RECT 110.425 146.745 110.715 146.790 ;
        RECT 72.245 146.590 72.535 146.635 ;
        RECT 71.770 146.450 72.535 146.590 ;
        RECT 71.770 146.390 72.090 146.450 ;
        RECT 72.245 146.405 72.535 146.450 ;
        RECT 74.545 146.405 74.835 146.635 ;
        RECT 78.670 146.590 78.990 146.650 ;
        RECT 80.510 146.590 80.830 146.650 ;
        RECT 78.670 146.450 80.830 146.590 ;
        RECT 78.670 146.390 78.990 146.450 ;
        RECT 80.510 146.390 80.830 146.450 ;
        RECT 81.430 146.590 81.750 146.650 ;
        RECT 81.905 146.590 82.195 146.635 ;
        RECT 81.430 146.450 82.195 146.590 ;
        RECT 81.430 146.390 81.750 146.450 ;
        RECT 81.905 146.405 82.195 146.450 ;
        RECT 82.350 146.390 82.670 146.650 ;
        RECT 92.930 146.390 93.250 146.650 ;
        RECT 95.245 146.590 95.535 146.635 ;
        RECT 103.050 146.590 103.370 146.650 ;
        RECT 95.245 146.450 103.370 146.590 ;
        RECT 95.245 146.405 95.535 146.450 ;
        RECT 103.050 146.390 103.370 146.450 ;
        RECT 109.965 146.590 110.255 146.635 ;
        RECT 111.330 146.590 111.650 146.650 ;
        RECT 109.965 146.450 111.650 146.590 ;
        RECT 112.800 146.590 112.940 147.085 ;
        RECT 113.630 147.070 113.950 147.330 ;
        RECT 118.230 147.070 118.550 147.330 ;
        RECT 120.160 147.270 120.300 147.765 ;
        RECT 121.925 147.270 122.215 147.315 ;
        RECT 120.160 147.130 122.215 147.270 ;
        RECT 121.925 147.085 122.215 147.130 ;
        RECT 117.310 146.590 117.630 146.650 ;
        RECT 117.785 146.590 118.075 146.635 ;
        RECT 112.800 146.450 118.075 146.590 ;
        RECT 109.965 146.405 110.255 146.450 ;
        RECT 111.330 146.390 111.650 146.450 ;
        RECT 117.310 146.390 117.630 146.450 ;
        RECT 117.785 146.405 118.075 146.450 ;
        RECT 122.845 146.590 123.135 146.635 ;
        RECT 124.210 146.590 124.530 146.650 ;
        RECT 122.845 146.450 124.530 146.590 ;
        RECT 122.845 146.405 123.135 146.450 ;
        RECT 124.210 146.390 124.530 146.450 ;
        RECT 14.660 145.770 127.820 146.250 ;
        RECT 18.425 145.570 18.715 145.615 ;
        RECT 21.630 145.570 21.950 145.630 ;
        RECT 18.425 145.430 21.950 145.570 ;
        RECT 18.425 145.385 18.715 145.430 ;
        RECT 21.630 145.370 21.950 145.430 ;
        RECT 27.610 145.370 27.930 145.630 ;
        RECT 43.800 145.430 48.080 145.570 ;
        RECT 19.330 145.230 19.650 145.290 ;
        RECT 19.905 145.230 20.195 145.275 ;
        RECT 23.145 145.230 23.795 145.275 ;
        RECT 19.330 145.090 23.795 145.230 ;
        RECT 19.330 145.030 19.650 145.090 ;
        RECT 19.905 145.045 20.495 145.090 ;
        RECT 23.145 145.045 23.795 145.090 ;
        RECT 29.105 145.230 29.395 145.275 ;
        RECT 32.345 145.230 32.995 145.275 ;
        RECT 29.105 145.090 32.995 145.230 ;
        RECT 29.105 145.045 29.695 145.090 ;
        RECT 32.345 145.045 32.995 145.090 ;
        RECT 17.045 144.890 17.335 144.935 ;
        RECT 17.045 144.750 20.020 144.890 ;
        RECT 17.045 144.705 17.335 144.750 ;
        RECT 19.880 144.610 20.020 144.750 ;
        RECT 20.205 144.730 20.495 145.045 ;
        RECT 21.285 144.890 21.575 144.935 ;
        RECT 24.865 144.890 25.155 144.935 ;
        RECT 26.700 144.890 26.990 144.935 ;
        RECT 21.285 144.750 26.990 144.890 ;
        RECT 21.285 144.705 21.575 144.750 ;
        RECT 24.865 144.705 25.155 144.750 ;
        RECT 26.700 144.705 26.990 144.750 ;
        RECT 29.405 144.890 29.695 145.045 ;
        RECT 34.970 145.030 35.290 145.290 ;
        RECT 36.810 145.230 37.130 145.290 ;
        RECT 39.585 145.230 39.875 145.275 ;
        RECT 36.810 145.090 43.480 145.230 ;
        RECT 36.810 145.030 37.130 145.090 ;
        RECT 39.585 145.045 39.875 145.090 ;
        RECT 29.910 144.890 30.230 144.950 ;
        RECT 29.405 144.750 30.230 144.890 ;
        RECT 29.405 144.730 29.695 144.750 ;
        RECT 29.910 144.690 30.230 144.750 ;
        RECT 30.485 144.890 30.775 144.935 ;
        RECT 34.065 144.890 34.355 144.935 ;
        RECT 35.900 144.890 36.190 144.935 ;
        RECT 30.485 144.750 36.190 144.890 ;
        RECT 30.485 144.705 30.775 144.750 ;
        RECT 34.065 144.705 34.355 144.750 ;
        RECT 35.900 144.705 36.190 144.750 ;
        RECT 39.110 144.690 39.430 144.950 ;
        RECT 42.345 144.890 42.635 144.935 ;
        RECT 42.790 144.890 43.110 144.950 ;
        RECT 43.340 144.935 43.480 145.090 ;
        RECT 43.800 144.935 43.940 145.430 ;
        RECT 46.025 145.230 46.315 145.275 ;
        RECT 46.470 145.230 46.790 145.290 ;
        RECT 46.025 145.090 46.790 145.230 ;
        RECT 46.025 145.045 46.315 145.090 ;
        RECT 46.470 145.030 46.790 145.090 ;
        RECT 47.940 145.230 48.080 145.430 ;
        RECT 63.490 145.370 63.810 145.630 ;
        RECT 65.345 145.570 65.635 145.615 ;
        RECT 68.090 145.570 68.410 145.630 ;
        RECT 65.345 145.430 68.410 145.570 ;
        RECT 65.345 145.385 65.635 145.430 ;
        RECT 68.090 145.370 68.410 145.430 ;
        RECT 86.490 145.370 86.810 145.630 ;
        RECT 53.370 145.230 53.690 145.290 ;
        RECT 47.940 145.090 53.690 145.230 ;
        RECT 47.940 144.950 48.080 145.090 ;
        RECT 53.370 145.030 53.690 145.090 ;
        RECT 55.325 145.230 55.615 145.275 ;
        RECT 56.130 145.230 56.450 145.290 ;
        RECT 58.565 145.230 59.215 145.275 ;
        RECT 55.325 145.090 59.215 145.230 ;
        RECT 55.325 145.045 55.915 145.090 ;
        RECT 42.345 144.750 43.110 144.890 ;
        RECT 42.345 144.705 42.635 144.750 ;
        RECT 42.790 144.690 43.110 144.750 ;
        RECT 43.265 144.705 43.555 144.935 ;
        RECT 43.725 144.705 44.015 144.935 ;
        RECT 44.185 144.890 44.475 144.935 ;
        RECT 45.550 144.890 45.870 144.950 ;
        RECT 47.390 144.890 47.710 144.950 ;
        RECT 44.185 144.750 47.710 144.890 ;
        RECT 44.185 144.705 44.475 144.750 ;
        RECT 45.550 144.690 45.870 144.750 ;
        RECT 47.390 144.690 47.710 144.750 ;
        RECT 47.850 144.690 48.170 144.950 ;
        RECT 48.325 144.705 48.615 144.935 ;
        RECT 49.245 144.890 49.535 144.935 ;
        RECT 49.690 144.890 50.010 144.950 ;
        RECT 49.245 144.750 50.010 144.890 ;
        RECT 49.245 144.705 49.535 144.750 ;
        RECT 19.790 144.350 20.110 144.610 ;
        RECT 25.770 144.350 26.090 144.610 ;
        RECT 27.165 144.550 27.455 144.595 ;
        RECT 28.070 144.550 28.390 144.610 ;
        RECT 36.365 144.550 36.655 144.595 ;
        RECT 27.165 144.410 36.655 144.550 ;
        RECT 27.165 144.365 27.455 144.410 ;
        RECT 28.070 144.350 28.390 144.410 ;
        RECT 36.365 144.365 36.655 144.410 ;
        RECT 36.810 144.550 37.130 144.610 ;
        RECT 38.205 144.550 38.495 144.595 ;
        RECT 48.400 144.550 48.540 144.705 ;
        RECT 49.690 144.690 50.010 144.750 ;
        RECT 55.625 144.730 55.915 145.045 ;
        RECT 56.130 145.030 56.450 145.090 ;
        RECT 58.565 145.045 59.215 145.090 ;
        RECT 61.190 145.030 61.510 145.290 ;
        RECT 79.130 145.230 79.450 145.290 ;
        RECT 86.580 145.230 86.720 145.370 ;
        RECT 79.130 145.090 82.120 145.230 ;
        RECT 79.130 145.030 79.450 145.090 ;
        RECT 56.705 144.890 56.995 144.935 ;
        RECT 60.285 144.890 60.575 144.935 ;
        RECT 62.120 144.890 62.410 144.935 ;
        RECT 56.705 144.750 62.410 144.890 ;
        RECT 56.705 144.705 56.995 144.750 ;
        RECT 60.285 144.705 60.575 144.750 ;
        RECT 62.120 144.705 62.410 144.750 ;
        RECT 63.030 144.890 63.350 144.950 ;
        RECT 67.645 144.890 67.935 144.935 ;
        RECT 68.550 144.890 68.870 144.950 ;
        RECT 63.030 144.750 68.870 144.890 ;
        RECT 63.030 144.690 63.350 144.750 ;
        RECT 67.645 144.705 67.935 144.750 ;
        RECT 68.550 144.690 68.870 144.750 ;
        RECT 69.470 144.690 69.790 144.950 ;
        RECT 81.980 144.935 82.120 145.090 ;
        RECT 85.660 145.090 86.720 145.230 ;
        RECT 91.500 145.230 91.790 145.275 ;
        RECT 92.930 145.230 93.250 145.290 ;
        RECT 94.760 145.230 95.050 145.275 ;
        RECT 91.500 145.090 95.050 145.230 ;
        RECT 81.445 144.705 81.735 144.935 ;
        RECT 81.905 144.705 82.195 144.935 ;
        RECT 82.365 144.890 82.655 144.935 ;
        RECT 82.810 144.890 83.130 144.950 ;
        RECT 82.365 144.750 83.130 144.890 ;
        RECT 82.365 144.705 82.655 144.750 ;
        RECT 36.810 144.410 38.495 144.550 ;
        RECT 17.965 144.210 18.255 144.255 ;
        RECT 20.710 144.210 21.030 144.270 ;
        RECT 17.965 144.070 21.030 144.210 ;
        RECT 17.965 144.025 18.255 144.070 ;
        RECT 20.710 144.010 21.030 144.070 ;
        RECT 21.285 144.210 21.575 144.255 ;
        RECT 24.405 144.210 24.695 144.255 ;
        RECT 26.295 144.210 26.585 144.255 ;
        RECT 21.285 144.070 26.585 144.210 ;
        RECT 21.285 144.025 21.575 144.070 ;
        RECT 24.405 144.025 24.695 144.070 ;
        RECT 26.295 144.025 26.585 144.070 ;
        RECT 30.485 144.210 30.775 144.255 ;
        RECT 33.605 144.210 33.895 144.255 ;
        RECT 35.495 144.210 35.785 144.255 ;
        RECT 30.485 144.070 35.785 144.210 ;
        RECT 36.440 144.210 36.580 144.365 ;
        RECT 36.810 144.350 37.130 144.410 ;
        RECT 38.205 144.365 38.495 144.410 ;
        RECT 40.580 144.410 48.540 144.550 ;
        RECT 62.585 144.550 62.875 144.595 ;
        RECT 65.330 144.550 65.650 144.610 ;
        RECT 62.585 144.410 65.650 144.550 ;
        RECT 37.270 144.210 37.590 144.270 ;
        RECT 36.440 144.070 37.590 144.210 ;
        RECT 30.485 144.025 30.775 144.070 ;
        RECT 33.605 144.025 33.895 144.070 ;
        RECT 35.495 144.025 35.785 144.070 ;
        RECT 37.270 144.010 37.590 144.070 ;
        RECT 22.550 143.870 22.870 143.930 ;
        RECT 40.580 143.870 40.720 144.410 ;
        RECT 62.585 144.365 62.875 144.410 ;
        RECT 65.330 144.350 65.650 144.410 ;
        RECT 65.805 144.365 66.095 144.595 ;
        RECT 56.705 144.210 56.995 144.255 ;
        RECT 59.825 144.210 60.115 144.255 ;
        RECT 61.715 144.210 62.005 144.255 ;
        RECT 65.880 144.210 66.020 144.365 ;
        RECT 66.710 144.350 67.030 144.610 ;
        RECT 81.520 144.550 81.660 144.705 ;
        RECT 82.810 144.690 83.130 144.750 ;
        RECT 83.285 144.890 83.575 144.935 ;
        RECT 83.730 144.890 84.050 144.950 ;
        RECT 83.285 144.750 84.050 144.890 ;
        RECT 83.285 144.705 83.575 144.750 ;
        RECT 83.730 144.690 84.050 144.750 ;
        RECT 85.660 144.595 85.800 145.090 ;
        RECT 91.500 145.045 91.790 145.090 ;
        RECT 92.930 145.030 93.250 145.090 ;
        RECT 94.760 145.045 95.050 145.090 ;
        RECT 95.680 145.230 95.970 145.275 ;
        RECT 97.540 145.230 97.830 145.275 ;
        RECT 95.680 145.090 97.830 145.230 ;
        RECT 95.680 145.045 95.970 145.090 ;
        RECT 97.540 145.045 97.830 145.090 ;
        RECT 104.905 145.230 105.195 145.275 ;
        RECT 107.665 145.230 107.955 145.275 ;
        RECT 110.410 145.230 110.730 145.290 ;
        RECT 104.905 145.090 107.955 145.230 ;
        RECT 104.905 145.045 105.195 145.090 ;
        RECT 107.665 145.045 107.955 145.090 ;
        RECT 108.660 145.090 110.730 145.230 ;
        RECT 86.490 144.690 86.810 144.950 ;
        RECT 93.360 144.890 93.650 144.935 ;
        RECT 95.680 144.890 95.895 145.045 ;
        RECT 93.360 144.750 95.895 144.890 ;
        RECT 99.370 144.890 99.690 144.950 ;
        RECT 106.285 144.890 106.575 144.935 ;
        RECT 108.660 144.890 108.800 145.090 ;
        RECT 110.410 145.030 110.730 145.090 ;
        RECT 115.945 145.230 116.235 145.275 ;
        RECT 119.100 145.230 119.390 145.275 ;
        RECT 122.360 145.230 122.650 145.275 ;
        RECT 115.945 145.090 122.650 145.230 ;
        RECT 115.945 145.045 116.235 145.090 ;
        RECT 119.100 145.045 119.390 145.090 ;
        RECT 122.360 145.045 122.650 145.090 ;
        RECT 123.280 145.230 123.570 145.275 ;
        RECT 125.140 145.230 125.430 145.275 ;
        RECT 123.280 145.090 125.430 145.230 ;
        RECT 123.280 145.045 123.570 145.090 ;
        RECT 125.140 145.045 125.430 145.090 ;
        RECT 99.370 144.750 106.040 144.890 ;
        RECT 93.360 144.705 93.650 144.750 ;
        RECT 99.370 144.690 99.690 144.750 ;
        RECT 81.520 144.410 82.120 144.550 ;
        RECT 81.980 144.270 82.120 144.410 ;
        RECT 85.585 144.365 85.875 144.595 ;
        RECT 86.030 144.550 86.350 144.610 ;
        RECT 89.495 144.550 89.785 144.595 ;
        RECT 91.090 144.550 91.410 144.610 ;
        RECT 86.030 144.410 91.410 144.550 ;
        RECT 86.030 144.350 86.350 144.410 ;
        RECT 89.495 144.365 89.785 144.410 ;
        RECT 91.090 144.350 91.410 144.410 ;
        RECT 96.610 144.350 96.930 144.610 ;
        RECT 98.450 144.350 98.770 144.610 ;
        RECT 104.890 144.550 105.210 144.610 ;
        RECT 105.365 144.550 105.655 144.595 ;
        RECT 104.890 144.410 105.655 144.550 ;
        RECT 105.900 144.550 106.040 144.750 ;
        RECT 106.285 144.750 108.800 144.890 ;
        RECT 106.285 144.705 106.575 144.750 ;
        RECT 109.045 144.705 109.335 144.935 ;
        RECT 109.505 144.705 109.795 144.935 ;
        RECT 109.120 144.550 109.260 144.705 ;
        RECT 105.900 144.410 109.260 144.550 ;
        RECT 104.890 144.350 105.210 144.410 ;
        RECT 105.365 144.365 105.655 144.410 ;
        RECT 74.070 144.210 74.390 144.270 ;
        RECT 56.705 144.070 62.005 144.210 ;
        RECT 56.705 144.025 56.995 144.070 ;
        RECT 59.825 144.025 60.115 144.070 ;
        RECT 61.715 144.025 62.005 144.070 ;
        RECT 65.420 144.070 66.020 144.210 ;
        RECT 66.800 144.070 74.390 144.210 ;
        RECT 22.550 143.730 40.720 143.870 ;
        RECT 22.550 143.670 22.870 143.730 ;
        RECT 41.410 143.670 41.730 143.930 ;
        RECT 45.565 143.870 45.855 143.915 ;
        RECT 50.150 143.870 50.470 143.930 ;
        RECT 45.565 143.730 50.470 143.870 ;
        RECT 45.565 143.685 45.855 143.730 ;
        RECT 50.150 143.670 50.470 143.730 ;
        RECT 53.845 143.870 54.135 143.915 ;
        RECT 58.430 143.870 58.750 143.930 ;
        RECT 65.420 143.870 65.560 144.070 ;
        RECT 53.845 143.730 65.560 143.870 ;
        RECT 65.790 143.870 66.110 143.930 ;
        RECT 66.800 143.870 66.940 144.070 ;
        RECT 74.070 144.010 74.390 144.070 ;
        RECT 81.890 144.010 82.210 144.270 ;
        RECT 93.360 144.210 93.650 144.255 ;
        RECT 96.140 144.210 96.430 144.255 ;
        RECT 98.000 144.210 98.290 144.255 ;
        RECT 93.360 144.070 98.290 144.210 ;
        RECT 93.360 144.025 93.650 144.070 ;
        RECT 96.140 144.025 96.430 144.070 ;
        RECT 98.000 144.025 98.290 144.070 ;
        RECT 106.730 144.210 107.050 144.270 ;
        RECT 109.580 144.210 109.720 144.705 ;
        RECT 109.950 144.690 110.270 144.950 ;
        RECT 110.870 144.690 111.190 144.950 ;
        RECT 111.805 144.705 112.095 144.935 ;
        RECT 113.185 144.890 113.475 144.935 ;
        RECT 113.630 144.890 113.950 144.950 ;
        RECT 113.185 144.750 113.950 144.890 ;
        RECT 113.185 144.705 113.475 144.750 ;
        RECT 111.880 144.550 112.020 144.705 ;
        RECT 113.630 144.690 113.950 144.750 ;
        RECT 115.470 144.690 115.790 144.950 ;
        RECT 117.310 144.935 117.630 144.950 ;
        RECT 117.095 144.705 117.630 144.935 ;
        RECT 120.960 144.890 121.250 144.935 ;
        RECT 123.280 144.890 123.495 145.045 ;
        RECT 120.960 144.750 123.495 144.890 ;
        RECT 120.960 144.705 121.250 144.750 ;
        RECT 117.310 144.690 117.630 144.705 ;
        RECT 124.210 144.690 124.530 144.950 ;
        RECT 119.610 144.550 119.930 144.610 ;
        RECT 111.880 144.410 119.930 144.550 ;
        RECT 119.610 144.350 119.930 144.410 ;
        RECT 126.050 144.350 126.370 144.610 ;
        RECT 112.250 144.210 112.570 144.270 ;
        RECT 106.730 144.070 112.570 144.210 ;
        RECT 106.730 144.010 107.050 144.070 ;
        RECT 112.250 144.010 112.570 144.070 ;
        RECT 120.960 144.210 121.250 144.255 ;
        RECT 123.740 144.210 124.030 144.255 ;
        RECT 125.600 144.210 125.890 144.255 ;
        RECT 120.960 144.070 125.890 144.210 ;
        RECT 120.960 144.025 121.250 144.070 ;
        RECT 123.740 144.025 124.030 144.070 ;
        RECT 125.600 144.025 125.890 144.070 ;
        RECT 65.790 143.730 66.940 143.870 ;
        RECT 53.845 143.685 54.135 143.730 ;
        RECT 58.430 143.670 58.750 143.730 ;
        RECT 65.790 143.670 66.110 143.730 ;
        RECT 68.090 143.670 68.410 143.930 ;
        RECT 70.390 143.670 70.710 143.930 ;
        RECT 78.210 143.870 78.530 143.930 ;
        RECT 80.065 143.870 80.355 143.915 ;
        RECT 78.210 143.730 80.355 143.870 ;
        RECT 78.210 143.670 78.530 143.730 ;
        RECT 80.065 143.685 80.355 143.730 ;
        RECT 88.330 143.670 88.650 143.930 ;
        RECT 105.350 143.670 105.670 143.930 ;
        RECT 106.270 143.870 106.590 143.930 ;
        RECT 107.205 143.870 107.495 143.915 ;
        RECT 106.270 143.730 107.495 143.870 ;
        RECT 106.270 143.670 106.590 143.730 ;
        RECT 107.205 143.685 107.495 143.730 ;
        RECT 14.660 143.050 127.820 143.530 ;
        RECT 19.330 142.650 19.650 142.910 ;
        RECT 19.790 142.850 20.110 142.910 ;
        RECT 20.265 142.850 20.555 142.895 ;
        RECT 19.790 142.710 20.555 142.850 ;
        RECT 19.790 142.650 20.110 142.710 ;
        RECT 20.265 142.665 20.555 142.710 ;
        RECT 25.770 142.850 26.090 142.910 ;
        RECT 26.245 142.850 26.535 142.895 ;
        RECT 25.770 142.710 26.535 142.850 ;
        RECT 25.770 142.650 26.090 142.710 ;
        RECT 26.245 142.665 26.535 142.710 ;
        RECT 29.910 142.650 30.230 142.910 ;
        RECT 31.305 142.850 31.595 142.895 ;
        RECT 32.670 142.850 32.990 142.910 ;
        RECT 31.305 142.710 32.990 142.850 ;
        RECT 31.305 142.665 31.595 142.710 ;
        RECT 32.670 142.650 32.990 142.710 ;
        RECT 37.270 142.850 37.590 142.910 ;
        RECT 45.550 142.850 45.870 142.910 ;
        RECT 37.270 142.710 41.640 142.850 ;
        RECT 37.270 142.650 37.590 142.710 ;
        RECT 35.085 142.510 35.375 142.555 ;
        RECT 38.205 142.510 38.495 142.555 ;
        RECT 40.095 142.510 40.385 142.555 ;
        RECT 23.560 142.370 32.900 142.510 ;
        RECT 22.550 141.970 22.870 142.230 ;
        RECT 23.560 142.215 23.700 142.370 ;
        RECT 23.485 141.985 23.775 142.215 ;
        RECT 32.210 141.970 32.530 142.230 ;
        RECT 32.760 142.170 32.900 142.370 ;
        RECT 35.085 142.370 40.385 142.510 ;
        RECT 35.085 142.325 35.375 142.370 ;
        RECT 38.205 142.325 38.495 142.370 ;
        RECT 40.095 142.325 40.385 142.370 ;
        RECT 36.350 142.170 36.670 142.230 ;
        RECT 32.760 142.030 36.670 142.170 ;
        RECT 36.350 141.970 36.670 142.030 ;
        RECT 37.730 142.170 38.050 142.230 ;
        RECT 39.585 142.170 39.875 142.215 ;
        RECT 37.730 142.030 39.875 142.170 ;
        RECT 37.730 141.970 38.050 142.030 ;
        RECT 39.585 141.985 39.875 142.030 ;
        RECT 40.965 142.170 41.255 142.215 ;
        RECT 41.500 142.170 41.640 142.710 ;
        RECT 40.965 142.030 41.640 142.170 ;
        RECT 45.180 142.710 45.870 142.850 ;
        RECT 40.965 141.985 41.255 142.030 ;
        RECT 19.805 141.645 20.095 141.875 ;
        RECT 19.880 141.490 20.020 141.645 ;
        RECT 25.310 141.630 25.630 141.890 ;
        RECT 29.465 141.830 29.755 141.875 ;
        RECT 30.830 141.830 31.150 141.890 ;
        RECT 29.465 141.690 31.150 141.830 ;
        RECT 29.465 141.645 29.755 141.690 ;
        RECT 20.250 141.490 20.570 141.550 ;
        RECT 29.540 141.490 29.680 141.645 ;
        RECT 30.830 141.630 31.150 141.690 ;
        RECT 32.670 141.490 32.990 141.550 ;
        RECT 34.005 141.535 34.295 141.850 ;
        RECT 35.085 141.830 35.375 141.875 ;
        RECT 38.665 141.830 38.955 141.875 ;
        RECT 40.500 141.830 40.790 141.875 ;
        RECT 35.085 141.690 40.790 141.830 ;
        RECT 35.085 141.645 35.375 141.690 ;
        RECT 38.665 141.645 38.955 141.690 ;
        RECT 40.500 141.645 40.790 141.690 ;
        RECT 41.410 141.830 41.730 141.890 ;
        RECT 42.345 141.830 42.635 141.875 ;
        RECT 41.410 141.690 42.635 141.830 ;
        RECT 41.410 141.630 41.730 141.690 ;
        RECT 42.345 141.645 42.635 141.690 ;
        RECT 42.790 141.630 43.110 141.890 ;
        RECT 43.710 141.630 44.030 141.890 ;
        RECT 44.185 141.645 44.475 141.875 ;
        RECT 44.645 141.830 44.935 141.875 ;
        RECT 45.180 141.830 45.320 142.710 ;
        RECT 45.550 142.650 45.870 142.710 ;
        RECT 51.070 142.650 51.390 142.910 ;
        RECT 69.470 142.850 69.790 142.910 ;
        RECT 68.640 142.710 69.790 142.850 ;
        RECT 46.025 142.510 46.315 142.555 ;
        RECT 45.640 142.370 46.315 142.510 ;
        RECT 45.640 142.230 45.780 142.370 ;
        RECT 46.025 142.325 46.315 142.370 ;
        RECT 64.425 142.510 64.715 142.555 ;
        RECT 68.640 142.510 68.780 142.710 ;
        RECT 69.470 142.650 69.790 142.710 ;
        RECT 78.670 142.650 78.990 142.910 ;
        RECT 81.445 142.850 81.735 142.895 ;
        RECT 83.270 142.850 83.590 142.910 ;
        RECT 81.445 142.710 83.590 142.850 ;
        RECT 81.445 142.665 81.735 142.710 ;
        RECT 83.270 142.650 83.590 142.710 ;
        RECT 93.865 142.850 94.155 142.895 ;
        RECT 96.610 142.850 96.930 142.910 ;
        RECT 112.710 142.850 113.030 142.910 ;
        RECT 93.865 142.710 96.930 142.850 ;
        RECT 93.865 142.665 94.155 142.710 ;
        RECT 96.610 142.650 96.930 142.710 ;
        RECT 107.740 142.710 113.030 142.850 ;
        RECT 64.425 142.370 68.780 142.510 ;
        RECT 68.980 142.510 69.270 142.555 ;
        RECT 71.760 142.510 72.050 142.555 ;
        RECT 73.620 142.510 73.910 142.555 ;
        RECT 68.980 142.370 73.910 142.510 ;
        RECT 64.425 142.325 64.715 142.370 ;
        RECT 68.980 142.325 69.270 142.370 ;
        RECT 71.760 142.325 72.050 142.370 ;
        RECT 73.620 142.325 73.910 142.370 ;
        RECT 45.550 141.970 45.870 142.230 ;
        RECT 46.930 142.170 47.250 142.230 ;
        RECT 49.690 142.170 50.010 142.230 ;
        RECT 46.560 142.030 50.010 142.170 ;
        RECT 46.560 141.875 46.700 142.030 ;
        RECT 46.930 141.970 47.250 142.030 ;
        RECT 49.690 141.970 50.010 142.030 ;
        RECT 50.150 142.170 50.470 142.230 ;
        RECT 51.085 142.170 51.375 142.215 ;
        RECT 50.150 142.030 51.375 142.170 ;
        RECT 50.150 141.970 50.470 142.030 ;
        RECT 51.085 141.985 51.375 142.030 ;
        RECT 61.665 142.170 61.955 142.215 ;
        RECT 65.790 142.170 66.110 142.230 ;
        RECT 66.710 142.170 67.030 142.230 ;
        RECT 61.665 142.030 67.030 142.170 ;
        RECT 61.665 141.985 61.955 142.030 ;
        RECT 65.790 141.970 66.110 142.030 ;
        RECT 66.710 141.970 67.030 142.030 ;
        RECT 70.390 142.170 70.710 142.230 ;
        RECT 72.245 142.170 72.535 142.215 ;
        RECT 70.390 142.030 72.535 142.170 ;
        RECT 70.390 141.970 70.710 142.030 ;
        RECT 72.245 141.985 72.535 142.030 ;
        RECT 74.070 141.970 74.390 142.230 ;
        RECT 78.210 141.970 78.530 142.230 ;
        RECT 80.510 141.970 80.830 142.230 ;
        RECT 88.330 142.170 88.650 142.230 ;
        RECT 105.810 142.170 106.130 142.230 ;
        RECT 107.740 142.215 107.880 142.710 ;
        RECT 112.710 142.650 113.030 142.710 ;
        RECT 109.950 142.510 110.270 142.570 ;
        RECT 115.255 142.510 115.545 142.555 ;
        RECT 116.850 142.510 117.170 142.570 ;
        RECT 109.120 142.370 117.170 142.510 ;
        RECT 107.665 142.170 107.955 142.215 ;
        RECT 88.330 142.030 93.160 142.170 ;
        RECT 88.330 141.970 88.650 142.030 ;
        RECT 44.645 141.690 45.320 141.830 ;
        RECT 44.645 141.645 44.935 141.690 ;
        RECT 46.485 141.645 46.775 141.875 ;
        RECT 33.705 141.490 34.295 141.535 ;
        RECT 36.945 141.490 37.595 141.535 ;
        RECT 19.880 141.350 29.680 141.490 ;
        RECT 31.840 141.350 32.440 141.490 ;
        RECT 20.250 141.290 20.570 141.350 ;
        RECT 21.630 141.150 21.950 141.210 ;
        RECT 22.105 141.150 22.395 141.195 ;
        RECT 31.840 141.150 31.980 141.350 ;
        RECT 21.630 141.010 31.980 141.150 ;
        RECT 32.300 141.150 32.440 141.350 ;
        RECT 32.670 141.350 37.595 141.490 ;
        RECT 44.260 141.490 44.400 141.645 ;
        RECT 47.390 141.630 47.710 141.890 ;
        RECT 47.850 141.630 48.170 141.890 ;
        RECT 48.325 141.830 48.615 141.875 ;
        RECT 48.770 141.830 49.090 141.890 ;
        RECT 48.325 141.690 49.090 141.830 ;
        RECT 48.325 141.645 48.615 141.690 ;
        RECT 48.770 141.630 49.090 141.690 ;
        RECT 52.005 141.830 52.295 141.875 ;
        RECT 52.450 141.830 52.770 141.890 ;
        RECT 52.005 141.690 52.770 141.830 ;
        RECT 52.005 141.645 52.295 141.690 ;
        RECT 52.450 141.630 52.770 141.690 ;
        RECT 57.510 141.630 57.830 141.890 ;
        RECT 57.985 141.645 58.275 141.875 ;
        RECT 44.260 141.350 44.860 141.490 ;
        RECT 32.670 141.290 32.990 141.350 ;
        RECT 33.705 141.305 33.995 141.350 ;
        RECT 36.945 141.305 37.595 141.350 ;
        RECT 37.730 141.150 38.050 141.210 ;
        RECT 32.300 141.010 38.050 141.150 ;
        RECT 21.630 140.950 21.950 141.010 ;
        RECT 22.105 140.965 22.395 141.010 ;
        RECT 37.730 140.950 38.050 141.010 ;
        RECT 38.190 141.150 38.510 141.210 ;
        RECT 41.425 141.150 41.715 141.195 ;
        RECT 38.190 141.010 41.715 141.150 ;
        RECT 44.720 141.150 44.860 141.350 ;
        RECT 47.940 141.150 48.080 141.630 ;
        RECT 50.625 141.490 50.915 141.535 ;
        RECT 56.145 141.490 56.435 141.535 ;
        RECT 50.625 141.350 56.435 141.490 ;
        RECT 50.625 141.305 50.915 141.350 ;
        RECT 56.145 141.305 56.435 141.350 ;
        RECT 44.720 141.010 48.080 141.150 ;
        RECT 38.190 140.950 38.510 141.010 ;
        RECT 41.425 140.965 41.715 141.010 ;
        RECT 49.690 140.950 50.010 141.210 ;
        RECT 52.925 141.150 53.215 141.195 ;
        RECT 54.290 141.150 54.610 141.210 ;
        RECT 52.925 141.010 54.610 141.150 ;
        RECT 58.060 141.150 58.200 141.645 ;
        RECT 58.430 141.630 58.750 141.890 ;
        RECT 59.365 141.830 59.655 141.875 ;
        RECT 60.730 141.830 61.050 141.890 ;
        RECT 59.365 141.690 61.050 141.830 ;
        RECT 59.365 141.645 59.655 141.690 ;
        RECT 60.730 141.630 61.050 141.690 ;
        RECT 68.980 141.830 69.270 141.875 ;
        RECT 76.370 141.830 76.690 141.890 ;
        RECT 77.305 141.830 77.595 141.875 ;
        RECT 68.980 141.690 71.515 141.830 ;
        RECT 68.980 141.645 69.270 141.690 ;
        RECT 58.520 141.490 58.660 141.630 ;
        RECT 62.585 141.490 62.875 141.535 ;
        RECT 58.520 141.350 62.875 141.490 ;
        RECT 62.585 141.305 62.875 141.350 ;
        RECT 67.120 141.490 67.410 141.535 ;
        RECT 68.090 141.490 68.410 141.550 ;
        RECT 71.300 141.535 71.515 141.690 ;
        RECT 76.370 141.690 77.595 141.830 ;
        RECT 76.370 141.630 76.690 141.690 ;
        RECT 77.305 141.645 77.595 141.690 ;
        RECT 80.050 141.630 80.370 141.890 ;
        RECT 81.445 141.830 81.735 141.875 ;
        RECT 82.350 141.830 82.670 141.890 ;
        RECT 81.445 141.690 82.670 141.830 ;
        RECT 81.445 141.645 81.735 141.690 ;
        RECT 82.350 141.630 82.670 141.690 ;
        RECT 82.810 141.830 83.130 141.890 ;
        RECT 83.285 141.830 83.575 141.875 ;
        RECT 82.810 141.690 83.575 141.830 ;
        RECT 82.810 141.630 83.130 141.690 ;
        RECT 83.285 141.645 83.575 141.690 ;
        RECT 83.730 141.630 84.050 141.890 ;
        RECT 84.205 141.645 84.495 141.875 ;
        RECT 85.125 141.830 85.415 141.875 ;
        RECT 86.030 141.830 86.350 141.890 ;
        RECT 85.125 141.690 86.350 141.830 ;
        RECT 85.125 141.645 85.415 141.690 ;
        RECT 70.380 141.490 70.670 141.535 ;
        RECT 67.120 141.350 70.670 141.490 ;
        RECT 67.120 141.305 67.410 141.350 ;
        RECT 68.090 141.290 68.410 141.350 ;
        RECT 70.380 141.305 70.670 141.350 ;
        RECT 71.300 141.490 71.590 141.535 ;
        RECT 73.160 141.490 73.450 141.535 ;
        RECT 71.300 141.350 73.450 141.490 ;
        RECT 71.300 141.305 71.590 141.350 ;
        RECT 73.160 141.305 73.450 141.350 ;
        RECT 78.685 141.490 78.975 141.535 ;
        RECT 81.905 141.490 82.195 141.535 ;
        RECT 78.685 141.350 82.195 141.490 ;
        RECT 84.280 141.490 84.420 141.645 ;
        RECT 86.030 141.630 86.350 141.690 ;
        RECT 91.090 141.830 91.410 141.890 ;
        RECT 93.020 141.875 93.160 142.030 ;
        RECT 105.810 142.030 107.955 142.170 ;
        RECT 105.810 141.970 106.130 142.030 ;
        RECT 107.665 141.985 107.955 142.030 ;
        RECT 109.120 141.875 109.260 142.370 ;
        RECT 109.950 142.310 110.270 142.370 ;
        RECT 115.255 142.325 115.545 142.370 ;
        RECT 116.850 142.310 117.170 142.370 ;
        RECT 119.120 142.510 119.410 142.555 ;
        RECT 121.900 142.510 122.190 142.555 ;
        RECT 123.760 142.510 124.050 142.555 ;
        RECT 119.120 142.370 124.050 142.510 ;
        RECT 119.120 142.325 119.410 142.370 ;
        RECT 121.900 142.325 122.190 142.370 ;
        RECT 123.760 142.325 124.050 142.370 ;
        RECT 112.710 142.170 113.030 142.230 ;
        RECT 112.710 142.030 122.140 142.170 ;
        RECT 112.710 141.970 113.030 142.030 ;
        RECT 91.565 141.830 91.855 141.875 ;
        RECT 91.090 141.690 91.855 141.830 ;
        RECT 91.090 141.630 91.410 141.690 ;
        RECT 91.565 141.645 91.855 141.690 ;
        RECT 92.945 141.645 93.235 141.875 ;
        RECT 109.045 141.645 109.335 141.875 ;
        RECT 113.645 141.830 113.935 141.875 ;
        RECT 115.470 141.830 115.790 141.890 ;
        RECT 113.645 141.690 115.790 141.830 ;
        RECT 113.645 141.645 113.935 141.690 ;
        RECT 115.470 141.630 115.790 141.690 ;
        RECT 119.120 141.830 119.410 141.875 ;
        RECT 122.000 141.830 122.140 142.030 ;
        RECT 122.370 141.970 122.690 142.230 ;
        RECT 124.225 141.830 124.515 141.875 ;
        RECT 126.050 141.830 126.370 141.890 ;
        RECT 119.120 141.690 121.655 141.830 ;
        RECT 122.000 141.690 126.370 141.830 ;
        RECT 119.120 141.645 119.410 141.690 ;
        RECT 86.490 141.490 86.810 141.550 ;
        RECT 89.710 141.490 90.030 141.550 ;
        RECT 121.440 141.535 121.655 141.690 ;
        RECT 124.225 141.645 124.515 141.690 ;
        RECT 126.050 141.630 126.370 141.690 ;
        RECT 84.280 141.350 90.030 141.490 ;
        RECT 78.685 141.305 78.975 141.350 ;
        RECT 81.905 141.305 82.195 141.350 ;
        RECT 86.490 141.290 86.810 141.350 ;
        RECT 89.710 141.290 90.030 141.350 ;
        RECT 114.105 141.490 114.395 141.535 ;
        RECT 117.260 141.490 117.550 141.535 ;
        RECT 120.520 141.490 120.810 141.535 ;
        RECT 114.105 141.350 120.810 141.490 ;
        RECT 114.105 141.305 114.395 141.350 ;
        RECT 117.260 141.305 117.550 141.350 ;
        RECT 120.520 141.305 120.810 141.350 ;
        RECT 121.440 141.490 121.730 141.535 ;
        RECT 123.300 141.490 123.590 141.535 ;
        RECT 121.440 141.350 123.590 141.490 ;
        RECT 121.440 141.305 121.730 141.350 ;
        RECT 123.300 141.305 123.590 141.350 ;
        RECT 135.635 141.220 136.775 165.470 ;
        RECT 59.350 141.150 59.670 141.210 ;
        RECT 58.060 141.010 59.670 141.150 ;
        RECT 52.925 140.965 53.215 141.010 ;
        RECT 54.290 140.950 54.610 141.010 ;
        RECT 59.350 140.950 59.670 141.010 ;
        RECT 62.125 141.150 62.415 141.195 ;
        RECT 63.950 141.150 64.270 141.210 ;
        RECT 65.115 141.150 65.405 141.195 ;
        RECT 62.125 141.010 65.405 141.150 ;
        RECT 62.125 140.965 62.415 141.010 ;
        RECT 63.950 140.950 64.270 141.010 ;
        RECT 65.115 140.965 65.405 141.010 ;
        RECT 75.910 141.150 76.230 141.210 ;
        RECT 76.385 141.150 76.675 141.195 ;
        RECT 75.910 141.010 76.675 141.150 ;
        RECT 75.910 140.950 76.230 141.010 ;
        RECT 76.385 140.965 76.675 141.010 ;
        RECT 79.145 141.150 79.435 141.195 ;
        RECT 79.590 141.150 79.910 141.210 ;
        RECT 79.145 141.010 79.910 141.150 ;
        RECT 79.145 140.965 79.435 141.010 ;
        RECT 79.590 140.950 79.910 141.010 ;
        RECT 92.485 141.150 92.775 141.195 ;
        RECT 96.610 141.150 96.930 141.210 ;
        RECT 92.485 141.010 96.930 141.150 ;
        RECT 92.485 140.965 92.775 141.010 ;
        RECT 96.610 140.950 96.930 141.010 ;
        RECT 104.890 141.150 105.210 141.210 ;
        RECT 108.585 141.150 108.875 141.195 ;
        RECT 104.890 141.010 108.875 141.150 ;
        RECT 104.890 140.950 105.210 141.010 ;
        RECT 108.585 140.965 108.875 141.010 ;
        RECT 109.950 141.150 110.270 141.210 ;
        RECT 110.885 141.150 111.175 141.195 ;
        RECT 109.950 141.010 111.175 141.150 ;
        RECT 109.950 140.950 110.270 141.010 ;
        RECT 110.885 140.965 111.175 141.010 ;
        RECT 14.660 140.330 127.820 140.810 ;
        RECT 135.580 140.230 136.830 141.220 ;
        RECT 33.145 140.130 33.435 140.175 ;
        RECT 34.050 140.130 34.370 140.190 ;
        RECT 33.145 139.990 34.370 140.130 ;
        RECT 33.145 139.945 33.435 139.990 ;
        RECT 34.050 139.930 34.370 139.990 ;
        RECT 42.790 140.130 43.110 140.190 ;
        RECT 43.265 140.130 43.555 140.175 ;
        RECT 42.790 139.990 43.555 140.130 ;
        RECT 42.790 139.930 43.110 139.990 ;
        RECT 43.265 139.945 43.555 139.990 ;
        RECT 47.850 140.130 48.170 140.190 ;
        RECT 53.370 140.130 53.690 140.190 ;
        RECT 89.710 140.175 90.030 140.190 ;
        RECT 47.850 139.990 53.690 140.130 ;
        RECT 47.850 139.930 48.170 139.990 ;
        RECT 53.370 139.930 53.690 139.990 ;
        RECT 89.495 139.945 90.030 140.175 ;
        RECT 89.710 139.930 90.030 139.945 ;
        RECT 116.850 139.930 117.170 140.190 ;
        RECT 117.310 139.930 117.630 140.190 ;
        RECT 119.165 140.130 119.455 140.175 ;
        RECT 121.005 140.130 121.295 140.175 ;
        RECT 122.370 140.130 122.690 140.190 ;
        RECT 135.635 140.155 136.775 140.230 ;
        RECT 119.165 139.990 120.300 140.130 ;
        RECT 119.165 139.945 119.455 139.990 ;
        RECT 27.610 139.790 27.930 139.850 ;
        RECT 35.445 139.790 35.735 139.835 ;
        RECT 43.710 139.790 44.030 139.850 ;
        RECT 27.610 139.650 44.030 139.790 ;
        RECT 27.610 139.590 27.930 139.650 ;
        RECT 35.445 139.605 35.735 139.650 ;
        RECT 43.710 139.590 44.030 139.650 ;
        RECT 45.565 139.790 45.855 139.835 ;
        RECT 57.525 139.790 57.815 139.835 ;
        RECT 45.565 139.650 57.815 139.790 ;
        RECT 45.565 139.605 45.855 139.650 ;
        RECT 57.525 139.605 57.815 139.650 ;
        RECT 57.970 139.790 58.290 139.850 ;
        RECT 71.770 139.790 72.090 139.850 ;
        RECT 81.890 139.790 82.210 139.850 ;
        RECT 82.810 139.790 83.130 139.850 ;
        RECT 57.970 139.650 83.130 139.790 ;
        RECT 57.970 139.590 58.290 139.650 ;
        RECT 32.210 139.450 32.530 139.510 ;
        RECT 34.985 139.450 35.275 139.495 ;
        RECT 39.110 139.450 39.430 139.510 ;
        RECT 32.210 139.310 43.940 139.450 ;
        RECT 32.210 139.250 32.530 139.310 ;
        RECT 34.985 139.265 35.275 139.310 ;
        RECT 39.110 139.250 39.430 139.310 ;
        RECT 36.350 138.910 36.670 139.170 ;
        RECT 43.800 139.110 43.940 139.310 ;
        RECT 44.170 139.250 44.490 139.510 ;
        RECT 44.720 139.310 47.160 139.450 ;
        RECT 44.720 139.110 44.860 139.310 ;
        RECT 43.800 138.970 44.860 139.110 ;
        RECT 45.105 139.110 45.395 139.155 ;
        RECT 46.025 139.110 46.315 139.155 ;
        RECT 45.105 138.970 46.315 139.110 ;
        RECT 47.020 139.110 47.160 139.310 ;
        RECT 47.390 139.250 47.710 139.510 ;
        RECT 47.850 139.250 48.170 139.510 ;
        RECT 48.325 139.265 48.615 139.495 ;
        RECT 49.245 139.450 49.535 139.495 ;
        RECT 50.150 139.450 50.470 139.510 ;
        RECT 58.980 139.495 59.120 139.650 ;
        RECT 71.770 139.590 72.090 139.650 ;
        RECT 81.890 139.590 82.210 139.650 ;
        RECT 82.810 139.590 83.130 139.650 ;
        RECT 91.500 139.790 91.790 139.835 ;
        RECT 93.850 139.790 94.170 139.850 ;
        RECT 94.760 139.790 95.050 139.835 ;
        RECT 91.500 139.650 95.050 139.790 ;
        RECT 91.500 139.605 91.790 139.650 ;
        RECT 93.850 139.590 94.170 139.650 ;
        RECT 94.760 139.605 95.050 139.650 ;
        RECT 95.680 139.790 95.970 139.835 ;
        RECT 97.540 139.790 97.830 139.835 ;
        RECT 95.680 139.650 97.830 139.790 ;
        RECT 95.680 139.605 95.970 139.650 ;
        RECT 97.540 139.605 97.830 139.650 ;
        RECT 105.760 139.790 106.050 139.835 ;
        RECT 107.190 139.790 107.510 139.850 ;
        RECT 109.020 139.790 109.310 139.835 ;
        RECT 105.760 139.650 109.310 139.790 ;
        RECT 105.760 139.605 106.050 139.650 ;
        RECT 49.245 139.310 50.470 139.450 ;
        RECT 49.245 139.265 49.535 139.310 ;
        RECT 48.400 139.110 48.540 139.265 ;
        RECT 50.150 139.250 50.470 139.310 ;
        RECT 58.905 139.265 59.195 139.495 ;
        RECT 59.350 139.250 59.670 139.510 ;
        RECT 59.825 139.265 60.115 139.495 ;
        RECT 47.020 138.970 48.540 139.110 ;
        RECT 58.430 139.110 58.750 139.170 ;
        RECT 59.440 139.110 59.580 139.250 ;
        RECT 58.430 138.970 59.580 139.110 ;
        RECT 59.900 139.110 60.040 139.265 ;
        RECT 60.730 139.250 61.050 139.510 ;
        RECT 68.550 139.250 68.870 139.510 ;
        RECT 69.010 139.250 69.330 139.510 ;
        RECT 69.470 139.450 69.790 139.510 ;
        RECT 71.325 139.450 71.615 139.495 ;
        RECT 69.470 139.310 71.615 139.450 ;
        RECT 69.470 139.250 69.790 139.310 ;
        RECT 71.325 139.265 71.615 139.310 ;
        RECT 93.360 139.450 93.650 139.495 ;
        RECT 95.680 139.450 95.895 139.605 ;
        RECT 107.190 139.590 107.510 139.650 ;
        RECT 109.020 139.605 109.310 139.650 ;
        RECT 109.940 139.790 110.230 139.835 ;
        RECT 111.800 139.790 112.090 139.835 ;
        RECT 109.940 139.650 112.090 139.790 ;
        RECT 109.940 139.605 110.230 139.650 ;
        RECT 111.800 139.605 112.090 139.650 ;
        RECT 93.360 139.310 95.895 139.450 ;
        RECT 93.360 139.265 93.650 139.310 ;
        RECT 96.610 139.250 96.930 139.510 ;
        RECT 98.450 139.250 98.770 139.510 ;
        RECT 107.620 139.450 107.910 139.495 ;
        RECT 109.940 139.450 110.155 139.605 ;
        RECT 120.160 139.495 120.300 139.990 ;
        RECT 121.005 139.990 122.690 140.130 ;
        RECT 121.005 139.945 121.295 139.990 ;
        RECT 122.370 139.930 122.690 139.990 ;
        RECT 107.620 139.310 110.155 139.450 ;
        RECT 107.620 139.265 107.910 139.310 ;
        RECT 120.085 139.265 120.375 139.495 ;
        RECT 129.090 139.190 134.150 139.405 ;
        RECT 143.370 139.390 144.510 223.840 ;
        RECT 137.240 139.380 144.510 139.390 ;
        RECT 136.210 139.190 144.510 139.380 ;
        RECT 63.950 139.110 64.270 139.170 ;
        RECT 59.900 138.970 64.270 139.110 ;
        RECT 45.105 138.925 45.395 138.970 ;
        RECT 46.025 138.925 46.315 138.970 ;
        RECT 58.430 138.910 58.750 138.970 ;
        RECT 63.950 138.910 64.270 138.970 ;
        RECT 110.870 138.910 111.190 139.170 ;
        RECT 112.710 138.910 113.030 139.170 ;
        RECT 113.170 139.110 113.490 139.170 ;
        RECT 115.945 139.110 116.235 139.155 ;
        RECT 113.170 138.970 116.235 139.110 ;
        RECT 113.170 138.910 113.490 138.970 ;
        RECT 115.945 138.925 116.235 138.970 ;
        RECT 93.360 138.770 93.650 138.815 ;
        RECT 96.140 138.770 96.430 138.815 ;
        RECT 98.000 138.770 98.290 138.815 ;
        RECT 93.360 138.630 98.290 138.770 ;
        RECT 93.360 138.585 93.650 138.630 ;
        RECT 96.140 138.585 96.430 138.630 ;
        RECT 98.000 138.585 98.290 138.630 ;
        RECT 107.620 138.770 107.910 138.815 ;
        RECT 110.400 138.770 110.690 138.815 ;
        RECT 112.260 138.770 112.550 138.815 ;
        RECT 107.620 138.630 112.550 138.770 ;
        RECT 107.620 138.585 107.910 138.630 ;
        RECT 110.400 138.585 110.690 138.630 ;
        RECT 112.260 138.585 112.550 138.630 ;
        RECT 129.090 138.530 144.510 139.190 ;
        RECT 44.170 138.230 44.490 138.490 ;
        RECT 72.245 138.430 72.535 138.475 ;
        RECT 73.610 138.430 73.930 138.490 ;
        RECT 72.245 138.290 73.930 138.430 ;
        RECT 72.245 138.245 72.535 138.290 ;
        RECT 73.610 138.230 73.930 138.290 ;
        RECT 99.370 138.430 99.690 138.490 ;
        RECT 100.290 138.430 100.610 138.490 ;
        RECT 103.755 138.430 104.045 138.475 ;
        RECT 104.890 138.430 105.210 138.490 ;
        RECT 99.370 138.290 105.210 138.430 ;
        RECT 99.370 138.230 99.690 138.290 ;
        RECT 100.290 138.230 100.610 138.290 ;
        RECT 103.755 138.245 104.045 138.290 ;
        RECT 104.890 138.230 105.210 138.290 ;
        RECT 129.090 138.225 134.150 138.530 ;
        RECT 136.210 138.250 144.510 138.530 ;
        RECT 136.210 138.240 138.350 138.250 ;
        RECT 14.660 137.610 127.820 138.090 ;
        RECT 49.230 137.210 49.550 137.470 ;
        RECT 82.365 137.410 82.655 137.455 ;
        RECT 82.810 137.410 83.130 137.470 ;
        RECT 82.365 137.270 83.130 137.410 ;
        RECT 82.365 137.225 82.655 137.270 ;
        RECT 82.810 137.210 83.130 137.270 ;
        RECT 91.090 137.410 91.410 137.470 ;
        RECT 92.025 137.410 92.315 137.455 ;
        RECT 91.090 137.270 92.315 137.410 ;
        RECT 91.090 137.210 91.410 137.270 ;
        RECT 92.025 137.225 92.315 137.270 ;
        RECT 92.945 137.410 93.235 137.455 ;
        RECT 93.850 137.410 94.170 137.470 ;
        RECT 105.810 137.410 106.130 137.470 ;
        RECT 92.945 137.270 94.170 137.410 ;
        RECT 92.945 137.225 93.235 137.270 ;
        RECT 93.850 137.210 94.170 137.270 ;
        RECT 98.080 137.270 106.130 137.410 ;
        RECT 65.805 137.070 66.095 137.115 ;
        RECT 69.470 137.070 69.790 137.130 ;
        RECT 65.805 136.930 69.790 137.070 ;
        RECT 65.805 136.885 66.095 136.930 ;
        RECT 69.470 136.870 69.790 136.930 ;
        RECT 70.360 137.070 70.650 137.115 ;
        RECT 73.140 137.070 73.430 137.115 ;
        RECT 75.000 137.070 75.290 137.115 ;
        RECT 70.360 136.930 75.290 137.070 ;
        RECT 70.360 136.885 70.650 136.930 ;
        RECT 73.140 136.885 73.430 136.930 ;
        RECT 75.000 136.885 75.290 136.930 ;
        RECT 63.045 136.730 63.335 136.775 ;
        RECT 72.690 136.730 73.010 136.790 ;
        RECT 63.045 136.590 66.020 136.730 ;
        RECT 63.045 136.545 63.335 136.590 ;
        RECT 65.880 136.450 66.020 136.590 ;
        RECT 72.690 136.590 73.380 136.730 ;
        RECT 72.690 136.530 73.010 136.590 ;
        RECT 29.450 136.390 29.770 136.450 ;
        RECT 47.405 136.390 47.695 136.435 ;
        RECT 29.450 136.250 47.695 136.390 ;
        RECT 29.450 136.190 29.770 136.250 ;
        RECT 47.405 136.205 47.695 136.250 ;
        RECT 48.325 136.390 48.615 136.435 ;
        RECT 51.990 136.390 52.310 136.450 ;
        RECT 48.325 136.250 52.310 136.390 ;
        RECT 48.325 136.205 48.615 136.250 ;
        RECT 51.990 136.190 52.310 136.250 ;
        RECT 63.950 136.190 64.270 136.450 ;
        RECT 65.790 136.190 66.110 136.450 ;
        RECT 70.360 136.390 70.650 136.435 ;
        RECT 73.240 136.390 73.380 136.590 ;
        RECT 73.610 136.530 73.930 136.790 ;
        RECT 74.070 136.730 74.390 136.790 ;
        RECT 75.465 136.730 75.755 136.775 ;
        RECT 74.070 136.590 75.755 136.730 ;
        RECT 74.070 136.530 74.390 136.590 ;
        RECT 75.465 136.545 75.755 136.590 ;
        RECT 80.970 136.730 81.290 136.790 ;
        RECT 81.445 136.730 81.735 136.775 ;
        RECT 80.970 136.590 81.735 136.730 ;
        RECT 80.970 136.530 81.290 136.590 ;
        RECT 81.445 136.545 81.735 136.590 ;
        RECT 86.950 136.730 87.270 136.790 ;
        RECT 88.805 136.730 89.095 136.775 ;
        RECT 86.950 136.590 89.095 136.730 ;
        RECT 86.950 136.530 87.270 136.590 ;
        RECT 88.805 136.545 89.095 136.590 ;
        RECT 82.365 136.390 82.655 136.435 ;
        RECT 70.360 136.250 72.895 136.390 ;
        RECT 73.240 136.250 82.655 136.390 ;
        RECT 88.880 136.390 89.020 136.545 ;
        RECT 89.710 136.530 90.030 136.790 ;
        RECT 98.080 136.775 98.220 137.270 ;
        RECT 105.810 137.210 106.130 137.270 ;
        RECT 107.190 137.210 107.510 137.470 ;
        RECT 110.870 137.210 111.190 137.470 ;
        RECT 101.225 136.885 101.515 137.115 ;
        RECT 98.005 136.730 98.295 136.775 ;
        RECT 90.260 136.590 98.295 136.730 ;
        RECT 90.260 136.450 90.400 136.590 ;
        RECT 98.005 136.545 98.295 136.590 ;
        RECT 90.170 136.390 90.490 136.450 ;
        RECT 88.880 136.250 90.490 136.390 ;
        RECT 70.360 136.205 70.650 136.250 ;
        RECT 68.500 136.050 68.790 136.095 ;
        RECT 69.010 136.050 69.330 136.110 ;
        RECT 72.680 136.095 72.895 136.250 ;
        RECT 82.365 136.205 82.655 136.250 ;
        RECT 90.170 136.190 90.490 136.250 ;
        RECT 93.405 136.390 93.695 136.435 ;
        RECT 94.310 136.390 94.630 136.450 ;
        RECT 93.405 136.250 94.630 136.390 ;
        RECT 93.405 136.205 93.695 136.250 ;
        RECT 94.310 136.190 94.630 136.250 ;
        RECT 99.370 136.190 99.690 136.450 ;
        RECT 101.300 136.390 101.440 136.885 ;
        RECT 103.985 136.390 104.275 136.435 ;
        RECT 101.300 136.250 104.275 136.390 ;
        RECT 103.985 136.205 104.275 136.250 ;
        RECT 106.745 136.205 107.035 136.435 ;
        RECT 71.760 136.050 72.050 136.095 ;
        RECT 68.500 135.910 72.050 136.050 ;
        RECT 68.500 135.865 68.790 135.910 ;
        RECT 69.010 135.850 69.330 135.910 ;
        RECT 71.760 135.865 72.050 135.910 ;
        RECT 72.680 136.050 72.970 136.095 ;
        RECT 74.540 136.050 74.830 136.095 ;
        RECT 72.680 135.910 74.830 136.050 ;
        RECT 72.680 135.865 72.970 135.910 ;
        RECT 74.540 135.865 74.830 135.910 ;
        RECT 80.970 135.850 81.290 136.110 ;
        RECT 94.400 136.050 94.540 136.190 ;
        RECT 106.820 136.050 106.960 136.205 ;
        RECT 109.950 136.190 110.270 136.450 ;
        RECT 113.630 136.050 113.950 136.110 ;
        RECT 94.400 135.910 113.950 136.050 ;
        RECT 113.630 135.850 113.950 135.910 ;
        RECT 63.505 135.710 63.795 135.755 ;
        RECT 66.495 135.710 66.785 135.755 ;
        RECT 67.170 135.710 67.490 135.770 ;
        RECT 63.505 135.570 67.490 135.710 ;
        RECT 63.505 135.525 63.795 135.570 ;
        RECT 66.495 135.525 66.785 135.570 ;
        RECT 67.170 135.510 67.490 135.570 ;
        RECT 83.285 135.710 83.575 135.755 ;
        RECT 84.190 135.710 84.510 135.770 ;
        RECT 83.285 135.570 84.510 135.710 ;
        RECT 83.285 135.525 83.575 135.570 ;
        RECT 84.190 135.510 84.510 135.570 ;
        RECT 89.710 135.710 90.030 135.770 ;
        RECT 90.185 135.710 90.475 135.755 ;
        RECT 89.710 135.570 90.475 135.710 ;
        RECT 89.710 135.510 90.030 135.570 ;
        RECT 90.185 135.525 90.475 135.570 ;
        RECT 97.530 135.710 97.850 135.770 ;
        RECT 98.925 135.710 99.215 135.755 ;
        RECT 97.530 135.570 99.215 135.710 ;
        RECT 97.530 135.510 97.850 135.570 ;
        RECT 98.925 135.525 99.215 135.570 ;
        RECT 104.890 135.510 105.210 135.770 ;
        RECT 14.660 134.890 127.820 135.370 ;
        RECT 42.345 134.690 42.635 134.735 ;
        RECT 44.170 134.690 44.490 134.750 ;
        RECT 42.345 134.550 44.490 134.690 ;
        RECT 42.345 134.505 42.635 134.550 ;
        RECT 44.170 134.490 44.490 134.550 ;
        RECT 44.630 134.490 44.950 134.750 ;
        RECT 45.090 134.490 45.410 134.750 ;
        RECT 46.010 134.690 46.330 134.750 ;
        RECT 48.770 134.690 49.090 134.750 ;
        RECT 46.010 134.550 49.090 134.690 ;
        RECT 46.010 134.490 46.330 134.550 ;
        RECT 48.770 134.490 49.090 134.550 ;
        RECT 80.970 134.690 81.290 134.750 ;
        RECT 82.825 134.690 83.115 134.735 ;
        RECT 80.970 134.550 83.115 134.690 ;
        RECT 80.970 134.490 81.290 134.550 ;
        RECT 82.825 134.505 83.115 134.550 ;
        RECT 109.490 134.490 109.810 134.750 ;
        RECT 111.790 134.490 112.110 134.750 ;
        RECT 112.710 134.490 113.030 134.750 ;
        RECT 26.180 134.350 26.470 134.395 ;
        RECT 26.690 134.350 27.010 134.410 ;
        RECT 29.440 134.350 29.730 134.395 ;
        RECT 26.180 134.210 29.730 134.350 ;
        RECT 26.180 134.165 26.470 134.210 ;
        RECT 26.690 134.150 27.010 134.210 ;
        RECT 29.440 134.165 29.730 134.210 ;
        RECT 30.360 134.350 30.650 134.395 ;
        RECT 32.220 134.350 32.510 134.395 ;
        RECT 30.360 134.210 32.510 134.350 ;
        RECT 30.360 134.165 30.650 134.210 ;
        RECT 32.220 134.165 32.510 134.210 ;
        RECT 47.405 134.350 47.695 134.395 ;
        RECT 57.525 134.350 57.815 134.395 ;
        RECT 47.405 134.210 57.815 134.350 ;
        RECT 47.405 134.165 47.695 134.210 ;
        RECT 57.525 134.165 57.815 134.210 ;
        RECT 58.430 134.350 58.750 134.410 ;
        RECT 97.530 134.395 97.850 134.410 ;
        RECT 91.105 134.350 91.395 134.395 ;
        RECT 97.315 134.350 97.850 134.395 ;
        RECT 58.430 134.210 59.580 134.350 ;
        RECT 28.040 134.010 28.330 134.055 ;
        RECT 30.360 134.010 30.575 134.165 ;
        RECT 58.430 134.150 58.750 134.210 ;
        RECT 59.440 134.070 59.580 134.210 ;
        RECT 80.600 134.210 84.880 134.350 ;
        RECT 28.040 133.870 30.575 134.010 ;
        RECT 28.040 133.825 28.330 133.870 ;
        RECT 34.970 133.810 35.290 134.070 ;
        RECT 40.950 134.010 41.270 134.070 ;
        RECT 41.425 134.010 41.715 134.055 ;
        RECT 40.950 133.870 41.715 134.010 ;
        RECT 40.950 133.810 41.270 133.870 ;
        RECT 41.425 133.825 41.715 133.870 ;
        RECT 43.250 133.810 43.570 134.070 ;
        RECT 43.725 134.010 44.015 134.055 ;
        RECT 46.025 134.010 46.315 134.055 ;
        RECT 43.725 133.870 46.315 134.010 ;
        RECT 43.725 133.825 44.015 133.870 ;
        RECT 23.470 133.670 23.790 133.730 ;
        RECT 24.175 133.670 24.465 133.715 ;
        RECT 29.450 133.670 29.770 133.730 ;
        RECT 23.470 133.530 29.770 133.670 ;
        RECT 23.470 133.470 23.790 133.530 ;
        RECT 24.175 133.485 24.465 133.530 ;
        RECT 29.450 133.470 29.770 133.530 ;
        RECT 31.290 133.470 31.610 133.730 ;
        RECT 33.145 133.670 33.435 133.715 ;
        RECT 34.050 133.670 34.370 133.730 ;
        RECT 33.145 133.530 34.370 133.670 ;
        RECT 33.145 133.485 33.435 133.530 ;
        RECT 34.050 133.470 34.370 133.530 ;
        RECT 40.505 133.485 40.795 133.715 ;
        RECT 28.040 133.330 28.330 133.375 ;
        RECT 30.820 133.330 31.110 133.375 ;
        RECT 32.680 133.330 32.970 133.375 ;
        RECT 40.580 133.330 40.720 133.485 ;
        RECT 28.040 133.190 32.970 133.330 ;
        RECT 28.040 133.145 28.330 133.190 ;
        RECT 30.820 133.145 31.110 133.190 ;
        RECT 32.680 133.145 32.970 133.190 ;
        RECT 33.220 133.190 40.720 133.330 ;
        RECT 45.180 133.330 45.320 133.870 ;
        RECT 46.025 133.825 46.315 133.870 ;
        RECT 46.930 133.810 47.250 134.070 ;
        RECT 48.770 133.810 49.090 134.070 ;
        RECT 57.970 134.010 58.290 134.070 ;
        RECT 58.890 134.010 59.210 134.070 ;
        RECT 57.970 133.870 59.210 134.010 ;
        RECT 57.970 133.810 58.290 133.870 ;
        RECT 58.890 133.810 59.210 133.870 ;
        RECT 59.350 133.810 59.670 134.070 ;
        RECT 59.825 133.825 60.115 134.055 ;
        RECT 60.730 134.010 61.050 134.070 ;
        RECT 80.600 134.055 80.740 134.210 ;
        RECT 84.740 134.070 84.880 134.210 ;
        RECT 85.200 134.210 97.850 134.350 ;
        RECT 79.145 134.010 79.435 134.055 ;
        RECT 60.730 133.870 79.435 134.010 ;
        RECT 45.550 133.670 45.870 133.730 ;
        RECT 47.865 133.670 48.155 133.715 ;
        RECT 45.550 133.530 48.155 133.670 ;
        RECT 45.550 133.470 45.870 133.530 ;
        RECT 47.865 133.485 48.155 133.530 ;
        RECT 55.670 133.670 55.990 133.730 ;
        RECT 59.440 133.670 59.580 133.810 ;
        RECT 55.670 133.530 59.580 133.670 ;
        RECT 59.900 133.670 60.040 133.825 ;
        RECT 60.730 133.810 61.050 133.870 ;
        RECT 79.145 133.825 79.435 133.870 ;
        RECT 80.065 133.825 80.355 134.055 ;
        RECT 80.525 133.825 80.815 134.055 ;
        RECT 80.985 134.010 81.275 134.055 ;
        RECT 81.890 134.010 82.210 134.070 ;
        RECT 84.205 134.010 84.495 134.055 ;
        RECT 80.985 133.870 84.495 134.010 ;
        RECT 80.985 133.825 81.275 133.870 ;
        RECT 67.170 133.670 67.490 133.730 ;
        RECT 59.900 133.530 67.490 133.670 ;
        RECT 55.670 133.470 55.990 133.530 ;
        RECT 67.170 133.470 67.490 133.530 ;
        RECT 51.990 133.330 52.310 133.390 ;
        RECT 45.180 133.190 52.310 133.330 ;
        RECT 79.220 133.330 79.360 133.825 ;
        RECT 80.140 133.670 80.280 133.825 ;
        RECT 81.890 133.810 82.210 133.870 ;
        RECT 84.205 133.825 84.495 133.870 ;
        RECT 84.650 133.810 84.970 134.070 ;
        RECT 85.200 134.055 85.340 134.210 ;
        RECT 91.105 134.165 91.395 134.210 ;
        RECT 97.315 134.165 97.850 134.210 ;
        RECT 99.320 134.350 99.610 134.395 ;
        RECT 100.750 134.350 101.070 134.410 ;
        RECT 102.580 134.350 102.870 134.395 ;
        RECT 99.320 134.210 102.870 134.350 ;
        RECT 99.320 134.165 99.610 134.210 ;
        RECT 97.530 134.150 97.850 134.165 ;
        RECT 100.750 134.150 101.070 134.210 ;
        RECT 102.580 134.165 102.870 134.210 ;
        RECT 103.500 134.350 103.790 134.395 ;
        RECT 105.360 134.350 105.650 134.395 ;
        RECT 112.800 134.350 112.940 134.490 ;
        RECT 135.660 134.480 136.800 134.510 ;
        RECT 103.500 134.210 105.650 134.350 ;
        RECT 103.500 134.165 103.790 134.210 ;
        RECT 105.360 134.165 105.650 134.210 ;
        RECT 106.360 134.210 112.940 134.350 ;
        RECT 85.125 133.825 85.415 134.055 ;
        RECT 86.030 133.810 86.350 134.070 ;
        RECT 89.710 134.010 90.030 134.070 ;
        RECT 90.645 134.010 90.935 134.055 ;
        RECT 93.405 134.010 93.695 134.055 ;
        RECT 89.710 133.870 90.935 134.010 ;
        RECT 89.710 133.810 90.030 133.870 ;
        RECT 90.645 133.825 90.935 133.870 ;
        RECT 93.020 133.870 93.695 134.010 ;
        RECT 89.800 133.670 89.940 133.810 ;
        RECT 80.140 133.530 89.940 133.670 ;
        RECT 90.170 133.470 90.490 133.730 ;
        RECT 86.030 133.330 86.350 133.390 ;
        RECT 93.020 133.375 93.160 133.870 ;
        RECT 93.405 133.825 93.695 133.870 ;
        RECT 101.180 134.010 101.470 134.055 ;
        RECT 103.500 134.010 103.715 134.165 ;
        RECT 101.180 133.870 103.715 134.010 ;
        RECT 104.445 134.010 104.735 134.055 ;
        RECT 104.890 134.010 105.210 134.070 ;
        RECT 104.445 133.870 105.210 134.010 ;
        RECT 101.180 133.825 101.470 133.870 ;
        RECT 104.445 133.825 104.735 133.870 ;
        RECT 104.890 133.810 105.210 133.870 ;
        RECT 106.360 133.715 106.500 134.210 ;
        RECT 107.190 134.010 107.510 134.070 ;
        RECT 110.425 134.010 110.715 134.055 ;
        RECT 107.190 133.870 110.715 134.010 ;
        RECT 107.190 133.810 107.510 133.870 ;
        RECT 110.425 133.825 110.715 133.870 ;
        RECT 111.345 134.010 111.635 134.055 ;
        RECT 112.250 134.010 112.570 134.070 ;
        RECT 111.345 133.870 112.570 134.010 ;
        RECT 111.345 133.825 111.635 133.870 ;
        RECT 106.285 133.485 106.575 133.715 ;
        RECT 110.500 133.670 110.640 133.825 ;
        RECT 112.250 133.810 112.570 133.870 ;
        RECT 112.725 133.825 113.015 134.055 ;
        RECT 112.800 133.670 112.940 133.825 ;
        RECT 113.170 133.670 113.490 133.730 ;
        RECT 110.500 133.530 113.490 133.670 ;
        RECT 113.170 133.470 113.490 133.530 ;
        RECT 113.645 133.670 113.935 133.715 ;
        RECT 116.850 133.670 117.170 133.730 ;
        RECT 113.645 133.530 117.170 133.670 ;
        RECT 113.645 133.485 113.935 133.530 ;
        RECT 116.850 133.470 117.170 133.530 ;
        RECT 135.590 133.400 136.850 134.480 ;
        RECT 79.220 133.190 86.350 133.330 ;
        RECT 28.530 132.990 28.850 133.050 ;
        RECT 33.220 132.990 33.360 133.190 ;
        RECT 51.990 133.130 52.310 133.190 ;
        RECT 86.030 133.130 86.350 133.190 ;
        RECT 92.945 133.145 93.235 133.375 ;
        RECT 101.180 133.330 101.470 133.375 ;
        RECT 103.960 133.330 104.250 133.375 ;
        RECT 105.820 133.330 106.110 133.375 ;
        RECT 101.180 133.190 106.110 133.330 ;
        RECT 101.180 133.145 101.470 133.190 ;
        RECT 103.960 133.145 104.250 133.190 ;
        RECT 105.820 133.145 106.110 133.190 ;
        RECT 28.530 132.850 33.360 132.990 ;
        RECT 28.530 132.790 28.850 132.850 ;
        RECT 35.430 132.790 35.750 133.050 ;
        RECT 46.010 132.990 46.330 133.050 ;
        RECT 47.405 132.990 47.695 133.035 ;
        RECT 46.010 132.850 47.695 132.990 ;
        RECT 46.010 132.790 46.330 132.850 ;
        RECT 47.405 132.805 47.695 132.850 ;
        RECT 49.705 132.990 49.995 133.035 ;
        RECT 50.150 132.990 50.470 133.050 ;
        RECT 49.705 132.850 50.470 132.990 ;
        RECT 49.705 132.805 49.995 132.850 ;
        RECT 50.150 132.790 50.470 132.850 ;
        RECT 82.350 132.790 82.670 133.050 ;
        RECT 94.325 132.990 94.615 133.035 ;
        RECT 95.230 132.990 95.550 133.050 ;
        RECT 94.325 132.850 95.550 132.990 ;
        RECT 94.325 132.805 94.615 132.850 ;
        RECT 95.230 132.790 95.550 132.850 ;
        RECT 14.660 132.170 127.820 132.650 ;
        RECT 21.720 131.830 26.460 131.970 ;
        RECT 21.720 131.630 21.860 131.830 ;
        RECT 21.260 131.490 21.860 131.630 ;
        RECT 21.260 131.335 21.400 131.490 ;
        RECT 23.945 131.445 24.235 131.675 ;
        RECT 26.320 131.630 26.460 131.830 ;
        RECT 26.690 131.770 27.010 132.030 ;
        RECT 29.910 131.970 30.230 132.030 ;
        RECT 27.240 131.830 41.180 131.970 ;
        RECT 27.240 131.630 27.380 131.830 ;
        RECT 29.910 131.770 30.230 131.830 ;
        RECT 34.970 131.630 35.290 131.690 ;
        RECT 26.320 131.490 27.380 131.630 ;
        RECT 28.160 131.490 35.290 131.630 ;
        RECT 21.185 131.105 21.475 131.335 ;
        RECT 21.645 131.290 21.935 131.335 ;
        RECT 23.470 131.290 23.790 131.350 ;
        RECT 21.645 131.150 23.790 131.290 ;
        RECT 21.645 131.105 21.935 131.150 ;
        RECT 23.470 131.090 23.790 131.150 ;
        RECT 19.805 130.950 20.095 130.995 ;
        RECT 24.020 130.950 24.160 131.445 ;
        RECT 25.785 130.950 26.075 130.995 ;
        RECT 19.805 130.810 20.480 130.950 ;
        RECT 24.020 130.810 26.075 130.950 ;
        RECT 19.805 130.765 20.095 130.810 ;
        RECT 20.340 130.670 20.480 130.810 ;
        RECT 25.785 130.765 26.075 130.810 ;
        RECT 26.245 130.950 26.535 130.995 ;
        RECT 28.160 130.950 28.300 131.490 ;
        RECT 34.970 131.430 35.290 131.490 ;
        RECT 35.860 131.630 36.150 131.675 ;
        RECT 38.640 131.630 38.930 131.675 ;
        RECT 40.500 131.630 40.790 131.675 ;
        RECT 35.860 131.490 40.790 131.630 ;
        RECT 35.860 131.445 36.150 131.490 ;
        RECT 38.640 131.445 38.930 131.490 ;
        RECT 40.500 131.445 40.790 131.490 ;
        RECT 28.545 131.105 28.835 131.335 ;
        RECT 29.005 131.290 29.295 131.335 ;
        RECT 31.995 131.290 32.285 131.335 ;
        RECT 34.050 131.290 34.370 131.350 ;
        RECT 29.005 131.150 33.820 131.290 ;
        RECT 29.005 131.105 29.295 131.150 ;
        RECT 31.995 131.105 32.285 131.150 ;
        RECT 26.245 130.810 28.300 130.950 ;
        RECT 26.245 130.765 26.535 130.810 ;
        RECT 20.250 130.610 20.570 130.670 ;
        RECT 26.320 130.610 26.460 130.765 ;
        RECT 20.250 130.470 26.460 130.610 ;
        RECT 28.620 130.610 28.760 131.105 ;
        RECT 29.450 130.750 29.770 131.010 ;
        RECT 29.910 130.610 30.230 130.670 ;
        RECT 28.620 130.470 30.230 130.610 ;
        RECT 20.250 130.410 20.570 130.470 ;
        RECT 29.910 130.410 30.230 130.470 ;
        RECT 19.330 130.070 19.650 130.330 ;
        RECT 22.105 130.270 22.395 130.315 ;
        RECT 22.550 130.270 22.870 130.330 ;
        RECT 22.105 130.130 22.870 130.270 ;
        RECT 22.105 130.085 22.395 130.130 ;
        RECT 22.550 130.070 22.870 130.130 ;
        RECT 23.930 130.270 24.250 130.330 ;
        RECT 24.865 130.270 25.155 130.315 ;
        RECT 23.930 130.130 25.155 130.270 ;
        RECT 23.930 130.070 24.250 130.130 ;
        RECT 24.865 130.085 25.155 130.130 ;
        RECT 31.305 130.270 31.595 130.315 ;
        RECT 33.130 130.270 33.450 130.330 ;
        RECT 31.305 130.130 33.450 130.270 ;
        RECT 33.680 130.270 33.820 131.150 ;
        RECT 34.050 131.150 38.880 131.290 ;
        RECT 34.050 131.090 34.370 131.150 ;
        RECT 35.860 130.950 36.150 130.995 ;
        RECT 38.740 130.950 38.880 131.150 ;
        RECT 39.110 131.090 39.430 131.350 ;
        RECT 41.040 131.290 41.180 131.830 ;
        RECT 47.865 131.785 48.155 132.015 ;
        RECT 43.710 131.630 44.030 131.690 ;
        RECT 47.940 131.630 48.080 131.785 ;
        RECT 50.610 131.770 50.930 132.030 ;
        RECT 55.210 131.970 55.530 132.030 ;
        RECT 58.890 131.970 59.210 132.030 ;
        RECT 55.210 131.830 59.210 131.970 ;
        RECT 55.210 131.770 55.530 131.830 ;
        RECT 58.890 131.770 59.210 131.830 ;
        RECT 81.890 131.770 82.210 132.030 ;
        RECT 88.115 131.970 88.405 132.015 ;
        RECT 89.710 131.970 90.030 132.030 ;
        RECT 88.115 131.830 90.030 131.970 ;
        RECT 88.115 131.785 88.405 131.830 ;
        RECT 89.710 131.770 90.030 131.830 ;
        RECT 100.750 131.770 101.070 132.030 ;
        RECT 103.970 131.770 104.290 132.030 ;
        RECT 105.350 131.970 105.670 132.030 ;
        RECT 106.285 131.970 106.575 132.015 ;
        RECT 105.350 131.830 106.575 131.970 ;
        RECT 105.350 131.770 105.670 131.830 ;
        RECT 106.285 131.785 106.575 131.830 ;
        RECT 109.030 131.970 109.350 132.030 ;
        RECT 112.725 131.970 113.015 132.015 ;
        RECT 109.030 131.830 113.015 131.970 ;
        RECT 109.030 131.770 109.350 131.830 ;
        RECT 112.725 131.785 113.015 131.830 ;
        RECT 91.980 131.630 92.270 131.675 ;
        RECT 94.760 131.630 95.050 131.675 ;
        RECT 96.620 131.630 96.910 131.675 ;
        RECT 43.710 131.490 48.080 131.630 ;
        RECT 55.760 131.490 70.160 131.630 ;
        RECT 43.710 131.430 44.030 131.490 ;
        RECT 45.105 131.290 45.395 131.335 ;
        RECT 48.785 131.290 49.075 131.335 ;
        RECT 49.690 131.290 50.010 131.350 ;
        RECT 51.990 131.290 52.310 131.350 ;
        RECT 55.760 131.290 55.900 131.490 ;
        RECT 61.190 131.290 61.510 131.350 ;
        RECT 41.040 131.150 48.540 131.290 ;
        RECT 45.105 131.105 45.395 131.150 ;
        RECT 40.965 130.950 41.255 130.995 ;
        RECT 35.860 130.810 38.395 130.950 ;
        RECT 38.740 130.810 41.255 130.950 ;
        RECT 35.860 130.765 36.150 130.810 ;
        RECT 34.000 130.610 34.290 130.655 ;
        RECT 35.430 130.610 35.750 130.670 ;
        RECT 38.180 130.655 38.395 130.810 ;
        RECT 40.965 130.765 41.255 130.810 ;
        RECT 46.930 130.750 47.250 131.010 ;
        RECT 47.850 130.750 48.170 131.010 ;
        RECT 48.400 130.950 48.540 131.150 ;
        RECT 48.785 131.150 50.010 131.290 ;
        RECT 48.785 131.105 49.075 131.150 ;
        RECT 49.690 131.090 50.010 131.150 ;
        RECT 51.620 131.150 55.900 131.290 ;
        RECT 56.220 131.150 61.510 131.290 ;
        RECT 50.610 130.950 50.930 131.010 ;
        RECT 51.620 130.995 51.760 131.150 ;
        RECT 51.990 131.090 52.310 131.150 ;
        RECT 48.400 130.810 50.930 130.950 ;
        RECT 50.610 130.750 50.930 130.810 ;
        RECT 51.545 130.765 51.835 130.995 ;
        RECT 52.450 130.750 52.770 131.010 ;
        RECT 55.210 130.750 55.530 131.010 ;
        RECT 55.670 130.750 55.990 131.010 ;
        RECT 56.220 130.995 56.360 131.150 ;
        RECT 61.190 131.090 61.510 131.150 ;
        RECT 65.790 131.090 66.110 131.350 ;
        RECT 56.145 130.765 56.435 130.995 ;
        RECT 57.065 130.950 57.355 130.995 ;
        RECT 57.065 130.810 58.660 130.950 ;
        RECT 57.065 130.765 57.355 130.810 ;
        RECT 37.260 130.610 37.550 130.655 ;
        RECT 34.000 130.470 37.550 130.610 ;
        RECT 34.000 130.425 34.290 130.470 ;
        RECT 35.430 130.410 35.750 130.470 ;
        RECT 37.260 130.425 37.550 130.470 ;
        RECT 38.180 130.610 38.470 130.655 ;
        RECT 40.040 130.610 40.330 130.655 ;
        RECT 43.250 130.610 43.570 130.670 ;
        RECT 44.185 130.610 44.475 130.655 ;
        RECT 47.020 130.610 47.160 130.750 ;
        RECT 38.180 130.470 40.330 130.610 ;
        RECT 38.180 130.425 38.470 130.470 ;
        RECT 40.040 130.425 40.330 130.470 ;
        RECT 40.580 130.470 44.475 130.610 ;
        RECT 40.580 130.270 40.720 130.470 ;
        RECT 43.250 130.410 43.570 130.470 ;
        RECT 44.185 130.425 44.475 130.470 ;
        RECT 45.640 130.470 47.160 130.610 ;
        RECT 49.245 130.610 49.535 130.655 ;
        RECT 57.525 130.610 57.815 130.655 ;
        RECT 49.245 130.470 57.815 130.610 ;
        RECT 45.640 130.330 45.780 130.470 ;
        RECT 49.245 130.425 49.535 130.470 ;
        RECT 57.525 130.425 57.815 130.470 ;
        RECT 33.680 130.130 40.720 130.270 ;
        RECT 31.305 130.085 31.595 130.130 ;
        RECT 33.130 130.070 33.450 130.130 ;
        RECT 42.330 130.070 42.650 130.330 ;
        RECT 44.645 130.270 44.935 130.315 ;
        RECT 45.550 130.270 45.870 130.330 ;
        RECT 44.645 130.130 45.870 130.270 ;
        RECT 44.645 130.085 44.935 130.130 ;
        RECT 45.550 130.070 45.870 130.130 ;
        RECT 46.945 130.270 47.235 130.315 ;
        RECT 51.990 130.270 52.310 130.330 ;
        RECT 46.945 130.130 52.310 130.270 ;
        RECT 46.945 130.085 47.235 130.130 ;
        RECT 51.990 130.070 52.310 130.130 ;
        RECT 53.830 130.070 54.150 130.330 ;
        RECT 58.520 130.270 58.660 130.810 ;
        RECT 58.890 130.750 59.210 131.010 ;
        RECT 59.350 130.750 59.670 131.010 ;
        RECT 59.825 130.765 60.115 130.995 ;
        RECT 59.900 130.610 60.040 130.765 ;
        RECT 60.730 130.750 61.050 131.010 ;
        RECT 67.170 130.750 67.490 131.010 ;
        RECT 69.485 130.950 69.775 130.995 ;
        RECT 69.100 130.810 69.775 130.950 ;
        RECT 59.900 130.470 65.560 130.610 ;
        RECT 65.420 130.330 65.560 130.470 ;
        RECT 60.730 130.270 61.050 130.330 ;
        RECT 58.520 130.130 61.050 130.270 ;
        RECT 60.730 130.070 61.050 130.130 ;
        RECT 65.330 130.270 65.650 130.330 ;
        RECT 69.100 130.315 69.240 130.810 ;
        RECT 69.485 130.765 69.775 130.810 ;
        RECT 70.020 130.610 70.160 131.490 ;
        RECT 91.980 131.490 96.910 131.630 ;
        RECT 91.980 131.445 92.270 131.490 ;
        RECT 94.760 131.445 95.050 131.490 ;
        RECT 96.620 131.445 96.910 131.490 ;
        RECT 112.250 131.630 112.570 131.690 ;
        RECT 115.930 131.630 116.250 131.690 ;
        RECT 112.250 131.490 117.080 131.630 ;
        RECT 112.250 131.430 112.570 131.490 ;
        RECT 115.930 131.430 116.250 131.490 ;
        RECT 81.430 131.090 81.750 131.350 ;
        RECT 95.230 131.090 95.550 131.350 ;
        RECT 97.085 131.290 97.375 131.335 ;
        RECT 98.450 131.290 98.770 131.350 ;
        RECT 109.505 131.290 109.795 131.335 ;
        RECT 109.950 131.290 110.270 131.350 ;
        RECT 116.940 131.335 117.080 131.490 ;
        RECT 116.405 131.290 116.695 131.335 ;
        RECT 97.085 131.150 98.770 131.290 ;
        RECT 97.085 131.105 97.375 131.150 ;
        RECT 98.450 131.090 98.770 131.150 ;
        RECT 104.980 131.150 106.500 131.290 ;
        RECT 70.850 130.750 71.170 131.010 ;
        RECT 71.310 130.950 71.630 131.010 ;
        RECT 71.785 130.950 72.075 130.995 ;
        RECT 73.625 130.950 73.915 130.995 ;
        RECT 75.450 130.950 75.770 131.010 ;
        RECT 71.310 130.810 75.770 130.950 ;
        RECT 71.310 130.750 71.630 130.810 ;
        RECT 71.785 130.765 72.075 130.810 ;
        RECT 73.625 130.765 73.915 130.810 ;
        RECT 75.450 130.750 75.770 130.810 ;
        RECT 80.970 130.750 81.290 131.010 ;
        RECT 82.350 130.750 82.670 131.010 ;
        RECT 91.980 130.950 92.270 130.995 ;
        RECT 94.770 130.950 95.090 131.010 ;
        RECT 98.910 130.950 99.230 131.010 ;
        RECT 104.980 130.995 105.120 131.150 ;
        RECT 100.305 130.950 100.595 130.995 ;
        RECT 91.980 130.810 94.515 130.950 ;
        RECT 91.980 130.765 92.270 130.810 ;
        RECT 93.390 130.655 93.710 130.670 ;
        RECT 72.705 130.610 72.995 130.655 ;
        RECT 90.120 130.610 90.410 130.655 ;
        RECT 93.380 130.610 93.710 130.655 ;
        RECT 70.020 130.470 85.110 130.610 ;
        RECT 72.705 130.425 72.995 130.470 ;
        RECT 66.725 130.270 67.015 130.315 ;
        RECT 65.330 130.130 67.015 130.270 ;
        RECT 65.330 130.070 65.650 130.130 ;
        RECT 66.725 130.085 67.015 130.130 ;
        RECT 69.025 130.085 69.315 130.315 ;
        RECT 70.405 130.270 70.695 130.315 ;
        RECT 72.230 130.270 72.550 130.330 ;
        RECT 70.405 130.130 72.550 130.270 ;
        RECT 70.405 130.085 70.695 130.130 ;
        RECT 72.230 130.070 72.550 130.130 ;
        RECT 80.065 130.270 80.355 130.315 ;
        RECT 81.430 130.270 81.750 130.330 ;
        RECT 80.065 130.130 81.750 130.270 ;
        RECT 84.970 130.270 85.110 130.470 ;
        RECT 90.120 130.470 93.710 130.610 ;
        RECT 90.120 130.425 90.410 130.470 ;
        RECT 93.380 130.425 93.710 130.470 ;
        RECT 94.300 130.655 94.515 130.810 ;
        RECT 94.770 130.810 100.595 130.950 ;
        RECT 94.770 130.750 95.090 130.810 ;
        RECT 98.910 130.750 99.230 130.810 ;
        RECT 100.305 130.765 100.595 130.810 ;
        RECT 104.905 130.765 105.195 130.995 ;
        RECT 105.825 130.765 106.115 130.995 ;
        RECT 106.360 130.950 106.500 131.150 ;
        RECT 109.505 131.150 116.695 131.290 ;
        RECT 109.505 131.105 109.795 131.150 ;
        RECT 109.950 131.090 110.270 131.150 ;
        RECT 116.405 131.105 116.695 131.150 ;
        RECT 116.865 131.105 117.155 131.335 ;
        RECT 107.190 130.950 107.510 131.010 ;
        RECT 106.360 130.810 107.510 130.950 ;
        RECT 94.300 130.610 94.590 130.655 ;
        RECT 96.160 130.610 96.450 130.655 ;
        RECT 104.980 130.610 105.120 130.765 ;
        RECT 94.300 130.470 96.450 130.610 ;
        RECT 94.300 130.425 94.590 130.470 ;
        RECT 96.160 130.425 96.450 130.470 ;
        RECT 100.380 130.470 105.120 130.610 ;
        RECT 105.900 130.610 106.040 130.765 ;
        RECT 107.190 130.750 107.510 130.810 ;
        RECT 108.125 130.950 108.415 130.995 ;
        RECT 109.030 130.950 109.350 131.010 ;
        RECT 110.425 130.950 110.715 130.995 ;
        RECT 108.125 130.810 110.715 130.950 ;
        RECT 108.125 130.765 108.415 130.810 ;
        RECT 109.030 130.750 109.350 130.810 ;
        RECT 110.425 130.765 110.715 130.810 ;
        RECT 113.170 130.950 113.490 131.010 ;
        RECT 113.645 130.950 113.935 130.995 ;
        RECT 113.170 130.810 113.935 130.950 ;
        RECT 113.170 130.750 113.490 130.810 ;
        RECT 113.645 130.765 113.935 130.810 ;
        RECT 114.565 130.950 114.855 130.995 ;
        RECT 117.310 130.950 117.630 131.010 ;
        RECT 114.565 130.810 117.630 130.950 ;
        RECT 114.565 130.765 114.855 130.810 ;
        RECT 109.490 130.610 109.810 130.670 ;
        RECT 105.900 130.470 109.810 130.610 ;
        RECT 93.390 130.410 93.710 130.425 ;
        RECT 100.380 130.330 100.520 130.470 ;
        RECT 109.490 130.410 109.810 130.470 ;
        RECT 109.965 130.610 110.255 130.655 ;
        RECT 114.640 130.610 114.780 130.765 ;
        RECT 117.310 130.750 117.630 130.810 ;
        RECT 109.965 130.470 114.780 130.610 ;
        RECT 109.965 130.425 110.255 130.470 ;
        RECT 100.290 130.270 100.610 130.330 ;
        RECT 84.970 130.130 100.610 130.270 ;
        RECT 80.065 130.085 80.355 130.130 ;
        RECT 81.430 130.070 81.750 130.130 ;
        RECT 100.290 130.070 100.610 130.130 ;
        RECT 111.790 130.270 112.110 130.330 ;
        RECT 112.265 130.270 112.555 130.315 ;
        RECT 111.790 130.130 112.555 130.270 ;
        RECT 111.790 130.070 112.110 130.130 ;
        RECT 112.265 130.085 112.555 130.130 ;
        RECT 116.850 130.270 117.170 130.330 ;
        RECT 117.325 130.270 117.615 130.315 ;
        RECT 116.850 130.130 117.615 130.270 ;
        RECT 116.850 130.070 117.170 130.130 ;
        RECT 117.325 130.085 117.615 130.130 ;
        RECT 119.150 130.070 119.470 130.330 ;
        RECT 14.660 129.450 127.820 129.930 ;
        RECT 16.815 129.250 17.105 129.295 ;
        RECT 22.550 129.250 22.870 129.310 ;
        RECT 31.290 129.250 31.610 129.310 ;
        RECT 32.225 129.250 32.515 129.295 ;
        RECT 16.815 129.110 31.060 129.250 ;
        RECT 16.815 129.065 17.105 129.110 ;
        RECT 22.550 129.050 22.870 129.110 ;
        RECT 18.820 128.910 19.110 128.955 ;
        RECT 19.330 128.910 19.650 128.970 ;
        RECT 22.080 128.910 22.370 128.955 ;
        RECT 18.820 128.770 22.370 128.910 ;
        RECT 18.820 128.725 19.110 128.770 ;
        RECT 19.330 128.710 19.650 128.770 ;
        RECT 22.080 128.725 22.370 128.770 ;
        RECT 23.000 128.910 23.290 128.955 ;
        RECT 24.860 128.910 25.150 128.955 ;
        RECT 23.000 128.770 25.150 128.910 ;
        RECT 30.920 128.910 31.060 129.110 ;
        RECT 31.290 129.110 32.515 129.250 ;
        RECT 31.290 129.050 31.610 129.110 ;
        RECT 32.225 129.065 32.515 129.110 ;
        RECT 39.110 129.250 39.430 129.310 ;
        RECT 41.425 129.250 41.715 129.295 ;
        RECT 39.110 129.110 41.715 129.250 ;
        RECT 39.110 129.050 39.430 129.110 ;
        RECT 41.425 129.065 41.715 129.110 ;
        RECT 44.630 129.050 44.950 129.310 ;
        RECT 49.230 129.250 49.550 129.310 ;
        RECT 49.705 129.250 49.995 129.295 ;
        RECT 73.610 129.250 73.930 129.310 ;
        RECT 74.545 129.250 74.835 129.295 ;
        RECT 49.230 129.110 49.995 129.250 ;
        RECT 49.230 129.050 49.550 129.110 ;
        RECT 49.705 129.065 49.995 129.110 ;
        RECT 55.760 129.110 74.835 129.250 ;
        RECT 47.405 128.910 47.695 128.955 ;
        RECT 53.830 128.910 54.150 128.970 ;
        RECT 55.760 128.955 55.900 129.110 ;
        RECT 73.610 129.050 73.930 129.110 ;
        RECT 74.545 129.065 74.835 129.110 ;
        RECT 82.365 129.250 82.655 129.295 ;
        RECT 82.810 129.250 83.130 129.310 ;
        RECT 82.365 129.110 83.130 129.250 ;
        RECT 82.365 129.065 82.655 129.110 ;
        RECT 82.810 129.050 83.130 129.110 ;
        RECT 92.945 129.250 93.235 129.295 ;
        RECT 93.390 129.250 93.710 129.310 ;
        RECT 92.945 129.110 93.710 129.250 ;
        RECT 92.945 129.065 93.235 129.110 ;
        RECT 93.390 129.050 93.710 129.110 ;
        RECT 97.990 129.250 98.310 129.310 ;
        RECT 116.850 129.295 117.170 129.310 ;
        RECT 99.385 129.250 99.675 129.295 ;
        RECT 97.990 129.110 99.675 129.250 ;
        RECT 97.990 129.050 98.310 129.110 ;
        RECT 99.385 129.065 99.675 129.110 ;
        RECT 116.635 129.065 117.170 129.295 ;
        RECT 116.850 129.050 117.170 129.065 ;
        RECT 30.920 128.770 43.020 128.910 ;
        RECT 23.000 128.725 23.290 128.770 ;
        RECT 24.860 128.725 25.150 128.770 ;
        RECT 20.680 128.570 20.970 128.615 ;
        RECT 23.000 128.570 23.215 128.725 ;
        RECT 20.680 128.430 23.215 128.570 ;
        RECT 20.680 128.385 20.970 128.430 ;
        RECT 23.930 128.370 24.250 128.630 ;
        RECT 33.130 128.370 33.450 128.630 ;
        RECT 42.330 128.370 42.650 128.630 ;
        RECT 42.880 128.615 43.020 128.770 ;
        RECT 47.405 128.770 54.150 128.910 ;
        RECT 47.405 128.725 47.695 128.770 ;
        RECT 53.830 128.710 54.150 128.770 ;
        RECT 55.685 128.725 55.975 128.955 ;
        RECT 59.810 128.910 60.130 128.970 ;
        RECT 58.980 128.770 60.130 128.910 ;
        RECT 42.805 128.385 43.095 128.615 ;
        RECT 43.250 128.570 43.570 128.630 ;
        RECT 43.725 128.570 44.015 128.615 ;
        RECT 43.250 128.430 44.015 128.570 ;
        RECT 43.250 128.370 43.570 128.430 ;
        RECT 43.725 128.385 44.015 128.430 ;
        RECT 46.025 128.385 46.315 128.615 ;
        RECT 25.785 128.230 26.075 128.275 ;
        RECT 30.370 128.230 30.690 128.290 ;
        RECT 34.050 128.230 34.370 128.290 ;
        RECT 25.785 128.090 34.370 128.230 ;
        RECT 25.785 128.045 26.075 128.090 ;
        RECT 30.370 128.030 30.690 128.090 ;
        RECT 34.050 128.030 34.370 128.090 ;
        RECT 41.870 128.230 42.190 128.290 ;
        RECT 46.100 128.230 46.240 128.385 ;
        RECT 46.470 128.370 46.790 128.630 ;
        RECT 50.625 128.570 50.915 128.615 ;
        RECT 51.070 128.570 51.390 128.630 ;
        RECT 50.625 128.430 51.390 128.570 ;
        RECT 50.625 128.385 50.915 128.430 ;
        RECT 51.070 128.370 51.390 128.430 ;
        RECT 52.005 128.385 52.295 128.615 ;
        RECT 41.870 128.090 46.240 128.230 ;
        RECT 41.870 128.030 42.190 128.090 ;
        RECT 51.545 128.045 51.835 128.275 ;
        RECT 52.080 128.230 52.220 128.385 ;
        RECT 58.430 128.370 58.750 128.630 ;
        RECT 58.980 128.615 59.120 128.770 ;
        RECT 59.810 128.710 60.130 128.770 ;
        RECT 62.125 128.910 62.415 128.955 ;
        RECT 67.120 128.910 67.410 128.955 ;
        RECT 70.380 128.910 70.670 128.955 ;
        RECT 62.125 128.770 70.670 128.910 ;
        RECT 62.125 128.725 62.415 128.770 ;
        RECT 67.120 128.725 67.410 128.770 ;
        RECT 70.380 128.725 70.670 128.770 ;
        RECT 71.300 128.910 71.590 128.955 ;
        RECT 73.160 128.910 73.450 128.955 ;
        RECT 71.300 128.770 73.450 128.910 ;
        RECT 71.300 128.725 71.590 128.770 ;
        RECT 73.160 128.725 73.450 128.770 ;
        RECT 112.265 128.910 112.555 128.955 ;
        RECT 112.710 128.910 113.030 128.970 ;
        RECT 112.265 128.770 113.030 128.910 ;
        RECT 112.265 128.725 112.555 128.770 ;
        RECT 58.905 128.385 59.195 128.615 ;
        RECT 59.365 128.385 59.655 128.615 ;
        RECT 60.285 128.570 60.575 128.615 ;
        RECT 60.730 128.570 61.050 128.630 ;
        RECT 65.330 128.615 65.650 128.630 ;
        RECT 60.285 128.430 61.050 128.570 ;
        RECT 60.285 128.385 60.575 128.430 ;
        RECT 57.065 128.230 57.355 128.275 ;
        RECT 52.080 128.090 57.355 128.230 ;
        RECT 57.065 128.045 57.355 128.090 ;
        RECT 20.680 127.890 20.970 127.935 ;
        RECT 23.460 127.890 23.750 127.935 ;
        RECT 25.320 127.890 25.610 127.935 ;
        RECT 20.680 127.750 25.610 127.890 ;
        RECT 20.680 127.705 20.970 127.750 ;
        RECT 23.460 127.705 23.750 127.750 ;
        RECT 25.320 127.705 25.610 127.750 ;
        RECT 45.090 127.690 45.410 127.950 ;
        RECT 51.620 127.890 51.760 128.045 ;
        RECT 52.910 127.890 53.230 127.950 ;
        RECT 51.620 127.750 53.230 127.890 ;
        RECT 59.440 127.890 59.580 128.385 ;
        RECT 60.730 128.370 61.050 128.430 ;
        RECT 61.665 128.570 61.955 128.615 ;
        RECT 63.505 128.570 63.795 128.615 ;
        RECT 61.665 128.430 63.795 128.570 ;
        RECT 61.665 128.385 61.955 128.430 ;
        RECT 63.505 128.385 63.795 128.430 ;
        RECT 65.115 128.385 65.650 128.615 ;
        RECT 68.980 128.570 69.270 128.615 ;
        RECT 71.300 128.570 71.515 128.725 ;
        RECT 112.710 128.710 113.030 128.770 ;
        RECT 113.645 128.910 113.935 128.955 ;
        RECT 118.640 128.910 118.930 128.955 ;
        RECT 121.900 128.910 122.190 128.955 ;
        RECT 113.645 128.770 122.190 128.910 ;
        RECT 113.645 128.725 113.935 128.770 ;
        RECT 118.640 128.725 118.930 128.770 ;
        RECT 121.900 128.725 122.190 128.770 ;
        RECT 122.820 128.910 123.110 128.955 ;
        RECT 124.680 128.910 124.970 128.955 ;
        RECT 122.820 128.770 124.970 128.910 ;
        RECT 122.820 128.725 123.110 128.770 ;
        RECT 124.680 128.725 124.970 128.770 ;
        RECT 68.980 128.430 71.515 128.570 ;
        RECT 68.980 128.385 69.270 128.430 ;
        RECT 63.580 128.230 63.720 128.385 ;
        RECT 65.330 128.370 65.650 128.385 ;
        RECT 72.230 128.370 72.550 128.630 ;
        RECT 74.070 128.370 74.390 128.630 ;
        RECT 75.450 128.370 75.770 128.630 ;
        RECT 82.350 128.570 82.670 128.630 ;
        RECT 83.285 128.570 83.575 128.615 ;
        RECT 82.350 128.430 83.575 128.570 ;
        RECT 82.350 128.370 82.670 128.430 ;
        RECT 83.285 128.385 83.575 128.430 ;
        RECT 83.730 128.370 84.050 128.630 ;
        RECT 93.405 128.570 93.695 128.615 ;
        RECT 94.310 128.570 94.630 128.630 ;
        RECT 93.405 128.430 94.630 128.570 ;
        RECT 93.405 128.385 93.695 128.430 ;
        RECT 94.310 128.370 94.630 128.430 ;
        RECT 100.290 128.370 100.610 128.630 ;
        RECT 103.510 128.370 103.830 128.630 ;
        RECT 68.550 128.230 68.870 128.290 ;
        RECT 63.580 128.090 68.870 128.230 ;
        RECT 68.550 128.030 68.870 128.090 ;
        RECT 74.990 128.230 75.310 128.290 ;
        RECT 76.370 128.230 76.690 128.290 ;
        RECT 74.990 128.090 76.690 128.230 ;
        RECT 74.990 128.030 75.310 128.090 ;
        RECT 76.370 128.030 76.690 128.090 ;
        RECT 101.210 128.030 101.530 128.290 ;
        RECT 112.800 128.230 112.940 128.710 ;
        RECT 113.170 128.570 113.490 128.630 ;
        RECT 115.025 128.570 115.315 128.615 ;
        RECT 113.170 128.430 115.315 128.570 ;
        RECT 113.170 128.370 113.490 128.430 ;
        RECT 115.025 128.385 115.315 128.430 ;
        RECT 120.500 128.570 120.790 128.615 ;
        RECT 122.820 128.570 123.035 128.725 ;
        RECT 120.500 128.430 123.035 128.570 ;
        RECT 123.765 128.570 124.055 128.615 ;
        RECT 125.130 128.570 125.450 128.630 ;
        RECT 123.765 128.430 125.450 128.570 ;
        RECT 120.500 128.385 120.790 128.430 ;
        RECT 123.765 128.385 124.055 128.430 ;
        RECT 125.130 128.370 125.450 128.430 ;
        RECT 124.210 128.230 124.530 128.290 ;
        RECT 125.605 128.230 125.895 128.275 ;
        RECT 112.800 128.090 125.895 128.230 ;
        RECT 124.210 128.030 124.530 128.090 ;
        RECT 125.605 128.045 125.895 128.090 ;
        RECT 64.870 127.890 65.190 127.950 ;
        RECT 59.440 127.750 65.190 127.890 ;
        RECT 52.910 127.690 53.230 127.750 ;
        RECT 64.870 127.690 65.190 127.750 ;
        RECT 68.980 127.890 69.270 127.935 ;
        RECT 71.760 127.890 72.050 127.935 ;
        RECT 73.620 127.890 73.910 127.935 ;
        RECT 68.980 127.750 73.910 127.890 ;
        RECT 68.980 127.705 69.270 127.750 ;
        RECT 71.760 127.705 72.050 127.750 ;
        RECT 73.620 127.705 73.910 127.750 ;
        RECT 120.500 127.890 120.790 127.935 ;
        RECT 123.280 127.890 123.570 127.935 ;
        RECT 125.140 127.890 125.430 127.935 ;
        RECT 120.500 127.750 125.430 127.890 ;
        RECT 120.500 127.705 120.790 127.750 ;
        RECT 123.280 127.705 123.570 127.750 ;
        RECT 125.140 127.705 125.430 127.750 ;
        RECT 41.410 127.550 41.730 127.610 ;
        RECT 46.025 127.550 46.315 127.595 ;
        RECT 41.410 127.410 46.315 127.550 ;
        RECT 41.410 127.350 41.730 127.410 ;
        RECT 46.025 127.365 46.315 127.410 ;
        RECT 49.690 127.550 50.010 127.610 ;
        RECT 50.625 127.550 50.915 127.595 ;
        RECT 49.690 127.410 50.915 127.550 ;
        RECT 49.690 127.350 50.010 127.410 ;
        RECT 50.625 127.365 50.915 127.410 ;
        RECT 51.070 127.550 51.390 127.610 ;
        RECT 54.305 127.550 54.595 127.595 ;
        RECT 51.070 127.410 54.595 127.550 ;
        RECT 51.070 127.350 51.390 127.410 ;
        RECT 54.305 127.365 54.595 127.410 ;
        RECT 63.965 127.550 64.255 127.595 ;
        RECT 64.410 127.550 64.730 127.610 ;
        RECT 63.965 127.410 64.730 127.550 ;
        RECT 63.965 127.365 64.255 127.410 ;
        RECT 64.410 127.350 64.730 127.410 ;
        RECT 115.470 127.350 115.790 127.610 ;
        RECT 14.660 126.730 127.820 127.210 ;
        RECT 34.140 126.390 42.560 126.530 ;
        RECT 22.550 125.650 22.870 125.910 ;
        RECT 23.485 125.850 23.775 125.895 ;
        RECT 24.390 125.850 24.710 125.910 ;
        RECT 29.005 125.850 29.295 125.895 ;
        RECT 29.910 125.850 30.230 125.910 ;
        RECT 31.290 125.850 31.610 125.910 ;
        RECT 33.605 125.850 33.895 125.895 ;
        RECT 23.485 125.710 33.895 125.850 ;
        RECT 23.485 125.665 23.775 125.710 ;
        RECT 24.390 125.650 24.710 125.710 ;
        RECT 29.005 125.665 29.295 125.710 ;
        RECT 29.910 125.650 30.230 125.710 ;
        RECT 31.290 125.650 31.610 125.710 ;
        RECT 33.605 125.665 33.895 125.710 ;
        RECT 18.885 125.510 19.175 125.555 ;
        RECT 22.105 125.510 22.395 125.555 ;
        RECT 28.085 125.510 28.375 125.555 ;
        RECT 28.530 125.510 28.850 125.570 ;
        RECT 18.885 125.370 20.480 125.510 ;
        RECT 18.885 125.325 19.175 125.370 ;
        RECT 19.330 124.830 19.650 124.890 ;
        RECT 20.340 124.875 20.480 125.370 ;
        RECT 22.105 125.370 23.010 125.510 ;
        RECT 22.105 125.325 22.395 125.370 ;
        RECT 22.870 125.170 23.010 125.370 ;
        RECT 28.085 125.370 28.850 125.510 ;
        RECT 28.085 125.325 28.375 125.370 ;
        RECT 23.470 125.170 23.790 125.230 ;
        RECT 28.160 125.170 28.300 125.325 ;
        RECT 28.530 125.310 28.850 125.370 ;
        RECT 22.870 125.030 28.300 125.170 ;
        RECT 23.470 124.970 23.790 125.030 ;
        RECT 19.805 124.830 20.095 124.875 ;
        RECT 19.330 124.690 20.095 124.830 ;
        RECT 19.330 124.630 19.650 124.690 ;
        RECT 19.805 124.645 20.095 124.690 ;
        RECT 20.265 124.645 20.555 124.875 ;
        RECT 23.010 124.830 23.330 124.890 ;
        RECT 25.785 124.830 26.075 124.875 ;
        RECT 23.010 124.690 26.075 124.830 ;
        RECT 23.010 124.630 23.330 124.690 ;
        RECT 25.785 124.645 26.075 124.690 ;
        RECT 27.625 124.830 27.915 124.875 ;
        RECT 29.910 124.830 30.230 124.890 ;
        RECT 34.140 124.830 34.280 126.390 ;
        RECT 36.350 126.190 36.670 126.250 ;
        RECT 42.420 126.190 42.560 126.390 ;
        RECT 43.710 126.330 44.030 126.590 ;
        RECT 49.690 126.330 50.010 126.590 ;
        RECT 81.890 126.530 82.210 126.590 ;
        RECT 82.365 126.530 82.655 126.575 ;
        RECT 81.890 126.390 82.655 126.530 ;
        RECT 81.890 126.330 82.210 126.390 ;
        RECT 82.365 126.345 82.655 126.390 ;
        RECT 125.130 126.330 125.450 126.590 ;
        RECT 65.300 126.190 65.590 126.235 ;
        RECT 68.080 126.190 68.370 126.235 ;
        RECT 69.940 126.190 70.230 126.235 ;
        RECT 36.350 126.050 42.100 126.190 ;
        RECT 42.420 126.050 44.400 126.190 ;
        RECT 36.350 125.990 36.670 126.050 ;
        RECT 35.430 125.850 35.750 125.910 ;
        RECT 39.585 125.850 39.875 125.895 ;
        RECT 34.600 125.710 39.875 125.850 ;
        RECT 34.600 125.555 34.740 125.710 ;
        RECT 35.430 125.650 35.750 125.710 ;
        RECT 39.585 125.665 39.875 125.710 ;
        RECT 41.410 125.650 41.730 125.910 ;
        RECT 41.960 125.895 42.100 126.050 ;
        RECT 44.260 125.895 44.400 126.050 ;
        RECT 65.300 126.050 70.230 126.190 ;
        RECT 65.300 126.005 65.590 126.050 ;
        RECT 68.080 126.005 68.370 126.050 ;
        RECT 69.940 126.005 70.230 126.050 ;
        RECT 70.850 126.190 71.170 126.250 ;
        RECT 108.080 126.190 108.370 126.235 ;
        RECT 110.860 126.190 111.150 126.235 ;
        RECT 112.720 126.190 113.010 126.235 ;
        RECT 70.850 126.050 81.660 126.190 ;
        RECT 70.850 125.990 71.170 126.050 ;
        RECT 41.885 125.665 42.175 125.895 ;
        RECT 44.185 125.665 44.475 125.895 ;
        RECT 46.470 125.850 46.790 125.910 ;
        RECT 47.865 125.850 48.155 125.895 ;
        RECT 70.940 125.850 71.080 125.990 ;
        RECT 74.070 125.850 74.390 125.910 ;
        RECT 46.470 125.710 48.155 125.850 ;
        RECT 46.470 125.650 46.790 125.710 ;
        RECT 47.865 125.665 48.155 125.710 ;
        RECT 48.860 125.710 71.080 125.850 ;
        RECT 71.400 125.710 74.390 125.850 ;
        RECT 34.525 125.325 34.815 125.555 ;
        RECT 40.505 125.510 40.795 125.555 ;
        RECT 40.950 125.510 41.270 125.570 ;
        RECT 42.805 125.510 43.095 125.555 ;
        RECT 43.250 125.510 43.570 125.570 ;
        RECT 45.105 125.510 45.395 125.555 ;
        RECT 40.505 125.370 45.395 125.510 ;
        RECT 40.505 125.325 40.795 125.370 ;
        RECT 40.950 125.310 41.270 125.370 ;
        RECT 42.805 125.325 43.095 125.370 ;
        RECT 43.250 125.310 43.570 125.370 ;
        RECT 45.105 125.325 45.395 125.370 ;
        RECT 45.180 125.170 45.320 125.325 ;
        RECT 46.010 125.310 46.330 125.570 ;
        RECT 48.860 125.555 49.000 125.710 ;
        RECT 71.400 125.570 71.540 125.710 ;
        RECT 74.070 125.650 74.390 125.710 ;
        RECT 48.785 125.325 49.075 125.555 ;
        RECT 65.300 125.510 65.590 125.555 ;
        RECT 68.565 125.510 68.855 125.555 ;
        RECT 70.405 125.510 70.695 125.555 ;
        RECT 71.310 125.510 71.630 125.570 ;
        RECT 65.300 125.370 67.835 125.510 ;
        RECT 65.300 125.325 65.590 125.370 ;
        RECT 48.860 125.170 49.000 125.325 ;
        RECT 45.180 125.030 49.000 125.170 ;
        RECT 61.190 125.215 61.510 125.230 ;
        RECT 61.190 124.985 61.725 125.215 ;
        RECT 63.440 125.170 63.730 125.215 ;
        RECT 64.410 125.170 64.730 125.230 ;
        RECT 67.620 125.215 67.835 125.370 ;
        RECT 68.565 125.370 70.160 125.510 ;
        RECT 68.565 125.325 68.855 125.370 ;
        RECT 66.700 125.170 66.990 125.215 ;
        RECT 63.440 125.030 66.990 125.170 ;
        RECT 63.440 124.985 63.730 125.030 ;
        RECT 61.190 124.970 61.510 124.985 ;
        RECT 64.410 124.970 64.730 125.030 ;
        RECT 66.700 124.985 66.990 125.030 ;
        RECT 67.620 125.170 67.910 125.215 ;
        RECT 69.480 125.170 69.770 125.215 ;
        RECT 67.620 125.030 69.770 125.170 ;
        RECT 67.620 124.985 67.910 125.030 ;
        RECT 69.480 124.985 69.770 125.030 ;
        RECT 27.625 124.690 34.280 124.830 ;
        RECT 34.510 124.830 34.830 124.890 ;
        RECT 34.985 124.830 35.275 124.875 ;
        RECT 34.510 124.690 35.275 124.830 ;
        RECT 27.625 124.645 27.915 124.690 ;
        RECT 29.910 124.630 30.230 124.690 ;
        RECT 34.510 124.630 34.830 124.690 ;
        RECT 34.985 124.645 35.275 124.690 ;
        RECT 36.825 124.830 37.115 124.875 ;
        RECT 37.730 124.830 38.050 124.890 ;
        RECT 36.825 124.690 38.050 124.830 ;
        RECT 70.020 124.830 70.160 125.370 ;
        RECT 70.405 125.370 71.630 125.510 ;
        RECT 70.405 125.325 70.695 125.370 ;
        RECT 71.310 125.310 71.630 125.370 ;
        RECT 71.770 125.310 72.090 125.570 ;
        RECT 73.610 125.310 73.930 125.570 ;
        RECT 79.220 125.555 79.360 126.050 ;
        RECT 80.050 125.650 80.370 125.910 ;
        RECT 81.520 125.850 81.660 126.050 ;
        RECT 108.080 126.050 113.010 126.190 ;
        RECT 108.080 126.005 108.370 126.050 ;
        RECT 110.860 126.005 111.150 126.050 ;
        RECT 112.720 126.005 113.010 126.050 ;
        RECT 113.645 126.005 113.935 126.235 ;
        RECT 119.580 126.190 119.870 126.235 ;
        RECT 122.360 126.190 122.650 126.235 ;
        RECT 124.220 126.190 124.510 126.235 ;
        RECT 119.580 126.050 124.510 126.190 ;
        RECT 119.580 126.005 119.870 126.050 ;
        RECT 122.360 126.005 122.650 126.050 ;
        RECT 124.220 126.005 124.510 126.050 ;
        RECT 82.350 125.850 82.670 125.910 ;
        RECT 81.520 125.710 83.960 125.850 ;
        RECT 79.145 125.325 79.435 125.555 ;
        RECT 79.590 125.510 79.910 125.570 ;
        RECT 81.520 125.555 81.660 125.710 ;
        RECT 82.350 125.650 82.670 125.710 ;
        RECT 80.525 125.510 80.815 125.555 ;
        RECT 79.590 125.370 80.815 125.510 ;
        RECT 79.590 125.310 79.910 125.370 ;
        RECT 80.525 125.325 80.815 125.370 ;
        RECT 81.445 125.325 81.735 125.555 ;
        RECT 82.825 125.510 83.115 125.555 ;
        RECT 83.270 125.510 83.590 125.570 ;
        RECT 83.820 125.555 83.960 125.710 ;
        RECT 84.650 125.650 84.970 125.910 ;
        RECT 113.720 125.850 113.860 126.005 ;
        RECT 112.340 125.710 113.860 125.850 ;
        RECT 115.715 125.850 116.005 125.895 ;
        RECT 117.310 125.850 117.630 125.910 ;
        RECT 115.715 125.710 117.630 125.850 ;
        RECT 82.825 125.370 83.590 125.510 ;
        RECT 82.825 125.325 83.115 125.370 ;
        RECT 83.270 125.310 83.590 125.370 ;
        RECT 83.745 125.325 84.035 125.555 ;
        RECT 95.690 125.510 96.010 125.570 ;
        RECT 96.625 125.510 96.915 125.555 ;
        RECT 95.690 125.370 96.915 125.510 ;
        RECT 95.690 125.310 96.010 125.370 ;
        RECT 96.625 125.325 96.915 125.370 ;
        RECT 98.910 125.510 99.230 125.570 ;
        RECT 102.590 125.510 102.910 125.570 ;
        RECT 98.910 125.370 102.910 125.510 ;
        RECT 98.910 125.310 99.230 125.370 ;
        RECT 102.590 125.310 102.910 125.370 ;
        RECT 108.080 125.510 108.370 125.555 ;
        RECT 111.345 125.510 111.635 125.555 ;
        RECT 112.340 125.510 112.480 125.710 ;
        RECT 115.715 125.665 116.005 125.710 ;
        RECT 117.310 125.650 117.630 125.710 ;
        RECT 122.830 125.650 123.150 125.910 ;
        RECT 108.080 125.370 110.615 125.510 ;
        RECT 108.080 125.325 108.370 125.370 ;
        RECT 75.450 124.970 75.770 125.230 ;
        RECT 110.400 125.215 110.615 125.370 ;
        RECT 111.345 125.370 112.480 125.510 ;
        RECT 112.710 125.510 113.030 125.570 ;
        RECT 113.185 125.510 113.475 125.555 ;
        RECT 112.710 125.370 113.475 125.510 ;
        RECT 111.345 125.325 111.635 125.370 ;
        RECT 112.710 125.310 113.030 125.370 ;
        RECT 113.185 125.325 113.475 125.370 ;
        RECT 114.565 125.325 114.855 125.555 ;
        RECT 119.580 125.510 119.870 125.555 ;
        RECT 124.210 125.510 124.530 125.570 ;
        RECT 124.685 125.510 124.975 125.555 ;
        RECT 119.580 125.370 122.115 125.510 ;
        RECT 119.580 125.325 119.870 125.370 ;
        RECT 103.065 125.170 103.355 125.215 ;
        RECT 106.220 125.170 106.510 125.215 ;
        RECT 109.480 125.170 109.770 125.215 ;
        RECT 103.065 125.030 109.770 125.170 ;
        RECT 103.065 124.985 103.355 125.030 ;
        RECT 106.220 124.985 106.510 125.030 ;
        RECT 109.480 124.985 109.770 125.030 ;
        RECT 110.400 125.170 110.690 125.215 ;
        RECT 112.260 125.170 112.550 125.215 ;
        RECT 110.400 125.030 112.550 125.170 ;
        RECT 110.400 124.985 110.690 125.030 ;
        RECT 112.260 124.985 112.550 125.030 ;
        RECT 70.865 124.830 71.155 124.875 ;
        RECT 70.020 124.690 71.155 124.830 ;
        RECT 36.825 124.645 37.115 124.690 ;
        RECT 37.730 124.630 38.050 124.690 ;
        RECT 70.865 124.645 71.155 124.690 ;
        RECT 78.225 124.830 78.515 124.875 ;
        RECT 79.130 124.830 79.450 124.890 ;
        RECT 78.225 124.690 79.450 124.830 ;
        RECT 78.225 124.645 78.515 124.690 ;
        RECT 79.130 124.630 79.450 124.690 ;
        RECT 97.530 124.630 97.850 124.890 ;
        RECT 104.215 124.830 104.505 124.875 ;
        RECT 109.030 124.830 109.350 124.890 ;
        RECT 104.215 124.690 109.350 124.830 ;
        RECT 104.215 124.645 104.505 124.690 ;
        RECT 109.030 124.630 109.350 124.690 ;
        RECT 111.790 124.830 112.110 124.890 ;
        RECT 114.640 124.830 114.780 125.325 ;
        RECT 115.470 125.170 115.790 125.230 ;
        RECT 121.900 125.215 122.115 125.370 ;
        RECT 124.210 125.370 124.975 125.510 ;
        RECT 124.210 125.310 124.530 125.370 ;
        RECT 124.685 125.325 124.975 125.370 ;
        RECT 126.065 125.325 126.355 125.555 ;
        RECT 117.720 125.170 118.010 125.215 ;
        RECT 120.980 125.170 121.270 125.215 ;
        RECT 115.470 125.030 121.270 125.170 ;
        RECT 115.470 124.970 115.790 125.030 ;
        RECT 117.720 124.985 118.010 125.030 ;
        RECT 120.980 124.985 121.270 125.030 ;
        RECT 121.900 125.170 122.190 125.215 ;
        RECT 123.760 125.170 124.050 125.215 ;
        RECT 121.900 125.030 124.050 125.170 ;
        RECT 121.900 124.985 122.190 125.030 ;
        RECT 123.760 124.985 124.050 125.030 ;
        RECT 111.790 124.690 114.780 124.830 ;
        RECT 119.150 124.830 119.470 124.890 ;
        RECT 126.140 124.830 126.280 125.325 ;
        RECT 119.150 124.690 126.280 124.830 ;
        RECT 111.790 124.630 112.110 124.690 ;
        RECT 119.150 124.630 119.470 124.690 ;
        RECT 14.660 124.010 127.820 124.490 ;
        RECT 16.355 123.810 16.645 123.855 ;
        RECT 23.470 123.810 23.790 123.870 ;
        RECT 16.355 123.670 23.790 123.810 ;
        RECT 16.355 123.625 16.645 123.670 ;
        RECT 23.470 123.610 23.790 123.670 ;
        RECT 30.370 123.610 30.690 123.870 ;
        RECT 34.510 123.810 34.830 123.870 ;
        RECT 46.470 123.810 46.790 123.870 ;
        RECT 52.465 123.810 52.755 123.855 ;
        RECT 34.510 123.670 52.755 123.810 ;
        RECT 34.510 123.610 34.830 123.670 ;
        RECT 46.470 123.610 46.790 123.670 ;
        RECT 52.465 123.625 52.755 123.670 ;
        RECT 61.190 123.810 61.510 123.870 ;
        RECT 63.950 123.810 64.270 123.870 ;
        RECT 64.885 123.810 65.175 123.855 ;
        RECT 61.190 123.670 65.175 123.810 ;
        RECT 61.190 123.610 61.510 123.670 ;
        RECT 63.950 123.610 64.270 123.670 ;
        RECT 64.885 123.625 65.175 123.670 ;
        RECT 65.330 123.610 65.650 123.870 ;
        RECT 67.185 123.810 67.475 123.855 ;
        RECT 71.770 123.810 72.090 123.870 ;
        RECT 67.185 123.670 72.090 123.810 ;
        RECT 67.185 123.625 67.475 123.670 ;
        RECT 71.770 123.610 72.090 123.670 ;
        RECT 83.730 123.810 84.050 123.870 ;
        RECT 93.865 123.810 94.155 123.855 ;
        RECT 83.730 123.670 94.155 123.810 ;
        RECT 83.730 123.610 84.050 123.670 ;
        RECT 93.865 123.625 94.155 123.670 ;
        RECT 95.690 123.610 96.010 123.870 ;
        RECT 101.210 123.810 101.530 123.870 ;
        RECT 107.665 123.810 107.955 123.855 ;
        RECT 98.080 123.670 107.955 123.810 ;
        RECT 18.360 123.470 18.650 123.515 ;
        RECT 19.790 123.470 20.110 123.530 ;
        RECT 21.620 123.470 21.910 123.515 ;
        RECT 18.360 123.330 21.910 123.470 ;
        RECT 18.360 123.285 18.650 123.330 ;
        RECT 19.790 123.270 20.110 123.330 ;
        RECT 21.620 123.285 21.910 123.330 ;
        RECT 22.540 123.470 22.830 123.515 ;
        RECT 24.400 123.470 24.690 123.515 ;
        RECT 22.540 123.330 24.690 123.470 ;
        RECT 22.540 123.285 22.830 123.330 ;
        RECT 24.400 123.285 24.690 123.330 ;
        RECT 20.220 123.130 20.510 123.175 ;
        RECT 22.540 123.130 22.755 123.285 ;
        RECT 20.220 122.990 22.755 123.130 ;
        RECT 24.850 123.130 25.170 123.190 ;
        RECT 25.325 123.130 25.615 123.175 ;
        RECT 30.460 123.130 30.600 123.610 ;
        RECT 79.130 123.470 79.450 123.530 ;
        RECT 80.050 123.470 80.370 123.530 ;
        RECT 79.130 123.330 80.370 123.470 ;
        RECT 79.130 123.270 79.450 123.330 ;
        RECT 80.050 123.270 80.370 123.330 ;
        RECT 24.850 122.990 30.600 123.130 ;
        RECT 20.220 122.945 20.510 122.990 ;
        RECT 24.850 122.930 25.170 122.990 ;
        RECT 25.325 122.945 25.615 122.990 ;
        RECT 36.810 122.930 37.130 123.190 ;
        RECT 52.450 123.130 52.770 123.190 ;
        RECT 52.925 123.130 53.215 123.175 ;
        RECT 52.450 122.990 53.215 123.130 ;
        RECT 52.450 122.930 52.770 122.990 ;
        RECT 52.925 122.945 53.215 122.990 ;
        RECT 58.445 123.130 58.735 123.175 ;
        RECT 60.270 123.130 60.590 123.190 ;
        RECT 58.445 122.990 60.590 123.130 ;
        RECT 58.445 122.945 58.735 122.990 ;
        RECT 60.270 122.930 60.590 122.990 ;
        RECT 61.190 123.130 61.510 123.190 ;
        RECT 61.665 123.130 61.955 123.175 ;
        RECT 71.310 123.130 71.630 123.190 ;
        RECT 84.205 123.130 84.495 123.175 ;
        RECT 61.190 122.990 71.630 123.130 ;
        RECT 61.190 122.930 61.510 122.990 ;
        RECT 61.665 122.945 61.955 122.990 ;
        RECT 71.310 122.930 71.630 122.990 ;
        RECT 79.680 122.990 84.495 123.130 ;
        RECT 79.680 122.850 79.820 122.990 ;
        RECT 84.205 122.945 84.495 122.990 ;
        RECT 90.630 122.930 90.950 123.190 ;
        RECT 93.405 123.130 93.695 123.175 ;
        RECT 96.395 123.130 96.685 123.175 ;
        RECT 98.080 123.130 98.220 123.670 ;
        RECT 101.210 123.610 101.530 123.670 ;
        RECT 107.665 123.625 107.955 123.670 ;
        RECT 108.125 123.810 108.415 123.855 ;
        RECT 109.030 123.810 109.350 123.870 ;
        RECT 108.125 123.670 109.350 123.810 ;
        RECT 108.125 123.625 108.415 123.670 ;
        RECT 109.030 123.610 109.350 123.670 ;
        RECT 116.850 123.610 117.170 123.870 ;
        RECT 117.310 123.610 117.630 123.870 ;
        RECT 119.165 123.625 119.455 123.855 ;
        RECT 121.925 123.810 122.215 123.855 ;
        RECT 122.830 123.810 123.150 123.870 ;
        RECT 121.925 123.670 123.150 123.810 ;
        RECT 121.925 123.625 122.215 123.670 ;
        RECT 98.400 123.470 98.690 123.515 ;
        RECT 98.910 123.470 99.230 123.530 ;
        RECT 101.660 123.470 101.950 123.515 ;
        RECT 98.400 123.330 101.950 123.470 ;
        RECT 98.400 123.285 98.690 123.330 ;
        RECT 98.910 123.270 99.230 123.330 ;
        RECT 101.660 123.285 101.950 123.330 ;
        RECT 102.580 123.470 102.870 123.515 ;
        RECT 104.440 123.470 104.730 123.515 ;
        RECT 102.580 123.330 104.730 123.470 ;
        RECT 102.580 123.285 102.870 123.330 ;
        RECT 104.440 123.285 104.730 123.330 ;
        RECT 93.405 122.990 98.220 123.130 ;
        RECT 100.260 123.130 100.550 123.175 ;
        RECT 102.580 123.130 102.795 123.285 ;
        RECT 100.260 122.990 102.795 123.130 ;
        RECT 93.405 122.945 93.695 122.990 ;
        RECT 96.395 122.945 96.685 122.990 ;
        RECT 100.260 122.945 100.550 122.990 ;
        RECT 103.510 122.930 103.830 123.190 ;
        RECT 112.265 123.130 112.555 123.175 ;
        RECT 112.710 123.130 113.030 123.190 ;
        RECT 112.265 122.990 113.030 123.130 ;
        RECT 119.240 123.130 119.380 123.625 ;
        RECT 122.830 123.610 123.150 123.670 ;
        RECT 121.005 123.130 121.295 123.175 ;
        RECT 119.240 122.990 121.295 123.130 ;
        RECT 112.265 122.945 112.555 122.990 ;
        RECT 112.710 122.930 113.030 122.990 ;
        RECT 121.005 122.945 121.295 122.990 ;
        RECT 19.330 122.790 19.650 122.850 ;
        RECT 23.485 122.790 23.775 122.835 ;
        RECT 19.330 122.650 23.775 122.790 ;
        RECT 19.330 122.590 19.650 122.650 ;
        RECT 23.485 122.605 23.775 122.650 ;
        RECT 50.610 122.790 50.930 122.850 ;
        RECT 51.545 122.790 51.835 122.835 ;
        RECT 50.610 122.650 51.835 122.790 ;
        RECT 50.610 122.590 50.930 122.650 ;
        RECT 51.545 122.605 51.835 122.650 ;
        RECT 53.830 122.790 54.150 122.850 ;
        RECT 57.065 122.790 57.355 122.835 ;
        RECT 53.830 122.650 57.355 122.790 ;
        RECT 53.830 122.590 54.150 122.650 ;
        RECT 57.065 122.605 57.355 122.650 ;
        RECT 64.410 122.790 64.730 122.850 ;
        RECT 65.790 122.790 66.110 122.850 ;
        RECT 64.410 122.650 66.110 122.790 ;
        RECT 64.410 122.590 64.730 122.650 ;
        RECT 65.790 122.590 66.110 122.650 ;
        RECT 75.450 122.790 75.770 122.850 ;
        RECT 78.685 122.790 78.975 122.835 ;
        RECT 75.450 122.650 78.975 122.790 ;
        RECT 75.450 122.590 75.770 122.650 ;
        RECT 78.685 122.605 78.975 122.650 ;
        RECT 20.220 122.450 20.510 122.495 ;
        RECT 23.000 122.450 23.290 122.495 ;
        RECT 24.860 122.450 25.150 122.495 ;
        RECT 20.220 122.310 25.150 122.450 ;
        RECT 78.760 122.450 78.900 122.605 ;
        RECT 79.590 122.590 79.910 122.850 ;
        RECT 82.825 122.790 83.115 122.835 ;
        RECT 90.170 122.790 90.490 122.850 ;
        RECT 92.485 122.790 92.775 122.835 ;
        RECT 82.825 122.650 92.775 122.790 ;
        RECT 82.825 122.605 83.115 122.650 ;
        RECT 82.900 122.450 83.040 122.605 ;
        RECT 90.170 122.590 90.490 122.650 ;
        RECT 92.485 122.605 92.775 122.650 ;
        RECT 98.450 122.790 98.770 122.850 ;
        RECT 105.365 122.790 105.655 122.835 ;
        RECT 98.450 122.650 105.655 122.790 ;
        RECT 98.450 122.590 98.770 122.650 ;
        RECT 105.365 122.605 105.655 122.650 ;
        RECT 108.570 122.790 108.890 122.850 ;
        RECT 109.950 122.790 110.270 122.850 ;
        RECT 115.945 122.790 116.235 122.835 ;
        RECT 108.570 122.650 116.235 122.790 ;
        RECT 108.570 122.590 108.890 122.650 ;
        RECT 109.950 122.590 110.270 122.650 ;
        RECT 115.945 122.605 116.235 122.650 ;
        RECT 78.760 122.310 83.040 122.450 ;
        RECT 100.260 122.450 100.550 122.495 ;
        RECT 103.040 122.450 103.330 122.495 ;
        RECT 104.900 122.450 105.190 122.495 ;
        RECT 100.260 122.310 105.190 122.450 ;
        RECT 20.220 122.265 20.510 122.310 ;
        RECT 23.000 122.265 23.290 122.310 ;
        RECT 24.860 122.265 25.150 122.310 ;
        RECT 100.260 122.265 100.550 122.310 ;
        RECT 103.040 122.265 103.330 122.310 ;
        RECT 104.900 122.265 105.190 122.310 ;
        RECT 54.765 122.110 55.055 122.155 ;
        RECT 55.670 122.110 55.990 122.170 ;
        RECT 54.765 121.970 55.990 122.110 ;
        RECT 54.765 121.925 55.055 121.970 ;
        RECT 55.670 121.910 55.990 121.970 ;
        RECT 81.905 122.110 82.195 122.155 ;
        RECT 82.810 122.110 83.130 122.170 ;
        RECT 81.905 121.970 83.130 122.110 ;
        RECT 81.905 121.925 82.195 121.970 ;
        RECT 82.810 121.910 83.130 121.970 ;
        RECT 86.045 122.110 86.335 122.155 ;
        RECT 88.790 122.110 89.110 122.170 ;
        RECT 86.045 121.970 89.110 122.110 ;
        RECT 86.045 121.925 86.335 121.970 ;
        RECT 88.790 121.910 89.110 121.970 ;
        RECT 91.090 121.910 91.410 122.170 ;
        RECT 105.810 121.910 106.130 122.170 ;
        RECT 14.660 121.290 127.820 121.770 ;
        RECT 19.790 120.890 20.110 121.150 ;
        RECT 35.430 121.090 35.750 121.150 ;
        RECT 36.135 121.090 36.425 121.135 ;
        RECT 35.430 120.950 36.425 121.090 ;
        RECT 35.430 120.890 35.750 120.950 ;
        RECT 36.135 120.905 36.425 120.950 ;
        RECT 40.490 121.090 40.810 121.150 ;
        RECT 78.455 121.090 78.745 121.135 ;
        RECT 79.590 121.090 79.910 121.150 ;
        RECT 40.490 120.950 71.310 121.090 ;
        RECT 40.490 120.890 40.810 120.950 ;
        RECT 25.330 120.750 25.620 120.795 ;
        RECT 27.190 120.750 27.480 120.795 ;
        RECT 29.970 120.750 30.260 120.795 ;
        RECT 25.330 120.610 30.260 120.750 ;
        RECT 25.330 120.565 25.620 120.610 ;
        RECT 27.190 120.565 27.480 120.610 ;
        RECT 29.970 120.565 30.260 120.610 ;
        RECT 40.000 120.750 40.290 120.795 ;
        RECT 42.780 120.750 43.070 120.795 ;
        RECT 44.640 120.750 44.930 120.795 ;
        RECT 50.610 120.750 50.930 120.810 ;
        RECT 40.000 120.610 44.930 120.750 ;
        RECT 40.000 120.565 40.290 120.610 ;
        RECT 42.780 120.565 43.070 120.610 ;
        RECT 44.640 120.565 44.930 120.610 ;
        RECT 47.020 120.610 50.930 120.750 ;
        RECT 24.850 120.210 25.170 120.470 ;
        RECT 33.590 120.455 33.910 120.470 ;
        RECT 33.590 120.410 34.125 120.455 ;
        RECT 36.350 120.410 36.670 120.470 ;
        RECT 33.590 120.270 36.670 120.410 ;
        RECT 33.590 120.225 34.125 120.270 ;
        RECT 33.590 120.210 33.910 120.225 ;
        RECT 36.350 120.210 36.670 120.270 ;
        RECT 40.490 120.410 40.810 120.470 ;
        RECT 47.020 120.455 47.160 120.610 ;
        RECT 50.610 120.550 50.930 120.610 ;
        RECT 67.185 120.565 67.475 120.795 ;
        RECT 43.265 120.410 43.555 120.455 ;
        RECT 40.490 120.270 43.555 120.410 ;
        RECT 40.490 120.210 40.810 120.270 ;
        RECT 43.265 120.225 43.555 120.270 ;
        RECT 46.945 120.225 47.235 120.455 ;
        RECT 47.405 120.410 47.695 120.455 ;
        RECT 52.450 120.410 52.770 120.470 ;
        RECT 47.405 120.270 52.770 120.410 ;
        RECT 47.405 120.225 47.695 120.270 ;
        RECT 52.450 120.210 52.770 120.270 ;
        RECT 61.190 120.210 61.510 120.470 ;
        RECT 64.410 120.210 64.730 120.470 ;
        RECT 64.870 120.210 65.190 120.470 ;
        RECT 20.250 119.870 20.570 120.130 ;
        RECT 23.010 119.870 23.330 120.130 ;
        RECT 26.690 119.870 27.010 120.130 ;
        RECT 29.970 120.070 30.260 120.115 ;
        RECT 27.725 119.930 30.260 120.070 ;
        RECT 22.550 119.730 22.870 119.790 ;
        RECT 27.725 119.775 27.940 119.930 ;
        RECT 29.970 119.885 30.260 119.930 ;
        RECT 34.525 120.070 34.815 120.115 ;
        RECT 35.890 120.070 36.210 120.130 ;
        RECT 34.525 119.930 36.210 120.070 ;
        RECT 34.525 119.885 34.815 119.930 ;
        RECT 35.890 119.870 36.210 119.930 ;
        RECT 40.000 120.070 40.290 120.115 ;
        RECT 45.105 120.070 45.395 120.115 ;
        RECT 46.470 120.070 46.790 120.130 ;
        RECT 40.000 119.930 42.535 120.070 ;
        RECT 40.000 119.885 40.290 119.930 ;
        RECT 25.790 119.730 26.080 119.775 ;
        RECT 27.650 119.730 27.940 119.775 ;
        RECT 22.550 119.590 24.620 119.730 ;
        RECT 22.550 119.530 22.870 119.590 ;
        RECT 23.930 119.190 24.250 119.450 ;
        RECT 24.480 119.390 24.620 119.590 ;
        RECT 25.790 119.590 27.940 119.730 ;
        RECT 25.790 119.545 26.080 119.590 ;
        RECT 27.650 119.545 27.940 119.590 ;
        RECT 28.530 119.775 28.850 119.790 ;
        RECT 28.530 119.730 28.860 119.775 ;
        RECT 31.830 119.730 32.120 119.775 ;
        RECT 28.530 119.590 32.120 119.730 ;
        RECT 28.530 119.545 28.860 119.590 ;
        RECT 31.830 119.545 32.120 119.590 ;
        RECT 34.050 119.730 34.370 119.790 ;
        RECT 42.320 119.775 42.535 119.930 ;
        RECT 45.105 119.930 46.790 120.070 ;
        RECT 45.105 119.885 45.395 119.930 ;
        RECT 46.470 119.870 46.790 119.930 ;
        RECT 52.910 119.870 53.230 120.130 ;
        RECT 63.950 120.070 64.270 120.130 ;
        RECT 65.345 120.070 65.635 120.115 ;
        RECT 63.950 119.930 65.635 120.070 ;
        RECT 67.260 120.070 67.400 120.565 ;
        RECT 68.105 120.070 68.395 120.115 ;
        RECT 67.260 119.930 68.395 120.070 ;
        RECT 71.170 120.070 71.310 120.950 ;
        RECT 78.455 120.950 79.910 121.090 ;
        RECT 78.455 120.905 78.745 120.950 ;
        RECT 79.590 120.890 79.910 120.950 ;
        RECT 83.730 121.090 84.050 121.150 ;
        RECT 89.955 121.090 90.245 121.135 ;
        RECT 83.730 120.950 90.245 121.090 ;
        RECT 83.730 120.890 84.050 120.950 ;
        RECT 89.955 120.905 90.245 120.950 ;
        RECT 103.510 121.090 103.830 121.150 ;
        RECT 103.985 121.090 104.275 121.135 ;
        RECT 103.510 120.950 104.275 121.090 ;
        RECT 103.510 120.890 103.830 120.950 ;
        RECT 103.985 120.905 104.275 120.950 ;
        RECT 82.320 120.750 82.610 120.795 ;
        RECT 85.100 120.750 85.390 120.795 ;
        RECT 86.960 120.750 87.250 120.795 ;
        RECT 82.320 120.610 87.250 120.750 ;
        RECT 82.320 120.565 82.610 120.610 ;
        RECT 85.100 120.565 85.390 120.610 ;
        RECT 86.960 120.565 87.250 120.610 ;
        RECT 93.820 120.750 94.110 120.795 ;
        RECT 96.600 120.750 96.890 120.795 ;
        RECT 98.460 120.750 98.750 120.795 ;
        RECT 93.820 120.610 98.750 120.750 ;
        RECT 93.820 120.565 94.110 120.610 ;
        RECT 96.600 120.565 96.890 120.610 ;
        RECT 98.460 120.565 98.750 120.610 ;
        RECT 86.030 120.410 86.350 120.470 ;
        RECT 87.425 120.410 87.715 120.455 ;
        RECT 97.085 120.410 97.375 120.455 ;
        RECT 97.530 120.410 97.850 120.470 ;
        RECT 86.030 120.270 96.840 120.410 ;
        RECT 86.030 120.210 86.350 120.270 ;
        RECT 87.425 120.225 87.715 120.270 ;
        RECT 76.845 120.070 77.135 120.115 ;
        RECT 71.170 119.930 77.135 120.070 ;
        RECT 63.950 119.870 64.270 119.930 ;
        RECT 65.345 119.885 65.635 119.930 ;
        RECT 68.105 119.885 68.395 119.930 ;
        RECT 76.845 119.885 77.135 119.930 ;
        RECT 82.320 120.070 82.610 120.115 ;
        RECT 85.585 120.070 85.875 120.115 ;
        RECT 82.320 119.930 84.855 120.070 ;
        RECT 82.320 119.885 82.610 119.930 ;
        RECT 38.140 119.730 38.430 119.775 ;
        RECT 41.400 119.730 41.690 119.775 ;
        RECT 34.050 119.590 41.690 119.730 ;
        RECT 28.530 119.530 28.850 119.545 ;
        RECT 34.050 119.530 34.370 119.590 ;
        RECT 38.140 119.545 38.430 119.590 ;
        RECT 41.400 119.545 41.690 119.590 ;
        RECT 42.320 119.730 42.610 119.775 ;
        RECT 44.180 119.730 44.470 119.775 ;
        RECT 42.320 119.590 44.470 119.730 ;
        RECT 42.320 119.545 42.610 119.590 ;
        RECT 44.180 119.545 44.470 119.590 ;
        RECT 29.910 119.390 30.230 119.450 ;
        RECT 24.480 119.250 30.230 119.390 ;
        RECT 29.910 119.190 30.230 119.250 ;
        RECT 34.970 119.190 35.290 119.450 ;
        RECT 45.550 119.390 45.870 119.450 ;
        RECT 47.865 119.390 48.155 119.435 ;
        RECT 45.550 119.250 48.155 119.390 ;
        RECT 45.550 119.190 45.870 119.250 ;
        RECT 47.865 119.205 48.155 119.250 ;
        RECT 49.690 119.190 50.010 119.450 ;
        RECT 69.010 119.190 69.330 119.450 ;
        RECT 76.920 119.390 77.060 119.885 ;
        RECT 84.640 119.775 84.855 119.930 ;
        RECT 85.585 119.930 88.100 120.070 ;
        RECT 85.585 119.885 85.875 119.930 ;
        RECT 77.305 119.730 77.595 119.775 ;
        RECT 80.460 119.730 80.750 119.775 ;
        RECT 83.720 119.730 84.010 119.775 ;
        RECT 77.305 119.590 84.010 119.730 ;
        RECT 77.305 119.545 77.595 119.590 ;
        RECT 80.460 119.545 80.750 119.590 ;
        RECT 83.720 119.545 84.010 119.590 ;
        RECT 84.640 119.730 84.930 119.775 ;
        RECT 86.500 119.730 86.790 119.775 ;
        RECT 84.640 119.590 86.790 119.730 ;
        RECT 84.640 119.545 84.930 119.590 ;
        RECT 86.500 119.545 86.790 119.590 ;
        RECT 87.410 119.390 87.730 119.450 ;
        RECT 87.960 119.435 88.100 119.930 ;
        RECT 88.790 119.870 89.110 120.130 ;
        RECT 93.820 120.070 94.110 120.115 ;
        RECT 96.700 120.070 96.840 120.270 ;
        RECT 97.085 120.270 97.850 120.410 ;
        RECT 97.085 120.225 97.375 120.270 ;
        RECT 97.530 120.210 97.850 120.270 ;
        RECT 98.450 120.070 98.770 120.130 ;
        RECT 98.925 120.070 99.215 120.115 ;
        RECT 100.305 120.070 100.595 120.115 ;
        RECT 93.820 119.930 96.355 120.070 ;
        RECT 96.700 119.930 100.595 120.070 ;
        RECT 93.820 119.885 94.110 119.930 ;
        RECT 91.090 119.730 91.410 119.790 ;
        RECT 96.140 119.775 96.355 119.930 ;
        RECT 98.450 119.870 98.770 119.930 ;
        RECT 98.925 119.885 99.215 119.930 ;
        RECT 100.305 119.885 100.595 119.930 ;
        RECT 104.905 120.070 105.195 120.115 ;
        RECT 105.810 120.070 106.130 120.130 ;
        RECT 104.905 119.930 106.130 120.070 ;
        RECT 104.905 119.885 105.195 119.930 ;
        RECT 105.810 119.870 106.130 119.930 ;
        RECT 113.170 120.070 113.490 120.130 ;
        RECT 118.245 120.070 118.535 120.115 ;
        RECT 113.170 119.930 118.535 120.070 ;
        RECT 113.170 119.870 113.490 119.930 ;
        RECT 118.245 119.885 118.535 119.930 ;
        RECT 119.625 119.885 119.915 120.115 ;
        RECT 91.960 119.730 92.250 119.775 ;
        RECT 95.220 119.730 95.510 119.775 ;
        RECT 91.090 119.590 95.510 119.730 ;
        RECT 91.090 119.530 91.410 119.590 ;
        RECT 91.960 119.545 92.250 119.590 ;
        RECT 95.220 119.545 95.510 119.590 ;
        RECT 96.140 119.730 96.430 119.775 ;
        RECT 98.000 119.730 98.290 119.775 ;
        RECT 96.140 119.590 98.290 119.730 ;
        RECT 96.140 119.545 96.430 119.590 ;
        RECT 98.000 119.545 98.290 119.590 ;
        RECT 114.090 119.730 114.410 119.790 ;
        RECT 119.700 119.730 119.840 119.885 ;
        RECT 114.090 119.590 119.840 119.730 ;
        RECT 114.090 119.530 114.410 119.590 ;
        RECT 76.920 119.250 87.730 119.390 ;
        RECT 87.410 119.190 87.730 119.250 ;
        RECT 87.885 119.205 88.175 119.435 ;
        RECT 90.170 119.390 90.490 119.450 ;
        RECT 105.810 119.390 106.130 119.450 ;
        RECT 108.570 119.390 108.890 119.450 ;
        RECT 90.170 119.250 108.890 119.390 ;
        RECT 90.170 119.190 90.490 119.250 ;
        RECT 105.810 119.190 106.130 119.250 ;
        RECT 108.570 119.190 108.890 119.250 ;
        RECT 118.690 119.190 119.010 119.450 ;
        RECT 120.545 119.390 120.835 119.435 ;
        RECT 122.370 119.390 122.690 119.450 ;
        RECT 120.545 119.250 122.690 119.390 ;
        RECT 120.545 119.205 120.835 119.250 ;
        RECT 122.370 119.190 122.690 119.250 ;
        RECT 14.660 118.570 127.820 119.050 ;
        RECT 19.805 118.370 20.095 118.415 ;
        RECT 32.225 118.370 32.515 118.415 ;
        RECT 34.050 118.370 34.370 118.430 ;
        RECT 19.805 118.230 30.600 118.370 ;
        RECT 19.805 118.185 20.095 118.230 ;
        RECT 19.345 118.030 19.635 118.075 ;
        RECT 22.550 118.030 22.870 118.090 ;
        RECT 25.770 118.075 26.090 118.090 ;
        RECT 19.345 117.890 22.870 118.030 ;
        RECT 19.345 117.845 19.635 117.890 ;
        RECT 22.550 117.830 22.870 117.890 ;
        RECT 23.030 118.030 23.320 118.075 ;
        RECT 24.890 118.030 25.180 118.075 ;
        RECT 23.030 117.890 25.180 118.030 ;
        RECT 23.030 117.845 23.320 117.890 ;
        RECT 24.890 117.845 25.180 117.890 ;
        RECT 23.930 117.490 24.250 117.750 ;
        RECT 24.965 117.690 25.180 117.845 ;
        RECT 25.770 118.030 26.100 118.075 ;
        RECT 29.070 118.030 29.360 118.075 ;
        RECT 25.770 117.890 29.360 118.030 ;
        RECT 25.770 117.845 26.100 117.890 ;
        RECT 29.070 117.845 29.360 117.890 ;
        RECT 25.770 117.830 26.090 117.845 ;
        RECT 29.910 117.830 30.230 118.090 ;
        RECT 30.460 118.030 30.600 118.230 ;
        RECT 32.225 118.230 34.370 118.370 ;
        RECT 32.225 118.185 32.515 118.230 ;
        RECT 34.050 118.170 34.370 118.230 ;
        RECT 34.985 118.370 35.275 118.415 ;
        RECT 35.430 118.370 35.750 118.430 ;
        RECT 34.985 118.230 35.750 118.370 ;
        RECT 34.985 118.185 35.275 118.230 ;
        RECT 35.430 118.170 35.750 118.230 ;
        RECT 40.030 118.170 40.350 118.430 ;
        RECT 40.735 118.370 41.025 118.415 ;
        RECT 45.550 118.370 45.870 118.430 ;
        RECT 98.450 118.370 98.770 118.430 ;
        RECT 40.735 118.230 45.870 118.370 ;
        RECT 40.735 118.185 41.025 118.230 ;
        RECT 45.550 118.170 45.870 118.230 ;
        RECT 98.080 118.230 98.770 118.370 ;
        RECT 33.590 118.030 33.910 118.090 ;
        RECT 34.525 118.030 34.815 118.075 ;
        RECT 30.460 117.890 34.815 118.030 ;
        RECT 33.590 117.830 33.910 117.890 ;
        RECT 34.525 117.845 34.815 117.890 ;
        RECT 35.890 118.030 36.210 118.090 ;
        RECT 46.010 118.075 46.330 118.090 ;
        RECT 42.740 118.030 43.030 118.075 ;
        RECT 46.000 118.030 46.330 118.075 ;
        RECT 35.890 117.890 39.800 118.030 ;
        RECT 35.890 117.830 36.210 117.890 ;
        RECT 27.210 117.690 27.500 117.735 ;
        RECT 24.965 117.550 27.500 117.690 ;
        RECT 30.000 117.690 30.140 117.830 ;
        RECT 31.075 117.690 31.365 117.735 ;
        RECT 30.000 117.550 31.365 117.690 ;
        RECT 27.210 117.505 27.500 117.550 ;
        RECT 31.075 117.505 31.365 117.550 ;
        RECT 31.765 117.690 32.055 117.735 ;
        RECT 35.980 117.690 36.120 117.830 ;
        RECT 31.765 117.550 36.120 117.690 ;
        RECT 31.765 117.505 32.055 117.550 ;
        RECT 18.870 117.150 19.190 117.410 ;
        RECT 22.105 117.350 22.395 117.395 ;
        RECT 24.850 117.350 25.170 117.410 ;
        RECT 29.910 117.350 30.230 117.410 ;
        RECT 22.105 117.210 30.230 117.350 ;
        RECT 22.105 117.165 22.395 117.210 ;
        RECT 24.850 117.150 25.170 117.210 ;
        RECT 29.910 117.150 30.230 117.210 ;
        RECT 30.370 117.350 30.690 117.410 ;
        RECT 31.840 117.350 31.980 117.505 ;
        RECT 37.730 117.490 38.050 117.750 ;
        RECT 39.125 117.505 39.415 117.735 ;
        RECT 30.370 117.210 31.980 117.350 ;
        RECT 30.370 117.150 30.690 117.210 ;
        RECT 33.605 117.165 33.895 117.395 ;
        RECT 39.200 117.350 39.340 117.505 ;
        RECT 36.900 117.210 39.340 117.350 ;
        RECT 22.570 117.010 22.860 117.055 ;
        RECT 24.430 117.010 24.720 117.055 ;
        RECT 27.210 117.010 27.500 117.055 ;
        RECT 22.570 116.870 27.500 117.010 ;
        RECT 22.570 116.825 22.860 116.870 ;
        RECT 24.430 116.825 24.720 116.870 ;
        RECT 27.210 116.825 27.500 116.870 ;
        RECT 31.290 117.010 31.610 117.070 ;
        RECT 33.680 117.010 33.820 117.165 ;
        RECT 36.900 117.055 37.040 117.210 ;
        RECT 31.290 116.870 33.820 117.010 ;
        RECT 31.290 116.810 31.610 116.870 ;
        RECT 36.825 116.825 37.115 117.055 ;
        RECT 21.645 116.670 21.935 116.715 ;
        RECT 27.610 116.670 27.930 116.730 ;
        RECT 21.645 116.530 27.930 116.670 ;
        RECT 21.645 116.485 21.935 116.530 ;
        RECT 27.610 116.470 27.930 116.530 ;
        RECT 38.650 116.470 38.970 116.730 ;
        RECT 39.660 116.670 39.800 117.890 ;
        RECT 42.740 117.890 46.330 118.030 ;
        RECT 42.740 117.845 43.030 117.890 ;
        RECT 46.000 117.845 46.330 117.890 ;
        RECT 46.010 117.830 46.330 117.845 ;
        RECT 46.920 118.030 47.210 118.075 ;
        RECT 48.780 118.030 49.070 118.075 ;
        RECT 46.920 117.890 49.070 118.030 ;
        RECT 46.920 117.845 47.210 117.890 ;
        RECT 48.780 117.845 49.070 117.890 ;
        RECT 52.400 118.030 52.690 118.075 ;
        RECT 52.910 118.030 53.230 118.090 ;
        RECT 69.930 118.075 70.250 118.090 ;
        RECT 55.660 118.030 55.950 118.075 ;
        RECT 52.400 117.890 55.950 118.030 ;
        RECT 52.400 117.845 52.690 117.890 ;
        RECT 44.600 117.690 44.890 117.735 ;
        RECT 46.920 117.690 47.135 117.845 ;
        RECT 52.910 117.830 53.230 117.890 ;
        RECT 55.660 117.845 55.950 117.890 ;
        RECT 56.580 118.030 56.870 118.075 ;
        RECT 58.440 118.030 58.730 118.075 ;
        RECT 56.580 117.890 58.730 118.030 ;
        RECT 56.580 117.845 56.870 117.890 ;
        RECT 58.440 117.845 58.730 117.890 ;
        RECT 66.660 118.030 66.950 118.075 ;
        RECT 69.920 118.030 70.250 118.075 ;
        RECT 66.660 117.890 70.250 118.030 ;
        RECT 66.660 117.845 66.950 117.890 ;
        RECT 69.920 117.845 70.250 117.890 ;
        RECT 44.600 117.550 47.135 117.690 ;
        RECT 47.865 117.690 48.155 117.735 ;
        RECT 53.370 117.690 53.690 117.750 ;
        RECT 47.865 117.550 53.690 117.690 ;
        RECT 44.600 117.505 44.890 117.550 ;
        RECT 47.865 117.505 48.155 117.550 ;
        RECT 53.370 117.490 53.690 117.550 ;
        RECT 54.260 117.690 54.550 117.735 ;
        RECT 56.580 117.690 56.795 117.845 ;
        RECT 69.930 117.830 70.250 117.845 ;
        RECT 70.840 118.030 71.130 118.075 ;
        RECT 72.700 118.030 72.990 118.075 ;
        RECT 70.840 117.890 72.990 118.030 ;
        RECT 70.840 117.845 71.130 117.890 ;
        RECT 72.700 117.845 72.990 117.890 ;
        RECT 78.620 118.030 78.910 118.075 ;
        RECT 80.050 118.030 80.370 118.090 ;
        RECT 81.880 118.030 82.170 118.075 ;
        RECT 78.620 117.890 82.170 118.030 ;
        RECT 78.620 117.845 78.910 117.890 ;
        RECT 54.260 117.550 56.795 117.690 ;
        RECT 59.365 117.690 59.655 117.735 ;
        RECT 61.190 117.690 61.510 117.750 ;
        RECT 59.365 117.550 61.510 117.690 ;
        RECT 54.260 117.505 54.550 117.550 ;
        RECT 59.365 117.505 59.655 117.550 ;
        RECT 61.190 117.490 61.510 117.550 ;
        RECT 68.520 117.690 68.810 117.735 ;
        RECT 70.840 117.690 71.055 117.845 ;
        RECT 80.050 117.830 80.370 117.890 ;
        RECT 81.880 117.845 82.170 117.890 ;
        RECT 82.800 118.030 83.090 118.075 ;
        RECT 84.660 118.030 84.950 118.075 ;
        RECT 82.800 117.890 84.950 118.030 ;
        RECT 82.800 117.845 83.090 117.890 ;
        RECT 84.660 117.845 84.950 117.890 ;
        RECT 68.520 117.550 71.055 117.690 ;
        RECT 73.625 117.690 73.915 117.735 ;
        RECT 74.070 117.690 74.390 117.750 ;
        RECT 73.625 117.550 74.390 117.690 ;
        RECT 68.520 117.505 68.810 117.550 ;
        RECT 73.625 117.505 73.915 117.550 ;
        RECT 74.070 117.490 74.390 117.550 ;
        RECT 80.480 117.690 80.770 117.735 ;
        RECT 82.800 117.690 83.015 117.845 ;
        RECT 89.250 117.830 89.570 118.090 ;
        RECT 98.080 118.075 98.220 118.230 ;
        RECT 98.450 118.170 98.770 118.230 ;
        RECT 98.910 118.170 99.230 118.430 ;
        RECT 106.730 118.370 107.050 118.430 ;
        RECT 109.490 118.370 109.810 118.430 ;
        RECT 111.805 118.370 112.095 118.415 ;
        RECT 106.730 118.230 112.095 118.370 ;
        RECT 106.730 118.170 107.050 118.230 ;
        RECT 109.490 118.170 109.810 118.230 ;
        RECT 111.805 118.185 112.095 118.230 ;
        RECT 114.090 118.170 114.410 118.430 ;
        RECT 115.255 118.370 115.545 118.415 ;
        RECT 115.930 118.370 116.250 118.430 ;
        RECT 114.640 118.230 116.250 118.370 ;
        RECT 98.005 117.845 98.295 118.075 ;
        RECT 112.265 118.030 112.555 118.075 ;
        RECT 114.640 118.030 114.780 118.230 ;
        RECT 115.255 118.185 115.545 118.230 ;
        RECT 115.930 118.170 116.250 118.230 ;
        RECT 112.265 117.890 114.780 118.030 ;
        RECT 117.260 118.030 117.550 118.075 ;
        RECT 118.690 118.030 119.010 118.090 ;
        RECT 120.520 118.030 120.810 118.075 ;
        RECT 117.260 117.890 120.810 118.030 ;
        RECT 112.265 117.845 112.555 117.890 ;
        RECT 117.260 117.845 117.550 117.890 ;
        RECT 118.690 117.830 119.010 117.890 ;
        RECT 120.520 117.845 120.810 117.890 ;
        RECT 121.440 118.030 121.730 118.075 ;
        RECT 123.300 118.030 123.590 118.075 ;
        RECT 121.440 117.890 123.590 118.030 ;
        RECT 121.440 117.845 121.730 117.890 ;
        RECT 123.300 117.845 123.590 117.890 ;
        RECT 80.480 117.550 83.015 117.690 ;
        RECT 85.585 117.690 85.875 117.735 ;
        RECT 86.030 117.690 86.350 117.750 ;
        RECT 85.585 117.550 86.350 117.690 ;
        RECT 80.480 117.505 80.770 117.550 ;
        RECT 85.585 117.505 85.875 117.550 ;
        RECT 86.030 117.490 86.350 117.550 ;
        RECT 87.410 117.690 87.730 117.750 ;
        RECT 90.630 117.690 90.950 117.750 ;
        RECT 98.465 117.690 98.755 117.735 ;
        RECT 87.410 117.550 98.755 117.690 ;
        RECT 87.410 117.490 87.730 117.550 ;
        RECT 90.630 117.490 90.950 117.550 ;
        RECT 98.465 117.505 98.755 117.550 ;
        RECT 102.590 117.690 102.910 117.750 ;
        RECT 103.525 117.690 103.815 117.735 ;
        RECT 106.285 117.690 106.575 117.735 ;
        RECT 102.590 117.550 103.815 117.690 ;
        RECT 102.590 117.490 102.910 117.550 ;
        RECT 103.525 117.505 103.815 117.550 ;
        RECT 104.060 117.550 106.575 117.690 ;
        RECT 46.470 117.350 46.790 117.410 ;
        RECT 49.705 117.350 49.995 117.395 ;
        RECT 46.470 117.210 49.995 117.350 ;
        RECT 46.470 117.150 46.790 117.210 ;
        RECT 49.705 117.165 49.995 117.210 ;
        RECT 50.395 117.350 50.685 117.395 ;
        RECT 52.450 117.350 52.770 117.410 ;
        RECT 50.395 117.210 52.770 117.350 ;
        RECT 50.395 117.165 50.685 117.210 ;
        RECT 52.450 117.150 52.770 117.210 ;
        RECT 57.510 117.150 57.830 117.410 ;
        RECT 71.770 117.150 72.090 117.410 ;
        RECT 83.730 117.150 84.050 117.410 ;
        RECT 84.650 117.350 84.970 117.410 ;
        RECT 104.060 117.350 104.200 117.550 ;
        RECT 106.285 117.505 106.575 117.550 ;
        RECT 119.120 117.690 119.410 117.735 ;
        RECT 121.440 117.690 121.655 117.845 ;
        RECT 119.120 117.550 121.655 117.690 ;
        RECT 119.120 117.505 119.410 117.550 ;
        RECT 122.370 117.490 122.690 117.750 ;
        RECT 84.650 117.210 104.200 117.350 ;
        RECT 105.810 117.350 106.130 117.410 ;
        RECT 110.885 117.350 111.175 117.395 ;
        RECT 105.810 117.210 111.175 117.350 ;
        RECT 84.650 117.150 84.970 117.210 ;
        RECT 105.810 117.150 106.130 117.210 ;
        RECT 110.885 117.165 111.175 117.210 ;
        RECT 124.210 117.150 124.530 117.410 ;
        RECT 44.600 117.010 44.890 117.055 ;
        RECT 47.380 117.010 47.670 117.055 ;
        RECT 49.240 117.010 49.530 117.055 ;
        RECT 44.600 116.870 49.530 117.010 ;
        RECT 44.600 116.825 44.890 116.870 ;
        RECT 47.380 116.825 47.670 116.870 ;
        RECT 49.240 116.825 49.530 116.870 ;
        RECT 54.260 117.010 54.550 117.055 ;
        RECT 57.040 117.010 57.330 117.055 ;
        RECT 58.900 117.010 59.190 117.055 ;
        RECT 54.260 116.870 59.190 117.010 ;
        RECT 54.260 116.825 54.550 116.870 ;
        RECT 57.040 116.825 57.330 116.870 ;
        RECT 58.900 116.825 59.190 116.870 ;
        RECT 68.520 117.010 68.810 117.055 ;
        RECT 71.300 117.010 71.590 117.055 ;
        RECT 73.160 117.010 73.450 117.055 ;
        RECT 68.520 116.870 73.450 117.010 ;
        RECT 68.520 116.825 68.810 116.870 ;
        RECT 71.300 116.825 71.590 116.870 ;
        RECT 73.160 116.825 73.450 116.870 ;
        RECT 80.480 117.010 80.770 117.055 ;
        RECT 83.260 117.010 83.550 117.055 ;
        RECT 85.120 117.010 85.410 117.055 ;
        RECT 80.480 116.870 85.410 117.010 ;
        RECT 80.480 116.825 80.770 116.870 ;
        RECT 83.260 116.825 83.550 116.870 ;
        RECT 85.120 116.825 85.410 116.870 ;
        RECT 119.120 117.010 119.410 117.055 ;
        RECT 121.900 117.010 122.190 117.055 ;
        RECT 123.760 117.010 124.050 117.055 ;
        RECT 119.120 116.870 124.050 117.010 ;
        RECT 119.120 116.825 119.410 116.870 ;
        RECT 121.900 116.825 122.190 116.870 ;
        RECT 123.760 116.825 124.050 116.870 ;
        RECT 53.830 116.670 54.150 116.730 ;
        RECT 39.660 116.530 54.150 116.670 ;
        RECT 53.830 116.470 54.150 116.530 ;
        RECT 64.655 116.670 64.945 116.715 ;
        RECT 66.250 116.670 66.570 116.730 ;
        RECT 64.655 116.530 66.570 116.670 ;
        RECT 64.655 116.485 64.945 116.530 ;
        RECT 66.250 116.470 66.570 116.530 ;
        RECT 76.615 116.670 76.905 116.715 ;
        RECT 79.130 116.670 79.450 116.730 ;
        RECT 76.615 116.530 79.450 116.670 ;
        RECT 76.615 116.485 76.905 116.530 ;
        RECT 79.130 116.470 79.450 116.530 ;
        RECT 87.870 116.470 88.190 116.730 ;
        RECT 103.970 116.470 104.290 116.730 ;
        RECT 108.585 116.670 108.875 116.715 ;
        RECT 109.490 116.670 109.810 116.730 ;
        RECT 108.585 116.530 109.810 116.670 ;
        RECT 108.585 116.485 108.875 116.530 ;
        RECT 109.490 116.470 109.810 116.530 ;
        RECT 14.660 115.850 127.820 116.330 ;
        RECT 25.325 115.650 25.615 115.695 ;
        RECT 25.770 115.650 26.090 115.710 ;
        RECT 25.325 115.510 26.090 115.650 ;
        RECT 25.325 115.465 25.615 115.510 ;
        RECT 25.770 115.450 26.090 115.510 ;
        RECT 26.690 115.450 27.010 115.710 ;
        RECT 32.455 115.650 32.745 115.695 ;
        RECT 34.510 115.650 34.830 115.710 ;
        RECT 32.455 115.510 34.830 115.650 ;
        RECT 32.455 115.465 32.745 115.510 ;
        RECT 34.510 115.450 34.830 115.510 ;
        RECT 46.010 115.650 46.330 115.710 ;
        RECT 51.545 115.650 51.835 115.695 ;
        RECT 46.010 115.510 51.835 115.650 ;
        RECT 46.010 115.450 46.330 115.510 ;
        RECT 51.545 115.465 51.835 115.510 ;
        RECT 52.910 115.450 53.230 115.710 ;
        RECT 53.370 115.650 53.690 115.710 ;
        RECT 53.845 115.650 54.135 115.695 ;
        RECT 53.370 115.510 54.135 115.650 ;
        RECT 53.370 115.450 53.690 115.510 ;
        RECT 53.845 115.465 54.135 115.510 ;
        RECT 56.605 115.650 56.895 115.695 ;
        RECT 57.510 115.650 57.830 115.710 ;
        RECT 56.605 115.510 57.830 115.650 ;
        RECT 56.605 115.465 56.895 115.510 ;
        RECT 57.510 115.450 57.830 115.510 ;
        RECT 62.815 115.650 63.105 115.695 ;
        RECT 64.870 115.650 65.190 115.710 ;
        RECT 62.815 115.510 65.190 115.650 ;
        RECT 62.815 115.465 63.105 115.510 ;
        RECT 64.870 115.450 65.190 115.510 ;
        RECT 69.930 115.650 70.250 115.710 ;
        RECT 72.705 115.650 72.995 115.695 ;
        RECT 69.930 115.510 72.995 115.650 ;
        RECT 69.930 115.450 70.250 115.510 ;
        RECT 72.705 115.465 72.995 115.510 ;
        RECT 80.050 115.450 80.370 115.710 ;
        RECT 83.730 115.450 84.050 115.710 ;
        RECT 84.650 115.650 84.970 115.710 ;
        RECT 88.115 115.650 88.405 115.695 ;
        RECT 84.650 115.510 88.405 115.650 ;
        RECT 84.650 115.450 84.970 115.510 ;
        RECT 88.115 115.465 88.405 115.510 ;
        RECT 104.675 115.650 104.965 115.695 ;
        RECT 106.730 115.650 107.050 115.710 ;
        RECT 104.675 115.510 107.050 115.650 ;
        RECT 104.675 115.465 104.965 115.510 ;
        RECT 106.730 115.450 107.050 115.510 ;
        RECT 23.025 115.310 23.315 115.355 ;
        RECT 28.530 115.310 28.850 115.370 ;
        RECT 23.025 115.170 28.850 115.310 ;
        RECT 23.025 115.125 23.315 115.170 ;
        RECT 28.530 115.110 28.850 115.170 ;
        RECT 36.320 115.310 36.610 115.355 ;
        RECT 39.100 115.310 39.390 115.355 ;
        RECT 40.960 115.310 41.250 115.355 ;
        RECT 36.320 115.170 41.250 115.310 ;
        RECT 36.320 115.125 36.610 115.170 ;
        RECT 39.100 115.125 39.390 115.170 ;
        RECT 40.960 115.125 41.250 115.170 ;
        RECT 66.680 115.310 66.970 115.355 ;
        RECT 69.460 115.310 69.750 115.355 ;
        RECT 71.320 115.310 71.610 115.355 ;
        RECT 66.680 115.170 71.610 115.310 ;
        RECT 66.680 115.125 66.970 115.170 ;
        RECT 69.460 115.125 69.750 115.170 ;
        RECT 71.320 115.125 71.610 115.170 ;
        RECT 91.980 115.310 92.270 115.355 ;
        RECT 94.760 115.310 95.050 115.355 ;
        RECT 96.620 115.310 96.910 115.355 ;
        RECT 91.980 115.170 96.910 115.310 ;
        RECT 91.980 115.125 92.270 115.170 ;
        RECT 94.760 115.125 95.050 115.170 ;
        RECT 96.620 115.125 96.910 115.170 ;
        RECT 108.540 115.310 108.830 115.355 ;
        RECT 111.320 115.310 111.610 115.355 ;
        RECT 113.180 115.310 113.470 115.355 ;
        RECT 108.540 115.170 113.470 115.310 ;
        RECT 108.540 115.125 108.830 115.170 ;
        RECT 111.320 115.125 111.610 115.170 ;
        RECT 113.180 115.125 113.470 115.170 ;
        RECT 18.870 114.970 19.190 115.030 ;
        RECT 24.390 114.970 24.710 115.030 ;
        RECT 30.370 114.970 30.690 115.030 ;
        RECT 18.870 114.830 24.710 114.970 ;
        RECT 18.870 114.770 19.190 114.830 ;
        RECT 24.390 114.770 24.710 114.830 ;
        RECT 24.940 114.830 30.690 114.970 ;
        RECT 20.250 114.630 20.570 114.690 ;
        RECT 24.940 114.675 25.080 114.830 ;
        RECT 30.370 114.770 30.690 114.830 ;
        RECT 38.650 114.970 38.970 115.030 ;
        RECT 39.585 114.970 39.875 115.015 ;
        RECT 38.650 114.830 39.875 114.970 ;
        RECT 38.650 114.770 38.970 114.830 ;
        RECT 39.585 114.785 39.875 114.830 ;
        RECT 49.690 114.970 50.010 115.030 ;
        RECT 69.010 114.970 69.330 115.030 ;
        RECT 69.945 114.970 70.235 115.015 ;
        RECT 49.690 114.830 54.980 114.970 ;
        RECT 49.690 114.770 50.010 114.830 ;
        RECT 22.565 114.630 22.855 114.675 ;
        RECT 24.865 114.630 25.155 114.675 ;
        RECT 20.250 114.490 25.155 114.630 ;
        RECT 20.250 114.430 20.570 114.490 ;
        RECT 22.565 114.445 22.855 114.490 ;
        RECT 24.865 114.445 25.155 114.490 ;
        RECT 27.610 114.430 27.930 114.690 ;
        RECT 36.320 114.630 36.610 114.675 ;
        RECT 41.425 114.630 41.715 114.675 ;
        RECT 46.470 114.630 46.790 114.690 ;
        RECT 36.320 114.490 38.855 114.630 ;
        RECT 36.320 114.445 36.610 114.490 ;
        RECT 34.460 114.290 34.750 114.335 ;
        RECT 34.970 114.290 35.290 114.350 ;
        RECT 38.640 114.335 38.855 114.490 ;
        RECT 41.425 114.490 46.790 114.630 ;
        RECT 41.425 114.445 41.715 114.490 ;
        RECT 46.470 114.430 46.790 114.490 ;
        RECT 52.005 114.630 52.295 114.675 ;
        RECT 52.465 114.630 52.755 114.675 ;
        RECT 53.830 114.630 54.150 114.690 ;
        RECT 54.840 114.675 54.980 114.830 ;
        RECT 69.010 114.830 70.235 114.970 ;
        RECT 69.010 114.770 69.330 114.830 ;
        RECT 69.945 114.785 70.235 114.830 ;
        RECT 71.785 114.970 72.075 115.015 ;
        RECT 74.070 114.970 74.390 115.030 ;
        RECT 87.410 114.970 87.730 115.030 ;
        RECT 71.785 114.830 74.390 114.970 ;
        RECT 71.785 114.785 72.075 114.830 ;
        RECT 74.070 114.770 74.390 114.830 ;
        RECT 79.680 114.830 87.730 114.970 ;
        RECT 52.005 114.490 54.150 114.630 ;
        RECT 52.005 114.445 52.295 114.490 ;
        RECT 52.465 114.445 52.755 114.490 ;
        RECT 53.830 114.430 54.150 114.490 ;
        RECT 54.765 114.445 55.055 114.675 ;
        RECT 55.670 114.430 55.990 114.690 ;
        RECT 60.270 114.630 60.590 114.690 ;
        RECT 61.205 114.630 61.495 114.675 ;
        RECT 60.270 114.490 61.495 114.630 ;
        RECT 60.270 114.430 60.590 114.490 ;
        RECT 61.205 114.445 61.495 114.490 ;
        RECT 66.680 114.630 66.970 114.675 ;
        RECT 66.680 114.490 69.215 114.630 ;
        RECT 66.680 114.445 66.970 114.490 ;
        RECT 69.000 114.335 69.215 114.490 ;
        RECT 73.150 114.430 73.470 114.690 ;
        RECT 79.680 114.675 79.820 114.830 ;
        RECT 87.410 114.770 87.730 114.830 ;
        RECT 97.085 114.970 97.375 115.015 ;
        RECT 98.450 114.970 98.770 115.030 ;
        RECT 97.085 114.830 98.770 114.970 ;
        RECT 97.085 114.785 97.375 114.830 ;
        RECT 98.450 114.770 98.770 114.830 ;
        RECT 113.645 114.970 113.935 115.015 ;
        RECT 124.210 114.970 124.530 115.030 ;
        RECT 113.645 114.830 124.530 114.970 ;
        RECT 113.645 114.785 113.935 114.830 ;
        RECT 124.210 114.770 124.530 114.830 ;
        RECT 79.605 114.445 79.895 114.675 ;
        RECT 82.810 114.430 83.130 114.690 ;
        RECT 91.980 114.630 92.270 114.675 ;
        RECT 91.980 114.490 94.515 114.630 ;
        RECT 91.980 114.445 92.270 114.490 ;
        RECT 37.720 114.290 38.010 114.335 ;
        RECT 34.460 114.150 38.010 114.290 ;
        RECT 34.460 114.105 34.750 114.150 ;
        RECT 34.970 114.090 35.290 114.150 ;
        RECT 37.720 114.105 38.010 114.150 ;
        RECT 38.640 114.290 38.930 114.335 ;
        RECT 40.500 114.290 40.790 114.335 ;
        RECT 38.640 114.150 40.790 114.290 ;
        RECT 38.640 114.105 38.930 114.150 ;
        RECT 40.500 114.105 40.790 114.150 ;
        RECT 61.665 114.290 61.955 114.335 ;
        RECT 64.820 114.290 65.110 114.335 ;
        RECT 68.080 114.290 68.370 114.335 ;
        RECT 61.665 114.150 68.370 114.290 ;
        RECT 61.665 114.105 61.955 114.150 ;
        RECT 64.820 114.105 65.110 114.150 ;
        RECT 68.080 114.105 68.370 114.150 ;
        RECT 69.000 114.290 69.290 114.335 ;
        RECT 70.860 114.290 71.150 114.335 ;
        RECT 69.000 114.150 71.150 114.290 ;
        RECT 69.000 114.105 69.290 114.150 ;
        RECT 70.860 114.105 71.150 114.150 ;
        RECT 87.870 114.290 88.190 114.350 ;
        RECT 94.300 114.335 94.515 114.490 ;
        RECT 95.230 114.430 95.550 114.690 ;
        RECT 108.540 114.630 108.830 114.675 ;
        RECT 108.540 114.490 111.075 114.630 ;
        RECT 108.540 114.445 108.830 114.490 ;
        RECT 90.120 114.290 90.410 114.335 ;
        RECT 93.380 114.290 93.670 114.335 ;
        RECT 87.870 114.150 93.670 114.290 ;
        RECT 87.870 114.090 88.190 114.150 ;
        RECT 90.120 114.105 90.410 114.150 ;
        RECT 93.380 114.105 93.670 114.150 ;
        RECT 94.300 114.290 94.590 114.335 ;
        RECT 96.160 114.290 96.450 114.335 ;
        RECT 94.300 114.150 96.450 114.290 ;
        RECT 94.300 114.105 94.590 114.150 ;
        RECT 96.160 114.105 96.450 114.150 ;
        RECT 103.970 114.290 104.290 114.350 ;
        RECT 110.860 114.335 111.075 114.490 ;
        RECT 111.790 114.430 112.110 114.690 ;
        RECT 106.680 114.290 106.970 114.335 ;
        RECT 109.940 114.290 110.230 114.335 ;
        RECT 103.970 114.150 110.230 114.290 ;
        RECT 103.970 114.090 104.290 114.150 ;
        RECT 106.680 114.105 106.970 114.150 ;
        RECT 109.940 114.105 110.230 114.150 ;
        RECT 110.860 114.290 111.150 114.335 ;
        RECT 112.720 114.290 113.010 114.335 ;
        RECT 110.860 114.150 113.010 114.290 ;
        RECT 110.860 114.105 111.150 114.150 ;
        RECT 112.720 114.105 113.010 114.150 ;
        RECT 14.660 113.130 127.820 113.610 ;
        RECT 37.730 112.930 38.050 112.990 ;
        RECT 43.265 112.930 43.555 112.975 ;
        RECT 37.730 112.790 43.555 112.930 ;
        RECT 37.730 112.730 38.050 112.790 ;
        RECT 43.265 112.745 43.555 112.790 ;
        RECT 66.250 112.730 66.570 112.990 ;
        RECT 68.565 112.930 68.855 112.975 ;
        RECT 70.405 112.930 70.695 112.975 ;
        RECT 71.770 112.930 72.090 112.990 ;
        RECT 68.565 112.790 69.700 112.930 ;
        RECT 68.565 112.745 68.855 112.790 ;
        RECT 21.285 112.590 21.575 112.635 ;
        RECT 22.090 112.590 22.410 112.650 ;
        RECT 24.525 112.590 25.175 112.635 ;
        RECT 21.285 112.450 25.175 112.590 ;
        RECT 21.285 112.405 21.875 112.450 ;
        RECT 21.585 112.090 21.875 112.405 ;
        RECT 22.090 112.390 22.410 112.450 ;
        RECT 24.525 112.405 25.175 112.450 ;
        RECT 64.870 112.590 65.190 112.650 ;
        RECT 66.725 112.590 67.015 112.635 ;
        RECT 64.870 112.450 67.015 112.590 ;
        RECT 64.870 112.390 65.190 112.450 ;
        RECT 66.725 112.405 67.015 112.450 ;
        RECT 22.665 112.250 22.955 112.295 ;
        RECT 26.245 112.250 26.535 112.295 ;
        RECT 28.080 112.250 28.370 112.295 ;
        RECT 22.665 112.110 28.370 112.250 ;
        RECT 22.665 112.065 22.955 112.110 ;
        RECT 26.245 112.065 26.535 112.110 ;
        RECT 28.080 112.065 28.370 112.110 ;
        RECT 28.545 112.250 28.835 112.295 ;
        RECT 29.910 112.250 30.230 112.310 ;
        RECT 28.545 112.110 30.230 112.250 ;
        RECT 28.545 112.065 28.835 112.110 ;
        RECT 29.910 112.050 30.230 112.110 ;
        RECT 34.510 112.050 34.830 112.310 ;
        RECT 34.970 112.050 35.290 112.310 ;
        RECT 36.825 112.250 37.115 112.295 ;
        RECT 39.570 112.250 39.890 112.310 ;
        RECT 36.825 112.110 39.890 112.250 ;
        RECT 36.825 112.065 37.115 112.110 ;
        RECT 39.570 112.050 39.890 112.110 ;
        RECT 44.170 112.050 44.490 112.310 ;
        RECT 45.090 112.250 45.410 112.310 ;
        RECT 69.560 112.295 69.700 112.790 ;
        RECT 70.405 112.790 72.090 112.930 ;
        RECT 70.405 112.745 70.695 112.790 ;
        RECT 71.770 112.730 72.090 112.790 ;
        RECT 79.130 112.930 79.450 112.990 ;
        RECT 90.645 112.930 90.935 112.975 ;
        RECT 79.130 112.790 90.935 112.930 ;
        RECT 79.130 112.730 79.450 112.790 ;
        RECT 90.645 112.745 90.935 112.790 ;
        RECT 92.945 112.930 93.235 112.975 ;
        RECT 94.325 112.930 94.615 112.975 ;
        RECT 95.230 112.930 95.550 112.990 ;
        RECT 92.945 112.790 93.620 112.930 ;
        RECT 92.945 112.745 93.235 112.790 ;
        RECT 84.650 112.590 84.970 112.650 ;
        RECT 91.105 112.590 91.395 112.635 ;
        RECT 84.650 112.450 91.395 112.590 ;
        RECT 84.650 112.390 84.970 112.450 ;
        RECT 91.105 112.405 91.395 112.450 ;
        RECT 45.565 112.250 45.855 112.295 ;
        RECT 45.090 112.110 45.855 112.250 ;
        RECT 45.090 112.050 45.410 112.110 ;
        RECT 45.565 112.065 45.855 112.110 ;
        RECT 69.485 112.065 69.775 112.295 ;
        RECT 80.510 112.050 80.830 112.310 ;
        RECT 93.480 112.295 93.620 112.790 ;
        RECT 94.325 112.790 95.550 112.930 ;
        RECT 94.325 112.745 94.615 112.790 ;
        RECT 95.230 112.730 95.550 112.790 ;
        RECT 110.425 112.930 110.715 112.975 ;
        RECT 111.790 112.930 112.110 112.990 ;
        RECT 110.425 112.790 112.110 112.930 ;
        RECT 110.425 112.745 110.715 112.790 ;
        RECT 111.790 112.730 112.110 112.790 ;
        RECT 121.925 112.745 122.215 112.975 ;
        RECT 117.310 112.590 117.630 112.650 ;
        RECT 122.000 112.590 122.140 112.745 ;
        RECT 117.310 112.450 122.140 112.590 ;
        RECT 117.310 112.390 117.630 112.450 ;
        RECT 93.405 112.065 93.695 112.295 ;
        RECT 109.490 112.050 109.810 112.310 ;
        RECT 118.690 112.250 119.010 112.310 ;
        RECT 119.165 112.250 119.455 112.295 ;
        RECT 118.690 112.110 119.455 112.250 ;
        RECT 118.690 112.050 119.010 112.110 ;
        RECT 119.165 112.065 119.455 112.110 ;
        RECT 120.070 112.250 120.390 112.310 ;
        RECT 120.545 112.250 120.835 112.295 ;
        RECT 120.070 112.110 120.835 112.250 ;
        RECT 120.070 112.050 120.390 112.110 ;
        RECT 120.545 112.065 120.835 112.110 ;
        RECT 120.990 112.250 121.310 112.310 ;
        RECT 122.845 112.250 123.135 112.295 ;
        RECT 120.990 112.110 123.135 112.250 ;
        RECT 120.990 112.050 121.310 112.110 ;
        RECT 122.845 112.065 123.135 112.110 ;
        RECT 18.425 111.910 18.715 111.955 ;
        RECT 20.250 111.910 20.570 111.970 ;
        RECT 18.425 111.770 20.570 111.910 ;
        RECT 30.000 111.910 30.140 112.050 ;
        RECT 35.890 111.910 36.210 111.970 ;
        RECT 30.000 111.770 36.210 111.910 ;
        RECT 18.425 111.725 18.715 111.770 ;
        RECT 20.250 111.710 20.570 111.770 ;
        RECT 35.890 111.710 36.210 111.770 ;
        RECT 64.410 111.910 64.730 111.970 ;
        RECT 65.345 111.910 65.635 111.955 ;
        RECT 64.410 111.770 65.635 111.910 ;
        RECT 64.410 111.710 64.730 111.770 ;
        RECT 65.345 111.725 65.635 111.770 ;
        RECT 80.050 111.710 80.370 111.970 ;
        RECT 90.170 111.710 90.490 111.970 ;
        RECT 119.610 111.710 119.930 111.970 ;
        RECT 22.665 111.570 22.955 111.615 ;
        RECT 25.785 111.570 26.075 111.615 ;
        RECT 27.675 111.570 27.965 111.615 ;
        RECT 22.665 111.430 27.965 111.570 ;
        RECT 22.665 111.385 22.955 111.430 ;
        RECT 25.785 111.385 26.075 111.430 ;
        RECT 27.675 111.385 27.965 111.430 ;
        RECT 27.150 111.275 27.470 111.290 ;
        RECT 27.150 111.045 27.520 111.275 ;
        RECT 34.050 111.230 34.370 111.290 ;
        RECT 35.905 111.230 36.195 111.275 ;
        RECT 34.050 111.090 36.195 111.230 ;
        RECT 27.150 111.030 27.470 111.045 ;
        RECT 34.050 111.030 34.370 111.090 ;
        RECT 35.905 111.045 36.195 111.090 ;
        RECT 46.010 111.230 46.330 111.290 ;
        RECT 46.485 111.230 46.775 111.275 ;
        RECT 46.010 111.090 46.775 111.230 ;
        RECT 46.010 111.030 46.330 111.090 ;
        RECT 46.485 111.045 46.775 111.090 ;
        RECT 60.270 111.230 60.590 111.290 ;
        RECT 73.150 111.230 73.470 111.290 ;
        RECT 77.750 111.230 78.070 111.290 ;
        RECT 60.270 111.090 78.070 111.230 ;
        RECT 60.270 111.030 60.590 111.090 ;
        RECT 73.150 111.030 73.470 111.090 ;
        RECT 77.750 111.030 78.070 111.090 ;
        RECT 121.465 111.230 121.755 111.275 ;
        RECT 124.670 111.230 124.990 111.290 ;
        RECT 121.465 111.090 124.990 111.230 ;
        RECT 121.465 111.045 121.755 111.090 ;
        RECT 124.670 111.030 124.990 111.090 ;
        RECT 14.660 110.410 127.820 110.890 ;
        RECT 42.790 110.210 43.110 110.270 ;
        RECT 76.370 110.210 76.690 110.270 ;
        RECT 77.305 110.210 77.595 110.255 ;
        RECT 42.790 110.070 47.160 110.210 ;
        RECT 42.790 110.010 43.110 110.070 ;
        RECT 29.105 109.870 29.395 109.915 ;
        RECT 32.225 109.870 32.515 109.915 ;
        RECT 34.115 109.870 34.405 109.915 ;
        RECT 29.105 109.730 34.405 109.870 ;
        RECT 29.105 109.685 29.395 109.730 ;
        RECT 32.225 109.685 32.515 109.730 ;
        RECT 34.115 109.685 34.405 109.730 ;
        RECT 40.605 109.870 40.895 109.915 ;
        RECT 43.725 109.870 44.015 109.915 ;
        RECT 45.615 109.870 45.905 109.915 ;
        RECT 40.605 109.730 45.905 109.870 ;
        RECT 40.605 109.685 40.895 109.730 ;
        RECT 43.725 109.685 44.015 109.730 ;
        RECT 45.615 109.685 45.905 109.730 ;
        RECT 14.270 109.530 14.590 109.590 ;
        RECT 24.865 109.530 25.155 109.575 ;
        RECT 14.270 109.390 25.155 109.530 ;
        RECT 14.270 109.330 14.590 109.390 ;
        RECT 24.865 109.345 25.155 109.390 ;
        RECT 46.470 109.330 46.790 109.590 ;
        RECT 47.020 109.530 47.160 110.070 ;
        RECT 76.370 110.070 77.595 110.210 ;
        RECT 76.370 110.010 76.690 110.070 ;
        RECT 77.305 110.025 77.595 110.070 ;
        RECT 98.910 110.210 99.230 110.270 ;
        RECT 124.210 110.210 124.530 110.270 ;
        RECT 98.910 110.070 101.440 110.210 ;
        RECT 98.910 110.010 99.230 110.070 ;
        RECT 54.290 109.870 54.610 109.930 ;
        RECT 95.345 109.870 95.635 109.915 ;
        RECT 98.465 109.870 98.755 109.915 ;
        RECT 100.355 109.870 100.645 109.915 ;
        RECT 54.290 109.730 68.320 109.870 ;
        RECT 54.290 109.670 54.610 109.730 ;
        RECT 47.020 109.390 60.960 109.530 ;
        RECT 23.025 109.190 23.315 109.235 ;
        RECT 23.470 109.190 23.790 109.250 ;
        RECT 23.025 109.050 23.790 109.190 ;
        RECT 23.025 109.005 23.315 109.050 ;
        RECT 23.470 108.990 23.790 109.050 ;
        RECT 20.710 108.850 21.030 108.910 ;
        RECT 28.025 108.895 28.315 109.210 ;
        RECT 29.105 109.190 29.395 109.235 ;
        RECT 32.685 109.190 32.975 109.235 ;
        RECT 34.520 109.190 34.810 109.235 ;
        RECT 29.105 109.050 34.810 109.190 ;
        RECT 29.105 109.005 29.395 109.050 ;
        RECT 32.685 109.005 32.975 109.050 ;
        RECT 34.520 109.005 34.810 109.050 ;
        RECT 34.985 109.190 35.275 109.235 ;
        RECT 35.890 109.190 36.210 109.250 ;
        RECT 34.985 109.050 36.210 109.190 ;
        RECT 34.985 109.005 35.275 109.050 ;
        RECT 35.890 108.990 36.210 109.050 ;
        RECT 36.365 109.190 36.655 109.235 ;
        RECT 38.190 109.190 38.510 109.250 ;
        RECT 36.365 109.050 38.510 109.190 ;
        RECT 36.365 109.005 36.655 109.050 ;
        RECT 38.190 108.990 38.510 109.050 ;
        RECT 27.725 108.850 28.315 108.895 ;
        RECT 30.965 108.850 31.615 108.895 ;
        RECT 20.710 108.710 31.615 108.850 ;
        RECT 20.710 108.650 21.030 108.710 ;
        RECT 27.725 108.665 28.015 108.710 ;
        RECT 30.965 108.665 31.615 108.710 ;
        RECT 33.605 108.665 33.895 108.895 ;
        RECT 35.430 108.850 35.750 108.910 ;
        RECT 39.525 108.895 39.815 109.210 ;
        RECT 40.605 109.190 40.895 109.235 ;
        RECT 44.185 109.190 44.475 109.235 ;
        RECT 46.020 109.190 46.310 109.235 ;
        RECT 40.605 109.050 46.310 109.190 ;
        RECT 40.605 109.005 40.895 109.050 ;
        RECT 44.185 109.005 44.475 109.050 ;
        RECT 46.020 109.005 46.310 109.050 ;
        RECT 47.865 109.190 48.155 109.235 ;
        RECT 49.230 109.190 49.550 109.250 ;
        RECT 47.865 109.050 49.550 109.190 ;
        RECT 47.865 109.005 48.155 109.050 ;
        RECT 49.230 108.990 49.550 109.050 ;
        RECT 50.150 109.190 50.470 109.250 ;
        RECT 55.225 109.190 55.515 109.235 ;
        RECT 50.150 109.050 55.515 109.190 ;
        RECT 50.150 108.990 50.470 109.050 ;
        RECT 55.225 109.005 55.515 109.050 ;
        RECT 60.270 108.990 60.590 109.250 ;
        RECT 60.820 109.190 60.960 109.390 ;
        RECT 68.180 109.235 68.320 109.730 ;
        RECT 95.345 109.730 100.645 109.870 ;
        RECT 95.345 109.685 95.635 109.730 ;
        RECT 98.465 109.685 98.755 109.730 ;
        RECT 100.355 109.685 100.645 109.730 ;
        RECT 75.910 109.530 76.230 109.590 ;
        RECT 84.190 109.530 84.510 109.590 ;
        RECT 91.105 109.530 91.395 109.575 ;
        RECT 97.990 109.530 98.310 109.590 ;
        RECT 101.300 109.575 101.440 110.070 ;
        RECT 116.480 110.070 124.530 110.210 ;
        RECT 104.890 109.870 105.210 109.930 ;
        RECT 109.505 109.870 109.795 109.915 ;
        RECT 104.890 109.730 109.795 109.870 ;
        RECT 104.890 109.670 105.210 109.730 ;
        RECT 109.505 109.685 109.795 109.730 ;
        RECT 75.910 109.390 82.580 109.530 ;
        RECT 75.910 109.330 76.230 109.390 ;
        RECT 63.505 109.190 63.795 109.235 ;
        RECT 60.820 109.050 63.795 109.190 ;
        RECT 63.505 109.005 63.795 109.050 ;
        RECT 68.105 109.005 68.395 109.235 ;
        RECT 75.465 109.005 75.755 109.235 ;
        RECT 76.370 109.190 76.690 109.250 ;
        RECT 77.765 109.190 78.055 109.235 ;
        RECT 76.370 109.050 78.055 109.190 ;
        RECT 39.225 108.850 39.815 108.895 ;
        RECT 42.465 108.850 43.115 108.895 ;
        RECT 35.430 108.710 43.115 108.850 ;
        RECT 23.945 108.510 24.235 108.555 ;
        RECT 33.680 108.510 33.820 108.665 ;
        RECT 35.430 108.650 35.750 108.710 ;
        RECT 39.225 108.665 39.515 108.710 ;
        RECT 42.465 108.665 43.115 108.710 ;
        RECT 45.105 108.850 45.395 108.895 ;
        RECT 59.810 108.850 60.130 108.910 ;
        RECT 61.665 108.850 61.955 108.895 ;
        RECT 45.105 108.710 47.160 108.850 ;
        RECT 45.105 108.665 45.395 108.710 ;
        RECT 47.020 108.555 47.160 108.710 ;
        RECT 59.810 108.710 61.955 108.850 ;
        RECT 75.540 108.850 75.680 109.005 ;
        RECT 76.370 108.990 76.690 109.050 ;
        RECT 77.765 109.005 78.055 109.050 ;
        RECT 78.210 108.990 78.530 109.250 ;
        RECT 79.605 109.005 79.895 109.235 ;
        RECT 79.680 108.850 79.820 109.005 ;
        RECT 80.970 108.990 81.290 109.250 ;
        RECT 82.440 109.235 82.580 109.390 ;
        RECT 84.190 109.390 89.940 109.530 ;
        RECT 84.190 109.330 84.510 109.390 ;
        RECT 89.800 109.235 89.940 109.390 ;
        RECT 91.105 109.390 98.310 109.530 ;
        RECT 91.105 109.345 91.395 109.390 ;
        RECT 97.990 109.330 98.310 109.390 ;
        RECT 101.225 109.345 101.515 109.575 ;
        RECT 115.945 109.530 116.235 109.575 ;
        RECT 116.480 109.530 116.620 110.070 ;
        RECT 124.210 110.010 124.530 110.070 ;
        RECT 116.815 109.870 117.105 109.915 ;
        RECT 118.705 109.870 118.995 109.915 ;
        RECT 121.825 109.870 122.115 109.915 ;
        RECT 116.815 109.730 122.115 109.870 ;
        RECT 116.815 109.685 117.105 109.730 ;
        RECT 118.705 109.685 118.995 109.730 ;
        RECT 121.825 109.685 122.115 109.730 ;
        RECT 115.945 109.390 116.620 109.530 ;
        RECT 115.945 109.345 116.235 109.390 ;
        RECT 117.310 109.330 117.630 109.590 ;
        RECT 82.365 109.005 82.655 109.235 ;
        RECT 88.345 109.005 88.635 109.235 ;
        RECT 89.725 109.005 90.015 109.235 ;
        RECT 80.510 108.850 80.830 108.910 ;
        RECT 84.190 108.850 84.510 108.910 ;
        RECT 88.420 108.850 88.560 109.005 ;
        RECT 94.265 108.895 94.555 109.210 ;
        RECT 95.345 109.190 95.635 109.235 ;
        RECT 98.925 109.190 99.215 109.235 ;
        RECT 100.760 109.190 101.050 109.235 ;
        RECT 95.345 109.050 101.050 109.190 ;
        RECT 95.345 109.005 95.635 109.050 ;
        RECT 98.925 109.005 99.215 109.050 ;
        RECT 100.760 109.005 101.050 109.050 ;
        RECT 103.050 108.990 103.370 109.250 ;
        RECT 105.365 109.005 105.655 109.235 ;
        RECT 106.270 109.190 106.590 109.250 ;
        RECT 106.745 109.190 107.035 109.235 ;
        RECT 106.270 109.050 107.035 109.190 ;
        RECT 97.530 108.895 97.850 108.910 ;
        RECT 93.965 108.850 94.555 108.895 ;
        RECT 97.205 108.850 97.855 108.895 ;
        RECT 75.540 108.710 91.320 108.850 ;
        RECT 59.810 108.650 60.130 108.710 ;
        RECT 61.665 108.665 61.955 108.710 ;
        RECT 80.510 108.650 80.830 108.710 ;
        RECT 84.190 108.650 84.510 108.710 ;
        RECT 23.945 108.370 33.820 108.510 ;
        RECT 23.945 108.325 24.235 108.370 ;
        RECT 46.945 108.325 47.235 108.555 ;
        RECT 56.145 108.510 56.435 108.555 ;
        RECT 60.270 108.510 60.590 108.570 ;
        RECT 56.145 108.370 60.590 108.510 ;
        RECT 56.145 108.325 56.435 108.370 ;
        RECT 60.270 108.310 60.590 108.370 ;
        RECT 64.425 108.510 64.715 108.555 ;
        RECT 67.170 108.510 67.490 108.570 ;
        RECT 64.425 108.370 67.490 108.510 ;
        RECT 64.425 108.325 64.715 108.370 ;
        RECT 67.170 108.310 67.490 108.370 ;
        RECT 69.025 108.510 69.315 108.555 ;
        RECT 72.230 108.510 72.550 108.570 ;
        RECT 69.025 108.370 72.550 108.510 ;
        RECT 69.025 108.325 69.315 108.370 ;
        RECT 72.230 108.310 72.550 108.370 ;
        RECT 75.005 108.510 75.295 108.555 ;
        RECT 79.590 108.510 79.910 108.570 ;
        RECT 75.005 108.370 79.910 108.510 ;
        RECT 75.005 108.325 75.295 108.370 ;
        RECT 79.590 108.310 79.910 108.370 ;
        RECT 81.890 108.310 82.210 108.570 ;
        RECT 83.270 108.310 83.590 108.570 ;
        RECT 88.790 108.310 89.110 108.570 ;
        RECT 90.630 108.310 90.950 108.570 ;
        RECT 91.180 108.510 91.320 108.710 ;
        RECT 93.965 108.710 97.855 108.850 ;
        RECT 93.965 108.665 94.255 108.710 ;
        RECT 97.205 108.665 97.855 108.710 ;
        RECT 99.845 108.665 100.135 108.895 ;
        RECT 100.290 108.850 100.610 108.910 ;
        RECT 105.440 108.850 105.580 109.005 ;
        RECT 106.270 108.990 106.590 109.050 ;
        RECT 106.745 109.005 107.035 109.050 ;
        RECT 110.425 109.190 110.715 109.235 ;
        RECT 111.330 109.190 111.650 109.250 ;
        RECT 110.425 109.050 111.650 109.190 ;
        RECT 110.425 109.005 110.715 109.050 ;
        RECT 111.330 108.990 111.650 109.050 ;
        RECT 114.550 108.990 114.870 109.250 ;
        RECT 116.410 109.190 116.700 109.235 ;
        RECT 118.245 109.190 118.535 109.235 ;
        RECT 121.825 109.190 122.115 109.235 ;
        RECT 116.410 109.050 122.115 109.190 ;
        RECT 116.410 109.005 116.700 109.050 ;
        RECT 118.245 109.005 118.535 109.050 ;
        RECT 121.825 109.005 122.115 109.050 ;
        RECT 112.710 108.850 113.030 108.910 ;
        RECT 119.610 108.895 119.930 108.910 ;
        RECT 122.905 108.895 123.195 109.210 ;
        RECT 100.290 108.710 113.030 108.850 ;
        RECT 97.530 108.650 97.850 108.665 ;
        RECT 99.370 108.510 99.690 108.570 ;
        RECT 91.180 108.370 99.690 108.510 ;
        RECT 99.920 108.510 100.060 108.665 ;
        RECT 100.290 108.650 100.610 108.710 ;
        RECT 112.710 108.650 113.030 108.710 ;
        RECT 119.605 108.850 120.255 108.895 ;
        RECT 122.905 108.850 123.495 108.895 ;
        RECT 119.605 108.710 123.495 108.850 ;
        RECT 119.605 108.665 120.255 108.710 ;
        RECT 123.205 108.665 123.495 108.710 ;
        RECT 126.065 108.850 126.355 108.895 ;
        RECT 127.890 108.850 128.210 108.910 ;
        RECT 126.065 108.710 128.210 108.850 ;
        RECT 126.065 108.665 126.355 108.710 ;
        RECT 119.610 108.650 119.930 108.665 ;
        RECT 127.890 108.650 128.210 108.710 ;
        RECT 102.145 108.510 102.435 108.555 ;
        RECT 99.920 108.370 102.435 108.510 ;
        RECT 99.370 108.310 99.690 108.370 ;
        RECT 102.145 108.325 102.435 108.370 ;
        RECT 104.905 108.510 105.195 108.555 ;
        RECT 105.350 108.510 105.670 108.570 ;
        RECT 104.905 108.370 105.670 108.510 ;
        RECT 104.905 108.325 105.195 108.370 ;
        RECT 105.350 108.310 105.670 108.370 ;
        RECT 107.665 108.510 107.955 108.555 ;
        RECT 109.030 108.510 109.350 108.570 ;
        RECT 107.665 108.370 109.350 108.510 ;
        RECT 107.665 108.325 107.955 108.370 ;
        RECT 109.030 108.310 109.350 108.370 ;
        RECT 115.470 108.310 115.790 108.570 ;
        RECT 14.660 107.690 127.820 108.170 ;
        RECT 20.710 107.290 21.030 107.550 ;
        RECT 22.090 107.490 22.410 107.550 ;
        RECT 23.025 107.490 23.315 107.535 ;
        RECT 22.090 107.350 23.315 107.490 ;
        RECT 22.090 107.290 22.410 107.350 ;
        RECT 23.025 107.305 23.315 107.350 ;
        RECT 34.985 107.490 35.275 107.535 ;
        RECT 35.430 107.490 35.750 107.550 ;
        RECT 45.550 107.490 45.870 107.550 ;
        RECT 34.985 107.350 35.750 107.490 ;
        RECT 34.985 107.305 35.275 107.350 ;
        RECT 35.430 107.290 35.750 107.350 ;
        RECT 35.980 107.350 45.870 107.490 ;
        RECT 26.805 107.150 27.095 107.195 ;
        RECT 30.045 107.150 30.695 107.195 ;
        RECT 26.805 107.010 30.695 107.150 ;
        RECT 26.805 106.965 27.395 107.010 ;
        RECT 30.045 106.965 30.695 107.010 ;
        RECT 32.685 107.150 32.975 107.195 ;
        RECT 34.050 107.150 34.370 107.210 ;
        RECT 32.685 107.010 34.370 107.150 ;
        RECT 32.685 106.965 32.975 107.010 ;
        RECT 21.185 106.810 21.475 106.855 ;
        RECT 23.485 106.810 23.775 106.855 ;
        RECT 27.105 106.810 27.395 106.965 ;
        RECT 34.050 106.950 34.370 107.010 ;
        RECT 21.185 106.670 23.775 106.810 ;
        RECT 21.185 106.625 21.475 106.670 ;
        RECT 23.485 106.625 23.775 106.670 ;
        RECT 26.780 106.670 27.395 106.810 ;
        RECT 23.560 106.130 23.700 106.625 ;
        RECT 26.780 106.530 26.920 106.670 ;
        RECT 27.105 106.650 27.395 106.670 ;
        RECT 28.185 106.810 28.475 106.855 ;
        RECT 31.765 106.810 32.055 106.855 ;
        RECT 33.600 106.810 33.890 106.855 ;
        RECT 28.185 106.670 33.890 106.810 ;
        RECT 28.185 106.625 28.475 106.670 ;
        RECT 31.765 106.625 32.055 106.670 ;
        RECT 33.600 106.625 33.890 106.670 ;
        RECT 34.525 106.810 34.815 106.855 ;
        RECT 34.970 106.810 35.290 106.870 ;
        RECT 35.980 106.855 36.120 107.350 ;
        RECT 45.550 107.290 45.870 107.350 ;
        RECT 46.010 107.290 46.330 107.550 ;
        RECT 68.090 107.490 68.410 107.550 ;
        RECT 64.500 107.350 68.410 107.490 ;
        RECT 41.065 107.150 41.355 107.195 ;
        RECT 44.305 107.150 44.955 107.195 ;
        RECT 41.065 107.010 44.955 107.150 ;
        RECT 46.100 107.150 46.240 107.290 ;
        RECT 46.910 107.150 47.200 107.195 ;
        RECT 46.100 107.010 47.200 107.150 ;
        RECT 41.065 106.965 41.655 107.010 ;
        RECT 44.305 106.965 44.955 107.010 ;
        RECT 46.910 106.965 47.200 107.010 ;
        RECT 54.405 107.150 54.695 107.195 ;
        RECT 56.590 107.150 56.910 107.210 ;
        RECT 57.645 107.150 58.295 107.195 ;
        RECT 54.405 107.010 58.295 107.150 ;
        RECT 54.405 106.965 54.995 107.010 ;
        RECT 35.905 106.810 36.195 106.855 ;
        RECT 34.525 106.670 36.195 106.810 ;
        RECT 34.525 106.625 34.815 106.670 ;
        RECT 34.970 106.610 35.290 106.670 ;
        RECT 35.905 106.625 36.195 106.670 ;
        RECT 36.365 106.810 36.655 106.855 ;
        RECT 41.365 106.810 41.655 106.965 ;
        RECT 36.365 106.670 41.655 106.810 ;
        RECT 36.365 106.625 36.655 106.670 ;
        RECT 41.365 106.650 41.655 106.670 ;
        RECT 42.445 106.810 42.735 106.855 ;
        RECT 46.025 106.810 46.315 106.855 ;
        RECT 47.860 106.810 48.150 106.855 ;
        RECT 42.445 106.670 48.150 106.810 ;
        RECT 42.445 106.625 42.735 106.670 ;
        RECT 46.025 106.625 46.315 106.670 ;
        RECT 47.860 106.625 48.150 106.670 ;
        RECT 49.690 106.610 50.010 106.870 ;
        RECT 51.085 106.810 51.375 106.855 ;
        RECT 51.990 106.810 52.310 106.870 ;
        RECT 51.085 106.670 52.310 106.810 ;
        RECT 51.085 106.625 51.375 106.670 ;
        RECT 51.990 106.610 52.310 106.670 ;
        RECT 54.705 106.650 54.995 106.965 ;
        RECT 56.590 106.950 56.910 107.010 ;
        RECT 57.645 106.965 58.295 107.010 ;
        RECT 60.270 106.950 60.590 107.210 ;
        RECT 63.505 107.150 63.795 107.195 ;
        RECT 64.500 107.150 64.640 107.350 ;
        RECT 68.090 107.290 68.410 107.350 ;
        RECT 82.350 107.490 82.670 107.550 ;
        RECT 88.790 107.490 89.110 107.550 ;
        RECT 120.530 107.490 120.850 107.550 ;
        RECT 82.350 107.350 87.180 107.490 ;
        RECT 82.350 107.290 82.670 107.350 ;
        RECT 63.505 107.010 64.640 107.150 ;
        RECT 64.870 107.150 65.190 107.210 ;
        RECT 66.365 107.150 66.655 107.195 ;
        RECT 69.605 107.150 70.255 107.195 ;
        RECT 64.870 107.010 70.255 107.150 ;
        RECT 63.505 106.965 63.795 107.010 ;
        RECT 64.870 106.950 65.190 107.010 ;
        RECT 66.365 106.965 66.955 107.010 ;
        RECT 69.605 106.965 70.255 107.010 ;
        RECT 55.785 106.810 56.075 106.855 ;
        RECT 59.365 106.810 59.655 106.855 ;
        RECT 61.200 106.810 61.490 106.855 ;
        RECT 55.785 106.670 61.490 106.810 ;
        RECT 55.785 106.625 56.075 106.670 ;
        RECT 59.365 106.625 59.655 106.670 ;
        RECT 61.200 106.625 61.490 106.670 ;
        RECT 66.665 106.650 66.955 106.965 ;
        RECT 72.230 106.950 72.550 107.210 ;
        RECT 77.865 107.150 78.155 107.195 ;
        RECT 80.050 107.150 80.370 107.210 ;
        RECT 81.105 107.150 81.755 107.195 ;
        RECT 77.865 107.010 81.755 107.150 ;
        RECT 77.865 106.965 78.455 107.010 ;
        RECT 67.745 106.810 68.035 106.855 ;
        RECT 71.325 106.810 71.615 106.855 ;
        RECT 73.160 106.810 73.450 106.855 ;
        RECT 67.745 106.670 73.450 106.810 ;
        RECT 67.745 106.625 68.035 106.670 ;
        RECT 71.325 106.625 71.615 106.670 ;
        RECT 73.160 106.625 73.450 106.670 ;
        RECT 73.625 106.810 73.915 106.855 ;
        RECT 74.070 106.810 74.390 106.870 ;
        RECT 73.625 106.670 74.390 106.810 ;
        RECT 73.625 106.625 73.915 106.670 ;
        RECT 74.070 106.610 74.390 106.670 ;
        RECT 78.165 106.650 78.455 106.965 ;
        RECT 80.050 106.950 80.370 107.010 ;
        RECT 81.105 106.965 81.755 107.010 ;
        RECT 83.270 107.150 83.590 107.210 ;
        RECT 83.745 107.150 84.035 107.195 ;
        RECT 83.270 107.010 84.035 107.150 ;
        RECT 83.270 106.950 83.590 107.010 ;
        RECT 83.745 106.965 84.035 107.010 ;
        RECT 84.190 107.150 84.510 107.210 ;
        RECT 84.190 107.010 85.800 107.150 ;
        RECT 84.190 106.950 84.510 107.010 ;
        RECT 85.660 106.855 85.800 107.010 ;
        RECT 87.040 106.855 87.180 107.350 ;
        RECT 88.790 107.350 91.320 107.490 ;
        RECT 88.790 107.290 89.110 107.350 ;
        RECT 90.630 106.950 90.950 107.210 ;
        RECT 91.180 107.150 91.320 107.350 ;
        RECT 116.020 107.350 120.850 107.490 ;
        RECT 92.925 107.150 93.575 107.195 ;
        RECT 96.525 107.150 96.815 107.195 ;
        RECT 91.180 107.010 96.815 107.150 ;
        RECT 92.925 106.965 93.575 107.010 ;
        RECT 96.225 106.965 96.815 107.010 ;
        RECT 103.165 107.150 103.455 107.195 ;
        RECT 105.350 107.150 105.670 107.210 ;
        RECT 106.405 107.150 107.055 107.195 ;
        RECT 103.165 107.010 107.055 107.150 ;
        RECT 103.165 106.965 103.755 107.010 ;
        RECT 79.245 106.810 79.535 106.855 ;
        RECT 82.825 106.810 83.115 106.855 ;
        RECT 84.660 106.810 84.950 106.855 ;
        RECT 79.245 106.670 84.950 106.810 ;
        RECT 79.245 106.625 79.535 106.670 ;
        RECT 82.825 106.625 83.115 106.670 ;
        RECT 84.660 106.625 84.950 106.670 ;
        RECT 85.585 106.625 85.875 106.855 ;
        RECT 86.965 106.625 87.255 106.855 ;
        RECT 89.730 106.810 90.020 106.855 ;
        RECT 91.565 106.810 91.855 106.855 ;
        RECT 95.145 106.810 95.435 106.855 ;
        RECT 89.730 106.670 95.435 106.810 ;
        RECT 89.730 106.625 90.020 106.670 ;
        RECT 91.565 106.625 91.855 106.670 ;
        RECT 95.145 106.625 95.435 106.670 ;
        RECT 96.225 106.650 96.515 106.965 ;
        RECT 103.465 106.650 103.755 106.965 ;
        RECT 105.350 106.950 105.670 107.010 ;
        RECT 106.405 106.965 107.055 107.010 ;
        RECT 109.030 106.950 109.350 107.210 ;
        RECT 116.020 107.195 116.160 107.350 ;
        RECT 120.530 107.290 120.850 107.350 ;
        RECT 115.945 106.965 116.235 107.195 ;
        RECT 118.805 107.150 119.095 107.195 ;
        RECT 122.045 107.150 122.695 107.195 ;
        RECT 118.805 107.010 122.695 107.150 ;
        RECT 118.805 106.965 119.395 107.010 ;
        RECT 122.045 106.965 122.695 107.010 ;
        RECT 119.105 106.870 119.395 106.965 ;
        RECT 124.670 106.950 124.990 107.210 ;
        RECT 104.545 106.810 104.835 106.855 ;
        RECT 108.125 106.810 108.415 106.855 ;
        RECT 109.960 106.810 110.250 106.855 ;
        RECT 104.545 106.670 110.250 106.810 ;
        RECT 104.545 106.625 104.835 106.670 ;
        RECT 108.125 106.625 108.415 106.670 ;
        RECT 109.960 106.625 110.250 106.670 ;
        RECT 111.805 106.810 112.095 106.855 ;
        RECT 112.710 106.810 113.030 106.870 ;
        RECT 113.185 106.810 113.475 106.855 ;
        RECT 118.230 106.810 118.550 106.870 ;
        RECT 111.805 106.670 118.550 106.810 ;
        RECT 111.805 106.625 112.095 106.670 ;
        RECT 112.710 106.610 113.030 106.670 ;
        RECT 113.185 106.625 113.475 106.670 ;
        RECT 118.230 106.610 118.550 106.670 ;
        RECT 119.105 106.650 119.470 106.870 ;
        RECT 119.150 106.610 119.470 106.650 ;
        RECT 120.185 106.810 120.475 106.855 ;
        RECT 123.765 106.810 124.055 106.855 ;
        RECT 125.600 106.810 125.890 106.855 ;
        RECT 120.185 106.670 125.890 106.810 ;
        RECT 135.660 106.690 136.800 133.400 ;
        RECT 120.185 106.625 120.475 106.670 ;
        RECT 123.765 106.625 124.055 106.670 ;
        RECT 125.600 106.625 125.890 106.670 ;
        RECT 133.100 106.600 136.850 106.690 ;
        RECT 23.945 106.470 24.235 106.515 ;
        RECT 26.230 106.470 26.550 106.530 ;
        RECT 23.945 106.330 26.550 106.470 ;
        RECT 23.945 106.285 24.235 106.330 ;
        RECT 26.230 106.270 26.550 106.330 ;
        RECT 26.690 106.270 27.010 106.530 ;
        RECT 34.065 106.470 34.355 106.515 ;
        RECT 38.205 106.470 38.495 106.515 ;
        RECT 44.170 106.470 44.490 106.530 ;
        RECT 34.065 106.330 36.120 106.470 ;
        RECT 34.065 106.285 34.355 106.330 ;
        RECT 35.980 106.190 36.120 106.330 ;
        RECT 38.205 106.330 44.490 106.470 ;
        RECT 38.205 106.285 38.495 106.330 ;
        RECT 44.170 106.270 44.490 106.330 ;
        RECT 46.470 106.470 46.790 106.530 ;
        RECT 48.325 106.470 48.615 106.515 ;
        RECT 46.470 106.330 48.615 106.470 ;
        RECT 46.470 106.270 46.790 106.330 ;
        RECT 48.325 106.285 48.615 106.330 ;
        RECT 51.545 106.470 51.835 106.515 ;
        RECT 54.290 106.470 54.610 106.530 ;
        RECT 51.545 106.330 54.610 106.470 ;
        RECT 51.545 106.285 51.835 106.330 ;
        RECT 54.290 106.270 54.610 106.330 ;
        RECT 61.665 106.470 61.955 106.515 ;
        RECT 63.950 106.470 64.270 106.530 ;
        RECT 61.665 106.330 64.270 106.470 ;
        RECT 61.665 106.285 61.955 106.330 ;
        RECT 63.950 106.270 64.270 106.330 ;
        RECT 75.005 106.470 75.295 106.515 ;
        RECT 80.050 106.470 80.370 106.530 ;
        RECT 75.005 106.330 80.370 106.470 ;
        RECT 75.005 106.285 75.295 106.330 ;
        RECT 80.050 106.270 80.370 106.330 ;
        RECT 85.125 106.470 85.415 106.515 ;
        RECT 89.250 106.470 89.570 106.530 ;
        RECT 85.125 106.330 89.570 106.470 ;
        RECT 85.125 106.285 85.415 106.330 ;
        RECT 89.250 106.270 89.570 106.330 ;
        RECT 93.850 106.470 94.170 106.530 ;
        RECT 99.385 106.470 99.675 106.515 ;
        RECT 93.850 106.330 99.675 106.470 ;
        RECT 93.850 106.270 94.170 106.330 ;
        RECT 99.385 106.285 99.675 106.330 ;
        RECT 100.305 106.470 100.595 106.515 ;
        RECT 103.970 106.470 104.290 106.530 ;
        RECT 100.305 106.330 104.290 106.470 ;
        RECT 100.305 106.285 100.595 106.330 ;
        RECT 103.970 106.270 104.290 106.330 ;
        RECT 110.425 106.470 110.715 106.515 ;
        RECT 124.210 106.470 124.530 106.530 ;
        RECT 126.065 106.470 126.355 106.515 ;
        RECT 110.425 106.330 126.355 106.470 ;
        RECT 110.425 106.285 110.715 106.330 ;
        RECT 124.210 106.270 124.530 106.330 ;
        RECT 126.065 106.285 126.355 106.330 ;
        RECT 28.185 106.130 28.475 106.175 ;
        RECT 31.305 106.130 31.595 106.175 ;
        RECT 33.195 106.130 33.485 106.175 ;
        RECT 23.560 105.990 27.840 106.130 ;
        RECT 27.700 105.850 27.840 105.990 ;
        RECT 28.185 105.990 33.485 106.130 ;
        RECT 28.185 105.945 28.475 105.990 ;
        RECT 31.305 105.945 31.595 105.990 ;
        RECT 33.195 105.945 33.485 105.990 ;
        RECT 35.890 105.930 36.210 106.190 ;
        RECT 42.445 106.130 42.735 106.175 ;
        RECT 45.565 106.130 45.855 106.175 ;
        RECT 47.455 106.130 47.745 106.175 ;
        RECT 50.165 106.130 50.455 106.175 ;
        RECT 42.445 105.990 47.745 106.130 ;
        RECT 42.445 105.945 42.735 105.990 ;
        RECT 45.565 105.945 45.855 105.990 ;
        RECT 47.455 105.945 47.745 105.990 ;
        RECT 47.940 105.990 50.455 106.130 ;
        RECT 27.610 105.790 27.930 105.850 ;
        RECT 34.970 105.790 35.290 105.850 ;
        RECT 27.610 105.650 35.290 105.790 ;
        RECT 27.610 105.590 27.930 105.650 ;
        RECT 34.970 105.590 35.290 105.650 ;
        RECT 40.950 105.790 41.270 105.850 ;
        RECT 47.940 105.790 48.080 105.990 ;
        RECT 50.165 105.945 50.455 105.990 ;
        RECT 55.785 106.130 56.075 106.175 ;
        RECT 58.905 106.130 59.195 106.175 ;
        RECT 60.795 106.130 61.085 106.175 ;
        RECT 55.785 105.990 61.085 106.130 ;
        RECT 55.785 105.945 56.075 105.990 ;
        RECT 58.905 105.945 59.195 105.990 ;
        RECT 60.795 105.945 61.085 105.990 ;
        RECT 67.745 106.130 68.035 106.175 ;
        RECT 70.865 106.130 71.155 106.175 ;
        RECT 72.755 106.130 73.045 106.175 ;
        RECT 67.745 105.990 73.045 106.130 ;
        RECT 67.745 105.945 68.035 105.990 ;
        RECT 70.865 105.945 71.155 105.990 ;
        RECT 72.755 105.945 73.045 105.990 ;
        RECT 79.245 106.130 79.535 106.175 ;
        RECT 82.365 106.130 82.655 106.175 ;
        RECT 84.255 106.130 84.545 106.175 ;
        RECT 79.245 105.990 84.545 106.130 ;
        RECT 79.245 105.945 79.535 105.990 ;
        RECT 82.365 105.945 82.655 105.990 ;
        RECT 84.255 105.945 84.545 105.990 ;
        RECT 90.135 106.130 90.425 106.175 ;
        RECT 92.025 106.130 92.315 106.175 ;
        RECT 95.145 106.130 95.435 106.175 ;
        RECT 90.135 105.990 95.435 106.130 ;
        RECT 90.135 105.945 90.425 105.990 ;
        RECT 92.025 105.945 92.315 105.990 ;
        RECT 95.145 105.945 95.435 105.990 ;
        RECT 104.545 106.130 104.835 106.175 ;
        RECT 107.665 106.130 107.955 106.175 ;
        RECT 109.555 106.130 109.845 106.175 ;
        RECT 104.545 105.990 109.845 106.130 ;
        RECT 104.545 105.945 104.835 105.990 ;
        RECT 107.665 105.945 107.955 105.990 ;
        RECT 109.555 105.945 109.845 105.990 ;
        RECT 120.185 106.130 120.475 106.175 ;
        RECT 123.305 106.130 123.595 106.175 ;
        RECT 125.195 106.130 125.485 106.175 ;
        RECT 120.185 105.990 125.485 106.130 ;
        RECT 120.185 105.945 120.475 105.990 ;
        RECT 123.305 105.945 123.595 105.990 ;
        RECT 125.195 105.945 125.485 105.990 ;
        RECT 40.950 105.650 48.080 105.790 ;
        RECT 40.950 105.590 41.270 105.650 ;
        RECT 49.230 105.590 49.550 105.850 ;
        RECT 86.045 105.790 86.335 105.835 ;
        RECT 87.410 105.790 87.730 105.850 ;
        RECT 86.045 105.650 87.730 105.790 ;
        RECT 86.045 105.605 86.335 105.650 ;
        RECT 87.410 105.590 87.730 105.650 ;
        RECT 87.870 105.590 88.190 105.850 ;
        RECT 111.330 105.590 111.650 105.850 ;
        RECT 113.645 105.790 113.935 105.835 ;
        RECT 116.390 105.790 116.710 105.850 ;
        RECT 113.645 105.650 116.710 105.790 ;
        RECT 113.645 105.605 113.935 105.650 ;
        RECT 116.390 105.590 116.710 105.650 ;
        RECT 129.700 105.630 136.850 106.600 ;
        RECT 133.100 105.500 136.850 105.630 ;
        RECT 14.660 104.970 127.820 105.450 ;
        RECT 26.690 104.570 27.010 104.830 ;
        RECT 27.150 104.770 27.470 104.830 ;
        RECT 27.625 104.770 27.915 104.815 ;
        RECT 27.150 104.630 27.915 104.770 ;
        RECT 27.150 104.570 27.470 104.630 ;
        RECT 27.625 104.585 27.915 104.630 ;
        RECT 35.890 104.770 36.210 104.830 ;
        RECT 46.470 104.770 46.790 104.830 ;
        RECT 35.890 104.630 46.790 104.770 ;
        RECT 35.890 104.570 36.210 104.630 ;
        RECT 33.245 104.430 33.535 104.475 ;
        RECT 36.365 104.430 36.655 104.475 ;
        RECT 38.255 104.430 38.545 104.475 ;
        RECT 33.245 104.290 38.545 104.430 ;
        RECT 33.245 104.245 33.535 104.290 ;
        RECT 36.365 104.245 36.655 104.290 ;
        RECT 38.255 104.245 38.545 104.290 ;
        RECT 37.730 103.890 38.050 104.150 ;
        RECT 39.125 104.090 39.415 104.135 ;
        RECT 39.585 104.090 39.875 104.135 ;
        RECT 40.120 104.090 40.260 104.630 ;
        RECT 46.470 104.570 46.790 104.630 ;
        RECT 56.145 104.770 56.435 104.815 ;
        RECT 56.590 104.770 56.910 104.830 ;
        RECT 56.145 104.630 56.910 104.770 ;
        RECT 56.145 104.585 56.435 104.630 ;
        RECT 56.590 104.570 56.910 104.630 ;
        RECT 64.410 104.770 64.730 104.830 ;
        RECT 89.250 104.770 89.570 104.830 ;
        RECT 97.530 104.770 97.850 104.830 ;
        RECT 98.925 104.770 99.215 104.815 ;
        RECT 64.410 104.630 68.320 104.770 ;
        RECT 64.410 104.570 64.730 104.630 ;
        RECT 40.455 104.430 40.745 104.475 ;
        RECT 42.345 104.430 42.635 104.475 ;
        RECT 45.465 104.430 45.755 104.475 ;
        RECT 40.455 104.290 45.755 104.430 ;
        RECT 40.455 104.245 40.745 104.290 ;
        RECT 42.345 104.245 42.635 104.290 ;
        RECT 45.465 104.245 45.755 104.290 ;
        RECT 62.685 104.430 62.975 104.475 ;
        RECT 65.805 104.430 66.095 104.475 ;
        RECT 67.695 104.430 67.985 104.475 ;
        RECT 62.685 104.290 67.985 104.430 ;
        RECT 62.685 104.245 62.975 104.290 ;
        RECT 65.805 104.245 66.095 104.290 ;
        RECT 67.695 104.245 67.985 104.290 ;
        RECT 39.125 103.950 40.260 104.090 ;
        RECT 39.125 103.905 39.415 103.950 ;
        RECT 39.585 103.905 39.875 103.950 ;
        RECT 40.950 103.890 41.270 104.150 ;
        RECT 49.690 103.890 50.010 104.150 ;
        RECT 67.170 103.890 67.490 104.150 ;
        RECT 68.180 104.090 68.320 104.630 ;
        RECT 89.250 104.630 97.300 104.770 ;
        RECT 89.250 104.570 89.570 104.630 ;
        RECT 80.625 104.430 80.915 104.475 ;
        RECT 83.745 104.430 84.035 104.475 ;
        RECT 85.635 104.430 85.925 104.475 ;
        RECT 89.340 104.430 89.480 104.570 ;
        RECT 80.625 104.290 85.925 104.430 ;
        RECT 80.625 104.245 80.915 104.290 ;
        RECT 83.745 104.245 84.035 104.290 ;
        RECT 85.635 104.245 85.925 104.290 ;
        RECT 86.580 104.290 89.480 104.430 ;
        RECT 91.205 104.430 91.495 104.475 ;
        RECT 94.325 104.430 94.615 104.475 ;
        RECT 96.215 104.430 96.505 104.475 ;
        RECT 91.205 104.290 96.505 104.430 ;
        RECT 68.565 104.090 68.855 104.135 ;
        RECT 74.070 104.090 74.390 104.150 ;
        RECT 68.180 103.950 74.390 104.090 ;
        RECT 68.565 103.905 68.855 103.950 ;
        RECT 74.070 103.890 74.390 103.950 ;
        RECT 81.890 104.090 82.210 104.150 ;
        RECT 86.580 104.135 86.720 104.290 ;
        RECT 91.205 104.245 91.495 104.290 ;
        RECT 94.325 104.245 94.615 104.290 ;
        RECT 96.215 104.245 96.505 104.290 ;
        RECT 85.125 104.090 85.415 104.135 ;
        RECT 81.890 103.950 85.415 104.090 ;
        RECT 81.890 103.890 82.210 103.950 ;
        RECT 85.125 103.905 85.415 103.950 ;
        RECT 86.505 103.905 86.795 104.135 ;
        RECT 87.870 104.090 88.190 104.150 ;
        RECT 97.160 104.135 97.300 104.630 ;
        RECT 97.530 104.630 99.215 104.770 ;
        RECT 97.530 104.570 97.850 104.630 ;
        RECT 98.925 104.585 99.215 104.630 ;
        RECT 104.395 104.430 104.685 104.475 ;
        RECT 106.285 104.430 106.575 104.475 ;
        RECT 109.405 104.430 109.695 104.475 ;
        RECT 104.395 104.290 109.695 104.430 ;
        RECT 104.395 104.245 104.685 104.290 ;
        RECT 106.285 104.245 106.575 104.290 ;
        RECT 109.405 104.245 109.695 104.290 ;
        RECT 118.345 104.430 118.635 104.475 ;
        RECT 121.465 104.430 121.755 104.475 ;
        RECT 123.355 104.430 123.645 104.475 ;
        RECT 118.345 104.290 123.645 104.430 ;
        RECT 118.345 104.245 118.635 104.290 ;
        RECT 121.465 104.245 121.755 104.290 ;
        RECT 123.355 104.245 123.645 104.290 ;
        RECT 95.705 104.090 95.995 104.135 ;
        RECT 87.870 103.950 95.995 104.090 ;
        RECT 87.870 103.890 88.190 103.950 ;
        RECT 95.705 103.905 95.995 103.950 ;
        RECT 97.085 104.090 97.375 104.135 ;
        RECT 98.910 104.090 99.230 104.150 ;
        RECT 103.525 104.090 103.815 104.135 ;
        RECT 97.085 103.950 103.815 104.090 ;
        RECT 97.085 103.905 97.375 103.950 ;
        RECT 98.910 103.890 99.230 103.950 ;
        RECT 103.525 103.905 103.815 103.950 ;
        RECT 104.890 103.890 105.210 104.150 ;
        RECT 109.950 104.090 110.270 104.150 ;
        RECT 113.645 104.090 113.935 104.135 ;
        RECT 109.950 103.950 113.935 104.090 ;
        RECT 109.950 103.890 110.270 103.950 ;
        RECT 113.645 103.905 113.935 103.950 ;
        RECT 115.470 104.090 115.790 104.150 ;
        RECT 122.845 104.090 123.135 104.135 ;
        RECT 115.470 103.950 123.135 104.090 ;
        RECT 115.470 103.890 115.790 103.950 ;
        RECT 122.845 103.905 123.135 103.950 ;
        RECT 124.210 103.890 124.530 104.150 ;
        RECT 26.245 103.750 26.535 103.795 ;
        RECT 27.610 103.750 27.930 103.810 ;
        RECT 26.245 103.610 27.930 103.750 ;
        RECT 26.245 103.565 26.535 103.610 ;
        RECT 27.610 103.550 27.930 103.610 ;
        RECT 28.530 103.550 28.850 103.810 ;
        RECT 29.005 103.410 29.295 103.455 ;
        RECT 30.370 103.410 30.690 103.470 ;
        RECT 32.165 103.455 32.455 103.770 ;
        RECT 33.245 103.750 33.535 103.795 ;
        RECT 36.825 103.750 37.115 103.795 ;
        RECT 38.660 103.750 38.950 103.795 ;
        RECT 33.245 103.610 38.950 103.750 ;
        RECT 33.245 103.565 33.535 103.610 ;
        RECT 36.825 103.565 37.115 103.610 ;
        RECT 38.660 103.565 38.950 103.610 ;
        RECT 40.050 103.750 40.340 103.795 ;
        RECT 41.885 103.750 42.175 103.795 ;
        RECT 45.465 103.750 45.755 103.795 ;
        RECT 40.050 103.610 45.755 103.750 ;
        RECT 40.050 103.565 40.340 103.610 ;
        RECT 41.885 103.565 42.175 103.610 ;
        RECT 45.465 103.565 45.755 103.610 ;
        RECT 29.005 103.270 30.690 103.410 ;
        RECT 29.005 103.225 29.295 103.270 ;
        RECT 30.370 103.210 30.690 103.270 ;
        RECT 31.865 103.410 32.455 103.455 ;
        RECT 34.510 103.410 34.830 103.470 ;
        RECT 46.545 103.455 46.835 103.770 ;
        RECT 49.780 103.750 49.920 103.890 ;
        RECT 56.605 103.750 56.895 103.795 ;
        RECT 59.810 103.750 60.130 103.810 ;
        RECT 49.780 103.610 60.130 103.750 ;
        RECT 56.605 103.565 56.895 103.610 ;
        RECT 59.810 103.550 60.130 103.610 ;
        RECT 35.105 103.410 35.755 103.455 ;
        RECT 31.865 103.270 35.755 103.410 ;
        RECT 31.865 103.225 32.155 103.270 ;
        RECT 34.510 103.210 34.830 103.270 ;
        RECT 35.105 103.225 35.755 103.270 ;
        RECT 43.245 103.410 43.895 103.455 ;
        RECT 46.545 103.410 47.135 103.455 ;
        RECT 49.230 103.410 49.550 103.470 ;
        RECT 43.245 103.270 49.550 103.410 ;
        RECT 43.245 103.225 43.895 103.270 ;
        RECT 46.845 103.225 47.135 103.270 ;
        RECT 49.230 103.210 49.550 103.270 ;
        RECT 49.690 103.210 50.010 103.470 ;
        RECT 58.445 103.410 58.735 103.455 ;
        RECT 60.730 103.410 61.050 103.470 ;
        RECT 61.605 103.455 61.895 103.770 ;
        RECT 62.685 103.750 62.975 103.795 ;
        RECT 66.265 103.750 66.555 103.795 ;
        RECT 68.100 103.750 68.390 103.795 ;
        RECT 79.590 103.770 79.910 103.810 ;
        RECT 62.685 103.610 68.390 103.750 ;
        RECT 62.685 103.565 62.975 103.610 ;
        RECT 66.265 103.565 66.555 103.610 ;
        RECT 68.100 103.565 68.390 103.610 ;
        RECT 79.545 103.550 79.910 103.770 ;
        RECT 80.625 103.750 80.915 103.795 ;
        RECT 84.205 103.750 84.495 103.795 ;
        RECT 86.040 103.750 86.330 103.795 ;
        RECT 80.625 103.610 86.330 103.750 ;
        RECT 80.625 103.565 80.915 103.610 ;
        RECT 84.205 103.565 84.495 103.610 ;
        RECT 86.040 103.565 86.330 103.610 ;
        RECT 58.445 103.270 61.050 103.410 ;
        RECT 58.445 103.225 58.735 103.270 ;
        RECT 60.730 103.210 61.050 103.270 ;
        RECT 61.305 103.410 61.895 103.455 ;
        RECT 62.110 103.410 62.430 103.470 ;
        RECT 64.545 103.410 65.195 103.455 ;
        RECT 61.305 103.270 65.195 103.410 ;
        RECT 61.305 103.225 61.595 103.270 ;
        RECT 62.110 103.210 62.430 103.270 ;
        RECT 64.545 103.225 65.195 103.270 ;
        RECT 74.070 103.410 74.390 103.470 ;
        RECT 79.545 103.455 79.835 103.550 ;
        RECT 76.385 103.410 76.675 103.455 ;
        RECT 74.070 103.270 76.675 103.410 ;
        RECT 74.070 103.210 74.390 103.270 ;
        RECT 76.385 103.225 76.675 103.270 ;
        RECT 79.245 103.410 79.835 103.455 ;
        RECT 82.485 103.410 83.135 103.455 ;
        RECT 79.245 103.270 83.135 103.410 ;
        RECT 79.245 103.225 79.535 103.270 ;
        RECT 82.485 103.225 83.135 103.270 ;
        RECT 86.965 103.225 87.255 103.455 ;
        RECT 87.410 103.410 87.730 103.470 ;
        RECT 90.125 103.455 90.415 103.770 ;
        RECT 91.205 103.750 91.495 103.795 ;
        RECT 94.785 103.750 95.075 103.795 ;
        RECT 96.620 103.750 96.910 103.795 ;
        RECT 91.205 103.610 96.910 103.750 ;
        RECT 91.205 103.565 91.495 103.610 ;
        RECT 94.785 103.565 95.075 103.610 ;
        RECT 96.620 103.565 96.910 103.610 ;
        RECT 99.385 103.750 99.675 103.795 ;
        RECT 100.290 103.750 100.610 103.810 ;
        RECT 99.385 103.610 100.610 103.750 ;
        RECT 99.385 103.565 99.675 103.610 ;
        RECT 100.290 103.550 100.610 103.610 ;
        RECT 103.990 103.750 104.280 103.795 ;
        RECT 105.825 103.750 106.115 103.795 ;
        RECT 109.405 103.750 109.695 103.795 ;
        RECT 103.990 103.610 109.695 103.750 ;
        RECT 103.990 103.565 104.280 103.610 ;
        RECT 105.825 103.565 106.115 103.610 ;
        RECT 109.405 103.565 109.695 103.610 ;
        RECT 110.485 103.455 110.775 103.770 ;
        RECT 89.825 103.410 90.415 103.455 ;
        RECT 93.065 103.410 93.715 103.455 ;
        RECT 87.410 103.270 93.715 103.410 ;
        RECT 86.030 103.070 86.350 103.130 ;
        RECT 87.040 103.070 87.180 103.225 ;
        RECT 87.410 103.210 87.730 103.270 ;
        RECT 89.825 103.225 90.115 103.270 ;
        RECT 93.065 103.225 93.715 103.270 ;
        RECT 107.185 103.410 107.835 103.455 ;
        RECT 110.485 103.410 111.075 103.455 ;
        RECT 111.330 103.410 111.650 103.470 ;
        RECT 107.185 103.270 111.650 103.410 ;
        RECT 107.185 103.225 107.835 103.270 ;
        RECT 110.785 103.225 111.075 103.270 ;
        RECT 111.330 103.210 111.650 103.270 ;
        RECT 114.105 103.410 114.395 103.455 ;
        RECT 115.930 103.410 116.250 103.470 ;
        RECT 114.105 103.270 116.250 103.410 ;
        RECT 114.105 103.225 114.395 103.270 ;
        RECT 115.930 103.210 116.250 103.270 ;
        RECT 116.390 103.410 116.710 103.470 ;
        RECT 117.265 103.455 117.555 103.770 ;
        RECT 118.345 103.750 118.635 103.795 ;
        RECT 121.925 103.750 122.215 103.795 ;
        RECT 123.760 103.750 124.050 103.795 ;
        RECT 118.345 103.610 124.050 103.750 ;
        RECT 118.345 103.565 118.635 103.610 ;
        RECT 121.925 103.565 122.215 103.610 ;
        RECT 123.760 103.565 124.050 103.610 ;
        RECT 126.050 103.550 126.370 103.810 ;
        RECT 116.965 103.410 117.555 103.455 ;
        RECT 120.205 103.410 120.855 103.455 ;
        RECT 116.390 103.270 120.855 103.410 ;
        RECT 116.390 103.210 116.710 103.270 ;
        RECT 116.965 103.225 117.255 103.270 ;
        RECT 120.205 103.225 120.855 103.270 ;
        RECT 86.030 102.930 87.180 103.070 ;
        RECT 86.030 102.870 86.350 102.930 ;
        RECT 125.130 102.870 125.450 103.130 ;
        RECT 14.660 102.250 127.820 102.730 ;
        RECT 62.110 101.850 62.430 102.110 ;
        RECT 64.870 101.850 65.190 102.110 ;
        RECT 119.150 102.050 119.470 102.110 ;
        RECT 119.625 102.050 119.915 102.095 ;
        RECT 119.150 101.910 119.915 102.050 ;
        RECT 119.150 101.850 119.470 101.910 ;
        RECT 119.625 101.865 119.915 101.910 ;
        RECT 76.370 101.710 76.690 101.770 ;
        RECT 125.130 101.710 125.450 101.770 ;
        RECT 76.370 101.570 125.450 101.710 ;
        RECT 76.370 101.510 76.690 101.570 ;
        RECT 125.130 101.510 125.450 101.570 ;
        RECT 59.810 101.370 60.130 101.430 ;
        RECT 61.665 101.370 61.955 101.415 ;
        RECT 64.425 101.370 64.715 101.415 ;
        RECT 59.810 101.230 64.715 101.370 ;
        RECT 59.810 101.170 60.130 101.230 ;
        RECT 61.665 101.185 61.955 101.230 ;
        RECT 64.425 101.185 64.715 101.230 ;
        RECT 118.690 101.370 119.010 101.430 ;
        RECT 119.165 101.370 119.455 101.415 ;
        RECT 118.690 101.230 119.455 101.370 ;
        RECT 118.690 101.170 119.010 101.230 ;
        RECT 119.165 101.185 119.455 101.230 ;
        RECT 14.660 99.530 127.820 100.010 ;
        RECT 133.330 76.630 136.060 77.830 ;
        RECT 137.920 77.810 143.450 77.960 ;
        RECT 21.115 74.380 23.065 74.390 ;
        RECT 19.415 73.240 23.065 74.380 ;
        RECT 19.415 73.230 21.125 73.240 ;
        RECT 28.135 73.230 30.305 74.410 ;
        RECT 32.315 74.390 34.265 74.400 ;
        RECT 30.615 73.250 34.265 74.390 ;
        RECT 30.615 73.240 32.325 73.250 ;
        RECT 39.425 73.200 41.595 74.380 ;
        RECT 43.535 74.360 45.485 74.370 ;
        RECT 41.835 73.220 45.485 74.360 ;
        RECT 54.785 74.340 56.735 74.350 ;
        RECT 41.835 73.210 43.545 73.220 ;
        RECT 3.910 73.080 6.100 73.190 ;
        RECT 50.005 73.140 52.175 74.320 ;
        RECT 53.085 73.200 56.735 74.340 ;
        RECT 53.085 73.190 54.795 73.200 ;
        RECT 61.425 73.170 63.595 74.350 ;
        RECT 66.005 74.330 67.955 74.340 ;
        RECT 64.305 73.190 67.955 74.330 ;
        RECT 64.305 73.180 66.015 73.190 ;
        RECT 72.535 73.180 74.705 74.360 ;
        RECT 77.245 74.320 79.195 74.330 ;
        RECT 75.545 73.180 79.195 74.320 ;
        RECT 75.545 73.170 77.255 73.180 ;
        RECT 83.805 73.170 85.975 74.350 ;
        RECT 88.495 74.330 90.445 74.340 ;
        RECT 86.795 73.190 90.445 74.330 ;
        RECT 99.775 74.320 101.725 74.330 ;
        RECT 86.795 73.180 88.505 73.190 ;
        RECT 94.995 73.110 97.165 74.290 ;
        RECT 98.075 73.180 101.725 74.320 ;
        RECT 98.075 73.170 99.785 73.180 ;
        RECT 106.405 73.160 108.575 74.340 ;
        RECT 111.045 74.320 112.995 74.330 ;
        RECT 109.345 73.180 112.995 74.320 ;
        RECT 109.345 73.170 111.055 73.180 ;
        RECT 117.605 73.160 119.775 74.340 ;
        RECT 122.295 74.320 124.245 74.330 ;
        RECT 120.595 73.180 124.245 74.320 ;
        RECT 129.455 73.240 131.625 74.420 ;
        RECT 120.595 73.170 122.305 73.180 ;
        RECT 3.910 72.820 12.240 73.080 ;
        RECT 29.635 72.840 43.235 72.850 ;
        RECT 18.435 72.820 43.235 72.840 ;
        RECT 3.910 72.800 54.455 72.820 ;
        RECT 3.910 72.790 65.705 72.800 ;
        RECT 133.960 72.790 135.640 76.630 ;
        RECT 137.190 76.610 143.450 77.810 ;
        RECT 137.920 75.460 143.450 76.610 ;
        RECT 3.910 72.780 76.925 72.790 ;
        RECT 85.815 72.780 99.415 72.790 ;
        RECT 132.085 72.780 140.600 72.790 ;
        RECT 3.910 71.700 140.600 72.780 ;
        RECT 3.910 71.690 32.035 71.700 ;
        RECT 3.910 71.670 19.135 71.690 ;
        RECT 40.855 71.670 140.600 71.700 ;
        RECT 3.910 71.500 12.240 71.670 ;
        RECT 52.105 71.650 140.600 71.670 ;
        RECT 63.325 71.640 140.600 71.650 ;
        RECT 74.565 71.630 88.165 71.640 ;
        RECT 97.095 71.630 133.215 71.640 ;
        RECT 3.910 71.370 6.100 71.500 ;
        RECT 10.800 71.180 11.950 71.500 ;
        RECT 10.800 69.480 11.915 71.180 ;
        RECT 29.635 71.170 43.285 71.180 ;
        RECT 15.510 71.155 17.040 71.160 ;
        RECT 18.435 71.155 43.285 71.170 ;
        RECT 12.285 71.150 43.285 71.155 ;
        RECT 12.285 71.130 54.505 71.150 ;
        RECT 141.810 71.140 143.230 75.460 ;
        RECT 12.285 71.120 65.755 71.130 ;
        RECT 12.285 71.110 76.975 71.120 ;
        RECT 85.815 71.110 99.465 71.120 ;
        RECT 140.220 71.110 143.240 71.140 ;
        RECT 12.285 70.030 143.240 71.110 ;
        RECT 12.285 70.020 32.085 70.030 ;
        RECT 12.285 70.005 19.375 70.020 ;
        RECT 10.800 13.800 11.950 69.480 ;
        RECT 12.320 15.450 13.470 70.005 ;
        RECT 15.510 68.660 17.040 70.005 ;
        RECT 40.855 70.000 143.240 70.030 ;
        RECT 52.105 69.980 143.240 70.000 ;
        RECT 63.325 69.970 143.240 69.980 ;
        RECT 74.565 69.960 88.215 69.970 ;
        RECT 97.095 69.960 143.240 69.970 ;
        RECT 140.220 69.910 143.240 69.960 ;
        RECT 29.645 69.670 43.315 69.680 ;
        RECT 18.445 69.650 43.315 69.670 ;
        RECT 18.445 69.630 54.535 69.650 ;
        RECT 18.445 69.620 65.785 69.630 ;
        RECT 139.590 69.620 150.610 69.640 ;
        RECT 18.445 69.610 77.005 69.620 ;
        RECT 85.825 69.610 99.495 69.620 ;
        RECT 132.155 69.610 150.610 69.620 ;
        RECT 18.445 69.570 150.610 69.610 ;
        RECT 18.445 68.530 150.740 69.570 ;
        RECT 18.445 68.520 32.115 68.530 ;
        RECT 40.865 68.500 150.740 68.530 ;
        RECT 52.115 68.490 143.320 68.500 ;
        RECT 52.115 68.480 140.670 68.490 ;
        RECT 63.335 68.470 140.670 68.480 ;
        RECT 74.575 68.460 88.245 68.470 ;
        RECT 97.105 68.460 133.295 68.470 ;
        RECT 141.080 68.450 142.300 68.490 ;
        RECT 149.360 68.470 150.740 68.500 ;
        RECT 29.655 68.100 43.325 68.110 ;
        RECT 13.950 68.080 43.325 68.100 ;
        RECT 13.950 68.060 54.545 68.080 ;
        RECT 13.950 68.050 65.795 68.060 ;
        RECT 13.950 68.040 77.015 68.050 ;
        RECT 85.835 68.040 99.505 68.050 ;
        RECT 139.530 68.040 143.320 68.060 ;
        RECT 13.950 66.960 152.870 68.040 ;
        RECT 13.950 66.950 32.125 66.960 ;
        RECT 13.950 18.530 15.100 66.950 ;
        RECT 40.875 66.930 152.870 66.960 ;
        RECT 52.125 66.910 152.870 66.930 ;
        RECT 63.345 66.900 152.870 66.910 ;
        RECT 74.585 66.890 88.255 66.900 ;
        RECT 97.115 66.890 143.320 66.900 ;
        RECT 141.030 66.770 142.490 66.890 ;
        RECT 21.405 65.510 26.555 65.790 ;
        RECT 27.815 65.490 28.965 65.800 ;
        RECT 32.605 65.520 37.755 65.800 ;
        RECT 39.015 65.500 40.165 65.810 ;
        RECT 43.825 65.490 48.975 65.770 ;
        RECT 50.235 65.470 51.385 65.780 ;
        RECT 149.460 65.760 150.600 65.780 ;
        RECT 55.075 65.470 60.225 65.750 ;
        RECT 61.485 65.450 62.635 65.760 ;
        RECT 66.295 65.460 71.445 65.740 ;
        RECT 72.705 65.440 73.855 65.750 ;
        RECT 77.535 65.450 82.685 65.730 ;
        RECT 83.945 65.430 85.095 65.740 ;
        RECT 88.785 65.460 93.935 65.740 ;
        RECT 95.195 65.440 96.345 65.750 ;
        RECT 100.065 65.450 105.215 65.730 ;
        RECT 106.475 65.430 107.625 65.740 ;
        RECT 111.335 65.450 116.485 65.730 ;
        RECT 117.745 65.430 118.895 65.740 ;
        RECT 122.585 65.450 127.735 65.730 ;
        RECT 128.995 65.430 130.145 65.740 ;
        RECT 133.315 65.430 138.455 65.690 ;
        RECT 21.205 65.140 21.435 65.320 ;
        RECT 26.495 65.190 26.725 65.320 ;
        RECT 21.125 55.220 21.485 65.140 ;
        RECT 26.435 55.240 26.805 65.190 ;
        RECT 27.635 65.150 27.865 65.320 ;
        RECT 27.565 55.200 27.935 65.150 ;
        RECT 28.925 65.140 29.155 65.320 ;
        RECT 32.405 65.150 32.635 65.330 ;
        RECT 37.695 65.200 37.925 65.330 ;
        RECT 28.835 55.250 29.255 65.140 ;
        RECT 32.325 55.230 32.685 65.150 ;
        RECT 37.635 55.250 38.005 65.200 ;
        RECT 38.835 65.160 39.065 65.330 ;
        RECT 38.765 55.210 39.135 65.160 ;
        RECT 40.125 65.150 40.355 65.330 ;
        RECT 40.035 55.260 40.455 65.150 ;
        RECT 43.625 65.120 43.855 65.300 ;
        RECT 48.915 65.170 49.145 65.300 ;
        RECT 43.545 55.200 43.905 65.120 ;
        RECT 48.855 55.220 49.225 65.170 ;
        RECT 50.055 65.130 50.285 65.300 ;
        RECT 49.985 55.180 50.355 65.130 ;
        RECT 51.345 65.120 51.575 65.300 ;
        RECT 51.255 55.230 51.675 65.120 ;
        RECT 54.875 65.100 55.105 65.280 ;
        RECT 60.165 65.150 60.395 65.280 ;
        RECT 54.795 55.180 55.155 65.100 ;
        RECT 60.105 55.200 60.475 65.150 ;
        RECT 61.305 65.110 61.535 65.280 ;
        RECT 61.235 55.160 61.605 65.110 ;
        RECT 62.595 65.100 62.825 65.280 ;
        RECT 62.505 55.210 62.925 65.100 ;
        RECT 66.095 65.090 66.325 65.270 ;
        RECT 71.385 65.140 71.615 65.270 ;
        RECT 66.015 55.170 66.375 65.090 ;
        RECT 71.325 55.190 71.695 65.140 ;
        RECT 72.525 65.100 72.755 65.270 ;
        RECT 72.455 55.150 72.825 65.100 ;
        RECT 73.815 65.090 74.045 65.270 ;
        RECT 73.725 55.200 74.145 65.090 ;
        RECT 77.335 65.080 77.565 65.260 ;
        RECT 82.625 65.130 82.855 65.260 ;
        RECT 77.255 55.160 77.615 65.080 ;
        RECT 82.565 55.180 82.935 65.130 ;
        RECT 83.765 65.090 83.995 65.260 ;
        RECT 83.695 55.140 84.065 65.090 ;
        RECT 85.055 65.080 85.285 65.260 ;
        RECT 88.585 65.090 88.815 65.270 ;
        RECT 93.875 65.140 94.105 65.270 ;
        RECT 84.965 55.190 85.385 65.080 ;
        RECT 88.505 55.170 88.865 65.090 ;
        RECT 93.815 55.190 94.185 65.140 ;
        RECT 95.015 65.100 95.245 65.270 ;
        RECT 94.945 55.150 95.315 65.100 ;
        RECT 96.305 65.090 96.535 65.270 ;
        RECT 96.215 55.200 96.635 65.090 ;
        RECT 99.865 65.080 100.095 65.260 ;
        RECT 105.155 65.130 105.385 65.260 ;
        RECT 99.785 55.160 100.145 65.080 ;
        RECT 105.095 55.180 105.465 65.130 ;
        RECT 106.295 65.090 106.525 65.260 ;
        RECT 106.225 55.140 106.595 65.090 ;
        RECT 107.585 65.080 107.815 65.260 ;
        RECT 111.135 65.080 111.365 65.260 ;
        RECT 116.425 65.130 116.655 65.260 ;
        RECT 107.495 55.190 107.915 65.080 ;
        RECT 111.055 55.160 111.415 65.080 ;
        RECT 116.365 55.180 116.735 65.130 ;
        RECT 117.565 65.090 117.795 65.260 ;
        RECT 117.495 55.140 117.865 65.090 ;
        RECT 118.855 65.080 119.085 65.260 ;
        RECT 122.385 65.080 122.615 65.260 ;
        RECT 127.675 65.130 127.905 65.260 ;
        RECT 118.765 55.190 119.185 65.080 ;
        RECT 122.305 55.160 122.665 65.080 ;
        RECT 127.615 55.180 127.985 65.130 ;
        RECT 128.815 65.090 129.045 65.260 ;
        RECT 128.745 55.140 129.115 65.090 ;
        RECT 130.105 65.080 130.335 65.260 ;
        RECT 133.135 65.130 133.365 65.230 ;
        RECT 130.015 55.190 130.435 65.080 ;
        RECT 133.005 55.240 133.405 65.130 ;
        RECT 138.425 65.100 138.655 65.230 ;
        RECT 133.135 55.230 133.365 55.240 ;
        RECT 138.345 55.130 138.725 65.100 ;
        RECT 149.340 64.660 150.720 65.760 ;
        RECT 20.815 54.230 25.555 54.530 ;
        RECT 32.015 54.240 36.755 54.540 ;
        RECT 43.235 54.210 47.975 54.510 ;
        RECT 54.485 54.190 59.225 54.490 ;
        RECT 65.705 54.180 70.445 54.480 ;
        RECT 76.945 54.170 81.685 54.470 ;
        RECT 88.195 54.180 92.935 54.480 ;
        RECT 99.475 54.170 104.215 54.470 ;
        RECT 110.745 54.170 115.485 54.470 ;
        RECT 121.995 54.170 126.735 54.470 ;
        RECT 21.655 52.320 22.115 52.550 ;
        RECT 25.625 52.280 26.255 52.560 ;
        RECT 25.735 52.240 26.195 52.280 ;
        RECT 27.665 52.240 28.125 52.470 ;
        RECT 32.855 52.330 33.315 52.560 ;
        RECT 36.825 52.290 37.455 52.570 ;
        RECT 36.935 52.250 37.395 52.290 ;
        RECT 38.865 52.250 39.325 52.480 ;
        RECT 44.075 52.300 44.535 52.530 ;
        RECT 48.045 52.260 48.675 52.540 ;
        RECT 48.155 52.220 48.615 52.260 ;
        RECT 50.085 52.220 50.545 52.450 ;
        RECT 55.325 52.280 55.785 52.510 ;
        RECT 59.295 52.240 59.925 52.520 ;
        RECT 59.405 52.200 59.865 52.240 ;
        RECT 61.335 52.200 61.795 52.430 ;
        RECT 66.545 52.270 67.005 52.500 ;
        RECT 70.515 52.230 71.145 52.510 ;
        RECT 70.625 52.190 71.085 52.230 ;
        RECT 72.555 52.190 73.015 52.420 ;
        RECT 77.785 52.260 78.245 52.490 ;
        RECT 81.755 52.220 82.385 52.500 ;
        RECT 81.865 52.180 82.325 52.220 ;
        RECT 83.795 52.180 84.255 52.410 ;
        RECT 89.035 52.270 89.495 52.500 ;
        RECT 93.005 52.230 93.635 52.510 ;
        RECT 93.115 52.190 93.575 52.230 ;
        RECT 95.045 52.190 95.505 52.420 ;
        RECT 100.315 52.260 100.775 52.490 ;
        RECT 104.285 52.220 104.915 52.500 ;
        RECT 104.395 52.180 104.855 52.220 ;
        RECT 106.325 52.180 106.785 52.410 ;
        RECT 111.585 52.260 112.045 52.490 ;
        RECT 115.555 52.220 116.185 52.500 ;
        RECT 115.665 52.180 116.125 52.220 ;
        RECT 117.595 52.180 118.055 52.410 ;
        RECT 122.835 52.260 123.295 52.490 ;
        RECT 126.805 52.220 127.435 52.500 ;
        RECT 126.915 52.180 127.375 52.220 ;
        RECT 128.845 52.180 129.305 52.410 ;
        RECT 21.375 52.010 21.605 52.115 ;
        RECT 21.245 50.290 21.615 52.010 ;
        RECT 22.165 51.890 22.395 52.115 ;
        RECT 25.455 51.980 25.685 52.035 ;
        RECT 21.375 50.115 21.605 50.290 ;
        RECT 22.155 50.210 22.525 51.890 ;
        RECT 22.165 50.115 22.395 50.210 ;
        RECT 21.525 49.670 22.245 49.930 ;
        RECT 19.295 46.650 20.065 47.720 ;
        RECT 21.385 47.490 22.105 47.750 ;
        RECT 21.225 47.200 21.455 47.340 ;
        RECT 21.085 46.430 21.475 47.200 ;
        RECT 22.015 47.190 22.245 47.340 ;
        RECT 22.005 46.450 22.375 47.190 ;
        RECT 25.305 47.010 25.735 51.980 ;
        RECT 26.245 51.970 26.475 52.035 ;
        RECT 27.385 51.970 27.615 52.035 ;
        RECT 26.185 46.970 26.585 51.970 ;
        RECT 27.265 46.970 27.665 51.970 ;
        RECT 28.175 51.940 28.405 52.035 ;
        RECT 32.575 52.020 32.805 52.125 ;
        RECT 28.115 46.970 28.545 51.940 ;
        RECT 32.445 50.300 32.815 52.020 ;
        RECT 33.365 51.900 33.595 52.125 ;
        RECT 36.655 51.990 36.885 52.045 ;
        RECT 32.575 50.125 32.805 50.300 ;
        RECT 33.355 50.220 33.725 51.900 ;
        RECT 33.365 50.125 33.595 50.220 ;
        RECT 32.725 49.680 33.445 49.940 ;
        RECT 25.735 46.600 26.195 46.830 ;
        RECT 27.665 46.710 28.125 46.830 ;
        RECT 27.515 46.600 28.125 46.710 ;
        RECT 30.495 46.660 31.265 47.730 ;
        RECT 32.585 47.500 33.305 47.760 ;
        RECT 32.425 47.210 32.655 47.350 ;
        RECT 21.225 46.340 21.455 46.430 ;
        RECT 22.015 46.340 22.245 46.450 ;
        RECT 27.515 46.430 28.095 46.600 ;
        RECT 32.285 46.440 32.675 47.210 ;
        RECT 33.215 47.200 33.445 47.350 ;
        RECT 33.205 46.460 33.575 47.200 ;
        RECT 36.505 47.020 36.935 51.990 ;
        RECT 37.445 51.980 37.675 52.045 ;
        RECT 38.585 51.980 38.815 52.045 ;
        RECT 37.385 46.980 37.785 51.980 ;
        RECT 38.465 46.980 38.865 51.980 ;
        RECT 39.375 51.950 39.605 52.045 ;
        RECT 43.795 51.990 44.025 52.095 ;
        RECT 39.315 46.980 39.745 51.950 ;
        RECT 43.665 50.270 44.035 51.990 ;
        RECT 44.585 51.870 44.815 52.095 ;
        RECT 47.875 51.960 48.105 52.015 ;
        RECT 43.795 50.095 44.025 50.270 ;
        RECT 44.575 50.190 44.945 51.870 ;
        RECT 44.585 50.095 44.815 50.190 ;
        RECT 43.945 49.650 44.665 49.910 ;
        RECT 36.935 46.610 37.395 46.840 ;
        RECT 38.865 46.720 39.325 46.840 ;
        RECT 38.715 46.610 39.325 46.720 ;
        RECT 41.715 46.630 42.485 47.700 ;
        RECT 43.805 47.470 44.525 47.730 ;
        RECT 43.645 47.180 43.875 47.320 ;
        RECT 32.425 46.350 32.655 46.440 ;
        RECT 33.215 46.350 33.445 46.460 ;
        RECT 38.715 46.440 39.295 46.610 ;
        RECT 43.505 46.410 43.895 47.180 ;
        RECT 44.435 47.170 44.665 47.320 ;
        RECT 44.425 46.430 44.795 47.170 ;
        RECT 47.725 46.990 48.155 51.960 ;
        RECT 48.665 51.950 48.895 52.015 ;
        RECT 49.805 51.950 50.035 52.015 ;
        RECT 48.605 46.950 49.005 51.950 ;
        RECT 49.685 46.950 50.085 51.950 ;
        RECT 50.595 51.920 50.825 52.015 ;
        RECT 55.045 51.970 55.275 52.075 ;
        RECT 50.535 46.950 50.965 51.920 ;
        RECT 54.915 50.250 55.285 51.970 ;
        RECT 55.835 51.850 56.065 52.075 ;
        RECT 59.125 51.940 59.355 51.995 ;
        RECT 55.045 50.075 55.275 50.250 ;
        RECT 55.825 50.170 56.195 51.850 ;
        RECT 55.835 50.075 56.065 50.170 ;
        RECT 55.195 49.630 55.915 49.890 ;
        RECT 48.155 46.580 48.615 46.810 ;
        RECT 50.085 46.690 50.545 46.810 ;
        RECT 49.935 46.580 50.545 46.690 ;
        RECT 52.965 46.610 53.735 47.680 ;
        RECT 55.055 47.450 55.775 47.710 ;
        RECT 54.895 47.160 55.125 47.300 ;
        RECT 43.645 46.320 43.875 46.410 ;
        RECT 44.435 46.320 44.665 46.430 ;
        RECT 49.935 46.410 50.515 46.580 ;
        RECT 54.755 46.390 55.145 47.160 ;
        RECT 55.685 47.150 55.915 47.300 ;
        RECT 55.675 46.410 56.045 47.150 ;
        RECT 58.975 46.970 59.405 51.940 ;
        RECT 59.915 51.930 60.145 51.995 ;
        RECT 61.055 51.930 61.285 51.995 ;
        RECT 59.855 46.930 60.255 51.930 ;
        RECT 60.935 46.930 61.335 51.930 ;
        RECT 61.845 51.900 62.075 51.995 ;
        RECT 66.265 51.960 66.495 52.065 ;
        RECT 61.785 46.930 62.215 51.900 ;
        RECT 66.135 50.240 66.505 51.960 ;
        RECT 67.055 51.840 67.285 52.065 ;
        RECT 70.345 51.930 70.575 51.985 ;
        RECT 66.265 50.065 66.495 50.240 ;
        RECT 67.045 50.160 67.415 51.840 ;
        RECT 67.055 50.065 67.285 50.160 ;
        RECT 66.415 49.620 67.135 49.880 ;
        RECT 59.405 46.560 59.865 46.790 ;
        RECT 61.335 46.670 61.795 46.790 ;
        RECT 61.185 46.560 61.795 46.670 ;
        RECT 64.185 46.600 64.955 47.670 ;
        RECT 66.275 47.440 66.995 47.700 ;
        RECT 66.115 47.150 66.345 47.290 ;
        RECT 54.895 46.300 55.125 46.390 ;
        RECT 55.685 46.300 55.915 46.410 ;
        RECT 61.185 46.390 61.765 46.560 ;
        RECT 65.975 46.380 66.365 47.150 ;
        RECT 66.905 47.140 67.135 47.290 ;
        RECT 66.895 46.400 67.265 47.140 ;
        RECT 70.195 46.960 70.625 51.930 ;
        RECT 71.135 51.920 71.365 51.985 ;
        RECT 72.275 51.920 72.505 51.985 ;
        RECT 71.075 46.920 71.475 51.920 ;
        RECT 72.155 46.920 72.555 51.920 ;
        RECT 73.065 51.890 73.295 51.985 ;
        RECT 77.505 51.950 77.735 52.055 ;
        RECT 73.005 46.920 73.435 51.890 ;
        RECT 77.375 50.230 77.745 51.950 ;
        RECT 78.295 51.830 78.525 52.055 ;
        RECT 81.585 51.920 81.815 51.975 ;
        RECT 77.505 50.055 77.735 50.230 ;
        RECT 78.285 50.150 78.655 51.830 ;
        RECT 78.295 50.055 78.525 50.150 ;
        RECT 77.655 49.610 78.375 49.870 ;
        RECT 70.625 46.550 71.085 46.780 ;
        RECT 72.555 46.660 73.015 46.780 ;
        RECT 72.405 46.550 73.015 46.660 ;
        RECT 75.425 46.590 76.195 47.660 ;
        RECT 77.515 47.430 78.235 47.690 ;
        RECT 77.355 47.140 77.585 47.280 ;
        RECT 66.115 46.290 66.345 46.380 ;
        RECT 66.905 46.290 67.135 46.400 ;
        RECT 72.405 46.380 72.985 46.550 ;
        RECT 77.215 46.370 77.605 47.140 ;
        RECT 78.145 47.130 78.375 47.280 ;
        RECT 78.135 46.390 78.505 47.130 ;
        RECT 81.435 46.950 81.865 51.920 ;
        RECT 82.375 51.910 82.605 51.975 ;
        RECT 83.515 51.910 83.745 51.975 ;
        RECT 82.315 46.910 82.715 51.910 ;
        RECT 83.395 46.910 83.795 51.910 ;
        RECT 84.305 51.880 84.535 51.975 ;
        RECT 88.755 51.960 88.985 52.065 ;
        RECT 84.245 46.910 84.675 51.880 ;
        RECT 88.625 50.240 88.995 51.960 ;
        RECT 89.545 51.840 89.775 52.065 ;
        RECT 92.835 51.930 93.065 51.985 ;
        RECT 88.755 50.065 88.985 50.240 ;
        RECT 89.535 50.160 89.905 51.840 ;
        RECT 89.545 50.065 89.775 50.160 ;
        RECT 88.905 49.620 89.625 49.880 ;
        RECT 81.865 46.540 82.325 46.770 ;
        RECT 83.795 46.650 84.255 46.770 ;
        RECT 83.645 46.540 84.255 46.650 ;
        RECT 86.675 46.600 87.445 47.670 ;
        RECT 88.765 47.440 89.485 47.700 ;
        RECT 88.605 47.150 88.835 47.290 ;
        RECT 77.355 46.280 77.585 46.370 ;
        RECT 78.145 46.280 78.375 46.390 ;
        RECT 83.645 46.370 84.225 46.540 ;
        RECT 88.465 46.380 88.855 47.150 ;
        RECT 89.395 47.140 89.625 47.290 ;
        RECT 89.385 46.400 89.755 47.140 ;
        RECT 92.685 46.960 93.115 51.930 ;
        RECT 93.625 51.920 93.855 51.985 ;
        RECT 94.765 51.920 94.995 51.985 ;
        RECT 93.565 46.920 93.965 51.920 ;
        RECT 94.645 46.920 95.045 51.920 ;
        RECT 95.555 51.890 95.785 51.985 ;
        RECT 100.035 51.950 100.265 52.055 ;
        RECT 95.495 46.920 95.925 51.890 ;
        RECT 99.905 50.230 100.275 51.950 ;
        RECT 100.825 51.830 101.055 52.055 ;
        RECT 104.115 51.920 104.345 51.975 ;
        RECT 100.035 50.055 100.265 50.230 ;
        RECT 100.815 50.150 101.185 51.830 ;
        RECT 100.825 50.055 101.055 50.150 ;
        RECT 100.185 49.610 100.905 49.870 ;
        RECT 93.115 46.550 93.575 46.780 ;
        RECT 95.045 46.660 95.505 46.780 ;
        RECT 94.895 46.550 95.505 46.660 ;
        RECT 97.955 46.590 98.725 47.660 ;
        RECT 100.045 47.430 100.765 47.690 ;
        RECT 99.885 47.140 100.115 47.280 ;
        RECT 88.605 46.290 88.835 46.380 ;
        RECT 89.395 46.290 89.625 46.400 ;
        RECT 94.895 46.380 95.475 46.550 ;
        RECT 99.745 46.370 100.135 47.140 ;
        RECT 100.675 47.130 100.905 47.280 ;
        RECT 100.665 46.390 101.035 47.130 ;
        RECT 103.965 46.950 104.395 51.920 ;
        RECT 104.905 51.910 105.135 51.975 ;
        RECT 106.045 51.910 106.275 51.975 ;
        RECT 104.845 46.910 105.245 51.910 ;
        RECT 105.925 46.910 106.325 51.910 ;
        RECT 106.835 51.880 107.065 51.975 ;
        RECT 111.305 51.950 111.535 52.055 ;
        RECT 106.775 46.910 107.205 51.880 ;
        RECT 111.175 50.230 111.545 51.950 ;
        RECT 112.095 51.830 112.325 52.055 ;
        RECT 115.385 51.920 115.615 51.975 ;
        RECT 111.305 50.055 111.535 50.230 ;
        RECT 112.085 50.150 112.455 51.830 ;
        RECT 112.095 50.055 112.325 50.150 ;
        RECT 111.455 49.610 112.175 49.870 ;
        RECT 104.395 46.540 104.855 46.770 ;
        RECT 106.325 46.650 106.785 46.770 ;
        RECT 106.175 46.540 106.785 46.650 ;
        RECT 109.225 46.590 109.995 47.660 ;
        RECT 111.315 47.430 112.035 47.690 ;
        RECT 111.155 47.140 111.385 47.280 ;
        RECT 99.885 46.280 100.115 46.370 ;
        RECT 100.675 46.280 100.905 46.390 ;
        RECT 106.175 46.370 106.755 46.540 ;
        RECT 111.015 46.370 111.405 47.140 ;
        RECT 111.945 47.130 112.175 47.280 ;
        RECT 111.935 46.390 112.305 47.130 ;
        RECT 115.235 46.950 115.665 51.920 ;
        RECT 116.175 51.910 116.405 51.975 ;
        RECT 117.315 51.910 117.545 51.975 ;
        RECT 116.115 46.910 116.515 51.910 ;
        RECT 117.195 46.910 117.595 51.910 ;
        RECT 118.105 51.880 118.335 51.975 ;
        RECT 122.555 51.950 122.785 52.055 ;
        RECT 118.045 46.910 118.475 51.880 ;
        RECT 122.425 50.230 122.795 51.950 ;
        RECT 123.345 51.830 123.575 52.055 ;
        RECT 126.635 51.920 126.865 51.975 ;
        RECT 122.555 50.055 122.785 50.230 ;
        RECT 123.335 50.150 123.705 51.830 ;
        RECT 123.345 50.055 123.575 50.150 ;
        RECT 122.705 49.610 123.425 49.870 ;
        RECT 115.665 46.540 116.125 46.770 ;
        RECT 117.595 46.650 118.055 46.770 ;
        RECT 117.445 46.540 118.055 46.650 ;
        RECT 120.475 46.590 121.245 47.660 ;
        RECT 122.565 47.430 123.285 47.690 ;
        RECT 122.405 47.140 122.635 47.280 ;
        RECT 111.155 46.280 111.385 46.370 ;
        RECT 111.945 46.280 112.175 46.390 ;
        RECT 117.445 46.370 118.025 46.540 ;
        RECT 122.265 46.370 122.655 47.140 ;
        RECT 123.195 47.130 123.425 47.280 ;
        RECT 123.185 46.390 123.555 47.130 ;
        RECT 126.485 46.950 126.915 51.920 ;
        RECT 127.425 51.910 127.655 51.975 ;
        RECT 128.565 51.910 128.795 51.975 ;
        RECT 127.365 46.910 127.765 51.910 ;
        RECT 128.445 46.910 128.845 51.910 ;
        RECT 129.355 51.880 129.585 51.975 ;
        RECT 129.295 46.910 129.725 51.880 ;
        RECT 126.915 46.540 127.375 46.770 ;
        RECT 128.845 46.650 129.305 46.770 ;
        RECT 128.695 46.540 129.305 46.650 ;
        RECT 122.405 46.280 122.635 46.370 ;
        RECT 123.195 46.280 123.425 46.390 ;
        RECT 128.695 46.370 129.275 46.540 ;
        RECT 21.505 45.950 21.965 46.180 ;
        RECT 32.705 45.960 33.165 46.190 ;
        RECT 43.925 45.930 44.385 46.160 ;
        RECT 55.175 45.910 55.635 46.140 ;
        RECT 66.395 45.900 66.855 46.130 ;
        RECT 77.635 45.890 78.095 46.120 ;
        RECT 88.885 45.900 89.345 46.130 ;
        RECT 100.165 45.890 100.625 46.120 ;
        RECT 111.435 45.890 111.895 46.120 ;
        RECT 122.685 45.890 123.145 46.120 ;
        RECT 29.055 45.020 41.225 45.030 ;
        RECT 17.855 45.005 41.225 45.020 ;
        RECT 15.900 45.000 41.225 45.005 ;
        RECT 15.900 44.980 52.445 45.000 ;
        RECT 15.900 44.970 63.695 44.980 ;
        RECT 15.900 44.960 74.915 44.970 ;
        RECT 85.235 44.960 97.405 44.970 ;
        RECT 15.900 43.880 131.205 44.960 ;
        RECT 15.900 43.870 30.025 43.880 ;
        RECT 15.900 43.855 18.690 43.870 ;
        RECT 15.900 41.620 17.050 43.855 ;
        RECT 40.275 43.850 131.205 43.880 ;
        RECT 51.525 43.830 131.205 43.850 ;
        RECT 62.745 43.820 131.205 43.830 ;
        RECT 73.985 43.810 86.155 43.820 ;
        RECT 96.515 43.810 131.205 43.820 ;
        RECT 29.015 43.330 41.185 43.340 ;
        RECT 17.815 43.310 41.185 43.330 ;
        RECT 142.830 43.320 144.150 43.340 ;
        RECT 17.815 43.290 52.405 43.310 ;
        RECT 140.750 43.300 144.150 43.320 ;
        RECT 17.815 43.280 63.655 43.290 ;
        RECT 119.895 43.280 144.150 43.300 ;
        RECT 17.815 43.270 74.875 43.280 ;
        RECT 85.195 43.270 97.365 43.280 ;
        RECT 108.685 43.270 144.150 43.280 ;
        RECT 17.815 42.180 144.150 43.270 ;
        RECT 18.755 42.150 144.150 42.180 ;
        RECT 18.755 42.120 131.165 42.150 ;
        RECT 18.755 42.090 109.655 42.120 ;
        RECT 18.755 42.080 98.445 42.090 ;
        RECT 41.325 42.070 98.445 42.080 ;
        RECT 142.830 42.070 144.150 42.150 ;
        RECT 41.325 42.060 87.205 42.070 ;
        RECT 75.035 42.050 87.205 42.060 ;
        RECT 15.900 41.540 19.685 41.620 ;
        RECT 142.070 41.610 146.210 41.640 ;
        RECT 119.855 41.590 146.210 41.610 ;
        RECT 108.645 41.550 146.210 41.590 ;
        RECT 15.900 41.520 42.165 41.540 ;
        RECT 97.445 41.530 146.210 41.550 ;
        RECT 15.900 41.510 75.875 41.520 ;
        RECT 86.235 41.510 146.210 41.530 ;
        RECT 15.900 40.500 146.210 41.510 ;
        RECT 15.900 40.480 142.320 40.500 ;
        RECT 15.900 40.470 140.920 40.480 ;
        RECT 18.715 40.460 140.920 40.470 ;
        RECT 142.070 40.460 142.250 40.480 ;
        RECT 18.715 40.440 120.815 40.460 ;
        RECT 18.715 40.400 109.615 40.440 ;
        RECT 18.715 40.390 98.405 40.400 ;
        RECT 41.285 40.380 98.405 40.390 ;
        RECT 41.285 40.370 87.165 40.380 ;
        RECT 74.995 40.360 87.165 40.370 ;
        RECT 26.775 39.230 27.235 39.460 ;
        RECT 38.055 39.230 38.515 39.460 ;
        RECT 49.345 39.210 49.805 39.440 ;
        RECT 60.565 39.210 61.025 39.440 ;
        RECT 71.765 39.210 72.225 39.440 ;
        RECT 83.055 39.200 83.515 39.430 ;
        RECT 94.295 39.220 94.755 39.450 ;
        RECT 105.505 39.240 105.965 39.470 ;
        RECT 116.705 39.280 117.165 39.510 ;
        RECT 127.915 39.300 128.375 39.530 ;
        RECT 20.645 38.810 21.225 38.980 ;
        RECT 26.495 38.960 26.725 39.070 ;
        RECT 27.285 38.980 27.515 39.070 ;
        RECT 20.615 38.700 21.225 38.810 ;
        RECT 20.615 38.580 21.075 38.700 ;
        RECT 22.545 38.580 23.005 38.810 ;
        RECT 20.195 33.470 20.625 38.440 ;
        RECT 20.335 33.375 20.565 33.470 ;
        RECT 21.075 33.440 21.475 38.440 ;
        RECT 22.155 33.440 22.555 38.440 ;
        RECT 21.125 33.375 21.355 33.440 ;
        RECT 22.265 33.375 22.495 33.440 ;
        RECT 23.005 33.430 23.435 38.400 ;
        RECT 26.365 38.220 26.735 38.960 ;
        RECT 26.495 38.070 26.725 38.220 ;
        RECT 27.265 38.210 27.655 38.980 ;
        RECT 31.925 38.810 32.505 38.980 ;
        RECT 37.775 38.960 38.005 39.070 ;
        RECT 38.565 38.980 38.795 39.070 ;
        RECT 27.285 38.070 27.515 38.210 ;
        RECT 26.635 37.660 27.355 37.920 ;
        RECT 28.675 37.690 29.445 38.760 ;
        RECT 31.895 38.700 32.505 38.810 ;
        RECT 31.895 38.580 32.355 38.700 ;
        RECT 33.825 38.580 34.285 38.810 ;
        RECT 26.495 35.480 27.215 35.740 ;
        RECT 26.345 35.200 26.575 35.295 ;
        RECT 26.215 33.520 26.585 35.200 ;
        RECT 27.135 35.120 27.365 35.295 ;
        RECT 23.055 33.375 23.285 33.430 ;
        RECT 26.345 33.295 26.575 33.520 ;
        RECT 27.125 33.400 27.495 35.120 ;
        RECT 31.475 33.470 31.905 38.440 ;
        RECT 27.135 33.295 27.365 33.400 ;
        RECT 31.615 33.375 31.845 33.470 ;
        RECT 32.355 33.440 32.755 38.440 ;
        RECT 33.435 33.440 33.835 38.440 ;
        RECT 32.405 33.375 32.635 33.440 ;
        RECT 33.545 33.375 33.775 33.440 ;
        RECT 34.285 33.430 34.715 38.400 ;
        RECT 37.645 38.220 38.015 38.960 ;
        RECT 37.775 38.070 38.005 38.220 ;
        RECT 38.545 38.210 38.935 38.980 ;
        RECT 43.215 38.790 43.795 38.960 ;
        RECT 49.065 38.940 49.295 39.050 ;
        RECT 49.855 38.960 50.085 39.050 ;
        RECT 38.565 38.070 38.795 38.210 ;
        RECT 37.915 37.660 38.635 37.920 ;
        RECT 39.955 37.690 40.725 38.760 ;
        RECT 43.185 38.680 43.795 38.790 ;
        RECT 43.185 38.560 43.645 38.680 ;
        RECT 45.115 38.560 45.575 38.790 ;
        RECT 37.775 35.480 38.495 35.740 ;
        RECT 37.625 35.200 37.855 35.295 ;
        RECT 37.495 33.520 37.865 35.200 ;
        RECT 38.415 35.120 38.645 35.295 ;
        RECT 34.335 33.375 34.565 33.430 ;
        RECT 37.625 33.295 37.855 33.520 ;
        RECT 38.405 33.400 38.775 35.120 ;
        RECT 42.765 33.450 43.195 38.420 ;
        RECT 38.415 33.295 38.645 33.400 ;
        RECT 42.905 33.355 43.135 33.450 ;
        RECT 43.645 33.420 44.045 38.420 ;
        RECT 44.725 33.420 45.125 38.420 ;
        RECT 43.695 33.355 43.925 33.420 ;
        RECT 44.835 33.355 45.065 33.420 ;
        RECT 45.575 33.410 46.005 38.380 ;
        RECT 48.935 38.200 49.305 38.940 ;
        RECT 49.065 38.050 49.295 38.200 ;
        RECT 49.835 38.190 50.225 38.960 ;
        RECT 54.435 38.790 55.015 38.960 ;
        RECT 60.285 38.940 60.515 39.050 ;
        RECT 61.075 38.960 61.305 39.050 ;
        RECT 49.855 38.050 50.085 38.190 ;
        RECT 49.205 37.640 49.925 37.900 ;
        RECT 51.245 37.670 52.015 38.740 ;
        RECT 54.405 38.680 55.015 38.790 ;
        RECT 54.405 38.560 54.865 38.680 ;
        RECT 56.335 38.560 56.795 38.790 ;
        RECT 49.065 35.460 49.785 35.720 ;
        RECT 48.915 35.180 49.145 35.275 ;
        RECT 48.785 33.500 49.155 35.180 ;
        RECT 49.705 35.100 49.935 35.275 ;
        RECT 45.625 33.355 45.855 33.410 ;
        RECT 48.915 33.275 49.145 33.500 ;
        RECT 49.695 33.380 50.065 35.100 ;
        RECT 53.985 33.450 54.415 38.420 ;
        RECT 49.705 33.275 49.935 33.380 ;
        RECT 54.125 33.355 54.355 33.450 ;
        RECT 54.865 33.420 55.265 38.420 ;
        RECT 55.945 33.420 56.345 38.420 ;
        RECT 54.915 33.355 55.145 33.420 ;
        RECT 56.055 33.355 56.285 33.420 ;
        RECT 56.795 33.410 57.225 38.380 ;
        RECT 60.155 38.200 60.525 38.940 ;
        RECT 60.285 38.050 60.515 38.200 ;
        RECT 61.055 38.190 61.445 38.960 ;
        RECT 65.635 38.790 66.215 38.960 ;
        RECT 71.485 38.940 71.715 39.050 ;
        RECT 72.275 38.960 72.505 39.050 ;
        RECT 61.075 38.050 61.305 38.190 ;
        RECT 60.425 37.640 61.145 37.900 ;
        RECT 62.465 37.670 63.235 38.740 ;
        RECT 65.605 38.680 66.215 38.790 ;
        RECT 65.605 38.560 66.065 38.680 ;
        RECT 67.535 38.560 67.995 38.790 ;
        RECT 60.285 35.460 61.005 35.720 ;
        RECT 60.135 35.180 60.365 35.275 ;
        RECT 60.005 33.500 60.375 35.180 ;
        RECT 60.925 35.100 61.155 35.275 ;
        RECT 56.845 33.355 57.075 33.410 ;
        RECT 60.135 33.275 60.365 33.500 ;
        RECT 60.915 33.380 61.285 35.100 ;
        RECT 65.185 33.450 65.615 38.420 ;
        RECT 60.925 33.275 61.155 33.380 ;
        RECT 65.325 33.355 65.555 33.450 ;
        RECT 66.065 33.420 66.465 38.420 ;
        RECT 67.145 33.420 67.545 38.420 ;
        RECT 66.115 33.355 66.345 33.420 ;
        RECT 67.255 33.355 67.485 33.420 ;
        RECT 67.995 33.410 68.425 38.380 ;
        RECT 71.355 38.200 71.725 38.940 ;
        RECT 71.485 38.050 71.715 38.200 ;
        RECT 72.255 38.190 72.645 38.960 ;
        RECT 76.925 38.780 77.505 38.950 ;
        RECT 82.775 38.930 83.005 39.040 ;
        RECT 83.565 38.950 83.795 39.040 ;
        RECT 72.275 38.050 72.505 38.190 ;
        RECT 71.625 37.640 72.345 37.900 ;
        RECT 73.665 37.670 74.435 38.740 ;
        RECT 76.895 38.670 77.505 38.780 ;
        RECT 76.895 38.550 77.355 38.670 ;
        RECT 78.825 38.550 79.285 38.780 ;
        RECT 71.485 35.460 72.205 35.720 ;
        RECT 71.335 35.180 71.565 35.275 ;
        RECT 71.205 33.500 71.575 35.180 ;
        RECT 72.125 35.100 72.355 35.275 ;
        RECT 68.045 33.355 68.275 33.410 ;
        RECT 71.335 33.275 71.565 33.500 ;
        RECT 72.115 33.380 72.485 35.100 ;
        RECT 76.475 33.440 76.905 38.410 ;
        RECT 72.125 33.275 72.355 33.380 ;
        RECT 76.615 33.345 76.845 33.440 ;
        RECT 77.355 33.410 77.755 38.410 ;
        RECT 78.435 33.410 78.835 38.410 ;
        RECT 77.405 33.345 77.635 33.410 ;
        RECT 78.545 33.345 78.775 33.410 ;
        RECT 79.285 33.400 79.715 38.370 ;
        RECT 82.645 38.190 83.015 38.930 ;
        RECT 82.775 38.040 83.005 38.190 ;
        RECT 83.545 38.180 83.935 38.950 ;
        RECT 88.165 38.800 88.745 38.970 ;
        RECT 94.015 38.950 94.245 39.060 ;
        RECT 94.805 38.970 95.035 39.060 ;
        RECT 83.565 38.040 83.795 38.180 ;
        RECT 82.915 37.630 83.635 37.890 ;
        RECT 84.955 37.660 85.725 38.730 ;
        RECT 88.135 38.690 88.745 38.800 ;
        RECT 88.135 38.570 88.595 38.690 ;
        RECT 90.065 38.570 90.525 38.800 ;
        RECT 82.775 35.450 83.495 35.710 ;
        RECT 82.625 35.170 82.855 35.265 ;
        RECT 82.495 33.490 82.865 35.170 ;
        RECT 83.415 35.090 83.645 35.265 ;
        RECT 79.335 33.345 79.565 33.400 ;
        RECT 82.625 33.265 82.855 33.490 ;
        RECT 83.405 33.370 83.775 35.090 ;
        RECT 87.715 33.460 88.145 38.430 ;
        RECT 83.415 33.265 83.645 33.370 ;
        RECT 87.855 33.365 88.085 33.460 ;
        RECT 88.595 33.430 88.995 38.430 ;
        RECT 89.675 33.430 90.075 38.430 ;
        RECT 88.645 33.365 88.875 33.430 ;
        RECT 89.785 33.365 90.015 33.430 ;
        RECT 90.525 33.420 90.955 38.390 ;
        RECT 93.885 38.210 94.255 38.950 ;
        RECT 94.015 38.060 94.245 38.210 ;
        RECT 94.785 38.200 95.175 38.970 ;
        RECT 99.375 38.820 99.955 38.990 ;
        RECT 105.225 38.970 105.455 39.080 ;
        RECT 106.015 38.990 106.245 39.080 ;
        RECT 94.805 38.060 95.035 38.200 ;
        RECT 94.155 37.650 94.875 37.910 ;
        RECT 96.195 37.680 96.965 38.750 ;
        RECT 99.345 38.710 99.955 38.820 ;
        RECT 99.345 38.590 99.805 38.710 ;
        RECT 101.275 38.590 101.735 38.820 ;
        RECT 94.015 35.470 94.735 35.730 ;
        RECT 93.865 35.190 94.095 35.285 ;
        RECT 93.735 33.510 94.105 35.190 ;
        RECT 94.655 35.110 94.885 35.285 ;
        RECT 90.575 33.365 90.805 33.420 ;
        RECT 93.865 33.285 94.095 33.510 ;
        RECT 94.645 33.390 95.015 35.110 ;
        RECT 98.925 33.480 99.355 38.450 ;
        RECT 94.655 33.285 94.885 33.390 ;
        RECT 99.065 33.385 99.295 33.480 ;
        RECT 99.805 33.450 100.205 38.450 ;
        RECT 100.885 33.450 101.285 38.450 ;
        RECT 99.855 33.385 100.085 33.450 ;
        RECT 100.995 33.385 101.225 33.450 ;
        RECT 101.735 33.440 102.165 38.410 ;
        RECT 105.095 38.230 105.465 38.970 ;
        RECT 105.225 38.080 105.455 38.230 ;
        RECT 105.995 38.220 106.385 38.990 ;
        RECT 110.575 38.860 111.155 39.030 ;
        RECT 116.425 39.010 116.655 39.120 ;
        RECT 117.215 39.030 117.445 39.120 ;
        RECT 106.015 38.080 106.245 38.220 ;
        RECT 105.365 37.670 106.085 37.930 ;
        RECT 107.405 37.700 108.175 38.770 ;
        RECT 110.545 38.750 111.155 38.860 ;
        RECT 110.545 38.630 111.005 38.750 ;
        RECT 112.475 38.630 112.935 38.860 ;
        RECT 105.225 35.490 105.945 35.750 ;
        RECT 105.075 35.210 105.305 35.305 ;
        RECT 104.945 33.530 105.315 35.210 ;
        RECT 105.865 35.130 106.095 35.305 ;
        RECT 101.785 33.385 102.015 33.440 ;
        RECT 105.075 33.305 105.305 33.530 ;
        RECT 105.855 33.410 106.225 35.130 ;
        RECT 110.125 33.520 110.555 38.490 ;
        RECT 110.265 33.425 110.495 33.520 ;
        RECT 111.005 33.490 111.405 38.490 ;
        RECT 112.085 33.490 112.485 38.490 ;
        RECT 111.055 33.425 111.285 33.490 ;
        RECT 112.195 33.425 112.425 33.490 ;
        RECT 112.935 33.480 113.365 38.450 ;
        RECT 116.295 38.270 116.665 39.010 ;
        RECT 116.425 38.120 116.655 38.270 ;
        RECT 117.195 38.260 117.585 39.030 ;
        RECT 121.785 38.880 122.365 39.050 ;
        RECT 127.635 39.030 127.865 39.140 ;
        RECT 128.425 39.050 128.655 39.140 ;
        RECT 117.215 38.120 117.445 38.260 ;
        RECT 116.565 37.710 117.285 37.970 ;
        RECT 118.605 37.740 119.375 38.810 ;
        RECT 121.755 38.770 122.365 38.880 ;
        RECT 121.755 38.650 122.215 38.770 ;
        RECT 123.685 38.650 124.145 38.880 ;
        RECT 116.425 35.530 117.145 35.790 ;
        RECT 116.275 35.250 116.505 35.345 ;
        RECT 116.145 33.570 116.515 35.250 ;
        RECT 117.065 35.170 117.295 35.345 ;
        RECT 112.985 33.425 113.215 33.480 ;
        RECT 105.865 33.305 106.095 33.410 ;
        RECT 116.275 33.345 116.505 33.570 ;
        RECT 117.055 33.450 117.425 35.170 ;
        RECT 121.335 33.540 121.765 38.510 ;
        RECT 117.065 33.345 117.295 33.450 ;
        RECT 121.475 33.445 121.705 33.540 ;
        RECT 122.215 33.510 122.615 38.510 ;
        RECT 123.295 33.510 123.695 38.510 ;
        RECT 122.265 33.445 122.495 33.510 ;
        RECT 123.405 33.445 123.635 33.510 ;
        RECT 124.145 33.500 124.575 38.470 ;
        RECT 127.505 38.290 127.875 39.030 ;
        RECT 127.635 38.140 127.865 38.290 ;
        RECT 128.405 38.280 128.795 39.050 ;
        RECT 128.425 38.140 128.655 38.280 ;
        RECT 127.775 37.730 128.495 37.990 ;
        RECT 129.815 37.760 130.585 38.830 ;
        RECT 142.850 37.630 144.170 38.900 ;
        RECT 127.635 35.550 128.355 35.810 ;
        RECT 127.485 35.270 127.715 35.365 ;
        RECT 127.355 33.590 127.725 35.270 ;
        RECT 128.275 35.190 128.505 35.365 ;
        RECT 124.195 33.445 124.425 33.500 ;
        RECT 127.485 33.365 127.715 33.590 ;
        RECT 128.265 33.470 128.635 35.190 ;
        RECT 128.275 33.365 128.505 33.470 ;
        RECT 20.615 32.940 21.075 33.170 ;
        RECT 22.545 33.130 23.005 33.170 ;
        RECT 22.485 32.850 23.115 33.130 ;
        RECT 26.625 32.860 27.085 33.090 ;
        RECT 31.895 32.940 32.355 33.170 ;
        RECT 33.825 33.130 34.285 33.170 ;
        RECT 33.765 32.850 34.395 33.130 ;
        RECT 37.905 32.860 38.365 33.090 ;
        RECT 43.185 32.920 43.645 33.150 ;
        RECT 45.115 33.110 45.575 33.150 ;
        RECT 45.055 32.830 45.685 33.110 ;
        RECT 49.195 32.840 49.655 33.070 ;
        RECT 54.405 32.920 54.865 33.150 ;
        RECT 56.335 33.110 56.795 33.150 ;
        RECT 56.275 32.830 56.905 33.110 ;
        RECT 60.415 32.840 60.875 33.070 ;
        RECT 65.605 32.920 66.065 33.150 ;
        RECT 67.535 33.110 67.995 33.150 ;
        RECT 67.475 32.830 68.105 33.110 ;
        RECT 71.615 32.840 72.075 33.070 ;
        RECT 76.895 32.910 77.355 33.140 ;
        RECT 78.825 33.100 79.285 33.140 ;
        RECT 78.765 32.820 79.395 33.100 ;
        RECT 82.905 32.830 83.365 33.060 ;
        RECT 88.135 32.930 88.595 33.160 ;
        RECT 90.065 33.120 90.525 33.160 ;
        RECT 90.005 32.840 90.635 33.120 ;
        RECT 94.145 32.850 94.605 33.080 ;
        RECT 99.345 32.950 99.805 33.180 ;
        RECT 101.275 33.140 101.735 33.180 ;
        RECT 101.215 32.860 101.845 33.140 ;
        RECT 105.355 32.870 105.815 33.100 ;
        RECT 110.545 32.990 111.005 33.220 ;
        RECT 112.475 33.180 112.935 33.220 ;
        RECT 112.415 32.900 113.045 33.180 ;
        RECT 116.555 32.910 117.015 33.140 ;
        RECT 121.755 33.010 122.215 33.240 ;
        RECT 123.685 33.200 124.145 33.240 ;
        RECT 123.625 32.920 124.255 33.200 ;
        RECT 127.765 32.930 128.225 33.160 ;
        RECT 23.185 30.880 27.925 31.180 ;
        RECT 34.465 30.880 39.205 31.180 ;
        RECT 45.755 30.860 50.495 31.160 ;
        RECT 56.975 30.860 61.715 31.160 ;
        RECT 68.175 30.860 72.915 31.160 ;
        RECT 79.465 30.850 84.205 31.150 ;
        RECT 90.705 30.870 95.445 31.170 ;
        RECT 101.915 30.890 106.655 31.190 ;
        RECT 113.115 30.930 117.855 31.230 ;
        RECT 124.325 30.950 129.065 31.250 ;
        RECT 19.485 20.270 19.905 30.160 ;
        RECT 19.585 20.090 19.815 20.270 ;
        RECT 20.805 20.260 21.175 30.210 ;
        RECT 20.875 20.090 21.105 20.260 ;
        RECT 21.935 20.220 22.305 30.170 ;
        RECT 27.255 20.270 27.615 30.190 ;
        RECT 30.765 20.270 31.185 30.160 ;
        RECT 22.015 20.090 22.245 20.220 ;
        RECT 27.305 20.090 27.535 20.270 ;
        RECT 30.865 20.090 31.095 20.270 ;
        RECT 32.085 20.260 32.455 30.210 ;
        RECT 32.155 20.090 32.385 20.260 ;
        RECT 33.215 20.220 33.585 30.170 ;
        RECT 38.535 20.270 38.895 30.190 ;
        RECT 33.295 20.090 33.525 20.220 ;
        RECT 38.585 20.090 38.815 20.270 ;
        RECT 42.055 20.250 42.475 30.140 ;
        RECT 42.155 20.070 42.385 20.250 ;
        RECT 43.375 20.240 43.745 30.190 ;
        RECT 43.445 20.070 43.675 20.240 ;
        RECT 44.505 20.200 44.875 30.150 ;
        RECT 49.825 20.250 50.185 30.170 ;
        RECT 53.275 20.250 53.695 30.140 ;
        RECT 44.585 20.070 44.815 20.200 ;
        RECT 49.875 20.070 50.105 20.250 ;
        RECT 53.375 20.070 53.605 20.250 ;
        RECT 54.595 20.240 54.965 30.190 ;
        RECT 54.665 20.070 54.895 20.240 ;
        RECT 55.725 20.200 56.095 30.150 ;
        RECT 61.045 20.250 61.405 30.170 ;
        RECT 64.475 20.250 64.895 30.140 ;
        RECT 55.805 20.070 56.035 20.200 ;
        RECT 61.095 20.070 61.325 20.250 ;
        RECT 64.575 20.070 64.805 20.250 ;
        RECT 65.795 20.240 66.165 30.190 ;
        RECT 65.865 20.070 66.095 20.240 ;
        RECT 66.925 20.200 67.295 30.150 ;
        RECT 72.245 20.250 72.605 30.170 ;
        RECT 67.005 20.070 67.235 20.200 ;
        RECT 72.295 20.070 72.525 20.250 ;
        RECT 75.765 20.240 76.185 30.130 ;
        RECT 75.865 20.060 76.095 20.240 ;
        RECT 77.085 20.230 77.455 30.180 ;
        RECT 77.155 20.060 77.385 20.230 ;
        RECT 78.215 20.190 78.585 30.140 ;
        RECT 83.535 20.240 83.895 30.160 ;
        RECT 87.005 20.260 87.425 30.150 ;
        RECT 78.295 20.060 78.525 20.190 ;
        RECT 83.585 20.060 83.815 20.240 ;
        RECT 87.105 20.080 87.335 20.260 ;
        RECT 88.325 20.250 88.695 30.200 ;
        RECT 88.395 20.080 88.625 20.250 ;
        RECT 89.455 20.210 89.825 30.160 ;
        RECT 94.775 20.260 95.135 30.180 ;
        RECT 98.215 20.280 98.635 30.170 ;
        RECT 89.535 20.080 89.765 20.210 ;
        RECT 94.825 20.080 95.055 20.260 ;
        RECT 98.315 20.100 98.545 20.280 ;
        RECT 99.535 20.270 99.905 30.220 ;
        RECT 99.605 20.100 99.835 20.270 ;
        RECT 100.665 20.230 101.035 30.180 ;
        RECT 105.985 20.280 106.345 30.200 ;
        RECT 109.415 20.320 109.835 30.210 ;
        RECT 100.745 20.100 100.975 20.230 ;
        RECT 106.035 20.100 106.265 20.280 ;
        RECT 109.515 20.140 109.745 20.320 ;
        RECT 110.735 20.310 111.105 30.260 ;
        RECT 110.805 20.140 111.035 20.310 ;
        RECT 111.865 20.270 112.235 30.220 ;
        RECT 117.185 20.320 117.545 30.240 ;
        RECT 120.625 20.340 121.045 30.230 ;
        RECT 111.945 20.140 112.175 20.270 ;
        RECT 117.235 20.140 117.465 20.320 ;
        RECT 120.725 20.160 120.955 20.340 ;
        RECT 121.945 20.330 122.315 30.280 ;
        RECT 122.015 20.160 122.245 20.330 ;
        RECT 123.075 20.290 123.445 30.240 ;
        RECT 128.395 20.340 128.755 30.260 ;
        RECT 123.155 20.160 123.385 20.290 ;
        RECT 128.445 20.160 128.675 20.340 ;
        RECT 132.345 20.170 132.755 30.180 ;
        RECT 137.735 30.120 137.965 30.130 ;
        RECT 132.445 20.130 132.675 20.170 ;
        RECT 137.665 20.080 138.055 30.120 ;
        RECT 19.775 19.610 20.925 19.920 ;
        RECT 22.185 19.620 27.335 19.900 ;
        RECT 31.055 19.610 32.205 19.920 ;
        RECT 33.465 19.620 38.615 19.900 ;
        RECT 42.345 19.590 43.495 19.900 ;
        RECT 44.755 19.600 49.905 19.880 ;
        RECT 53.565 19.590 54.715 19.900 ;
        RECT 55.975 19.600 61.125 19.880 ;
        RECT 64.765 19.590 65.915 19.900 ;
        RECT 67.175 19.600 72.325 19.880 ;
        RECT 76.055 19.580 77.205 19.890 ;
        RECT 78.465 19.590 83.615 19.870 ;
        RECT 87.295 19.600 88.445 19.910 ;
        RECT 89.705 19.610 94.855 19.890 ;
        RECT 98.505 19.620 99.655 19.930 ;
        RECT 100.915 19.630 106.065 19.910 ;
        RECT 109.705 19.660 110.855 19.970 ;
        RECT 112.115 19.670 117.265 19.950 ;
        RECT 120.915 19.680 122.065 19.990 ;
        RECT 123.325 19.690 128.475 19.970 ;
        RECT 132.635 19.640 138.025 19.930 ;
        RECT 142.940 19.110 144.080 37.630 ;
        RECT 13.940 18.460 17.635 18.530 ;
        RECT 117.755 18.510 131.425 18.530 ;
        RECT 106.545 18.470 131.425 18.510 ;
        RECT 13.940 18.440 41.565 18.460 ;
        RECT 95.345 18.450 131.425 18.470 ;
        RECT 13.940 18.430 75.275 18.440 ;
        RECT 84.135 18.430 131.425 18.450 ;
        RECT 13.940 17.380 131.425 18.430 ;
        RECT 142.890 17.990 144.140 19.110 ;
        RECT 145.070 18.880 146.210 40.500 ;
        RECT 145.030 17.960 146.250 18.880 ;
        RECT 13.950 17.370 15.100 17.380 ;
        RECT 16.615 17.360 120.215 17.380 ;
        RECT 16.615 17.320 109.015 17.360 ;
        RECT 16.615 17.310 97.805 17.320 ;
        RECT 39.185 17.300 97.805 17.310 ;
        RECT 39.185 17.290 86.565 17.300 ;
        RECT 72.895 17.280 86.565 17.290 ;
        RECT 117.765 16.950 140.620 16.960 ;
        RECT 142.040 16.950 148.010 16.980 ;
        RECT 117.765 16.940 148.010 16.950 ;
        RECT 106.555 16.900 148.010 16.940 ;
        RECT 16.625 16.870 41.575 16.890 ;
        RECT 95.355 16.880 148.010 16.900 ;
        RECT 16.625 16.860 75.285 16.870 ;
        RECT 84.145 16.860 148.010 16.880 ;
        RECT 16.625 15.840 148.010 16.860 ;
        RECT 16.625 15.820 142.660 15.840 ;
        RECT 16.625 15.810 140.620 15.820 ;
        RECT 142.040 15.810 142.660 15.820 ;
        RECT 16.625 15.790 120.225 15.810 ;
        RECT 16.625 15.750 109.025 15.790 ;
        RECT 16.625 15.740 97.815 15.750 ;
        RECT 39.195 15.730 97.815 15.740 ;
        RECT 39.195 15.720 86.575 15.730 ;
        RECT 72.905 15.710 86.575 15.720 ;
        RECT 131.215 15.460 132.585 15.470 ;
        RECT 12.290 15.390 17.625 15.450 ;
        RECT 117.795 15.440 132.785 15.460 ;
        RECT 106.585 15.400 132.785 15.440 ;
        RECT 12.290 15.370 41.585 15.390 ;
        RECT 95.385 15.380 132.785 15.400 ;
        RECT 12.290 15.360 75.295 15.370 ;
        RECT 84.175 15.360 132.785 15.380 ;
        RECT 12.290 14.320 132.785 15.360 ;
        RECT 142.905 15.040 144.045 15.050 ;
        RECT 12.290 14.310 131.445 14.320 ;
        RECT 12.290 14.300 120.235 14.310 ;
        RECT 12.320 14.280 13.470 14.300 ;
        RECT 16.655 14.290 120.235 14.300 ;
        RECT 16.655 14.250 109.035 14.290 ;
        RECT 16.655 14.240 97.825 14.250 ;
        RECT 39.225 14.230 97.825 14.240 ;
        RECT 39.225 14.220 86.585 14.230 ;
        RECT 72.935 14.210 86.585 14.220 ;
        RECT 142.850 13.920 144.100 15.040 ;
        RECT 145.020 14.870 146.160 14.980 ;
        RECT 144.980 13.950 146.200 14.870 ;
        RECT 16.965 13.800 17.435 13.810 ;
        RECT 10.800 13.780 17.435 13.800 ;
        RECT 10.800 13.720 17.555 13.780 ;
        RECT 117.845 13.770 131.445 13.790 ;
        RECT 106.635 13.730 131.445 13.770 ;
        RECT 10.800 13.700 41.585 13.720 ;
        RECT 95.435 13.710 131.445 13.730 ;
        RECT 10.800 13.690 75.295 13.700 ;
        RECT 84.225 13.690 131.445 13.710 ;
        RECT 10.800 12.650 131.445 13.690 ;
        RECT 16.705 12.640 131.445 12.650 ;
        RECT 16.705 12.620 120.235 12.640 ;
        RECT 16.705 12.580 109.035 12.620 ;
        RECT 16.705 12.570 97.825 12.580 ;
        RECT 39.275 12.560 97.825 12.570 ;
        RECT 39.275 12.550 86.585 12.560 ;
        RECT 72.985 12.540 86.585 12.550 ;
        RECT 128.755 12.240 130.465 12.250 ;
        RECT 117.545 12.220 119.255 12.230 ;
        RECT 106.345 12.180 108.055 12.190 ;
        RECT 27.615 12.170 29.325 12.180 ;
        RECT 38.895 12.170 40.605 12.180 ;
        RECT 25.675 11.030 29.325 12.170 ;
        RECT 36.955 11.030 40.605 12.170 ;
        RECT 95.135 12.160 96.845 12.170 ;
        RECT 50.185 12.150 51.895 12.160 ;
        RECT 61.405 12.150 63.115 12.160 ;
        RECT 72.605 12.150 74.315 12.160 ;
        RECT 25.675 11.020 27.625 11.030 ;
        RECT 36.955 11.020 38.905 11.030 ;
        RECT 48.245 11.010 51.895 12.150 ;
        RECT 59.465 11.010 63.115 12.150 ;
        RECT 70.665 11.010 74.315 12.150 ;
        RECT 83.895 12.140 85.605 12.150 ;
        RECT 48.245 11.000 50.195 11.010 ;
        RECT 59.465 11.000 61.415 11.010 ;
        RECT 70.665 11.000 72.615 11.010 ;
        RECT 81.955 11.000 85.605 12.140 ;
        RECT 93.195 11.020 96.845 12.160 ;
        RECT 104.405 11.040 108.055 12.180 ;
        RECT 115.605 11.080 119.255 12.220 ;
        RECT 126.815 11.100 130.465 12.240 ;
        RECT 126.815 11.090 128.765 11.100 ;
        RECT 115.605 11.070 117.555 11.080 ;
        RECT 104.405 11.030 106.355 11.040 ;
        RECT 93.195 11.010 95.145 11.020 ;
        RECT 81.955 10.990 83.905 11.000 ;
        RECT 142.905 8.580 144.045 13.920 ;
        RECT 74.420 7.440 144.045 8.580 ;
        RECT 74.420 1.410 75.560 7.440 ;
        RECT 145.020 6.630 146.160 13.950 ;
        RECT 93.650 5.490 146.160 6.630 ;
        RECT 93.650 1.480 94.790 5.490 ;
        RECT 146.870 4.560 148.010 15.840 ;
        RECT 113.130 3.420 148.010 4.560 ;
        RECT 113.130 1.610 114.270 3.420 ;
        RECT 149.460 2.770 150.600 64.660 ;
        RECT 131.940 1.880 150.600 2.770 ;
        RECT 131.800 1.630 150.600 1.880 ;
        RECT 74.290 0.160 75.680 1.410 ;
        RECT 93.500 0.230 94.890 1.480 ;
        RECT 112.900 0.360 114.290 1.610 ;
        RECT 131.800 1.380 133.490 1.630 ;
        RECT 151.730 1.420 152.870 66.900 ;
        RECT 131.800 0.430 133.540 1.380 ;
        RECT 113.130 0.330 114.270 0.360 ;
        RECT 151.600 0.300 152.970 1.420 ;
        RECT 93.650 0.150 94.790 0.230 ;
      LAYER met2 ;
        RECT 135.390 223.830 136.740 225.230 ;
        RECT 138.180 223.760 139.530 225.160 ;
        RECT 143.230 223.790 144.580 225.190 ;
        RECT 16.880 211.105 18.760 211.475 ;
        RECT 46.880 211.105 48.760 211.475 ;
        RECT 76.880 211.105 78.760 211.475 ;
        RECT 106.880 211.105 108.760 211.475 ;
        RECT 31.880 208.385 33.760 208.755 ;
        RECT 61.880 208.385 63.760 208.755 ;
        RECT 91.880 208.385 93.760 208.755 ;
        RECT 121.880 208.385 123.760 208.755 ;
        RECT 16.880 205.665 18.760 206.035 ;
        RECT 46.880 205.665 48.760 206.035 ;
        RECT 76.880 205.665 78.760 206.035 ;
        RECT 106.880 205.665 108.760 206.035 ;
        RECT 63.980 204.500 64.240 204.820 ;
        RECT 61.220 203.480 61.480 203.800 ;
        RECT 31.880 202.945 33.760 203.315 ;
        RECT 61.280 202.100 61.420 203.480 ;
        RECT 61.880 202.945 63.760 203.315 ;
        RECT 61.220 201.780 61.480 202.100 ;
        RECT 16.880 200.225 18.760 200.595 ;
        RECT 46.880 200.225 48.760 200.595 ;
        RECT 31.880 197.505 33.760 197.875 ;
        RECT 61.880 197.505 63.760 197.875 ;
        RECT 64.040 196.320 64.180 204.500 ;
        RECT 73.180 204.160 73.440 204.480 ;
        RECT 74.560 204.160 74.820 204.480 ;
        RECT 67.200 203.480 67.460 203.800 ;
        RECT 66.740 199.060 67.000 199.380 ;
        RECT 66.800 197.340 66.940 199.060 ;
        RECT 65.820 197.020 66.080 197.340 ;
        RECT 66.740 197.020 67.000 197.340 ;
        RECT 63.980 196.000 64.240 196.320 ;
        RECT 61.680 195.320 61.940 195.640 ;
        RECT 16.880 194.785 18.760 195.155 ;
        RECT 46.880 194.785 48.760 195.155 ;
        RECT 61.740 194.280 61.880 195.320 ;
        RECT 55.240 194.020 55.500 194.280 ;
        RECT 55.240 193.960 55.900 194.020 ;
        RECT 61.680 193.960 61.940 194.280 ;
        RECT 55.300 193.880 55.900 193.960 ;
        RECT 46.040 192.600 46.300 192.920 ;
        RECT 52.940 192.600 53.200 192.920 ;
        RECT 31.880 192.065 33.760 192.435 ;
        RECT 42.820 190.900 43.080 191.220 ;
        RECT 16.880 189.345 18.760 189.715 ;
        RECT 42.880 188.500 43.020 190.900 ;
        RECT 46.100 190.540 46.240 192.600 ;
        RECT 49.260 190.560 49.520 190.880 ;
        RECT 46.040 190.220 46.300 190.540 ;
        RECT 46.880 189.345 48.760 189.715 ;
        RECT 42.820 188.180 43.080 188.500 ;
        RECT 41.900 187.840 42.160 188.160 ;
        RECT 31.880 186.625 33.760 186.995 ;
        RECT 41.960 185.780 42.100 187.840 ;
        RECT 31.320 185.460 31.580 185.780 ;
        RECT 41.900 185.460 42.160 185.780 ;
        RECT 42.360 185.460 42.620 185.780 ;
        RECT 16.880 183.905 18.760 184.275 ;
        RECT 31.380 183.740 31.520 185.460 ;
        RECT 34.080 185.120 34.340 185.440 ;
        RECT 32.700 184.440 32.960 184.760 ;
        RECT 31.320 183.420 31.580 183.740 ;
        RECT 30.400 182.400 30.660 182.720 ;
        RECT 23.040 179.680 23.300 180.000 ;
        RECT 16.880 178.465 18.760 178.835 ;
        RECT 23.100 173.940 23.240 179.680 ;
        RECT 26.260 179.340 26.520 179.660 ;
        RECT 26.320 178.300 26.460 179.340 ;
        RECT 30.460 179.320 30.600 182.400 ;
        RECT 30.400 179.000 30.660 179.320 ;
        RECT 30.860 179.000 31.120 179.320 ;
        RECT 26.260 177.980 26.520 178.300 ;
        RECT 29.940 176.620 30.200 176.940 ;
        RECT 30.000 175.580 30.140 176.620 ;
        RECT 29.940 175.260 30.200 175.580 ;
        RECT 29.940 174.580 30.200 174.900 ;
        RECT 22.640 173.800 23.240 173.940 ;
        RECT 16.880 173.025 18.760 173.395 ;
        RECT 22.640 171.840 22.780 173.800 ;
        RECT 22.580 171.520 22.840 171.840 ;
        RECT 22.640 169.120 22.780 171.520 ;
        RECT 30.000 169.460 30.140 174.580 ;
        RECT 30.460 171.840 30.600 179.000 ;
        RECT 30.920 177.280 31.060 179.000 ;
        RECT 31.380 177.620 31.520 183.420 ;
        RECT 32.760 183.400 32.900 184.440 ;
        RECT 32.700 183.080 32.960 183.400 ;
        RECT 31.880 181.185 33.760 181.555 ;
        RECT 34.140 180.000 34.280 185.120 ;
        RECT 36.380 184.440 36.640 184.760 ;
        RECT 35.460 183.080 35.720 183.400 ;
        RECT 35.920 183.080 36.180 183.400 ;
        RECT 35.520 180.680 35.660 183.080 ;
        RECT 35.980 181.020 36.120 183.080 ;
        RECT 35.920 180.700 36.180 181.020 ;
        RECT 35.460 180.360 35.720 180.680 ;
        RECT 36.440 180.000 36.580 184.440 ;
        RECT 34.080 179.680 34.340 180.000 ;
        RECT 35.920 179.680 36.180 180.000 ;
        RECT 36.380 179.680 36.640 180.000 ;
        RECT 31.320 177.300 31.580 177.620 ;
        RECT 30.860 176.960 31.120 177.280 ;
        RECT 30.920 174.560 31.060 176.960 ;
        RECT 30.860 174.240 31.120 174.560 ;
        RECT 30.400 171.520 30.660 171.840 ;
        RECT 29.940 169.140 30.200 169.460 ;
        RECT 22.580 168.800 22.840 169.120 ;
        RECT 22.120 168.120 22.380 168.440 ;
        RECT 16.880 167.585 18.760 167.955 ;
        RECT 22.180 167.080 22.320 168.120 ;
        RECT 22.120 166.760 22.380 167.080 ;
        RECT 17.980 165.400 18.240 165.720 ;
        RECT 21.660 165.400 21.920 165.720 ;
        RECT 18.040 164.700 18.180 165.400 ;
        RECT 17.980 164.380 18.240 164.700 ;
        RECT 21.200 163.930 21.460 164.020 ;
        RECT 21.720 163.930 21.860 165.400 ;
        RECT 21.200 163.790 21.860 163.930 ;
        RECT 21.200 163.700 21.460 163.790 ;
        RECT 16.880 162.145 18.760 162.515 ;
        RECT 17.980 161.320 18.240 161.640 ;
        RECT 18.040 159.260 18.180 161.320 ;
        RECT 17.980 158.940 18.240 159.260 ;
        RECT 21.260 158.580 21.400 163.700 ;
        RECT 22.640 163.340 22.780 168.800 ;
        RECT 28.560 166.420 28.820 166.740 ;
        RECT 25.340 166.080 25.600 166.400 ;
        RECT 25.400 164.700 25.540 166.080 ;
        RECT 25.340 164.380 25.600 164.700 ;
        RECT 22.580 163.020 22.840 163.340 ;
        RECT 21.660 162.680 21.920 163.000 ;
        RECT 21.720 160.280 21.860 162.680 ;
        RECT 21.660 159.960 21.920 160.280 ;
        RECT 21.200 158.260 21.460 158.580 ;
        RECT 19.820 157.240 20.080 157.560 ;
        RECT 16.880 156.705 18.760 157.075 ;
        RECT 19.880 155.860 20.020 157.240 ;
        RECT 19.820 155.540 20.080 155.860 ;
        RECT 21.260 153.140 21.400 158.260 ;
        RECT 21.720 157.560 21.860 159.960 ;
        RECT 22.640 158.240 22.780 163.020 ;
        RECT 28.620 161.980 28.760 166.420 ;
        RECT 30.000 163.680 30.140 169.140 ;
        RECT 30.460 166.740 30.600 171.520 ;
        RECT 30.400 166.420 30.660 166.740 ;
        RECT 30.920 166.060 31.060 174.240 ;
        RECT 30.860 165.740 31.120 166.060 ;
        RECT 29.940 163.360 30.200 163.680 ;
        RECT 31.380 163.000 31.520 177.300 ;
        RECT 31.880 175.745 33.760 176.115 ;
        RECT 35.980 174.900 36.120 179.680 ;
        RECT 41.960 177.280 42.100 185.460 ;
        RECT 42.420 185.100 42.560 185.460 ;
        RECT 42.880 185.100 43.020 188.180 ;
        RECT 49.320 186.460 49.460 190.560 ;
        RECT 53.000 190.540 53.140 192.600 ;
        RECT 52.940 190.220 53.200 190.540 ;
        RECT 51.100 189.880 51.360 190.200 ;
        RECT 51.160 188.500 51.300 189.880 ;
        RECT 55.760 188.500 55.900 193.880 ;
        RECT 56.620 193.280 56.880 193.600 ;
        RECT 56.680 191.220 56.820 193.280 ;
        RECT 61.880 192.065 63.760 192.435 ;
        RECT 56.620 190.900 56.880 191.220 ;
        RECT 58.000 190.900 58.260 191.220 ;
        RECT 51.100 188.180 51.360 188.500 ;
        RECT 53.400 188.180 53.660 188.500 ;
        RECT 55.700 188.180 55.960 188.500 ;
        RECT 49.260 186.140 49.520 186.460 ;
        RECT 42.360 184.780 42.620 185.100 ;
        RECT 42.820 184.780 43.080 185.100 ;
        RECT 42.420 182.040 42.560 184.780 ;
        RECT 42.360 181.720 42.620 182.040 ;
        RECT 41.900 176.960 42.160 177.280 ;
        RECT 40.060 175.260 40.320 175.580 ;
        RECT 35.920 174.580 36.180 174.900 ;
        RECT 36.840 174.580 37.100 174.900 ;
        RECT 32.700 173.900 32.960 174.220 ;
        RECT 32.760 171.840 32.900 173.900 ;
        RECT 33.620 173.560 33.880 173.880 ;
        RECT 33.680 172.180 33.820 173.560 ;
        RECT 36.900 172.860 37.040 174.580 ;
        RECT 40.120 172.860 40.260 175.260 ;
        RECT 36.840 172.540 37.100 172.860 ;
        RECT 40.060 172.540 40.320 172.860 ;
        RECT 33.620 171.860 33.880 172.180 ;
        RECT 32.700 171.520 32.960 171.840 ;
        RECT 36.380 171.180 36.640 171.500 ;
        RECT 31.880 170.305 33.760 170.675 ;
        RECT 34.990 168.605 35.270 168.975 ;
        RECT 31.880 164.865 33.760 165.235 ;
        RECT 30.400 162.680 30.660 163.000 ;
        RECT 31.320 162.680 31.580 163.000 ;
        RECT 28.560 161.660 28.820 161.980 ;
        RECT 26.720 160.980 26.980 161.300 ;
        RECT 24.420 160.640 24.680 160.960 ;
        RECT 24.480 159.260 24.620 160.640 ;
        RECT 24.420 158.940 24.680 159.260 ;
        RECT 22.580 157.920 22.840 158.240 ;
        RECT 21.660 157.240 21.920 157.560 ;
        RECT 22.580 157.240 22.840 157.560 ;
        RECT 21.720 154.840 21.860 157.240 ;
        RECT 22.640 155.520 22.780 157.240 ;
        RECT 26.780 155.520 26.920 160.980 ;
        RECT 30.460 157.900 30.600 162.680 ;
        RECT 35.060 161.640 35.200 168.605 ;
        RECT 36.440 167.080 36.580 171.180 ;
        RECT 36.380 166.760 36.640 167.080 ;
        RECT 40.120 166.820 40.260 172.540 ;
        RECT 41.960 171.840 42.100 176.960 ;
        RECT 41.900 171.520 42.160 171.840 ;
        RECT 41.900 169.820 42.160 170.140 ;
        RECT 41.960 169.120 42.100 169.820 ;
        RECT 41.900 168.800 42.160 169.120 ;
        RECT 40.120 166.740 40.720 166.820 ;
        RECT 37.760 166.420 38.020 166.740 ;
        RECT 40.120 166.680 40.780 166.740 ;
        RECT 40.520 166.420 40.780 166.680 ;
        RECT 41.440 166.420 41.700 166.740 ;
        RECT 35.920 165.400 36.180 165.720 ;
        RECT 35.000 161.320 35.260 161.640 ;
        RECT 35.980 160.620 36.120 165.400 ;
        RECT 36.380 163.700 36.640 164.020 ;
        RECT 36.440 161.640 36.580 163.700 ;
        RECT 37.820 161.980 37.960 166.420 ;
        RECT 40.980 165.740 41.240 166.060 ;
        RECT 38.680 165.400 38.940 165.720 ;
        RECT 38.740 164.020 38.880 165.400 ;
        RECT 39.600 164.380 39.860 164.700 ;
        RECT 38.680 163.700 38.940 164.020 ;
        RECT 39.660 161.980 39.800 164.380 ;
        RECT 41.040 163.680 41.180 165.740 ;
        RECT 41.500 164.360 41.640 166.420 ;
        RECT 41.440 164.040 41.700 164.360 ;
        RECT 40.060 163.360 40.320 163.680 ;
        RECT 40.980 163.360 41.240 163.680 ;
        RECT 37.760 161.660 38.020 161.980 ;
        RECT 39.600 161.660 39.860 161.980 ;
        RECT 36.380 161.320 36.640 161.640 ;
        RECT 35.920 160.300 36.180 160.620 ;
        RECT 31.880 159.425 33.760 159.795 ;
        RECT 34.080 158.490 34.340 158.580 ;
        RECT 34.080 158.350 34.740 158.490 ;
        RECT 34.080 158.260 34.340 158.350 ;
        RECT 30.400 157.580 30.660 157.900 ;
        RECT 28.100 155.540 28.360 155.860 ;
        RECT 29.020 155.540 29.280 155.860 ;
        RECT 22.580 155.200 22.840 155.520 ;
        RECT 26.720 155.200 26.980 155.520 ;
        RECT 21.660 154.520 21.920 154.840 ;
        RECT 21.200 152.820 21.460 153.140 ;
        RECT 16.880 151.265 18.760 151.635 ;
        RECT 18.900 150.440 19.160 150.760 ;
        RECT 18.960 148.380 19.100 150.440 ;
        RECT 20.740 149.760 21.000 150.080 ;
        RECT 18.900 148.060 19.160 148.380 ;
        RECT 20.280 147.040 20.540 147.360 ;
        RECT 16.880 145.825 18.760 146.195 ;
        RECT 19.360 145.000 19.620 145.320 ;
        RECT 19.420 142.940 19.560 145.000 ;
        RECT 19.820 144.320 20.080 144.640 ;
        RECT 19.880 142.940 20.020 144.320 ;
        RECT 19.360 142.620 19.620 142.940 ;
        RECT 19.820 142.620 20.080 142.940 ;
        RECT 20.340 141.580 20.480 147.040 ;
        RECT 20.800 144.300 20.940 149.760 ;
        RECT 21.260 147.700 21.400 152.820 ;
        RECT 22.640 152.460 22.780 155.200 ;
        RECT 22.580 152.140 22.840 152.460 ;
        RECT 22.120 151.800 22.380 152.120 ;
        RECT 22.180 149.400 22.320 151.800 ;
        RECT 24.420 150.780 24.680 151.100 ;
        RECT 22.120 149.310 22.380 149.400 ;
        RECT 22.120 149.170 22.780 149.310 ;
        RECT 22.120 149.080 22.380 149.170 ;
        RECT 21.200 147.380 21.460 147.700 ;
        RECT 21.660 146.360 21.920 146.680 ;
        RECT 21.720 145.660 21.860 146.360 ;
        RECT 21.660 145.340 21.920 145.660 ;
        RECT 20.740 143.980 21.000 144.300 ;
        RECT 20.280 141.260 20.540 141.580 ;
        RECT 21.720 141.240 21.860 145.340 ;
        RECT 22.640 143.960 22.780 149.170 ;
        RECT 22.580 143.640 22.840 143.960 ;
        RECT 22.640 142.260 22.780 143.640 ;
        RECT 22.580 141.940 22.840 142.260 ;
        RECT 21.660 140.920 21.920 141.240 ;
        RECT 16.880 140.385 18.760 140.755 ;
        RECT 16.880 134.945 18.760 135.315 ;
        RECT 23.500 133.440 23.760 133.760 ;
        RECT 23.560 131.380 23.700 133.440 ;
        RECT 23.500 131.060 23.760 131.380 ;
        RECT 20.280 130.380 20.540 130.700 ;
        RECT 19.360 130.040 19.620 130.360 ;
        RECT 16.880 129.505 18.760 129.875 ;
        RECT 19.420 129.000 19.560 130.040 ;
        RECT 19.360 128.680 19.620 129.000 ;
        RECT 19.360 124.600 19.620 124.920 ;
        RECT 16.880 124.065 18.760 124.435 ;
        RECT 19.420 122.880 19.560 124.600 ;
        RECT 19.820 123.240 20.080 123.560 ;
        RECT 19.360 122.560 19.620 122.880 ;
        RECT 19.880 121.180 20.020 123.240 ;
        RECT 19.820 120.860 20.080 121.180 ;
        RECT 20.340 120.160 20.480 130.380 ;
        RECT 22.580 130.040 22.840 130.360 ;
        RECT 23.960 130.040 24.220 130.360 ;
        RECT 22.640 129.340 22.780 130.040 ;
        RECT 22.580 129.020 22.840 129.340 ;
        RECT 22.640 125.940 22.780 129.020 ;
        RECT 24.020 128.660 24.160 130.040 ;
        RECT 23.960 128.340 24.220 128.660 ;
        RECT 24.480 128.060 24.620 150.780 ;
        RECT 26.780 150.080 26.920 155.200 ;
        RECT 28.160 153.820 28.300 155.540 ;
        RECT 28.100 153.500 28.360 153.820 ;
        RECT 26.720 149.760 26.980 150.080 ;
        RECT 28.100 149.760 28.360 150.080 ;
        RECT 27.640 146.700 27.900 147.020 ;
        RECT 25.340 146.360 25.600 146.680 ;
        RECT 25.400 141.920 25.540 146.360 ;
        RECT 27.700 145.660 27.840 146.700 ;
        RECT 27.640 145.340 27.900 145.660 ;
        RECT 25.800 144.320 26.060 144.640 ;
        RECT 25.860 142.940 26.000 144.320 ;
        RECT 25.800 142.620 26.060 142.940 ;
        RECT 25.340 141.600 25.600 141.920 ;
        RECT 27.700 139.880 27.840 145.340 ;
        RECT 28.160 144.640 28.300 149.760 ;
        RECT 28.100 144.320 28.360 144.640 ;
        RECT 27.640 139.560 27.900 139.880 ;
        RECT 26.720 134.120 26.980 134.440 ;
        RECT 26.780 132.060 26.920 134.120 ;
        RECT 28.560 132.760 28.820 133.080 ;
        RECT 26.720 131.740 26.980 132.060 ;
        RECT 24.020 127.920 24.620 128.060 ;
        RECT 22.580 125.620 22.840 125.940 ;
        RECT 23.500 124.940 23.760 125.260 ;
        RECT 23.040 124.600 23.300 124.920 ;
        RECT 23.100 120.160 23.240 124.600 ;
        RECT 23.560 123.900 23.700 124.940 ;
        RECT 23.500 123.580 23.760 123.900 ;
        RECT 24.020 123.300 24.160 127.920 ;
        RECT 24.420 125.620 24.680 125.940 ;
        RECT 23.560 123.160 24.160 123.300 ;
        RECT 20.280 119.840 20.540 120.160 ;
        RECT 23.040 119.840 23.300 120.160 ;
        RECT 16.880 118.625 18.760 118.995 ;
        RECT 18.900 117.120 19.160 117.440 ;
        RECT 18.960 115.060 19.100 117.120 ;
        RECT 18.900 114.740 19.160 115.060 ;
        RECT 20.340 114.720 20.480 119.840 ;
        RECT 22.580 119.500 22.840 119.820 ;
        RECT 22.640 118.120 22.780 119.500 ;
        RECT 22.580 117.800 22.840 118.120 ;
        RECT 20.280 114.400 20.540 114.720 ;
        RECT 16.880 113.185 18.760 113.555 ;
        RECT 22.120 112.360 22.380 112.680 ;
        RECT 20.280 111.680 20.540 112.000 ;
        RECT 14.300 109.300 14.560 109.620 ;
        RECT 14.360 89.420 14.500 109.300 ;
        RECT 16.880 107.745 18.760 108.115 ;
        RECT 16.880 102.305 18.760 102.675 ;
        RECT 20.340 89.850 20.480 111.680 ;
        RECT 20.740 108.620 21.000 108.940 ;
        RECT 20.800 107.580 20.940 108.620 ;
        RECT 22.180 107.580 22.320 112.360 ;
        RECT 23.560 109.280 23.700 123.160 ;
        RECT 23.960 119.160 24.220 119.480 ;
        RECT 24.020 117.780 24.160 119.160 ;
        RECT 23.960 117.460 24.220 117.780 ;
        RECT 24.480 115.060 24.620 125.620 ;
        RECT 28.620 125.600 28.760 132.760 ;
        RECT 28.560 125.280 28.820 125.600 ;
        RECT 24.880 122.900 25.140 123.220 ;
        RECT 24.940 120.500 25.080 122.900 ;
        RECT 24.880 120.180 25.140 120.500 ;
        RECT 24.940 117.440 25.080 120.180 ;
        RECT 26.720 119.840 26.980 120.160 ;
        RECT 25.800 117.800 26.060 118.120 ;
        RECT 24.880 117.120 25.140 117.440 ;
        RECT 25.860 115.740 26.000 117.800 ;
        RECT 26.780 115.740 26.920 119.840 ;
        RECT 28.560 119.500 28.820 119.820 ;
        RECT 27.640 116.440 27.900 116.760 ;
        RECT 25.800 115.420 26.060 115.740 ;
        RECT 26.720 115.420 26.980 115.740 ;
        RECT 24.420 114.740 24.680 115.060 ;
        RECT 27.700 114.720 27.840 116.440 ;
        RECT 28.620 115.400 28.760 119.500 ;
        RECT 28.560 115.080 28.820 115.400 ;
        RECT 27.640 114.400 27.900 114.720 ;
        RECT 29.080 111.840 29.220 155.540 ;
        RECT 34.600 155.520 34.740 158.350 ;
        RECT 35.000 155.880 35.260 156.200 ;
        RECT 35.060 155.520 35.200 155.880 ;
        RECT 34.540 155.200 34.800 155.520 ;
        RECT 35.000 155.200 35.260 155.520 ;
        RECT 31.880 153.985 33.760 154.355 ;
        RECT 34.600 152.120 34.740 155.200 ;
        RECT 35.980 155.180 36.120 160.300 ;
        RECT 36.440 155.520 36.580 161.320 ;
        RECT 39.660 159.260 39.800 161.660 ;
        RECT 40.120 161.300 40.260 163.360 ;
        RECT 40.060 160.980 40.320 161.300 ;
        RECT 39.600 158.940 39.860 159.260 ;
        RECT 40.120 158.580 40.260 160.980 ;
        RECT 40.060 158.260 40.320 158.580 ;
        RECT 40.980 157.920 41.240 158.240 ;
        RECT 41.040 156.540 41.180 157.920 ;
        RECT 40.980 156.220 41.240 156.540 ;
        RECT 36.380 155.200 36.640 155.520 ;
        RECT 35.920 154.860 36.180 155.180 ;
        RECT 35.980 153.050 36.120 154.860 ;
        RECT 36.380 153.050 36.640 153.140 ;
        RECT 35.980 152.910 36.640 153.050 ;
        RECT 36.380 152.820 36.640 152.910 ;
        RECT 39.140 152.820 39.400 153.140 ;
        RECT 39.600 152.820 39.860 153.140 ;
        RECT 34.540 151.800 34.800 152.120 ;
        RECT 34.540 150.440 34.800 150.760 ;
        RECT 31.880 148.545 33.760 148.915 ;
        RECT 34.600 148.380 34.740 150.440 ;
        RECT 34.540 148.060 34.800 148.380 ;
        RECT 34.080 147.040 34.340 147.360 ;
        RECT 30.860 146.700 31.120 147.020 ;
        RECT 29.940 144.660 30.200 144.980 ;
        RECT 30.000 142.940 30.140 144.660 ;
        RECT 29.940 142.620 30.200 142.940 ;
        RECT 30.920 141.920 31.060 146.700 ;
        RECT 31.880 143.105 33.760 143.475 ;
        RECT 32.700 142.620 32.960 142.940 ;
        RECT 32.240 141.940 32.500 142.260 ;
        RECT 30.860 141.600 31.120 141.920 ;
        RECT 32.300 139.540 32.440 141.940 ;
        RECT 32.760 141.580 32.900 142.620 ;
        RECT 32.700 141.260 32.960 141.580 ;
        RECT 34.140 140.220 34.280 147.040 ;
        RECT 35.000 146.360 35.260 146.680 ;
        RECT 35.060 145.320 35.200 146.360 ;
        RECT 35.000 145.000 35.260 145.320 ;
        RECT 36.440 144.380 36.580 152.820 ;
        RECT 36.840 152.480 37.100 152.800 ;
        RECT 36.900 149.400 37.040 152.480 ;
        RECT 39.200 150.420 39.340 152.820 ;
        RECT 39.140 150.100 39.400 150.420 ;
        RECT 36.840 149.080 37.100 149.400 ;
        RECT 36.900 145.320 37.040 149.080 ;
        RECT 36.840 145.000 37.100 145.320 ;
        RECT 39.140 144.660 39.400 144.980 ;
        RECT 36.840 144.380 37.100 144.640 ;
        RECT 36.440 144.320 37.100 144.380 ;
        RECT 36.440 144.240 37.040 144.320 ;
        RECT 36.440 142.260 36.580 144.240 ;
        RECT 37.300 143.980 37.560 144.300 ;
        RECT 37.360 142.940 37.500 143.980 ;
        RECT 37.300 142.620 37.560 142.940 ;
        RECT 36.380 141.940 36.640 142.260 ;
        RECT 37.760 142.170 38.020 142.260 ;
        RECT 37.760 142.030 38.420 142.170 ;
        RECT 37.760 141.940 38.020 142.030 ;
        RECT 34.080 139.900 34.340 140.220 ;
        RECT 32.240 139.220 32.500 139.540 ;
        RECT 36.440 139.200 36.580 141.940 ;
        RECT 37.750 141.405 38.030 141.775 ;
        RECT 37.820 141.240 37.960 141.405 ;
        RECT 38.280 141.240 38.420 142.030 ;
        RECT 37.760 140.920 38.020 141.240 ;
        RECT 38.220 140.920 38.480 141.240 ;
        RECT 39.200 139.540 39.340 144.660 ;
        RECT 39.140 139.220 39.400 139.540 ;
        RECT 36.380 138.880 36.640 139.200 ;
        RECT 31.880 137.665 33.760 138.035 ;
        RECT 29.480 136.160 29.740 136.480 ;
        RECT 29.540 133.760 29.680 136.160 ;
        RECT 35.000 133.780 35.260 134.100 ;
        RECT 29.480 133.440 29.740 133.760 ;
        RECT 31.320 133.440 31.580 133.760 ;
        RECT 34.080 133.440 34.340 133.760 ;
        RECT 29.540 131.040 29.680 133.440 ;
        RECT 29.940 131.740 30.200 132.060 ;
        RECT 29.480 130.720 29.740 131.040 ;
        RECT 30.000 130.700 30.140 131.740 ;
        RECT 29.940 130.380 30.200 130.700 ;
        RECT 30.000 125.940 30.140 130.380 ;
        RECT 31.380 129.340 31.520 133.440 ;
        RECT 31.880 132.225 33.760 132.595 ;
        RECT 34.140 131.380 34.280 133.440 ;
        RECT 35.060 131.720 35.200 133.780 ;
        RECT 35.460 132.760 35.720 133.080 ;
        RECT 35.000 131.400 35.260 131.720 ;
        RECT 34.080 131.060 34.340 131.380 ;
        RECT 33.160 130.040 33.420 130.360 ;
        RECT 31.320 129.020 31.580 129.340 ;
        RECT 33.220 128.660 33.360 130.040 ;
        RECT 33.160 128.340 33.420 128.660 ;
        RECT 34.140 128.320 34.280 131.060 ;
        RECT 35.520 130.700 35.660 132.760 ;
        RECT 39.140 131.060 39.400 131.380 ;
        RECT 35.460 130.380 35.720 130.700 ;
        RECT 39.200 129.340 39.340 131.060 ;
        RECT 39.140 129.020 39.400 129.340 ;
        RECT 30.400 128.000 30.660 128.320 ;
        RECT 34.080 128.000 34.340 128.320 ;
        RECT 29.940 125.620 30.200 125.940 ;
        RECT 29.940 124.600 30.200 124.920 ;
        RECT 30.000 119.480 30.140 124.600 ;
        RECT 30.460 123.900 30.600 128.000 ;
        RECT 31.880 126.785 33.760 127.155 ;
        RECT 36.380 125.960 36.640 126.280 ;
        RECT 31.320 125.620 31.580 125.940 ;
        RECT 35.460 125.620 35.720 125.940 ;
        RECT 30.400 123.580 30.660 123.900 ;
        RECT 29.940 119.160 30.200 119.480 ;
        RECT 30.000 118.120 30.140 119.160 ;
        RECT 29.940 117.800 30.200 118.120 ;
        RECT 29.940 117.120 30.200 117.440 ;
        RECT 30.400 117.120 30.660 117.440 ;
        RECT 30.000 112.340 30.140 117.120 ;
        RECT 30.460 115.060 30.600 117.120 ;
        RECT 31.380 117.100 31.520 125.620 ;
        RECT 34.540 124.600 34.800 124.920 ;
        RECT 34.600 123.900 34.740 124.600 ;
        RECT 34.540 123.580 34.800 123.900 ;
        RECT 31.880 121.345 33.760 121.715 ;
        RECT 33.620 120.180 33.880 120.500 ;
        RECT 33.680 118.120 33.820 120.180 ;
        RECT 34.080 119.500 34.340 119.820 ;
        RECT 34.140 118.460 34.280 119.500 ;
        RECT 34.080 118.140 34.340 118.460 ;
        RECT 33.620 117.800 33.880 118.120 ;
        RECT 31.320 116.780 31.580 117.100 ;
        RECT 31.880 115.905 33.760 116.275 ;
        RECT 34.600 115.740 34.740 123.580 ;
        RECT 35.520 121.180 35.660 125.620 ;
        RECT 35.460 120.860 35.720 121.180 ;
        RECT 35.000 119.160 35.260 119.480 ;
        RECT 34.540 115.420 34.800 115.740 ;
        RECT 30.400 114.740 30.660 115.060 ;
        RECT 35.060 114.380 35.200 119.160 ;
        RECT 35.520 118.460 35.660 120.860 ;
        RECT 36.440 120.500 36.580 125.960 ;
        RECT 37.760 124.600 38.020 124.920 ;
        RECT 36.840 122.900 37.100 123.220 ;
        RECT 36.900 120.695 37.040 122.900 ;
        RECT 36.380 120.180 36.640 120.500 ;
        RECT 36.830 120.325 37.110 120.695 ;
        RECT 35.920 119.840 36.180 120.160 ;
        RECT 35.460 118.140 35.720 118.460 ;
        RECT 35.980 118.120 36.120 119.840 ;
        RECT 35.920 117.800 36.180 118.120 ;
        RECT 37.820 117.780 37.960 124.600 ;
        RECT 37.760 117.460 38.020 117.780 ;
        RECT 38.680 116.440 38.940 116.760 ;
        RECT 38.740 115.060 38.880 116.440 ;
        RECT 38.680 114.740 38.940 115.060 ;
        RECT 35.000 114.060 35.260 114.380 ;
        RECT 37.760 112.700 38.020 113.020 ;
        RECT 29.940 112.020 30.200 112.340 ;
        RECT 34.540 112.020 34.800 112.340 ;
        RECT 35.000 112.020 35.260 112.340 ;
        RECT 28.620 111.700 29.220 111.840 ;
        RECT 27.180 111.000 27.440 111.320 ;
        RECT 23.500 108.960 23.760 109.280 ;
        RECT 20.740 107.260 21.000 107.580 ;
        RECT 22.120 107.260 22.380 107.580 ;
        RECT 26.260 106.240 26.520 106.560 ;
        RECT 26.720 106.240 26.980 106.560 ;
        RECT 13.920 85.550 15.140 89.420 ;
        RECT 19.910 85.980 21.130 89.850 ;
        RECT 26.320 89.170 26.460 106.240 ;
        RECT 26.780 104.860 26.920 106.240 ;
        RECT 27.240 104.860 27.380 111.000 ;
        RECT 27.640 105.560 27.900 105.880 ;
        RECT 26.720 104.540 26.980 104.860 ;
        RECT 27.180 104.540 27.440 104.860 ;
        RECT 27.700 103.840 27.840 105.560 ;
        RECT 28.620 103.840 28.760 111.700 ;
        RECT 34.080 111.000 34.340 111.320 ;
        RECT 31.880 110.465 33.760 110.835 ;
        RECT 34.140 107.240 34.280 111.000 ;
        RECT 34.080 106.920 34.340 107.240 ;
        RECT 31.880 105.025 33.760 105.395 ;
        RECT 27.640 103.520 27.900 103.840 ;
        RECT 28.560 103.520 28.820 103.840 ;
        RECT 34.600 103.500 34.740 112.020 ;
        RECT 35.060 106.900 35.200 112.020 ;
        RECT 35.920 111.680 36.180 112.000 ;
        RECT 35.980 109.280 36.120 111.680 ;
        RECT 35.920 108.960 36.180 109.280 ;
        RECT 35.460 108.620 35.720 108.940 ;
        RECT 35.520 107.580 35.660 108.620 ;
        RECT 35.460 107.260 35.720 107.580 ;
        RECT 35.000 106.580 35.260 106.900 ;
        RECT 35.060 105.880 35.200 106.580 ;
        RECT 35.980 106.220 36.120 108.960 ;
        RECT 35.920 105.900 36.180 106.220 ;
        RECT 35.000 105.560 35.260 105.880 ;
        RECT 35.980 104.860 36.120 105.900 ;
        RECT 35.920 104.540 36.180 104.860 ;
        RECT 37.820 104.180 37.960 112.700 ;
        RECT 39.660 112.340 39.800 152.820 ;
        RECT 41.960 147.360 42.100 168.800 ;
        RECT 42.420 164.700 42.560 181.720 ;
        RECT 42.880 169.800 43.020 184.780 ;
        RECT 43.280 184.440 43.540 184.760 ;
        RECT 43.340 180.000 43.480 184.440 ;
        RECT 46.880 183.905 48.760 184.275 ;
        RECT 45.120 182.400 45.380 182.720 ;
        RECT 45.180 181.020 45.320 182.400 ;
        RECT 45.120 180.700 45.380 181.020 ;
        RECT 43.280 179.680 43.540 180.000 ;
        RECT 49.260 179.000 49.520 179.320 ;
        RECT 46.880 178.465 48.760 178.835 ;
        RECT 49.320 178.300 49.460 179.000 ;
        RECT 49.260 177.980 49.520 178.300 ;
        RECT 50.640 176.960 50.900 177.280 ;
        RECT 46.960 176.280 47.220 176.600 ;
        RECT 47.020 174.900 47.160 176.280 ;
        RECT 50.700 175.580 50.840 176.960 ;
        RECT 50.640 175.260 50.900 175.580 ;
        RECT 46.500 174.580 46.760 174.900 ;
        RECT 46.960 174.580 47.220 174.900 ;
        RECT 44.200 174.240 44.460 174.560 ;
        RECT 44.260 172.860 44.400 174.240 ;
        RECT 44.200 172.540 44.460 172.860 ;
        RECT 43.740 171.860 44.000 172.180 ;
        RECT 42.820 169.480 43.080 169.800 ;
        RECT 43.800 169.120 43.940 171.860 ;
        RECT 46.560 171.840 46.700 174.580 ;
        RECT 49.720 173.900 49.980 174.220 ;
        RECT 46.880 173.025 48.760 173.395 ;
        RECT 46.500 171.520 46.760 171.840 ;
        RECT 43.740 168.800 44.000 169.120 ;
        RECT 45.580 168.800 45.840 169.120 ;
        RECT 45.120 168.460 45.380 168.780 ;
        RECT 44.200 168.120 44.460 168.440 ;
        RECT 44.260 167.080 44.400 168.120 ;
        RECT 44.200 166.760 44.460 167.080 ;
        RECT 43.280 166.310 43.540 166.400 ;
        RECT 42.880 166.170 43.540 166.310 ;
        RECT 42.880 165.720 43.020 166.170 ;
        RECT 43.280 166.080 43.540 166.170 ;
        RECT 42.820 165.400 43.080 165.720 ;
        RECT 43.280 165.400 43.540 165.720 ;
        RECT 42.360 164.380 42.620 164.700 ;
        RECT 41.900 147.040 42.160 147.360 ;
        RECT 40.520 146.700 40.780 147.020 ;
        RECT 40.580 121.180 40.720 146.700 ;
        RECT 43.340 146.590 43.480 165.400 ;
        RECT 44.260 163.680 44.400 166.760 ;
        RECT 45.180 166.740 45.320 168.460 ;
        RECT 45.640 166.740 45.780 168.800 ;
        RECT 46.040 168.295 46.300 168.440 ;
        RECT 46.030 167.925 46.310 168.295 ;
        RECT 46.500 168.120 46.760 168.440 ;
        RECT 49.260 168.120 49.520 168.440 ;
        RECT 45.120 166.420 45.380 166.740 ;
        RECT 45.580 166.420 45.840 166.740 ;
        RECT 45.180 164.360 45.320 166.420 ;
        RECT 46.040 165.400 46.300 165.720 ;
        RECT 45.580 164.380 45.840 164.700 ;
        RECT 45.120 164.040 45.380 164.360 ;
        RECT 44.200 163.360 44.460 163.680 ;
        RECT 45.180 163.340 45.320 164.040 ;
        RECT 45.640 163.680 45.780 164.380 ;
        RECT 45.580 163.360 45.840 163.680 ;
        RECT 45.120 163.020 45.380 163.340 ;
        RECT 44.200 162.680 44.460 163.000 ;
        RECT 43.740 155.540 44.000 155.860 ;
        RECT 43.800 155.375 43.940 155.540 ;
        RECT 43.730 155.005 44.010 155.375 ;
        RECT 43.740 150.440 44.000 150.760 ;
        RECT 41.960 146.450 43.480 146.590 ;
        RECT 41.440 143.640 41.700 143.960 ;
        RECT 41.500 141.920 41.640 143.640 ;
        RECT 41.440 141.600 41.700 141.920 ;
        RECT 40.980 133.780 41.240 134.100 ;
        RECT 41.040 125.600 41.180 133.780 ;
        RECT 41.960 128.320 42.100 146.450 ;
        RECT 42.820 144.660 43.080 144.980 ;
        RECT 42.880 142.455 43.020 144.660 ;
        RECT 42.810 142.085 43.090 142.455 ;
        RECT 43.800 142.340 43.940 150.440 ;
        RECT 43.340 142.200 43.940 142.340 ;
        RECT 42.880 141.920 43.020 142.085 ;
        RECT 42.820 141.600 43.080 141.920 ;
        RECT 42.820 139.900 43.080 140.220 ;
        RECT 42.360 130.040 42.620 130.360 ;
        RECT 42.420 128.660 42.560 130.040 ;
        RECT 42.360 128.340 42.620 128.660 ;
        RECT 41.900 128.000 42.160 128.320 ;
        RECT 41.440 127.320 41.700 127.640 ;
        RECT 41.500 125.940 41.640 127.320 ;
        RECT 41.440 125.620 41.700 125.940 ;
        RECT 40.980 125.280 41.240 125.600 ;
        RECT 40.520 120.860 40.780 121.180 ;
        RECT 40.520 120.180 40.780 120.500 ;
        RECT 40.580 119.900 40.720 120.180 ;
        RECT 40.120 119.760 40.720 119.900 ;
        RECT 40.120 118.460 40.260 119.760 ;
        RECT 40.060 118.140 40.320 118.460 ;
        RECT 39.600 112.020 39.860 112.340 ;
        RECT 42.880 110.300 43.020 139.900 ;
        RECT 43.340 138.940 43.480 142.200 ;
        RECT 43.740 141.600 44.000 141.920 ;
        RECT 43.800 139.880 43.940 141.600 ;
        RECT 43.740 139.560 44.000 139.880 ;
        RECT 44.260 139.540 44.400 162.680 ;
        RECT 44.660 159.960 44.920 160.280 ;
        RECT 44.720 155.520 44.860 159.960 ;
        RECT 45.580 157.240 45.840 157.560 ;
        RECT 44.660 155.200 44.920 155.520 ;
        RECT 44.660 154.520 44.920 154.840 ;
        RECT 44.200 139.220 44.460 139.540 ;
        RECT 43.340 138.800 43.940 138.940 ;
        RECT 43.800 134.180 43.940 138.800 ;
        RECT 44.200 138.200 44.460 138.520 ;
        RECT 44.260 134.780 44.400 138.200 ;
        RECT 44.720 134.780 44.860 154.520 ;
        RECT 45.120 153.500 45.380 153.820 ;
        RECT 45.180 134.780 45.320 153.500 ;
        RECT 45.640 153.140 45.780 157.240 ;
        RECT 45.580 152.820 45.840 153.140 ;
        RECT 45.570 152.285 45.850 152.655 ;
        RECT 45.640 144.980 45.780 152.285 ;
        RECT 45.580 144.660 45.840 144.980 ;
        RECT 45.640 142.940 45.780 144.660 ;
        RECT 45.580 142.620 45.840 142.940 ;
        RECT 45.580 141.940 45.840 142.260 ;
        RECT 44.200 134.460 44.460 134.780 ;
        RECT 44.660 134.460 44.920 134.780 ;
        RECT 45.120 134.460 45.380 134.780 ;
        RECT 43.280 133.780 43.540 134.100 ;
        RECT 43.800 134.040 44.400 134.180 ;
        RECT 43.340 130.700 43.480 133.780 ;
        RECT 43.740 131.400 44.000 131.720 ;
        RECT 43.280 130.380 43.540 130.700 ;
        RECT 43.280 128.340 43.540 128.660 ;
        RECT 43.340 125.600 43.480 128.340 ;
        RECT 43.800 126.620 43.940 131.400 ;
        RECT 43.740 126.300 44.000 126.620 ;
        RECT 43.280 125.280 43.540 125.600 ;
        RECT 44.260 112.340 44.400 134.040 ;
        RECT 44.650 133.925 44.930 134.295 ;
        RECT 44.720 129.340 44.860 133.925 ;
        RECT 45.640 133.760 45.780 141.940 ;
        RECT 46.100 134.780 46.240 165.400 ;
        RECT 46.560 150.420 46.700 168.120 ;
        RECT 46.880 167.585 48.760 167.955 ;
        RECT 49.320 166.740 49.460 168.120 ;
        RECT 46.960 166.420 47.220 166.740 ;
        RECT 49.260 166.420 49.520 166.740 ;
        RECT 47.020 163.680 47.160 166.420 ;
        RECT 49.780 166.400 49.920 173.900 ;
        RECT 50.640 171.860 50.900 172.180 ;
        RECT 50.700 168.975 50.840 171.860 ;
        RECT 50.630 168.605 50.910 168.975 ;
        RECT 50.170 166.565 50.450 166.935 ;
        RECT 49.720 166.080 49.980 166.400 ;
        RECT 50.240 163.680 50.380 166.565 ;
        RECT 50.640 165.400 50.900 165.720 ;
        RECT 46.960 163.360 47.220 163.680 ;
        RECT 50.180 163.360 50.440 163.680 ;
        RECT 46.880 162.145 48.760 162.515 ;
        RECT 49.720 161.210 49.980 161.300 ;
        RECT 50.240 161.210 50.380 163.360 ;
        RECT 49.720 161.070 50.380 161.210 ;
        RECT 49.720 160.980 49.980 161.070 ;
        RECT 50.700 158.490 50.840 165.400 ;
        RECT 51.160 161.980 51.300 188.180 ;
        RECT 51.560 187.160 51.820 187.480 ;
        RECT 51.620 185.440 51.760 187.160 ;
        RECT 51.560 185.120 51.820 185.440 ;
        RECT 53.460 184.760 53.600 188.180 ;
        RECT 53.400 184.440 53.660 184.760 ;
        RECT 53.460 180.000 53.600 184.440 ;
        RECT 55.760 180.680 55.900 188.180 ;
        RECT 56.160 187.840 56.420 188.160 ;
        RECT 56.220 185.100 56.360 187.840 ;
        RECT 56.160 184.780 56.420 185.100 ;
        RECT 56.680 184.760 56.820 190.900 ;
        RECT 58.060 189.180 58.200 190.900 ;
        RECT 64.040 189.180 64.180 196.000 ;
        RECT 65.880 193.600 66.020 197.020 ;
        RECT 65.820 193.280 66.080 193.600 ;
        RECT 65.880 191.900 66.020 193.280 ;
        RECT 65.820 191.580 66.080 191.900 ;
        RECT 64.900 190.220 65.160 190.540 ;
        RECT 58.000 188.860 58.260 189.180 ;
        RECT 63.980 188.860 64.240 189.180 ;
        RECT 61.880 186.625 63.760 186.995 ;
        RECT 64.960 185.780 65.100 190.220 ;
        RECT 67.260 188.840 67.400 203.480 ;
        RECT 73.240 202.780 73.380 204.160 ;
        RECT 73.180 202.460 73.440 202.780 ;
        RECT 68.580 201.440 68.840 201.760 ;
        RECT 69.960 201.440 70.220 201.760 ;
        RECT 74.100 201.440 74.360 201.760 ;
        RECT 67.660 201.100 67.920 201.420 ;
        RECT 67.720 200.060 67.860 201.100 ;
        RECT 67.660 199.740 67.920 200.060 ;
        RECT 68.640 190.880 68.780 201.440 ;
        RECT 69.500 200.760 69.760 201.080 ;
        RECT 69.040 196.680 69.300 197.000 ;
        RECT 69.100 193.940 69.240 196.680 ;
        RECT 69.560 196.660 69.700 200.760 ;
        RECT 70.020 200.060 70.160 201.440 ;
        RECT 69.960 199.740 70.220 200.060 ;
        RECT 70.420 199.400 70.680 199.720 ;
        RECT 73.180 199.400 73.440 199.720 ;
        RECT 69.960 198.720 70.220 199.040 ;
        RECT 69.500 196.340 69.760 196.660 ;
        RECT 69.040 193.620 69.300 193.940 ;
        RECT 69.500 192.600 69.760 192.920 ;
        RECT 68.580 190.560 68.840 190.880 ;
        RECT 69.040 189.880 69.300 190.200 ;
        RECT 67.200 188.520 67.460 188.840 ;
        RECT 65.820 187.840 66.080 188.160 ;
        RECT 64.900 185.460 65.160 185.780 ;
        RECT 59.840 185.120 60.100 185.440 ;
        RECT 56.620 184.440 56.880 184.760 ;
        RECT 56.680 182.720 56.820 184.440 ;
        RECT 59.900 183.740 60.040 185.120 ;
        RECT 65.880 185.100 66.020 187.840 ;
        RECT 66.280 185.800 66.540 186.120 ;
        RECT 65.820 184.780 66.080 185.100 ;
        RECT 59.840 183.420 60.100 183.740 ;
        RECT 58.000 182.740 58.260 183.060 ;
        RECT 56.620 182.400 56.880 182.720 ;
        RECT 55.700 180.360 55.960 180.680 ;
        RECT 54.780 180.020 55.040 180.340 ;
        RECT 53.400 179.680 53.660 180.000 ;
        RECT 52.480 168.800 52.740 169.120 ;
        RECT 52.020 168.120 52.280 168.440 ;
        RECT 51.560 166.080 51.820 166.400 ;
        RECT 51.100 161.660 51.360 161.980 ;
        RECT 50.240 158.350 50.840 158.490 ;
        RECT 49.720 158.095 49.980 158.240 ;
        RECT 49.710 157.725 49.990 158.095 ;
        RECT 49.260 157.240 49.520 157.560 ;
        RECT 46.880 156.705 48.760 157.075 ;
        RECT 46.960 155.540 47.220 155.860 ;
        RECT 47.420 155.540 47.680 155.860 ;
        RECT 47.020 153.335 47.160 155.540 ;
        RECT 47.480 154.840 47.620 155.540 ;
        RECT 47.420 154.520 47.680 154.840 ;
        RECT 46.950 152.965 47.230 153.335 ;
        RECT 49.320 152.800 49.460 157.240 ;
        RECT 49.780 156.200 49.920 157.725 ;
        RECT 49.720 155.880 49.980 156.200 ;
        RECT 50.240 153.820 50.380 158.350 ;
        RECT 50.640 157.580 50.900 157.900 ;
        RECT 50.700 155.860 50.840 157.580 ;
        RECT 51.100 157.240 51.360 157.560 ;
        RECT 51.160 155.860 51.300 157.240 ;
        RECT 50.640 155.540 50.900 155.860 ;
        RECT 51.100 155.540 51.360 155.860 ;
        RECT 50.180 153.500 50.440 153.820 ;
        RECT 49.720 153.335 49.980 153.480 ;
        RECT 49.710 152.965 49.990 153.335 ;
        RECT 46.960 152.655 47.220 152.800 ;
        RECT 46.950 152.285 47.230 152.655 ;
        RECT 49.260 152.480 49.520 152.800 ;
        RECT 49.710 152.285 49.990 152.655 ;
        RECT 50.180 152.370 50.440 152.460 ;
        RECT 50.700 152.370 50.840 155.540 ;
        RECT 51.100 154.520 51.360 154.840 ;
        RECT 49.260 151.975 49.520 152.120 ;
        RECT 46.880 151.265 48.760 151.635 ;
        RECT 49.250 151.605 49.530 151.975 ;
        RECT 46.500 150.100 46.760 150.420 ;
        RECT 49.260 149.080 49.520 149.400 ;
        RECT 46.880 145.825 48.760 146.195 ;
        RECT 46.500 145.000 46.760 145.320 ;
        RECT 46.040 134.460 46.300 134.780 ;
        RECT 45.580 133.440 45.840 133.760 ;
        RECT 46.040 132.760 46.300 133.080 ;
        RECT 45.580 130.040 45.840 130.360 ;
        RECT 44.660 129.020 44.920 129.340 ;
        RECT 45.120 127.660 45.380 127.980 ;
        RECT 45.180 112.340 45.320 127.660 ;
        RECT 45.640 119.480 45.780 130.040 ;
        RECT 46.100 125.600 46.240 132.760 ;
        RECT 46.560 128.660 46.700 145.000 ;
        RECT 47.410 144.805 47.690 145.175 ;
        RECT 47.420 144.660 47.680 144.805 ;
        RECT 47.880 144.660 48.140 144.980 ;
        RECT 48.790 144.805 49.070 145.175 ;
        RECT 46.950 142.085 47.230 142.455 ;
        RECT 46.960 141.940 47.220 142.085 ;
        RECT 47.940 141.920 48.080 144.660 ;
        RECT 48.860 141.920 49.000 144.805 ;
        RECT 47.420 141.775 47.680 141.920 ;
        RECT 47.410 141.405 47.690 141.775 ;
        RECT 47.880 141.600 48.140 141.920 ;
        RECT 48.800 141.775 49.060 141.920 ;
        RECT 48.790 141.405 49.070 141.775 ;
        RECT 46.880 140.385 48.760 140.755 ;
        RECT 47.880 139.900 48.140 140.220 ;
        RECT 47.410 139.365 47.690 139.735 ;
        RECT 47.940 139.540 48.080 139.900 ;
        RECT 47.420 139.220 47.680 139.365 ;
        RECT 47.880 139.220 48.140 139.540 ;
        RECT 49.320 137.500 49.460 149.080 ;
        RECT 49.780 148.040 49.920 152.285 ;
        RECT 50.180 152.230 50.840 152.370 ;
        RECT 50.180 152.140 50.440 152.230 ;
        RECT 51.160 150.080 51.300 154.520 ;
        RECT 51.100 149.760 51.360 150.080 ;
        RECT 50.640 149.080 50.900 149.400 ;
        RECT 49.720 147.720 49.980 148.040 ;
        RECT 49.780 144.980 49.920 147.720 ;
        RECT 49.720 144.660 49.980 144.980 ;
        RECT 49.780 142.260 49.920 144.660 ;
        RECT 50.180 143.640 50.440 143.960 ;
        RECT 50.240 142.260 50.380 143.640 ;
        RECT 49.720 141.940 49.980 142.260 ;
        RECT 50.180 141.940 50.440 142.260 ;
        RECT 49.780 141.660 49.920 141.940 ;
        RECT 49.780 141.520 50.380 141.660 ;
        RECT 49.720 140.920 49.980 141.240 ;
        RECT 49.260 137.180 49.520 137.500 ;
        RECT 46.880 134.945 48.760 135.315 ;
        RECT 48.800 134.460 49.060 134.780 ;
        RECT 48.860 134.100 49.000 134.460 ;
        RECT 46.960 133.780 47.220 134.100 ;
        RECT 48.800 133.780 49.060 134.100 ;
        RECT 47.020 131.040 47.160 133.780 ;
        RECT 47.870 131.885 48.150 132.255 ;
        RECT 47.940 131.040 48.080 131.885 ;
        RECT 49.780 131.380 49.920 140.920 ;
        RECT 50.240 139.540 50.380 141.520 ;
        RECT 50.180 139.220 50.440 139.540 ;
        RECT 50.180 132.760 50.440 133.080 ;
        RECT 49.720 131.060 49.980 131.380 ;
        RECT 46.960 130.720 47.220 131.040 ;
        RECT 47.880 130.720 48.140 131.040 ;
        RECT 46.880 129.505 48.760 129.875 ;
        RECT 49.260 129.020 49.520 129.340 ;
        RECT 46.500 128.340 46.760 128.660 ;
        RECT 46.500 125.620 46.760 125.940 ;
        RECT 46.040 125.280 46.300 125.600 ;
        RECT 46.560 123.900 46.700 125.620 ;
        RECT 46.880 124.065 48.760 124.435 ;
        RECT 46.500 123.580 46.760 123.900 ;
        RECT 46.500 119.840 46.760 120.160 ;
        RECT 45.580 119.160 45.840 119.480 ;
        RECT 45.640 118.460 45.780 119.160 ;
        RECT 45.580 118.140 45.840 118.460 ;
        RECT 46.040 117.800 46.300 118.120 ;
        RECT 46.100 115.740 46.240 117.800 ;
        RECT 46.560 117.440 46.700 119.840 ;
        RECT 46.880 118.625 48.760 118.995 ;
        RECT 46.500 117.120 46.760 117.440 ;
        RECT 46.040 115.420 46.300 115.740 ;
        RECT 46.560 114.720 46.700 117.120 ;
        RECT 46.500 114.400 46.760 114.720 ;
        RECT 44.200 112.020 44.460 112.340 ;
        RECT 45.120 112.020 45.380 112.340 ;
        RECT 46.040 111.000 46.300 111.320 ;
        RECT 42.820 109.980 43.080 110.300 ;
        RECT 38.220 108.960 38.480 109.280 ;
        RECT 37.760 103.860 38.020 104.180 ;
        RECT 30.400 103.180 30.660 103.500 ;
        RECT 34.540 103.180 34.800 103.500 ;
        RECT 26.250 88.990 26.530 89.170 ;
        RECT 25.730 85.120 26.950 88.990 ;
        RECT 30.460 88.620 30.600 103.180 ;
        RECT 31.880 99.585 33.760 99.955 ;
        RECT 31.780 88.620 33.000 89.380 ;
        RECT 38.280 89.290 38.420 108.960 ;
        RECT 46.100 107.580 46.240 111.000 ;
        RECT 46.560 109.620 46.700 114.400 ;
        RECT 46.880 113.185 48.760 113.555 ;
        RECT 46.500 109.300 46.760 109.620 ;
        RECT 45.580 107.260 45.840 107.580 ;
        RECT 46.040 107.260 46.300 107.580 ;
        RECT 45.640 107.095 45.780 107.260 ;
        RECT 45.570 106.725 45.850 107.095 ;
        RECT 46.560 106.560 46.700 109.300 ;
        RECT 49.320 109.280 49.460 129.020 ;
        RECT 49.720 127.320 49.980 127.640 ;
        RECT 49.780 126.620 49.920 127.320 ;
        RECT 49.720 126.300 49.980 126.620 ;
        RECT 49.720 119.160 49.980 119.480 ;
        RECT 49.780 115.060 49.920 119.160 ;
        RECT 49.720 114.740 49.980 115.060 ;
        RECT 50.240 109.280 50.380 132.760 ;
        RECT 50.700 132.060 50.840 149.080 ;
        RECT 51.100 142.620 51.360 142.940 ;
        RECT 51.160 134.295 51.300 142.620 ;
        RECT 51.090 133.925 51.370 134.295 ;
        RECT 50.640 131.740 50.900 132.060 ;
        RECT 50.640 130.720 50.900 131.040 ;
        RECT 50.700 127.380 50.840 130.720 ;
        RECT 51.100 128.570 51.360 128.660 ;
        RECT 51.620 128.570 51.760 166.080 ;
        RECT 52.080 150.420 52.220 168.120 ;
        RECT 52.540 166.740 52.680 168.800 ;
        RECT 52.940 167.100 53.200 167.420 ;
        RECT 52.480 166.420 52.740 166.740 ;
        RECT 53.000 163.340 53.140 167.100 ;
        RECT 53.460 166.740 53.600 179.680 ;
        RECT 54.320 179.340 54.580 179.660 ;
        RECT 54.380 176.600 54.520 179.340 ;
        RECT 54.320 176.280 54.580 176.600 ;
        RECT 54.380 173.880 54.520 176.280 ;
        RECT 54.840 174.900 54.980 180.020 ;
        RECT 55.240 179.000 55.500 179.320 ;
        RECT 55.300 177.960 55.440 179.000 ;
        RECT 55.240 177.640 55.500 177.960 ;
        RECT 54.780 174.580 55.040 174.900 ;
        RECT 54.320 173.560 54.580 173.880 ;
        RECT 54.380 169.120 54.520 173.560 ;
        RECT 54.840 172.860 54.980 174.580 ;
        RECT 54.780 172.540 55.040 172.860 ;
        RECT 55.240 169.480 55.500 169.800 ;
        RECT 55.300 169.120 55.440 169.480 ;
        RECT 53.860 168.800 54.120 169.120 ;
        RECT 54.320 168.800 54.580 169.120 ;
        RECT 55.240 168.800 55.500 169.120 ;
        RECT 53.400 166.420 53.660 166.740 ;
        RECT 53.920 166.400 54.060 168.800 ;
        RECT 55.300 167.080 55.440 168.800 ;
        RECT 55.240 166.760 55.500 167.080 ;
        RECT 55.760 166.740 55.900 180.360 ;
        RECT 56.680 177.280 56.820 182.400 ;
        RECT 58.060 181.020 58.200 182.740 ;
        RECT 66.340 182.460 66.480 185.800 ;
        RECT 67.260 185.780 67.400 188.520 ;
        RECT 67.660 188.180 67.920 188.500 ;
        RECT 67.200 185.460 67.460 185.780 ;
        RECT 66.740 184.440 67.000 184.760 ;
        RECT 66.800 183.060 66.940 184.440 ;
        RECT 67.260 183.740 67.400 185.460 ;
        RECT 67.720 185.440 67.860 188.180 ;
        RECT 69.100 188.160 69.240 189.880 ;
        RECT 69.040 187.840 69.300 188.160 ;
        RECT 67.660 185.120 67.920 185.440 ;
        RECT 67.200 183.420 67.460 183.740 ;
        RECT 69.100 183.400 69.240 187.840 ;
        RECT 69.040 183.080 69.300 183.400 ;
        RECT 66.740 182.740 67.000 183.060 ;
        RECT 65.880 182.320 66.480 182.460 ;
        RECT 61.880 181.185 63.760 181.555 ;
        RECT 58.000 180.700 58.260 181.020 ;
        RECT 58.000 179.680 58.260 180.000 ;
        RECT 63.980 179.680 64.240 180.000 ;
        RECT 56.620 176.960 56.880 177.280 ;
        RECT 56.680 172.520 56.820 176.960 ;
        RECT 58.060 175.580 58.200 179.680 ;
        RECT 60.300 179.000 60.560 179.320 ;
        RECT 60.360 177.620 60.500 179.000 ;
        RECT 60.300 177.300 60.560 177.620 ;
        RECT 61.880 175.745 63.760 176.115 ;
        RECT 58.000 175.260 58.260 175.580 ;
        RECT 56.620 172.200 56.880 172.520 ;
        RECT 55.700 166.420 55.960 166.740 ;
        RECT 53.860 166.080 54.120 166.400 ;
        RECT 52.940 163.020 53.200 163.340 ;
        RECT 52.480 162.680 52.740 163.000 ;
        RECT 52.020 150.100 52.280 150.420 ;
        RECT 52.540 141.920 52.680 162.680 ;
        RECT 53.000 160.960 53.140 163.020 ;
        RECT 53.860 160.980 54.120 161.300 ;
        RECT 52.940 160.640 53.200 160.960 ;
        RECT 53.920 158.095 54.060 160.980 ;
        RECT 53.850 157.725 54.130 158.095 ;
        RECT 53.400 154.860 53.660 155.180 ;
        RECT 53.460 153.820 53.600 154.860 ;
        RECT 53.400 153.500 53.660 153.820 ;
        RECT 52.930 152.965 53.210 153.335 ;
        RECT 52.480 141.600 52.740 141.920 ;
        RECT 52.020 136.160 52.280 136.480 ;
        RECT 52.080 133.420 52.220 136.160 ;
        RECT 52.020 133.100 52.280 133.420 ;
        RECT 52.080 131.380 52.220 133.100 ;
        RECT 52.020 131.060 52.280 131.380 ;
        RECT 52.480 130.720 52.740 131.040 ;
        RECT 52.020 130.040 52.280 130.360 ;
        RECT 51.100 128.430 51.760 128.570 ;
        RECT 51.100 128.340 51.360 128.430 ;
        RECT 51.100 127.380 51.360 127.640 ;
        RECT 50.700 127.320 51.360 127.380 ;
        RECT 50.700 127.240 51.300 127.320 ;
        RECT 50.700 122.880 50.840 127.240 ;
        RECT 50.640 122.560 50.900 122.880 ;
        RECT 50.700 120.840 50.840 122.560 ;
        RECT 50.640 120.520 50.900 120.840 ;
        RECT 49.260 108.960 49.520 109.280 ;
        RECT 50.180 108.960 50.440 109.280 ;
        RECT 46.880 107.745 48.760 108.115 ;
        RECT 49.710 106.725 49.990 107.095 ;
        RECT 52.080 106.900 52.220 130.040 ;
        RECT 52.540 123.220 52.680 130.720 ;
        RECT 53.000 127.980 53.140 152.965 ;
        RECT 53.460 145.320 53.600 153.500 ;
        RECT 53.920 152.800 54.060 157.725 ;
        RECT 54.320 153.160 54.580 153.480 ;
        RECT 53.860 152.480 54.120 152.800 ;
        RECT 53.860 151.975 54.120 152.120 ;
        RECT 53.850 151.605 54.130 151.975 ;
        RECT 54.380 149.740 54.520 153.160 ;
        RECT 54.320 149.420 54.580 149.740 ;
        RECT 55.760 147.360 55.900 166.420 ;
        RECT 56.680 164.020 56.820 172.200 ;
        RECT 61.880 170.305 63.760 170.675 ;
        RECT 64.040 170.140 64.180 179.680 ;
        RECT 64.900 172.540 65.160 172.860 ;
        RECT 57.080 169.820 57.340 170.140 ;
        RECT 63.980 169.820 64.240 170.140 ;
        RECT 57.140 168.780 57.280 169.820 ;
        RECT 57.080 168.460 57.340 168.780 ;
        RECT 57.140 166.740 57.280 168.460 ;
        RECT 59.380 166.760 59.640 167.080 ;
        RECT 57.080 166.420 57.340 166.740 ;
        RECT 58.460 166.420 58.720 166.740 ;
        RECT 56.620 163.700 56.880 164.020 ;
        RECT 58.520 161.300 58.660 166.420 ;
        RECT 59.440 163.340 59.580 166.760 ;
        RECT 64.040 166.740 64.180 169.820 ;
        RECT 64.960 169.460 65.100 172.540 ;
        RECT 64.900 169.140 65.160 169.460 ;
        RECT 65.880 169.120 66.020 182.320 ;
        RECT 66.280 181.720 66.540 182.040 ;
        RECT 65.820 168.800 66.080 169.120 ;
        RECT 65.880 166.740 66.020 168.800 ;
        RECT 63.980 166.420 64.240 166.740 ;
        RECT 65.820 166.420 66.080 166.740 ;
        RECT 61.220 165.400 61.480 165.720 ;
        RECT 61.280 163.340 61.420 165.400 ;
        RECT 61.880 164.865 63.760 165.235 ;
        RECT 59.380 163.020 59.640 163.340 ;
        RECT 61.220 163.020 61.480 163.340 ;
        RECT 58.460 160.980 58.720 161.300 ;
        RECT 58.000 159.960 58.260 160.280 ;
        RECT 58.520 160.140 58.660 160.980 ;
        RECT 58.520 160.000 59.120 160.140 ;
        RECT 57.540 158.940 57.800 159.260 ;
        RECT 56.160 150.780 56.420 151.100 ;
        RECT 56.220 150.420 56.360 150.780 ;
        RECT 57.600 150.420 57.740 158.940 ;
        RECT 58.060 157.900 58.200 159.960 ;
        RECT 58.980 158.240 59.120 160.000 ;
        RECT 58.920 157.920 59.180 158.240 ;
        RECT 58.000 157.580 58.260 157.900 ;
        RECT 58.000 156.220 58.260 156.540 ;
        RECT 58.060 150.420 58.200 156.220 ;
        RECT 56.160 150.100 56.420 150.420 ;
        RECT 57.540 150.100 57.800 150.420 ;
        RECT 58.000 150.100 58.260 150.420 ;
        RECT 55.700 147.040 55.960 147.360 ;
        RECT 56.160 146.360 56.420 146.680 ;
        RECT 56.220 145.320 56.360 146.360 ;
        RECT 53.400 145.000 53.660 145.320 ;
        RECT 56.160 145.000 56.420 145.320 ;
        RECT 53.460 140.220 53.600 145.000 ;
        RECT 58.460 143.640 58.720 143.960 ;
        RECT 58.520 141.920 58.660 143.640 ;
        RECT 57.540 141.600 57.800 141.920 ;
        RECT 58.460 141.600 58.720 141.920 ;
        RECT 54.320 140.920 54.580 141.240 ;
        RECT 53.400 139.900 53.660 140.220 ;
        RECT 53.860 130.040 54.120 130.360 ;
        RECT 53.920 129.000 54.060 130.040 ;
        RECT 53.860 128.680 54.120 129.000 ;
        RECT 52.940 127.660 53.200 127.980 ;
        RECT 52.930 125.085 53.210 125.455 ;
        RECT 52.480 122.900 52.740 123.220 ;
        RECT 52.540 120.500 52.680 122.900 ;
        RECT 53.000 120.695 53.140 125.085 ;
        RECT 53.860 122.560 54.120 122.880 ;
        RECT 52.480 120.180 52.740 120.500 ;
        RECT 52.930 120.325 53.210 120.695 ;
        RECT 52.540 117.440 52.680 120.180 ;
        RECT 53.000 120.160 53.140 120.325 ;
        RECT 52.940 119.840 53.200 120.160 ;
        RECT 52.940 117.800 53.200 118.120 ;
        RECT 52.480 117.120 52.740 117.440 ;
        RECT 53.000 115.740 53.140 117.800 ;
        RECT 53.400 117.460 53.660 117.780 ;
        RECT 53.460 115.740 53.600 117.460 ;
        RECT 53.920 116.760 54.060 122.560 ;
        RECT 53.860 116.440 54.120 116.760 ;
        RECT 52.940 115.420 53.200 115.740 ;
        RECT 53.400 115.420 53.660 115.740 ;
        RECT 53.920 114.720 54.060 116.440 ;
        RECT 53.860 114.400 54.120 114.720 ;
        RECT 54.380 109.960 54.520 140.920 ;
        RECT 57.600 140.300 57.740 141.600 ;
        RECT 57.600 140.160 58.200 140.300 ;
        RECT 58.060 139.880 58.200 140.160 ;
        RECT 58.000 139.560 58.260 139.880 ;
        RECT 58.060 134.100 58.200 139.560 ;
        RECT 58.460 138.880 58.720 139.200 ;
        RECT 58.520 134.440 58.660 138.880 ;
        RECT 58.980 134.860 59.120 157.920 ;
        RECT 59.440 155.860 59.580 163.020 ;
        RECT 60.300 162.680 60.560 163.000 ;
        RECT 60.360 160.960 60.500 162.680 ;
        RECT 60.760 160.980 61.020 161.300 ;
        RECT 64.900 160.980 65.160 161.300 ;
        RECT 65.360 160.980 65.620 161.300 ;
        RECT 60.300 160.640 60.560 160.960 ;
        RECT 59.380 155.540 59.640 155.860 ;
        RECT 59.830 155.685 60.110 156.055 ;
        RECT 60.360 155.860 60.500 160.640 ;
        RECT 59.900 152.800 60.040 155.685 ;
        RECT 60.300 155.540 60.560 155.860 ;
        RECT 60.820 155.260 60.960 160.980 ;
        RECT 61.220 160.300 61.480 160.620 ;
        RECT 61.280 158.920 61.420 160.300 ;
        RECT 64.960 160.280 65.100 160.980 ;
        RECT 64.900 159.960 65.160 160.280 ;
        RECT 61.880 159.425 63.760 159.795 ;
        RECT 61.220 158.600 61.480 158.920 ;
        RECT 61.680 157.920 61.940 158.240 ;
        RECT 61.210 155.685 61.490 156.055 ;
        RECT 61.740 155.860 61.880 157.920 ;
        RECT 61.220 155.540 61.480 155.685 ;
        RECT 61.680 155.540 61.940 155.860 ;
        RECT 62.600 155.375 62.860 155.520 ;
        RECT 60.820 155.180 61.420 155.260 ;
        RECT 60.300 154.860 60.560 155.180 ;
        RECT 60.820 155.120 61.480 155.180 ;
        RECT 60.360 152.800 60.500 154.860 ;
        RECT 60.820 152.800 60.960 155.120 ;
        RECT 61.220 154.860 61.480 155.120 ;
        RECT 62.590 155.005 62.870 155.375 ;
        RECT 63.980 154.520 64.240 154.840 ;
        RECT 61.880 153.985 63.760 154.355 ;
        RECT 64.040 152.800 64.180 154.520 ;
        RECT 64.960 153.140 65.100 159.960 ;
        RECT 65.420 155.520 65.560 160.980 ;
        RECT 65.820 159.960 66.080 160.280 ;
        RECT 66.340 160.140 66.480 181.720 ;
        RECT 69.100 175.580 69.240 183.080 ;
        RECT 69.560 177.530 69.700 192.600 ;
        RECT 70.020 188.500 70.160 198.720 ;
        RECT 70.480 195.640 70.620 199.400 ;
        RECT 70.880 197.020 71.140 197.340 ;
        RECT 70.420 195.320 70.680 195.640 ;
        RECT 70.420 193.280 70.680 193.600 ;
        RECT 70.480 190.880 70.620 193.280 ;
        RECT 70.420 190.560 70.680 190.880 ;
        RECT 69.960 188.180 70.220 188.500 ;
        RECT 70.480 187.820 70.620 190.560 ;
        RECT 70.940 190.200 71.080 197.020 ;
        RECT 72.260 196.340 72.520 196.660 ;
        RECT 71.800 196.000 72.060 196.320 ;
        RECT 71.860 194.620 72.000 196.000 ;
        RECT 71.800 194.300 72.060 194.620 ;
        RECT 72.320 190.880 72.460 196.340 ;
        RECT 73.240 194.620 73.380 199.400 ;
        RECT 73.640 198.040 73.900 198.360 ;
        RECT 74.160 198.100 74.300 201.440 ;
        RECT 74.620 199.040 74.760 204.160 ;
        RECT 91.880 202.945 93.760 203.315 ;
        RECT 121.880 202.945 123.760 203.315 ;
        RECT 103.080 201.780 103.340 202.100 ;
        RECT 75.940 201.440 76.200 201.760 ;
        RECT 99.400 201.440 99.660 201.760 ;
        RECT 100.780 201.440 101.040 201.760 ;
        RECT 75.020 199.740 75.280 200.060 ;
        RECT 74.560 198.720 74.820 199.040 ;
        RECT 75.080 198.100 75.220 199.740 ;
        RECT 76.000 199.720 76.140 201.440 ;
        RECT 76.880 200.225 78.760 200.595 ;
        RECT 99.460 200.060 99.600 201.440 ;
        RECT 99.400 199.740 99.660 200.060 ;
        RECT 75.940 199.400 76.200 199.720 ;
        RECT 79.620 199.400 79.880 199.720 ;
        RECT 96.640 199.400 96.900 199.720 ;
        RECT 75.940 198.720 76.200 199.040 ;
        RECT 73.700 196.660 73.840 198.040 ;
        RECT 74.160 197.960 75.220 198.100 ;
        RECT 73.640 196.340 73.900 196.660 ;
        RECT 73.640 195.660 73.900 195.980 ;
        RECT 73.180 194.300 73.440 194.620 ;
        RECT 73.700 193.600 73.840 195.660 ;
        RECT 73.640 193.280 73.900 193.600 ;
        RECT 72.260 190.560 72.520 190.880 ;
        RECT 70.880 189.880 71.140 190.200 ;
        RECT 70.420 187.500 70.680 187.820 ;
        RECT 69.960 177.530 70.220 177.620 ;
        RECT 69.560 177.390 70.220 177.530 ;
        RECT 69.960 177.300 70.220 177.390 ;
        RECT 69.040 175.260 69.300 175.580 ;
        RECT 67.200 173.900 67.460 174.220 ;
        RECT 67.260 172.180 67.400 173.900 ;
        RECT 70.020 172.180 70.160 177.300 ;
        RECT 70.480 175.240 70.620 187.500 ;
        RECT 70.940 187.480 71.080 189.880 ;
        RECT 70.880 187.160 71.140 187.480 ;
        RECT 70.940 182.380 71.080 187.160 ;
        RECT 72.320 183.400 72.460 190.560 ;
        RECT 74.160 189.180 74.300 197.960 ;
        RECT 75.020 196.340 75.280 196.660 ;
        RECT 74.560 195.320 74.820 195.640 ;
        RECT 74.620 193.940 74.760 195.320 ;
        RECT 75.080 194.620 75.220 196.340 ;
        RECT 75.020 194.300 75.280 194.620 ;
        RECT 74.560 193.620 74.820 193.940 ;
        RECT 74.100 188.860 74.360 189.180 ;
        RECT 74.620 188.500 74.760 193.620 ;
        RECT 74.560 188.180 74.820 188.500 ;
        RECT 76.000 187.480 76.140 198.720 ;
        RECT 79.680 197.340 79.820 199.400 ;
        RECT 91.120 198.040 91.380 198.360 ;
        RECT 79.620 197.020 79.880 197.340 ;
        RECT 91.180 197.250 91.320 198.040 ;
        RECT 91.880 197.505 93.760 197.875 ;
        RECT 96.700 197.340 96.840 199.400 ;
        RECT 98.940 198.040 99.200 198.360 ;
        RECT 91.180 197.110 91.780 197.250 ;
        RECT 91.640 196.660 91.780 197.110 ;
        RECT 96.640 197.020 96.900 197.340 ;
        RECT 91.580 196.340 91.840 196.660 ;
        RECT 99.000 195.980 99.140 198.040 ;
        RECT 98.940 195.660 99.200 195.980 ;
        RECT 86.060 195.320 86.320 195.640 ;
        RECT 76.880 194.785 78.760 195.155 ;
        RECT 84.220 193.620 84.480 193.940 ;
        RECT 82.840 190.900 83.100 191.220 ;
        RECT 76.880 189.345 78.760 189.715 ;
        RECT 76.400 188.860 76.660 189.180 ;
        RECT 74.100 187.160 74.360 187.480 ;
        RECT 75.940 187.160 76.200 187.480 ;
        RECT 74.160 185.780 74.300 187.160 ;
        RECT 76.000 185.780 76.140 187.160 ;
        RECT 74.100 185.460 74.360 185.780 ;
        RECT 75.940 185.460 76.200 185.780 ;
        RECT 76.460 183.400 76.600 188.860 ;
        RECT 80.080 184.780 80.340 185.100 ;
        RECT 76.880 183.905 78.760 184.275 ;
        RECT 72.260 183.310 72.520 183.400 ;
        RECT 72.260 183.170 72.920 183.310 ;
        RECT 72.260 183.080 72.520 183.170 ;
        RECT 70.880 182.060 71.140 182.380 ;
        RECT 70.940 178.300 71.080 182.060 ;
        RECT 72.260 179.340 72.520 179.660 ;
        RECT 70.880 177.980 71.140 178.300 ;
        RECT 71.340 176.280 71.600 176.600 ;
        RECT 70.420 174.920 70.680 175.240 ;
        RECT 70.480 174.560 70.620 174.920 ;
        RECT 70.420 174.240 70.680 174.560 ;
        RECT 67.200 171.860 67.460 172.180 ;
        RECT 68.580 171.860 68.840 172.180 ;
        RECT 69.960 171.860 70.220 172.180 ;
        RECT 67.200 170.840 67.460 171.160 ;
        RECT 66.740 168.120 67.000 168.440 ;
        RECT 66.800 167.420 66.940 168.120 ;
        RECT 66.740 167.100 67.000 167.420 ;
        RECT 67.260 166.935 67.400 170.840 ;
        RECT 68.640 169.120 68.780 171.860 ;
        RECT 69.500 171.520 69.760 171.840 ;
        RECT 69.560 170.140 69.700 171.520 ;
        RECT 70.420 170.840 70.680 171.160 ;
        RECT 69.500 169.820 69.760 170.140 ;
        RECT 70.480 169.460 70.620 170.840 ;
        RECT 70.420 169.140 70.680 169.460 ;
        RECT 68.580 168.800 68.840 169.120 ;
        RECT 67.190 166.565 67.470 166.935 ;
        RECT 67.200 166.080 67.460 166.400 ;
        RECT 67.260 165.720 67.400 166.080 ;
        RECT 67.200 165.400 67.460 165.720 ;
        RECT 67.260 164.700 67.400 165.400 ;
        RECT 67.200 164.380 67.460 164.700 ;
        RECT 67.200 163.930 67.460 164.020 ;
        RECT 66.800 163.790 67.460 163.930 ;
        RECT 66.800 161.980 66.940 163.790 ;
        RECT 67.200 163.700 67.460 163.790 ;
        RECT 67.660 163.360 67.920 163.680 ;
        RECT 66.740 161.660 67.000 161.980 ;
        RECT 66.340 160.000 67.400 160.140 ;
        RECT 65.880 158.580 66.020 159.960 ;
        RECT 65.820 158.260 66.080 158.580 ;
        RECT 65.360 155.200 65.620 155.520 ;
        RECT 64.900 152.820 65.160 153.140 ;
        RECT 66.740 152.820 67.000 153.140 ;
        RECT 67.260 153.050 67.400 160.000 ;
        RECT 67.720 158.580 67.860 163.360 ;
        RECT 68.120 160.980 68.380 161.300 ;
        RECT 68.180 159.260 68.320 160.980 ;
        RECT 68.120 158.940 68.380 159.260 ;
        RECT 70.880 158.940 71.140 159.260 ;
        RECT 67.660 158.260 67.920 158.580 ;
        RECT 67.660 153.050 67.920 153.140 ;
        RECT 67.260 152.910 67.920 153.050 ;
        RECT 67.660 152.820 67.920 152.910 ;
        RECT 59.840 152.480 60.100 152.800 ;
        RECT 60.300 152.480 60.560 152.800 ;
        RECT 60.760 152.480 61.020 152.800 ;
        RECT 61.680 152.480 61.940 152.800 ;
        RECT 63.980 152.480 64.240 152.800 ;
        RECT 59.900 151.100 60.040 152.480 ;
        RECT 59.840 150.780 60.100 151.100 ;
        RECT 59.900 150.420 60.040 150.780 ;
        RECT 60.360 150.420 60.500 152.480 ;
        RECT 61.740 150.420 61.880 152.480 ;
        RECT 66.280 151.800 66.540 152.120 ;
        RECT 59.840 150.100 60.100 150.420 ;
        RECT 60.300 150.100 60.560 150.420 ;
        RECT 61.680 150.100 61.940 150.420 ;
        RECT 66.340 150.080 66.480 151.800 ;
        RECT 66.280 149.760 66.540 150.080 ;
        RECT 64.900 149.255 65.160 149.400 ;
        RECT 61.880 148.545 63.760 148.915 ;
        RECT 64.890 148.885 65.170 149.255 ;
        RECT 63.060 147.040 63.320 147.360 ;
        RECT 63.520 147.040 63.780 147.360 ;
        RECT 59.380 146.700 59.640 147.020 ;
        RECT 59.440 141.240 59.580 146.700 ;
        RECT 61.220 146.360 61.480 146.680 ;
        RECT 61.280 145.320 61.420 146.360 ;
        RECT 61.220 145.000 61.480 145.320 ;
        RECT 63.120 144.980 63.260 147.040 ;
        RECT 63.580 145.660 63.720 147.040 ;
        RECT 63.520 145.340 63.780 145.660 ;
        RECT 63.060 144.660 63.320 144.980 ;
        RECT 65.360 144.320 65.620 144.640 ;
        RECT 65.420 143.870 65.560 144.320 ;
        RECT 65.820 143.870 66.080 143.960 ;
        RECT 65.420 143.730 66.080 143.870 ;
        RECT 65.820 143.640 66.080 143.730 ;
        RECT 61.880 143.105 63.760 143.475 ;
        RECT 65.820 141.940 66.080 142.260 ;
        RECT 60.760 141.600 61.020 141.920 ;
        RECT 59.380 140.920 59.640 141.240 ;
        RECT 59.440 139.540 59.580 140.920 ;
        RECT 60.820 139.540 60.960 141.600 ;
        RECT 63.980 140.920 64.240 141.240 ;
        RECT 59.380 139.220 59.640 139.540 ;
        RECT 60.760 139.220 61.020 139.540 ;
        RECT 58.980 134.720 60.500 134.860 ;
        RECT 58.460 134.120 58.720 134.440 ;
        RECT 58.000 133.780 58.260 134.100 ;
        RECT 58.920 133.780 59.180 134.100 ;
        RECT 59.380 133.780 59.640 134.100 ;
        RECT 55.700 133.440 55.960 133.760 ;
        RECT 55.240 131.740 55.500 132.060 ;
        RECT 55.300 131.040 55.440 131.740 ;
        RECT 55.760 131.040 55.900 133.440 ;
        RECT 58.980 132.060 59.120 133.780 ;
        RECT 58.920 131.740 59.180 132.060 ;
        RECT 58.980 131.040 59.120 131.740 ;
        RECT 59.440 131.040 59.580 133.780 ;
        RECT 55.240 130.720 55.500 131.040 ;
        RECT 55.700 130.720 55.960 131.040 ;
        RECT 58.920 130.720 59.180 131.040 ;
        RECT 59.380 130.950 59.640 131.040 ;
        RECT 59.380 130.810 60.040 130.950 ;
        RECT 59.380 130.720 59.640 130.810 ;
        RECT 58.460 128.570 58.720 128.660 ;
        RECT 58.980 128.570 59.120 130.720 ;
        RECT 59.900 129.000 60.040 130.810 ;
        RECT 59.840 128.680 60.100 129.000 ;
        RECT 58.460 128.430 59.120 128.570 ;
        RECT 58.460 128.340 58.720 128.430 ;
        RECT 60.360 123.220 60.500 134.720 ;
        RECT 60.820 134.100 60.960 139.220 ;
        RECT 64.040 139.200 64.180 140.920 ;
        RECT 63.980 138.880 64.240 139.200 ;
        RECT 61.880 137.665 63.760 138.035 ;
        RECT 64.040 136.480 64.180 138.880 ;
        RECT 65.880 136.480 66.020 141.940 ;
        RECT 63.980 136.160 64.240 136.480 ;
        RECT 65.820 136.160 66.080 136.480 ;
        RECT 60.760 133.780 61.020 134.100 ;
        RECT 60.820 131.040 60.960 133.780 ;
        RECT 61.880 132.225 63.760 132.595 ;
        RECT 65.880 131.380 66.020 136.160 ;
        RECT 61.220 131.060 61.480 131.380 ;
        RECT 65.820 131.060 66.080 131.380 ;
        RECT 60.760 130.720 61.020 131.040 ;
        RECT 60.820 130.360 60.960 130.720 ;
        RECT 60.760 130.040 61.020 130.360 ;
        RECT 60.820 128.660 60.960 130.040 ;
        RECT 60.760 128.340 61.020 128.660 ;
        RECT 61.280 125.260 61.420 131.060 ;
        RECT 65.360 130.040 65.620 130.360 ;
        RECT 65.420 128.660 65.560 130.040 ;
        RECT 65.360 128.340 65.620 128.660 ;
        RECT 64.900 127.660 65.160 127.980 ;
        RECT 64.440 127.320 64.700 127.640 ;
        RECT 61.880 126.785 63.760 127.155 ;
        RECT 64.500 125.260 64.640 127.320 ;
        RECT 61.220 124.940 61.480 125.260 ;
        RECT 64.440 124.940 64.700 125.260 ;
        RECT 61.280 123.900 61.420 124.940 ;
        RECT 61.220 123.580 61.480 123.900 ;
        RECT 63.980 123.580 64.240 123.900 ;
        RECT 60.300 122.900 60.560 123.220 ;
        RECT 61.220 122.900 61.480 123.220 ;
        RECT 55.700 121.880 55.960 122.200 ;
        RECT 55.760 114.720 55.900 121.880 ;
        RECT 57.540 117.120 57.800 117.440 ;
        RECT 57.600 115.740 57.740 117.120 ;
        RECT 57.540 115.420 57.800 115.740 ;
        RECT 60.360 114.720 60.500 122.900 ;
        RECT 61.280 120.500 61.420 122.900 ;
        RECT 61.880 121.345 63.760 121.715 ;
        RECT 61.220 120.180 61.480 120.500 ;
        RECT 61.280 117.780 61.420 120.180 ;
        RECT 64.040 120.160 64.180 123.580 ;
        RECT 64.440 122.560 64.700 122.880 ;
        RECT 64.500 120.500 64.640 122.560 ;
        RECT 64.960 120.500 65.100 127.660 ;
        RECT 65.420 123.900 65.560 128.340 ;
        RECT 65.360 123.580 65.620 123.900 ;
        RECT 65.880 122.880 66.020 131.060 ;
        RECT 65.820 122.560 66.080 122.880 ;
        RECT 64.440 120.180 64.700 120.500 ;
        RECT 64.900 120.180 65.160 120.500 ;
        RECT 63.980 119.840 64.240 120.160 ;
        RECT 61.220 117.460 61.480 117.780 ;
        RECT 61.880 115.905 63.760 116.275 ;
        RECT 55.700 114.400 55.960 114.720 ;
        RECT 60.300 114.400 60.560 114.720 ;
        RECT 60.360 111.320 60.500 114.400 ;
        RECT 64.500 112.000 64.640 120.180 ;
        RECT 64.960 115.740 65.100 120.180 ;
        RECT 66.340 116.760 66.480 149.760 ;
        RECT 66.800 144.640 66.940 152.820 ;
        RECT 68.180 145.660 68.320 158.940 ;
        RECT 69.500 157.240 69.760 157.560 ;
        RECT 69.560 156.540 69.700 157.240 ;
        RECT 69.500 156.220 69.760 156.540 ;
        RECT 70.940 153.480 71.080 158.940 ;
        RECT 70.880 153.160 71.140 153.480 ;
        RECT 70.880 152.480 71.140 152.800 ;
        RECT 70.940 150.080 71.080 152.480 ;
        RECT 70.880 149.760 71.140 150.080 ;
        RECT 70.940 147.360 71.080 149.760 ;
        RECT 70.880 147.040 71.140 147.360 ;
        RECT 68.120 145.340 68.380 145.660 ;
        RECT 68.580 144.660 68.840 144.980 ;
        RECT 69.500 144.660 69.760 144.980 ;
        RECT 66.740 144.320 67.000 144.640 ;
        RECT 66.800 142.260 66.940 144.320 ;
        RECT 68.120 143.640 68.380 143.960 ;
        RECT 66.740 141.940 67.000 142.260 ;
        RECT 68.180 141.580 68.320 143.640 ;
        RECT 68.120 141.260 68.380 141.580 ;
        RECT 68.640 139.540 68.780 144.660 ;
        RECT 69.560 142.940 69.700 144.660 ;
        RECT 70.420 143.640 70.680 143.960 ;
        RECT 69.500 142.620 69.760 142.940 ;
        RECT 70.480 142.260 70.620 143.640 ;
        RECT 70.420 141.940 70.680 142.260 ;
        RECT 68.580 139.220 68.840 139.540 ;
        RECT 69.040 139.220 69.300 139.540 ;
        RECT 69.500 139.220 69.760 139.540 ;
        RECT 67.200 135.480 67.460 135.800 ;
        RECT 67.260 133.760 67.400 135.480 ;
        RECT 67.200 133.440 67.460 133.760 ;
        RECT 67.260 131.040 67.400 133.440 ;
        RECT 67.200 130.720 67.460 131.040 ;
        RECT 68.640 128.320 68.780 139.220 ;
        RECT 69.100 136.140 69.240 139.220 ;
        RECT 69.560 137.160 69.700 139.220 ;
        RECT 69.500 136.840 69.760 137.160 ;
        RECT 69.040 135.820 69.300 136.140 ;
        RECT 71.400 131.040 71.540 176.280 ;
        RECT 71.800 174.580 72.060 174.900 ;
        RECT 71.860 173.880 72.000 174.580 ;
        RECT 71.800 173.560 72.060 173.880 ;
        RECT 71.800 170.840 72.060 171.160 ;
        RECT 71.860 169.120 72.000 170.840 ;
        RECT 71.800 168.800 72.060 169.120 ;
        RECT 71.860 157.900 72.000 168.800 ;
        RECT 72.320 160.140 72.460 179.340 ;
        RECT 72.780 176.940 72.920 183.170 ;
        RECT 76.400 183.080 76.660 183.400 ;
        RECT 75.020 182.740 75.280 183.060 ;
        RECT 75.080 180.000 75.220 182.740 ;
        RECT 80.140 182.040 80.280 184.780 ;
        RECT 82.380 184.440 82.640 184.760 ;
        RECT 82.440 183.400 82.580 184.440 ;
        RECT 82.380 183.080 82.640 183.400 ;
        RECT 80.080 181.720 80.340 182.040 ;
        RECT 75.020 179.680 75.280 180.000 ;
        RECT 80.140 179.320 80.280 181.720 ;
        RECT 80.540 180.020 80.800 180.340 ;
        RECT 80.080 179.000 80.340 179.320 ;
        RECT 76.880 178.465 78.760 178.835 ;
        RECT 73.180 177.980 73.440 178.300 ;
        RECT 73.240 177.280 73.380 177.980 ;
        RECT 73.640 177.300 73.900 177.620 ;
        RECT 79.610 177.445 79.890 177.815 ;
        RECT 79.620 177.300 79.880 177.445 ;
        RECT 73.180 176.960 73.440 177.280 ;
        RECT 72.720 176.620 72.980 176.940 ;
        RECT 72.780 174.220 72.920 176.620 ;
        RECT 72.720 173.900 72.980 174.220 ;
        RECT 72.780 172.180 72.920 173.900 ;
        RECT 73.240 173.880 73.380 176.960 ;
        RECT 73.700 174.900 73.840 177.300 ;
        RECT 74.560 175.260 74.820 175.580 ;
        RECT 74.100 174.920 74.360 175.240 ;
        RECT 73.640 174.580 73.900 174.900 ;
        RECT 73.180 173.560 73.440 173.880 ;
        RECT 73.240 172.180 73.380 173.560 ;
        RECT 73.700 172.180 73.840 174.580 ;
        RECT 74.160 172.180 74.300 174.920 ;
        RECT 72.720 171.860 72.980 172.180 ;
        RECT 73.180 171.860 73.440 172.180 ;
        RECT 73.640 171.860 73.900 172.180 ;
        RECT 74.100 171.860 74.360 172.180 ;
        RECT 74.100 169.480 74.360 169.800 ;
        RECT 74.160 169.120 74.300 169.480 ;
        RECT 74.100 168.800 74.360 169.120 ;
        RECT 74.160 161.640 74.300 168.800 ;
        RECT 74.620 168.780 74.760 175.260 ;
        RECT 79.680 174.415 79.820 177.300 ;
        RECT 75.940 173.900 76.200 174.220 ;
        RECT 77.780 174.130 78.040 174.220 ;
        RECT 76.460 173.990 78.040 174.130 ;
        RECT 79.610 174.045 79.890 174.415 ;
        RECT 75.480 168.800 75.740 169.120 ;
        RECT 74.560 168.460 74.820 168.780 ;
        RECT 74.620 161.980 74.760 168.460 ;
        RECT 75.540 166.740 75.680 168.800 ;
        RECT 75.480 166.420 75.740 166.740 ;
        RECT 75.020 164.380 75.280 164.700 ;
        RECT 74.560 161.660 74.820 161.980 ;
        RECT 74.100 161.380 74.360 161.640 ;
        RECT 74.100 161.320 74.760 161.380 ;
        RECT 74.160 161.240 74.760 161.320 ;
        RECT 74.100 160.640 74.360 160.960 ;
        RECT 72.320 160.000 73.840 160.140 ;
        RECT 71.800 157.580 72.060 157.900 ;
        RECT 72.720 157.240 72.980 157.560 ;
        RECT 72.260 150.100 72.520 150.420 ;
        RECT 71.800 146.360 72.060 146.680 ;
        RECT 72.320 146.535 72.460 150.100 ;
        RECT 71.860 139.880 72.000 146.360 ;
        RECT 72.250 146.165 72.530 146.535 ;
        RECT 71.800 139.560 72.060 139.880 ;
        RECT 72.780 136.820 72.920 157.240 ;
        RECT 73.700 155.940 73.840 160.000 ;
        RECT 74.160 158.580 74.300 160.640 ;
        RECT 74.100 158.260 74.360 158.580 ;
        RECT 73.700 155.800 74.300 155.940 ;
        RECT 73.640 155.200 73.900 155.520 ;
        RECT 73.180 153.500 73.440 153.820 ;
        RECT 73.240 148.040 73.380 153.500 ;
        RECT 73.700 152.120 73.840 155.200 ;
        RECT 73.640 151.800 73.900 152.120 ;
        RECT 74.160 151.860 74.300 155.800 ;
        RECT 74.620 152.540 74.760 161.240 ;
        RECT 75.080 157.560 75.220 164.380 ;
        RECT 75.540 163.680 75.680 166.420 ;
        RECT 75.480 163.360 75.740 163.680 ;
        RECT 75.540 158.240 75.680 163.360 ;
        RECT 75.480 157.920 75.740 158.240 ;
        RECT 75.020 157.240 75.280 157.560 ;
        RECT 75.540 156.200 75.680 157.920 ;
        RECT 75.480 155.880 75.740 156.200 ;
        RECT 75.540 152.800 75.680 155.880 ;
        RECT 76.000 153.820 76.140 173.900 ;
        RECT 76.460 172.520 76.600 173.990 ;
        RECT 77.780 173.900 78.040 173.990 ;
        RECT 76.880 173.025 78.760 173.395 ;
        RECT 76.400 172.200 76.660 172.520 ;
        RECT 76.460 170.140 76.600 172.200 ;
        RECT 79.160 170.840 79.420 171.160 ;
        RECT 76.400 169.820 76.660 170.140 ;
        RECT 76.880 167.585 78.760 167.955 ;
        RECT 77.320 166.650 77.580 166.740 ;
        RECT 79.220 166.650 79.360 170.840 ;
        RECT 77.320 166.510 79.360 166.650 ;
        RECT 79.610 166.565 79.890 166.935 ;
        RECT 77.320 166.420 77.580 166.510 ;
        RECT 79.620 166.420 79.880 166.565 ;
        RECT 80.140 166.140 80.280 179.000 ;
        RECT 80.600 175.580 80.740 180.020 ;
        RECT 80.540 175.260 80.800 175.580 ;
        RECT 80.540 167.330 80.800 167.420 ;
        RECT 80.540 167.190 81.200 167.330 ;
        RECT 80.540 167.100 80.800 167.190 ;
        RECT 78.700 165.740 78.960 166.060 ;
        RECT 79.680 166.000 80.280 166.140 ;
        RECT 81.060 166.650 81.200 167.190 ;
        RECT 81.460 166.650 81.720 166.740 ;
        RECT 81.060 166.510 81.720 166.650 ;
        RECT 81.910 166.565 82.190 166.935 ;
        RECT 78.760 163.680 78.900 165.740 ;
        RECT 79.680 165.460 79.820 166.000 ;
        RECT 79.220 165.320 79.820 165.460 ;
        RECT 80.080 165.400 80.340 165.720 ;
        RECT 78.700 163.360 78.960 163.680 ;
        RECT 76.400 162.680 76.660 163.000 ;
        RECT 75.940 153.500 76.200 153.820 ;
        RECT 74.620 152.400 75.220 152.540 ;
        RECT 75.480 152.480 75.740 152.800 ;
        RECT 75.080 152.120 75.220 152.400 ;
        RECT 74.160 151.720 74.760 151.860 ;
        RECT 75.020 151.800 75.280 152.120 ;
        RECT 74.620 150.760 74.760 151.720 ;
        RECT 74.560 150.440 74.820 150.760 ;
        RECT 73.180 147.720 73.440 148.040 ;
        RECT 74.100 143.980 74.360 144.300 ;
        RECT 74.160 142.260 74.300 143.980 ;
        RECT 74.100 141.940 74.360 142.260 ;
        RECT 73.640 138.200 73.900 138.520 ;
        RECT 73.700 136.820 73.840 138.200 ;
        RECT 74.160 136.820 74.300 141.940 ;
        RECT 72.720 136.500 72.980 136.820 ;
        RECT 73.640 136.500 73.900 136.820 ;
        RECT 74.100 136.500 74.360 136.820 ;
        RECT 70.880 130.720 71.140 131.040 ;
        RECT 71.340 130.720 71.600 131.040 ;
        RECT 68.580 128.000 68.840 128.320 ;
        RECT 70.940 126.280 71.080 130.720 ;
        RECT 72.260 130.040 72.520 130.360 ;
        RECT 72.320 128.660 72.460 130.040 ;
        RECT 73.640 129.020 73.900 129.340 ;
        RECT 72.260 128.340 72.520 128.660 ;
        RECT 70.880 125.960 71.140 126.280 ;
        RECT 73.700 125.600 73.840 129.020 ;
        RECT 74.160 128.660 74.300 136.500 ;
        RECT 74.100 128.340 74.360 128.660 ;
        RECT 74.160 125.940 74.300 128.340 ;
        RECT 75.080 128.320 75.220 151.800 ;
        RECT 75.540 147.700 75.680 152.480 ;
        RECT 76.000 150.420 76.140 153.500 ;
        RECT 75.940 150.100 76.200 150.420 ;
        RECT 75.480 147.380 75.740 147.700 ;
        RECT 76.000 147.360 76.140 150.100 ;
        RECT 75.940 147.040 76.200 147.360 ;
        RECT 76.460 141.920 76.600 162.680 ;
        RECT 76.880 162.145 78.760 162.515 ;
        RECT 79.220 160.140 79.360 165.320 ;
        RECT 79.620 163.360 79.880 163.680 ;
        RECT 79.680 161.300 79.820 163.360 ;
        RECT 79.620 160.980 79.880 161.300 ;
        RECT 79.220 160.000 79.820 160.140 ;
        RECT 77.310 157.725 77.590 158.095 ;
        RECT 77.380 157.560 77.520 157.725 ;
        RECT 77.320 157.240 77.580 157.560 ;
        RECT 76.880 156.705 78.760 157.075 ;
        RECT 77.320 155.540 77.580 155.860 ;
        RECT 77.380 152.800 77.520 155.540 ;
        RECT 79.160 153.160 79.420 153.480 ;
        RECT 77.780 152.820 78.040 153.140 ;
        RECT 77.320 152.480 77.580 152.800 ;
        RECT 77.840 152.120 77.980 152.820 ;
        RECT 77.780 151.800 78.040 152.120 ;
        RECT 76.880 151.265 78.760 151.635 ;
        RECT 79.220 150.760 79.360 153.160 ;
        RECT 79.160 150.440 79.420 150.760 ;
        RECT 77.320 150.100 77.580 150.420 ;
        RECT 76.860 149.255 77.120 149.400 ;
        RECT 76.850 148.885 77.130 149.255 ;
        RECT 77.380 147.700 77.520 150.100 ;
        RECT 78.700 149.420 78.960 149.740 ;
        RECT 77.320 147.380 77.580 147.700 ;
        RECT 78.760 146.680 78.900 149.420 ;
        RECT 79.220 147.700 79.360 150.440 ;
        RECT 79.160 147.380 79.420 147.700 ;
        RECT 78.700 146.360 78.960 146.680 ;
        RECT 76.880 145.825 78.760 146.195 ;
        RECT 79.220 145.320 79.360 147.380 ;
        RECT 79.680 147.360 79.820 160.000 ;
        RECT 79.620 147.040 79.880 147.360 ;
        RECT 79.160 145.000 79.420 145.320 ;
        RECT 78.240 143.640 78.500 143.960 ;
        RECT 78.300 142.260 78.440 143.640 ;
        RECT 78.700 142.850 78.960 142.940 ;
        RECT 78.700 142.710 79.360 142.850 ;
        RECT 78.700 142.620 78.960 142.710 ;
        RECT 78.240 141.940 78.500 142.260 ;
        RECT 76.400 141.600 76.660 141.920 ;
        RECT 75.940 140.920 76.200 141.240 ;
        RECT 75.480 130.720 75.740 131.040 ;
        RECT 75.540 128.660 75.680 130.720 ;
        RECT 75.480 128.340 75.740 128.660 ;
        RECT 75.020 128.000 75.280 128.320 ;
        RECT 74.100 125.620 74.360 125.940 ;
        RECT 71.340 125.280 71.600 125.600 ;
        RECT 71.800 125.280 72.060 125.600 ;
        RECT 73.640 125.280 73.900 125.600 ;
        RECT 71.400 123.220 71.540 125.280 ;
        RECT 71.860 123.900 72.000 125.280 ;
        RECT 71.800 123.580 72.060 123.900 ;
        RECT 71.340 122.900 71.600 123.220 ;
        RECT 69.040 119.160 69.300 119.480 ;
        RECT 66.280 116.440 66.540 116.760 ;
        RECT 64.900 115.420 65.160 115.740 ;
        RECT 64.960 112.680 65.100 115.420 ;
        RECT 66.340 113.020 66.480 116.440 ;
        RECT 69.100 115.060 69.240 119.160 ;
        RECT 69.960 117.800 70.220 118.120 ;
        RECT 70.020 115.740 70.160 117.800 ;
        RECT 74.160 117.780 74.300 125.620 ;
        RECT 75.480 124.940 75.740 125.260 ;
        RECT 75.540 122.880 75.680 124.940 ;
        RECT 75.480 122.560 75.740 122.880 ;
        RECT 74.100 117.460 74.360 117.780 ;
        RECT 71.800 117.120 72.060 117.440 ;
        RECT 69.960 115.420 70.220 115.740 ;
        RECT 69.040 114.740 69.300 115.060 ;
        RECT 71.860 113.020 72.000 117.120 ;
        RECT 74.160 115.060 74.300 117.460 ;
        RECT 74.100 114.740 74.360 115.060 ;
        RECT 73.180 114.400 73.440 114.720 ;
        RECT 66.280 112.700 66.540 113.020 ;
        RECT 71.800 112.700 72.060 113.020 ;
        RECT 64.900 112.360 65.160 112.680 ;
        RECT 64.440 111.680 64.700 112.000 ;
        RECT 73.240 111.320 73.380 114.400 ;
        RECT 60.300 111.000 60.560 111.320 ;
        RECT 73.180 111.000 73.440 111.320 ;
        RECT 54.320 109.640 54.580 109.960 ;
        RECT 60.360 109.280 60.500 111.000 ;
        RECT 61.880 110.465 63.760 110.835 ;
        RECT 60.300 108.960 60.560 109.280 ;
        RECT 59.840 108.620 60.100 108.940 ;
        RECT 56.620 106.920 56.880 107.240 ;
        RECT 49.720 106.580 49.980 106.725 ;
        RECT 52.020 106.580 52.280 106.900 ;
        RECT 44.200 106.240 44.460 106.560 ;
        RECT 46.500 106.240 46.760 106.560 ;
        RECT 40.980 105.560 41.240 105.880 ;
        RECT 41.040 104.180 41.180 105.560 ;
        RECT 40.980 103.860 41.240 104.180 ;
        RECT 44.260 89.530 44.400 106.240 ;
        RECT 46.560 104.860 46.700 106.240 ;
        RECT 49.260 105.560 49.520 105.880 ;
        RECT 46.500 104.540 46.760 104.860 ;
        RECT 49.320 103.500 49.460 105.560 ;
        RECT 49.780 104.180 49.920 106.580 ;
        RECT 54.320 106.240 54.580 106.560 ;
        RECT 49.720 103.860 49.980 104.180 ;
        RECT 49.260 103.180 49.520 103.500 ;
        RECT 49.720 103.180 49.980 103.500 ;
        RECT 46.880 102.305 48.760 102.675 ;
        RECT 37.750 88.780 38.970 89.290 ;
        RECT 30.460 88.480 33.000 88.620 ;
        RECT 31.780 85.510 33.000 88.480 ;
        RECT 37.680 88.620 38.970 88.780 ;
        RECT 43.810 88.630 45.030 89.530 ;
        RECT 49.780 89.040 49.920 103.180 ;
        RECT 50.170 89.040 50.450 89.170 ;
        RECT 49.740 88.640 50.960 89.040 ;
        RECT 37.680 86.810 39.070 88.620 ;
        RECT 37.750 85.420 38.970 86.810 ;
        RECT 43.810 86.720 45.140 88.630 ;
        RECT 49.740 86.920 51.010 88.640 ;
        RECT 54.380 88.620 54.520 106.240 ;
        RECT 56.680 104.860 56.820 106.920 ;
        RECT 56.620 104.540 56.880 104.860 ;
        RECT 59.900 103.840 60.040 108.620 ;
        RECT 60.300 108.280 60.560 108.600 ;
        RECT 67.200 108.280 67.460 108.600 ;
        RECT 72.260 108.280 72.520 108.600 ;
        RECT 60.360 107.240 60.500 108.280 ;
        RECT 60.300 106.920 60.560 107.240 ;
        RECT 64.900 106.920 65.160 107.240 ;
        RECT 63.980 106.240 64.240 106.560 ;
        RECT 61.880 105.025 63.760 105.395 ;
        RECT 64.040 104.940 64.180 106.240 ;
        RECT 64.040 104.860 64.640 104.940 ;
        RECT 64.040 104.800 64.700 104.860 ;
        RECT 64.440 104.540 64.700 104.800 ;
        RECT 59.840 103.520 60.100 103.840 ;
        RECT 59.900 101.460 60.040 103.520 ;
        RECT 60.760 103.180 61.020 103.500 ;
        RECT 62.140 103.180 62.400 103.500 ;
        RECT 59.840 101.140 60.100 101.460 ;
        RECT 55.530 88.620 56.750 89.190 ;
        RECT 54.380 88.480 56.750 88.620 ;
        RECT 60.820 88.620 60.960 103.180 ;
        RECT 62.200 102.140 62.340 103.180 ;
        RECT 64.960 102.140 65.100 106.920 ;
        RECT 67.260 104.180 67.400 108.280 ;
        RECT 68.120 107.260 68.380 107.580 ;
        RECT 67.200 103.860 67.460 104.180 ;
        RECT 62.140 101.820 62.400 102.140 ;
        RECT 64.900 101.820 65.160 102.140 ;
        RECT 61.880 99.585 63.760 99.955 ;
        RECT 68.180 89.840 68.320 107.260 ;
        RECT 72.320 107.240 72.460 108.280 ;
        RECT 72.260 106.920 72.520 107.240 ;
        RECT 74.160 106.900 74.300 114.740 ;
        RECT 76.000 109.620 76.140 140.920 ;
        RECT 76.880 140.385 78.760 140.755 ;
        RECT 76.880 134.945 78.760 135.315 ;
        RECT 76.880 129.505 78.760 129.875 ;
        RECT 76.400 128.000 76.660 128.320 ;
        RECT 76.460 110.300 76.600 128.000 ;
        RECT 79.220 124.920 79.360 142.710 ;
        RECT 80.140 141.920 80.280 165.400 ;
        RECT 81.060 163.680 81.200 166.510 ;
        RECT 81.460 166.420 81.720 166.510 ;
        RECT 81.920 166.420 82.180 166.565 ;
        RECT 80.540 163.360 80.800 163.680 ;
        RECT 81.000 163.360 81.260 163.680 ;
        RECT 80.600 161.210 80.740 163.360 ;
        RECT 81.060 161.980 81.200 163.360 ;
        RECT 81.000 161.660 81.260 161.980 ;
        RECT 81.980 161.300 82.120 166.420 ;
        RECT 81.920 161.210 82.180 161.300 ;
        RECT 80.600 161.070 82.180 161.210 ;
        RECT 81.920 160.980 82.180 161.070 ;
        RECT 82.900 160.140 83.040 190.900 ;
        RECT 83.300 190.560 83.560 190.880 ;
        RECT 83.360 185.440 83.500 190.560 ;
        RECT 83.760 189.880 84.020 190.200 ;
        RECT 83.820 188.840 83.960 189.880 ;
        RECT 83.760 188.520 84.020 188.840 ;
        RECT 84.280 188.160 84.420 193.620 ;
        RECT 86.120 193.600 86.260 195.320 ;
        RECT 99.460 193.940 99.600 199.740 ;
        RECT 100.840 199.720 100.980 201.440 ;
        RECT 100.780 199.400 101.040 199.720 ;
        RECT 103.140 194.280 103.280 201.780 ;
        RECT 112.740 201.670 113.000 201.760 ;
        RECT 112.340 201.530 113.000 201.670 ;
        RECT 109.060 201.100 109.320 201.420 ;
        RECT 111.360 201.100 111.620 201.420 ;
        RECT 106.880 200.225 108.760 200.595 ;
        RECT 109.120 200.060 109.260 201.100 ;
        RECT 109.060 199.740 109.320 200.060 ;
        RECT 108.600 199.060 108.860 199.380 ;
        RECT 108.660 197.340 108.800 199.060 ;
        RECT 111.420 197.340 111.560 201.100 ;
        RECT 112.340 199.040 112.480 201.530 ;
        RECT 112.740 201.440 113.000 201.530 ;
        RECT 112.280 198.720 112.540 199.040 ;
        RECT 108.600 197.020 108.860 197.340 ;
        RECT 111.360 197.020 111.620 197.340 ;
        RECT 105.380 196.340 105.640 196.660 ;
        RECT 104.920 195.660 105.180 195.980 ;
        RECT 103.080 193.960 103.340 194.280 ;
        RECT 99.400 193.620 99.660 193.940 ;
        RECT 102.620 193.620 102.880 193.940 ;
        RECT 85.140 193.280 85.400 193.600 ;
        RECT 86.060 193.280 86.320 193.600 ;
        RECT 84.220 187.840 84.480 188.160 ;
        RECT 83.300 185.120 83.560 185.440 ;
        RECT 83.360 180.000 83.500 185.120 ;
        RECT 84.280 184.760 84.420 187.840 ;
        RECT 85.200 185.780 85.340 193.280 ;
        RECT 86.120 191.220 86.260 193.280 ;
        RECT 90.660 192.600 90.920 192.920 ;
        RECT 90.720 191.220 90.860 192.600 ;
        RECT 91.880 192.065 93.760 192.435 ;
        RECT 86.060 190.900 86.320 191.220 ;
        RECT 90.660 190.900 90.920 191.220 ;
        RECT 93.420 190.560 93.680 190.880 ;
        RECT 90.200 188.180 90.460 188.500 ;
        RECT 87.440 187.160 87.700 187.480 ;
        RECT 85.140 185.460 85.400 185.780 ;
        RECT 84.220 184.615 84.480 184.760 ;
        RECT 84.210 184.245 84.490 184.615 ;
        RECT 85.200 180.340 85.340 185.460 ;
        RECT 86.520 183.080 86.780 183.400 ;
        RECT 85.140 180.020 85.400 180.340 ;
        RECT 83.300 179.680 83.560 180.000 ;
        RECT 83.360 174.900 83.500 179.680 ;
        RECT 83.760 179.000 84.020 179.320 ;
        RECT 84.220 179.000 84.480 179.320 ;
        RECT 83.300 174.580 83.560 174.900 ;
        RECT 83.820 174.560 83.960 179.000 ;
        RECT 84.280 178.300 84.420 179.000 ;
        RECT 84.220 177.980 84.480 178.300 ;
        RECT 85.200 177.280 85.340 180.020 ;
        RECT 85.140 176.960 85.400 177.280 ;
        RECT 86.580 175.580 86.720 183.080 ;
        RECT 87.500 183.060 87.640 187.160 ;
        RECT 90.260 186.460 90.400 188.180 ;
        RECT 93.480 188.160 93.620 190.560 ;
        RECT 93.420 187.840 93.680 188.160 ;
        RECT 99.400 187.160 99.660 187.480 ;
        RECT 91.880 186.625 93.760 186.995 ;
        RECT 90.200 186.140 90.460 186.460 ;
        RECT 99.460 185.440 99.600 187.160 ;
        RECT 99.400 185.120 99.660 185.440 ;
        RECT 102.160 185.120 102.420 185.440 ;
        RECT 99.860 184.440 100.120 184.760 ;
        RECT 87.440 182.740 87.700 183.060 ;
        RECT 90.660 182.740 90.920 183.060 ;
        RECT 87.500 179.320 87.640 182.740 ;
        RECT 87.900 179.340 88.160 179.660 ;
        RECT 87.440 179.000 87.700 179.320 ;
        RECT 87.500 177.960 87.640 179.000 ;
        RECT 87.440 177.640 87.700 177.960 ;
        RECT 87.960 175.580 88.100 179.340 ;
        RECT 90.720 178.300 90.860 182.740 ;
        RECT 99.920 182.040 100.060 184.440 ;
        RECT 100.320 183.420 100.580 183.740 ;
        RECT 100.380 182.040 100.520 183.420 ;
        RECT 101.240 183.080 101.500 183.400 ;
        RECT 100.780 182.400 101.040 182.720 ;
        RECT 91.120 181.720 91.380 182.040 ;
        RECT 99.860 181.720 100.120 182.040 ;
        RECT 100.320 181.720 100.580 182.040 ;
        RECT 91.180 180.340 91.320 181.720 ;
        RECT 91.880 181.185 93.760 181.555 ;
        RECT 91.120 180.020 91.380 180.340 ;
        RECT 91.120 179.000 91.380 179.320 ;
        RECT 90.660 177.980 90.920 178.300 ;
        RECT 86.520 175.260 86.780 175.580 ;
        RECT 87.900 175.260 88.160 175.580 ;
        RECT 91.180 174.560 91.320 179.000 ;
        RECT 99.920 177.620 100.060 181.720 ;
        RECT 100.380 177.620 100.520 181.720 ;
        RECT 100.840 180.000 100.980 182.400 ;
        RECT 100.780 179.680 101.040 180.000 ;
        RECT 99.860 177.300 100.120 177.620 ;
        RECT 100.320 177.300 100.580 177.620 ;
        RECT 99.400 176.280 99.660 176.600 ;
        RECT 91.880 175.745 93.760 176.115 ;
        RECT 99.460 174.560 99.600 176.280 ;
        RECT 83.760 174.240 84.020 174.560 ;
        RECT 91.120 174.240 91.380 174.560 ;
        RECT 99.400 174.240 99.660 174.560 ;
        RECT 84.680 172.200 84.940 172.520 ;
        RECT 84.220 170.840 84.480 171.160 ;
        RECT 84.280 169.120 84.420 170.840 ;
        RECT 84.740 170.140 84.880 172.200 ;
        RECT 91.180 172.180 91.320 174.240 ;
        RECT 94.340 173.900 94.600 174.220 ;
        RECT 94.400 172.520 94.540 173.900 ;
        RECT 98.020 172.540 98.280 172.860 ;
        RECT 94.340 172.200 94.600 172.520 ;
        RECT 91.120 171.860 91.380 172.180 ;
        RECT 93.880 171.860 94.140 172.180 ;
        RECT 85.140 171.520 85.400 171.840 ;
        RECT 89.280 171.520 89.540 171.840 ;
        RECT 84.680 169.820 84.940 170.140 ;
        RECT 85.200 169.800 85.340 171.520 ;
        RECT 89.340 170.140 89.480 171.520 ;
        RECT 91.880 170.305 93.760 170.675 ;
        RECT 89.280 169.820 89.540 170.140 ;
        RECT 85.140 169.480 85.400 169.800 ;
        RECT 86.980 169.480 87.240 169.800 ;
        RECT 84.220 168.800 84.480 169.120 ;
        RECT 87.040 168.440 87.180 169.480 ;
        RECT 87.440 168.800 87.700 169.120 ;
        RECT 85.140 168.120 85.400 168.440 ;
        RECT 86.980 168.120 87.240 168.440 ;
        RECT 85.200 166.400 85.340 168.120 ;
        RECT 86.060 166.420 86.320 166.740 ;
        RECT 85.140 166.080 85.400 166.400 ;
        RECT 83.300 165.400 83.560 165.720 ;
        RECT 84.220 165.400 84.480 165.720 ;
        RECT 83.360 164.700 83.500 165.400 ;
        RECT 83.300 164.380 83.560 164.700 ;
        RECT 83.760 162.680 84.020 163.000 ;
        RECT 83.820 161.640 83.960 162.680 ;
        RECT 83.760 161.320 84.020 161.640 ;
        RECT 84.280 161.300 84.420 165.400 ;
        RECT 85.200 164.020 85.340 166.080 ;
        RECT 85.140 163.700 85.400 164.020 ;
        RECT 85.600 163.700 85.860 164.020 ;
        RECT 85.660 161.980 85.800 163.700 ;
        RECT 86.120 163.000 86.260 166.420 ;
        RECT 87.040 166.400 87.180 168.120 ;
        RECT 87.500 167.420 87.640 168.800 ;
        RECT 91.120 168.120 91.380 168.440 ;
        RECT 87.440 167.100 87.700 167.420 ;
        RECT 86.980 166.080 87.240 166.400 ;
        RECT 86.520 163.020 86.780 163.340 ;
        RECT 86.060 162.680 86.320 163.000 ;
        RECT 85.600 161.660 85.860 161.980 ;
        RECT 84.220 160.980 84.480 161.300 ;
        RECT 83.300 160.815 83.560 160.960 ;
        RECT 83.290 160.445 83.570 160.815 ;
        RECT 86.120 160.620 86.260 162.680 ;
        RECT 86.580 161.980 86.720 163.020 ;
        RECT 86.520 161.660 86.780 161.980 ;
        RECT 87.500 161.300 87.640 167.100 ;
        RECT 91.180 163.680 91.320 168.120 ;
        RECT 91.880 164.865 93.760 165.235 ;
        RECT 93.940 164.020 94.080 171.860 ;
        RECT 97.560 171.520 97.820 171.840 ;
        RECT 97.620 169.460 97.760 171.520 ;
        RECT 97.560 169.140 97.820 169.460 ;
        RECT 98.080 167.420 98.220 172.540 ;
        RECT 98.480 168.120 98.740 168.440 ;
        RECT 98.020 167.100 98.280 167.420 ;
        RECT 94.340 166.420 94.600 166.740 ;
        RECT 94.400 164.700 94.540 166.420 ;
        RECT 94.800 166.080 95.060 166.400 ;
        RECT 94.340 164.380 94.600 164.700 ;
        RECT 93.880 163.700 94.140 164.020 ;
        RECT 91.120 163.360 91.380 163.680 ;
        RECT 87.440 160.980 87.700 161.300 ;
        RECT 86.060 160.300 86.320 160.620 ;
        RECT 87.500 160.140 87.640 160.980 ;
        RECT 93.940 160.960 94.080 163.700 ;
        RECT 94.860 163.680 95.000 166.080 ;
        RECT 96.640 165.400 96.900 165.720 ;
        RECT 94.800 163.360 95.060 163.680 ;
        RECT 96.180 162.680 96.440 163.000 ;
        RECT 93.880 160.640 94.140 160.960 ;
        RECT 82.900 160.000 83.500 160.140 ;
        RECT 80.540 157.580 80.800 157.900 ;
        RECT 80.600 150.420 80.740 157.580 ;
        RECT 81.460 154.520 81.720 154.840 ;
        RECT 80.540 150.100 80.800 150.420 ;
        RECT 80.600 147.360 80.740 150.100 ;
        RECT 81.520 149.740 81.660 154.520 ;
        RECT 83.360 150.420 83.500 160.000 ;
        RECT 87.040 160.000 87.640 160.140 ;
        RECT 87.040 152.800 87.180 160.000 ;
        RECT 91.880 159.425 93.760 159.795 ;
        RECT 93.880 155.540 94.140 155.860 ;
        RECT 91.880 153.985 93.760 154.355 ;
        RECT 86.980 152.480 87.240 152.800 ;
        RECT 86.520 152.140 86.780 152.460 ;
        RECT 83.300 150.100 83.560 150.420 ;
        RECT 83.760 150.100 84.020 150.420 ;
        RECT 81.000 149.420 81.260 149.740 ;
        RECT 81.460 149.420 81.720 149.740 ;
        RECT 80.540 147.040 80.800 147.360 ;
        RECT 80.540 146.360 80.800 146.680 ;
        RECT 80.600 142.260 80.740 146.360 ;
        RECT 80.540 141.940 80.800 142.260 ;
        RECT 80.080 141.600 80.340 141.920 ;
        RECT 79.620 141.095 79.880 141.240 ;
        RECT 79.610 140.725 79.890 141.095 ;
        RECT 81.060 136.820 81.200 149.420 ;
        RECT 82.380 149.255 82.640 149.400 ;
        RECT 82.370 148.885 82.650 149.255 ;
        RECT 83.820 148.040 83.960 150.100 ;
        RECT 86.580 150.080 86.720 152.140 ;
        RECT 88.360 151.800 88.620 152.120 ;
        RECT 88.420 150.760 88.560 151.800 ;
        RECT 93.940 151.100 94.080 155.540 ;
        RECT 95.720 154.520 95.980 154.840 ;
        RECT 95.780 153.140 95.920 154.520 ;
        RECT 95.720 152.820 95.980 153.140 ;
        RECT 93.880 150.780 94.140 151.100 ;
        RECT 88.360 150.440 88.620 150.760 ;
        RECT 91.120 150.100 91.380 150.420 ;
        RECT 86.520 149.760 86.780 150.080 ;
        RECT 85.600 148.060 85.860 148.380 ;
        RECT 83.760 147.720 84.020 148.040 ;
        RECT 81.920 147.040 82.180 147.360 ;
        RECT 83.300 147.040 83.560 147.360 ;
        RECT 81.460 146.360 81.720 146.680 ;
        RECT 81.000 136.500 81.260 136.820 ;
        RECT 81.000 135.820 81.260 136.140 ;
        RECT 81.060 134.780 81.200 135.820 ;
        RECT 81.000 134.460 81.260 134.780 ;
        RECT 80.990 131.885 81.270 132.255 ;
        RECT 81.060 131.040 81.200 131.885 ;
        RECT 81.520 131.380 81.660 146.360 ;
        RECT 81.980 145.175 82.120 147.040 ;
        RECT 82.380 146.360 82.640 146.680 ;
        RECT 81.910 144.805 82.190 145.175 ;
        RECT 81.980 144.300 82.120 144.805 ;
        RECT 81.920 143.980 82.180 144.300 ;
        RECT 82.440 141.920 82.580 146.360 ;
        RECT 82.830 145.485 83.110 145.855 ;
        RECT 82.900 144.980 83.040 145.485 ;
        RECT 82.840 144.660 83.100 144.980 ;
        RECT 83.360 144.380 83.500 147.040 ;
        RECT 83.820 144.980 83.960 147.720 ;
        RECT 85.660 147.360 85.800 148.060 ;
        RECT 84.220 147.040 84.480 147.360 ;
        RECT 85.600 147.040 85.860 147.360 ;
        RECT 83.760 144.660 84.020 144.980 ;
        RECT 82.900 144.240 83.500 144.380 ;
        RECT 82.900 141.920 83.040 144.240 ;
        RECT 83.300 142.620 83.560 142.940 ;
        RECT 82.380 141.600 82.640 141.920 ;
        RECT 82.840 141.600 83.100 141.920 ;
        RECT 82.900 139.880 83.040 141.600 ;
        RECT 81.920 139.560 82.180 139.880 ;
        RECT 82.840 139.560 83.100 139.880 ;
        RECT 81.980 134.100 82.120 139.560 ;
        RECT 82.840 137.180 83.100 137.500 ;
        RECT 81.920 133.780 82.180 134.100 ;
        RECT 82.380 132.760 82.640 133.080 ;
        RECT 81.920 131.740 82.180 132.060 ;
        RECT 81.460 131.060 81.720 131.380 ;
        RECT 81.000 130.720 81.260 131.040 ;
        RECT 81.460 130.040 81.720 130.360 ;
        RECT 80.080 125.620 80.340 125.940 ;
        RECT 79.620 125.280 79.880 125.600 ;
        RECT 79.160 124.600 79.420 124.920 ;
        RECT 76.880 124.065 78.760 124.435 ;
        RECT 79.160 123.240 79.420 123.560 ;
        RECT 76.880 118.625 78.760 118.995 ;
        RECT 79.220 116.760 79.360 123.240 ;
        RECT 79.680 122.880 79.820 125.280 ;
        RECT 80.140 123.560 80.280 125.620 ;
        RECT 80.080 123.240 80.340 123.560 ;
        RECT 79.620 122.560 79.880 122.880 ;
        RECT 79.680 121.180 79.820 122.560 ;
        RECT 79.620 120.860 79.880 121.180 ;
        RECT 80.080 117.800 80.340 118.120 ;
        RECT 79.160 116.440 79.420 116.760 ;
        RECT 76.880 113.185 78.760 113.555 ;
        RECT 79.220 113.020 79.360 116.440 ;
        RECT 80.140 115.740 80.280 117.800 ;
        RECT 80.080 115.420 80.340 115.740 ;
        RECT 79.160 112.700 79.420 113.020 ;
        RECT 80.540 112.020 80.800 112.340 ;
        RECT 80.080 111.680 80.340 112.000 ;
        RECT 77.780 111.000 78.040 111.320 ;
        RECT 76.400 109.980 76.660 110.300 ;
        RECT 75.940 109.300 76.200 109.620 ;
        RECT 76.400 108.960 76.660 109.280 ;
        RECT 77.840 109.190 77.980 111.000 ;
        RECT 78.240 109.190 78.500 109.280 ;
        RECT 77.840 109.050 78.500 109.190 ;
        RECT 78.240 108.960 78.500 109.050 ;
        RECT 74.100 106.580 74.360 106.900 ;
        RECT 74.160 104.180 74.300 106.580 ;
        RECT 74.100 103.860 74.360 104.180 ;
        RECT 74.100 103.180 74.360 103.500 ;
        RECT 67.730 89.640 68.670 89.840 ;
        RECT 62.130 88.870 62.410 89.170 ;
        RECT 61.720 88.640 62.940 88.870 ;
        RECT 61.720 88.620 63.130 88.640 ;
        RECT 60.820 88.480 63.130 88.620 ;
        RECT 43.810 85.660 45.030 86.720 ;
        RECT 49.740 85.170 50.960 86.920 ;
        RECT 55.530 85.320 56.750 88.480 ;
        RECT 61.720 86.600 63.130 88.480 ;
        RECT 61.720 85.000 62.940 86.600 ;
        RECT 67.580 85.770 68.800 89.640 ;
        RECT 74.160 89.170 74.300 103.180 ;
        RECT 76.460 101.800 76.600 108.960 ;
        RECT 79.620 108.280 79.880 108.600 ;
        RECT 76.880 107.745 78.760 108.115 ;
        RECT 79.680 103.840 79.820 108.280 ;
        RECT 80.140 107.240 80.280 111.680 ;
        RECT 80.600 108.940 80.740 112.020 ;
        RECT 80.990 111.485 81.270 111.855 ;
        RECT 81.520 111.840 81.660 130.040 ;
        RECT 81.980 126.620 82.120 131.740 ;
        RECT 82.440 131.040 82.580 132.760 ;
        RECT 82.380 130.720 82.640 131.040 ;
        RECT 82.900 129.340 83.040 137.180 ;
        RECT 82.840 129.020 83.100 129.340 ;
        RECT 82.380 128.340 82.640 128.660 ;
        RECT 81.920 126.300 82.180 126.620 ;
        RECT 82.440 125.940 82.580 128.340 ;
        RECT 82.380 125.620 82.640 125.940 ;
        RECT 83.360 125.600 83.500 142.620 ;
        RECT 83.760 141.830 84.020 141.920 ;
        RECT 84.280 141.830 84.420 147.040 ;
        RECT 85.660 143.700 85.800 147.040 ;
        RECT 86.060 146.700 86.320 147.020 ;
        RECT 86.120 144.640 86.260 146.700 ;
        RECT 86.580 145.740 86.720 149.760 ;
        RECT 86.580 145.660 87.180 145.740 ;
        RECT 86.520 145.600 87.180 145.660 ;
        RECT 86.520 145.340 86.780 145.600 ;
        RECT 86.520 144.660 86.780 144.980 ;
        RECT 86.060 144.320 86.320 144.640 ;
        RECT 85.660 143.560 86.260 143.700 ;
        RECT 86.120 141.920 86.260 143.560 ;
        RECT 83.760 141.690 84.880 141.830 ;
        RECT 83.760 141.600 84.020 141.690 ;
        RECT 84.220 135.480 84.480 135.800 ;
        RECT 83.760 128.340 84.020 128.660 ;
        RECT 83.300 125.280 83.560 125.600 ;
        RECT 83.820 123.900 83.960 128.340 ;
        RECT 83.760 123.580 84.020 123.900 ;
        RECT 82.840 121.880 83.100 122.200 ;
        RECT 82.900 114.720 83.040 121.880 ;
        RECT 83.820 121.180 83.960 123.580 ;
        RECT 83.760 120.860 84.020 121.180 ;
        RECT 83.760 117.120 84.020 117.440 ;
        RECT 83.820 115.740 83.960 117.120 ;
        RECT 83.760 115.420 84.020 115.740 ;
        RECT 82.840 114.400 83.100 114.720 ;
        RECT 81.520 111.700 82.580 111.840 ;
        RECT 81.060 109.280 81.200 111.485 ;
        RECT 81.000 108.960 81.260 109.280 ;
        RECT 80.540 108.620 80.800 108.940 ;
        RECT 81.920 108.280 82.180 108.600 ;
        RECT 80.080 106.920 80.340 107.240 ;
        RECT 80.080 106.240 80.340 106.560 ;
        RECT 79.620 103.520 79.880 103.840 ;
        RECT 76.880 102.305 78.760 102.675 ;
        RECT 76.400 101.480 76.660 101.800 ;
        RECT 80.140 89.170 80.280 106.240 ;
        RECT 81.980 104.180 82.120 108.280 ;
        RECT 82.440 107.580 82.580 111.700 ;
        RECT 84.280 109.620 84.420 135.480 ;
        RECT 84.740 134.100 84.880 141.690 ;
        RECT 86.060 141.600 86.320 141.920 ;
        RECT 86.120 134.100 86.260 141.600 ;
        RECT 86.580 141.580 86.720 144.660 ;
        RECT 86.520 141.260 86.780 141.580 ;
        RECT 87.040 136.820 87.180 145.600 ;
        RECT 91.180 144.640 91.320 150.100 ;
        RECT 91.880 148.545 93.760 148.915 ;
        RECT 96.240 147.360 96.380 162.680 ;
        RECT 96.700 161.300 96.840 165.400 ;
        RECT 98.080 163.680 98.220 167.100 ;
        RECT 98.540 166.400 98.680 168.120 ;
        RECT 98.480 166.080 98.740 166.400 ;
        RECT 98.020 163.360 98.280 163.680 ;
        RECT 96.640 160.980 96.900 161.300 ;
        RECT 97.100 160.640 97.360 160.960 ;
        RECT 97.160 155.520 97.300 160.640 ;
        RECT 99.400 159.960 99.660 160.280 ;
        RECT 99.460 159.260 99.600 159.960 ;
        RECT 99.400 158.940 99.660 159.260 ;
        RECT 99.920 155.860 100.060 177.300 ;
        RECT 100.380 175.580 100.520 177.300 ;
        RECT 101.300 175.580 101.440 183.080 ;
        RECT 101.690 177.445 101.970 177.815 ;
        RECT 101.700 177.300 101.960 177.445 ;
        RECT 100.320 175.260 100.580 175.580 ;
        RECT 101.240 175.260 101.500 175.580 ;
        RECT 101.300 172.860 101.440 175.260 ;
        RECT 101.240 172.770 101.500 172.860 ;
        RECT 101.240 172.630 101.900 172.770 ;
        RECT 101.240 172.540 101.500 172.630 ;
        RECT 101.760 169.460 101.900 172.630 ;
        RECT 101.700 169.140 101.960 169.460 ;
        RECT 101.700 168.460 101.960 168.780 ;
        RECT 100.320 168.180 100.580 168.440 ;
        RECT 101.760 168.180 101.900 168.460 ;
        RECT 100.320 168.120 101.900 168.180 ;
        RECT 100.380 168.040 101.900 168.120 ;
        RECT 100.380 163.680 100.520 168.040 ;
        RECT 100.320 163.360 100.580 163.680 ;
        RECT 101.240 163.360 101.500 163.680 ;
        RECT 101.300 161.980 101.440 163.360 ;
        RECT 101.240 161.660 101.500 161.980 ;
        RECT 101.700 160.980 101.960 161.300 ;
        RECT 101.760 158.240 101.900 160.980 ;
        RECT 101.700 157.920 101.960 158.240 ;
        RECT 101.760 155.860 101.900 157.920 ;
        RECT 102.220 155.860 102.360 185.120 ;
        RECT 102.680 185.100 102.820 193.620 ;
        RECT 102.620 184.780 102.880 185.100 ;
        RECT 102.620 172.540 102.880 172.860 ;
        RECT 102.680 170.140 102.820 172.540 ;
        RECT 102.620 169.820 102.880 170.140 ;
        RECT 99.860 155.540 100.120 155.860 ;
        RECT 101.700 155.540 101.960 155.860 ;
        RECT 102.160 155.540 102.420 155.860 ;
        RECT 97.100 155.200 97.360 155.520 ;
        RECT 97.160 153.140 97.300 155.200 ;
        RECT 97.560 154.520 97.820 154.840 ;
        RECT 97.100 152.820 97.360 153.140 ;
        RECT 97.620 147.700 97.760 154.520 ;
        RECT 101.760 152.800 101.900 155.540 ;
        RECT 103.140 152.800 103.280 193.960 ;
        RECT 103.540 192.940 103.800 193.260 ;
        RECT 103.600 190.200 103.740 192.940 ;
        RECT 104.000 192.600 104.260 192.920 ;
        RECT 104.060 190.540 104.200 192.600 ;
        RECT 104.000 190.220 104.260 190.540 ;
        RECT 103.540 189.880 103.800 190.200 ;
        RECT 103.600 185.180 103.740 189.880 ;
        RECT 104.460 188.520 104.720 188.840 ;
        RECT 104.520 186.120 104.660 188.520 ;
        RECT 104.460 185.800 104.720 186.120 ;
        RECT 103.600 185.040 104.200 185.180 ;
        RECT 104.060 184.760 104.200 185.040 ;
        RECT 103.540 184.440 103.800 184.760 ;
        RECT 104.000 184.440 104.260 184.760 ;
        RECT 103.600 183.060 103.740 184.440 ;
        RECT 103.540 182.740 103.800 183.060 ;
        RECT 104.060 182.460 104.200 184.440 ;
        RECT 103.600 182.320 104.200 182.460 ;
        RECT 103.600 160.140 103.740 182.320 ;
        RECT 104.000 168.120 104.260 168.440 ;
        RECT 104.060 166.740 104.200 168.120 ;
        RECT 104.000 166.420 104.260 166.740 ;
        RECT 104.980 161.980 105.120 195.660 ;
        RECT 105.440 193.600 105.580 196.340 ;
        RECT 105.840 196.060 106.100 196.320 ;
        RECT 105.840 196.000 106.500 196.060 ;
        RECT 105.900 195.920 106.500 196.000 ;
        RECT 105.840 195.320 106.100 195.640 ;
        RECT 105.900 194.280 106.040 195.320 ;
        RECT 105.840 193.960 106.100 194.280 ;
        RECT 105.380 193.280 105.640 193.600 ;
        RECT 105.440 185.780 105.580 193.280 ;
        RECT 105.380 185.460 105.640 185.780 ;
        RECT 105.840 171.860 106.100 172.180 ;
        RECT 105.900 169.120 106.040 171.860 ;
        RECT 106.360 169.655 106.500 195.920 ;
        RECT 106.880 194.785 108.760 195.155 ;
        RECT 110.900 192.600 111.160 192.920 ;
        RECT 110.960 191.220 111.100 192.600 ;
        RECT 110.900 190.900 111.160 191.220 ;
        RECT 112.340 190.880 112.480 198.720 ;
        RECT 121.880 197.505 123.760 197.875 ;
        RECT 121.880 192.065 123.760 192.435 ;
        RECT 112.280 190.560 112.540 190.880 ;
        RECT 113.660 190.560 113.920 190.880 ;
        RECT 106.880 189.345 108.760 189.715 ;
        RECT 112.340 188.160 112.480 190.560 ;
        RECT 112.280 187.840 112.540 188.160 ;
        RECT 108.140 187.160 108.400 187.480 ;
        RECT 108.200 186.460 108.340 187.160 ;
        RECT 108.140 186.140 108.400 186.460 ;
        RECT 113.720 185.440 113.860 190.560 ;
        RECT 118.720 189.880 118.980 190.200 ;
        RECT 118.780 188.840 118.920 189.880 ;
        RECT 118.720 188.520 118.980 188.840 ;
        RECT 125.620 187.840 125.880 188.160 ;
        RECT 117.340 187.160 117.600 187.480 ;
        RECT 124.240 187.160 124.500 187.480 ;
        RECT 116.880 185.800 117.140 186.120 ;
        RECT 113.660 185.120 113.920 185.440 ;
        RECT 106.880 183.905 108.760 184.275 ;
        RECT 109.060 182.740 109.320 183.060 ;
        RECT 108.140 181.720 108.400 182.040 ;
        RECT 108.200 179.660 108.340 181.720 ;
        RECT 109.120 180.340 109.260 182.740 ;
        RECT 113.720 182.380 113.860 185.120 ;
        RECT 116.940 183.060 117.080 185.800 ;
        RECT 116.880 182.740 117.140 183.060 ;
        RECT 113.660 182.060 113.920 182.380 ;
        RECT 113.200 181.720 113.460 182.040 ;
        RECT 109.060 180.020 109.320 180.340 ;
        RECT 108.140 179.340 108.400 179.660 ;
        RECT 109.120 179.320 109.260 180.020 ;
        RECT 109.060 179.000 109.320 179.320 ;
        RECT 106.880 178.465 108.760 178.835 ;
        RECT 106.880 173.025 108.760 173.395 ;
        RECT 106.290 169.285 106.570 169.655 ;
        RECT 105.840 168.800 106.100 169.120 ;
        RECT 106.760 168.860 107.020 169.120 ;
        RECT 106.360 168.800 107.020 168.860 ;
        RECT 105.380 168.120 105.640 168.440 ;
        RECT 104.920 161.660 105.180 161.980 ;
        RECT 104.000 160.980 104.260 161.300 ;
        RECT 104.920 160.980 105.180 161.300 ;
        RECT 104.060 160.700 104.200 160.980 ;
        RECT 104.060 160.560 104.660 160.700 ;
        RECT 103.600 160.000 104.200 160.140 ;
        RECT 104.060 158.240 104.200 160.000 ;
        RECT 104.520 159.260 104.660 160.560 ;
        RECT 104.460 158.940 104.720 159.260 ;
        RECT 104.520 158.240 104.660 158.940 ;
        RECT 104.980 158.240 105.120 160.980 ;
        RECT 104.000 157.920 104.260 158.240 ;
        RECT 104.460 157.920 104.720 158.240 ;
        RECT 104.920 157.920 105.180 158.240 ;
        RECT 103.540 157.580 103.800 157.900 ;
        RECT 103.600 156.540 103.740 157.580 ;
        RECT 103.540 156.220 103.800 156.540 ;
        RECT 103.600 155.860 103.740 156.220 ;
        RECT 104.520 156.200 104.660 157.920 ;
        RECT 104.460 155.940 104.720 156.200 ;
        RECT 104.060 155.880 104.720 155.940 ;
        RECT 103.540 155.540 103.800 155.860 ;
        RECT 104.060 155.800 104.660 155.880 ;
        RECT 103.600 153.480 103.740 155.540 ;
        RECT 103.540 153.160 103.800 153.480 ;
        RECT 104.060 152.800 104.200 155.800 ;
        RECT 104.460 154.860 104.720 155.180 ;
        RECT 99.390 152.285 99.670 152.655 ;
        RECT 101.700 152.480 101.960 152.800 ;
        RECT 103.080 152.480 103.340 152.800 ;
        RECT 104.000 152.480 104.260 152.800 ;
        RECT 99.460 150.080 99.600 152.285 ;
        RECT 99.860 152.140 100.120 152.460 ;
        RECT 99.400 149.760 99.660 150.080 ;
        RECT 98.020 148.060 98.280 148.380 ;
        RECT 97.560 147.380 97.820 147.700 ;
        RECT 94.340 147.040 94.600 147.360 ;
        RECT 96.180 147.040 96.440 147.360 ;
        RECT 92.960 146.360 93.220 146.680 ;
        RECT 93.020 145.320 93.160 146.360 ;
        RECT 92.960 145.000 93.220 145.320 ;
        RECT 91.120 144.320 91.380 144.640 ;
        RECT 88.360 143.640 88.620 143.960 ;
        RECT 88.420 142.260 88.560 143.640 ;
        RECT 91.880 143.105 93.760 143.475 ;
        RECT 88.360 141.940 88.620 142.260 ;
        RECT 91.120 141.600 91.380 141.920 ;
        RECT 89.740 141.260 90.000 141.580 ;
        RECT 89.800 140.220 89.940 141.260 ;
        RECT 89.740 139.900 90.000 140.220 ;
        RECT 89.800 136.820 89.940 139.900 ;
        RECT 91.180 137.500 91.320 141.600 ;
        RECT 93.880 139.560 94.140 139.880 ;
        RECT 91.880 137.665 93.760 138.035 ;
        RECT 93.940 137.500 94.080 139.560 ;
        RECT 91.120 137.180 91.380 137.500 ;
        RECT 93.880 137.180 94.140 137.500 ;
        RECT 86.980 136.500 87.240 136.820 ;
        RECT 89.740 136.500 90.000 136.820 ;
        RECT 94.400 136.480 94.540 147.040 ;
        RECT 96.640 144.320 96.900 144.640 ;
        RECT 96.700 142.940 96.840 144.320 ;
        RECT 96.640 142.620 96.900 142.940 ;
        RECT 96.640 140.920 96.900 141.240 ;
        RECT 96.700 139.540 96.840 140.920 ;
        RECT 96.640 139.220 96.900 139.540 ;
        RECT 90.200 136.160 90.460 136.480 ;
        RECT 94.340 136.160 94.600 136.480 ;
        RECT 89.740 135.480 90.000 135.800 ;
        RECT 89.800 134.100 89.940 135.480 ;
        RECT 84.680 133.780 84.940 134.100 ;
        RECT 86.060 133.780 86.320 134.100 ;
        RECT 89.740 133.780 90.000 134.100 ;
        RECT 86.120 133.420 86.260 133.780 ;
        RECT 86.060 133.100 86.320 133.420 ;
        RECT 89.800 132.060 89.940 133.780 ;
        RECT 90.260 133.760 90.400 136.160 ;
        RECT 90.200 133.440 90.460 133.760 ;
        RECT 91.880 132.225 93.760 132.595 ;
        RECT 89.740 131.740 90.000 132.060 ;
        RECT 94.400 130.950 94.540 136.160 ;
        RECT 97.560 135.480 97.820 135.800 ;
        RECT 97.620 134.440 97.760 135.480 ;
        RECT 97.560 134.120 97.820 134.440 ;
        RECT 95.260 132.760 95.520 133.080 ;
        RECT 95.320 131.380 95.460 132.760 ;
        RECT 95.260 131.060 95.520 131.380 ;
        RECT 94.800 130.950 95.060 131.040 ;
        RECT 94.400 130.810 95.060 130.950 ;
        RECT 93.420 130.380 93.680 130.700 ;
        RECT 93.480 129.340 93.620 130.380 ;
        RECT 93.420 129.020 93.680 129.340 ;
        RECT 94.400 128.660 94.540 130.810 ;
        RECT 94.800 130.720 95.060 130.810 ;
        RECT 98.080 129.340 98.220 148.060 ;
        RECT 99.460 147.360 99.600 149.760 ;
        RECT 99.920 149.400 100.060 152.140 ;
        RECT 104.000 151.800 104.260 152.120 ;
        RECT 104.060 150.760 104.200 151.800 ;
        RECT 104.000 150.440 104.260 150.760 ;
        RECT 104.520 150.080 104.660 154.860 ;
        RECT 104.920 154.520 105.180 154.840 ;
        RECT 104.460 149.760 104.720 150.080 ;
        RECT 101.240 149.420 101.500 149.740 ;
        RECT 99.860 149.080 100.120 149.400 ;
        RECT 99.920 147.360 100.060 149.080 ;
        RECT 101.300 147.360 101.440 149.420 ;
        RECT 104.000 149.080 104.260 149.400 ;
        RECT 99.400 147.040 99.660 147.360 ;
        RECT 99.860 147.040 100.120 147.360 ;
        RECT 100.320 147.040 100.580 147.360 ;
        RECT 101.240 147.040 101.500 147.360 ;
        RECT 99.460 144.980 99.600 147.040 ;
        RECT 99.400 144.660 99.660 144.980 ;
        RECT 98.480 144.320 98.740 144.640 ;
        RECT 98.540 139.540 98.680 144.320 ;
        RECT 98.480 139.220 98.740 139.540 ;
        RECT 98.540 131.380 98.680 139.220 ;
        RECT 100.380 138.520 100.520 147.040 ;
        RECT 103.080 146.360 103.340 146.680 ;
        RECT 99.400 138.200 99.660 138.520 ;
        RECT 100.320 138.200 100.580 138.520 ;
        RECT 99.460 136.480 99.600 138.200 ;
        RECT 99.400 136.160 99.660 136.480 ;
        RECT 100.780 134.120 101.040 134.440 ;
        RECT 100.840 132.060 100.980 134.120 ;
        RECT 100.780 131.740 101.040 132.060 ;
        RECT 98.480 131.060 98.740 131.380 ;
        RECT 98.020 129.020 98.280 129.340 ;
        RECT 94.340 128.340 94.600 128.660 ;
        RECT 91.880 126.785 93.760 127.155 ;
        RECT 84.680 125.620 84.940 125.940 ;
        RECT 84.740 117.440 84.880 125.620 ;
        RECT 95.720 125.280 95.980 125.600 ;
        RECT 95.780 123.900 95.920 125.280 ;
        RECT 97.560 124.600 97.820 124.920 ;
        RECT 95.720 123.580 95.980 123.900 ;
        RECT 90.660 122.900 90.920 123.220 ;
        RECT 90.200 122.560 90.460 122.880 ;
        RECT 88.820 121.880 89.080 122.200 ;
        RECT 86.060 120.180 86.320 120.500 ;
        RECT 86.120 117.780 86.260 120.180 ;
        RECT 88.880 120.160 89.020 121.880 ;
        RECT 88.820 119.840 89.080 120.160 ;
        RECT 90.260 119.480 90.400 122.560 ;
        RECT 87.440 119.160 87.700 119.480 ;
        RECT 90.200 119.160 90.460 119.480 ;
        RECT 87.500 117.780 87.640 119.160 ;
        RECT 89.270 118.285 89.550 118.655 ;
        RECT 89.340 118.120 89.480 118.285 ;
        RECT 89.280 117.800 89.540 118.120 ;
        RECT 86.060 117.460 86.320 117.780 ;
        RECT 87.440 117.460 87.700 117.780 ;
        RECT 84.680 117.120 84.940 117.440 ;
        RECT 84.740 115.740 84.880 117.120 ;
        RECT 84.680 115.420 84.940 115.740 ;
        RECT 84.740 112.680 84.880 115.420 ;
        RECT 87.500 115.060 87.640 117.460 ;
        RECT 87.900 116.440 88.160 116.760 ;
        RECT 87.440 114.740 87.700 115.060 ;
        RECT 87.960 114.380 88.100 116.440 ;
        RECT 87.900 114.060 88.160 114.380 ;
        RECT 84.680 112.360 84.940 112.680 ;
        RECT 90.260 112.000 90.400 119.160 ;
        RECT 90.720 117.780 90.860 122.900 ;
        RECT 91.120 121.880 91.380 122.200 ;
        RECT 91.180 119.820 91.320 121.880 ;
        RECT 91.880 121.345 93.760 121.715 ;
        RECT 97.620 120.500 97.760 124.600 ;
        RECT 98.540 122.880 98.680 131.060 ;
        RECT 98.940 130.720 99.200 131.040 ;
        RECT 99.000 125.600 99.140 130.720 ;
        RECT 100.320 130.040 100.580 130.360 ;
        RECT 100.380 128.660 100.520 130.040 ;
        RECT 100.320 128.340 100.580 128.660 ;
        RECT 101.240 128.000 101.500 128.320 ;
        RECT 98.940 125.280 99.200 125.600 ;
        RECT 101.300 123.900 101.440 128.000 ;
        RECT 102.620 125.280 102.880 125.600 ;
        RECT 101.240 123.580 101.500 123.900 ;
        RECT 98.940 123.240 99.200 123.560 ;
        RECT 98.480 122.560 98.740 122.880 ;
        RECT 97.560 120.180 97.820 120.500 ;
        RECT 98.540 120.160 98.680 122.560 ;
        RECT 98.480 119.840 98.740 120.160 ;
        RECT 91.120 119.500 91.380 119.820 ;
        RECT 98.540 118.460 98.680 119.840 ;
        RECT 99.000 118.460 99.140 123.240 ;
        RECT 98.480 118.140 98.740 118.460 ;
        RECT 98.940 118.140 99.200 118.460 ;
        RECT 90.660 117.460 90.920 117.780 ;
        RECT 91.880 115.905 93.760 116.275 ;
        RECT 98.540 115.060 98.680 118.140 ;
        RECT 102.680 117.780 102.820 125.280 ;
        RECT 102.620 117.460 102.880 117.780 ;
        RECT 98.480 114.740 98.740 115.060 ;
        RECT 95.260 114.400 95.520 114.720 ;
        RECT 95.320 113.020 95.460 114.400 ;
        RECT 95.260 112.700 95.520 113.020 ;
        RECT 90.200 111.680 90.460 112.000 ;
        RECT 98.540 111.740 98.680 114.740 ;
        RECT 98.540 111.600 99.140 111.740 ;
        RECT 91.880 110.465 93.760 110.835 ;
        RECT 99.000 110.300 99.140 111.600 ;
        RECT 98.940 109.980 99.200 110.300 ;
        RECT 84.220 109.300 84.480 109.620 ;
        RECT 98.020 109.300 98.280 109.620 ;
        RECT 84.220 108.620 84.480 108.940 ;
        RECT 97.560 108.620 97.820 108.940 ;
        RECT 83.300 108.280 83.560 108.600 ;
        RECT 82.380 107.260 82.640 107.580 ;
        RECT 83.360 107.240 83.500 108.280 ;
        RECT 84.280 107.240 84.420 108.620 ;
        RECT 88.820 108.280 89.080 108.600 ;
        RECT 90.660 108.280 90.920 108.600 ;
        RECT 88.880 107.580 89.020 108.280 ;
        RECT 88.820 107.260 89.080 107.580 ;
        RECT 90.720 107.240 90.860 108.280 ;
        RECT 83.300 106.920 83.560 107.240 ;
        RECT 84.220 106.920 84.480 107.240 ;
        RECT 90.660 106.920 90.920 107.240 ;
        RECT 89.280 106.240 89.540 106.560 ;
        RECT 93.880 106.240 94.140 106.560 ;
        RECT 87.440 105.560 87.700 105.880 ;
        RECT 87.900 105.560 88.160 105.880 ;
        RECT 81.920 103.860 82.180 104.180 ;
        RECT 87.500 103.500 87.640 105.560 ;
        RECT 87.960 104.180 88.100 105.560 ;
        RECT 89.340 104.860 89.480 106.240 ;
        RECT 91.880 105.025 93.760 105.395 ;
        RECT 89.280 104.540 89.540 104.860 ;
        RECT 87.900 103.860 88.160 104.180 ;
        RECT 87.440 103.180 87.700 103.500 ;
        RECT 86.060 102.840 86.320 103.160 ;
        RECT 86.120 89.170 86.260 102.840 ;
        RECT 91.880 99.585 93.760 99.955 ;
        RECT 74.090 88.160 74.370 89.170 ;
        RECT 80.070 88.180 80.350 89.170 ;
        RECT 73.850 84.290 75.070 88.160 ;
        RECT 79.730 84.310 80.950 88.180 ;
        RECT 86.050 87.970 86.330 89.170 ;
        RECT 92.030 88.620 92.310 89.170 ;
        RECT 93.940 88.620 94.080 106.240 ;
        RECT 97.620 104.860 97.760 108.620 ;
        RECT 97.560 104.540 97.820 104.860 ;
        RECT 98.080 89.170 98.220 109.300 ;
        RECT 99.000 104.180 99.140 109.980 ;
        RECT 103.140 109.280 103.280 146.360 ;
        RECT 104.060 132.060 104.200 149.080 ;
        RECT 104.980 144.640 105.120 154.520 ;
        RECT 105.440 150.420 105.580 168.120 ;
        RECT 105.900 167.420 106.040 168.800 ;
        RECT 106.360 168.720 106.960 168.800 ;
        RECT 105.840 167.100 106.100 167.420 ;
        RECT 105.830 166.565 106.110 166.935 ;
        RECT 105.900 162.740 106.040 166.565 ;
        RECT 106.360 163.340 106.500 168.720 ;
        RECT 106.880 167.585 108.760 167.955 ;
        RECT 108.600 167.100 108.860 167.420 ;
        RECT 108.660 166.740 108.800 167.100 ;
        RECT 108.600 166.420 108.860 166.740 ;
        RECT 108.660 164.700 108.800 166.420 ;
        RECT 108.600 164.380 108.860 164.700 ;
        RECT 108.660 163.680 108.800 164.380 ;
        RECT 109.120 164.020 109.260 179.000 ;
        RECT 113.260 177.620 113.400 181.720 ;
        RECT 113.200 177.300 113.460 177.620 ;
        RECT 111.820 176.960 112.080 177.280 ;
        RECT 111.880 174.560 112.020 176.960 ;
        RECT 113.720 175.240 113.860 182.060 ;
        RECT 115.960 179.340 116.220 179.660 ;
        RECT 114.580 179.000 114.840 179.320 ;
        RECT 113.660 174.920 113.920 175.240 ;
        RECT 111.820 174.240 112.080 174.560 ;
        RECT 112.280 171.860 112.540 172.180 ;
        RECT 114.120 171.860 114.380 172.180 ;
        RECT 109.980 171.520 110.240 171.840 ;
        RECT 109.520 170.840 109.780 171.160 ;
        RECT 109.060 163.700 109.320 164.020 ;
        RECT 108.600 163.360 108.860 163.680 ;
        RECT 106.300 163.020 106.560 163.340 ;
        RECT 105.900 162.600 106.500 162.740 ;
        RECT 109.060 162.680 109.320 163.000 ;
        RECT 105.840 159.960 106.100 160.280 ;
        RECT 105.900 158.580 106.040 159.960 ;
        RECT 105.840 158.260 106.100 158.580 ;
        RECT 105.840 157.240 106.100 157.560 ;
        RECT 105.900 155.260 106.040 157.240 ;
        RECT 106.360 155.860 106.500 162.600 ;
        RECT 106.880 162.145 108.760 162.515 ;
        RECT 109.120 158.240 109.260 162.680 ;
        RECT 109.060 157.920 109.320 158.240 ;
        RECT 106.880 156.705 108.760 157.075 ;
        RECT 106.300 155.540 106.560 155.860 ;
        RECT 108.600 155.540 108.860 155.860 ;
        RECT 105.900 155.120 106.500 155.260 ;
        RECT 105.840 152.140 106.100 152.460 ;
        RECT 105.900 150.420 106.040 152.140 ;
        RECT 105.380 150.100 105.640 150.420 ;
        RECT 105.840 150.100 106.100 150.420 ;
        RECT 106.360 147.700 106.500 155.120 ;
        RECT 108.660 152.800 108.800 155.540 ;
        RECT 107.680 152.655 107.940 152.800 ;
        RECT 108.600 152.710 108.860 152.800 ;
        RECT 107.670 152.285 107.950 152.655 ;
        RECT 108.600 152.570 109.260 152.710 ;
        RECT 108.600 152.480 108.860 152.570 ;
        RECT 106.880 151.265 108.760 151.635 ;
        RECT 109.120 151.100 109.260 152.570 ;
        RECT 109.060 150.780 109.320 151.100 ;
        RECT 109.060 148.060 109.320 148.380 ;
        RECT 106.300 147.380 106.560 147.700 ;
        RECT 106.300 146.700 106.560 147.020 ;
        RECT 104.920 144.320 105.180 144.640 ;
        RECT 106.360 144.380 106.500 146.700 ;
        RECT 106.880 145.825 108.760 146.195 ;
        RECT 106.360 144.300 106.960 144.380 ;
        RECT 106.360 144.240 107.020 144.300 ;
        RECT 106.760 143.980 107.020 144.240 ;
        RECT 105.380 143.640 105.640 143.960 ;
        RECT 106.300 143.640 106.560 143.960 ;
        RECT 104.920 140.920 105.180 141.240 ;
        RECT 104.980 138.520 105.120 140.920 ;
        RECT 104.920 138.200 105.180 138.520 ;
        RECT 104.920 135.480 105.180 135.800 ;
        RECT 104.980 134.100 105.120 135.480 ;
        RECT 104.920 133.780 105.180 134.100 ;
        RECT 105.440 132.060 105.580 143.640 ;
        RECT 105.840 141.940 106.100 142.260 ;
        RECT 105.900 137.500 106.040 141.940 ;
        RECT 105.840 137.180 106.100 137.500 ;
        RECT 104.000 131.740 104.260 132.060 ;
        RECT 105.380 131.740 105.640 132.060 ;
        RECT 103.540 128.340 103.800 128.660 ;
        RECT 103.600 126.135 103.740 128.340 ;
        RECT 103.530 125.765 103.810 126.135 ;
        RECT 103.540 122.900 103.800 123.220 ;
        RECT 103.600 121.180 103.740 122.900 ;
        RECT 105.840 121.880 106.100 122.200 ;
        RECT 103.540 120.860 103.800 121.180 ;
        RECT 105.900 120.160 106.040 121.880 ;
        RECT 105.840 119.840 106.100 120.160 ;
        RECT 105.840 119.160 106.100 119.480 ;
        RECT 105.900 117.440 106.040 119.160 ;
        RECT 105.840 117.120 106.100 117.440 ;
        RECT 104.000 116.440 104.260 116.760 ;
        RECT 104.060 114.380 104.200 116.440 ;
        RECT 104.000 114.060 104.260 114.380 ;
        RECT 104.920 109.640 105.180 109.960 ;
        RECT 103.080 108.960 103.340 109.280 ;
        RECT 100.320 108.620 100.580 108.940 ;
        RECT 99.400 108.340 99.660 108.600 ;
        RECT 100.380 108.340 100.520 108.620 ;
        RECT 99.400 108.280 100.520 108.340 ;
        RECT 99.460 108.200 100.520 108.280 ;
        RECT 98.940 103.860 99.200 104.180 ;
        RECT 100.380 103.840 100.520 108.200 ;
        RECT 104.000 106.240 104.260 106.560 ;
        RECT 100.320 103.520 100.580 103.840 ;
        RECT 104.060 89.170 104.200 106.240 ;
        RECT 104.980 104.180 105.120 109.640 ;
        RECT 106.360 109.280 106.500 143.640 ;
        RECT 106.880 140.385 108.760 140.755 ;
        RECT 107.220 139.560 107.480 139.880 ;
        RECT 107.280 137.500 107.420 139.560 ;
        RECT 107.220 137.180 107.480 137.500 ;
        RECT 106.880 134.945 108.760 135.315 ;
        RECT 107.220 133.780 107.480 134.100 ;
        RECT 107.280 131.040 107.420 133.780 ;
        RECT 109.120 132.060 109.260 148.060 ;
        RECT 109.580 147.360 109.720 170.840 ;
        RECT 110.040 166.740 110.180 171.520 ;
        RECT 110.440 171.180 110.700 171.500 ;
        RECT 110.500 168.440 110.640 171.180 ;
        RECT 112.340 169.120 112.480 171.860 ;
        RECT 114.180 170.140 114.320 171.860 ;
        RECT 114.120 169.820 114.380 170.140 ;
        RECT 110.900 168.800 111.160 169.120 ;
        RECT 112.280 168.800 112.540 169.120 ;
        RECT 110.440 168.120 110.700 168.440 ;
        RECT 110.500 166.740 110.640 168.120 ;
        RECT 109.980 166.420 110.240 166.740 ;
        RECT 110.440 166.420 110.700 166.740 ;
        RECT 110.960 166.650 111.100 168.800 ;
        RECT 111.360 166.650 111.620 166.740 ;
        RECT 110.960 166.510 111.620 166.650 ;
        RECT 111.360 166.420 111.620 166.510 ;
        RECT 110.040 163.680 110.180 166.420 ;
        RECT 110.440 165.400 110.700 165.720 ;
        RECT 109.980 163.360 110.240 163.680 ;
        RECT 109.980 158.940 110.240 159.260 ;
        RECT 109.520 147.040 109.780 147.360 ;
        RECT 110.040 146.420 110.180 158.940 ;
        RECT 109.580 146.280 110.180 146.420 ;
        RECT 109.580 134.780 109.720 146.280 ;
        RECT 110.500 145.320 110.640 165.400 ;
        RECT 111.420 164.360 111.560 166.420 ;
        RECT 112.280 164.380 112.540 164.700 ;
        RECT 111.360 164.040 111.620 164.360 ;
        RECT 112.340 163.680 112.480 164.380 ;
        RECT 114.640 163.680 114.780 179.000 ;
        RECT 116.020 178.300 116.160 179.340 ;
        RECT 116.940 179.320 117.080 182.740 ;
        RECT 117.400 182.720 117.540 187.160 ;
        RECT 121.880 186.625 123.760 186.995 ;
        RECT 124.300 186.460 124.440 187.160 ;
        RECT 124.240 186.140 124.500 186.460 ;
        RECT 125.680 185.780 125.820 187.840 ;
        RECT 125.620 185.460 125.880 185.780 ;
        RECT 124.240 185.120 124.500 185.440 ;
        RECT 122.400 184.780 122.660 185.100 ;
        RECT 118.720 184.440 118.980 184.760 ;
        RECT 118.780 183.740 118.920 184.440 ;
        RECT 122.460 183.740 122.600 184.780 ;
        RECT 118.720 183.420 118.980 183.740 ;
        RECT 122.400 183.420 122.660 183.740 ;
        RECT 119.640 182.740 119.900 183.060 ;
        RECT 117.340 182.400 117.600 182.720 ;
        RECT 116.880 179.000 117.140 179.320 ;
        RECT 115.960 177.980 116.220 178.300 ;
        RECT 115.960 177.300 116.220 177.620 ;
        RECT 116.020 174.900 116.160 177.300 ;
        RECT 115.960 174.580 116.220 174.900 ;
        RECT 116.020 169.800 116.160 174.580 ;
        RECT 117.400 174.560 117.540 182.400 ;
        RECT 118.260 182.060 118.520 182.380 ;
        RECT 118.320 180.340 118.460 182.060 ;
        RECT 119.700 181.020 119.840 182.740 ;
        RECT 121.880 181.185 123.760 181.555 ;
        RECT 119.640 180.700 119.900 181.020 ;
        RECT 118.260 180.020 118.520 180.340 ;
        RECT 118.320 177.620 118.460 180.020 ;
        RECT 124.300 179.660 124.440 185.120 ;
        RECT 124.240 179.340 124.500 179.660 ;
        RECT 118.260 177.300 118.520 177.620 ;
        RECT 121.880 175.745 123.760 176.115 ;
        RECT 118.720 174.580 118.980 174.900 ;
        RECT 117.340 174.240 117.600 174.560 ;
        RECT 116.880 173.560 117.140 173.880 ;
        RECT 116.940 171.500 117.080 173.560 ;
        RECT 117.400 172.520 117.540 174.240 ;
        RECT 117.340 172.200 117.600 172.520 ;
        RECT 118.780 172.180 118.920 174.580 ;
        RECT 124.300 174.220 124.440 179.340 ;
        RECT 124.240 173.900 124.500 174.220 ;
        RECT 122.860 173.560 123.120 173.880 ;
        RECT 119.640 172.540 119.900 172.860 ;
        RECT 118.720 171.860 118.980 172.180 ;
        RECT 116.880 171.180 117.140 171.500 ;
        RECT 116.420 170.840 116.680 171.160 ;
        RECT 115.960 169.480 116.220 169.800 ;
        RECT 116.480 169.460 116.620 170.840 ;
        RECT 116.420 169.140 116.680 169.460 ;
        RECT 116.880 168.460 117.140 168.780 ;
        RECT 116.940 167.080 117.080 168.460 ;
        RECT 119.700 168.440 119.840 172.540 ;
        RECT 122.920 172.520 123.060 173.560 ;
        RECT 122.860 172.200 123.120 172.520 ;
        RECT 124.300 171.840 124.440 173.900 ;
        RECT 135.630 173.380 136.780 174.600 ;
        RECT 124.240 171.520 124.500 171.840 ;
        RECT 121.880 170.305 123.760 170.675 ;
        RECT 124.300 169.120 124.440 171.520 ;
        RECT 130.210 171.325 130.490 171.695 ;
        RECT 130.280 169.120 130.420 171.325 ;
        RECT 133.970 170.540 134.710 172.220 ;
        RECT 124.240 168.800 124.500 169.120 ;
        RECT 130.220 168.800 130.480 169.120 ;
        RECT 119.640 168.120 119.900 168.440 ;
        RECT 116.880 166.760 117.140 167.080 ;
        RECT 119.700 166.740 119.840 168.120 ;
        RECT 118.720 166.420 118.980 166.740 ;
        RECT 119.640 166.420 119.900 166.740 ;
        RECT 112.280 163.360 112.540 163.680 ;
        RECT 114.580 163.360 114.840 163.680 ;
        RECT 110.900 162.680 111.160 163.000 ;
        RECT 110.960 150.420 111.100 162.680 ;
        RECT 118.780 161.300 118.920 166.420 ;
        RECT 115.500 160.980 115.760 161.300 ;
        RECT 118.720 160.980 118.980 161.300 ;
        RECT 113.200 158.260 113.460 158.580 ;
        RECT 112.280 157.920 112.540 158.240 ;
        RECT 111.820 157.240 112.080 157.560 ;
        RECT 111.880 156.540 112.020 157.240 ;
        RECT 111.820 156.220 112.080 156.540 ;
        RECT 112.340 152.800 112.480 157.920 ;
        RECT 112.740 155.200 113.000 155.520 ;
        RECT 112.800 153.480 112.940 155.200 ;
        RECT 112.740 153.160 113.000 153.480 ;
        RECT 111.360 152.480 111.620 152.800 ;
        RECT 112.280 152.480 112.540 152.800 ;
        RECT 110.900 150.100 111.160 150.420 ;
        RECT 111.420 150.080 111.560 152.480 ;
        RECT 111.360 149.820 111.620 150.080 ;
        RECT 110.960 149.760 111.620 149.820 ;
        RECT 110.960 149.680 111.560 149.760 ;
        RECT 110.440 145.000 110.700 145.320 ;
        RECT 110.960 144.980 111.100 149.680 ;
        RECT 111.820 149.080 112.080 149.400 ;
        RECT 111.360 146.360 111.620 146.680 ;
        RECT 109.980 144.660 110.240 144.980 ;
        RECT 110.900 144.660 111.160 144.980 ;
        RECT 110.040 142.600 110.180 144.660 ;
        RECT 109.980 142.280 110.240 142.600 ;
        RECT 109.980 140.920 110.240 141.240 ;
        RECT 110.040 136.480 110.180 140.920 ;
        RECT 110.900 138.880 111.160 139.200 ;
        RECT 110.960 137.500 111.100 138.880 ;
        RECT 110.900 137.180 111.160 137.500 ;
        RECT 109.980 136.160 110.240 136.480 ;
        RECT 109.520 134.460 109.780 134.780 ;
        RECT 109.060 131.740 109.320 132.060 ;
        RECT 109.980 131.060 110.240 131.380 ;
        RECT 107.220 130.720 107.480 131.040 ;
        RECT 109.060 130.720 109.320 131.040 ;
        RECT 106.880 129.505 108.760 129.875 ;
        RECT 109.120 124.920 109.260 130.720 ;
        RECT 109.520 130.380 109.780 130.700 ;
        RECT 109.060 124.600 109.320 124.920 ;
        RECT 106.880 124.065 108.760 124.435 ;
        RECT 109.120 123.900 109.260 124.600 ;
        RECT 109.060 123.580 109.320 123.900 ;
        RECT 108.600 122.560 108.860 122.880 ;
        RECT 108.660 119.480 108.800 122.560 ;
        RECT 108.600 119.160 108.860 119.480 ;
        RECT 106.880 118.625 108.760 118.995 ;
        RECT 109.580 118.460 109.720 130.380 ;
        RECT 110.040 122.880 110.180 131.060 ;
        RECT 109.980 122.560 110.240 122.880 ;
        RECT 106.760 118.140 107.020 118.460 ;
        RECT 109.520 118.140 109.780 118.460 ;
        RECT 106.820 115.740 106.960 118.140 ;
        RECT 109.520 116.440 109.780 116.760 ;
        RECT 106.760 115.420 107.020 115.740 ;
        RECT 106.880 113.185 108.760 113.555 ;
        RECT 109.580 112.340 109.720 116.440 ;
        RECT 109.520 112.020 109.780 112.340 ;
        RECT 111.420 109.280 111.560 146.360 ;
        RECT 111.880 134.780 112.020 149.080 ;
        RECT 112.340 147.360 112.480 152.480 ;
        RECT 112.800 148.040 112.940 153.160 ;
        RECT 113.260 152.460 113.400 158.260 ;
        RECT 113.660 157.920 113.920 158.240 ;
        RECT 113.200 152.140 113.460 152.460 ;
        RECT 112.740 147.720 113.000 148.040 ;
        RECT 112.280 147.040 112.540 147.360 ;
        RECT 112.340 144.300 112.480 147.040 ;
        RECT 112.280 143.980 112.540 144.300 ;
        RECT 112.800 142.940 112.940 147.720 ;
        RECT 113.260 147.700 113.400 152.140 ;
        RECT 113.720 150.080 113.860 157.920 ;
        RECT 115.560 155.860 115.700 160.980 ;
        RECT 119.180 159.960 119.440 160.280 ;
        RECT 119.240 157.900 119.380 159.960 ;
        RECT 119.180 157.580 119.440 157.900 ;
        RECT 118.260 157.240 118.520 157.560 ;
        RECT 115.500 155.540 115.760 155.860 ;
        RECT 114.120 151.800 114.380 152.120 ;
        RECT 114.180 150.760 114.320 151.800 ;
        RECT 114.580 150.780 114.840 151.100 ;
        RECT 114.120 150.440 114.380 150.760 ;
        RECT 113.660 149.760 113.920 150.080 ;
        RECT 113.200 147.380 113.460 147.700 ;
        RECT 113.720 147.360 113.860 149.760 ;
        RECT 113.660 147.040 113.920 147.360 ;
        RECT 113.660 144.660 113.920 144.980 ;
        RECT 112.740 142.850 113.000 142.940 ;
        RECT 112.740 142.710 113.400 142.850 ;
        RECT 112.740 142.620 113.000 142.710 ;
        RECT 112.740 141.940 113.000 142.260 ;
        RECT 112.800 139.200 112.940 141.940 ;
        RECT 113.260 139.200 113.400 142.710 ;
        RECT 112.740 138.880 113.000 139.200 ;
        RECT 113.200 138.880 113.460 139.200 ;
        RECT 112.800 134.780 112.940 138.880 ;
        RECT 113.720 136.140 113.860 144.660 ;
        RECT 113.660 135.820 113.920 136.140 ;
        RECT 111.820 134.460 112.080 134.780 ;
        RECT 112.740 134.460 113.000 134.780 ;
        RECT 112.280 133.780 112.540 134.100 ;
        RECT 112.340 131.720 112.480 133.780 ;
        RECT 112.280 131.400 112.540 131.720 ;
        RECT 111.820 130.040 112.080 130.360 ;
        RECT 111.880 124.920 112.020 130.040 ;
        RECT 112.800 129.000 112.940 134.460 ;
        RECT 113.200 133.440 113.460 133.760 ;
        RECT 113.260 131.040 113.400 133.440 ;
        RECT 113.200 130.720 113.460 131.040 ;
        RECT 112.740 128.680 113.000 129.000 ;
        RECT 112.800 125.600 112.940 128.680 ;
        RECT 113.200 128.570 113.460 128.660 ;
        RECT 113.720 128.570 113.860 135.820 ;
        RECT 113.200 128.430 113.860 128.570 ;
        RECT 113.200 128.340 113.460 128.430 ;
        RECT 112.740 125.280 113.000 125.600 ;
        RECT 111.820 124.600 112.080 124.920 ;
        RECT 112.800 123.220 112.940 125.280 ;
        RECT 112.740 122.900 113.000 123.220 ;
        RECT 113.260 120.160 113.400 128.340 ;
        RECT 113.200 119.840 113.460 120.160 ;
        RECT 114.120 119.500 114.380 119.820 ;
        RECT 114.180 118.460 114.320 119.500 ;
        RECT 114.120 118.140 114.380 118.460 ;
        RECT 111.820 114.400 112.080 114.720 ;
        RECT 111.880 113.020 112.020 114.400 ;
        RECT 111.820 112.700 112.080 113.020 ;
        RECT 114.640 109.280 114.780 150.780 ;
        RECT 115.560 144.980 115.700 155.540 ;
        RECT 117.800 154.860 118.060 155.180 ;
        RECT 117.860 153.820 118.000 154.860 ;
        RECT 117.800 153.500 118.060 153.820 ;
        RECT 117.860 151.860 118.000 153.500 ;
        RECT 118.320 152.800 118.460 157.240 ;
        RECT 118.720 154.520 118.980 154.840 ;
        RECT 118.780 152.800 118.920 154.520 ;
        RECT 118.260 152.480 118.520 152.800 ;
        RECT 118.720 152.480 118.980 152.800 ;
        RECT 118.260 151.860 118.520 152.120 ;
        RECT 117.860 151.800 118.520 151.860 ;
        RECT 117.860 151.720 118.460 151.800 ;
        RECT 118.320 147.360 118.460 151.720 ;
        RECT 118.260 147.040 118.520 147.360 ;
        RECT 117.340 146.360 117.600 146.680 ;
        RECT 117.400 144.980 117.540 146.360 ;
        RECT 115.500 144.660 115.760 144.980 ;
        RECT 117.340 144.660 117.600 144.980 ;
        RECT 115.560 141.920 115.700 144.660 ;
        RECT 116.880 142.280 117.140 142.600 ;
        RECT 115.500 141.600 115.760 141.920 ;
        RECT 116.940 140.220 117.080 142.280 ;
        RECT 117.400 140.220 117.540 144.660 ;
        RECT 119.700 144.640 119.840 166.420 ;
        RECT 124.300 166.400 124.440 168.800 ;
        RECT 135.630 166.640 136.740 173.380 ;
        RECT 124.240 166.080 124.500 166.400 ;
        RECT 121.880 164.865 123.760 165.235 ;
        RECT 121.880 159.425 123.760 159.795 ;
        RECT 120.100 158.260 120.360 158.580 ;
        RECT 119.640 144.320 119.900 144.640 ;
        RECT 116.880 139.900 117.140 140.220 ;
        RECT 117.340 139.900 117.600 140.220 ;
        RECT 116.880 133.440 117.140 133.760 ;
        RECT 115.960 131.400 116.220 131.720 ;
        RECT 115.500 127.320 115.760 127.640 ;
        RECT 115.560 125.260 115.700 127.320 ;
        RECT 115.500 124.940 115.760 125.260 ;
        RECT 116.020 118.460 116.160 131.400 ;
        RECT 116.940 130.360 117.080 133.440 ;
        RECT 117.340 130.720 117.600 131.040 ;
        RECT 116.880 130.040 117.140 130.360 ;
        RECT 116.940 129.340 117.080 130.040 ;
        RECT 116.880 129.020 117.140 129.340 ;
        RECT 116.940 123.900 117.080 129.020 ;
        RECT 117.400 125.940 117.540 130.720 ;
        RECT 119.180 130.040 119.440 130.360 ;
        RECT 117.340 125.620 117.600 125.940 ;
        RECT 117.400 123.900 117.540 125.620 ;
        RECT 119.240 124.920 119.380 130.040 ;
        RECT 119.180 124.600 119.440 124.920 ;
        RECT 116.880 123.580 117.140 123.900 ;
        RECT 117.340 123.580 117.600 123.900 ;
        RECT 118.720 119.160 118.980 119.480 ;
        RECT 115.960 118.140 116.220 118.460 ;
        RECT 118.780 118.120 118.920 119.160 ;
        RECT 118.720 117.800 118.980 118.120 ;
        RECT 117.340 112.360 117.600 112.680 ;
        RECT 117.400 109.620 117.540 112.360 ;
        RECT 120.160 112.340 120.300 158.260 ;
        RECT 124.300 158.240 124.440 166.080 ;
        RECT 135.630 165.420 136.780 166.640 ;
        RECT 124.240 157.920 124.500 158.240 ;
        RECT 126.080 157.920 126.340 158.240 ;
        RECT 121.480 157.580 121.740 157.900 ;
        RECT 121.540 153.820 121.680 157.580 ;
        RECT 126.140 155.860 126.280 157.920 ;
        RECT 126.080 155.540 126.340 155.860 ;
        RECT 124.240 155.200 124.500 155.520 ;
        RECT 121.880 153.985 123.760 154.355 ;
        RECT 124.300 153.820 124.440 155.200 ;
        RECT 121.480 153.500 121.740 153.820 ;
        RECT 124.240 153.500 124.500 153.820 ;
        RECT 121.020 149.420 121.280 149.740 ;
        RECT 121.080 112.340 121.220 149.420 ;
        RECT 121.880 148.545 123.760 148.915 ;
        RECT 124.240 146.360 124.500 146.680 ;
        RECT 124.300 144.980 124.440 146.360 ;
        RECT 124.240 144.660 124.500 144.980 ;
        RECT 126.080 144.320 126.340 144.640 ;
        RECT 121.880 143.105 123.760 143.475 ;
        RECT 122.400 141.940 122.660 142.260 ;
        RECT 122.460 140.220 122.600 141.940 ;
        RECT 126.140 141.920 126.280 144.320 ;
        RECT 126.080 141.600 126.340 141.920 ;
        RECT 135.630 141.200 136.780 141.270 ;
        RECT 122.400 139.900 122.660 140.220 ;
        RECT 135.630 140.180 136.800 141.200 ;
        RECT 129.140 138.175 134.100 139.455 ;
        RECT 121.880 137.665 123.760 138.035 ;
        RECT 135.640 133.320 136.800 140.180 ;
        RECT 121.880 132.225 123.760 132.595 ;
        RECT 125.160 128.340 125.420 128.660 ;
        RECT 124.240 128.000 124.500 128.320 ;
        RECT 121.880 126.785 123.760 127.155 ;
        RECT 122.860 125.620 123.120 125.940 ;
        RECT 122.920 123.900 123.060 125.620 ;
        RECT 124.300 125.600 124.440 128.000 ;
        RECT 125.220 126.620 125.360 128.340 ;
        RECT 125.160 126.300 125.420 126.620 ;
        RECT 124.240 125.280 124.500 125.600 ;
        RECT 122.860 123.580 123.120 123.900 ;
        RECT 121.880 121.345 123.760 121.715 ;
        RECT 122.400 119.160 122.660 119.480 ;
        RECT 122.460 117.780 122.600 119.160 ;
        RECT 122.400 117.460 122.660 117.780 ;
        RECT 124.300 117.440 124.440 125.280 ;
        RECT 124.240 117.120 124.500 117.440 ;
        RECT 121.880 115.905 123.760 116.275 ;
        RECT 124.300 115.060 124.440 117.120 ;
        RECT 124.240 114.740 124.500 115.060 ;
        RECT 118.720 112.020 118.980 112.340 ;
        RECT 120.100 112.020 120.360 112.340 ;
        RECT 121.020 112.020 121.280 112.340 ;
        RECT 117.340 109.300 117.600 109.620 ;
        RECT 106.300 108.960 106.560 109.280 ;
        RECT 111.360 108.960 111.620 109.280 ;
        RECT 114.580 108.960 114.840 109.280 ;
        RECT 112.740 108.620 113.000 108.940 ;
        RECT 105.380 108.280 105.640 108.600 ;
        RECT 109.060 108.280 109.320 108.600 ;
        RECT 105.440 107.240 105.580 108.280 ;
        RECT 106.880 107.745 108.760 108.115 ;
        RECT 109.120 107.240 109.260 108.280 ;
        RECT 105.380 106.920 105.640 107.240 ;
        RECT 109.060 106.920 109.320 107.240 ;
        RECT 112.800 106.900 112.940 108.620 ;
        RECT 115.500 108.280 115.760 108.600 ;
        RECT 112.740 106.580 113.000 106.900 ;
        RECT 111.360 105.560 111.620 105.880 ;
        RECT 104.920 103.860 105.180 104.180 ;
        RECT 109.980 103.860 110.240 104.180 ;
        RECT 106.880 102.305 108.760 102.675 ;
        RECT 110.040 89.290 110.180 103.860 ;
        RECT 111.420 103.500 111.560 105.560 ;
        RECT 115.560 104.180 115.700 108.280 ;
        RECT 118.780 106.980 118.920 112.020 ;
        RECT 119.640 111.680 119.900 112.000 ;
        RECT 119.700 108.940 119.840 111.680 ;
        RECT 121.880 110.465 123.760 110.835 ;
        RECT 124.300 110.300 124.440 114.740 ;
        RECT 124.700 111.000 124.960 111.320 ;
        RECT 124.240 109.980 124.500 110.300 ;
        RECT 119.640 108.620 119.900 108.940 ;
        RECT 120.560 107.260 120.820 107.580 ;
        RECT 118.320 106.900 118.920 106.980 ;
        RECT 118.260 106.840 118.920 106.900 ;
        RECT 118.260 106.580 118.520 106.840 ;
        RECT 116.420 105.560 116.680 105.880 ;
        RECT 115.500 103.860 115.760 104.180 ;
        RECT 116.480 103.500 116.620 105.560 ;
        RECT 111.360 103.180 111.620 103.500 ;
        RECT 115.960 103.180 116.220 103.500 ;
        RECT 116.420 103.180 116.680 103.500 ;
        RECT 116.020 89.570 116.160 103.180 ;
        RECT 118.780 101.460 118.920 106.840 ;
        RECT 119.180 106.580 119.440 106.900 ;
        RECT 119.240 102.140 119.380 106.580 ;
        RECT 119.180 101.820 119.440 102.140 ;
        RECT 118.720 101.140 118.980 101.460 ;
        RECT 92.030 88.480 94.080 88.620 ;
        RECT 98.010 88.500 98.290 89.170 ;
        RECT 103.990 88.610 104.270 89.170 ;
        RECT 92.030 88.320 92.310 88.480 ;
        RECT 74.090 80.440 74.370 84.290 ;
        RECT 20.140 80.160 74.370 80.440 ;
        RECT 20.140 75.650 20.420 80.160 ;
        RECT 80.070 79.800 80.350 84.310 ;
        RECT 85.470 84.100 86.690 87.970 ;
        RECT 91.460 84.500 92.680 88.320 ;
        RECT 97.600 84.630 98.820 88.500 ;
        RECT 103.650 84.740 104.870 88.610 ;
        RECT 109.620 85.420 110.840 89.290 ;
        RECT 115.740 85.700 116.960 89.570 ;
        RECT 120.620 88.620 120.760 107.260 ;
        RECT 124.300 106.560 124.440 109.980 ;
        RECT 124.760 107.240 124.900 111.000 ;
        RECT 127.920 108.620 128.180 108.940 ;
        RECT 124.700 106.920 124.960 107.240 ;
        RECT 124.240 106.240 124.500 106.560 ;
        RECT 121.880 105.025 123.760 105.395 ;
        RECT 124.300 104.180 124.440 106.240 ;
        RECT 126.070 106.045 126.350 106.415 ;
        RECT 124.240 103.860 124.500 104.180 ;
        RECT 126.140 103.840 126.280 106.045 ;
        RECT 126.080 103.520 126.340 103.840 ;
        RECT 125.160 102.840 125.420 103.160 ;
        RECT 125.220 101.800 125.360 102.840 ;
        RECT 125.160 101.480 125.420 101.800 ;
        RECT 121.880 99.585 123.760 99.955 ;
        RECT 121.520 88.620 122.740 89.570 ;
        RECT 127.980 89.380 128.120 108.620 ;
        RECT 129.750 105.580 133.160 106.650 ;
        RECT 120.620 88.480 122.740 88.620 ;
        RECT 121.520 85.700 122.740 88.480 ;
        RECT 31.380 79.520 80.350 79.800 ;
        RECT 31.380 75.850 31.660 79.520 ;
        RECT 86.050 79.170 86.330 84.100 ;
        RECT 42.510 78.890 86.330 79.170 ;
        RECT 3.960 71.320 6.050 73.240 ;
        RECT 19.330 73.120 21.890 75.650 ;
        RECT 28.185 73.180 30.255 74.460 ;
        RECT 30.670 73.320 33.230 75.850 ;
        RECT 42.510 75.750 42.790 78.890 ;
        RECT 92.030 78.570 92.310 84.500 ;
        RECT 53.830 78.290 92.310 78.570 ;
        RECT 53.830 75.820 54.110 78.290 ;
        RECT 98.010 77.990 98.290 84.630 ;
        RECT 64.900 77.710 98.290 77.990 ;
        RECT 19.005 71.800 19.865 72.640 ;
        RECT 15.560 68.610 16.990 71.210 ;
        RECT 19.305 68.570 19.845 71.800 ;
        RECT 20.145 70.600 20.555 73.120 ;
        RECT 30.205 71.810 31.065 72.650 ;
        RECT 19.325 47.770 19.825 68.570 ;
        RECT 20.165 49.090 20.555 70.600 ;
        RECT 20.955 70.010 21.845 70.740 ;
        RECT 21.055 65.190 21.315 70.010 ;
        RECT 22.695 68.620 25.405 69.470 ;
        RECT 22.895 65.840 24.825 68.620 ;
        RECT 30.505 68.580 31.045 71.810 ;
        RECT 31.345 70.610 31.755 73.320 ;
        RECT 39.475 73.150 41.545 74.430 ;
        RECT 41.910 73.220 44.470 75.750 ;
        RECT 41.425 71.780 42.285 72.620 ;
        RECT 27.795 67.130 28.915 67.810 ;
        RECT 28.075 65.850 28.745 67.130 ;
        RECT 21.455 65.460 26.505 65.840 ;
        RECT 27.865 65.440 28.915 65.850 ;
        RECT 21.055 63.640 21.435 65.190 ;
        RECT 21.175 55.800 21.435 63.640 ;
        RECT 26.485 63.200 26.755 65.240 ;
        RECT 27.615 63.200 27.885 65.200 ;
        RECT 26.485 56.510 27.885 63.200 ;
        RECT 21.085 55.290 21.445 55.800 ;
        RECT 21.065 54.860 21.445 55.290 ;
        RECT 26.485 55.190 26.755 56.510 ;
        RECT 27.615 55.150 27.885 56.510 ;
        RECT 28.885 55.260 29.205 65.190 ;
        RECT 28.885 55.200 29.215 55.260 ;
        RECT 21.065 54.580 21.315 54.860 ;
        RECT 20.865 54.180 25.505 54.580 ;
        RECT 26.405 54.290 27.535 54.300 ;
        RECT 28.895 54.290 29.215 55.200 ;
        RECT 21.065 52.060 21.315 54.180 ;
        RECT 25.765 53.490 26.125 54.110 ;
        RECT 25.845 52.610 26.105 53.490 ;
        RECT 26.385 53.240 29.215 54.290 ;
        RECT 25.675 52.230 26.205 52.610 ;
        RECT 21.065 51.970 21.565 52.060 ;
        RECT 21.055 51.240 21.565 51.970 ;
        RECT 21.295 50.240 21.565 51.240 ;
        RECT 22.205 50.990 22.475 51.940 ;
        RECT 22.205 50.840 22.675 50.990 ;
        RECT 22.205 50.160 22.765 50.840 ;
        RECT 22.285 50.150 22.765 50.160 ;
        RECT 21.575 49.620 22.195 49.980 ;
        RECT 21.615 49.090 22.045 49.620 ;
        RECT 20.165 48.670 22.045 49.090 ;
        RECT 22.535 48.960 22.765 50.150 ;
        RECT 21.615 47.800 22.045 48.670 ;
        RECT 22.455 48.360 22.835 48.960 ;
        RECT 19.325 47.060 20.015 47.770 ;
        RECT 21.435 47.440 22.055 47.800 ;
        RECT 21.135 47.060 21.425 47.250 ;
        RECT 19.325 46.620 21.425 47.060 ;
        RECT 19.325 46.600 20.015 46.620 ;
        RECT 21.135 46.380 21.425 46.620 ;
        RECT 22.055 46.990 22.325 47.240 ;
        RECT 22.535 46.990 22.765 48.360 ;
        RECT 25.355 47.010 25.685 52.030 ;
        RECT 26.405 52.020 27.535 53.240 ;
        RECT 28.895 53.220 29.215 53.240 ;
        RECT 22.055 46.880 22.765 46.990 ;
        RECT 25.345 46.960 25.685 47.010 ;
        RECT 26.235 47.780 27.615 52.020 ;
        RECT 22.055 46.570 22.715 46.880 ;
        RECT 22.055 46.400 22.325 46.570 ;
        RECT 25.345 45.000 25.625 46.960 ;
        RECT 26.235 46.920 26.535 47.780 ;
        RECT 27.315 46.920 27.615 47.780 ;
        RECT 28.165 46.920 28.495 51.990 ;
        RECT 27.565 46.380 28.045 46.760 ;
        RECT 27.665 45.760 27.915 46.380 ;
        RECT 27.565 45.160 27.945 45.760 ;
        RECT 24.825 44.230 25.925 45.000 ;
        RECT 28.215 44.930 28.495 46.920 ;
        RECT 30.525 47.780 31.025 68.580 ;
        RECT 31.365 49.100 31.755 70.610 ;
        RECT 32.155 70.020 33.045 70.750 ;
        RECT 32.255 65.200 32.515 70.020 ;
        RECT 33.895 68.630 36.605 69.480 ;
        RECT 34.095 65.850 36.025 68.630 ;
        RECT 41.725 68.550 42.265 71.780 ;
        RECT 42.565 70.580 42.975 73.220 ;
        RECT 50.055 73.090 52.125 74.370 ;
        RECT 53.150 73.290 55.710 75.820 ;
        RECT 64.900 75.810 65.180 77.710 ;
        RECT 103.990 77.230 104.270 84.740 ;
        RECT 76.140 76.950 104.270 77.230 ;
        RECT 52.675 71.760 53.535 72.600 ;
        RECT 38.995 67.140 40.115 67.820 ;
        RECT 39.275 65.860 39.945 67.140 ;
        RECT 32.655 65.470 37.705 65.850 ;
        RECT 39.065 65.450 40.115 65.860 ;
        RECT 32.255 63.650 32.635 65.200 ;
        RECT 32.375 55.810 32.635 63.650 ;
        RECT 37.685 63.210 37.955 65.250 ;
        RECT 38.815 63.210 39.085 65.210 ;
        RECT 37.685 56.520 39.085 63.210 ;
        RECT 32.285 55.300 32.645 55.810 ;
        RECT 32.265 54.870 32.645 55.300 ;
        RECT 37.685 55.200 37.955 56.520 ;
        RECT 38.815 55.160 39.085 56.520 ;
        RECT 40.085 55.270 40.405 65.200 ;
        RECT 40.085 55.210 40.415 55.270 ;
        RECT 32.265 54.590 32.515 54.870 ;
        RECT 32.065 54.190 36.705 54.590 ;
        RECT 37.605 54.300 38.735 54.310 ;
        RECT 40.095 54.300 40.415 55.210 ;
        RECT 32.265 52.070 32.515 54.190 ;
        RECT 36.965 53.500 37.325 54.120 ;
        RECT 37.045 52.620 37.305 53.500 ;
        RECT 37.585 53.250 40.415 54.300 ;
        RECT 36.875 52.240 37.405 52.620 ;
        RECT 32.265 51.980 32.765 52.070 ;
        RECT 32.255 51.250 32.765 51.980 ;
        RECT 32.495 50.250 32.765 51.250 ;
        RECT 33.405 51.000 33.675 51.950 ;
        RECT 33.405 50.850 33.875 51.000 ;
        RECT 33.405 50.170 33.965 50.850 ;
        RECT 33.485 50.160 33.965 50.170 ;
        RECT 32.775 49.630 33.395 49.990 ;
        RECT 32.815 49.100 33.245 49.630 ;
        RECT 31.365 48.680 33.245 49.100 ;
        RECT 33.735 48.970 33.965 50.160 ;
        RECT 32.815 47.810 33.245 48.680 ;
        RECT 33.655 48.370 34.035 48.970 ;
        RECT 30.525 47.070 31.215 47.780 ;
        RECT 32.635 47.450 33.255 47.810 ;
        RECT 32.335 47.070 32.625 47.260 ;
        RECT 30.525 46.630 32.625 47.070 ;
        RECT 30.525 46.610 31.215 46.630 ;
        RECT 32.335 46.390 32.625 46.630 ;
        RECT 33.255 47.000 33.525 47.250 ;
        RECT 33.735 47.000 33.965 48.370 ;
        RECT 36.555 47.020 36.885 52.040 ;
        RECT 37.605 52.030 38.735 53.250 ;
        RECT 40.095 53.230 40.415 53.250 ;
        RECT 33.255 46.890 33.965 47.000 ;
        RECT 36.545 46.970 36.885 47.020 ;
        RECT 37.435 47.790 38.815 52.030 ;
        RECT 33.255 46.580 33.915 46.890 ;
        RECT 33.255 46.410 33.525 46.580 ;
        RECT 36.545 45.010 36.825 46.970 ;
        RECT 37.435 46.930 37.735 47.790 ;
        RECT 38.515 46.930 38.815 47.790 ;
        RECT 39.365 46.930 39.695 52.000 ;
        RECT 38.765 46.390 39.245 46.770 ;
        RECT 38.865 45.770 39.115 46.390 ;
        RECT 38.765 45.170 39.145 45.770 ;
        RECT 28.215 43.200 28.515 44.930 ;
        RECT 36.025 44.240 37.125 45.010 ;
        RECT 39.415 44.940 39.695 46.930 ;
        RECT 41.745 47.750 42.245 68.550 ;
        RECT 42.585 49.070 42.975 70.580 ;
        RECT 43.375 69.990 44.265 70.720 ;
        RECT 43.475 65.170 43.735 69.990 ;
        RECT 45.115 68.600 47.825 69.450 ;
        RECT 45.315 65.820 47.245 68.600 ;
        RECT 52.975 68.530 53.515 71.760 ;
        RECT 53.815 70.560 54.225 73.290 ;
        RECT 61.475 73.120 63.545 74.400 ;
        RECT 64.400 73.280 66.960 75.810 ;
        RECT 76.140 75.740 76.420 76.950 ;
        RECT 109.970 76.610 110.250 85.420 ;
        RECT 87.580 76.330 110.250 76.610 ;
        RECT 87.580 75.760 87.860 76.330 ;
        RECT 115.950 76.030 116.230 85.700 ;
        RECT 98.850 75.840 116.230 76.030 ;
        RECT 63.895 71.750 64.755 72.590 ;
        RECT 50.215 67.110 51.335 67.790 ;
        RECT 50.495 65.830 51.165 67.110 ;
        RECT 43.875 65.440 48.925 65.820 ;
        RECT 50.285 65.420 51.335 65.830 ;
        RECT 43.475 63.620 43.855 65.170 ;
        RECT 43.595 55.780 43.855 63.620 ;
        RECT 48.905 63.180 49.175 65.220 ;
        RECT 50.035 63.180 50.305 65.180 ;
        RECT 48.905 56.490 50.305 63.180 ;
        RECT 43.505 55.270 43.865 55.780 ;
        RECT 43.485 54.840 43.865 55.270 ;
        RECT 48.905 55.170 49.175 56.490 ;
        RECT 50.035 55.130 50.305 56.490 ;
        RECT 51.305 55.240 51.625 65.170 ;
        RECT 51.305 55.180 51.635 55.240 ;
        RECT 43.485 54.560 43.735 54.840 ;
        RECT 43.285 54.160 47.925 54.560 ;
        RECT 48.825 54.270 49.955 54.280 ;
        RECT 51.315 54.270 51.635 55.180 ;
        RECT 43.485 52.040 43.735 54.160 ;
        RECT 48.185 53.470 48.545 54.090 ;
        RECT 48.265 52.590 48.525 53.470 ;
        RECT 48.805 53.220 51.635 54.270 ;
        RECT 48.095 52.210 48.625 52.590 ;
        RECT 43.485 51.950 43.985 52.040 ;
        RECT 43.475 51.220 43.985 51.950 ;
        RECT 43.715 50.220 43.985 51.220 ;
        RECT 44.625 50.970 44.895 51.920 ;
        RECT 44.625 50.820 45.095 50.970 ;
        RECT 44.625 50.140 45.185 50.820 ;
        RECT 44.705 50.130 45.185 50.140 ;
        RECT 43.995 49.600 44.615 49.960 ;
        RECT 44.035 49.070 44.465 49.600 ;
        RECT 42.585 48.650 44.465 49.070 ;
        RECT 44.955 48.940 45.185 50.130 ;
        RECT 44.035 47.780 44.465 48.650 ;
        RECT 44.875 48.340 45.255 48.940 ;
        RECT 41.745 47.040 42.435 47.750 ;
        RECT 43.855 47.420 44.475 47.780 ;
        RECT 43.555 47.040 43.845 47.230 ;
        RECT 41.745 46.600 43.845 47.040 ;
        RECT 41.745 46.580 42.435 46.600 ;
        RECT 43.555 46.360 43.845 46.600 ;
        RECT 44.475 46.970 44.745 47.220 ;
        RECT 44.955 46.970 45.185 48.340 ;
        RECT 47.775 46.990 48.105 52.010 ;
        RECT 48.825 52.000 49.955 53.220 ;
        RECT 51.315 53.200 51.635 53.220 ;
        RECT 44.475 46.860 45.185 46.970 ;
        RECT 47.765 46.940 48.105 46.990 ;
        RECT 48.655 47.760 50.035 52.000 ;
        RECT 44.475 46.550 45.135 46.860 ;
        RECT 44.475 46.380 44.745 46.550 ;
        RECT 47.765 44.980 48.045 46.940 ;
        RECT 48.655 46.900 48.955 47.760 ;
        RECT 49.735 46.900 50.035 47.760 ;
        RECT 50.585 46.900 50.915 51.970 ;
        RECT 49.985 46.360 50.465 46.740 ;
        RECT 50.085 45.740 50.335 46.360 ;
        RECT 49.985 45.140 50.365 45.740 ;
        RECT 39.415 43.210 39.715 44.940 ;
        RECT 47.245 44.210 48.345 44.980 ;
        RECT 50.635 44.910 50.915 46.900 ;
        RECT 52.995 47.730 53.495 68.530 ;
        RECT 53.835 49.050 54.225 70.560 ;
        RECT 54.625 69.970 55.515 70.700 ;
        RECT 54.725 65.150 54.985 69.970 ;
        RECT 56.365 68.580 59.075 69.430 ;
        RECT 56.565 65.800 58.495 68.580 ;
        RECT 64.195 68.520 64.735 71.750 ;
        RECT 65.035 70.550 65.445 73.280 ;
        RECT 72.585 73.130 74.655 74.410 ;
        RECT 75.550 73.210 78.110 75.740 ;
        RECT 75.135 71.740 75.995 72.580 ;
        RECT 61.465 67.090 62.585 67.770 ;
        RECT 61.745 65.810 62.415 67.090 ;
        RECT 55.125 65.420 60.175 65.800 ;
        RECT 61.535 65.400 62.585 65.810 ;
        RECT 54.725 63.600 55.105 65.150 ;
        RECT 54.845 55.760 55.105 63.600 ;
        RECT 60.155 63.160 60.425 65.200 ;
        RECT 61.285 63.160 61.555 65.160 ;
        RECT 60.155 56.470 61.555 63.160 ;
        RECT 54.755 55.250 55.115 55.760 ;
        RECT 54.735 54.820 55.115 55.250 ;
        RECT 60.155 55.150 60.425 56.470 ;
        RECT 61.285 55.110 61.555 56.470 ;
        RECT 62.555 55.220 62.875 65.150 ;
        RECT 62.555 55.160 62.885 55.220 ;
        RECT 54.735 54.540 54.985 54.820 ;
        RECT 54.535 54.140 59.175 54.540 ;
        RECT 60.075 54.250 61.205 54.260 ;
        RECT 62.565 54.250 62.885 55.160 ;
        RECT 54.735 52.020 54.985 54.140 ;
        RECT 59.435 53.450 59.795 54.070 ;
        RECT 59.515 52.570 59.775 53.450 ;
        RECT 60.055 53.200 62.885 54.250 ;
        RECT 59.345 52.190 59.875 52.570 ;
        RECT 54.735 51.930 55.235 52.020 ;
        RECT 54.725 51.200 55.235 51.930 ;
        RECT 54.965 50.200 55.235 51.200 ;
        RECT 55.875 50.950 56.145 51.900 ;
        RECT 55.875 50.800 56.345 50.950 ;
        RECT 55.875 50.120 56.435 50.800 ;
        RECT 55.955 50.110 56.435 50.120 ;
        RECT 55.245 49.580 55.865 49.940 ;
        RECT 55.285 49.050 55.715 49.580 ;
        RECT 53.835 48.630 55.715 49.050 ;
        RECT 56.205 48.920 56.435 50.110 ;
        RECT 55.285 47.760 55.715 48.630 ;
        RECT 56.125 48.320 56.505 48.920 ;
        RECT 52.995 47.020 53.685 47.730 ;
        RECT 55.105 47.400 55.725 47.760 ;
        RECT 54.805 47.020 55.095 47.210 ;
        RECT 52.995 46.580 55.095 47.020 ;
        RECT 52.995 46.560 53.685 46.580 ;
        RECT 54.805 46.340 55.095 46.580 ;
        RECT 55.725 46.950 55.995 47.200 ;
        RECT 56.205 46.950 56.435 48.320 ;
        RECT 59.025 46.970 59.355 51.990 ;
        RECT 60.075 51.980 61.205 53.200 ;
        RECT 62.565 53.180 62.885 53.200 ;
        RECT 55.725 46.840 56.435 46.950 ;
        RECT 59.015 46.920 59.355 46.970 ;
        RECT 59.905 47.740 61.285 51.980 ;
        RECT 55.725 46.530 56.385 46.840 ;
        RECT 55.725 46.360 55.995 46.530 ;
        RECT 59.015 44.960 59.295 46.920 ;
        RECT 59.905 46.880 60.205 47.740 ;
        RECT 60.985 46.880 61.285 47.740 ;
        RECT 61.835 46.880 62.165 51.950 ;
        RECT 61.235 46.340 61.715 46.720 ;
        RECT 61.335 45.720 61.585 46.340 ;
        RECT 61.235 45.120 61.615 45.720 ;
        RECT 19.865 42.210 21.245 42.780 ;
        RECT 27.495 42.630 28.875 43.200 ;
        RECT 31.145 42.210 32.525 42.780 ;
        RECT 38.695 42.640 40.075 43.210 ;
        RECT 50.635 43.180 50.935 44.910 ;
        RECT 58.495 44.190 59.595 44.960 ;
        RECT 61.885 44.890 62.165 46.880 ;
        RECT 64.215 47.720 64.715 68.520 ;
        RECT 65.055 49.040 65.445 70.550 ;
        RECT 65.845 69.960 66.735 70.690 ;
        RECT 65.945 65.140 66.205 69.960 ;
        RECT 67.585 68.570 70.295 69.420 ;
        RECT 67.785 65.790 69.715 68.570 ;
        RECT 75.435 68.510 75.975 71.740 ;
        RECT 76.275 70.540 76.685 73.210 ;
        RECT 83.855 73.120 85.925 74.400 ;
        RECT 86.850 73.230 89.410 75.760 ;
        RECT 98.150 75.750 116.230 75.840 ;
        RECT 86.385 71.750 87.245 72.590 ;
        RECT 72.685 67.080 73.805 67.760 ;
        RECT 72.965 65.800 73.635 67.080 ;
        RECT 66.345 65.410 71.395 65.790 ;
        RECT 72.755 65.390 73.805 65.800 ;
        RECT 65.945 63.590 66.325 65.140 ;
        RECT 66.065 55.750 66.325 63.590 ;
        RECT 71.375 63.150 71.645 65.190 ;
        RECT 72.505 63.150 72.775 65.150 ;
        RECT 71.375 56.460 72.775 63.150 ;
        RECT 65.975 55.240 66.335 55.750 ;
        RECT 65.955 54.810 66.335 55.240 ;
        RECT 71.375 55.140 71.645 56.460 ;
        RECT 72.505 55.100 72.775 56.460 ;
        RECT 73.775 55.210 74.095 65.140 ;
        RECT 73.775 55.150 74.105 55.210 ;
        RECT 65.955 54.530 66.205 54.810 ;
        RECT 65.755 54.130 70.395 54.530 ;
        RECT 71.295 54.240 72.425 54.250 ;
        RECT 73.785 54.240 74.105 55.150 ;
        RECT 65.955 52.010 66.205 54.130 ;
        RECT 70.655 53.440 71.015 54.060 ;
        RECT 70.735 52.560 70.995 53.440 ;
        RECT 71.275 53.190 74.105 54.240 ;
        RECT 70.565 52.180 71.095 52.560 ;
        RECT 65.955 51.920 66.455 52.010 ;
        RECT 65.945 51.190 66.455 51.920 ;
        RECT 66.185 50.190 66.455 51.190 ;
        RECT 67.095 50.940 67.365 51.890 ;
        RECT 67.095 50.790 67.565 50.940 ;
        RECT 67.095 50.110 67.655 50.790 ;
        RECT 67.175 50.100 67.655 50.110 ;
        RECT 66.465 49.570 67.085 49.930 ;
        RECT 66.505 49.040 66.935 49.570 ;
        RECT 65.055 48.620 66.935 49.040 ;
        RECT 67.425 48.910 67.655 50.100 ;
        RECT 66.505 47.750 66.935 48.620 ;
        RECT 67.345 48.310 67.725 48.910 ;
        RECT 64.215 47.010 64.905 47.720 ;
        RECT 66.325 47.390 66.945 47.750 ;
        RECT 66.025 47.010 66.315 47.200 ;
        RECT 64.215 46.570 66.315 47.010 ;
        RECT 64.215 46.550 64.905 46.570 ;
        RECT 66.025 46.330 66.315 46.570 ;
        RECT 66.945 46.940 67.215 47.190 ;
        RECT 67.425 46.940 67.655 48.310 ;
        RECT 70.245 46.960 70.575 51.980 ;
        RECT 71.295 51.970 72.425 53.190 ;
        RECT 73.785 53.170 74.105 53.190 ;
        RECT 66.945 46.830 67.655 46.940 ;
        RECT 70.235 46.910 70.575 46.960 ;
        RECT 71.125 47.730 72.505 51.970 ;
        RECT 66.945 46.520 67.605 46.830 ;
        RECT 66.945 46.350 67.215 46.520 ;
        RECT 70.235 44.950 70.515 46.910 ;
        RECT 71.125 46.870 71.425 47.730 ;
        RECT 72.205 46.870 72.505 47.730 ;
        RECT 73.055 46.870 73.385 51.940 ;
        RECT 72.455 46.330 72.935 46.710 ;
        RECT 72.555 45.710 72.805 46.330 ;
        RECT 72.455 45.110 72.835 45.710 ;
        RECT 20.225 40.480 20.525 42.210 ;
        RECT 20.245 38.490 20.525 40.480 ;
        RECT 22.815 40.410 23.915 41.180 ;
        RECT 31.505 40.480 31.805 42.210 ;
        RECT 42.435 42.190 43.815 42.760 ;
        RECT 49.915 42.610 51.295 43.180 ;
        RECT 61.885 43.160 62.185 44.890 ;
        RECT 69.715 44.180 70.815 44.950 ;
        RECT 73.105 44.880 73.385 46.870 ;
        RECT 75.455 47.710 75.955 68.510 ;
        RECT 76.295 49.030 76.685 70.540 ;
        RECT 77.085 69.950 77.975 70.680 ;
        RECT 77.185 65.130 77.445 69.950 ;
        RECT 78.825 68.560 81.535 69.410 ;
        RECT 79.025 65.780 80.955 68.560 ;
        RECT 86.685 68.520 87.225 71.750 ;
        RECT 87.525 70.550 87.935 73.230 ;
        RECT 95.045 73.060 97.115 74.340 ;
        RECT 98.150 73.310 100.710 75.750 ;
        RECT 109.390 75.480 111.950 75.560 ;
        RECT 121.930 75.480 122.210 85.700 ;
        RECT 127.550 85.510 128.770 89.380 ;
        RECT 127.910 76.040 128.190 85.510 ;
        RECT 133.380 76.580 136.010 77.880 ;
        RECT 137.240 76.560 139.870 77.860 ;
        RECT 109.390 75.200 122.210 75.480 ;
        RECT 97.665 71.740 98.525 72.580 ;
        RECT 83.925 67.070 85.045 67.750 ;
        RECT 84.205 65.790 84.875 67.070 ;
        RECT 77.585 65.400 82.635 65.780 ;
        RECT 83.995 65.380 85.045 65.790 ;
        RECT 77.185 63.580 77.565 65.130 ;
        RECT 77.305 55.740 77.565 63.580 ;
        RECT 82.615 63.140 82.885 65.180 ;
        RECT 83.745 63.140 84.015 65.140 ;
        RECT 82.615 56.450 84.015 63.140 ;
        RECT 77.215 55.230 77.575 55.740 ;
        RECT 77.195 54.800 77.575 55.230 ;
        RECT 82.615 55.130 82.885 56.450 ;
        RECT 83.745 55.090 84.015 56.450 ;
        RECT 85.015 55.200 85.335 65.130 ;
        RECT 85.015 55.140 85.345 55.200 ;
        RECT 77.195 54.520 77.445 54.800 ;
        RECT 76.995 54.120 81.635 54.520 ;
        RECT 82.535 54.230 83.665 54.240 ;
        RECT 85.025 54.230 85.345 55.140 ;
        RECT 77.195 52.000 77.445 54.120 ;
        RECT 81.895 53.430 82.255 54.050 ;
        RECT 81.975 52.550 82.235 53.430 ;
        RECT 82.515 53.180 85.345 54.230 ;
        RECT 81.805 52.170 82.335 52.550 ;
        RECT 77.195 51.910 77.695 52.000 ;
        RECT 77.185 51.180 77.695 51.910 ;
        RECT 77.425 50.180 77.695 51.180 ;
        RECT 78.335 50.930 78.605 51.880 ;
        RECT 78.335 50.780 78.805 50.930 ;
        RECT 78.335 50.100 78.895 50.780 ;
        RECT 78.415 50.090 78.895 50.100 ;
        RECT 77.705 49.560 78.325 49.920 ;
        RECT 77.745 49.030 78.175 49.560 ;
        RECT 76.295 48.610 78.175 49.030 ;
        RECT 78.665 48.900 78.895 50.090 ;
        RECT 77.745 47.740 78.175 48.610 ;
        RECT 78.585 48.300 78.965 48.900 ;
        RECT 75.455 47.000 76.145 47.710 ;
        RECT 77.565 47.380 78.185 47.740 ;
        RECT 77.265 47.000 77.555 47.190 ;
        RECT 75.455 46.560 77.555 47.000 ;
        RECT 75.455 46.540 76.145 46.560 ;
        RECT 77.265 46.320 77.555 46.560 ;
        RECT 78.185 46.930 78.455 47.180 ;
        RECT 78.665 46.930 78.895 48.300 ;
        RECT 81.485 46.950 81.815 51.970 ;
        RECT 82.535 51.960 83.665 53.180 ;
        RECT 85.025 53.160 85.345 53.180 ;
        RECT 78.185 46.820 78.895 46.930 ;
        RECT 81.475 46.900 81.815 46.950 ;
        RECT 82.365 47.720 83.745 51.960 ;
        RECT 78.185 46.510 78.845 46.820 ;
        RECT 78.185 46.340 78.455 46.510 ;
        RECT 81.475 44.940 81.755 46.900 ;
        RECT 82.365 46.860 82.665 47.720 ;
        RECT 83.445 46.860 83.745 47.720 ;
        RECT 84.295 46.860 84.625 51.930 ;
        RECT 83.695 46.320 84.175 46.700 ;
        RECT 83.795 45.700 84.045 46.320 ;
        RECT 83.695 45.100 84.075 45.700 ;
        RECT 53.655 42.190 55.035 42.760 ;
        RECT 61.165 42.590 62.545 43.160 ;
        RECT 73.105 43.150 73.405 44.880 ;
        RECT 80.955 44.170 82.055 44.940 ;
        RECT 84.345 44.870 84.625 46.860 ;
        RECT 86.705 47.720 87.205 68.520 ;
        RECT 87.545 49.040 87.935 70.550 ;
        RECT 88.335 69.960 89.225 70.690 ;
        RECT 88.435 65.140 88.695 69.960 ;
        RECT 90.075 68.570 92.785 69.420 ;
        RECT 90.275 65.790 92.205 68.570 ;
        RECT 97.965 68.510 98.505 71.740 ;
        RECT 98.805 70.540 99.215 73.310 ;
        RECT 106.455 73.110 108.525 74.390 ;
        RECT 109.390 73.030 111.950 75.200 ;
        RECT 125.760 74.810 128.190 76.040 ;
        RECT 121.290 74.790 128.190 74.810 ;
        RECT 120.600 74.530 128.190 74.790 ;
        RECT 117.655 73.110 119.725 74.390 ;
        RECT 120.600 73.180 128.160 74.530 ;
        RECT 129.505 73.190 131.575 74.470 ;
        RECT 120.600 73.110 126.160 73.180 ;
        RECT 108.935 71.740 109.795 72.580 ;
        RECT 95.175 67.080 96.295 67.760 ;
        RECT 95.455 65.800 96.125 67.080 ;
        RECT 88.835 65.410 93.885 65.790 ;
        RECT 95.245 65.390 96.295 65.800 ;
        RECT 88.435 63.590 88.815 65.140 ;
        RECT 88.555 55.750 88.815 63.590 ;
        RECT 93.865 63.150 94.135 65.190 ;
        RECT 94.995 63.150 95.265 65.150 ;
        RECT 93.865 56.460 95.265 63.150 ;
        RECT 88.465 55.240 88.825 55.750 ;
        RECT 88.445 54.810 88.825 55.240 ;
        RECT 93.865 55.140 94.135 56.460 ;
        RECT 94.995 55.100 95.265 56.460 ;
        RECT 96.265 55.210 96.585 65.140 ;
        RECT 96.265 55.150 96.595 55.210 ;
        RECT 88.445 54.530 88.695 54.810 ;
        RECT 88.245 54.130 92.885 54.530 ;
        RECT 93.785 54.240 94.915 54.250 ;
        RECT 96.275 54.240 96.595 55.150 ;
        RECT 88.445 52.010 88.695 54.130 ;
        RECT 93.145 53.440 93.505 54.060 ;
        RECT 93.225 52.560 93.485 53.440 ;
        RECT 93.765 53.190 96.595 54.240 ;
        RECT 93.055 52.180 93.585 52.560 ;
        RECT 88.445 51.920 88.945 52.010 ;
        RECT 88.435 51.190 88.945 51.920 ;
        RECT 88.675 50.190 88.945 51.190 ;
        RECT 89.585 50.940 89.855 51.890 ;
        RECT 89.585 50.790 90.055 50.940 ;
        RECT 89.585 50.110 90.145 50.790 ;
        RECT 89.665 50.100 90.145 50.110 ;
        RECT 88.955 49.570 89.575 49.930 ;
        RECT 88.995 49.040 89.425 49.570 ;
        RECT 87.545 48.620 89.425 49.040 ;
        RECT 89.915 48.910 90.145 50.100 ;
        RECT 88.995 47.750 89.425 48.620 ;
        RECT 89.835 48.310 90.215 48.910 ;
        RECT 86.705 47.010 87.395 47.720 ;
        RECT 88.815 47.390 89.435 47.750 ;
        RECT 88.515 47.010 88.805 47.200 ;
        RECT 86.705 46.570 88.805 47.010 ;
        RECT 86.705 46.550 87.395 46.570 ;
        RECT 88.515 46.330 88.805 46.570 ;
        RECT 89.435 46.940 89.705 47.190 ;
        RECT 89.915 46.940 90.145 48.310 ;
        RECT 92.735 46.960 93.065 51.980 ;
        RECT 93.785 51.970 94.915 53.190 ;
        RECT 96.275 53.170 96.595 53.190 ;
        RECT 89.435 46.830 90.145 46.940 ;
        RECT 92.725 46.910 93.065 46.960 ;
        RECT 93.615 47.730 94.995 51.970 ;
        RECT 89.435 46.520 90.095 46.830 ;
        RECT 89.435 46.350 89.705 46.520 ;
        RECT 92.725 44.950 93.005 46.910 ;
        RECT 93.615 46.870 93.915 47.730 ;
        RECT 94.695 46.870 94.995 47.730 ;
        RECT 95.545 46.870 95.875 51.940 ;
        RECT 94.945 46.330 95.425 46.710 ;
        RECT 95.045 45.710 95.295 46.330 ;
        RECT 94.945 45.110 95.325 45.710 ;
        RECT 64.855 42.190 66.235 42.760 ;
        RECT 72.385 42.580 73.765 43.150 ;
        RECT 84.345 43.140 84.645 44.870 ;
        RECT 92.205 44.180 93.305 44.950 ;
        RECT 95.595 44.880 95.875 46.870 ;
        RECT 97.985 47.710 98.485 68.510 ;
        RECT 98.825 49.030 99.215 70.540 ;
        RECT 99.615 69.950 100.505 70.680 ;
        RECT 99.715 65.130 99.975 69.950 ;
        RECT 101.355 68.560 104.065 69.410 ;
        RECT 101.555 65.780 103.485 68.560 ;
        RECT 109.235 68.510 109.775 71.740 ;
        RECT 110.075 70.540 110.485 73.030 ;
        RECT 120.185 71.740 121.045 72.580 ;
        RECT 106.455 67.070 107.575 67.750 ;
        RECT 106.735 65.790 107.405 67.070 ;
        RECT 100.115 65.400 105.165 65.780 ;
        RECT 106.525 65.380 107.575 65.790 ;
        RECT 99.715 63.580 100.095 65.130 ;
        RECT 99.835 55.740 100.095 63.580 ;
        RECT 105.145 63.140 105.415 65.180 ;
        RECT 106.275 63.140 106.545 65.140 ;
        RECT 105.145 56.450 106.545 63.140 ;
        RECT 99.745 55.230 100.105 55.740 ;
        RECT 99.725 54.800 100.105 55.230 ;
        RECT 105.145 55.130 105.415 56.450 ;
        RECT 106.275 55.090 106.545 56.450 ;
        RECT 107.545 55.200 107.865 65.130 ;
        RECT 107.545 55.140 107.875 55.200 ;
        RECT 99.725 54.520 99.975 54.800 ;
        RECT 99.525 54.120 104.165 54.520 ;
        RECT 105.065 54.230 106.195 54.240 ;
        RECT 107.555 54.230 107.875 55.140 ;
        RECT 99.725 52.000 99.975 54.120 ;
        RECT 104.425 53.430 104.785 54.050 ;
        RECT 104.505 52.550 104.765 53.430 ;
        RECT 105.045 53.180 107.875 54.230 ;
        RECT 104.335 52.170 104.865 52.550 ;
        RECT 99.725 51.910 100.225 52.000 ;
        RECT 99.715 51.180 100.225 51.910 ;
        RECT 99.955 50.180 100.225 51.180 ;
        RECT 100.865 50.930 101.135 51.880 ;
        RECT 100.865 50.780 101.335 50.930 ;
        RECT 100.865 50.100 101.425 50.780 ;
        RECT 100.945 50.090 101.425 50.100 ;
        RECT 100.235 49.560 100.855 49.920 ;
        RECT 100.275 49.030 100.705 49.560 ;
        RECT 98.825 48.610 100.705 49.030 ;
        RECT 101.195 48.900 101.425 50.090 ;
        RECT 100.275 47.740 100.705 48.610 ;
        RECT 101.115 48.300 101.495 48.900 ;
        RECT 97.985 47.000 98.675 47.710 ;
        RECT 100.095 47.380 100.715 47.740 ;
        RECT 99.795 47.000 100.085 47.190 ;
        RECT 97.985 46.560 100.085 47.000 ;
        RECT 97.985 46.540 98.675 46.560 ;
        RECT 99.795 46.320 100.085 46.560 ;
        RECT 100.715 46.930 100.985 47.180 ;
        RECT 101.195 46.930 101.425 48.300 ;
        RECT 104.015 46.950 104.345 51.970 ;
        RECT 105.065 51.960 106.195 53.180 ;
        RECT 107.555 53.160 107.875 53.180 ;
        RECT 100.715 46.820 101.425 46.930 ;
        RECT 104.005 46.900 104.345 46.950 ;
        RECT 104.895 47.720 106.275 51.960 ;
        RECT 100.715 46.510 101.375 46.820 ;
        RECT 100.715 46.340 100.985 46.510 ;
        RECT 104.005 44.940 104.285 46.900 ;
        RECT 104.895 46.860 105.195 47.720 ;
        RECT 105.975 46.860 106.275 47.720 ;
        RECT 106.825 46.860 107.155 51.930 ;
        RECT 106.225 46.320 106.705 46.700 ;
        RECT 106.325 45.700 106.575 46.320 ;
        RECT 106.225 45.100 106.605 45.700 ;
        RECT 95.595 43.150 95.895 44.880 ;
        RECT 103.485 44.170 104.585 44.940 ;
        RECT 106.875 44.870 107.155 46.860 ;
        RECT 109.255 47.710 109.755 68.510 ;
        RECT 110.095 49.030 110.485 70.540 ;
        RECT 110.885 69.950 111.775 70.680 ;
        RECT 110.985 65.130 111.245 69.950 ;
        RECT 112.625 68.560 115.335 69.410 ;
        RECT 112.825 65.780 114.755 68.560 ;
        RECT 120.485 68.510 121.025 71.740 ;
        RECT 121.325 70.540 121.735 73.110 ;
        RECT 132.925 70.810 133.225 70.900 ;
        RECT 117.725 67.070 118.845 67.750 ;
        RECT 118.005 65.790 118.675 67.070 ;
        RECT 111.385 65.400 116.435 65.780 ;
        RECT 117.795 65.380 118.845 65.790 ;
        RECT 110.985 63.580 111.365 65.130 ;
        RECT 111.105 55.740 111.365 63.580 ;
        RECT 116.415 63.140 116.685 65.180 ;
        RECT 117.545 63.140 117.815 65.140 ;
        RECT 116.415 56.450 117.815 63.140 ;
        RECT 111.015 55.230 111.375 55.740 ;
        RECT 110.995 54.800 111.375 55.230 ;
        RECT 116.415 55.130 116.685 56.450 ;
        RECT 117.545 55.090 117.815 56.450 ;
        RECT 118.815 55.200 119.135 65.130 ;
        RECT 118.815 55.140 119.145 55.200 ;
        RECT 110.995 54.520 111.245 54.800 ;
        RECT 110.795 54.120 115.435 54.520 ;
        RECT 116.335 54.230 117.465 54.240 ;
        RECT 118.825 54.230 119.145 55.140 ;
        RECT 110.995 52.000 111.245 54.120 ;
        RECT 115.695 53.430 116.055 54.050 ;
        RECT 115.775 52.550 116.035 53.430 ;
        RECT 116.315 53.180 119.145 54.230 ;
        RECT 115.605 52.170 116.135 52.550 ;
        RECT 110.995 51.910 111.495 52.000 ;
        RECT 110.985 51.180 111.495 51.910 ;
        RECT 111.225 50.180 111.495 51.180 ;
        RECT 112.135 50.930 112.405 51.880 ;
        RECT 112.135 50.780 112.605 50.930 ;
        RECT 112.135 50.100 112.695 50.780 ;
        RECT 112.215 50.090 112.695 50.100 ;
        RECT 111.505 49.560 112.125 49.920 ;
        RECT 111.545 49.030 111.975 49.560 ;
        RECT 110.095 48.610 111.975 49.030 ;
        RECT 112.465 48.900 112.695 50.090 ;
        RECT 111.545 47.740 111.975 48.610 ;
        RECT 112.385 48.300 112.765 48.900 ;
        RECT 109.255 47.000 109.945 47.710 ;
        RECT 111.365 47.380 111.985 47.740 ;
        RECT 111.065 47.000 111.355 47.190 ;
        RECT 109.255 46.560 111.355 47.000 ;
        RECT 109.255 46.540 109.945 46.560 ;
        RECT 111.065 46.320 111.355 46.560 ;
        RECT 111.985 46.930 112.255 47.180 ;
        RECT 112.465 46.930 112.695 48.300 ;
        RECT 115.285 46.950 115.615 51.970 ;
        RECT 116.335 51.960 117.465 53.180 ;
        RECT 118.825 53.160 119.145 53.180 ;
        RECT 111.985 46.820 112.695 46.930 ;
        RECT 115.275 46.900 115.615 46.950 ;
        RECT 116.165 47.720 117.545 51.960 ;
        RECT 111.985 46.510 112.645 46.820 ;
        RECT 111.985 46.340 112.255 46.510 ;
        RECT 115.275 44.940 115.555 46.900 ;
        RECT 116.165 46.860 116.465 47.720 ;
        RECT 117.245 46.860 117.545 47.720 ;
        RECT 118.095 46.860 118.425 51.930 ;
        RECT 117.495 46.320 117.975 46.700 ;
        RECT 117.595 45.700 117.845 46.320 ;
        RECT 117.495 45.100 117.875 45.700 ;
        RECT 20.795 39.650 21.175 40.250 ;
        RECT 20.825 39.030 21.075 39.650 ;
        RECT 20.695 38.650 21.175 39.030 ;
        RECT 20.245 33.420 20.575 38.490 ;
        RECT 21.125 37.630 21.425 38.490 ;
        RECT 22.205 37.630 22.505 38.490 ;
        RECT 23.115 38.450 23.395 40.410 ;
        RECT 26.415 38.840 26.685 39.010 ;
        RECT 26.025 38.530 26.685 38.840 ;
        RECT 21.125 33.390 22.505 37.630 ;
        RECT 23.055 38.400 23.395 38.450 ;
        RECT 25.975 38.420 26.685 38.530 ;
        RECT 19.525 32.170 19.845 32.190 ;
        RECT 21.205 32.170 22.335 33.390 ;
        RECT 23.055 33.380 23.385 38.400 ;
        RECT 25.975 37.050 26.205 38.420 ;
        RECT 26.415 38.170 26.685 38.420 ;
        RECT 27.315 38.790 27.605 39.030 ;
        RECT 28.725 38.790 29.415 38.810 ;
        RECT 27.315 38.350 29.415 38.790 ;
        RECT 27.315 38.160 27.605 38.350 ;
        RECT 26.685 37.610 27.305 37.970 ;
        RECT 28.725 37.640 29.415 38.350 ;
        RECT 25.905 36.450 26.285 37.050 ;
        RECT 26.695 36.740 27.125 37.610 ;
        RECT 25.975 35.260 26.205 36.450 ;
        RECT 26.695 36.320 28.575 36.740 ;
        RECT 26.695 35.790 27.125 36.320 ;
        RECT 26.545 35.430 27.165 35.790 ;
        RECT 25.975 35.250 26.455 35.260 ;
        RECT 25.975 34.570 26.535 35.250 ;
        RECT 26.065 34.420 26.535 34.570 ;
        RECT 26.265 33.470 26.535 34.420 ;
        RECT 27.175 34.170 27.445 35.170 ;
        RECT 27.175 33.440 27.685 34.170 ;
        RECT 27.175 33.350 27.675 33.440 ;
        RECT 22.535 32.800 23.065 33.180 ;
        RECT 19.525 31.120 22.355 32.170 ;
        RECT 22.635 31.920 22.895 32.800 ;
        RECT 22.615 31.300 22.975 31.920 ;
        RECT 27.425 31.230 27.675 33.350 ;
        RECT 19.525 30.210 19.845 31.120 ;
        RECT 21.205 31.110 22.335 31.120 ;
        RECT 23.235 30.830 27.875 31.230 ;
        RECT 27.425 30.550 27.675 30.830 ;
        RECT 19.525 30.150 19.855 30.210 ;
        RECT 19.535 20.220 19.855 30.150 ;
        RECT 20.855 28.900 21.125 30.260 ;
        RECT 21.985 28.900 22.255 30.220 ;
        RECT 27.295 30.120 27.675 30.550 ;
        RECT 27.295 29.610 27.655 30.120 ;
        RECT 20.855 22.210 22.255 28.900 ;
        RECT 20.855 20.210 21.125 22.210 ;
        RECT 21.985 20.170 22.255 22.210 ;
        RECT 27.305 21.770 27.565 29.610 ;
        RECT 27.305 20.220 27.685 21.770 ;
        RECT 19.825 19.560 20.875 19.970 ;
        RECT 22.235 19.570 27.285 19.950 ;
        RECT 19.995 18.280 20.665 19.560 ;
        RECT 19.825 17.600 20.945 18.280 ;
        RECT 23.915 16.790 25.845 19.570 ;
        RECT 23.335 15.940 26.045 16.790 ;
        RECT 27.425 15.400 27.685 20.220 ;
        RECT 26.895 14.670 27.785 15.400 ;
        RECT 28.185 14.810 28.575 36.320 ;
        RECT 28.915 16.840 29.415 37.640 ;
        RECT 31.525 38.490 31.805 40.480 ;
        RECT 34.095 40.410 35.195 41.180 ;
        RECT 42.795 40.460 43.095 42.190 ;
        RECT 32.075 39.650 32.455 40.250 ;
        RECT 32.105 39.030 32.355 39.650 ;
        RECT 31.975 38.650 32.455 39.030 ;
        RECT 31.525 33.420 31.855 38.490 ;
        RECT 32.405 37.630 32.705 38.490 ;
        RECT 33.485 37.630 33.785 38.490 ;
        RECT 34.395 38.450 34.675 40.410 ;
        RECT 37.695 38.840 37.965 39.010 ;
        RECT 37.305 38.530 37.965 38.840 ;
        RECT 32.405 33.390 33.785 37.630 ;
        RECT 34.335 38.400 34.675 38.450 ;
        RECT 37.255 38.420 37.965 38.530 ;
        RECT 30.805 32.170 31.125 32.190 ;
        RECT 32.485 32.170 33.615 33.390 ;
        RECT 34.335 33.380 34.665 38.400 ;
        RECT 37.255 37.050 37.485 38.420 ;
        RECT 37.695 38.170 37.965 38.420 ;
        RECT 38.595 38.790 38.885 39.030 ;
        RECT 40.005 38.790 40.695 38.810 ;
        RECT 38.595 38.350 40.695 38.790 ;
        RECT 38.595 38.160 38.885 38.350 ;
        RECT 37.965 37.610 38.585 37.970 ;
        RECT 40.005 37.640 40.695 38.350 ;
        RECT 37.185 36.450 37.565 37.050 ;
        RECT 37.975 36.740 38.405 37.610 ;
        RECT 37.255 35.260 37.485 36.450 ;
        RECT 37.975 36.320 39.855 36.740 ;
        RECT 37.975 35.790 38.405 36.320 ;
        RECT 37.825 35.430 38.445 35.790 ;
        RECT 37.255 35.250 37.735 35.260 ;
        RECT 37.255 34.570 37.815 35.250 ;
        RECT 37.345 34.420 37.815 34.570 ;
        RECT 37.545 33.470 37.815 34.420 ;
        RECT 38.455 34.170 38.725 35.170 ;
        RECT 38.455 33.440 38.965 34.170 ;
        RECT 38.455 33.350 38.955 33.440 ;
        RECT 33.815 32.800 34.345 33.180 ;
        RECT 30.805 31.120 33.635 32.170 ;
        RECT 33.915 31.920 34.175 32.800 ;
        RECT 33.895 31.300 34.255 31.920 ;
        RECT 38.705 31.230 38.955 33.350 ;
        RECT 30.805 30.210 31.125 31.120 ;
        RECT 32.485 31.110 33.615 31.120 ;
        RECT 34.515 30.830 39.155 31.230 ;
        RECT 38.705 30.550 38.955 30.830 ;
        RECT 30.805 30.150 31.135 30.210 ;
        RECT 30.815 20.220 31.135 30.150 ;
        RECT 32.135 28.900 32.405 30.260 ;
        RECT 33.265 28.900 33.535 30.220 ;
        RECT 38.575 30.120 38.955 30.550 ;
        RECT 38.575 29.610 38.935 30.120 ;
        RECT 32.135 22.210 33.535 28.900 ;
        RECT 32.135 20.210 32.405 22.210 ;
        RECT 33.265 20.170 33.535 22.210 ;
        RECT 38.585 21.770 38.845 29.610 ;
        RECT 38.585 20.220 38.965 21.770 ;
        RECT 31.105 19.560 32.155 19.970 ;
        RECT 33.515 19.570 38.565 19.950 ;
        RECT 31.275 18.280 31.945 19.560 ;
        RECT 31.105 17.600 32.225 18.280 ;
        RECT 28.185 12.290 28.595 14.810 ;
        RECT 28.895 13.610 29.435 16.840 ;
        RECT 35.195 16.790 37.125 19.570 ;
        RECT 34.615 15.940 37.325 16.790 ;
        RECT 38.705 15.400 38.965 20.220 ;
        RECT 38.175 14.670 39.065 15.400 ;
        RECT 39.465 14.810 39.855 36.320 ;
        RECT 40.195 16.840 40.695 37.640 ;
        RECT 42.815 38.470 43.095 40.460 ;
        RECT 45.385 40.390 46.485 41.160 ;
        RECT 54.015 40.460 54.315 42.190 ;
        RECT 43.365 39.630 43.745 40.230 ;
        RECT 43.395 39.010 43.645 39.630 ;
        RECT 43.265 38.630 43.745 39.010 ;
        RECT 42.815 33.400 43.145 38.470 ;
        RECT 43.695 37.610 43.995 38.470 ;
        RECT 44.775 37.610 45.075 38.470 ;
        RECT 45.685 38.430 45.965 40.390 ;
        RECT 48.985 38.820 49.255 38.990 ;
        RECT 48.595 38.510 49.255 38.820 ;
        RECT 43.695 33.370 45.075 37.610 ;
        RECT 45.625 38.380 45.965 38.430 ;
        RECT 48.545 38.400 49.255 38.510 ;
        RECT 42.095 32.150 42.415 32.170 ;
        RECT 43.775 32.150 44.905 33.370 ;
        RECT 45.625 33.360 45.955 38.380 ;
        RECT 48.545 37.030 48.775 38.400 ;
        RECT 48.985 38.150 49.255 38.400 ;
        RECT 49.885 38.770 50.175 39.010 ;
        RECT 51.295 38.770 51.985 38.790 ;
        RECT 49.885 38.330 51.985 38.770 ;
        RECT 49.885 38.140 50.175 38.330 ;
        RECT 49.255 37.590 49.875 37.950 ;
        RECT 51.295 37.620 51.985 38.330 ;
        RECT 48.475 36.430 48.855 37.030 ;
        RECT 49.265 36.720 49.695 37.590 ;
        RECT 48.545 35.240 48.775 36.430 ;
        RECT 49.265 36.300 51.145 36.720 ;
        RECT 49.265 35.770 49.695 36.300 ;
        RECT 49.115 35.410 49.735 35.770 ;
        RECT 48.545 35.230 49.025 35.240 ;
        RECT 48.545 34.550 49.105 35.230 ;
        RECT 48.635 34.400 49.105 34.550 ;
        RECT 48.835 33.450 49.105 34.400 ;
        RECT 49.745 34.150 50.015 35.150 ;
        RECT 49.745 33.420 50.255 34.150 ;
        RECT 49.745 33.330 50.245 33.420 ;
        RECT 45.105 32.780 45.635 33.160 ;
        RECT 42.095 31.100 44.925 32.150 ;
        RECT 45.205 31.900 45.465 32.780 ;
        RECT 45.185 31.280 45.545 31.900 ;
        RECT 49.995 31.210 50.245 33.330 ;
        RECT 42.095 30.190 42.415 31.100 ;
        RECT 43.775 31.090 44.905 31.100 ;
        RECT 45.805 30.810 50.445 31.210 ;
        RECT 49.995 30.530 50.245 30.810 ;
        RECT 42.095 30.130 42.425 30.190 ;
        RECT 42.105 20.200 42.425 30.130 ;
        RECT 43.425 28.880 43.695 30.240 ;
        RECT 44.555 28.880 44.825 30.200 ;
        RECT 49.865 30.100 50.245 30.530 ;
        RECT 49.865 29.590 50.225 30.100 ;
        RECT 43.425 22.190 44.825 28.880 ;
        RECT 43.425 20.190 43.695 22.190 ;
        RECT 44.555 20.150 44.825 22.190 ;
        RECT 49.875 21.750 50.135 29.590 ;
        RECT 49.875 20.200 50.255 21.750 ;
        RECT 42.395 19.540 43.445 19.950 ;
        RECT 44.805 19.550 49.855 19.930 ;
        RECT 42.565 18.260 43.235 19.540 ;
        RECT 42.395 17.580 43.515 18.260 ;
        RECT 28.875 12.770 29.735 13.610 ;
        RECT 28.185 11.950 30.415 12.290 ;
        RECT 39.465 11.990 39.875 14.810 ;
        RECT 40.175 13.610 40.715 16.840 ;
        RECT 46.485 16.770 48.415 19.550 ;
        RECT 45.905 15.920 48.615 16.770 ;
        RECT 49.995 15.380 50.255 20.200 ;
        RECT 49.465 14.650 50.355 15.380 ;
        RECT 50.755 14.790 51.145 36.300 ;
        RECT 51.485 16.820 51.985 37.620 ;
        RECT 54.035 38.470 54.315 40.460 ;
        RECT 56.605 40.390 57.705 41.160 ;
        RECT 65.215 40.460 65.515 42.190 ;
        RECT 76.145 42.180 77.525 42.750 ;
        RECT 83.625 42.570 85.005 43.140 ;
        RECT 87.385 42.200 88.765 42.770 ;
        RECT 94.875 42.580 96.255 43.150 ;
        RECT 106.875 43.140 107.175 44.870 ;
        RECT 114.755 44.170 115.855 44.940 ;
        RECT 118.145 44.870 118.425 46.860 ;
        RECT 120.505 47.710 121.005 68.510 ;
        RECT 121.345 49.030 121.735 70.540 ;
        RECT 122.135 69.950 123.025 70.680 ;
        RECT 132.615 70.040 134.265 70.810 ;
        RECT 122.235 65.130 122.495 69.950 ;
        RECT 123.875 68.560 126.585 69.410 ;
        RECT 124.075 65.780 126.005 68.560 ;
        RECT 128.975 67.070 130.095 67.750 ;
        RECT 129.255 65.790 129.925 67.070 ;
        RECT 122.635 65.400 127.685 65.780 ;
        RECT 129.045 65.380 130.095 65.790 ;
        RECT 132.925 65.180 133.225 70.040 ;
        RECT 137.675 68.690 139.075 69.460 ;
        RECT 138.385 65.740 138.645 68.690 ;
        RECT 149.410 68.420 150.690 69.620 ;
        RECT 149.480 65.810 150.640 68.420 ;
        RECT 133.365 65.380 138.645 65.740 ;
        RECT 122.235 63.580 122.615 65.130 ;
        RECT 122.355 55.740 122.615 63.580 ;
        RECT 127.665 63.140 127.935 65.180 ;
        RECT 128.795 63.140 129.065 65.140 ;
        RECT 127.665 56.450 129.065 63.140 ;
        RECT 122.265 55.230 122.625 55.740 ;
        RECT 122.245 54.800 122.625 55.230 ;
        RECT 127.665 55.130 127.935 56.450 ;
        RECT 128.795 55.090 129.065 56.450 ;
        RECT 130.065 55.200 130.385 65.130 ;
        RECT 132.925 61.010 133.355 65.180 ;
        RECT 138.385 65.150 138.645 65.380 ;
        RECT 138.385 64.770 138.675 65.150 ;
        RECT 130.065 55.140 130.395 55.200 ;
        RECT 133.055 55.190 133.355 61.010 ;
        RECT 122.245 54.520 122.495 54.800 ;
        RECT 122.045 54.120 126.685 54.520 ;
        RECT 127.585 54.230 128.715 54.240 ;
        RECT 130.075 54.230 130.395 55.140 ;
        RECT 138.395 55.080 138.675 64.770 ;
        RECT 149.390 64.610 150.670 65.810 ;
        RECT 122.245 52.000 122.495 54.120 ;
        RECT 126.945 53.430 127.305 54.050 ;
        RECT 127.025 52.550 127.285 53.430 ;
        RECT 127.565 53.180 130.395 54.230 ;
        RECT 126.855 52.170 127.385 52.550 ;
        RECT 122.245 51.910 122.745 52.000 ;
        RECT 122.235 51.180 122.745 51.910 ;
        RECT 122.475 50.180 122.745 51.180 ;
        RECT 123.385 50.930 123.655 51.880 ;
        RECT 123.385 50.780 123.855 50.930 ;
        RECT 123.385 50.100 123.945 50.780 ;
        RECT 123.465 50.090 123.945 50.100 ;
        RECT 122.755 49.560 123.375 49.920 ;
        RECT 122.795 49.030 123.225 49.560 ;
        RECT 121.345 48.610 123.225 49.030 ;
        RECT 123.715 48.900 123.945 50.090 ;
        RECT 122.795 47.740 123.225 48.610 ;
        RECT 123.635 48.300 124.015 48.900 ;
        RECT 120.505 47.000 121.195 47.710 ;
        RECT 122.615 47.380 123.235 47.740 ;
        RECT 122.315 47.000 122.605 47.190 ;
        RECT 120.505 46.560 122.605 47.000 ;
        RECT 120.505 46.540 121.195 46.560 ;
        RECT 122.315 46.320 122.605 46.560 ;
        RECT 123.235 46.930 123.505 47.180 ;
        RECT 123.715 46.930 123.945 48.300 ;
        RECT 126.535 46.950 126.865 51.970 ;
        RECT 127.585 51.960 128.715 53.180 ;
        RECT 130.075 53.160 130.395 53.180 ;
        RECT 123.235 46.820 123.945 46.930 ;
        RECT 126.525 46.900 126.865 46.950 ;
        RECT 127.415 47.720 128.795 51.960 ;
        RECT 123.235 46.510 123.895 46.820 ;
        RECT 123.235 46.340 123.505 46.510 ;
        RECT 126.525 44.940 126.805 46.900 ;
        RECT 127.415 46.860 127.715 47.720 ;
        RECT 128.495 46.860 128.795 47.720 ;
        RECT 129.345 46.860 129.675 51.930 ;
        RECT 128.745 46.320 129.225 46.700 ;
        RECT 128.845 45.700 129.095 46.320 ;
        RECT 128.745 45.100 129.125 45.700 ;
        RECT 118.145 43.140 118.445 44.870 ;
        RECT 126.005 44.170 127.105 44.940 ;
        RECT 129.395 44.870 129.675 46.860 ;
        RECT 129.395 43.140 129.695 44.870 ;
        RECT 98.595 42.220 99.975 42.790 ;
        RECT 106.155 42.570 107.535 43.140 ;
        RECT 109.795 42.260 111.175 42.830 ;
        RECT 117.425 42.570 118.805 43.140 ;
        RECT 121.005 42.280 122.385 42.850 ;
        RECT 128.675 42.570 130.055 43.140 ;
        RECT 54.585 39.630 54.965 40.230 ;
        RECT 54.615 39.010 54.865 39.630 ;
        RECT 54.485 38.630 54.965 39.010 ;
        RECT 54.035 33.400 54.365 38.470 ;
        RECT 54.915 37.610 55.215 38.470 ;
        RECT 55.995 37.610 56.295 38.470 ;
        RECT 56.905 38.430 57.185 40.390 ;
        RECT 60.205 38.820 60.475 38.990 ;
        RECT 59.815 38.510 60.475 38.820 ;
        RECT 54.915 33.370 56.295 37.610 ;
        RECT 56.845 38.380 57.185 38.430 ;
        RECT 59.765 38.400 60.475 38.510 ;
        RECT 53.315 32.150 53.635 32.170 ;
        RECT 54.995 32.150 56.125 33.370 ;
        RECT 56.845 33.360 57.175 38.380 ;
        RECT 59.765 37.030 59.995 38.400 ;
        RECT 60.205 38.150 60.475 38.400 ;
        RECT 61.105 38.770 61.395 39.010 ;
        RECT 62.515 38.770 63.205 38.790 ;
        RECT 61.105 38.330 63.205 38.770 ;
        RECT 61.105 38.140 61.395 38.330 ;
        RECT 60.475 37.590 61.095 37.950 ;
        RECT 62.515 37.620 63.205 38.330 ;
        RECT 59.695 36.430 60.075 37.030 ;
        RECT 60.485 36.720 60.915 37.590 ;
        RECT 59.765 35.240 59.995 36.430 ;
        RECT 60.485 36.300 62.365 36.720 ;
        RECT 60.485 35.770 60.915 36.300 ;
        RECT 60.335 35.410 60.955 35.770 ;
        RECT 59.765 35.230 60.245 35.240 ;
        RECT 59.765 34.550 60.325 35.230 ;
        RECT 59.855 34.400 60.325 34.550 ;
        RECT 60.055 33.450 60.325 34.400 ;
        RECT 60.965 34.150 61.235 35.150 ;
        RECT 60.965 33.420 61.475 34.150 ;
        RECT 60.965 33.330 61.465 33.420 ;
        RECT 56.325 32.780 56.855 33.160 ;
        RECT 53.315 31.100 56.145 32.150 ;
        RECT 56.425 31.900 56.685 32.780 ;
        RECT 56.405 31.280 56.765 31.900 ;
        RECT 61.215 31.210 61.465 33.330 ;
        RECT 53.315 30.190 53.635 31.100 ;
        RECT 54.995 31.090 56.125 31.100 ;
        RECT 57.025 30.810 61.665 31.210 ;
        RECT 61.215 30.530 61.465 30.810 ;
        RECT 53.315 30.130 53.645 30.190 ;
        RECT 53.325 20.200 53.645 30.130 ;
        RECT 54.645 28.880 54.915 30.240 ;
        RECT 55.775 28.880 56.045 30.200 ;
        RECT 61.085 30.100 61.465 30.530 ;
        RECT 61.085 29.590 61.445 30.100 ;
        RECT 54.645 22.190 56.045 28.880 ;
        RECT 54.645 20.190 54.915 22.190 ;
        RECT 55.775 20.150 56.045 22.190 ;
        RECT 61.095 21.750 61.355 29.590 ;
        RECT 61.095 20.200 61.475 21.750 ;
        RECT 53.615 19.540 54.665 19.950 ;
        RECT 56.025 19.550 61.075 19.930 ;
        RECT 53.785 18.260 54.455 19.540 ;
        RECT 53.615 17.580 54.735 18.260 ;
        RECT 40.155 12.770 41.015 13.610 ;
        RECT 50.755 12.170 51.165 14.790 ;
        RECT 51.465 13.590 52.005 16.820 ;
        RECT 57.705 16.770 59.635 19.550 ;
        RECT 57.125 15.920 59.835 16.770 ;
        RECT 61.215 15.380 61.475 20.200 ;
        RECT 60.685 14.650 61.575 15.380 ;
        RECT 61.975 14.790 62.365 36.300 ;
        RECT 62.705 16.820 63.205 37.620 ;
        RECT 65.235 38.470 65.515 40.460 ;
        RECT 67.805 40.390 68.905 41.160 ;
        RECT 76.505 40.450 76.805 42.180 ;
        RECT 65.785 39.630 66.165 40.230 ;
        RECT 65.815 39.010 66.065 39.630 ;
        RECT 65.685 38.630 66.165 39.010 ;
        RECT 65.235 33.400 65.565 38.470 ;
        RECT 66.115 37.610 66.415 38.470 ;
        RECT 67.195 37.610 67.495 38.470 ;
        RECT 68.105 38.430 68.385 40.390 ;
        RECT 71.405 38.820 71.675 38.990 ;
        RECT 71.015 38.510 71.675 38.820 ;
        RECT 66.115 33.370 67.495 37.610 ;
        RECT 68.045 38.380 68.385 38.430 ;
        RECT 70.965 38.400 71.675 38.510 ;
        RECT 64.515 32.150 64.835 32.170 ;
        RECT 66.195 32.150 67.325 33.370 ;
        RECT 68.045 33.360 68.375 38.380 ;
        RECT 70.965 37.030 71.195 38.400 ;
        RECT 71.405 38.150 71.675 38.400 ;
        RECT 72.305 38.770 72.595 39.010 ;
        RECT 73.715 38.770 74.405 38.790 ;
        RECT 72.305 38.330 74.405 38.770 ;
        RECT 72.305 38.140 72.595 38.330 ;
        RECT 71.675 37.590 72.295 37.950 ;
        RECT 73.715 37.620 74.405 38.330 ;
        RECT 70.895 36.430 71.275 37.030 ;
        RECT 71.685 36.720 72.115 37.590 ;
        RECT 70.965 35.240 71.195 36.430 ;
        RECT 71.685 36.300 73.565 36.720 ;
        RECT 71.685 35.770 72.115 36.300 ;
        RECT 71.535 35.410 72.155 35.770 ;
        RECT 70.965 35.230 71.445 35.240 ;
        RECT 70.965 34.550 71.525 35.230 ;
        RECT 71.055 34.400 71.525 34.550 ;
        RECT 71.255 33.450 71.525 34.400 ;
        RECT 72.165 34.150 72.435 35.150 ;
        RECT 72.165 33.420 72.675 34.150 ;
        RECT 72.165 33.330 72.665 33.420 ;
        RECT 67.525 32.780 68.055 33.160 ;
        RECT 64.515 31.100 67.345 32.150 ;
        RECT 67.625 31.900 67.885 32.780 ;
        RECT 67.605 31.280 67.965 31.900 ;
        RECT 72.415 31.210 72.665 33.330 ;
        RECT 64.515 30.190 64.835 31.100 ;
        RECT 66.195 31.090 67.325 31.100 ;
        RECT 68.225 30.810 72.865 31.210 ;
        RECT 72.415 30.530 72.665 30.810 ;
        RECT 64.515 30.130 64.845 30.190 ;
        RECT 64.525 20.200 64.845 30.130 ;
        RECT 65.845 28.880 66.115 30.240 ;
        RECT 66.975 28.880 67.245 30.200 ;
        RECT 72.285 30.100 72.665 30.530 ;
        RECT 72.285 29.590 72.645 30.100 ;
        RECT 65.845 22.190 67.245 28.880 ;
        RECT 65.845 20.190 66.115 22.190 ;
        RECT 66.975 20.150 67.245 22.190 ;
        RECT 72.295 21.750 72.555 29.590 ;
        RECT 72.295 20.200 72.675 21.750 ;
        RECT 64.815 19.540 65.865 19.950 ;
        RECT 67.225 19.550 72.275 19.930 ;
        RECT 64.985 18.260 65.655 19.540 ;
        RECT 64.815 17.580 65.935 18.260 ;
        RECT 51.445 12.750 52.305 13.590 ;
        RECT 27.865 11.130 30.415 11.950 ;
        RECT 28.395 11.090 30.415 11.130 ;
        RECT 39.115 10.980 41.565 11.990 ;
        RECT 50.335 10.970 52.355 12.170 ;
        RECT 61.975 12.160 62.385 14.790 ;
        RECT 62.685 13.590 63.225 16.820 ;
        RECT 68.905 16.770 70.835 19.550 ;
        RECT 68.325 15.920 71.035 16.770 ;
        RECT 72.415 15.380 72.675 20.200 ;
        RECT 71.885 14.650 72.775 15.380 ;
        RECT 73.175 14.790 73.565 36.300 ;
        RECT 73.905 16.820 74.405 37.620 ;
        RECT 76.525 38.460 76.805 40.450 ;
        RECT 79.095 40.380 80.195 41.150 ;
        RECT 87.745 40.470 88.045 42.200 ;
        RECT 77.075 39.620 77.455 40.220 ;
        RECT 77.105 39.000 77.355 39.620 ;
        RECT 76.975 38.620 77.455 39.000 ;
        RECT 76.525 33.390 76.855 38.460 ;
        RECT 77.405 37.600 77.705 38.460 ;
        RECT 78.485 37.600 78.785 38.460 ;
        RECT 79.395 38.420 79.675 40.380 ;
        RECT 82.695 38.810 82.965 38.980 ;
        RECT 82.305 38.500 82.965 38.810 ;
        RECT 77.405 33.360 78.785 37.600 ;
        RECT 79.335 38.370 79.675 38.420 ;
        RECT 82.255 38.390 82.965 38.500 ;
        RECT 75.805 32.140 76.125 32.160 ;
        RECT 77.485 32.140 78.615 33.360 ;
        RECT 79.335 33.350 79.665 38.370 ;
        RECT 82.255 37.020 82.485 38.390 ;
        RECT 82.695 38.140 82.965 38.390 ;
        RECT 83.595 38.760 83.885 39.000 ;
        RECT 85.005 38.760 85.695 38.780 ;
        RECT 83.595 38.320 85.695 38.760 ;
        RECT 83.595 38.130 83.885 38.320 ;
        RECT 82.965 37.580 83.585 37.940 ;
        RECT 85.005 37.610 85.695 38.320 ;
        RECT 82.185 36.420 82.565 37.020 ;
        RECT 82.975 36.710 83.405 37.580 ;
        RECT 82.255 35.230 82.485 36.420 ;
        RECT 82.975 36.290 84.855 36.710 ;
        RECT 82.975 35.760 83.405 36.290 ;
        RECT 82.825 35.400 83.445 35.760 ;
        RECT 82.255 35.220 82.735 35.230 ;
        RECT 82.255 34.540 82.815 35.220 ;
        RECT 82.345 34.390 82.815 34.540 ;
        RECT 82.545 33.440 82.815 34.390 ;
        RECT 83.455 34.140 83.725 35.140 ;
        RECT 83.455 33.410 83.965 34.140 ;
        RECT 83.455 33.320 83.955 33.410 ;
        RECT 78.815 32.770 79.345 33.150 ;
        RECT 75.805 31.090 78.635 32.140 ;
        RECT 78.915 31.890 79.175 32.770 ;
        RECT 78.895 31.270 79.255 31.890 ;
        RECT 83.705 31.200 83.955 33.320 ;
        RECT 75.805 30.180 76.125 31.090 ;
        RECT 77.485 31.080 78.615 31.090 ;
        RECT 79.515 30.800 84.155 31.200 ;
        RECT 83.705 30.520 83.955 30.800 ;
        RECT 75.805 30.120 76.135 30.180 ;
        RECT 75.815 20.190 76.135 30.120 ;
        RECT 77.135 28.870 77.405 30.230 ;
        RECT 78.265 28.870 78.535 30.190 ;
        RECT 83.575 30.090 83.955 30.520 ;
        RECT 83.575 29.580 83.935 30.090 ;
        RECT 77.135 22.180 78.535 28.870 ;
        RECT 77.135 20.180 77.405 22.180 ;
        RECT 78.265 20.140 78.535 22.180 ;
        RECT 83.585 21.740 83.845 29.580 ;
        RECT 83.585 20.190 83.965 21.740 ;
        RECT 76.105 19.530 77.155 19.940 ;
        RECT 78.515 19.540 83.565 19.920 ;
        RECT 76.275 18.250 76.945 19.530 ;
        RECT 76.105 17.570 77.225 18.250 ;
        RECT 62.665 12.750 63.525 13.590 ;
        RECT 73.175 12.190 73.585 14.790 ;
        RECT 73.885 13.590 74.425 16.820 ;
        RECT 80.195 16.760 82.125 19.540 ;
        RECT 79.615 15.910 82.325 16.760 ;
        RECT 83.705 15.370 83.965 20.190 ;
        RECT 83.175 14.640 84.065 15.370 ;
        RECT 84.465 14.780 84.855 36.290 ;
        RECT 85.195 16.810 85.695 37.610 ;
        RECT 87.765 38.480 88.045 40.470 ;
        RECT 90.335 40.400 91.435 41.170 ;
        RECT 98.955 40.490 99.255 42.220 ;
        RECT 88.315 39.640 88.695 40.240 ;
        RECT 88.345 39.020 88.595 39.640 ;
        RECT 88.215 38.640 88.695 39.020 ;
        RECT 87.765 33.410 88.095 38.480 ;
        RECT 88.645 37.620 88.945 38.480 ;
        RECT 89.725 37.620 90.025 38.480 ;
        RECT 90.635 38.440 90.915 40.400 ;
        RECT 93.935 38.830 94.205 39.000 ;
        RECT 93.545 38.520 94.205 38.830 ;
        RECT 88.645 33.380 90.025 37.620 ;
        RECT 90.575 38.390 90.915 38.440 ;
        RECT 93.495 38.410 94.205 38.520 ;
        RECT 87.045 32.160 87.365 32.180 ;
        RECT 88.725 32.160 89.855 33.380 ;
        RECT 90.575 33.370 90.905 38.390 ;
        RECT 93.495 37.040 93.725 38.410 ;
        RECT 93.935 38.160 94.205 38.410 ;
        RECT 94.835 38.780 95.125 39.020 ;
        RECT 96.245 38.780 96.935 38.800 ;
        RECT 94.835 38.340 96.935 38.780 ;
        RECT 94.835 38.150 95.125 38.340 ;
        RECT 94.205 37.600 94.825 37.960 ;
        RECT 96.245 37.630 96.935 38.340 ;
        RECT 93.425 36.440 93.805 37.040 ;
        RECT 94.215 36.730 94.645 37.600 ;
        RECT 93.495 35.250 93.725 36.440 ;
        RECT 94.215 36.310 96.095 36.730 ;
        RECT 94.215 35.780 94.645 36.310 ;
        RECT 94.065 35.420 94.685 35.780 ;
        RECT 93.495 35.240 93.975 35.250 ;
        RECT 93.495 34.560 94.055 35.240 ;
        RECT 93.585 34.410 94.055 34.560 ;
        RECT 93.785 33.460 94.055 34.410 ;
        RECT 94.695 34.160 94.965 35.160 ;
        RECT 94.695 33.430 95.205 34.160 ;
        RECT 94.695 33.340 95.195 33.430 ;
        RECT 90.055 32.790 90.585 33.170 ;
        RECT 87.045 31.110 89.875 32.160 ;
        RECT 90.155 31.910 90.415 32.790 ;
        RECT 90.135 31.290 90.495 31.910 ;
        RECT 94.945 31.220 95.195 33.340 ;
        RECT 87.045 30.200 87.365 31.110 ;
        RECT 88.725 31.100 89.855 31.110 ;
        RECT 90.755 30.820 95.395 31.220 ;
        RECT 94.945 30.540 95.195 30.820 ;
        RECT 87.045 30.140 87.375 30.200 ;
        RECT 87.055 20.210 87.375 30.140 ;
        RECT 88.375 28.890 88.645 30.250 ;
        RECT 89.505 28.890 89.775 30.210 ;
        RECT 94.815 30.110 95.195 30.540 ;
        RECT 94.815 29.600 95.175 30.110 ;
        RECT 88.375 22.200 89.775 28.890 ;
        RECT 88.375 20.200 88.645 22.200 ;
        RECT 89.505 20.160 89.775 22.200 ;
        RECT 94.825 21.760 95.085 29.600 ;
        RECT 94.825 20.210 95.205 21.760 ;
        RECT 87.345 19.550 88.395 19.960 ;
        RECT 89.755 19.560 94.805 19.940 ;
        RECT 87.515 18.270 88.185 19.550 ;
        RECT 87.345 17.590 88.465 18.270 ;
        RECT 73.865 12.750 74.725 13.590 ;
        RECT 61.415 10.960 63.435 12.160 ;
        RECT 72.725 10.990 74.745 12.190 ;
        RECT 84.465 12.180 84.875 14.780 ;
        RECT 85.175 13.580 85.715 16.810 ;
        RECT 91.435 16.780 93.365 19.560 ;
        RECT 90.855 15.930 93.565 16.780 ;
        RECT 94.945 15.390 95.205 20.210 ;
        RECT 94.415 14.660 95.305 15.390 ;
        RECT 95.705 14.800 96.095 36.310 ;
        RECT 96.435 16.830 96.935 37.630 ;
        RECT 98.975 38.500 99.255 40.490 ;
        RECT 101.545 40.420 102.645 41.190 ;
        RECT 110.155 40.530 110.455 42.260 ;
        RECT 99.525 39.660 99.905 40.260 ;
        RECT 99.555 39.040 99.805 39.660 ;
        RECT 99.425 38.660 99.905 39.040 ;
        RECT 98.975 33.430 99.305 38.500 ;
        RECT 99.855 37.640 100.155 38.500 ;
        RECT 100.935 37.640 101.235 38.500 ;
        RECT 101.845 38.460 102.125 40.420 ;
        RECT 105.145 38.850 105.415 39.020 ;
        RECT 104.755 38.540 105.415 38.850 ;
        RECT 99.855 33.400 101.235 37.640 ;
        RECT 101.785 38.410 102.125 38.460 ;
        RECT 104.705 38.430 105.415 38.540 ;
        RECT 98.255 32.180 98.575 32.200 ;
        RECT 99.935 32.180 101.065 33.400 ;
        RECT 101.785 33.390 102.115 38.410 ;
        RECT 104.705 37.060 104.935 38.430 ;
        RECT 105.145 38.180 105.415 38.430 ;
        RECT 106.045 38.800 106.335 39.040 ;
        RECT 107.455 38.800 108.145 38.820 ;
        RECT 106.045 38.360 108.145 38.800 ;
        RECT 106.045 38.170 106.335 38.360 ;
        RECT 105.415 37.620 106.035 37.980 ;
        RECT 107.455 37.650 108.145 38.360 ;
        RECT 104.635 36.460 105.015 37.060 ;
        RECT 105.425 36.750 105.855 37.620 ;
        RECT 104.705 35.270 104.935 36.460 ;
        RECT 105.425 36.330 107.305 36.750 ;
        RECT 105.425 35.800 105.855 36.330 ;
        RECT 105.275 35.440 105.895 35.800 ;
        RECT 104.705 35.260 105.185 35.270 ;
        RECT 104.705 34.580 105.265 35.260 ;
        RECT 104.795 34.430 105.265 34.580 ;
        RECT 104.995 33.480 105.265 34.430 ;
        RECT 105.905 34.180 106.175 35.180 ;
        RECT 105.905 33.450 106.415 34.180 ;
        RECT 105.905 33.360 106.405 33.450 ;
        RECT 101.265 32.810 101.795 33.190 ;
        RECT 98.255 31.130 101.085 32.180 ;
        RECT 101.365 31.930 101.625 32.810 ;
        RECT 101.345 31.310 101.705 31.930 ;
        RECT 106.155 31.240 106.405 33.360 ;
        RECT 98.255 30.220 98.575 31.130 ;
        RECT 99.935 31.120 101.065 31.130 ;
        RECT 101.965 30.840 106.605 31.240 ;
        RECT 106.155 30.560 106.405 30.840 ;
        RECT 98.255 30.160 98.585 30.220 ;
        RECT 98.265 20.230 98.585 30.160 ;
        RECT 99.585 28.910 99.855 30.270 ;
        RECT 100.715 28.910 100.985 30.230 ;
        RECT 106.025 30.130 106.405 30.560 ;
        RECT 106.025 29.620 106.385 30.130 ;
        RECT 99.585 22.220 100.985 28.910 ;
        RECT 99.585 20.220 99.855 22.220 ;
        RECT 100.715 20.180 100.985 22.220 ;
        RECT 106.035 21.780 106.295 29.620 ;
        RECT 106.035 20.230 106.415 21.780 ;
        RECT 98.555 19.570 99.605 19.980 ;
        RECT 100.965 19.580 106.015 19.960 ;
        RECT 98.725 18.290 99.395 19.570 ;
        RECT 98.555 17.610 99.675 18.290 ;
        RECT 85.155 12.740 86.015 13.580 ;
        RECT 95.705 12.180 96.115 14.800 ;
        RECT 96.415 13.600 96.955 16.830 ;
        RECT 102.645 16.800 104.575 19.580 ;
        RECT 102.065 15.950 104.775 16.800 ;
        RECT 106.155 15.410 106.415 20.230 ;
        RECT 105.625 14.680 106.515 15.410 ;
        RECT 106.915 14.820 107.305 36.330 ;
        RECT 107.645 16.850 108.145 37.650 ;
        RECT 110.175 38.540 110.455 40.530 ;
        RECT 112.745 40.460 113.845 41.230 ;
        RECT 121.365 40.550 121.665 42.280 ;
        RECT 142.880 42.020 144.100 43.390 ;
        RECT 110.725 39.700 111.105 40.300 ;
        RECT 110.755 39.080 111.005 39.700 ;
        RECT 110.625 38.700 111.105 39.080 ;
        RECT 110.175 33.470 110.505 38.540 ;
        RECT 111.055 37.680 111.355 38.540 ;
        RECT 112.135 37.680 112.435 38.540 ;
        RECT 113.045 38.500 113.325 40.460 ;
        RECT 116.345 38.890 116.615 39.060 ;
        RECT 115.955 38.580 116.615 38.890 ;
        RECT 111.055 33.440 112.435 37.680 ;
        RECT 112.985 38.450 113.325 38.500 ;
        RECT 115.905 38.470 116.615 38.580 ;
        RECT 109.455 32.220 109.775 32.240 ;
        RECT 111.135 32.220 112.265 33.440 ;
        RECT 112.985 33.430 113.315 38.450 ;
        RECT 115.905 37.100 116.135 38.470 ;
        RECT 116.345 38.220 116.615 38.470 ;
        RECT 117.245 38.840 117.535 39.080 ;
        RECT 118.655 38.840 119.345 38.860 ;
        RECT 117.245 38.400 119.345 38.840 ;
        RECT 117.245 38.210 117.535 38.400 ;
        RECT 116.615 37.660 117.235 38.020 ;
        RECT 118.655 37.690 119.345 38.400 ;
        RECT 115.835 36.500 116.215 37.100 ;
        RECT 116.625 36.790 117.055 37.660 ;
        RECT 115.905 35.310 116.135 36.500 ;
        RECT 116.625 36.370 118.505 36.790 ;
        RECT 116.625 35.840 117.055 36.370 ;
        RECT 116.475 35.480 117.095 35.840 ;
        RECT 115.905 35.300 116.385 35.310 ;
        RECT 115.905 34.620 116.465 35.300 ;
        RECT 115.995 34.470 116.465 34.620 ;
        RECT 116.195 33.520 116.465 34.470 ;
        RECT 117.105 34.220 117.375 35.220 ;
        RECT 117.105 33.490 117.615 34.220 ;
        RECT 117.105 33.400 117.605 33.490 ;
        RECT 112.465 32.850 112.995 33.230 ;
        RECT 109.455 31.170 112.285 32.220 ;
        RECT 112.565 31.970 112.825 32.850 ;
        RECT 112.545 31.350 112.905 31.970 ;
        RECT 117.355 31.280 117.605 33.400 ;
        RECT 109.455 30.260 109.775 31.170 ;
        RECT 111.135 31.160 112.265 31.170 ;
        RECT 113.165 30.880 117.805 31.280 ;
        RECT 117.355 30.600 117.605 30.880 ;
        RECT 109.455 30.200 109.785 30.260 ;
        RECT 109.465 20.270 109.785 30.200 ;
        RECT 110.785 28.950 111.055 30.310 ;
        RECT 111.915 28.950 112.185 30.270 ;
        RECT 117.225 30.170 117.605 30.600 ;
        RECT 117.225 29.660 117.585 30.170 ;
        RECT 110.785 22.260 112.185 28.950 ;
        RECT 110.785 20.260 111.055 22.260 ;
        RECT 111.915 20.220 112.185 22.260 ;
        RECT 117.235 21.820 117.495 29.660 ;
        RECT 117.235 20.270 117.615 21.820 ;
        RECT 109.755 19.610 110.805 20.020 ;
        RECT 112.165 19.620 117.215 20.000 ;
        RECT 109.925 18.330 110.595 19.610 ;
        RECT 109.755 17.650 110.875 18.330 ;
        RECT 96.395 12.760 97.255 13.600 ;
        RECT 106.915 12.230 107.325 14.820 ;
        RECT 107.625 13.620 108.165 16.850 ;
        RECT 113.845 16.840 115.775 19.620 ;
        RECT 113.265 15.990 115.975 16.840 ;
        RECT 117.355 15.450 117.615 20.270 ;
        RECT 116.825 14.720 117.715 15.450 ;
        RECT 118.115 14.860 118.505 36.370 ;
        RECT 118.845 16.890 119.345 37.690 ;
        RECT 121.385 38.560 121.665 40.550 ;
        RECT 123.955 40.480 125.055 41.250 ;
        RECT 121.935 39.720 122.315 40.320 ;
        RECT 121.965 39.100 122.215 39.720 ;
        RECT 121.835 38.720 122.315 39.100 ;
        RECT 121.385 33.490 121.715 38.560 ;
        RECT 122.265 37.700 122.565 38.560 ;
        RECT 123.345 37.700 123.645 38.560 ;
        RECT 124.255 38.520 124.535 40.480 ;
        RECT 127.555 38.910 127.825 39.080 ;
        RECT 127.165 38.600 127.825 38.910 ;
        RECT 122.265 33.460 123.645 37.700 ;
        RECT 124.195 38.470 124.535 38.520 ;
        RECT 127.115 38.490 127.825 38.600 ;
        RECT 120.665 32.240 120.985 32.260 ;
        RECT 122.345 32.240 123.475 33.460 ;
        RECT 124.195 33.450 124.525 38.470 ;
        RECT 127.115 37.120 127.345 38.490 ;
        RECT 127.555 38.240 127.825 38.490 ;
        RECT 128.455 38.860 128.745 39.100 ;
        RECT 142.940 38.950 144.100 42.020 ;
        RECT 129.865 38.860 130.555 38.880 ;
        RECT 128.455 38.420 130.555 38.860 ;
        RECT 128.455 38.230 128.745 38.420 ;
        RECT 127.825 37.680 128.445 38.040 ;
        RECT 129.865 37.710 130.555 38.420 ;
        RECT 127.045 36.520 127.425 37.120 ;
        RECT 127.835 36.810 128.265 37.680 ;
        RECT 127.115 35.330 127.345 36.520 ;
        RECT 127.835 36.390 129.715 36.810 ;
        RECT 127.835 35.860 128.265 36.390 ;
        RECT 127.685 35.500 128.305 35.860 ;
        RECT 127.115 35.320 127.595 35.330 ;
        RECT 127.115 34.640 127.675 35.320 ;
        RECT 127.205 34.490 127.675 34.640 ;
        RECT 127.405 33.540 127.675 34.490 ;
        RECT 128.315 34.240 128.585 35.240 ;
        RECT 128.315 33.510 128.825 34.240 ;
        RECT 128.315 33.420 128.815 33.510 ;
        RECT 123.675 32.870 124.205 33.250 ;
        RECT 120.665 31.190 123.495 32.240 ;
        RECT 123.775 31.990 124.035 32.870 ;
        RECT 123.755 31.370 124.115 31.990 ;
        RECT 128.565 31.300 128.815 33.420 ;
        RECT 120.665 30.280 120.985 31.190 ;
        RECT 122.345 31.180 123.475 31.190 ;
        RECT 124.375 30.900 129.015 31.300 ;
        RECT 128.565 30.620 128.815 30.900 ;
        RECT 120.665 30.220 120.995 30.280 ;
        RECT 120.675 20.290 120.995 30.220 ;
        RECT 121.995 28.970 122.265 30.330 ;
        RECT 123.125 28.970 123.395 30.290 ;
        RECT 128.435 30.190 128.815 30.620 ;
        RECT 128.435 29.680 128.795 30.190 ;
        RECT 121.995 22.280 123.395 28.970 ;
        RECT 121.995 20.280 122.265 22.280 ;
        RECT 123.125 20.240 123.395 22.280 ;
        RECT 128.445 21.840 128.705 29.680 ;
        RECT 128.445 20.290 128.825 21.840 ;
        RECT 120.965 19.630 122.015 20.040 ;
        RECT 123.375 19.640 128.425 20.020 ;
        RECT 121.135 18.350 121.805 19.630 ;
        RECT 120.965 17.670 122.085 18.350 ;
        RECT 107.605 12.780 108.465 13.620 ;
        RECT 118.115 12.230 118.525 14.860 ;
        RECT 118.825 13.660 119.365 16.890 ;
        RECT 125.055 16.860 126.985 19.640 ;
        RECT 124.475 16.010 127.185 16.860 ;
        RECT 128.565 15.470 128.825 20.290 ;
        RECT 128.035 14.740 128.925 15.470 ;
        RECT 129.325 14.880 129.715 36.390 ;
        RECT 130.055 16.910 130.555 37.710 ;
        RECT 142.900 37.580 144.120 38.950 ;
        RECT 132.395 24.340 132.705 30.230 ;
        RECT 132.195 20.120 132.705 24.340 ;
        RECT 118.805 12.820 119.665 13.660 ;
        RECT 129.325 12.260 129.735 14.880 ;
        RECT 130.035 13.680 130.575 16.910 ;
        RECT 132.195 15.510 132.505 20.120 ;
        RECT 137.715 19.980 138.005 30.170 ;
        RECT 132.685 19.590 138.005 19.980 ;
        RECT 137.715 16.940 138.005 19.590 ;
        RECT 142.940 17.940 144.090 19.160 ;
        RECT 145.080 18.760 146.200 18.930 ;
        RECT 137.395 15.890 138.295 16.940 ;
        RECT 137.715 15.720 138.005 15.890 ;
        RECT 131.975 14.270 132.735 15.510 ;
        RECT 142.940 15.090 144.050 17.940 ;
        RECT 142.900 13.870 144.050 15.090 ;
        RECT 145.070 14.920 146.200 18.760 ;
        RECT 145.030 13.970 146.200 14.920 ;
        RECT 145.030 13.900 146.150 13.970 ;
        RECT 130.015 12.840 130.875 13.680 ;
        RECT 83.845 10.980 85.865 12.180 ;
        RECT 95.145 10.980 97.165 12.180 ;
        RECT 106.335 11.030 108.355 12.230 ;
        RECT 117.565 11.030 119.585 12.230 ;
        RECT 128.865 11.060 130.885 12.260 ;
        RECT 74.340 0.110 75.630 1.460 ;
        RECT 93.550 0.180 94.840 1.530 ;
        RECT 112.950 0.310 114.240 1.660 ;
        RECT 131.850 0.380 133.490 1.930 ;
        RECT 151.650 0.250 152.920 1.470 ;
      LAYER met3 ;
        RECT 135.340 223.855 136.790 225.205 ;
        RECT 138.130 223.785 139.580 225.135 ;
        RECT 143.180 223.815 144.630 225.165 ;
        RECT 16.830 211.125 18.810 211.455 ;
        RECT 46.830 211.125 48.810 211.455 ;
        RECT 76.830 211.125 78.810 211.455 ;
        RECT 106.830 211.125 108.810 211.455 ;
        RECT 31.830 208.405 33.810 208.735 ;
        RECT 61.830 208.405 63.810 208.735 ;
        RECT 91.830 208.405 93.810 208.735 ;
        RECT 121.830 208.405 123.810 208.735 ;
        RECT 16.830 205.685 18.810 206.015 ;
        RECT 46.830 205.685 48.810 206.015 ;
        RECT 76.830 205.685 78.810 206.015 ;
        RECT 106.830 205.685 108.810 206.015 ;
        RECT 31.830 202.965 33.810 203.295 ;
        RECT 61.830 202.965 63.810 203.295 ;
        RECT 91.830 202.965 93.810 203.295 ;
        RECT 121.830 202.965 123.810 203.295 ;
        RECT 16.830 200.245 18.810 200.575 ;
        RECT 46.830 200.245 48.810 200.575 ;
        RECT 76.830 200.245 78.810 200.575 ;
        RECT 106.830 200.245 108.810 200.575 ;
        RECT 31.830 197.525 33.810 197.855 ;
        RECT 61.830 197.525 63.810 197.855 ;
        RECT 91.830 197.525 93.810 197.855 ;
        RECT 121.830 197.525 123.810 197.855 ;
        RECT 16.830 194.805 18.810 195.135 ;
        RECT 46.830 194.805 48.810 195.135 ;
        RECT 76.830 194.805 78.810 195.135 ;
        RECT 106.830 194.805 108.810 195.135 ;
        RECT 31.830 192.085 33.810 192.415 ;
        RECT 61.830 192.085 63.810 192.415 ;
        RECT 91.830 192.085 93.810 192.415 ;
        RECT 121.830 192.085 123.810 192.415 ;
        RECT 16.830 189.365 18.810 189.695 ;
        RECT 46.830 189.365 48.810 189.695 ;
        RECT 76.830 189.365 78.810 189.695 ;
        RECT 106.830 189.365 108.810 189.695 ;
        RECT 31.830 186.645 33.810 186.975 ;
        RECT 61.830 186.645 63.810 186.975 ;
        RECT 91.830 186.645 93.810 186.975 ;
        RECT 121.830 186.645 123.810 186.975 ;
        RECT 84.185 184.590 84.515 184.595 ;
        RECT 83.930 184.580 84.515 184.590 ;
        RECT 83.930 184.280 84.740 184.580 ;
        RECT 83.930 184.270 84.515 184.280 ;
        RECT 84.185 184.265 84.515 184.270 ;
        RECT 16.830 183.925 18.810 184.255 ;
        RECT 46.830 183.925 48.810 184.255 ;
        RECT 76.830 183.925 78.810 184.255 ;
        RECT 106.830 183.925 108.810 184.255 ;
        RECT 31.830 181.205 33.810 181.535 ;
        RECT 61.830 181.205 63.810 181.535 ;
        RECT 91.830 181.205 93.810 181.535 ;
        RECT 121.830 181.205 123.810 181.535 ;
        RECT 16.830 178.485 18.810 178.815 ;
        RECT 46.830 178.485 48.810 178.815 ;
        RECT 76.830 178.485 78.810 178.815 ;
        RECT 106.830 178.485 108.810 178.815 ;
        RECT 79.585 177.780 79.915 177.795 ;
        RECT 101.665 177.780 101.995 177.795 ;
        RECT 79.585 177.480 101.995 177.780 ;
        RECT 79.585 177.465 79.915 177.480 ;
        RECT 101.665 177.465 101.995 177.480 ;
        RECT 31.830 175.765 33.810 176.095 ;
        RECT 61.830 175.765 63.810 176.095 ;
        RECT 91.830 175.765 93.810 176.095 ;
        RECT 121.830 175.765 123.810 176.095 ;
        RECT 64.610 174.380 64.990 174.390 ;
        RECT 79.585 174.380 79.915 174.395 ;
        RECT 64.610 174.080 79.915 174.380 ;
        RECT 64.610 174.070 64.990 174.080 ;
        RECT 79.585 174.065 79.915 174.080 ;
        RECT 16.830 173.045 18.810 173.375 ;
        RECT 46.830 173.045 48.810 173.375 ;
        RECT 76.830 173.045 78.810 173.375 ;
        RECT 106.830 173.045 108.810 173.375 ;
        RECT 133.920 172.090 134.760 172.195 ;
        RECT 130.230 171.675 134.830 172.090 ;
        RECT 130.185 171.345 134.830 171.675 ;
        RECT 31.830 170.325 33.810 170.655 ;
        RECT 61.830 170.325 63.810 170.655 ;
        RECT 91.830 170.325 93.810 170.655 ;
        RECT 121.830 170.325 123.810 170.655 ;
        RECT 130.230 170.500 134.830 171.345 ;
        RECT 106.265 169.620 106.595 169.635 ;
        RECT 106.050 169.305 106.595 169.620 ;
        RECT 34.965 168.940 35.295 168.955 ;
        RECT 50.605 168.940 50.935 168.955 ;
        RECT 64.610 168.940 64.990 168.950 ;
        RECT 34.965 168.640 64.990 168.940 ;
        RECT 34.965 168.625 35.295 168.640 ;
        RECT 50.605 168.625 50.935 168.640 ;
        RECT 64.610 168.630 64.990 168.640 ;
        RECT 45.290 168.260 45.670 168.270 ;
        RECT 46.005 168.260 46.335 168.275 ;
        RECT 45.290 167.960 46.335 168.260 ;
        RECT 45.290 167.950 45.670 167.960 ;
        RECT 46.005 167.945 46.335 167.960 ;
        RECT 16.830 167.605 18.810 167.935 ;
        RECT 46.830 167.605 48.810 167.935 ;
        RECT 76.830 167.605 78.810 167.935 ;
        RECT 106.050 166.915 106.350 169.305 ;
        RECT 106.830 167.605 108.810 167.935 ;
        RECT 50.145 166.900 50.475 166.915 ;
        RECT 67.165 166.900 67.495 166.915 ;
        RECT 79.585 166.900 79.915 166.915 ;
        RECT 81.885 166.900 82.215 166.915 ;
        RECT 50.145 166.600 82.215 166.900 ;
        RECT 50.145 166.585 50.475 166.600 ;
        RECT 67.165 166.585 67.495 166.600 ;
        RECT 79.585 166.585 79.915 166.600 ;
        RECT 81.885 166.585 82.215 166.600 ;
        RECT 105.805 166.600 106.350 166.915 ;
        RECT 105.805 166.585 106.135 166.600 ;
        RECT 31.830 164.885 33.810 165.215 ;
        RECT 61.830 164.885 63.810 165.215 ;
        RECT 91.830 164.885 93.810 165.215 ;
        RECT 121.830 164.885 123.810 165.215 ;
        RECT 16.830 162.165 18.810 162.495 ;
        RECT 46.830 162.165 48.810 162.495 ;
        RECT 76.830 162.165 78.810 162.495 ;
        RECT 106.830 162.165 108.810 162.495 ;
        RECT 82.090 160.780 82.470 160.790 ;
        RECT 83.265 160.780 83.595 160.795 ;
        RECT 82.090 160.480 83.595 160.780 ;
        RECT 82.090 160.470 82.470 160.480 ;
        RECT 83.265 160.465 83.595 160.480 ;
        RECT 31.830 159.445 33.810 159.775 ;
        RECT 61.830 159.445 63.810 159.775 ;
        RECT 91.830 159.445 93.810 159.775 ;
        RECT 121.830 159.445 123.810 159.775 ;
        RECT 49.685 158.060 50.015 158.075 ;
        RECT 53.825 158.060 54.155 158.075 ;
        RECT 77.285 158.060 77.615 158.075 ;
        RECT 49.685 157.760 77.615 158.060 ;
        RECT 49.685 157.745 50.015 157.760 ;
        RECT 53.825 157.745 54.155 157.760 ;
        RECT 77.285 157.745 77.615 157.760 ;
        RECT 16.830 156.725 18.810 157.055 ;
        RECT 46.830 156.725 48.810 157.055 ;
        RECT 76.830 156.725 78.810 157.055 ;
        RECT 106.830 156.725 108.810 157.055 ;
        RECT 59.805 156.020 60.135 156.035 ;
        RECT 61.185 156.020 61.515 156.035 ;
        RECT 59.805 155.720 61.515 156.020 ;
        RECT 59.805 155.705 60.135 155.720 ;
        RECT 61.185 155.705 61.515 155.720 ;
        RECT 43.705 155.340 44.035 155.355 ;
        RECT 62.565 155.340 62.895 155.355 ;
        RECT 43.705 155.040 62.895 155.340 ;
        RECT 43.705 155.025 44.035 155.040 ;
        RECT 62.565 155.025 62.895 155.040 ;
        RECT 31.830 154.005 33.810 154.335 ;
        RECT 61.830 154.005 63.810 154.335 ;
        RECT 91.830 154.005 93.810 154.335 ;
        RECT 121.830 154.005 123.810 154.335 ;
        RECT 46.925 153.300 47.255 153.315 ;
        RECT 46.250 153.000 47.255 153.300 ;
        RECT 45.545 152.620 45.875 152.635 ;
        RECT 46.250 152.620 46.550 153.000 ;
        RECT 46.925 152.985 47.255 153.000 ;
        RECT 49.685 153.300 50.015 153.315 ;
        RECT 52.905 153.300 53.235 153.315 ;
        RECT 49.685 153.000 53.235 153.300 ;
        RECT 49.685 152.985 50.015 153.000 ;
        RECT 52.905 152.985 53.235 153.000 ;
        RECT 45.545 152.320 46.550 152.620 ;
        RECT 46.925 152.620 47.255 152.635 ;
        RECT 49.685 152.620 50.015 152.635 ;
        RECT 46.925 152.320 50.015 152.620 ;
        RECT 45.545 152.305 45.875 152.320 ;
        RECT 46.925 152.305 47.255 152.320 ;
        RECT 49.685 152.305 50.015 152.320 ;
        RECT 99.365 152.620 99.695 152.635 ;
        RECT 107.645 152.620 107.975 152.635 ;
        RECT 99.365 152.320 107.975 152.620 ;
        RECT 99.365 152.305 99.695 152.320 ;
        RECT 107.645 152.305 107.975 152.320 ;
        RECT 49.225 151.940 49.555 151.955 ;
        RECT 53.825 151.940 54.155 151.955 ;
        RECT 49.225 151.640 54.155 151.940 ;
        RECT 49.225 151.625 49.555 151.640 ;
        RECT 53.825 151.625 54.155 151.640 ;
        RECT 16.830 151.285 18.810 151.615 ;
        RECT 46.830 151.285 48.810 151.615 ;
        RECT 76.830 151.285 78.810 151.615 ;
        RECT 106.830 151.285 108.810 151.615 ;
        RECT 64.865 149.230 65.195 149.235 ;
        RECT 64.610 149.220 65.195 149.230 ;
        RECT 76.825 149.220 77.155 149.235 ;
        RECT 82.345 149.220 82.675 149.235 ;
        RECT 64.610 148.920 65.420 149.220 ;
        RECT 76.825 148.920 82.675 149.220 ;
        RECT 64.610 148.910 65.195 148.920 ;
        RECT 64.865 148.905 65.195 148.910 ;
        RECT 76.825 148.905 77.155 148.920 ;
        RECT 82.345 148.905 82.675 148.920 ;
        RECT 31.830 148.565 33.810 148.895 ;
        RECT 61.830 148.565 63.810 148.895 ;
        RECT 91.830 148.565 93.810 148.895 ;
        RECT 121.830 148.565 123.810 148.895 ;
        RECT 72.225 146.500 72.555 146.515 ;
        RECT 75.650 146.500 76.030 146.510 ;
        RECT 72.225 146.200 76.030 146.500 ;
        RECT 72.225 146.185 72.555 146.200 ;
        RECT 75.650 146.190 76.030 146.200 ;
        RECT 16.830 145.845 18.810 146.175 ;
        RECT 46.830 145.845 48.810 146.175 ;
        RECT 76.830 145.845 78.810 146.175 ;
        RECT 106.830 145.845 108.810 146.175 ;
        RECT 82.805 145.820 83.135 145.835 ;
        RECT 83.930 145.820 84.310 145.830 ;
        RECT 82.805 145.520 84.310 145.820 ;
        RECT 82.805 145.505 83.135 145.520 ;
        RECT 83.930 145.510 84.310 145.520 ;
        RECT 47.385 145.140 47.715 145.155 ;
        RECT 48.765 145.140 49.095 145.155 ;
        RECT 81.885 145.140 82.215 145.155 ;
        RECT 47.385 144.840 82.215 145.140 ;
        RECT 47.385 144.825 47.715 144.840 ;
        RECT 48.765 144.825 49.095 144.840 ;
        RECT 81.885 144.825 82.215 144.840 ;
        RECT 31.830 143.125 33.810 143.455 ;
        RECT 61.830 143.125 63.810 143.455 ;
        RECT 91.830 143.125 93.810 143.455 ;
        RECT 121.830 143.125 123.810 143.455 ;
        RECT 42.785 142.420 43.115 142.435 ;
        RECT 46.925 142.420 47.255 142.435 ;
        RECT 42.785 142.120 47.255 142.420 ;
        RECT 42.785 142.105 43.115 142.120 ;
        RECT 46.925 142.105 47.255 142.120 ;
        RECT 37.725 141.740 38.055 141.755 ;
        RECT 47.385 141.740 47.715 141.755 ;
        RECT 37.725 141.440 47.715 141.740 ;
        RECT 37.725 141.425 38.055 141.440 ;
        RECT 47.385 141.425 47.715 141.440 ;
        RECT 48.765 141.740 49.095 141.755 ;
        RECT 48.765 141.440 50.230 141.740 ;
        RECT 48.765 141.425 49.095 141.440 ;
        RECT 16.830 140.405 18.810 140.735 ;
        RECT 46.830 140.405 48.810 140.735 ;
        RECT 47.385 139.700 47.715 139.715 ;
        RECT 49.930 139.700 50.230 141.440 ;
        RECT 79.585 141.060 79.915 141.075 ;
        RECT 80.250 141.060 80.630 141.070 ;
        RECT 79.585 140.760 80.630 141.060 ;
        RECT 79.585 140.745 79.915 140.760 ;
        RECT 80.250 140.750 80.630 140.760 ;
        RECT 76.830 140.405 78.810 140.735 ;
        RECT 106.830 140.405 108.810 140.735 ;
        RECT 47.385 139.400 50.230 139.700 ;
        RECT 47.385 139.385 47.715 139.400 ;
        RECT 75.650 139.020 76.030 139.030 ;
        RECT 129.090 139.020 134.150 139.430 ;
        RECT 75.650 138.720 134.150 139.020 ;
        RECT 75.650 138.710 76.030 138.720 ;
        RECT 129.090 138.200 134.150 138.720 ;
        RECT 31.830 137.685 33.810 138.015 ;
        RECT 61.830 137.685 63.810 138.015 ;
        RECT 91.830 137.685 93.810 138.015 ;
        RECT 121.830 137.685 123.810 138.015 ;
        RECT 16.830 134.965 18.810 135.295 ;
        RECT 46.830 134.965 48.810 135.295 ;
        RECT 76.830 134.965 78.810 135.295 ;
        RECT 106.830 134.965 108.810 135.295 ;
        RECT 44.625 134.260 44.955 134.275 ;
        RECT 51.065 134.260 51.395 134.275 ;
        RECT 44.625 133.960 51.395 134.260 ;
        RECT 44.625 133.945 44.955 133.960 ;
        RECT 51.065 133.945 51.395 133.960 ;
        RECT 31.830 132.245 33.810 132.575 ;
        RECT 61.830 132.245 63.810 132.575 ;
        RECT 91.830 132.245 93.810 132.575 ;
        RECT 121.830 132.245 123.810 132.575 ;
        RECT 45.290 132.220 45.670 132.230 ;
        RECT 47.845 132.220 48.175 132.235 ;
        RECT 45.290 131.920 48.175 132.220 ;
        RECT 45.290 131.910 45.670 131.920 ;
        RECT 47.845 131.905 48.175 131.920 ;
        RECT 80.965 132.220 81.295 132.235 ;
        RECT 82.090 132.220 82.470 132.230 ;
        RECT 80.965 131.920 82.470 132.220 ;
        RECT 80.965 131.905 81.295 131.920 ;
        RECT 82.090 131.910 82.470 131.920 ;
        RECT 16.830 129.525 18.810 129.855 ;
        RECT 46.830 129.525 48.810 129.855 ;
        RECT 76.830 129.525 78.810 129.855 ;
        RECT 106.830 129.525 108.810 129.855 ;
        RECT 31.830 126.805 33.810 127.135 ;
        RECT 61.830 126.805 63.810 127.135 ;
        RECT 91.830 126.805 93.810 127.135 ;
        RECT 121.830 126.805 123.810 127.135 ;
        RECT 89.450 126.100 89.830 126.110 ;
        RECT 103.505 126.100 103.835 126.115 ;
        RECT 89.450 125.800 103.835 126.100 ;
        RECT 89.450 125.790 89.830 125.800 ;
        RECT 52.905 125.420 53.235 125.435 ;
        RECT 64.610 125.420 64.990 125.430 ;
        RECT 89.490 125.420 89.790 125.790 ;
        RECT 103.505 125.785 103.835 125.800 ;
        RECT 52.905 125.120 89.790 125.420 ;
        RECT 52.905 125.105 53.235 125.120 ;
        RECT 64.610 125.110 64.990 125.120 ;
        RECT 16.830 124.085 18.810 124.415 ;
        RECT 46.830 124.085 48.810 124.415 ;
        RECT 76.830 124.085 78.810 124.415 ;
        RECT 106.830 124.085 108.810 124.415 ;
        RECT 31.830 121.365 33.810 121.695 ;
        RECT 61.830 121.365 63.810 121.695 ;
        RECT 91.830 121.365 93.810 121.695 ;
        RECT 121.830 121.365 123.810 121.695 ;
        RECT 36.805 120.660 37.135 120.675 ;
        RECT 52.905 120.660 53.235 120.675 ;
        RECT 36.805 120.360 53.235 120.660 ;
        RECT 36.805 120.345 37.135 120.360 ;
        RECT 52.905 120.345 53.235 120.360 ;
        RECT 16.830 118.645 18.810 118.975 ;
        RECT 46.830 118.645 48.810 118.975 ;
        RECT 76.830 118.645 78.810 118.975 ;
        RECT 106.830 118.645 108.810 118.975 ;
        RECT 89.245 118.630 89.575 118.635 ;
        RECT 89.245 118.620 89.830 118.630 ;
        RECT 89.020 118.320 89.830 118.620 ;
        RECT 89.245 118.310 89.830 118.320 ;
        RECT 89.245 118.305 89.575 118.310 ;
        RECT 31.830 115.925 33.810 116.255 ;
        RECT 61.830 115.925 63.810 116.255 ;
        RECT 91.830 115.925 93.810 116.255 ;
        RECT 121.830 115.925 123.810 116.255 ;
        RECT 16.830 113.205 18.810 113.535 ;
        RECT 46.830 113.205 48.810 113.535 ;
        RECT 76.830 113.205 78.810 113.535 ;
        RECT 106.830 113.205 108.810 113.535 ;
        RECT 80.250 111.820 80.630 111.830 ;
        RECT 80.965 111.820 81.295 111.835 ;
        RECT 80.250 111.520 81.295 111.820 ;
        RECT 80.250 111.510 80.630 111.520 ;
        RECT 80.965 111.505 81.295 111.520 ;
        RECT 31.830 110.485 33.810 110.815 ;
        RECT 61.830 110.485 63.810 110.815 ;
        RECT 91.830 110.485 93.810 110.815 ;
        RECT 121.830 110.485 123.810 110.815 ;
        RECT 16.830 107.765 18.810 108.095 ;
        RECT 46.830 107.765 48.810 108.095 ;
        RECT 76.830 107.765 78.810 108.095 ;
        RECT 106.830 107.765 108.810 108.095 ;
        RECT 45.545 107.060 45.875 107.075 ;
        RECT 49.685 107.060 50.015 107.075 ;
        RECT 45.545 106.760 50.015 107.060 ;
        RECT 45.545 106.745 45.875 106.760 ;
        RECT 49.685 106.745 50.015 106.760 ;
        RECT 129.700 106.530 133.210 106.625 ;
        RECT 126.045 106.380 126.375 106.395 ;
        RECT 129.700 106.380 133.340 106.530 ;
        RECT 126.045 106.080 133.340 106.380 ;
        RECT 126.045 106.065 126.375 106.080 ;
        RECT 129.700 105.930 133.340 106.080 ;
        RECT 129.700 105.605 133.210 105.930 ;
        RECT 31.830 105.045 33.810 105.375 ;
        RECT 61.830 105.045 63.810 105.375 ;
        RECT 91.830 105.045 93.810 105.375 ;
        RECT 121.830 105.045 123.810 105.375 ;
        RECT 16.830 102.325 18.810 102.655 ;
        RECT 46.830 102.325 48.810 102.655 ;
        RECT 76.830 102.325 78.810 102.655 ;
        RECT 106.830 102.325 108.810 102.655 ;
        RECT 31.830 99.605 33.810 99.935 ;
        RECT 61.830 99.605 63.810 99.935 ;
        RECT 91.830 99.605 93.810 99.935 ;
        RECT 121.830 99.605 123.810 99.935 ;
        RECT 37.630 88.620 38.970 88.755 ;
        RECT 13.950 87.980 14.980 88.515 ;
        RECT 13.950 87.500 14.990 87.980 ;
        RECT 13.950 87.175 14.980 87.500 ;
        RECT 14.070 86.570 14.810 87.175 ;
        RECT 20.050 87.105 20.920 88.515 ;
        RECT 14.070 75.715 14.700 86.570 ;
        RECT 20.170 77.115 20.800 87.105 ;
        RECT 25.910 87.055 26.860 88.515 ;
        RECT 26.070 78.385 26.700 87.055 ;
        RECT 31.730 86.965 32.910 88.585 ;
        RECT 32.005 79.615 32.635 86.965 ;
        RECT 37.630 86.835 39.120 88.620 ;
        RECT 38.060 81.125 38.690 86.835 ;
        RECT 43.790 86.745 45.190 88.605 ;
        RECT 49.710 86.945 51.060 88.615 ;
        RECT 44.175 82.625 44.805 86.745 ;
        RECT 50.070 83.875 50.700 86.945 ;
        RECT 55.530 86.785 56.750 88.545 ;
        RECT 55.825 85.115 56.455 86.785 ;
        RECT 61.670 86.625 63.180 88.615 ;
        RECT 67.680 88.305 68.720 89.815 ;
        RECT 67.885 87.225 68.515 88.305 ;
        RECT 62.110 86.175 62.740 86.625 ;
        RECT 67.885 86.595 130.605 87.225 ;
        RECT 62.110 85.545 118.855 86.175 ;
        RECT 55.825 84.485 107.605 85.115 ;
        RECT 50.070 83.245 96.285 83.875 ;
        RECT 44.175 81.995 85.055 82.625 ;
        RECT 38.060 80.495 73.765 81.125 ;
        RECT 32.005 78.985 62.635 79.615 ;
        RECT 26.070 77.755 51.245 78.385 ;
        RECT 20.170 76.485 40.645 77.115 ;
        RECT 14.070 75.660 29.295 75.715 ;
        RECT 40.015 75.710 40.645 76.485 ;
        RECT 14.070 75.085 30.410 75.660 ;
        RECT 27.850 74.670 30.410 75.085 ;
        RECT 3.910 71.345 6.100 73.215 ;
        RECT 27.850 73.120 30.450 74.670 ;
        RECT 39.060 74.510 41.620 75.710 ;
        RECT 50.615 75.580 51.245 77.755 ;
        RECT 62.005 75.690 62.635 78.985 ;
        RECT 49.930 74.650 52.490 75.580 ;
        RECT 0.970 70.330 3.070 70.430 ;
        RECT 15.510 70.330 17.040 71.185 ;
        RECT 0.960 68.750 17.040 70.330 ;
        RECT 0.970 68.710 3.070 68.750 ;
        RECT 15.510 68.635 17.040 68.750 ;
        RECT 20.145 54.060 20.605 54.135 ;
        RECT 25.715 54.060 26.175 54.085 ;
        RECT 20.145 53.620 26.175 54.060 ;
        RECT 20.145 53.565 20.605 53.620 ;
        RECT 25.715 53.515 26.175 53.620 ;
        RECT 22.405 48.870 22.885 48.935 ;
        RECT 22.405 48.550 24.205 48.870 ;
        RECT 22.405 48.385 22.885 48.550 ;
        RECT 23.635 45.710 24.195 48.550 ;
        RECT 27.515 45.710 27.995 45.735 ;
        RECT 23.635 45.290 27.995 45.710 ;
        RECT 23.635 45.280 24.195 45.290 ;
        RECT 27.515 45.185 27.995 45.290 ;
        RECT 20.745 40.120 21.225 40.225 ;
        RECT 24.545 40.120 25.105 40.130 ;
        RECT 20.745 39.700 25.105 40.120 ;
        RECT 20.745 39.675 21.225 39.700 ;
        RECT 24.545 36.860 25.105 39.700 ;
        RECT 25.855 36.860 26.335 37.025 ;
        RECT 24.535 36.540 26.335 36.860 ;
        RECT 25.855 36.475 26.335 36.540 ;
        RECT 22.565 31.790 23.025 31.895 ;
        RECT 28.135 31.790 28.595 31.845 ;
        RECT 22.565 31.350 28.595 31.790 ;
        RECT 22.565 31.325 23.025 31.350 ;
        RECT 28.135 31.275 28.595 31.350 ;
        RECT 29.765 12.265 30.255 73.120 ;
        RECT 38.960 73.080 41.730 74.510 ;
        RECT 31.345 54.070 31.805 54.145 ;
        RECT 36.915 54.070 37.375 54.095 ;
        RECT 31.345 53.630 37.375 54.070 ;
        RECT 31.345 53.575 31.805 53.630 ;
        RECT 36.915 53.525 37.375 53.630 ;
        RECT 33.605 48.880 34.085 48.945 ;
        RECT 33.605 48.560 35.405 48.880 ;
        RECT 33.605 48.395 34.085 48.560 ;
        RECT 34.835 45.720 35.395 48.560 ;
        RECT 38.715 45.720 39.195 45.745 ;
        RECT 34.835 45.300 39.195 45.720 ;
        RECT 34.835 45.290 35.395 45.300 ;
        RECT 38.715 45.195 39.195 45.300 ;
        RECT 32.025 40.120 32.505 40.225 ;
        RECT 35.825 40.120 36.385 40.130 ;
        RECT 32.025 39.700 36.385 40.120 ;
        RECT 32.025 39.675 32.505 39.700 ;
        RECT 35.825 36.860 36.385 39.700 ;
        RECT 37.135 36.860 37.615 37.025 ;
        RECT 35.815 36.540 37.615 36.860 ;
        RECT 37.135 36.475 37.615 36.540 ;
        RECT 33.845 31.790 34.305 31.895 ;
        RECT 39.415 31.790 39.875 31.845 ;
        RECT 33.845 31.350 39.875 31.790 ;
        RECT 33.845 31.325 34.305 31.350 ;
        RECT 39.415 31.275 39.875 31.350 ;
        RECT 41.055 12.360 41.545 73.080 ;
        RECT 49.930 73.030 52.530 74.650 ;
        RECT 61.330 74.530 63.890 75.690 ;
        RECT 73.135 75.580 73.765 80.495 ;
        RECT 84.425 75.690 85.055 81.995 ;
        RECT 72.340 74.980 74.900 75.580 ;
        RECT 42.565 54.040 43.025 54.115 ;
        RECT 48.135 54.040 48.595 54.065 ;
        RECT 42.565 53.600 48.595 54.040 ;
        RECT 42.565 53.545 43.025 53.600 ;
        RECT 48.135 53.495 48.595 53.600 ;
        RECT 44.825 48.850 45.305 48.915 ;
        RECT 44.825 48.530 46.625 48.850 ;
        RECT 44.825 48.365 45.305 48.530 ;
        RECT 46.055 45.690 46.615 48.530 ;
        RECT 49.935 45.690 50.415 45.715 ;
        RECT 46.055 45.270 50.415 45.690 ;
        RECT 46.055 45.260 46.615 45.270 ;
        RECT 49.935 45.165 50.415 45.270 ;
        RECT 43.315 40.100 43.795 40.205 ;
        RECT 47.115 40.100 47.675 40.110 ;
        RECT 43.315 39.680 47.675 40.100 ;
        RECT 43.315 39.655 43.795 39.680 ;
        RECT 47.115 36.840 47.675 39.680 ;
        RECT 48.425 36.840 48.905 37.005 ;
        RECT 47.105 36.520 48.905 36.840 ;
        RECT 48.425 36.455 48.905 36.520 ;
        RECT 45.135 31.770 45.595 31.875 ;
        RECT 50.705 31.770 51.165 31.825 ;
        RECT 45.135 31.330 51.165 31.770 ;
        RECT 45.135 31.305 45.595 31.330 ;
        RECT 50.705 31.255 51.165 31.330 ;
        RECT 41.055 12.350 41.555 12.360 ;
        RECT 28.345 11.115 30.465 12.265 ;
        RECT 41.065 11.965 41.555 12.350 ;
        RECT 51.635 12.145 52.125 73.030 ;
        RECT 61.260 73.010 64.060 74.530 ;
        RECT 72.340 73.050 75.020 74.980 ;
        RECT 83.730 74.540 86.290 75.690 ;
        RECT 95.655 75.580 96.285 83.245 ;
        RECT 106.975 75.640 107.605 84.485 ;
        RECT 118.225 75.650 118.855 85.545 ;
        RECT 129.975 75.650 130.605 86.595 ;
        RECT 133.330 76.605 136.060 77.855 ;
        RECT 137.190 76.585 139.920 77.835 ;
        RECT 53.815 54.020 54.275 54.095 ;
        RECT 59.385 54.020 59.845 54.045 ;
        RECT 53.815 53.580 59.845 54.020 ;
        RECT 53.815 53.525 54.275 53.580 ;
        RECT 59.385 53.475 59.845 53.580 ;
        RECT 56.075 48.830 56.555 48.895 ;
        RECT 56.075 48.510 57.875 48.830 ;
        RECT 56.075 48.345 56.555 48.510 ;
        RECT 57.305 45.670 57.865 48.510 ;
        RECT 61.185 45.670 61.665 45.695 ;
        RECT 57.305 45.250 61.665 45.670 ;
        RECT 57.305 45.240 57.865 45.250 ;
        RECT 61.185 45.145 61.665 45.250 ;
        RECT 54.535 40.100 55.015 40.205 ;
        RECT 58.335 40.100 58.895 40.110 ;
        RECT 54.535 39.680 58.895 40.100 ;
        RECT 54.535 39.655 55.015 39.680 ;
        RECT 58.335 36.840 58.895 39.680 ;
        RECT 59.645 36.840 60.125 37.005 ;
        RECT 58.325 36.520 60.125 36.840 ;
        RECT 59.645 36.455 60.125 36.520 ;
        RECT 56.355 31.770 56.815 31.875 ;
        RECT 61.925 31.770 62.385 31.825 ;
        RECT 56.355 31.330 62.385 31.770 ;
        RECT 56.355 31.305 56.815 31.330 ;
        RECT 61.925 31.255 62.385 31.330 ;
        RECT 29.765 11.100 30.255 11.115 ;
        RECT 39.065 11.005 41.615 11.965 ;
        RECT 50.285 10.995 52.405 12.145 ;
        RECT 62.915 12.135 63.405 73.010 ;
        RECT 65.035 54.010 65.495 54.085 ;
        RECT 70.605 54.010 71.065 54.035 ;
        RECT 65.035 53.570 71.065 54.010 ;
        RECT 65.035 53.515 65.495 53.570 ;
        RECT 70.605 53.465 71.065 53.570 ;
        RECT 67.295 48.820 67.775 48.885 ;
        RECT 67.295 48.500 69.095 48.820 ;
        RECT 67.295 48.335 67.775 48.500 ;
        RECT 68.525 45.660 69.085 48.500 ;
        RECT 72.405 45.660 72.885 45.685 ;
        RECT 68.525 45.240 72.885 45.660 ;
        RECT 68.525 45.230 69.085 45.240 ;
        RECT 72.405 45.135 72.885 45.240 ;
        RECT 65.735 40.100 66.215 40.205 ;
        RECT 69.535 40.100 70.095 40.110 ;
        RECT 65.735 39.680 70.095 40.100 ;
        RECT 65.735 39.655 66.215 39.680 ;
        RECT 69.535 36.840 70.095 39.680 ;
        RECT 70.845 36.840 71.325 37.005 ;
        RECT 69.525 36.520 71.325 36.840 ;
        RECT 70.845 36.455 71.325 36.520 ;
        RECT 67.555 31.770 68.015 31.875 ;
        RECT 73.125 31.770 73.585 31.825 ;
        RECT 67.555 31.330 73.585 31.770 ;
        RECT 67.555 31.305 68.015 31.330 ;
        RECT 73.125 31.255 73.585 31.330 ;
        RECT 74.055 12.165 74.545 73.050 ;
        RECT 83.690 73.000 86.290 74.540 ;
        RECT 94.960 74.710 97.520 75.580 ;
        RECT 94.960 73.020 97.570 74.710 ;
        RECT 106.340 74.460 108.900 75.640 ;
        RECT 117.470 74.720 120.030 75.650 ;
        RECT 76.275 54.000 76.735 54.075 ;
        RECT 81.845 54.000 82.305 54.025 ;
        RECT 76.275 53.560 82.305 54.000 ;
        RECT 76.275 53.505 76.735 53.560 ;
        RECT 81.845 53.455 82.305 53.560 ;
        RECT 78.535 48.810 79.015 48.875 ;
        RECT 78.535 48.490 80.335 48.810 ;
        RECT 78.535 48.325 79.015 48.490 ;
        RECT 79.765 45.650 80.325 48.490 ;
        RECT 83.645 45.650 84.125 45.675 ;
        RECT 79.765 45.230 84.125 45.650 ;
        RECT 79.765 45.220 80.325 45.230 ;
        RECT 83.645 45.125 84.125 45.230 ;
        RECT 77.025 40.090 77.505 40.195 ;
        RECT 80.825 40.090 81.385 40.100 ;
        RECT 77.025 39.670 81.385 40.090 ;
        RECT 77.025 39.645 77.505 39.670 ;
        RECT 80.825 36.830 81.385 39.670 ;
        RECT 82.135 36.830 82.615 36.995 ;
        RECT 80.815 36.510 82.615 36.830 ;
        RECT 82.135 36.445 82.615 36.510 ;
        RECT 78.845 31.760 79.305 31.865 ;
        RECT 84.415 31.760 84.875 31.815 ;
        RECT 78.845 31.320 84.875 31.760 ;
        RECT 78.845 31.295 79.305 31.320 ;
        RECT 84.415 31.245 84.875 31.320 ;
        RECT 61.365 10.985 63.485 12.135 ;
        RECT 72.675 11.015 74.795 12.165 ;
        RECT 85.375 12.155 85.865 73.000 ;
        RECT 87.525 54.010 87.985 54.085 ;
        RECT 93.095 54.010 93.555 54.035 ;
        RECT 87.525 53.570 93.555 54.010 ;
        RECT 87.525 53.515 87.985 53.570 ;
        RECT 93.095 53.465 93.555 53.570 ;
        RECT 89.785 48.820 90.265 48.885 ;
        RECT 89.785 48.500 91.585 48.820 ;
        RECT 89.785 48.335 90.265 48.500 ;
        RECT 91.015 45.660 91.575 48.500 ;
        RECT 94.895 45.660 95.375 45.685 ;
        RECT 91.015 45.240 95.375 45.660 ;
        RECT 91.015 45.230 91.575 45.240 ;
        RECT 94.895 45.135 95.375 45.240 ;
        RECT 88.265 40.110 88.745 40.215 ;
        RECT 92.065 40.110 92.625 40.120 ;
        RECT 88.265 39.690 92.625 40.110 ;
        RECT 88.265 39.665 88.745 39.690 ;
        RECT 92.065 36.850 92.625 39.690 ;
        RECT 93.375 36.850 93.855 37.015 ;
        RECT 92.055 36.530 93.855 36.850 ;
        RECT 93.375 36.465 93.855 36.530 ;
        RECT 90.085 31.780 90.545 31.885 ;
        RECT 95.655 31.780 96.115 31.835 ;
        RECT 90.085 31.340 96.115 31.780 ;
        RECT 90.085 31.315 90.545 31.340 ;
        RECT 95.655 31.265 96.115 31.340 ;
        RECT 96.605 12.155 97.095 73.020 ;
        RECT 106.150 73.000 109.060 74.460 ;
        RECT 117.470 73.070 120.000 74.720 ;
        RECT 129.290 74.650 131.850 75.650 ;
        RECT 129.300 73.140 131.820 74.650 ;
        RECT 98.805 54.000 99.265 54.075 ;
        RECT 104.375 54.000 104.835 54.025 ;
        RECT 98.805 53.560 104.835 54.000 ;
        RECT 98.805 53.505 99.265 53.560 ;
        RECT 104.375 53.455 104.835 53.560 ;
        RECT 101.065 48.810 101.545 48.875 ;
        RECT 101.065 48.490 102.865 48.810 ;
        RECT 101.065 48.325 101.545 48.490 ;
        RECT 102.295 45.650 102.855 48.490 ;
        RECT 106.175 45.650 106.655 45.675 ;
        RECT 102.295 45.230 106.655 45.650 ;
        RECT 102.295 45.220 102.855 45.230 ;
        RECT 106.175 45.125 106.655 45.230 ;
        RECT 99.475 40.130 99.955 40.235 ;
        RECT 103.275 40.130 103.835 40.140 ;
        RECT 99.475 39.710 103.835 40.130 ;
        RECT 99.475 39.685 99.955 39.710 ;
        RECT 103.275 36.870 103.835 39.710 ;
        RECT 104.585 36.870 105.065 37.035 ;
        RECT 103.265 36.550 105.065 36.870 ;
        RECT 104.585 36.485 105.065 36.550 ;
        RECT 101.295 31.800 101.755 31.905 ;
        RECT 106.865 31.800 107.325 31.855 ;
        RECT 101.295 31.360 107.325 31.800 ;
        RECT 101.295 31.335 101.755 31.360 ;
        RECT 106.865 31.285 107.325 31.360 ;
        RECT 107.865 12.205 108.355 73.000 ;
        RECT 110.075 54.000 110.535 54.075 ;
        RECT 115.645 54.000 116.105 54.025 ;
        RECT 110.075 53.560 116.105 54.000 ;
        RECT 110.075 53.505 110.535 53.560 ;
        RECT 115.645 53.455 116.105 53.560 ;
        RECT 112.335 48.810 112.815 48.875 ;
        RECT 112.335 48.490 114.135 48.810 ;
        RECT 112.335 48.325 112.815 48.490 ;
        RECT 113.565 45.650 114.125 48.490 ;
        RECT 117.445 45.650 117.925 45.675 ;
        RECT 113.565 45.230 117.925 45.650 ;
        RECT 113.565 45.220 114.125 45.230 ;
        RECT 117.445 45.125 117.925 45.230 ;
        RECT 110.675 40.170 111.155 40.275 ;
        RECT 114.475 40.170 115.035 40.180 ;
        RECT 110.675 39.750 115.035 40.170 ;
        RECT 110.675 39.725 111.155 39.750 ;
        RECT 114.475 36.910 115.035 39.750 ;
        RECT 115.785 36.910 116.265 37.075 ;
        RECT 114.465 36.590 116.265 36.910 ;
        RECT 115.785 36.525 116.265 36.590 ;
        RECT 112.495 31.840 112.955 31.945 ;
        RECT 118.065 31.840 118.525 31.895 ;
        RECT 112.495 31.400 118.525 31.840 ;
        RECT 112.495 31.375 112.955 31.400 ;
        RECT 118.065 31.325 118.525 31.400 ;
        RECT 119.085 12.205 119.575 73.070 ;
        RECT 121.325 54.000 121.785 54.075 ;
        RECT 126.895 54.000 127.355 54.025 ;
        RECT 121.325 53.560 127.355 54.000 ;
        RECT 121.325 53.505 121.785 53.560 ;
        RECT 126.895 53.455 127.355 53.560 ;
        RECT 123.585 48.810 124.065 48.875 ;
        RECT 123.585 48.490 125.385 48.810 ;
        RECT 123.585 48.325 124.065 48.490 ;
        RECT 124.815 45.650 125.375 48.490 ;
        RECT 128.695 45.650 129.175 45.675 ;
        RECT 124.815 45.230 129.175 45.650 ;
        RECT 124.815 45.220 125.375 45.230 ;
        RECT 128.695 45.125 129.175 45.230 ;
        RECT 121.885 40.190 122.365 40.295 ;
        RECT 125.685 40.190 126.245 40.200 ;
        RECT 121.885 39.770 126.245 40.190 ;
        RECT 121.885 39.745 122.365 39.770 ;
        RECT 125.685 36.930 126.245 39.770 ;
        RECT 126.995 36.930 127.475 37.095 ;
        RECT 125.675 36.610 127.475 36.930 ;
        RECT 126.995 36.545 127.475 36.610 ;
        RECT 123.705 31.860 124.165 31.965 ;
        RECT 129.275 31.860 129.735 31.915 ;
        RECT 123.705 31.420 129.735 31.860 ;
        RECT 123.705 31.395 124.165 31.420 ;
        RECT 129.275 31.345 129.735 31.420 ;
        RECT 130.335 12.235 130.825 73.140 ;
        RECT 74.055 11.010 74.545 11.015 ;
        RECT 83.795 11.005 85.915 12.155 ;
        RECT 95.095 11.005 97.215 12.155 ;
        RECT 106.285 11.055 108.405 12.205 ;
        RECT 117.515 11.055 119.635 12.205 ;
        RECT 128.815 11.085 130.935 12.235 ;
        RECT 107.865 11.010 108.355 11.055 ;
        RECT 119.085 11.050 119.575 11.055 ;
        RECT 85.375 11.000 85.865 11.005 ;
        RECT 96.605 10.980 97.095 11.005 ;
        RECT 74.290 0.135 75.680 1.435 ;
        RECT 93.500 0.205 94.890 1.505 ;
        RECT 112.900 0.335 114.290 1.635 ;
        RECT 131.800 0.405 133.540 1.905 ;
        RECT 151.600 0.275 152.970 1.445 ;
      LAYER met4 ;
        RECT 30.420 225.130 30.670 225.140 ;
        RECT 30.300 224.760 30.670 225.130 ;
        RECT 30.970 224.760 33.430 225.140 ;
        RECT 33.730 224.760 36.190 225.140 ;
        RECT 36.490 224.760 38.950 225.140 ;
        RECT 39.250 224.760 41.710 225.140 ;
        RECT 42.010 224.760 44.470 225.140 ;
        RECT 44.770 224.760 47.230 225.140 ;
        RECT 47.530 224.760 49.990 225.140 ;
        RECT 50.290 224.760 52.750 225.140 ;
        RECT 53.050 224.760 55.510 225.140 ;
        RECT 55.810 224.760 58.270 225.140 ;
        RECT 58.570 224.760 61.030 225.140 ;
        RECT 61.330 224.760 63.790 225.140 ;
        RECT 64.090 224.760 66.550 225.140 ;
        RECT 66.850 224.760 69.310 225.140 ;
        RECT 69.610 224.760 72.070 225.140 ;
        RECT 72.370 224.760 74.830 225.140 ;
        RECT 75.130 224.760 77.590 225.140 ;
        RECT 77.890 224.760 80.350 225.140 ;
        RECT 80.650 224.760 83.110 225.140 ;
        RECT 83.410 224.760 85.870 225.140 ;
        RECT 86.170 224.760 88.630 225.140 ;
        RECT 88.930 224.760 91.390 225.140 ;
        RECT 91.690 224.760 94.150 225.140 ;
        RECT 94.450 224.760 96.910 225.140 ;
        RECT 97.210 224.760 99.670 225.140 ;
        RECT 99.970 224.760 102.430 225.140 ;
        RECT 102.730 224.760 105.190 225.140 ;
        RECT 105.490 224.760 107.950 225.140 ;
        RECT 108.250 224.760 110.710 225.140 ;
        RECT 111.010 224.760 113.470 225.140 ;
        RECT 113.770 224.760 116.230 225.140 ;
        RECT 116.530 224.760 118.990 225.140 ;
        RECT 119.290 224.760 121.750 225.140 ;
        RECT 122.050 224.760 124.510 225.140 ;
        RECT 124.810 224.760 127.270 225.140 ;
        RECT 127.570 224.760 130.030 225.140 ;
        RECT 130.330 224.760 132.790 225.140 ;
        RECT 133.090 224.760 133.520 225.140 ;
        RECT 30.300 224.240 133.520 224.760 ;
        RECT 135.385 224.760 135.550 225.185 ;
        RECT 135.850 224.760 136.745 225.185 ;
        RECT 30.300 219.100 31.660 224.240 ;
        RECT 135.385 223.875 136.745 224.760 ;
        RECT 138.175 224.760 138.310 225.115 ;
        RECT 138.610 224.760 139.535 225.115 ;
        RECT 138.175 223.805 139.535 224.760 ;
        RECT 143.225 224.760 143.830 225.145 ;
        RECT 144.130 224.760 144.585 225.145 ;
        RECT 143.225 223.835 144.585 224.760 ;
        RECT 6.000 218.040 31.660 219.100 ;
        RECT 30.300 217.960 31.660 218.040 ;
        RECT 16.820 99.530 18.820 211.530 ;
        RECT 31.820 99.530 33.820 211.530 ;
        RECT 45.315 167.945 45.645 168.275 ;
        RECT 45.330 132.235 45.630 167.945 ;
        RECT 45.315 131.905 45.645 132.235 ;
        RECT 46.820 99.530 48.820 211.530 ;
        RECT 61.820 99.530 63.820 211.530 ;
        RECT 64.635 174.065 64.965 174.395 ;
        RECT 64.650 168.955 64.950 174.065 ;
        RECT 64.635 168.625 64.965 168.955 ;
        RECT 64.650 149.235 64.950 168.625 ;
        RECT 64.635 148.905 64.965 149.235 ;
        RECT 64.650 125.435 64.950 148.905 ;
        RECT 75.675 146.185 76.005 146.515 ;
        RECT 75.690 139.035 75.990 146.185 ;
        RECT 75.675 138.705 76.005 139.035 ;
        RECT 64.635 125.105 64.965 125.435 ;
        RECT 76.820 99.530 78.820 211.530 ;
        RECT 83.955 184.265 84.285 184.595 ;
        RECT 82.115 160.465 82.445 160.795 ;
        RECT 80.275 140.745 80.605 141.075 ;
        RECT 80.290 111.835 80.590 140.745 ;
        RECT 82.130 132.235 82.430 160.465 ;
        RECT 83.970 145.835 84.270 184.265 ;
        RECT 83.955 145.505 84.285 145.835 ;
        RECT 82.115 131.905 82.445 132.235 ;
        RECT 89.475 125.785 89.805 126.115 ;
        RECT 89.490 118.635 89.790 125.785 ;
        RECT 89.475 118.305 89.805 118.635 ;
        RECT 80.275 111.505 80.605 111.835 ;
        RECT 91.820 99.530 93.820 211.530 ;
        RECT 106.820 99.530 108.820 211.530 ;
        RECT 121.820 99.720 123.820 211.530 ;
        RECT 118.110 97.700 120.130 99.670 ;
        RECT 121.810 97.750 123.830 99.720 ;
        RECT 118.130 93.980 120.130 97.700 ;
        RECT 121.820 96.830 123.820 97.750 ;
        RECT 121.820 94.830 139.410 96.830 ;
        RECT 118.130 91.980 135.580 93.980 ;
        RECT 133.580 77.835 135.580 91.980 ;
        RECT 133.375 76.625 136.015 77.835 ;
        RECT 137.410 77.815 139.410 94.830 ;
        RECT 137.235 76.605 139.875 77.815 ;
        RECT 3.955 71.365 4.000 73.195 ;
        RECT 6.000 71.365 6.055 73.195 ;
        RECT 3.000 68.705 3.025 70.435 ;
        RECT 15.555 68.655 16.995 71.165 ;
        RECT 74.335 1.000 75.635 1.415 ;
        RECT 74.335 0.155 74.530 1.000 ;
        RECT 75.430 0.155 75.635 1.000 ;
        RECT 93.545 1.000 94.845 1.485 ;
        RECT 93.545 0.225 93.850 1.000 ;
        RECT 94.750 0.225 94.845 1.000 ;
        RECT 112.945 1.000 114.245 1.615 ;
        RECT 112.945 0.355 113.170 1.000 ;
        RECT 114.070 0.355 114.245 1.000 ;
        RECT 131.845 1.000 133.495 1.885 ;
        RECT 131.845 0.425 132.490 1.000 ;
        RECT 133.390 0.425 133.495 1.000 ;
        RECT 151.645 1.000 152.925 1.425 ;
        RECT 151.645 0.295 151.810 1.000 ;
        RECT 152.710 0.295 152.925 1.000 ;
  END
END tt_um_08_sws
END LIBRARY

