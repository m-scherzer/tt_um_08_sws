VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_08_sws
  CLASS BLOCK ;
  FOREIGN tt_um_08_sws ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    ANTENNAGATEAREA 200.000000 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    ANTENNAGATEAREA 550.000000 ;
    ANTENNADIFFAREA 2.900000 ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    ANTENNAGATEAREA 550.000000 ;
    ANTENNADIFFAREA 2.900000 ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    ANTENNADIFFAREA 29.000000 ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    ANTENNADIFFAREA 29.000000 ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    ANTENNADIFFAREA 394.109192 ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 20.785 211.185 20.955 211.375 ;
        RECT 22.220 211.235 22.340 211.345 ;
        RECT 24.005 211.185 24.175 211.375 ;
        RECT 25.845 211.185 26.015 211.375 ;
        RECT 31.365 211.185 31.535 211.375 ;
        RECT 36.885 211.185 37.055 211.375 ;
        RECT 38.725 211.185 38.895 211.375 ;
        RECT 44.245 211.185 44.415 211.375 ;
        RECT 49.765 211.185 49.935 211.375 ;
        RECT 51.605 211.185 51.775 211.375 ;
        RECT 57.125 211.185 57.295 211.375 ;
        RECT 62.645 211.185 62.815 211.375 ;
        RECT 64.485 211.185 64.655 211.375 ;
        RECT 70.005 211.185 70.175 211.375 ;
        RECT 75.525 211.185 75.695 211.375 ;
        RECT 77.365 211.185 77.535 211.375 ;
        RECT 82.885 211.185 83.055 211.375 ;
        RECT 88.405 211.185 88.575 211.375 ;
        RECT 90.245 211.185 90.415 211.375 ;
        RECT 95.765 211.185 95.935 211.375 ;
        RECT 101.285 211.185 101.455 211.375 ;
        RECT 103.125 211.185 103.295 211.375 ;
        RECT 108.645 211.185 108.815 211.375 ;
        RECT 114.165 211.185 114.335 211.375 ;
        RECT 115.140 211.235 115.260 211.345 ;
        RECT 120.605 211.185 120.775 211.375 ;
        RECT 126.125 211.185 126.295 211.375 ;
        RECT 127.505 211.185 127.675 211.375 ;
        RECT 20.645 210.375 22.015 211.185 ;
        RECT 22.485 210.375 24.315 211.185 ;
        RECT 24.335 210.315 24.765 211.100 ;
        RECT 24.785 210.375 26.155 211.185 ;
        RECT 26.165 210.375 31.675 211.185 ;
        RECT 31.685 210.375 37.195 211.185 ;
        RECT 37.215 210.315 37.645 211.100 ;
        RECT 37.665 210.375 39.035 211.185 ;
        RECT 39.045 210.375 44.555 211.185 ;
        RECT 44.565 210.375 50.075 211.185 ;
        RECT 50.095 210.315 50.525 211.100 ;
        RECT 50.545 210.375 51.915 211.185 ;
        RECT 51.925 210.375 57.435 211.185 ;
        RECT 57.445 210.375 62.955 211.185 ;
        RECT 62.975 210.315 63.405 211.100 ;
        RECT 63.425 210.375 64.795 211.185 ;
        RECT 64.805 210.375 70.315 211.185 ;
        RECT 70.325 210.375 75.835 211.185 ;
        RECT 75.855 210.315 76.285 211.100 ;
        RECT 76.305 210.375 77.675 211.185 ;
        RECT 77.685 210.375 83.195 211.185 ;
        RECT 83.205 210.375 88.715 211.185 ;
        RECT 88.735 210.315 89.165 211.100 ;
        RECT 89.185 210.375 90.555 211.185 ;
        RECT 90.565 210.375 96.075 211.185 ;
        RECT 96.085 210.375 101.595 211.185 ;
        RECT 101.615 210.315 102.045 211.100 ;
        RECT 102.065 210.375 103.435 211.185 ;
        RECT 103.445 210.375 108.955 211.185 ;
        RECT 108.965 210.375 114.475 211.185 ;
        RECT 114.495 210.315 114.925 211.100 ;
        RECT 115.405 210.375 120.915 211.185 ;
        RECT 120.925 210.375 126.435 211.185 ;
        RECT 126.445 210.375 127.815 211.185 ;
      LAYER nwell ;
        RECT 20.450 207.155 128.010 209.985 ;
      LAYER pwell ;
        RECT 20.645 205.955 22.015 206.765 ;
        RECT 22.485 205.955 24.315 206.765 ;
        RECT 24.335 206.040 24.765 206.825 ;
        RECT 25.245 205.955 27.995 206.765 ;
        RECT 28.005 205.955 33.515 206.765 ;
        RECT 33.525 205.955 39.035 206.765 ;
        RECT 39.045 205.955 44.555 206.765 ;
        RECT 44.565 205.955 50.075 206.765 ;
        RECT 50.095 206.040 50.525 206.825 ;
        RECT 51.005 205.955 53.755 206.765 ;
        RECT 53.765 205.955 59.275 206.765 ;
        RECT 59.285 205.955 64.795 206.765 ;
        RECT 64.805 205.955 70.315 206.765 ;
        RECT 70.325 205.955 75.835 206.765 ;
        RECT 75.855 206.040 76.285 206.825 ;
        RECT 76.765 205.955 79.515 206.765 ;
        RECT 79.525 205.955 85.035 206.765 ;
        RECT 85.045 205.955 90.555 206.765 ;
        RECT 90.565 205.955 96.075 206.765 ;
        RECT 96.085 205.955 101.595 206.765 ;
        RECT 101.615 206.040 102.045 206.825 ;
        RECT 102.525 205.955 104.355 206.765 ;
        RECT 104.365 205.955 109.875 206.765 ;
        RECT 109.885 205.955 115.395 206.765 ;
        RECT 115.405 205.955 120.915 206.765 ;
        RECT 120.925 205.955 126.435 206.765 ;
        RECT 126.445 205.955 127.815 206.765 ;
        RECT 20.785 205.745 20.955 205.955 ;
        RECT 22.220 205.795 22.340 205.905 ;
        RECT 24.005 205.765 24.175 205.955 ;
        RECT 24.980 205.795 25.100 205.905 ;
        RECT 25.845 205.745 26.015 205.935 ;
        RECT 27.685 205.765 27.855 205.955 ;
        RECT 31.365 205.745 31.535 205.935 ;
        RECT 33.205 205.765 33.375 205.955 ;
        RECT 36.885 205.745 37.055 205.935 ;
        RECT 37.860 205.795 37.980 205.905 ;
        RECT 38.725 205.765 38.895 205.955 ;
        RECT 40.565 205.745 40.735 205.935 ;
        RECT 44.245 205.765 44.415 205.955 ;
        RECT 46.085 205.745 46.255 205.935 ;
        RECT 49.765 205.765 49.935 205.955 ;
        RECT 50.740 205.795 50.860 205.905 ;
        RECT 51.605 205.745 51.775 205.935 ;
        RECT 53.445 205.765 53.615 205.955 ;
        RECT 57.125 205.745 57.295 205.935 ;
        RECT 58.965 205.765 59.135 205.955 ;
        RECT 62.645 205.745 62.815 205.935 ;
        RECT 63.620 205.795 63.740 205.905 ;
        RECT 64.485 205.765 64.655 205.955 ;
        RECT 66.325 205.745 66.495 205.935 ;
        RECT 70.005 205.765 70.175 205.955 ;
        RECT 71.845 205.745 72.015 205.935 ;
        RECT 75.525 205.765 75.695 205.955 ;
        RECT 76.500 205.795 76.620 205.905 ;
        RECT 77.365 205.745 77.535 205.935 ;
        RECT 79.205 205.765 79.375 205.955 ;
        RECT 82.885 205.745 83.055 205.935 ;
        RECT 84.725 205.765 84.895 205.955 ;
        RECT 88.405 205.745 88.575 205.935 ;
        RECT 89.380 205.795 89.500 205.905 ;
        RECT 90.245 205.765 90.415 205.955 ;
        RECT 92.085 205.745 92.255 205.935 ;
        RECT 95.765 205.765 95.935 205.955 ;
        RECT 97.605 205.745 97.775 205.935 ;
        RECT 101.285 205.765 101.455 205.955 ;
        RECT 102.260 205.795 102.380 205.905 ;
        RECT 103.125 205.745 103.295 205.935 ;
        RECT 104.045 205.765 104.215 205.955 ;
        RECT 108.645 205.745 108.815 205.935 ;
        RECT 109.565 205.765 109.735 205.955 ;
        RECT 114.165 205.745 114.335 205.935 ;
        RECT 115.085 205.905 115.255 205.955 ;
        RECT 115.085 205.795 115.260 205.905 ;
        RECT 115.085 205.765 115.255 205.795 ;
        RECT 120.605 205.745 120.775 205.955 ;
        RECT 126.125 205.745 126.295 205.955 ;
        RECT 127.505 205.745 127.675 205.955 ;
        RECT 20.645 204.935 22.015 205.745 ;
        RECT 22.485 204.935 26.155 205.745 ;
        RECT 26.165 204.935 31.675 205.745 ;
        RECT 31.685 204.935 37.195 205.745 ;
        RECT 37.215 204.875 37.645 205.660 ;
        RECT 38.125 204.935 40.875 205.745 ;
        RECT 40.885 204.935 46.395 205.745 ;
        RECT 46.405 204.935 51.915 205.745 ;
        RECT 51.925 204.935 57.435 205.745 ;
        RECT 57.445 204.935 62.955 205.745 ;
        RECT 62.975 204.875 63.405 205.660 ;
        RECT 63.885 204.935 66.635 205.745 ;
        RECT 66.645 204.935 72.155 205.745 ;
        RECT 72.165 204.935 77.675 205.745 ;
        RECT 77.685 204.935 83.195 205.745 ;
        RECT 83.205 204.935 88.715 205.745 ;
        RECT 88.735 204.875 89.165 205.660 ;
        RECT 89.645 204.935 92.395 205.745 ;
        RECT 92.405 204.935 97.915 205.745 ;
        RECT 97.925 204.935 103.435 205.745 ;
        RECT 103.445 204.935 108.955 205.745 ;
        RECT 108.965 204.935 114.475 205.745 ;
        RECT 114.495 204.875 114.925 205.660 ;
        RECT 115.405 204.935 120.915 205.745 ;
        RECT 120.925 204.935 126.435 205.745 ;
        RECT 126.445 204.935 127.815 205.745 ;
      LAYER nwell ;
        RECT 20.450 201.715 128.010 204.545 ;
      LAYER pwell ;
        RECT 20.645 200.515 22.015 201.325 ;
        RECT 22.485 200.515 24.315 201.325 ;
        RECT 24.335 200.600 24.765 201.385 ;
        RECT 25.245 200.515 27.995 201.325 ;
        RECT 28.005 200.515 33.515 201.325 ;
        RECT 33.525 200.515 39.035 201.325 ;
        RECT 39.045 200.515 44.555 201.325 ;
        RECT 44.565 200.515 50.075 201.325 ;
        RECT 50.095 200.600 50.525 201.385 ;
        RECT 51.005 200.515 53.755 201.325 ;
        RECT 53.765 200.515 59.275 201.325 ;
        RECT 59.285 200.515 64.795 201.325 ;
        RECT 64.805 200.515 70.315 201.325 ;
        RECT 70.325 200.515 73.435 201.425 ;
        RECT 74.005 200.515 75.835 201.325 ;
        RECT 75.855 200.600 76.285 201.385 ;
        RECT 76.765 200.515 79.515 201.325 ;
        RECT 79.525 200.515 85.035 201.325 ;
        RECT 85.045 200.515 90.555 201.325 ;
        RECT 90.565 200.515 96.075 201.325 ;
        RECT 96.085 200.515 101.595 201.325 ;
        RECT 101.615 200.600 102.045 201.385 ;
        RECT 102.525 200.515 104.355 201.325 ;
        RECT 104.365 200.515 109.875 201.325 ;
        RECT 109.885 200.515 115.395 201.325 ;
        RECT 115.405 200.515 120.915 201.325 ;
        RECT 120.925 200.515 126.435 201.325 ;
        RECT 126.445 200.515 127.815 201.325 ;
        RECT 20.785 200.305 20.955 200.515 ;
        RECT 22.220 200.355 22.340 200.465 ;
        RECT 24.005 200.325 24.175 200.515 ;
        RECT 24.980 200.355 25.100 200.465 ;
        RECT 25.845 200.305 26.015 200.495 ;
        RECT 27.685 200.325 27.855 200.515 ;
        RECT 31.365 200.305 31.535 200.495 ;
        RECT 33.205 200.325 33.375 200.515 ;
        RECT 36.885 200.305 37.055 200.495 ;
        RECT 38.725 200.325 38.895 200.515 ;
        RECT 40.105 200.305 40.275 200.495 ;
        RECT 44.245 200.325 44.415 200.515 ;
        RECT 45.625 200.305 45.795 200.495 ;
        RECT 46.085 200.305 46.255 200.495 ;
        RECT 49.765 200.325 49.935 200.515 ;
        RECT 50.740 200.355 50.860 200.465 ;
        RECT 53.445 200.325 53.615 200.515 ;
        RECT 55.745 200.350 55.905 200.460 ;
        RECT 58.965 200.325 59.135 200.515 ;
        RECT 61.265 200.305 61.435 200.495 ;
        RECT 62.645 200.305 62.815 200.495 ;
        RECT 63.565 200.305 63.735 200.495 ;
        RECT 64.485 200.325 64.655 200.515 ;
        RECT 70.005 200.325 70.175 200.515 ;
        RECT 73.225 200.325 73.395 200.515 ;
        RECT 73.740 200.355 73.860 200.465 ;
        RECT 75.525 200.325 75.695 200.515 ;
        RECT 20.645 199.495 22.015 200.305 ;
        RECT 22.485 199.495 26.155 200.305 ;
        RECT 26.165 199.495 31.675 200.305 ;
        RECT 31.685 199.495 37.195 200.305 ;
        RECT 37.215 199.435 37.645 200.220 ;
        RECT 37.665 199.495 40.415 200.305 ;
        RECT 40.425 199.495 45.935 200.305 ;
        RECT 45.945 199.625 55.135 200.305 ;
        RECT 50.455 199.405 51.385 199.625 ;
        RECT 54.215 199.395 55.135 199.625 ;
        RECT 56.065 199.495 61.575 200.305 ;
        RECT 61.595 199.395 62.945 200.305 ;
        RECT 62.975 199.435 63.405 200.220 ;
        RECT 63.425 199.625 73.035 200.305 ;
        RECT 67.935 199.405 68.865 199.625 ;
        RECT 71.695 199.395 73.035 199.625 ;
        RECT 73.085 200.275 74.030 200.305 ;
        RECT 75.985 200.275 76.155 200.495 ;
        RECT 76.500 200.355 76.620 200.465 ;
        RECT 78.285 200.305 78.455 200.495 ;
        RECT 78.745 200.305 78.915 200.495 ;
        RECT 79.205 200.325 79.375 200.515 ;
        RECT 80.125 200.305 80.295 200.495 ;
        RECT 84.725 200.325 84.895 200.515 ;
        RECT 88.405 200.305 88.575 200.495 ;
        RECT 90.245 200.325 90.415 200.515 ;
        RECT 92.545 200.305 92.715 200.495 ;
        RECT 95.765 200.325 95.935 200.515 ;
        RECT 98.065 200.305 98.235 200.495 ;
        RECT 101.285 200.325 101.455 200.515 ;
        RECT 102.260 200.355 102.380 200.465 ;
        RECT 104.045 200.325 104.215 200.515 ;
        RECT 107.265 200.305 107.435 200.495 ;
        RECT 109.565 200.325 109.735 200.515 ;
        RECT 110.025 200.305 110.195 200.495 ;
        RECT 113.890 200.305 114.060 200.495 ;
        RECT 115.085 200.325 115.255 200.515 ;
        RECT 120.605 200.325 120.775 200.515 ;
        RECT 123.825 200.305 123.995 200.495 ;
        RECT 124.340 200.355 124.460 200.465 ;
        RECT 126.125 200.305 126.295 200.515 ;
        RECT 127.505 200.305 127.675 200.515 ;
        RECT 73.085 200.075 76.155 200.275 ;
        RECT 73.085 199.595 76.295 200.075 ;
        RECT 73.085 199.395 74.030 199.595 ;
        RECT 75.365 199.395 76.295 199.595 ;
        RECT 76.765 199.495 78.595 200.305 ;
        RECT 78.615 199.395 79.965 200.305 ;
        RECT 80.085 199.395 83.195 200.305 ;
        RECT 83.205 199.495 88.715 200.305 ;
        RECT 88.735 199.435 89.165 200.220 ;
        RECT 89.185 199.495 92.855 200.305 ;
        RECT 92.865 199.495 98.375 200.305 ;
        RECT 98.385 199.625 107.575 200.305 ;
        RECT 98.385 199.395 99.305 199.625 ;
        RECT 102.135 199.405 103.065 199.625 ;
        RECT 107.585 199.495 110.335 200.305 ;
        RECT 110.575 199.625 114.475 200.305 ;
        RECT 113.545 199.395 114.475 199.625 ;
        RECT 114.495 199.435 114.925 200.220 ;
        RECT 114.945 199.625 124.135 200.305 ;
        RECT 114.945 199.395 115.865 199.625 ;
        RECT 118.695 199.405 119.625 199.625 ;
        RECT 124.605 199.495 126.435 200.305 ;
        RECT 126.445 199.495 127.815 200.305 ;
      LAYER nwell ;
        RECT 20.450 196.275 128.010 199.105 ;
      LAYER pwell ;
        RECT 20.645 195.075 22.015 195.885 ;
        RECT 22.485 195.075 24.315 195.885 ;
        RECT 24.335 195.160 24.765 195.945 ;
        RECT 25.245 195.075 27.995 195.885 ;
        RECT 28.005 195.075 33.515 195.885 ;
        RECT 33.535 195.075 34.885 195.985 ;
        RECT 34.905 195.075 36.735 195.885 ;
        RECT 36.745 195.075 42.255 195.885 ;
        RECT 42.275 195.075 43.625 195.985 ;
        RECT 43.645 195.075 45.475 195.885 ;
        RECT 48.685 195.755 49.615 195.985 ;
        RECT 45.715 195.075 49.615 195.755 ;
        RECT 50.095 195.160 50.525 195.945 ;
        RECT 51.465 195.075 55.135 195.885 ;
        RECT 58.345 195.755 59.275 195.985 ;
        RECT 55.375 195.075 59.275 195.755 ;
        RECT 59.745 195.075 61.115 195.855 ;
        RECT 61.125 195.075 66.635 195.885 ;
        RECT 66.655 195.075 68.005 195.985 ;
        RECT 70.315 195.755 71.235 195.985 ;
        RECT 68.945 195.075 71.235 195.755 ;
        RECT 71.245 195.075 74.165 195.985 ;
        RECT 74.465 195.075 75.835 195.885 ;
        RECT 75.855 195.160 76.285 195.945 ;
        RECT 77.225 195.755 78.145 195.985 ;
        RECT 80.975 195.755 81.905 195.975 ;
        RECT 88.245 195.755 89.165 195.975 ;
        RECT 95.245 195.875 96.165 195.985 ;
        RECT 93.830 195.755 96.165 195.875 ;
        RECT 77.225 195.075 86.415 195.755 ;
        RECT 86.885 195.075 96.165 195.755 ;
        RECT 96.545 195.075 100.215 195.885 ;
        RECT 100.235 195.075 101.585 195.985 ;
        RECT 101.615 195.160 102.045 195.945 ;
        RECT 102.985 195.075 104.355 195.855 ;
        RECT 104.365 195.075 108.035 195.885 ;
        RECT 108.055 195.075 109.405 195.985 ;
        RECT 109.425 195.755 110.345 195.985 ;
        RECT 113.175 195.755 114.105 195.975 ;
        RECT 109.425 195.075 118.615 195.755 ;
        RECT 118.625 195.075 119.995 195.855 ;
        RECT 120.925 195.075 126.435 195.885 ;
        RECT 126.445 195.075 127.815 195.885 ;
        RECT 20.785 194.865 20.955 195.075 ;
        RECT 22.220 194.915 22.340 195.025 ;
        RECT 24.005 194.885 24.175 195.075 ;
        RECT 24.980 194.915 25.100 195.025 ;
        RECT 27.685 194.865 27.855 195.075 ;
        RECT 28.145 194.865 28.315 195.055 ;
        RECT 33.205 194.885 33.375 195.075 ;
        RECT 34.585 194.885 34.755 195.075 ;
        RECT 36.425 194.885 36.595 195.075 ;
        RECT 38.725 194.865 38.895 195.055 ;
        RECT 41.945 194.885 42.115 195.075 ;
        RECT 42.405 194.885 42.575 195.075 ;
        RECT 45.165 194.885 45.335 195.075 ;
        RECT 48.385 194.865 48.555 195.055 ;
        RECT 49.030 194.885 49.200 195.075 ;
        RECT 49.765 195.025 49.935 195.055 ;
        RECT 49.765 194.915 49.940 195.025 ;
        RECT 49.765 194.865 49.935 194.915 ;
        RECT 51.145 194.865 51.315 195.055 ;
        RECT 52.525 194.865 52.695 195.055 ;
        RECT 53.445 194.910 53.605 195.020 ;
        RECT 54.825 194.885 54.995 195.075 ;
        RECT 58.690 194.885 58.860 195.075 ;
        RECT 59.480 194.915 59.600 195.025 ;
        RECT 59.885 194.885 60.055 195.075 ;
        RECT 62.645 194.865 62.815 195.055 ;
        RECT 66.325 194.885 66.495 195.075 ;
        RECT 66.785 194.885 66.955 195.075 ;
        RECT 68.625 194.920 68.785 195.030 ;
        RECT 69.085 194.885 69.255 195.075 ;
        RECT 71.390 194.885 71.560 195.075 ;
        RECT 73.685 194.865 73.855 195.055 ;
        RECT 75.525 194.885 75.695 195.075 ;
        RECT 20.645 194.055 22.015 194.865 ;
        RECT 22.485 194.055 27.995 194.865 ;
        RECT 28.005 194.185 37.195 194.865 ;
        RECT 32.515 193.965 33.445 194.185 ;
        RECT 36.275 193.955 37.195 194.185 ;
        RECT 37.215 193.995 37.645 194.780 ;
        RECT 37.665 194.055 39.035 194.865 ;
        RECT 39.415 194.185 48.695 194.865 ;
        RECT 39.415 194.065 41.750 194.185 ;
        RECT 39.415 193.955 40.335 194.065 ;
        RECT 46.415 193.965 47.335 194.185 ;
        RECT 48.705 194.085 50.075 194.865 ;
        RECT 50.085 194.085 51.455 194.865 ;
        RECT 51.475 193.955 52.825 194.865 ;
        RECT 53.765 194.185 62.955 194.865 ;
        RECT 53.765 193.955 54.685 194.185 ;
        RECT 57.515 193.965 58.445 194.185 ;
        RECT 62.975 193.995 63.405 194.780 ;
        RECT 63.625 194.185 73.995 194.865 ;
        RECT 74.005 194.835 74.950 194.865 ;
        RECT 76.905 194.835 77.075 195.055 ;
        RECT 79.205 194.885 79.375 195.055 ;
        RECT 79.205 194.865 79.370 194.885 ;
        RECT 79.665 194.865 79.835 195.055 ;
        RECT 82.430 194.865 82.600 195.055 ;
        RECT 84.265 194.865 84.435 195.055 ;
        RECT 84.725 194.865 84.895 195.055 ;
        RECT 86.105 194.885 86.275 195.075 ;
        RECT 86.620 194.915 86.740 195.025 ;
        RECT 87.025 194.865 87.195 195.075 ;
        RECT 87.485 194.865 87.655 195.055 ;
        RECT 98.525 194.865 98.695 195.055 ;
        RECT 99.905 194.885 100.075 195.075 ;
        RECT 100.365 194.885 100.535 195.075 ;
        RECT 102.390 194.865 102.560 195.055 ;
        RECT 102.665 194.920 102.825 195.030 ;
        RECT 103.125 194.885 103.295 195.075 ;
        RECT 104.505 194.865 104.675 195.055 ;
        RECT 107.725 194.885 107.895 195.075 ;
        RECT 108.185 194.885 108.355 195.075 ;
        RECT 110.025 194.865 110.195 195.055 ;
        RECT 113.890 194.865 114.060 195.055 ;
        RECT 115.545 194.910 115.705 195.020 ;
        RECT 116.005 194.865 116.175 195.055 ;
        RECT 118.305 194.885 118.475 195.075 ;
        RECT 118.765 194.865 118.935 195.055 ;
        RECT 119.225 194.865 119.395 195.055 ;
        RECT 119.685 194.885 119.855 195.075 ;
        RECT 120.605 195.025 120.765 195.030 ;
        RECT 120.605 194.920 120.780 195.025 ;
        RECT 120.660 194.915 120.780 194.920 ;
        RECT 126.125 194.865 126.295 195.075 ;
        RECT 127.505 194.865 127.675 195.075 ;
        RECT 74.005 194.635 77.075 194.835 ;
        RECT 63.625 193.955 65.835 194.185 ;
        RECT 68.555 193.965 69.485 194.185 ;
        RECT 74.005 194.155 77.215 194.635 ;
        RECT 74.005 193.955 74.950 194.155 ;
        RECT 76.285 193.955 77.215 194.155 ;
        RECT 77.535 194.185 79.370 194.865 ;
        RECT 79.525 194.185 81.355 194.865 ;
        RECT 77.535 193.955 78.465 194.185 ;
        RECT 80.010 193.955 81.355 194.185 ;
        RECT 81.365 193.955 82.715 194.865 ;
        RECT 82.745 194.055 84.575 194.865 ;
        RECT 84.585 194.085 85.955 194.865 ;
        RECT 85.975 193.955 87.325 194.865 ;
        RECT 87.355 193.955 88.705 194.865 ;
        RECT 88.735 193.995 89.165 194.780 ;
        RECT 89.555 194.185 98.835 194.865 ;
        RECT 99.075 194.185 102.975 194.865 ;
        RECT 89.555 194.065 91.890 194.185 ;
        RECT 89.555 193.955 90.475 194.065 ;
        RECT 96.555 193.965 97.475 194.185 ;
        RECT 102.045 193.955 102.975 194.185 ;
        RECT 102.985 194.055 104.815 194.865 ;
        RECT 104.825 194.055 110.335 194.865 ;
        RECT 110.575 194.185 114.475 194.865 ;
        RECT 113.545 193.955 114.475 194.185 ;
        RECT 114.495 193.995 114.925 194.780 ;
        RECT 115.875 193.955 117.225 194.865 ;
        RECT 117.245 194.055 119.075 194.865 ;
        RECT 119.085 194.085 120.455 194.865 ;
        RECT 120.925 194.055 126.435 194.865 ;
        RECT 126.445 194.055 127.815 194.865 ;
      LAYER nwell ;
        RECT 20.450 190.835 128.010 193.665 ;
      LAYER pwell ;
        RECT 20.645 189.635 22.015 190.445 ;
        RECT 22.485 189.635 24.315 190.445 ;
        RECT 24.335 189.720 24.765 190.505 ;
        RECT 24.785 189.635 26.155 190.445 ;
        RECT 26.165 189.635 31.675 190.445 ;
        RECT 31.695 189.635 33.045 190.545 ;
        RECT 33.985 189.635 35.355 190.415 ;
        RECT 35.365 190.315 36.295 190.545 ;
        RECT 35.365 189.635 39.265 190.315 ;
        RECT 39.505 189.635 42.255 190.445 ;
        RECT 45.465 190.315 46.395 190.545 ;
        RECT 42.495 189.635 46.395 190.315 ;
        RECT 46.405 189.635 50.075 190.445 ;
        RECT 50.095 189.720 50.525 190.505 ;
        RECT 51.005 189.635 52.835 190.445 ;
        RECT 52.855 189.635 54.205 190.545 ;
        RECT 54.225 189.635 55.595 190.445 ;
        RECT 55.605 189.635 56.975 190.415 ;
        RECT 56.995 189.635 58.345 190.545 ;
        RECT 58.365 189.635 59.735 190.445 ;
        RECT 59.745 189.635 65.255 190.445 ;
        RECT 65.265 189.635 70.775 190.445 ;
        RECT 70.785 189.635 72.155 190.415 ;
        RECT 72.165 189.635 73.535 190.445 ;
        RECT 73.545 189.635 75.835 190.545 ;
        RECT 75.855 189.720 76.285 190.505 ;
        RECT 78.135 190.315 79.055 190.545 ;
        RECT 76.765 189.635 79.055 190.315 ;
        RECT 79.065 189.635 80.435 190.415 ;
        RECT 80.905 189.635 83.655 190.445 ;
        RECT 83.665 189.635 89.175 190.445 ;
        RECT 89.185 190.315 90.115 190.545 ;
        RECT 89.185 189.635 93.085 190.315 ;
        RECT 93.325 189.635 94.695 190.415 ;
        RECT 94.705 189.635 96.075 190.445 ;
        RECT 96.085 189.635 101.595 190.445 ;
        RECT 101.615 189.720 102.045 190.505 ;
        RECT 102.985 189.635 108.495 190.445 ;
        RECT 108.505 190.315 109.425 190.545 ;
        RECT 112.255 190.315 113.185 190.535 ;
        RECT 108.505 189.635 117.695 190.315 ;
        RECT 117.705 189.635 120.455 190.445 ;
        RECT 120.465 189.635 121.835 190.415 ;
        RECT 122.765 189.635 126.435 190.445 ;
        RECT 126.445 189.635 127.815 190.445 ;
        RECT 20.785 189.425 20.955 189.635 ;
        RECT 22.220 189.475 22.340 189.585 ;
        RECT 24.005 189.445 24.175 189.635 ;
        RECT 25.845 189.445 26.015 189.635 ;
        RECT 27.685 189.425 27.855 189.615 ;
        RECT 28.145 189.425 28.315 189.615 ;
        RECT 31.365 189.445 31.535 189.635 ;
        RECT 31.825 189.445 31.995 189.635 ;
        RECT 33.665 189.480 33.825 189.590 ;
        RECT 35.045 189.445 35.215 189.635 ;
        RECT 35.780 189.445 35.950 189.635 ;
        RECT 37.860 189.475 37.980 189.585 ;
        RECT 41.945 189.445 42.115 189.635 ;
        RECT 43.325 189.425 43.495 189.615 ;
        RECT 45.810 189.445 45.980 189.635 ;
        RECT 48.845 189.425 49.015 189.615 ;
        RECT 49.765 189.445 49.935 189.635 ;
        RECT 50.740 189.475 50.860 189.585 ;
        RECT 52.525 189.445 52.695 189.635 ;
        RECT 53.905 189.445 54.075 189.635 ;
        RECT 55.285 189.445 55.455 189.635 ;
        RECT 55.745 189.445 55.915 189.635 ;
        RECT 58.045 189.425 58.215 189.635 ;
        RECT 59.425 189.425 59.595 189.635 ;
        RECT 59.940 189.475 60.060 189.585 ;
        RECT 62.645 189.425 62.815 189.615 ;
        RECT 63.620 189.475 63.740 189.585 ;
        RECT 64.945 189.445 65.115 189.635 ;
        RECT 66.325 189.425 66.495 189.615 ;
        RECT 70.465 189.445 70.635 189.635 ;
        RECT 70.925 189.445 71.095 189.635 ;
        RECT 71.845 189.425 72.015 189.615 ;
        RECT 72.305 189.425 72.475 189.615 ;
        RECT 73.225 189.445 73.395 189.635 ;
        RECT 75.520 189.445 75.690 189.635 ;
        RECT 76.500 189.475 76.620 189.585 ;
        RECT 76.905 189.445 77.075 189.635 ;
        RECT 79.205 189.445 79.375 189.635 ;
        RECT 80.640 189.475 80.760 189.585 ;
        RECT 82.425 189.425 82.595 189.615 ;
        RECT 83.345 189.445 83.515 189.635 ;
        RECT 84.265 189.425 84.435 189.615 ;
        RECT 88.130 189.425 88.300 189.615 ;
        RECT 88.865 189.445 89.035 189.635 ;
        RECT 89.600 189.445 89.770 189.635 ;
        RECT 90.245 189.425 90.415 189.615 ;
        RECT 91.625 189.425 91.795 189.615 ;
        RECT 92.545 189.470 92.705 189.580 ;
        RECT 93.465 189.445 93.635 189.635 ;
        RECT 95.765 189.445 95.935 189.635 ;
        RECT 98.065 189.425 98.235 189.615 ;
        RECT 98.525 189.425 98.695 189.615 ;
        RECT 101.285 189.445 101.455 189.635 ;
        RECT 102.665 189.480 102.825 189.590 ;
        RECT 108.185 189.445 108.355 189.635 ;
        RECT 108.645 189.425 108.815 189.615 ;
        RECT 110.025 189.425 110.195 189.615 ;
        RECT 110.945 189.470 111.105 189.580 ;
        RECT 112.325 189.425 112.495 189.615 ;
        RECT 112.840 189.475 112.960 189.585 ;
        RECT 113.245 189.425 113.415 189.615 ;
        RECT 115.545 189.470 115.705 189.580 ;
        RECT 117.385 189.445 117.555 189.635 ;
        RECT 120.145 189.445 120.315 189.635 ;
        RECT 120.605 189.445 120.775 189.635 ;
        RECT 122.445 189.480 122.605 189.590 ;
        RECT 124.745 189.425 124.915 189.615 ;
        RECT 126.125 189.425 126.295 189.635 ;
        RECT 127.505 189.425 127.675 189.635 ;
        RECT 20.645 188.615 22.015 189.425 ;
        RECT 22.485 188.615 27.995 189.425 ;
        RECT 28.005 188.745 37.195 189.425 ;
        RECT 32.515 188.525 33.445 188.745 ;
        RECT 36.275 188.515 37.195 188.745 ;
        RECT 37.215 188.555 37.645 189.340 ;
        RECT 38.125 188.615 43.635 189.425 ;
        RECT 43.645 188.615 49.155 189.425 ;
        RECT 49.165 188.745 58.355 189.425 ;
        RECT 49.165 188.515 50.085 188.745 ;
        RECT 52.915 188.525 53.845 188.745 ;
        RECT 58.375 188.515 59.725 189.425 ;
        RECT 60.205 188.615 62.955 189.425 ;
        RECT 62.975 188.555 63.405 189.340 ;
        RECT 63.885 188.615 66.635 189.425 ;
        RECT 66.645 188.615 72.155 189.425 ;
        RECT 72.175 188.515 73.525 189.425 ;
        RECT 73.545 188.745 82.735 189.425 ;
        RECT 73.545 188.515 74.465 188.745 ;
        RECT 77.295 188.525 78.225 188.745 ;
        RECT 82.745 188.615 84.575 189.425 ;
        RECT 84.815 188.745 88.715 189.425 ;
        RECT 87.785 188.515 88.715 188.745 ;
        RECT 88.735 188.555 89.165 189.340 ;
        RECT 89.185 188.615 90.555 189.425 ;
        RECT 90.575 188.515 91.925 189.425 ;
        RECT 92.865 188.615 98.375 189.425 ;
        RECT 98.395 188.515 99.745 189.425 ;
        RECT 99.765 188.745 108.955 189.425 ;
        RECT 99.765 188.515 100.685 188.745 ;
        RECT 103.515 188.525 104.445 188.745 ;
        RECT 108.965 188.645 110.335 189.425 ;
        RECT 111.275 188.515 112.625 189.425 ;
        RECT 113.115 188.515 114.465 189.425 ;
        RECT 114.495 188.555 114.925 189.340 ;
        RECT 115.865 188.745 125.055 189.425 ;
        RECT 115.865 188.515 116.785 188.745 ;
        RECT 119.615 188.525 120.545 188.745 ;
        RECT 125.065 188.615 126.435 189.425 ;
        RECT 126.445 188.615 127.815 189.425 ;
      LAYER nwell ;
        RECT 20.450 185.395 128.010 188.225 ;
      LAYER pwell ;
        RECT 20.645 184.195 22.015 185.005 ;
        RECT 22.485 184.195 24.315 185.005 ;
        RECT 24.335 184.280 24.765 185.065 ;
        RECT 25.705 184.195 31.215 185.005 ;
        RECT 31.235 184.195 32.585 185.105 ;
        RECT 33.065 184.195 34.435 184.975 ;
        RECT 34.445 184.875 35.375 185.105 ;
        RECT 34.445 184.195 38.345 184.875 ;
        RECT 38.585 184.195 39.955 185.005 ;
        RECT 39.965 184.195 43.635 185.005 ;
        RECT 43.655 184.195 45.005 185.105 ;
        RECT 49.145 184.875 50.075 185.105 ;
        RECT 46.175 184.195 50.075 184.875 ;
        RECT 50.095 184.280 50.525 185.065 ;
        RECT 54.205 184.875 55.135 185.105 ;
        RECT 51.235 184.195 55.135 184.875 ;
        RECT 55.145 184.875 56.065 185.105 ;
        RECT 58.895 184.875 59.825 185.095 ;
        RECT 55.145 184.195 64.335 184.875 ;
        RECT 64.805 184.195 68.475 185.005 ;
        RECT 70.325 184.875 71.670 185.105 ;
        RECT 72.165 184.875 73.095 185.105 ;
        RECT 68.485 184.195 70.315 184.875 ;
        RECT 70.325 184.195 72.155 184.875 ;
        RECT 72.165 184.195 75.835 184.875 ;
        RECT 75.855 184.280 76.285 185.065 ;
        RECT 76.305 184.875 77.225 185.105 ;
        RECT 80.055 184.875 80.985 185.095 ;
        RECT 76.305 184.195 85.495 184.875 ;
        RECT 85.505 184.195 87.335 185.005 ;
        RECT 87.345 184.875 88.265 185.105 ;
        RECT 91.095 184.875 92.025 185.095 ;
        RECT 100.205 184.875 101.135 185.105 ;
        RECT 87.345 184.195 96.535 184.875 ;
        RECT 97.235 184.195 101.135 184.875 ;
        RECT 101.615 184.280 102.045 185.065 ;
        RECT 102.065 184.195 103.895 185.005 ;
        RECT 107.105 184.875 108.035 185.105 ;
        RECT 104.135 184.195 108.035 184.875 ;
        RECT 108.505 184.195 111.255 185.005 ;
        RECT 114.465 184.875 115.395 185.105 ;
        RECT 118.605 184.875 119.535 185.105 ;
        RECT 111.495 184.195 115.395 184.875 ;
        RECT 115.635 184.195 119.535 184.875 ;
        RECT 119.545 184.195 120.915 185.005 ;
        RECT 120.925 184.195 126.435 185.005 ;
        RECT 126.445 184.195 127.815 185.005 ;
        RECT 20.785 183.985 20.955 184.195 ;
        RECT 22.220 184.035 22.340 184.145 ;
        RECT 24.005 184.005 24.175 184.195 ;
        RECT 25.385 184.040 25.545 184.150 ;
        RECT 27.685 183.985 27.855 184.175 ;
        RECT 28.145 183.985 28.315 184.175 ;
        RECT 30.905 184.005 31.075 184.195 ;
        RECT 31.365 184.005 31.535 184.195 ;
        RECT 32.800 184.035 32.920 184.145 ;
        RECT 34.125 184.005 34.295 184.195 ;
        RECT 34.860 184.005 35.030 184.195 ;
        RECT 39.645 184.005 39.815 184.195 ;
        RECT 40.105 183.985 40.275 184.175 ;
        RECT 43.325 184.005 43.495 184.195 ;
        RECT 44.705 184.005 44.875 184.195 ;
        RECT 45.625 184.040 45.785 184.150 ;
        RECT 49.305 183.985 49.475 184.175 ;
        RECT 49.490 184.005 49.660 184.195 ;
        RECT 50.685 184.145 50.855 184.175 ;
        RECT 50.685 184.035 50.860 184.145 ;
        RECT 51.200 184.035 51.320 184.145 ;
        RECT 50.685 183.985 50.855 184.035 ;
        RECT 54.550 184.005 54.720 184.195 ;
        RECT 54.825 183.985 54.995 184.175 ;
        RECT 60.345 183.985 60.515 184.175 ;
        RECT 60.805 183.985 60.975 184.175 ;
        RECT 62.645 184.030 62.805 184.140 ;
        RECT 64.025 184.005 64.195 184.195 ;
        RECT 64.540 184.035 64.660 184.145 ;
        RECT 65.865 183.985 66.035 184.175 ;
        RECT 68.165 184.005 68.335 184.195 ;
        RECT 68.625 184.005 68.795 184.195 ;
        RECT 71.385 183.985 71.555 184.175 ;
        RECT 71.845 184.005 72.015 184.195 ;
        RECT 75.525 184.005 75.695 184.195 ;
        RECT 75.985 183.985 76.155 184.175 ;
        RECT 76.500 184.035 76.620 184.145 ;
        RECT 76.905 183.985 77.075 184.175 ;
        RECT 78.745 184.030 78.905 184.140 ;
        RECT 79.205 183.985 79.375 184.175 ;
        RECT 83.805 183.985 83.975 184.175 ;
        RECT 84.270 183.985 84.440 184.175 ;
        RECT 85.185 184.005 85.355 184.195 ;
        RECT 87.025 184.005 87.195 184.195 ;
        RECT 88.405 183.985 88.575 184.175 ;
        RECT 89.380 184.035 89.500 184.145 ;
        RECT 93.190 183.985 93.360 184.175 ;
        RECT 96.225 184.005 96.395 184.195 ;
        RECT 96.740 184.035 96.860 184.145 ;
        RECT 100.550 184.005 100.720 184.195 ;
        RECT 101.340 184.035 101.460 184.145 ;
        RECT 102.665 183.985 102.835 184.175 ;
        RECT 103.585 184.005 103.755 184.195 ;
        RECT 104.045 183.985 104.215 184.175 ;
        RECT 107.450 184.005 107.620 184.195 ;
        RECT 108.240 184.035 108.360 184.145 ;
        RECT 109.565 183.985 109.735 184.175 ;
        RECT 110.030 183.985 110.200 184.175 ;
        RECT 110.945 184.005 111.115 184.195 ;
        RECT 114.165 184.030 114.325 184.140 ;
        RECT 114.810 184.005 114.980 184.195 ;
        RECT 115.085 183.985 115.255 184.175 ;
        RECT 116.925 184.030 117.085 184.140 ;
        RECT 118.950 184.005 119.120 184.195 ;
        RECT 120.605 183.985 120.775 184.195 ;
        RECT 126.125 183.985 126.295 184.195 ;
        RECT 127.505 183.985 127.675 184.195 ;
        RECT 20.645 183.175 22.015 183.985 ;
        RECT 22.485 183.175 27.995 183.985 ;
        RECT 28.005 183.305 37.195 183.985 ;
        RECT 32.515 183.085 33.445 183.305 ;
        RECT 36.275 183.075 37.195 183.305 ;
        RECT 37.215 183.115 37.645 183.900 ;
        RECT 37.665 183.175 40.415 183.985 ;
        RECT 40.425 183.305 49.615 183.985 ;
        RECT 40.425 183.075 41.345 183.305 ;
        RECT 44.175 183.085 45.105 183.305 ;
        RECT 49.625 183.205 50.995 183.985 ;
        RECT 51.465 183.175 55.135 183.985 ;
        RECT 55.145 183.175 60.655 183.985 ;
        RECT 60.665 183.205 62.035 183.985 ;
        RECT 62.975 183.115 63.405 183.900 ;
        RECT 63.425 183.175 66.175 183.985 ;
        RECT 66.185 183.175 71.695 183.985 ;
        RECT 71.715 183.945 72.635 183.985 ;
        RECT 71.705 183.755 72.635 183.945 ;
        RECT 74.725 183.755 76.295 183.985 ;
        RECT 71.705 183.395 76.295 183.755 ;
        RECT 71.715 183.305 76.295 183.395 ;
        RECT 71.715 183.075 74.715 183.305 ;
        RECT 76.775 183.075 78.125 183.985 ;
        RECT 79.075 183.075 80.425 183.985 ;
        RECT 80.445 183.175 84.115 183.985 ;
        RECT 84.125 183.075 86.735 183.985 ;
        RECT 86.885 183.175 88.715 183.985 ;
        RECT 88.735 183.115 89.165 183.900 ;
        RECT 89.875 183.305 93.775 183.985 ;
        RECT 92.845 183.075 93.775 183.305 ;
        RECT 93.785 183.305 102.975 183.985 ;
        RECT 93.785 183.075 94.705 183.305 ;
        RECT 97.535 183.085 98.465 183.305 ;
        RECT 102.985 183.175 104.355 183.985 ;
        RECT 104.365 183.175 109.875 183.985 ;
        RECT 109.885 183.075 113.360 183.985 ;
        RECT 114.495 183.115 114.925 183.900 ;
        RECT 114.945 183.205 116.315 183.985 ;
        RECT 117.245 183.175 120.915 183.985 ;
        RECT 120.925 183.175 126.435 183.985 ;
        RECT 126.445 183.175 127.815 183.985 ;
      LAYER nwell ;
        RECT 20.450 179.955 128.010 182.785 ;
      LAYER pwell ;
        RECT 20.645 178.755 22.015 179.565 ;
        RECT 22.485 178.755 24.315 179.565 ;
        RECT 24.335 178.840 24.765 179.625 ;
        RECT 24.785 178.755 26.155 179.565 ;
        RECT 26.165 178.755 29.835 179.565 ;
        RECT 29.845 178.755 35.355 179.565 ;
        RECT 35.365 178.755 36.735 179.535 ;
        RECT 36.745 179.435 37.675 179.665 ;
        RECT 36.745 178.755 40.645 179.435 ;
        RECT 40.885 178.755 46.395 179.565 ;
        RECT 46.405 178.755 49.880 179.665 ;
        RECT 50.095 178.840 50.525 179.625 ;
        RECT 51.005 178.755 52.835 179.565 ;
        RECT 56.045 179.435 56.975 179.665 ;
        RECT 60.185 179.435 61.115 179.665 ;
        RECT 53.075 178.755 56.975 179.435 ;
        RECT 57.215 178.755 61.115 179.435 ;
        RECT 61.135 178.755 63.875 179.435 ;
        RECT 63.885 178.755 67.555 179.565 ;
        RECT 67.565 179.435 68.910 179.665 ;
        RECT 69.890 179.435 71.235 179.665 ;
        RECT 67.565 178.755 69.395 179.435 ;
        RECT 69.405 178.755 71.235 179.435 ;
        RECT 72.165 178.755 75.835 179.565 ;
        RECT 75.855 178.840 76.285 179.625 ;
        RECT 76.765 178.755 80.435 179.565 ;
        RECT 80.445 178.755 83.185 179.435 ;
        RECT 83.205 178.755 86.680 179.665 ;
        RECT 87.805 178.755 93.315 179.565 ;
        RECT 93.325 178.755 94.695 179.535 ;
        RECT 94.705 178.755 96.535 179.565 ;
        RECT 96.555 178.755 97.905 179.665 ;
        RECT 98.385 178.755 100.215 179.565 ;
        RECT 100.225 178.755 101.595 179.535 ;
        RECT 101.615 178.840 102.045 179.625 ;
        RECT 102.075 178.755 103.425 179.665 ;
        RECT 103.905 178.755 106.655 179.565 ;
        RECT 106.665 178.755 110.140 179.665 ;
        RECT 110.540 178.755 114.015 179.665 ;
        RECT 114.025 178.755 115.855 179.565 ;
        RECT 115.875 178.755 117.225 179.665 ;
        RECT 117.245 179.435 118.165 179.665 ;
        RECT 120.995 179.435 121.925 179.655 ;
        RECT 117.245 178.755 126.435 179.435 ;
        RECT 126.445 178.755 127.815 179.565 ;
        RECT 20.785 178.545 20.955 178.755 ;
        RECT 22.220 178.595 22.340 178.705 ;
        RECT 24.005 178.565 24.175 178.755 ;
        RECT 25.845 178.545 26.015 178.755 ;
        RECT 29.525 178.565 29.695 178.755 ;
        RECT 31.365 178.545 31.535 178.735 ;
        RECT 35.045 178.565 35.215 178.755 ;
        RECT 36.425 178.565 36.595 178.755 ;
        RECT 36.885 178.545 37.055 178.735 ;
        RECT 37.160 178.565 37.330 178.755 ;
        RECT 38.725 178.545 38.895 178.735 ;
        RECT 42.400 178.545 42.570 178.735 ;
        RECT 42.870 178.545 43.040 178.735 ;
        RECT 46.085 178.565 46.255 178.755 ;
        RECT 46.550 178.565 46.720 178.755 ;
        RECT 49.760 178.545 49.930 178.735 ;
        RECT 50.740 178.595 50.860 178.705 ;
        RECT 52.525 178.565 52.695 178.755 ;
        RECT 53.440 178.545 53.610 178.735 ;
        RECT 56.390 178.565 56.560 178.755 ;
        RECT 60.530 178.565 60.700 178.755 ;
        RECT 62.645 178.545 62.815 178.735 ;
        RECT 63.565 178.565 63.735 178.755 ;
        RECT 64.485 178.545 64.655 178.735 ;
        RECT 65.405 178.590 65.565 178.700 ;
        RECT 67.245 178.545 67.415 178.755 ;
        RECT 67.705 178.565 67.875 178.735 ;
        RECT 69.085 178.565 69.255 178.755 ;
        RECT 69.545 178.565 69.715 178.755 ;
        RECT 70.925 178.565 71.095 178.735 ;
        RECT 71.845 178.600 72.005 178.710 ;
        RECT 67.805 178.545 67.875 178.565 ;
        RECT 71.025 178.545 71.095 178.565 ;
        RECT 74.145 178.545 74.315 178.735 ;
        RECT 75.525 178.565 75.695 178.755 ;
        RECT 76.500 178.595 76.620 178.705 ;
        RECT 79.205 178.545 79.375 178.735 ;
        RECT 79.670 178.545 79.840 178.735 ;
        RECT 80.125 178.565 80.295 178.755 ;
        RECT 80.585 178.565 80.755 178.755 ;
        RECT 83.350 178.545 83.520 178.755 ;
        RECT 87.485 178.600 87.645 178.710 ;
        RECT 88.405 178.545 88.575 178.735 ;
        RECT 89.330 178.545 89.500 178.735 ;
        RECT 93.005 178.565 93.175 178.755 ;
        RECT 93.465 178.565 93.635 178.755 ;
        RECT 95.305 178.545 95.475 178.735 ;
        RECT 96.225 178.565 96.395 178.755 ;
        RECT 97.605 178.565 97.775 178.755 ;
        RECT 98.120 178.595 98.240 178.705 ;
        RECT 98.980 178.545 99.150 178.735 ;
        RECT 99.905 178.565 100.075 178.755 ;
        RECT 100.365 178.565 100.535 178.755 ;
        RECT 103.125 178.565 103.295 178.755 ;
        RECT 103.640 178.595 103.760 178.705 ;
        RECT 106.345 178.565 106.515 178.755 ;
        RECT 106.810 178.565 106.980 178.755 ;
        RECT 108.185 178.545 108.355 178.735 ;
        RECT 108.650 178.545 108.820 178.735 ;
        RECT 112.380 178.595 112.500 178.705 ;
        RECT 113.700 178.565 113.870 178.755 ;
        RECT 114.165 178.545 114.335 178.735 ;
        RECT 115.545 178.565 115.715 178.755 ;
        RECT 116.005 178.565 116.175 178.755 ;
        RECT 118.305 178.545 118.475 178.735 ;
        RECT 118.765 178.545 118.935 178.735 ;
        RECT 120.200 178.595 120.320 178.705 ;
        RECT 121.985 178.545 122.155 178.735 ;
        RECT 122.445 178.545 122.615 178.735 ;
        RECT 126.125 178.545 126.295 178.755 ;
        RECT 127.505 178.545 127.675 178.755 ;
        RECT 20.645 177.735 22.015 178.545 ;
        RECT 22.485 177.735 26.155 178.545 ;
        RECT 26.165 177.735 31.675 178.545 ;
        RECT 31.685 177.735 37.195 178.545 ;
        RECT 37.215 177.675 37.645 178.460 ;
        RECT 37.665 177.735 39.035 178.545 ;
        RECT 39.240 177.635 42.715 178.545 ;
        RECT 42.725 177.635 46.200 178.545 ;
        RECT 46.600 177.635 50.075 178.545 ;
        RECT 50.280 177.635 53.755 178.545 ;
        RECT 53.765 177.865 62.955 178.545 ;
        RECT 53.765 177.635 54.685 177.865 ;
        RECT 57.515 177.645 58.445 177.865 ;
        RECT 62.975 177.675 63.405 178.460 ;
        RECT 63.425 177.765 64.795 178.545 ;
        RECT 65.725 177.865 67.555 178.545 ;
        RECT 67.805 178.315 70.075 178.545 ;
        RECT 71.025 178.315 73.295 178.545 ;
        RECT 65.725 177.635 67.070 177.865 ;
        RECT 67.805 177.635 70.560 178.315 ;
        RECT 71.025 177.635 73.780 178.315 ;
        RECT 74.005 177.865 75.835 178.545 ;
        RECT 74.490 177.635 75.835 177.865 ;
        RECT 75.845 177.735 79.515 178.545 ;
        RECT 79.525 177.635 83.000 178.545 ;
        RECT 83.205 177.635 86.680 178.545 ;
        RECT 86.885 177.735 88.715 178.545 ;
        RECT 88.735 177.675 89.165 178.460 ;
        RECT 89.185 177.635 91.795 178.545 ;
        RECT 91.945 177.735 95.615 178.545 ;
        RECT 95.820 177.635 99.295 178.545 ;
        RECT 99.305 177.865 108.495 178.545 ;
        RECT 99.305 177.635 100.225 177.865 ;
        RECT 103.055 177.645 103.985 177.865 ;
        RECT 108.505 177.635 111.980 178.545 ;
        RECT 112.645 177.735 114.475 178.545 ;
        RECT 114.495 177.675 114.925 178.460 ;
        RECT 114.945 177.735 118.615 178.545 ;
        RECT 118.635 177.635 119.985 178.545 ;
        RECT 120.465 177.735 122.295 178.545 ;
        RECT 122.305 177.765 123.675 178.545 ;
        RECT 123.685 177.735 126.435 178.545 ;
        RECT 126.445 177.735 127.815 178.545 ;
      LAYER nwell ;
        RECT 20.450 174.515 128.010 177.345 ;
      LAYER pwell ;
        RECT 20.645 173.315 22.015 174.125 ;
        RECT 22.485 173.315 24.315 174.125 ;
        RECT 24.335 173.400 24.765 174.185 ;
        RECT 29.295 173.995 30.225 174.215 ;
        RECT 33.055 173.995 33.975 174.225 ;
        RECT 24.785 173.315 33.975 173.995 ;
        RECT 34.445 173.315 36.275 174.125 ;
        RECT 36.285 173.315 39.760 174.225 ;
        RECT 40.160 173.315 43.635 174.225 ;
        RECT 44.565 173.315 50.075 174.125 ;
        RECT 50.095 173.400 50.525 174.185 ;
        RECT 50.545 173.315 53.295 174.125 ;
        RECT 53.305 173.315 56.780 174.225 ;
        RECT 56.985 173.315 60.460 174.225 ;
        RECT 60.675 173.315 62.025 174.225 ;
        RECT 62.505 173.315 68.015 174.125 ;
        RECT 68.025 173.995 69.370 174.225 ;
        RECT 68.025 173.315 69.855 173.995 ;
        RECT 69.905 173.315 74.455 174.225 ;
        RECT 74.475 173.315 75.825 174.225 ;
        RECT 75.855 173.400 76.285 174.185 ;
        RECT 76.545 173.545 79.300 174.225 ;
        RECT 76.545 173.315 78.815 173.545 ;
        RECT 79.985 173.315 81.815 174.125 ;
        RECT 81.825 173.315 85.300 174.225 ;
        RECT 86.865 173.995 87.785 174.215 ;
        RECT 93.865 174.115 94.785 174.225 ;
        RECT 92.450 173.995 94.785 174.115 ;
        RECT 85.505 173.315 94.785 173.995 ;
        RECT 95.625 173.315 97.455 174.125 ;
        RECT 100.665 173.995 101.595 174.225 ;
        RECT 97.695 173.315 101.595 173.995 ;
        RECT 101.615 173.400 102.045 174.185 ;
        RECT 102.525 173.315 104.355 174.125 ;
        RECT 104.365 173.315 105.735 174.095 ;
        RECT 106.205 173.315 108.035 174.125 ;
        RECT 108.240 173.315 111.715 174.225 ;
        RECT 114.925 173.995 115.855 174.225 ;
        RECT 111.955 173.315 115.855 173.995 ;
        RECT 115.865 173.995 116.785 174.225 ;
        RECT 119.615 173.995 120.545 174.215 ;
        RECT 115.865 173.315 125.055 173.995 ;
        RECT 125.065 173.315 126.435 174.125 ;
        RECT 126.445 173.315 127.815 174.125 ;
        RECT 20.785 173.105 20.955 173.315 ;
        RECT 22.220 173.155 22.340 173.265 ;
        RECT 23.545 173.105 23.715 173.295 ;
        RECT 24.005 173.125 24.175 173.315 ;
        RECT 24.925 173.105 25.095 173.315 ;
        RECT 25.385 173.105 25.555 173.295 ;
        RECT 34.180 173.155 34.300 173.265 ;
        RECT 35.505 173.105 35.675 173.295 ;
        RECT 35.965 173.125 36.135 173.315 ;
        RECT 36.430 173.125 36.600 173.315 ;
        RECT 36.885 173.105 37.055 173.295 ;
        RECT 38.265 173.150 38.425 173.260 ;
        RECT 41.945 173.105 42.115 173.295 ;
        RECT 42.405 173.105 42.575 173.295 ;
        RECT 43.320 173.125 43.490 173.315 ;
        RECT 43.790 173.105 43.960 173.295 ;
        RECT 44.245 173.160 44.405 173.270 ;
        RECT 47.465 173.105 47.635 173.295 ;
        RECT 49.765 173.125 49.935 173.315 ;
        RECT 52.985 173.125 53.155 173.315 ;
        RECT 53.450 173.125 53.620 173.315 ;
        RECT 57.130 173.260 57.300 173.315 ;
        RECT 57.125 173.150 57.300 173.260 ;
        RECT 57.130 173.125 57.300 173.150 ;
        RECT 61.725 173.125 61.895 173.315 ;
        RECT 62.240 173.155 62.360 173.265 ;
        RECT 62.645 173.105 62.815 173.295 ;
        RECT 63.620 173.155 63.740 173.265 ;
        RECT 67.705 173.125 67.875 173.315 ;
        RECT 69.085 173.105 69.255 173.295 ;
        RECT 69.545 173.125 69.715 173.315 ;
        RECT 72.305 173.125 72.475 173.295 ;
        RECT 72.305 173.105 72.375 173.125 ;
        RECT 72.765 173.105 72.935 173.295 ;
        RECT 74.145 173.125 74.315 173.315 ;
        RECT 75.525 173.125 75.695 173.315 ;
        RECT 76.545 173.295 76.615 173.315 ;
        RECT 76.445 173.125 76.615 173.295 ;
        RECT 77.420 173.155 77.540 173.265 ;
        RECT 79.720 173.155 79.840 173.265 ;
        RECT 81.505 173.125 81.675 173.315 ;
        RECT 81.970 173.125 82.140 173.315 ;
        RECT 82.885 173.105 83.055 173.295 ;
        RECT 83.345 173.105 83.515 173.295 ;
        RECT 85.000 173.105 85.170 173.295 ;
        RECT 85.645 173.125 85.815 173.315 ;
        RECT 89.785 173.150 89.945 173.260 ;
        RECT 91.165 173.105 91.335 173.295 ;
        RECT 93.005 173.105 93.175 173.295 ;
        RECT 94.385 173.105 94.555 173.295 ;
        RECT 94.900 173.155 95.020 173.265 ;
        RECT 95.360 173.155 95.480 173.265 ;
        RECT 97.145 173.125 97.315 173.315 ;
        RECT 98.525 173.105 98.695 173.295 ;
        RECT 98.985 173.105 99.155 173.295 ;
        RECT 101.010 173.125 101.180 173.315 ;
        RECT 102.260 173.155 102.380 173.265 ;
        RECT 104.045 173.125 104.215 173.315 ;
        RECT 104.505 173.125 104.675 173.315 ;
        RECT 105.940 173.155 106.060 173.265 ;
        RECT 107.725 173.125 107.895 173.315 ;
        RECT 108.645 173.150 108.805 173.260 ;
        RECT 111.400 173.125 111.570 173.315 ;
        RECT 114.165 173.105 114.335 173.295 ;
        RECT 115.270 173.125 115.440 173.315 ;
        RECT 115.545 173.150 115.705 173.260 ;
        RECT 119.410 173.105 119.580 173.295 ;
        RECT 120.200 173.155 120.320 173.265 ;
        RECT 120.605 173.105 120.775 173.295 ;
        RECT 123.365 173.105 123.535 173.295 ;
        RECT 124.745 173.125 124.915 173.315 ;
        RECT 126.125 173.105 126.295 173.315 ;
        RECT 127.505 173.105 127.675 173.315 ;
        RECT 20.645 172.295 22.015 173.105 ;
        RECT 22.025 172.295 23.855 173.105 ;
        RECT 23.875 172.195 25.225 173.105 ;
        RECT 25.255 172.195 26.605 173.105 ;
        RECT 26.625 172.425 35.815 173.105 ;
        RECT 26.625 172.195 27.545 172.425 ;
        RECT 30.375 172.205 31.305 172.425 ;
        RECT 35.825 172.295 37.195 173.105 ;
        RECT 37.215 172.235 37.645 173.020 ;
        RECT 38.585 172.295 42.255 173.105 ;
        RECT 42.275 172.195 43.625 173.105 ;
        RECT 43.645 172.195 47.120 173.105 ;
        RECT 47.325 172.425 56.430 173.105 ;
        RECT 57.445 172.295 62.955 173.105 ;
        RECT 62.975 172.235 63.405 173.020 ;
        RECT 63.885 172.295 69.395 173.105 ;
        RECT 70.105 172.875 72.375 173.105 ;
        RECT 69.620 172.195 72.375 172.875 ;
        RECT 72.625 172.875 74.195 173.105 ;
        RECT 76.285 173.065 77.205 173.105 ;
        RECT 76.285 172.875 77.215 173.065 ;
        RECT 72.625 172.515 77.215 172.875 ;
        RECT 72.625 172.425 77.205 172.515 ;
        RECT 74.205 172.195 77.205 172.425 ;
        RECT 77.685 172.295 83.195 173.105 ;
        RECT 83.205 172.325 84.575 173.105 ;
        RECT 84.585 172.425 88.485 173.105 ;
        RECT 84.585 172.195 85.515 172.425 ;
        RECT 88.735 172.235 89.165 173.020 ;
        RECT 90.115 172.195 91.465 173.105 ;
        RECT 91.485 172.295 93.315 173.105 ;
        RECT 93.335 172.195 94.685 173.105 ;
        RECT 95.165 172.295 98.835 173.105 ;
        RECT 98.845 172.425 107.950 173.105 ;
        RECT 108.965 172.295 114.475 173.105 ;
        RECT 114.495 172.235 114.925 173.020 ;
        RECT 116.095 172.425 119.995 173.105 ;
        RECT 119.065 172.195 119.995 172.425 ;
        RECT 120.465 172.325 121.835 173.105 ;
        RECT 121.845 172.425 123.675 173.105 ;
        RECT 123.685 172.295 126.435 173.105 ;
        RECT 126.445 172.295 127.815 173.105 ;
      LAYER nwell ;
        RECT 20.450 169.075 128.010 171.905 ;
      LAYER pwell ;
        RECT 20.645 167.875 22.015 168.685 ;
        RECT 22.945 167.875 24.315 168.655 ;
        RECT 24.335 167.960 24.765 168.745 ;
        RECT 33.985 168.555 34.905 168.785 ;
        RECT 37.735 168.555 38.665 168.775 ;
        RECT 49.145 168.555 50.075 168.785 ;
        RECT 24.870 167.875 33.975 168.555 ;
        RECT 33.985 167.875 43.175 168.555 ;
        RECT 43.185 167.875 44.550 168.555 ;
        RECT 46.175 167.875 50.075 168.555 ;
        RECT 50.095 167.960 50.525 168.745 ;
        RECT 50.555 167.875 53.295 168.555 ;
        RECT 53.685 167.875 56.110 168.555 ;
        RECT 57.585 167.875 60.195 168.785 ;
        RECT 60.345 167.875 62.955 168.785 ;
        RECT 62.975 167.875 65.715 168.555 ;
        RECT 66.185 167.875 68.015 168.685 ;
        RECT 68.025 167.875 73.535 168.685 ;
        RECT 73.545 168.555 74.890 168.785 ;
        RECT 73.545 167.875 75.375 168.555 ;
        RECT 75.855 167.960 76.285 168.745 ;
        RECT 76.305 167.875 78.135 168.685 ;
        RECT 78.145 167.875 80.885 168.555 ;
        RECT 80.905 167.875 83.655 168.685 ;
        RECT 86.865 168.555 87.795 168.785 ;
        RECT 83.895 167.875 87.795 168.555 ;
        RECT 87.890 167.875 96.995 168.555 ;
        RECT 97.005 167.875 98.835 168.685 ;
        RECT 98.855 167.875 100.205 168.785 ;
        RECT 100.225 167.875 101.595 168.685 ;
        RECT 101.615 167.960 102.045 168.745 ;
        RECT 102.065 167.875 103.435 168.655 ;
        RECT 103.455 167.875 104.805 168.785 ;
        RECT 105.295 167.875 108.035 168.555 ;
        RECT 108.045 167.875 109.875 168.685 ;
        RECT 109.895 167.875 111.245 168.785 ;
        RECT 114.465 168.555 115.395 168.785 ;
        RECT 111.495 167.875 115.395 168.555 ;
        RECT 115.405 167.875 116.775 168.685 ;
        RECT 116.795 167.875 118.145 168.785 ;
        RECT 118.305 167.875 120.915 168.785 ;
        RECT 120.925 167.875 126.435 168.685 ;
        RECT 126.445 167.875 127.815 168.685 ;
        RECT 20.785 167.665 20.955 167.875 ;
        RECT 22.625 167.720 22.785 167.830 ;
        RECT 23.085 167.685 23.255 167.875 ;
        RECT 27.225 167.665 27.395 167.855 ;
        RECT 27.960 167.665 28.130 167.855 ;
        RECT 32.285 167.710 32.445 167.820 ;
        RECT 33.020 167.665 33.190 167.855 ;
        RECT 33.665 167.685 33.835 167.875 ;
        RECT 36.940 167.715 37.060 167.825 ;
        RECT 38.725 167.665 38.895 167.855 ;
        RECT 39.185 167.665 39.355 167.855 ;
        RECT 42.865 167.685 43.035 167.875 ;
        RECT 44.705 167.685 44.875 167.855 ;
        RECT 45.625 167.720 45.785 167.830 ;
        RECT 49.305 167.665 49.475 167.855 ;
        RECT 49.490 167.685 49.660 167.875 ;
        RECT 52.985 167.685 53.155 167.875 ;
        RECT 59.880 167.855 60.050 167.875 ;
        RECT 56.205 167.685 56.375 167.855 ;
        RECT 57.125 167.720 57.285 167.830 ;
        RECT 58.505 167.665 58.675 167.855 ;
        RECT 59.880 167.685 60.055 167.855 ;
        RECT 59.885 167.665 60.055 167.685 ;
        RECT 60.350 167.665 60.520 167.855 ;
        RECT 62.640 167.685 62.810 167.875 ;
        RECT 64.025 167.710 64.185 167.820 ;
        RECT 64.485 167.665 64.655 167.855 ;
        RECT 65.405 167.685 65.575 167.875 ;
        RECT 65.920 167.715 66.040 167.825 ;
        RECT 67.705 167.685 67.875 167.875 ;
        RECT 68.625 167.665 68.795 167.855 ;
        RECT 73.225 167.685 73.395 167.875 ;
        RECT 74.145 167.665 74.315 167.855 ;
        RECT 74.605 167.665 74.775 167.855 ;
        RECT 75.065 167.685 75.235 167.875 ;
        RECT 75.580 167.715 75.700 167.825 ;
        RECT 77.825 167.685 77.995 167.875 ;
        RECT 78.285 167.685 78.455 167.875 ;
        RECT 78.745 167.665 78.915 167.855 ;
        RECT 83.345 167.685 83.515 167.875 ;
        RECT 87.210 167.685 87.380 167.875 ;
        RECT 88.405 167.665 88.575 167.855 ;
        RECT 90.245 167.665 90.415 167.855 ;
        RECT 91.625 167.665 91.795 167.855 ;
        RECT 92.085 167.665 92.255 167.855 ;
        RECT 93.520 167.715 93.640 167.825 ;
        RECT 95.305 167.685 95.475 167.855 ;
        RECT 96.685 167.685 96.855 167.875 ;
        RECT 98.525 167.685 98.695 167.875 ;
        RECT 98.985 167.685 99.155 167.875 ;
        RECT 101.285 167.685 101.455 167.875 ;
        RECT 102.205 167.685 102.375 167.875 ;
        RECT 103.585 167.685 103.755 167.875 ;
        RECT 104.965 167.825 105.135 167.855 ;
        RECT 104.965 167.715 105.140 167.825 ;
        RECT 104.965 167.665 105.135 167.715 ;
        RECT 107.725 167.685 107.895 167.875 ;
        RECT 109.565 167.685 109.735 167.875 ;
        RECT 110.945 167.685 111.115 167.875 ;
        RECT 114.165 167.665 114.335 167.855 ;
        RECT 114.810 167.685 114.980 167.875 ;
        RECT 115.140 167.715 115.260 167.825 ;
        RECT 116.465 167.685 116.635 167.875 ;
        RECT 116.925 167.685 117.095 167.875 ;
        RECT 120.600 167.685 120.770 167.875 ;
        RECT 124.285 167.665 124.455 167.855 ;
        RECT 126.125 167.665 126.295 167.875 ;
        RECT 127.505 167.665 127.675 167.875 ;
        RECT 20.645 166.855 22.015 167.665 ;
        RECT 22.025 166.855 27.535 167.665 ;
        RECT 27.545 166.985 31.445 167.665 ;
        RECT 32.605 166.985 36.505 167.665 ;
        RECT 27.545 166.755 28.475 166.985 ;
        RECT 32.605 166.755 33.535 166.985 ;
        RECT 37.215 166.795 37.645 167.580 ;
        RECT 37.665 166.855 39.035 167.665 ;
        RECT 39.045 166.885 40.415 167.665 ;
        RECT 40.425 166.985 49.615 167.665 ;
        RECT 49.625 166.985 58.815 167.665 ;
        RECT 40.425 166.755 41.345 166.985 ;
        RECT 44.175 166.765 45.105 166.985 ;
        RECT 49.625 166.755 50.545 166.985 ;
        RECT 53.375 166.765 54.305 166.985 ;
        RECT 58.825 166.855 60.195 167.665 ;
        RECT 60.205 166.755 62.815 167.665 ;
        RECT 62.975 166.795 63.405 167.580 ;
        RECT 64.345 166.885 65.715 167.665 ;
        RECT 66.185 166.855 68.935 167.665 ;
        RECT 68.945 166.855 74.455 167.665 ;
        RECT 74.465 166.755 77.185 167.665 ;
        RECT 77.225 166.855 79.055 167.665 ;
        RECT 79.435 166.985 88.715 167.665 ;
        RECT 79.435 166.865 81.770 166.985 ;
        RECT 79.435 166.755 80.355 166.865 ;
        RECT 86.435 166.765 87.355 166.985 ;
        RECT 88.735 166.795 89.165 167.580 ;
        RECT 89.185 166.885 90.555 167.665 ;
        RECT 90.575 166.755 91.925 167.665 ;
        RECT 91.945 166.885 93.315 167.665 ;
        RECT 93.785 166.985 95.150 167.665 ;
        RECT 95.995 166.985 105.275 167.665 ;
        RECT 105.285 166.985 114.475 167.665 ;
        RECT 95.995 166.865 98.330 166.985 ;
        RECT 95.995 166.755 96.915 166.865 ;
        RECT 102.995 166.765 103.915 166.985 ;
        RECT 105.285 166.755 106.205 166.985 ;
        RECT 109.035 166.765 109.965 166.985 ;
        RECT 114.495 166.795 114.925 167.580 ;
        RECT 115.405 166.985 124.595 167.665 ;
        RECT 115.405 166.755 116.325 166.985 ;
        RECT 119.155 166.765 120.085 166.985 ;
        RECT 124.605 166.855 126.435 167.665 ;
        RECT 126.445 166.855 127.815 167.665 ;
      LAYER nwell ;
        RECT 20.450 163.635 128.010 166.465 ;
      LAYER pwell ;
        RECT 20.645 162.435 22.015 163.245 ;
        RECT 22.485 162.435 24.315 163.245 ;
        RECT 24.335 162.520 24.765 163.305 ;
        RECT 25.255 162.435 26.605 163.345 ;
        RECT 29.825 163.115 30.755 163.345 ;
        RECT 26.855 162.435 30.755 163.115 ;
        RECT 31.225 162.435 32.595 163.215 ;
        RECT 32.615 162.435 33.965 163.345 ;
        RECT 33.985 162.435 39.495 163.245 ;
        RECT 39.505 163.115 40.435 163.345 ;
        RECT 39.505 162.435 43.405 163.115 ;
        RECT 43.645 162.435 45.015 163.245 ;
        RECT 45.025 162.435 48.695 163.245 ;
        RECT 48.705 162.435 50.075 163.215 ;
        RECT 50.095 162.520 50.525 163.305 ;
        RECT 51.005 162.435 52.835 163.245 ;
        RECT 52.855 162.435 54.205 163.345 ;
        RECT 54.225 162.435 55.595 163.215 ;
        RECT 55.605 162.435 56.975 163.245 ;
        RECT 56.995 162.435 58.345 163.345 ;
        RECT 58.735 163.235 59.655 163.345 ;
        RECT 58.735 163.115 61.070 163.235 ;
        RECT 65.735 163.115 66.655 163.335 ;
        RECT 58.735 162.435 68.015 163.115 ;
        RECT 68.025 162.435 70.775 163.245 ;
        RECT 70.785 163.115 72.130 163.345 ;
        RECT 73.110 163.115 74.455 163.345 ;
        RECT 70.785 162.435 72.615 163.115 ;
        RECT 72.625 162.435 74.455 163.115 ;
        RECT 74.465 162.435 75.835 163.245 ;
        RECT 75.855 162.520 76.285 163.305 ;
        RECT 76.765 162.435 82.275 163.245 ;
        RECT 85.485 163.115 86.415 163.345 ;
        RECT 82.515 162.435 86.415 163.115 ;
        RECT 86.795 163.235 87.715 163.345 ;
        RECT 86.795 163.115 89.130 163.235 ;
        RECT 93.795 163.115 94.715 163.335 ;
        RECT 86.795 162.435 96.075 163.115 ;
        RECT 96.085 162.435 97.455 163.245 ;
        RECT 100.665 163.115 101.595 163.345 ;
        RECT 97.695 162.435 101.595 163.115 ;
        RECT 101.615 162.520 102.045 163.305 ;
        RECT 102.435 163.235 103.355 163.345 ;
        RECT 102.435 163.115 104.770 163.235 ;
        RECT 109.435 163.115 110.355 163.335 ;
        RECT 102.435 162.435 111.715 163.115 ;
        RECT 112.185 162.435 114.015 163.245 ;
        RECT 114.025 162.435 115.395 163.215 ;
        RECT 118.605 163.115 119.535 163.345 ;
        RECT 115.635 162.435 119.535 163.115 ;
        RECT 120.465 162.435 121.835 163.215 ;
        RECT 122.765 162.435 126.435 163.245 ;
        RECT 126.445 162.435 127.815 163.245 ;
        RECT 20.785 162.225 20.955 162.435 ;
        RECT 22.220 162.275 22.340 162.385 ;
        RECT 22.625 162.270 22.785 162.380 ;
        RECT 24.005 162.245 24.175 162.435 ;
        RECT 24.980 162.275 25.100 162.385 ;
        RECT 26.305 162.245 26.475 162.435 ;
        RECT 30.170 162.245 30.340 162.435 ;
        RECT 30.960 162.275 31.080 162.385 ;
        RECT 31.365 162.245 31.535 162.435 ;
        RECT 32.285 162.225 32.455 162.415 ;
        RECT 32.745 162.245 32.915 162.435 ;
        RECT 33.665 162.225 33.835 162.415 ;
        RECT 35.505 162.225 35.675 162.415 ;
        RECT 35.965 162.225 36.135 162.415 ;
        RECT 39.185 162.245 39.355 162.435 ;
        RECT 39.920 162.245 40.090 162.435 ;
        RECT 44.705 162.415 44.875 162.435 ;
        RECT 48.385 162.415 48.555 162.435 ;
        RECT 41.020 162.225 41.190 162.415 ;
        RECT 44.700 162.245 44.875 162.415 ;
        RECT 48.380 162.245 48.555 162.415 ;
        RECT 49.765 162.245 49.935 162.435 ;
        RECT 50.740 162.275 50.860 162.385 ;
        RECT 44.700 162.225 44.870 162.245 ;
        RECT 48.380 162.225 48.550 162.245 ;
        RECT 52.250 162.225 52.420 162.415 ;
        RECT 52.525 162.245 52.695 162.435 ;
        RECT 53.040 162.275 53.160 162.385 ;
        RECT 53.905 162.245 54.075 162.435 ;
        RECT 54.365 162.245 54.535 162.435 ;
        RECT 56.665 162.245 56.835 162.435 ;
        RECT 57.125 162.245 57.295 162.435 ;
        RECT 58.505 162.225 58.675 162.415 ;
        RECT 62.370 162.225 62.540 162.415 ;
        RECT 63.620 162.275 63.740 162.385 ;
        RECT 65.405 162.225 65.575 162.415 ;
        RECT 65.865 162.225 66.035 162.415 ;
        RECT 67.705 162.245 67.875 162.435 ;
        RECT 68.625 162.225 68.795 162.415 ;
        RECT 70.465 162.225 70.635 162.435 ;
        RECT 72.305 162.225 72.475 162.435 ;
        RECT 72.765 162.225 72.935 162.435 ;
        RECT 75.525 162.245 75.695 162.435 ;
        RECT 75.985 162.225 76.155 162.415 ;
        RECT 76.500 162.275 76.620 162.385 ;
        RECT 76.905 162.270 77.065 162.380 ;
        RECT 80.585 162.225 80.755 162.415 ;
        RECT 81.050 162.225 81.220 162.415 ;
        RECT 81.965 162.245 82.135 162.435 ;
        RECT 84.780 162.275 84.900 162.385 ;
        RECT 85.830 162.245 86.000 162.435 ;
        RECT 88.405 162.225 88.575 162.415 ;
        RECT 89.380 162.275 89.500 162.385 ;
        RECT 91.165 162.225 91.335 162.415 ;
        RECT 95.765 162.245 95.935 162.435 ;
        RECT 96.685 162.225 96.855 162.415 ;
        RECT 97.145 162.245 97.315 162.435 ;
        RECT 101.010 162.245 101.180 162.435 ;
        RECT 102.205 162.225 102.375 162.415 ;
        RECT 102.665 162.225 102.835 162.415 ;
        RECT 104.320 162.225 104.490 162.415 ;
        RECT 108.645 162.270 108.805 162.380 ;
        RECT 111.405 162.245 111.575 162.435 ;
        RECT 111.920 162.275 112.040 162.385 ;
        RECT 113.705 162.245 113.875 162.435 ;
        RECT 114.165 162.225 114.335 162.415 ;
        RECT 115.085 162.245 115.255 162.435 ;
        RECT 116.005 162.225 116.175 162.415 ;
        RECT 116.470 162.225 116.640 162.415 ;
        RECT 118.950 162.245 119.120 162.435 ;
        RECT 120.145 162.280 120.305 162.390 ;
        RECT 120.605 162.225 120.775 162.435 ;
        RECT 122.445 162.280 122.605 162.390 ;
        RECT 126.125 162.225 126.295 162.435 ;
        RECT 127.505 162.225 127.675 162.435 ;
        RECT 20.645 161.415 22.015 162.225 ;
        RECT 23.315 161.545 32.595 162.225 ;
        RECT 23.315 161.425 25.650 161.545 ;
        RECT 23.315 161.315 24.235 161.425 ;
        RECT 30.315 161.325 31.235 161.545 ;
        RECT 32.605 161.445 33.975 162.225 ;
        RECT 33.985 161.415 35.815 162.225 ;
        RECT 35.835 161.315 37.185 162.225 ;
        RECT 37.215 161.355 37.645 162.140 ;
        RECT 37.860 161.315 41.335 162.225 ;
        RECT 41.540 161.315 45.015 162.225 ;
        RECT 45.220 161.315 48.695 162.225 ;
        RECT 48.935 161.545 52.835 162.225 ;
        RECT 51.905 161.315 52.835 161.545 ;
        RECT 53.305 161.415 58.815 162.225 ;
        RECT 59.055 161.545 62.955 162.225 ;
        RECT 62.025 161.315 62.955 161.545 ;
        RECT 62.975 161.355 63.405 162.140 ;
        RECT 63.885 161.415 65.715 162.225 ;
        RECT 65.735 161.315 67.085 162.225 ;
        RECT 67.105 161.415 68.935 162.225 ;
        RECT 68.945 161.545 70.775 162.225 ;
        RECT 70.785 161.545 72.615 162.225 ;
        RECT 72.625 161.545 74.455 162.225 ;
        RECT 68.945 161.315 70.290 161.545 ;
        RECT 70.785 161.315 72.130 161.545 ;
        RECT 73.110 161.315 74.455 161.545 ;
        RECT 74.465 161.545 76.295 162.225 ;
        RECT 74.465 161.315 75.810 161.545 ;
        RECT 77.225 161.415 80.895 162.225 ;
        RECT 80.905 161.315 84.380 162.225 ;
        RECT 85.045 161.415 88.715 162.225 ;
        RECT 88.735 161.355 89.165 162.140 ;
        RECT 89.645 161.415 91.475 162.225 ;
        RECT 91.485 161.415 96.995 162.225 ;
        RECT 97.005 161.415 102.515 162.225 ;
        RECT 102.525 161.445 103.895 162.225 ;
        RECT 103.905 161.545 107.805 162.225 ;
        RECT 103.905 161.315 104.835 161.545 ;
        RECT 108.965 161.415 114.475 162.225 ;
        RECT 114.495 161.355 114.925 162.140 ;
        RECT 114.945 161.415 116.315 162.225 ;
        RECT 116.325 161.315 118.935 162.225 ;
        RECT 119.085 161.415 120.915 162.225 ;
        RECT 120.925 161.415 126.435 162.225 ;
        RECT 126.445 161.415 127.815 162.225 ;
      LAYER nwell ;
        RECT 20.450 158.195 128.010 161.025 ;
      LAYER pwell ;
        RECT 20.645 156.995 22.015 157.805 ;
        RECT 22.485 156.995 24.315 157.805 ;
        RECT 24.335 157.080 24.765 157.865 ;
        RECT 25.715 156.995 27.065 157.905 ;
        RECT 30.285 157.675 31.215 157.905 ;
        RECT 27.315 156.995 31.215 157.675 ;
        RECT 31.225 156.995 33.975 157.805 ;
        RECT 34.355 157.795 35.275 157.905 ;
        RECT 34.355 157.675 36.690 157.795 ;
        RECT 41.355 157.675 42.275 157.895 ;
        RECT 34.355 156.995 43.635 157.675 ;
        RECT 43.645 156.995 46.395 157.805 ;
        RECT 46.600 156.995 50.075 157.905 ;
        RECT 50.095 157.080 50.525 157.865 ;
        RECT 50.545 156.995 54.020 157.905 ;
        RECT 54.685 156.995 57.435 157.805 ;
        RECT 57.455 156.995 58.805 157.905 ;
        RECT 62.025 157.675 62.955 157.905 ;
        RECT 59.055 156.995 62.955 157.675 ;
        RECT 63.335 157.795 64.255 157.905 ;
        RECT 63.335 157.675 65.670 157.795 ;
        RECT 70.335 157.675 71.255 157.895 ;
        RECT 63.335 156.995 72.615 157.675 ;
        RECT 73.085 156.995 75.805 157.905 ;
        RECT 75.855 157.080 76.285 157.865 ;
        RECT 77.225 156.995 80.700 157.905 ;
        RECT 80.905 156.995 84.380 157.905 ;
        RECT 84.585 156.995 87.335 157.805 ;
        RECT 87.345 156.995 92.855 157.805 ;
        RECT 92.875 156.995 94.225 157.905 ;
        RECT 94.245 156.995 96.075 157.805 ;
        RECT 96.085 156.995 101.595 157.805 ;
        RECT 101.615 157.080 102.045 157.865 ;
        RECT 102.065 156.995 103.435 157.805 ;
        RECT 103.445 156.995 107.115 157.805 ;
        RECT 107.320 156.995 110.795 157.905 ;
        RECT 110.805 156.995 114.280 157.905 ;
        RECT 115.405 156.995 120.915 157.805 ;
        RECT 120.925 156.995 126.435 157.805 ;
        RECT 126.445 156.995 127.815 157.805 ;
        RECT 20.785 156.785 20.955 156.995 ;
        RECT 22.220 156.835 22.340 156.945 ;
        RECT 22.625 156.830 22.785 156.940 ;
        RECT 24.005 156.805 24.175 156.995 ;
        RECT 25.385 156.840 25.545 156.950 ;
        RECT 26.765 156.805 26.935 156.995 ;
        RECT 30.630 156.805 30.800 156.995 ;
        RECT 32.285 156.785 32.455 156.975 ;
        RECT 33.665 156.785 33.835 156.995 ;
        RECT 34.180 156.835 34.300 156.945 ;
        RECT 36.885 156.785 37.055 156.975 ;
        RECT 41.210 156.785 41.380 156.975 ;
        RECT 42.865 156.785 43.035 156.975 ;
        RECT 43.325 156.805 43.495 156.995 ;
        RECT 44.705 156.785 44.875 156.975 ;
        RECT 46.085 156.805 46.255 156.995 ;
        RECT 48.380 156.785 48.550 156.975 ;
        RECT 49.305 156.830 49.465 156.940 ;
        RECT 49.760 156.805 49.930 156.995 ;
        RECT 50.690 156.805 50.860 156.995 ;
        RECT 52.985 156.785 53.155 156.975 ;
        RECT 54.420 156.835 54.540 156.945 ;
        RECT 57.125 156.805 57.295 156.995 ;
        RECT 58.505 156.805 58.675 156.995 ;
        RECT 62.370 156.805 62.540 156.995 ;
        RECT 62.645 156.785 62.815 156.975 ;
        RECT 64.485 156.785 64.655 156.975 ;
        RECT 66.325 156.785 66.495 156.975 ;
        RECT 66.785 156.785 66.955 156.975 ;
        RECT 69.545 156.785 69.715 156.975 ;
        RECT 71.385 156.785 71.555 156.975 ;
        RECT 72.305 156.805 72.475 156.995 ;
        RECT 72.820 156.835 72.940 156.945 ;
        RECT 73.225 156.805 73.395 156.995 ;
        RECT 75.065 156.785 75.235 156.975 ;
        RECT 75.525 156.785 75.695 156.975 ;
        RECT 76.905 156.840 77.065 156.950 ;
        RECT 77.370 156.805 77.540 156.995 ;
        RECT 78.285 156.785 78.455 156.975 ;
        RECT 78.745 156.785 78.915 156.975 ;
        RECT 81.050 156.805 81.220 156.995 ;
        RECT 81.510 156.785 81.680 156.975 ;
        RECT 87.025 156.805 87.195 156.995 ;
        RECT 88.405 156.785 88.575 156.975 ;
        RECT 92.545 156.805 92.715 156.995 ;
        RECT 93.925 156.805 94.095 156.995 ;
        RECT 95.765 156.805 95.935 156.995 ;
        RECT 98.525 156.785 98.695 156.975 ;
        RECT 99.040 156.835 99.160 156.945 ;
        RECT 99.450 156.785 99.620 156.975 ;
        RECT 101.285 156.805 101.455 156.995 ;
        RECT 103.125 156.945 103.295 156.995 ;
        RECT 103.125 156.835 103.300 156.945 ;
        RECT 103.125 156.805 103.295 156.835 ;
        RECT 105.885 156.785 106.055 156.975 ;
        RECT 106.350 156.785 106.520 156.975 ;
        RECT 106.805 156.805 106.975 156.995 ;
        RECT 110.030 156.785 110.200 156.975 ;
        RECT 110.480 156.805 110.650 156.995 ;
        RECT 110.950 156.805 111.120 156.995 ;
        RECT 114.165 156.830 114.325 156.940 ;
        RECT 115.085 156.840 115.245 156.950 ;
        RECT 115.545 156.830 115.705 156.940 ;
        RECT 116.005 156.785 116.175 156.975 ;
        RECT 120.605 156.805 120.775 156.995 ;
        RECT 126.125 156.785 126.295 156.995 ;
        RECT 127.505 156.785 127.675 156.995 ;
        RECT 20.645 155.975 22.015 156.785 ;
        RECT 23.315 156.105 32.595 156.785 ;
        RECT 23.315 155.985 25.650 156.105 ;
        RECT 23.315 155.875 24.235 155.985 ;
        RECT 30.315 155.885 31.235 156.105 ;
        RECT 32.605 156.005 33.975 156.785 ;
        RECT 34.445 155.975 37.195 156.785 ;
        RECT 37.215 155.915 37.645 156.700 ;
        RECT 37.895 156.105 41.795 156.785 ;
        RECT 40.865 155.875 41.795 156.105 ;
        RECT 41.805 156.005 43.175 156.785 ;
        RECT 43.185 155.975 45.015 156.785 ;
        RECT 45.220 155.875 48.695 156.785 ;
        RECT 49.625 155.975 53.295 156.785 ;
        RECT 53.675 156.105 62.955 156.785 ;
        RECT 53.675 155.985 56.010 156.105 ;
        RECT 53.675 155.875 54.595 155.985 ;
        RECT 60.675 155.885 61.595 156.105 ;
        RECT 62.975 155.915 63.405 156.700 ;
        RECT 63.425 156.005 64.795 156.785 ;
        RECT 64.805 155.975 66.635 156.785 ;
        RECT 66.645 156.005 68.015 156.785 ;
        RECT 68.025 156.105 69.855 156.785 ;
        RECT 69.865 156.105 71.695 156.785 ;
        RECT 72.635 156.105 75.375 156.785 ;
        RECT 75.385 156.105 77.215 156.785 ;
        RECT 68.025 155.875 69.370 156.105 ;
        RECT 69.865 155.875 71.210 156.105 ;
        RECT 75.870 155.875 77.215 156.105 ;
        RECT 77.225 155.975 78.595 156.785 ;
        RECT 78.605 156.105 81.345 156.785 ;
        RECT 81.365 155.875 84.840 156.785 ;
        RECT 85.045 155.975 88.715 156.785 ;
        RECT 88.735 155.915 89.165 156.700 ;
        RECT 89.555 156.105 98.835 156.785 ;
        RECT 89.555 155.985 91.890 156.105 ;
        RECT 89.555 155.875 90.475 155.985 ;
        RECT 96.555 155.885 97.475 156.105 ;
        RECT 99.305 155.875 102.780 156.785 ;
        RECT 103.445 155.975 106.195 156.785 ;
        RECT 106.205 155.875 109.680 156.785 ;
        RECT 109.885 155.875 113.360 156.785 ;
        RECT 114.495 155.915 114.925 156.700 ;
        RECT 115.875 155.875 117.225 156.785 ;
        RECT 117.245 156.105 126.435 156.785 ;
        RECT 117.245 155.875 118.165 156.105 ;
        RECT 120.995 155.885 121.925 156.105 ;
        RECT 126.445 155.975 127.815 156.785 ;
      LAYER nwell ;
        RECT 20.450 152.755 128.010 155.585 ;
      LAYER pwell ;
        RECT 20.645 151.555 22.015 152.365 ;
        RECT 22.485 151.555 24.315 152.365 ;
        RECT 24.335 151.640 24.765 152.425 ;
        RECT 25.705 151.555 27.075 152.335 ;
        RECT 27.085 152.235 28.015 152.465 ;
        RECT 27.085 151.555 30.985 152.235 ;
        RECT 31.685 151.555 37.195 152.365 ;
        RECT 37.205 151.555 42.715 152.365 ;
        RECT 42.725 151.555 46.200 152.465 ;
        RECT 47.325 152.265 48.270 152.465 ;
        RECT 47.325 151.585 50.075 152.265 ;
        RECT 50.095 151.640 50.525 152.425 ;
        RECT 50.545 152.265 51.490 152.465 ;
        RECT 50.545 151.585 53.295 152.265 ;
        RECT 47.325 151.555 48.270 151.585 ;
        RECT 20.785 151.345 20.955 151.555 ;
        RECT 22.220 151.395 22.340 151.505 ;
        RECT 24.005 151.365 24.175 151.555 ;
        RECT 25.385 151.400 25.545 151.510 ;
        RECT 25.845 151.365 26.015 151.555 ;
        RECT 27.500 151.365 27.670 151.555 ;
        RECT 31.365 151.505 31.535 151.535 ;
        RECT 31.365 151.395 31.540 151.505 ;
        RECT 31.365 151.345 31.535 151.395 ;
        RECT 35.230 151.345 35.400 151.535 ;
        RECT 36.885 151.345 37.055 151.555 ;
        RECT 39.185 151.345 39.355 151.535 ;
        RECT 39.650 151.345 39.820 151.535 ;
        RECT 42.405 151.365 42.575 151.555 ;
        RECT 42.870 151.365 43.040 151.555 ;
        RECT 43.330 151.345 43.500 151.535 ;
        RECT 47.005 151.400 47.165 151.510 ;
        RECT 47.925 151.345 48.095 151.535 ;
        RECT 49.760 151.365 49.930 151.585 ;
        RECT 50.545 151.555 51.490 151.585 ;
        RECT 51.605 151.345 51.775 151.535 ;
        RECT 52.980 151.365 53.150 151.585 ;
        RECT 53.305 151.555 56.780 152.465 ;
        RECT 56.985 151.555 60.460 152.465 ;
        RECT 64.325 152.235 65.255 152.465 ;
        RECT 61.355 151.555 65.255 152.235 ;
        RECT 65.350 151.555 74.455 152.235 ;
        RECT 74.465 151.555 75.835 152.365 ;
        RECT 75.855 151.640 76.285 152.425 ;
        RECT 76.790 152.235 78.135 152.465 ;
        RECT 76.305 151.555 78.135 152.235 ;
        RECT 78.145 151.555 79.975 152.365 ;
        RECT 79.985 152.265 80.930 152.465 ;
        RECT 79.985 151.585 82.735 152.265 ;
        RECT 79.985 151.555 80.930 151.585 ;
        RECT 53.450 151.365 53.620 151.555 ;
        RECT 57.130 151.535 57.300 151.555 ;
        RECT 57.125 151.365 57.300 151.535 ;
        RECT 60.860 151.395 60.980 151.505 ;
        RECT 57.125 151.345 57.295 151.365 ;
        RECT 62.645 151.345 62.815 151.535 ;
        RECT 63.620 151.395 63.740 151.505 ;
        RECT 64.670 151.365 64.840 151.555 ;
        RECT 66.325 151.345 66.495 151.535 ;
        RECT 66.785 151.345 66.955 151.535 ;
        RECT 68.220 151.395 68.340 151.505 ;
        RECT 70.005 151.345 70.175 151.535 ;
        RECT 70.465 151.345 70.635 151.535 ;
        RECT 73.225 151.345 73.395 151.535 ;
        RECT 73.685 151.345 73.855 151.535 ;
        RECT 74.145 151.365 74.315 151.555 ;
        RECT 75.525 151.365 75.695 151.555 ;
        RECT 76.445 151.365 76.615 151.555 ;
        RECT 77.825 151.345 77.995 151.535 ;
        RECT 79.665 151.365 79.835 151.555 ;
        RECT 20.645 150.535 22.015 151.345 ;
        RECT 22.395 150.665 31.675 151.345 ;
        RECT 31.915 150.665 35.815 151.345 ;
        RECT 22.395 150.545 24.730 150.665 ;
        RECT 22.395 150.435 23.315 150.545 ;
        RECT 29.395 150.445 30.315 150.665 ;
        RECT 34.885 150.435 35.815 150.665 ;
        RECT 35.825 150.565 37.195 151.345 ;
        RECT 37.215 150.475 37.645 151.260 ;
        RECT 37.665 150.535 39.495 151.345 ;
        RECT 39.505 150.435 42.980 151.345 ;
        RECT 43.185 150.435 46.660 151.345 ;
        RECT 46.865 150.535 48.235 151.345 ;
        RECT 48.245 150.535 51.915 151.345 ;
        RECT 51.925 150.535 57.435 151.345 ;
        RECT 57.445 150.535 62.955 151.345 ;
        RECT 62.975 150.475 63.405 151.260 ;
        RECT 63.885 150.535 66.635 151.345 ;
        RECT 66.655 150.435 68.005 151.345 ;
        RECT 68.485 150.535 70.315 151.345 ;
        RECT 70.325 150.565 71.695 151.345 ;
        RECT 71.705 150.665 73.535 151.345 ;
        RECT 73.545 150.665 75.375 151.345 ;
        RECT 71.705 150.435 73.050 150.665 ;
        RECT 74.030 150.435 75.375 150.665 ;
        RECT 75.385 150.535 78.135 151.345 ;
        RECT 78.145 151.315 79.090 151.345 ;
        RECT 80.580 151.315 80.750 151.535 ;
        RECT 81.050 151.345 81.220 151.535 ;
        RECT 82.420 151.365 82.590 151.585 ;
        RECT 82.745 151.555 86.220 152.465 ;
        RECT 86.435 151.555 87.785 152.465 ;
        RECT 88.175 152.355 89.095 152.465 ;
        RECT 88.175 152.235 90.510 152.355 ;
        RECT 95.175 152.235 96.095 152.455 ;
        RECT 100.665 152.235 101.595 152.465 ;
        RECT 88.175 151.555 97.455 152.235 ;
        RECT 97.695 151.555 101.595 152.235 ;
        RECT 101.615 151.640 102.045 152.425 ;
        RECT 102.075 151.555 103.425 152.465 ;
        RECT 103.445 151.555 104.815 152.335 ;
        RECT 105.480 151.555 108.955 152.465 ;
        RECT 109.160 151.555 112.635 152.465 ;
        RECT 115.845 152.235 116.775 152.465 ;
        RECT 119.985 152.235 120.915 152.465 ;
        RECT 112.875 151.555 116.775 152.235 ;
        RECT 117.015 151.555 120.915 152.235 ;
        RECT 120.925 151.555 122.295 152.335 ;
        RECT 122.305 151.555 123.675 152.335 ;
        RECT 123.685 151.555 126.435 152.365 ;
        RECT 126.445 151.555 127.815 152.365 ;
        RECT 82.890 151.365 83.060 151.555 ;
        RECT 87.485 151.365 87.655 151.555 ;
        RECT 88.130 151.345 88.300 151.535 ;
        RECT 92.730 151.345 92.900 151.535 ;
        RECT 93.465 151.345 93.635 151.535 ;
        RECT 94.845 151.345 95.015 151.535 ;
        RECT 96.280 151.395 96.400 151.505 ;
        RECT 97.145 151.365 97.315 151.555 ;
        RECT 98.065 151.345 98.235 151.535 ;
        RECT 101.010 151.365 101.180 151.555 ;
        RECT 103.125 151.365 103.295 151.555 ;
        RECT 103.585 151.365 103.755 151.555 ;
        RECT 108.640 151.535 108.810 151.555 ;
        RECT 105.020 151.395 105.140 151.505 ;
        RECT 107.265 151.345 107.435 151.535 ;
        RECT 108.640 151.365 108.815 151.535 ;
        RECT 108.645 151.345 108.815 151.365 ;
        RECT 109.110 151.345 109.280 151.535 ;
        RECT 112.320 151.365 112.490 151.555 ;
        RECT 114.165 151.345 114.335 151.535 ;
        RECT 116.190 151.365 116.360 151.555 ;
        RECT 116.465 151.345 116.635 151.535 ;
        RECT 120.330 151.365 120.500 151.555 ;
        RECT 121.065 151.365 121.235 151.555 ;
        RECT 122.445 151.365 122.615 151.555 ;
        RECT 126.125 151.345 126.295 151.555 ;
        RECT 127.505 151.345 127.675 151.555 ;
        RECT 78.145 150.635 80.895 151.315 ;
        RECT 78.145 150.435 79.090 150.635 ;
        RECT 80.905 150.435 84.380 151.345 ;
        RECT 84.815 150.665 88.715 151.345 ;
        RECT 87.785 150.435 88.715 150.665 ;
        RECT 88.735 150.475 89.165 151.260 ;
        RECT 89.415 150.665 93.315 151.345 ;
        RECT 92.385 150.435 93.315 150.665 ;
        RECT 93.325 150.565 94.695 151.345 ;
        RECT 94.705 150.565 96.075 151.345 ;
        RECT 96.545 150.535 98.375 151.345 ;
        RECT 98.385 150.665 107.575 151.345 ;
        RECT 98.385 150.435 99.305 150.665 ;
        RECT 102.135 150.445 103.065 150.665 ;
        RECT 107.585 150.535 108.955 151.345 ;
        RECT 108.965 150.435 112.440 151.345 ;
        RECT 112.645 150.535 114.475 151.345 ;
        RECT 114.495 150.475 114.925 151.260 ;
        RECT 114.945 150.535 116.775 151.345 ;
        RECT 117.155 150.665 126.435 151.345 ;
        RECT 117.155 150.545 119.490 150.665 ;
        RECT 117.155 150.435 118.075 150.545 ;
        RECT 124.155 150.445 125.075 150.665 ;
        RECT 126.445 150.535 127.815 151.345 ;
      LAYER nwell ;
        RECT 20.450 147.315 128.010 150.145 ;
      LAYER pwell ;
        RECT 20.645 146.115 22.015 146.925 ;
        RECT 22.485 146.115 24.315 146.925 ;
        RECT 24.335 146.200 24.765 146.985 ;
        RECT 25.255 146.115 26.605 147.025 ;
        RECT 26.995 146.915 27.915 147.025 ;
        RECT 26.995 146.795 29.330 146.915 ;
        RECT 33.995 146.795 34.915 147.015 ;
        RECT 26.995 146.115 36.275 146.795 ;
        RECT 36.745 146.115 39.495 146.925 ;
        RECT 39.505 146.115 42.980 147.025 ;
        RECT 43.185 146.115 44.555 146.925 ;
        RECT 44.565 146.115 50.075 146.925 ;
        RECT 50.095 146.200 50.525 146.985 ;
        RECT 51.005 146.825 51.950 147.025 ;
        RECT 51.005 146.145 53.755 146.825 ;
        RECT 51.005 146.115 51.950 146.145 ;
        RECT 20.785 145.905 20.955 146.115 ;
        RECT 22.220 145.955 22.340 146.065 ;
        RECT 24.005 145.905 24.175 146.115 ;
        RECT 24.980 145.955 25.100 146.065 ;
        RECT 26.305 145.925 26.475 146.115 ;
        RECT 29.525 145.905 29.695 146.095 ;
        RECT 29.985 145.905 30.155 146.095 ;
        RECT 31.420 145.955 31.540 146.065 ;
        RECT 35.965 145.925 36.135 146.115 ;
        RECT 36.480 145.955 36.600 146.065 ;
        RECT 36.885 145.905 37.055 146.095 ;
        RECT 39.185 145.905 39.355 146.115 ;
        RECT 39.650 145.925 39.820 146.115 ;
        RECT 20.645 145.095 22.015 145.905 ;
        RECT 22.485 145.095 24.315 145.905 ;
        RECT 24.325 145.095 29.835 145.905 ;
        RECT 29.855 144.995 31.205 145.905 ;
        RECT 31.685 145.095 37.195 145.905 ;
        RECT 37.215 145.035 37.645 145.820 ;
        RECT 37.665 145.095 39.495 145.905 ;
        RECT 39.505 145.875 40.450 145.905 ;
        RECT 41.940 145.875 42.110 146.095 ;
        RECT 44.245 145.925 44.415 146.115 ;
        RECT 42.265 145.875 43.210 145.905 ;
        RECT 44.700 145.875 44.870 146.095 ;
        RECT 45.025 145.875 45.970 145.905 ;
        RECT 47.460 145.875 47.630 146.095 ;
        RECT 49.765 145.925 49.935 146.115 ;
        RECT 47.785 145.875 48.730 145.905 ;
        RECT 50.220 145.875 50.390 146.095 ;
        RECT 50.690 145.905 50.860 146.095 ;
        RECT 53.440 145.925 53.610 146.145 ;
        RECT 53.765 146.115 57.240 147.025 ;
        RECT 57.445 146.115 60.920 147.025 ;
        RECT 61.135 146.115 62.485 147.025 ;
        RECT 62.505 146.115 65.255 146.925 ;
        RECT 65.265 146.795 66.185 147.025 ;
        RECT 69.015 146.795 69.945 147.015 ;
        RECT 65.265 146.115 74.455 146.795 ;
        RECT 74.465 146.115 75.835 146.925 ;
        RECT 75.855 146.200 76.285 146.985 ;
        RECT 76.305 146.115 77.675 146.925 ;
        RECT 77.685 146.115 81.355 146.925 ;
        RECT 83.170 146.825 84.115 147.025 ;
        RECT 81.365 146.145 84.115 146.825 ;
        RECT 53.910 145.925 54.080 146.115 ;
        RECT 54.370 145.905 54.540 146.095 ;
        RECT 57.590 145.925 57.760 146.115 ;
        RECT 58.505 145.950 58.665 146.060 ;
        RECT 62.185 145.925 62.355 146.115 ;
        RECT 62.370 145.905 62.540 146.095 ;
        RECT 64.025 145.950 64.185 146.060 ;
        RECT 64.490 145.905 64.660 146.095 ;
        RECT 64.945 145.925 65.115 146.115 ;
        RECT 71.570 145.905 71.740 146.095 ;
        RECT 73.225 145.905 73.395 146.095 ;
        RECT 74.145 145.925 74.315 146.115 ;
        RECT 74.605 145.905 74.775 146.095 ;
        RECT 75.525 145.925 75.695 146.115 ;
        RECT 77.365 145.925 77.535 146.115 ;
        RECT 78.285 145.905 78.455 146.095 ;
        RECT 81.045 145.925 81.215 146.115 ;
        RECT 81.510 145.925 81.680 146.145 ;
        RECT 83.170 146.115 84.115 146.145 ;
        RECT 85.045 146.115 90.555 146.925 ;
        RECT 90.565 146.115 96.075 146.925 ;
        RECT 96.085 146.115 101.595 146.925 ;
        RECT 101.615 146.200 102.045 146.985 ;
        RECT 102.065 146.115 105.735 146.925 ;
        RECT 105.745 146.825 106.690 147.025 ;
        RECT 108.505 146.825 109.450 147.025 ;
        RECT 105.745 146.145 108.495 146.825 ;
        RECT 108.505 146.145 111.255 146.825 ;
        RECT 105.745 146.115 106.690 146.145 ;
        RECT 81.960 145.905 82.130 146.095 ;
        RECT 82.430 145.905 82.600 146.095 ;
        RECT 84.725 145.960 84.885 146.070 ;
        RECT 88.405 145.905 88.575 146.095 ;
        RECT 89.785 145.950 89.945 146.060 ;
        RECT 90.245 145.925 90.415 146.115 ;
        RECT 93.465 145.905 93.635 146.095 ;
        RECT 95.765 145.925 95.935 146.115 ;
        RECT 98.985 145.905 99.155 146.095 ;
        RECT 101.285 145.925 101.455 146.115 ;
        RECT 104.505 145.905 104.675 146.095 ;
        RECT 105.425 145.925 105.595 146.115 ;
        RECT 108.180 145.925 108.350 146.145 ;
        RECT 108.505 146.115 109.450 146.145 ;
        RECT 110.025 145.905 110.195 146.095 ;
        RECT 39.505 145.195 42.255 145.875 ;
        RECT 42.265 145.195 45.015 145.875 ;
        RECT 45.025 145.195 47.775 145.875 ;
        RECT 47.785 145.195 50.535 145.875 ;
        RECT 39.505 144.995 40.450 145.195 ;
        RECT 42.265 144.995 43.210 145.195 ;
        RECT 45.025 144.995 45.970 145.195 ;
        RECT 47.785 144.995 48.730 145.195 ;
        RECT 50.545 144.995 54.020 145.905 ;
        RECT 54.225 144.995 57.700 145.905 ;
        RECT 59.055 145.225 62.955 145.905 ;
        RECT 62.025 144.995 62.955 145.225 ;
        RECT 62.975 145.035 63.405 145.820 ;
        RECT 64.345 144.995 67.820 145.905 ;
        RECT 68.255 145.225 72.155 145.905 ;
        RECT 71.225 144.995 72.155 145.225 ;
        RECT 72.175 144.995 73.525 145.905 ;
        RECT 73.545 145.095 74.915 145.905 ;
        RECT 74.925 145.095 78.595 145.905 ;
        RECT 78.800 144.995 82.275 145.905 ;
        RECT 82.285 144.995 85.760 145.905 ;
        RECT 85.965 145.095 88.715 145.905 ;
        RECT 88.735 145.035 89.165 145.820 ;
        RECT 90.105 145.095 93.775 145.905 ;
        RECT 93.785 145.095 99.295 145.905 ;
        RECT 99.305 145.095 104.815 145.905 ;
        RECT 104.825 145.095 110.335 145.905 ;
        RECT 110.490 145.875 110.660 146.095 ;
        RECT 110.940 145.925 111.110 146.145 ;
        RECT 111.265 146.115 114.740 147.025 ;
        RECT 114.945 146.115 116.315 146.925 ;
        RECT 116.325 146.115 119.995 146.925 ;
        RECT 120.015 146.115 121.365 147.025 ;
        RECT 121.385 146.115 122.755 146.925 ;
        RECT 122.765 146.115 126.435 146.925 ;
        RECT 126.445 146.115 127.815 146.925 ;
        RECT 111.410 145.925 111.580 146.115 ;
        RECT 114.165 145.905 114.335 146.095 ;
        RECT 116.005 145.925 116.175 146.115 ;
        RECT 117.385 145.905 117.555 146.095 ;
        RECT 117.845 145.905 118.015 146.095 ;
        RECT 119.280 145.955 119.400 146.065 ;
        RECT 119.685 145.905 119.855 146.115 ;
        RECT 120.145 145.925 120.315 146.115 ;
        RECT 122.445 145.925 122.615 146.115 ;
        RECT 126.125 145.905 126.295 146.115 ;
        RECT 127.505 145.905 127.675 146.115 ;
        RECT 112.150 145.875 113.095 145.905 ;
        RECT 110.345 145.195 113.095 145.875 ;
        RECT 112.150 144.995 113.095 145.195 ;
        RECT 113.105 145.095 114.475 145.905 ;
        RECT 114.495 145.035 114.925 145.820 ;
        RECT 114.945 145.095 117.695 145.905 ;
        RECT 117.715 144.995 119.065 145.905 ;
        RECT 119.555 144.995 120.905 145.905 ;
        RECT 120.925 145.095 126.435 145.905 ;
        RECT 126.445 145.095 127.815 145.905 ;
      LAYER nwell ;
        RECT 20.450 141.875 128.010 144.705 ;
      LAYER pwell ;
        RECT 20.645 140.675 22.015 141.485 ;
        RECT 22.485 140.675 24.315 141.485 ;
        RECT 24.335 140.760 24.765 141.545 ;
        RECT 25.245 140.675 30.755 141.485 ;
        RECT 30.765 140.675 36.275 141.485 ;
        RECT 36.285 140.675 41.795 141.485 ;
        RECT 41.805 141.385 42.750 141.585 ;
        RECT 45.705 141.495 46.655 141.585 ;
        RECT 41.805 140.705 44.555 141.385 ;
        RECT 41.805 140.675 42.750 140.705 ;
        RECT 20.785 140.465 20.955 140.675 ;
        RECT 22.220 140.515 22.340 140.625 ;
        RECT 22.625 140.510 22.785 140.620 ;
        RECT 24.005 140.485 24.175 140.675 ;
        RECT 24.980 140.515 25.100 140.625 ;
        RECT 30.445 140.485 30.615 140.675 ;
        RECT 32.285 140.465 32.455 140.655 ;
        RECT 33.665 140.465 33.835 140.655 ;
        RECT 35.045 140.465 35.215 140.655 ;
        RECT 35.505 140.465 35.675 140.655 ;
        RECT 35.965 140.485 36.135 140.675 ;
        RECT 36.940 140.515 37.060 140.625 ;
        RECT 37.860 140.515 37.980 140.625 ;
        RECT 40.565 140.465 40.735 140.655 ;
        RECT 41.485 140.485 41.655 140.675 ;
        RECT 41.945 140.465 42.115 140.655 ;
        RECT 42.405 140.485 42.575 140.655 ;
        RECT 44.240 140.485 44.410 140.705 ;
        RECT 44.725 140.675 46.655 141.495 ;
        RECT 47.325 140.675 50.075 141.485 ;
        RECT 50.095 140.760 50.525 141.545 ;
        RECT 50.545 140.675 56.055 141.485 ;
        RECT 56.435 141.475 57.355 141.585 ;
        RECT 56.435 141.355 58.770 141.475 ;
        RECT 63.435 141.355 64.355 141.575 ;
        RECT 66.555 141.475 67.475 141.585 ;
        RECT 66.555 141.355 68.890 141.475 ;
        RECT 73.555 141.355 74.475 141.575 ;
        RECT 56.435 140.675 65.715 141.355 ;
        RECT 66.555 140.675 75.835 141.355 ;
        RECT 75.855 140.760 76.285 141.545 ;
        RECT 76.765 140.675 79.515 141.485 ;
        RECT 79.525 141.385 80.470 141.585 ;
        RECT 79.525 140.705 82.275 141.385 ;
        RECT 85.485 141.355 86.415 141.585 ;
        RECT 79.525 140.675 80.470 140.705 ;
        RECT 44.725 140.655 44.875 140.675 ;
        RECT 44.705 140.485 44.875 140.655 ;
        RECT 47.060 140.515 47.180 140.625 ;
        RECT 42.425 140.465 42.575 140.485 ;
        RECT 44.725 140.465 44.875 140.485 ;
        RECT 49.305 140.465 49.475 140.655 ;
        RECT 49.765 140.485 49.935 140.675 ;
        RECT 51.605 140.485 51.775 140.655 ;
        RECT 53.905 140.485 54.075 140.655 ;
        RECT 51.605 140.465 51.755 140.485 ;
        RECT 53.905 140.465 54.055 140.485 ;
        RECT 55.745 140.465 55.915 140.675 ;
        RECT 61.265 140.465 61.435 140.655 ;
        RECT 61.725 140.465 61.895 140.655 ;
        RECT 65.405 140.485 65.575 140.675 ;
        RECT 65.865 140.625 66.035 140.655 ;
        RECT 65.865 140.515 66.040 140.625 ;
        RECT 65.865 140.465 66.035 140.515 ;
        RECT 66.330 140.465 66.500 140.655 ;
        RECT 70.005 140.465 70.175 140.655 ;
        RECT 73.280 140.515 73.400 140.625 ;
        RECT 75.065 140.465 75.235 140.655 ;
        RECT 75.525 140.485 75.695 140.675 ;
        RECT 76.500 140.515 76.620 140.625 ;
        RECT 79.205 140.485 79.375 140.675 ;
        RECT 80.585 140.465 80.755 140.655 ;
        RECT 81.045 140.485 81.215 140.655 ;
        RECT 81.960 140.485 82.130 140.705 ;
        RECT 82.515 140.675 86.415 141.355 ;
        RECT 86.795 141.475 87.715 141.585 ;
        RECT 86.795 141.355 89.130 141.475 ;
        RECT 93.795 141.355 94.715 141.575 ;
        RECT 86.795 140.675 96.075 141.355 ;
        RECT 96.545 140.675 97.915 141.455 ;
        RECT 98.120 140.675 101.595 141.585 ;
        RECT 101.615 140.760 102.045 141.545 ;
        RECT 102.075 140.675 103.425 141.585 ;
        RECT 107.105 141.355 108.035 141.585 ;
        RECT 104.135 140.675 108.035 141.355 ;
        RECT 109.160 140.675 112.635 141.585 ;
        RECT 115.845 141.355 116.775 141.585 ;
        RECT 112.875 140.675 116.775 141.355 ;
        RECT 117.155 141.475 118.075 141.585 ;
        RECT 117.155 141.355 119.490 141.475 ;
        RECT 124.155 141.355 125.075 141.575 ;
        RECT 117.155 140.675 126.435 141.355 ;
        RECT 126.445 140.675 127.815 141.485 ;
        RECT 83.400 140.515 83.520 140.625 ;
        RECT 85.830 140.485 86.000 140.675 ;
        RECT 81.065 140.465 81.215 140.485 ;
        RECT 87.025 140.465 87.195 140.655 ;
        RECT 87.485 140.465 87.655 140.655 ;
        RECT 89.380 140.515 89.500 140.625 ;
        RECT 95.765 140.485 95.935 140.675 ;
        RECT 96.280 140.515 96.400 140.625 ;
        RECT 97.605 140.485 97.775 140.675 ;
        RECT 98.985 140.465 99.155 140.655 ;
        RECT 101.280 140.485 101.450 140.675 ;
        RECT 102.205 140.485 102.375 140.675 ;
        RECT 103.640 140.515 103.760 140.625 ;
        RECT 107.450 140.485 107.620 140.675 ;
        RECT 108.645 140.465 108.815 140.655 ;
        RECT 110.025 140.465 110.195 140.655 ;
        RECT 112.320 140.485 112.490 140.675 ;
        RECT 113.890 140.465 114.060 140.655 ;
        RECT 116.190 140.485 116.360 140.675 ;
        RECT 124.285 140.465 124.455 140.655 ;
        RECT 126.125 140.465 126.295 140.675 ;
        RECT 127.505 140.465 127.675 140.675 ;
        RECT 20.645 139.655 22.015 140.465 ;
        RECT 23.315 139.785 32.595 140.465 ;
        RECT 23.315 139.665 25.650 139.785 ;
        RECT 23.315 139.555 24.235 139.665 ;
        RECT 30.315 139.565 31.235 139.785 ;
        RECT 32.605 139.685 33.975 140.465 ;
        RECT 33.985 139.655 35.355 140.465 ;
        RECT 35.375 139.555 36.725 140.465 ;
        RECT 37.215 139.595 37.645 140.380 ;
        RECT 38.125 139.655 40.875 140.465 ;
        RECT 40.885 139.685 42.255 140.465 ;
        RECT 42.425 139.645 44.355 140.465 ;
        RECT 44.725 139.645 46.655 140.465 ;
        RECT 46.865 139.655 49.615 140.465 ;
        RECT 43.405 139.555 44.355 139.645 ;
        RECT 45.705 139.555 46.655 139.645 ;
        RECT 49.825 139.645 51.755 140.465 ;
        RECT 52.125 139.645 54.055 140.465 ;
        RECT 54.225 139.655 56.055 140.465 ;
        RECT 56.065 139.655 61.575 140.465 ;
        RECT 61.585 139.685 62.955 140.465 ;
        RECT 49.825 139.555 50.775 139.645 ;
        RECT 52.125 139.555 53.075 139.645 ;
        RECT 62.975 139.595 63.405 140.380 ;
        RECT 63.425 139.655 66.175 140.465 ;
        RECT 66.185 139.555 69.660 140.465 ;
        RECT 69.865 139.555 73.075 140.465 ;
        RECT 73.545 139.655 75.375 140.465 ;
        RECT 75.385 139.655 80.895 140.465 ;
        RECT 81.065 139.645 82.995 140.465 ;
        RECT 83.665 139.655 87.335 140.465 ;
        RECT 82.045 139.555 82.995 139.645 ;
        RECT 87.355 139.555 88.705 140.465 ;
        RECT 88.735 139.595 89.165 140.380 ;
        RECT 90.015 139.785 99.295 140.465 ;
        RECT 99.675 139.785 108.955 140.465 ;
        RECT 90.015 139.665 92.350 139.785 ;
        RECT 90.015 139.555 90.935 139.665 ;
        RECT 97.015 139.565 97.935 139.785 ;
        RECT 99.675 139.665 102.010 139.785 ;
        RECT 99.675 139.555 100.595 139.665 ;
        RECT 106.675 139.565 107.595 139.785 ;
        RECT 108.965 139.685 110.335 140.465 ;
        RECT 110.575 139.785 114.475 140.465 ;
        RECT 113.545 139.555 114.475 139.785 ;
        RECT 114.495 139.595 114.925 140.380 ;
        RECT 115.315 139.785 124.595 140.465 ;
        RECT 115.315 139.665 117.650 139.785 ;
        RECT 115.315 139.555 116.235 139.665 ;
        RECT 122.315 139.565 123.235 139.785 ;
        RECT 124.605 139.655 126.435 140.465 ;
        RECT 126.445 139.655 127.815 140.465 ;
      LAYER nwell ;
        RECT 20.450 136.435 128.010 139.265 ;
      LAYER pwell ;
        RECT 20.645 135.235 22.015 136.045 ;
        RECT 22.485 135.235 24.315 136.045 ;
        RECT 24.335 135.320 24.765 136.105 ;
        RECT 24.785 135.235 26.615 136.045 ;
        RECT 26.635 135.235 27.985 136.145 ;
        RECT 31.205 135.915 32.135 136.145 ;
        RECT 28.235 135.235 32.135 135.915 ;
        RECT 32.515 136.035 33.435 136.145 ;
        RECT 32.515 135.915 34.850 136.035 ;
        RECT 39.515 135.915 40.435 136.135 ;
        RECT 41.805 135.915 42.735 136.145 ;
        RECT 32.515 135.235 41.795 135.915 ;
        RECT 41.805 135.235 45.705 135.915 ;
        RECT 46.405 135.235 48.235 136.045 ;
        RECT 48.255 135.235 49.605 136.145 ;
        RECT 50.095 135.320 50.525 136.105 ;
        RECT 52.585 136.055 53.535 136.145 ;
        RECT 51.005 135.235 52.375 136.015 ;
        RECT 52.585 135.235 54.515 136.055 ;
        RECT 55.155 135.235 57.895 135.915 ;
        RECT 58.825 135.235 64.335 136.045 ;
        RECT 64.345 135.235 67.820 136.145 ;
        RECT 68.945 135.235 72.615 136.045 ;
        RECT 72.625 135.235 74.455 135.915 ;
        RECT 74.465 135.235 75.835 136.045 ;
        RECT 75.855 135.320 76.285 136.105 ;
        RECT 79.285 136.055 80.235 136.145 ;
        RECT 76.305 135.235 78.135 136.045 ;
        RECT 78.305 135.235 80.235 136.055 ;
        RECT 80.645 136.055 81.595 136.145 ;
        RECT 82.945 136.055 83.895 136.145 ;
        RECT 80.645 135.235 82.575 136.055 ;
        RECT 82.945 135.235 84.875 136.055 ;
        RECT 85.045 135.235 86.415 136.015 ;
        RECT 86.885 135.235 90.555 136.045 ;
        RECT 90.575 135.235 91.925 136.145 ;
        RECT 91.945 135.235 93.315 136.015 ;
        RECT 97.445 135.915 98.375 136.145 ;
        RECT 94.475 135.235 98.375 135.915 ;
        RECT 98.385 135.945 99.330 136.145 ;
        RECT 98.385 135.265 101.135 135.945 ;
        RECT 101.615 135.320 102.045 136.105 ;
        RECT 98.385 135.235 99.330 135.265 ;
        RECT 20.785 135.025 20.955 135.235 ;
        RECT 22.220 135.075 22.340 135.185 ;
        RECT 24.005 135.045 24.175 135.235 ;
        RECT 26.305 135.045 26.475 135.235 ;
        RECT 27.685 135.045 27.855 135.235 ;
        RECT 31.365 135.025 31.535 135.215 ;
        RECT 31.550 135.045 31.720 135.235 ;
        RECT 32.745 135.025 32.915 135.215 ;
        RECT 34.125 135.025 34.295 135.215 ;
        RECT 20.645 134.215 22.015 135.025 ;
        RECT 22.395 134.345 31.675 135.025 ;
        RECT 22.395 134.225 24.730 134.345 ;
        RECT 22.395 134.115 23.315 134.225 ;
        RECT 29.395 134.125 30.315 134.345 ;
        RECT 31.685 134.245 33.055 135.025 ;
        RECT 33.065 134.215 34.435 135.025 ;
        RECT 34.445 134.995 35.390 135.025 ;
        RECT 36.880 134.995 37.050 135.215 ;
        RECT 39.185 135.045 39.355 135.215 ;
        RECT 41.485 135.045 41.655 135.235 ;
        RECT 34.445 134.315 37.195 134.995 ;
        RECT 34.445 134.115 35.390 134.315 ;
        RECT 37.215 134.155 37.645 134.940 ;
        RECT 37.665 134.345 39.030 135.025 ;
        RECT 39.505 134.995 40.450 135.025 ;
        RECT 41.940 134.995 42.110 135.215 ;
        RECT 42.220 135.045 42.390 135.235 ;
        RECT 42.865 135.070 43.025 135.180 ;
        RECT 43.325 135.025 43.495 135.215 ;
        RECT 46.140 135.075 46.260 135.185 ;
        RECT 47.925 135.045 48.095 135.235 ;
        RECT 49.305 135.045 49.475 135.235 ;
        RECT 49.820 135.075 49.940 135.185 ;
        RECT 50.740 135.075 50.860 135.185 ;
        RECT 52.065 135.045 52.235 135.235 ;
        RECT 54.365 135.215 54.515 135.235 ;
        RECT 52.800 135.025 52.970 135.215 ;
        RECT 54.365 135.045 54.535 135.215 ;
        RECT 54.880 135.075 55.000 135.185 ;
        RECT 57.585 135.025 57.755 135.235 ;
        RECT 58.505 135.070 58.665 135.190 ;
        RECT 62.370 135.025 62.540 135.215 ;
        RECT 64.025 135.045 64.195 135.235 ;
        RECT 64.490 135.215 64.660 135.235 ;
        RECT 64.485 135.045 64.660 135.215 ;
        RECT 64.485 135.025 64.655 135.045 ;
        RECT 64.950 135.025 65.120 135.215 ;
        RECT 68.625 135.080 68.785 135.190 ;
        RECT 70.925 135.025 71.095 135.215 ;
        RECT 72.305 135.045 72.475 135.235 ;
        RECT 72.765 135.025 72.935 135.215 ;
        RECT 74.145 135.045 74.315 135.235 ;
        RECT 75.065 135.045 75.235 135.215 ;
        RECT 75.525 135.185 75.695 135.235 ;
        RECT 75.525 135.075 75.700 135.185 ;
        RECT 75.525 135.045 75.695 135.075 ;
        RECT 77.825 135.045 77.995 135.235 ;
        RECT 78.305 135.215 78.455 135.235 ;
        RECT 75.065 135.025 75.215 135.045 ;
        RECT 78.285 135.025 78.455 135.215 ;
        RECT 82.425 135.215 82.575 135.235 ;
        RECT 84.725 135.215 84.875 135.235 ;
        RECT 82.425 135.045 82.595 135.215 ;
        RECT 84.725 135.045 84.895 135.215 ;
        RECT 85.185 135.045 85.355 135.235 ;
        RECT 86.620 135.075 86.740 135.185 ;
        RECT 87.945 135.025 88.115 135.215 ;
        RECT 88.460 135.075 88.580 135.185 ;
        RECT 89.785 135.070 89.945 135.180 ;
        RECT 90.245 135.045 90.415 135.235 ;
        RECT 90.705 135.045 90.875 135.235 ;
        RECT 92.085 135.045 92.255 135.235 ;
        RECT 93.925 135.080 94.085 135.190 ;
        RECT 95.305 135.025 95.475 135.215 ;
        RECT 97.790 135.045 97.960 135.235 ;
        RECT 100.820 135.215 100.990 135.265 ;
        RECT 102.065 135.235 104.815 136.045 ;
        RECT 104.825 135.945 105.770 136.145 ;
        RECT 104.825 135.265 107.575 135.945 ;
        RECT 104.825 135.235 105.770 135.265 ;
        RECT 100.820 135.045 100.995 135.215 ;
        RECT 101.340 135.075 101.460 135.185 ;
        RECT 104.505 135.045 104.675 135.235 ;
        RECT 100.825 135.025 100.995 135.045 ;
        RECT 106.345 135.025 106.515 135.215 ;
        RECT 106.805 135.045 106.975 135.215 ;
        RECT 107.260 135.045 107.430 135.265 ;
        RECT 107.585 135.235 111.060 136.145 ;
        RECT 111.265 135.945 112.210 136.145 ;
        RECT 111.265 135.265 114.015 135.945 ;
        RECT 111.265 135.235 112.210 135.265 ;
        RECT 107.730 135.045 107.900 135.235 ;
        RECT 113.700 135.215 113.870 135.265 ;
        RECT 114.025 135.235 119.535 136.045 ;
        RECT 119.545 135.235 120.915 136.015 ;
        RECT 121.845 135.235 123.215 136.015 ;
        RECT 123.685 135.235 126.435 136.045 ;
        RECT 126.445 135.235 127.815 136.045 ;
        RECT 110.945 135.045 111.115 135.215 ;
        RECT 111.460 135.075 111.580 135.185 ;
        RECT 113.700 135.045 113.875 135.215 ;
        RECT 114.220 135.075 114.340 135.185 ;
        RECT 115.140 135.075 115.260 135.185 ;
        RECT 119.225 135.045 119.395 135.235 ;
        RECT 119.685 135.045 119.855 135.235 ;
        RECT 106.825 135.025 106.975 135.045 ;
        RECT 110.945 135.025 111.095 135.045 ;
        RECT 113.705 135.025 113.855 135.045 ;
        RECT 120.605 135.025 120.775 135.215 ;
        RECT 121.525 135.080 121.685 135.190 ;
        RECT 121.985 135.045 122.155 135.235 ;
        RECT 123.420 135.075 123.540 135.185 ;
        RECT 126.125 135.025 126.295 135.235 ;
        RECT 127.505 135.025 127.675 135.235 ;
        RECT 39.505 134.315 42.255 134.995 ;
        RECT 43.185 134.345 52.290 135.025 ;
        RECT 52.385 134.345 56.285 135.025 ;
        RECT 39.505 134.115 40.450 134.315 ;
        RECT 52.385 134.115 53.315 134.345 ;
        RECT 56.525 134.245 57.895 135.025 ;
        RECT 59.055 134.345 62.955 135.025 ;
        RECT 62.025 134.115 62.955 134.345 ;
        RECT 62.975 134.155 63.405 134.940 ;
        RECT 63.425 134.215 64.795 135.025 ;
        RECT 64.805 134.115 68.280 135.025 ;
        RECT 68.485 134.215 71.235 135.025 ;
        RECT 71.245 134.345 73.075 135.025 ;
        RECT 73.285 134.205 75.215 135.025 ;
        RECT 75.845 134.215 78.595 135.025 ;
        RECT 78.975 134.345 88.255 135.025 ;
        RECT 78.975 134.225 81.310 134.345 ;
        RECT 73.285 134.115 74.235 134.205 ;
        RECT 78.975 134.115 79.895 134.225 ;
        RECT 85.975 134.125 86.895 134.345 ;
        RECT 88.735 134.155 89.165 134.940 ;
        RECT 90.105 134.215 95.615 135.025 ;
        RECT 95.625 134.215 101.135 135.025 ;
        RECT 101.145 134.215 106.655 135.025 ;
        RECT 106.825 134.205 108.755 135.025 ;
        RECT 107.805 134.115 108.755 134.205 ;
        RECT 109.165 134.205 111.095 135.025 ;
        RECT 111.925 134.205 113.855 135.025 ;
        RECT 109.165 134.115 110.115 134.205 ;
        RECT 111.925 134.115 112.875 134.205 ;
        RECT 114.495 134.155 114.925 134.940 ;
        RECT 115.405 134.215 120.915 135.025 ;
        RECT 120.925 134.215 126.435 135.025 ;
        RECT 126.445 134.215 127.815 135.025 ;
      LAYER nwell ;
        RECT 20.450 130.995 128.010 133.825 ;
      LAYER pwell ;
        RECT 20.645 129.795 22.015 130.605 ;
        RECT 22.485 129.795 24.315 130.605 ;
        RECT 24.335 129.880 24.765 130.665 ;
        RECT 25.715 129.795 27.065 130.705 ;
        RECT 30.285 130.475 31.215 130.705 ;
        RECT 40.795 130.595 41.715 130.705 ;
        RECT 40.795 130.475 43.130 130.595 ;
        RECT 47.795 130.475 48.715 130.695 ;
        RECT 27.315 129.795 31.215 130.475 ;
        RECT 31.310 129.795 40.415 130.475 ;
        RECT 40.795 129.795 50.075 130.475 ;
        RECT 50.095 129.880 50.525 130.665 ;
        RECT 51.015 129.795 52.365 130.705 ;
        RECT 55.585 130.475 56.515 130.705 ;
        RECT 52.615 129.795 56.515 130.475 ;
        RECT 56.905 129.795 59.330 130.475 ;
        RECT 59.745 129.795 63.415 130.605 ;
        RECT 63.425 129.795 64.795 130.575 ;
        RECT 65.265 129.795 68.015 130.605 ;
        RECT 71.225 130.475 72.155 130.705 ;
        RECT 68.255 129.795 72.155 130.475 ;
        RECT 73.085 129.795 75.825 130.475 ;
        RECT 75.855 129.880 76.285 130.665 ;
        RECT 76.315 129.795 77.665 130.705 ;
        RECT 77.685 130.475 78.615 130.705 ;
        RECT 85.025 130.475 85.955 130.705 ;
        RECT 77.685 129.795 81.585 130.475 ;
        RECT 82.055 129.795 85.955 130.475 ;
        RECT 85.965 129.795 87.795 130.605 ;
        RECT 87.805 129.795 93.315 130.605 ;
        RECT 93.335 129.795 94.685 130.705 ;
        RECT 97.905 130.475 98.835 130.705 ;
        RECT 94.935 129.795 98.835 130.475 ;
        RECT 98.845 129.795 100.215 130.575 ;
        RECT 100.225 129.795 101.595 130.605 ;
        RECT 101.615 129.880 102.045 130.665 ;
        RECT 106.405 130.615 107.355 130.705 ;
        RECT 102.065 129.795 103.435 130.605 ;
        RECT 103.455 129.795 106.195 130.475 ;
        RECT 106.405 129.795 108.335 130.615 ;
        RECT 108.505 129.795 110.335 130.605 ;
        RECT 113.545 130.475 114.475 130.705 ;
        RECT 110.575 129.795 114.475 130.475 ;
        RECT 114.485 129.795 118.155 130.605 ;
        RECT 118.175 129.795 119.525 130.705 ;
        RECT 120.465 129.795 121.835 130.575 ;
        RECT 122.765 129.795 126.435 130.605 ;
        RECT 126.445 129.795 127.815 130.605 ;
        RECT 20.785 129.585 20.955 129.795 ;
        RECT 22.220 129.635 22.340 129.745 ;
        RECT 24.005 129.605 24.175 129.795 ;
        RECT 25.385 129.640 25.545 129.750 ;
        RECT 26.765 129.605 26.935 129.795 ;
        RECT 27.685 129.585 27.855 129.775 ;
        RECT 30.630 129.605 30.800 129.795 ;
        RECT 31.550 129.585 31.720 129.775 ;
        RECT 32.340 129.635 32.460 129.745 ;
        RECT 32.745 129.605 32.915 129.775 ;
        RECT 35.045 129.605 35.215 129.775 ;
        RECT 37.860 129.635 37.980 129.745 ;
        RECT 32.765 129.585 32.915 129.605 ;
        RECT 35.065 129.585 35.215 129.605 ;
        RECT 40.105 129.605 40.275 129.795 ;
        RECT 41.025 129.630 41.185 129.740 ;
        RECT 41.485 129.605 41.655 129.775 ;
        RECT 49.765 129.605 49.935 129.795 ;
        RECT 50.740 129.635 50.860 129.745 ;
        RECT 52.065 129.605 52.235 129.795 ;
        RECT 40.105 129.585 40.255 129.605 ;
        RECT 20.645 128.775 22.015 129.585 ;
        RECT 22.485 128.775 27.995 129.585 ;
        RECT 28.235 128.905 32.135 129.585 ;
        RECT 31.205 128.675 32.135 128.905 ;
        RECT 32.765 128.765 34.695 129.585 ;
        RECT 35.065 128.765 36.995 129.585 ;
        RECT 33.745 128.675 34.695 128.765 ;
        RECT 36.045 128.675 36.995 128.765 ;
        RECT 37.215 128.715 37.645 129.500 ;
        RECT 38.325 128.765 40.255 129.585 ;
        RECT 41.505 129.585 41.655 129.605 ;
        RECT 52.985 129.585 53.155 129.775 ;
        RECT 55.930 129.605 56.100 129.795 ;
        RECT 59.425 129.605 59.595 129.775 ;
        RECT 62.645 129.585 62.815 129.775 ;
        RECT 63.105 129.605 63.275 129.795 ;
        RECT 64.485 129.585 64.655 129.795 ;
        RECT 65.000 129.635 65.120 129.745 ;
        RECT 66.785 129.585 66.955 129.775 ;
        RECT 67.705 129.605 67.875 129.795 ;
        RECT 71.570 129.605 71.740 129.795 ;
        RECT 72.765 129.640 72.925 129.750 ;
        RECT 73.225 129.605 73.395 129.795 ;
        RECT 76.445 129.585 76.615 129.795 ;
        RECT 78.100 129.605 78.270 129.795 ;
        RECT 79.205 129.585 79.375 129.775 ;
        RECT 79.665 129.585 79.835 129.775 ;
        RECT 85.370 129.605 85.540 129.795 ;
        RECT 87.485 129.605 87.655 129.795 ;
        RECT 89.380 129.635 89.500 129.745 ;
        RECT 92.085 129.585 92.255 129.775 ;
        RECT 92.545 129.585 92.715 129.775 ;
        RECT 93.005 129.605 93.175 129.795 ;
        RECT 93.465 129.605 93.635 129.795 ;
        RECT 98.250 129.605 98.420 129.795 ;
        RECT 99.905 129.605 100.075 129.795 ;
        RECT 101.285 129.605 101.455 129.795 ;
        RECT 102.205 129.585 102.375 129.775 ;
        RECT 103.125 129.605 103.295 129.795 ;
        RECT 105.885 129.605 106.055 129.795 ;
        RECT 108.185 129.775 108.335 129.795 ;
        RECT 108.185 129.605 108.355 129.775 ;
        RECT 110.025 129.605 110.195 129.795 ;
        RECT 111.405 129.605 111.575 129.775 ;
        RECT 113.890 129.605 114.060 129.795 ;
        RECT 114.165 129.630 114.325 129.740 ;
        RECT 115.140 129.635 115.260 129.745 ;
        RECT 117.845 129.605 118.015 129.795 ;
        RECT 118.305 129.605 118.475 129.795 ;
        RECT 120.145 129.640 120.305 129.750 ;
        RECT 120.605 129.605 120.775 129.795 ;
        RECT 122.445 129.640 122.605 129.750 ;
        RECT 111.425 129.585 111.575 129.605 ;
        RECT 124.745 129.585 124.915 129.775 ;
        RECT 126.125 129.585 126.295 129.795 ;
        RECT 127.505 129.585 127.675 129.795 ;
        RECT 41.505 128.765 43.435 129.585 ;
        RECT 38.325 128.675 39.275 128.765 ;
        RECT 42.485 128.675 43.435 128.765 ;
        RECT 44.015 128.905 53.295 129.585 ;
        RECT 53.675 128.905 62.955 129.585 ;
        RECT 44.015 128.785 46.350 128.905 ;
        RECT 44.015 128.675 44.935 128.785 ;
        RECT 51.015 128.685 51.935 128.905 ;
        RECT 53.675 128.785 56.010 128.905 ;
        RECT 53.675 128.675 54.595 128.785 ;
        RECT 60.675 128.685 61.595 128.905 ;
        RECT 62.975 128.715 63.405 129.500 ;
        RECT 63.435 128.675 64.785 129.585 ;
        RECT 65.265 128.775 67.095 129.585 ;
        RECT 67.475 128.905 76.755 129.585 ;
        RECT 67.475 128.785 69.810 128.905 ;
        RECT 67.475 128.675 68.395 128.785 ;
        RECT 74.475 128.685 75.395 128.905 ;
        RECT 76.765 128.775 79.515 129.585 ;
        RECT 79.525 128.905 88.630 129.585 ;
        RECT 88.735 128.715 89.165 129.500 ;
        RECT 89.645 128.775 92.395 129.585 ;
        RECT 92.405 128.905 101.685 129.585 ;
        RECT 102.065 128.905 111.170 129.585 ;
        RECT 93.765 128.685 94.685 128.905 ;
        RECT 99.350 128.785 101.685 128.905 ;
        RECT 100.765 128.675 101.685 128.785 ;
        RECT 111.425 128.765 113.355 129.585 ;
        RECT 112.405 128.675 113.355 128.765 ;
        RECT 114.495 128.715 114.925 129.500 ;
        RECT 115.775 128.905 125.055 129.585 ;
        RECT 115.775 128.785 118.110 128.905 ;
        RECT 115.775 128.675 116.695 128.785 ;
        RECT 122.775 128.685 123.695 128.905 ;
        RECT 125.065 128.775 126.435 129.585 ;
        RECT 126.445 128.775 127.815 129.585 ;
      LAYER nwell ;
        RECT 20.450 125.555 128.010 128.385 ;
      LAYER pwell ;
        RECT 20.645 124.355 22.015 125.165 ;
        RECT 22.955 124.355 24.305 125.265 ;
        RECT 24.335 124.440 24.765 125.225 ;
        RECT 24.795 124.355 26.145 125.265 ;
        RECT 26.165 124.355 27.535 125.135 ;
        RECT 27.545 125.035 28.475 125.265 ;
        RECT 32.975 125.155 33.895 125.265 ;
        RECT 32.975 125.035 35.310 125.155 ;
        RECT 39.975 125.035 40.895 125.255 ;
        RECT 45.925 125.035 46.855 125.265 ;
        RECT 27.545 124.355 31.445 125.035 ;
        RECT 32.975 124.355 42.255 125.035 ;
        RECT 42.955 124.355 46.855 125.035 ;
        RECT 47.325 124.355 50.075 125.165 ;
        RECT 50.095 124.440 50.525 125.225 ;
        RECT 53.745 125.035 54.675 125.265 ;
        RECT 50.775 124.355 54.675 125.035 ;
        RECT 55.605 124.355 61.115 125.165 ;
        RECT 64.325 125.035 65.255 125.265 ;
        RECT 61.355 124.355 65.255 125.035 ;
        RECT 65.265 124.355 66.635 125.165 ;
        RECT 69.845 125.035 70.775 125.265 ;
        RECT 66.875 124.355 70.775 125.035 ;
        RECT 70.795 124.355 72.145 125.265 ;
        RECT 72.625 124.355 73.995 125.135 ;
        RECT 74.465 124.355 75.835 125.135 ;
        RECT 75.855 124.440 76.285 125.225 ;
        RECT 77.235 124.355 78.585 125.265 ;
        RECT 78.975 125.155 79.895 125.265 ;
        RECT 78.975 125.035 81.310 125.155 ;
        RECT 85.975 125.035 86.895 125.255 ;
        RECT 78.975 124.355 88.255 125.035 ;
        RECT 89.195 124.355 90.545 125.265 ;
        RECT 90.565 125.035 91.495 125.265 ;
        RECT 90.565 124.355 94.465 125.035 ;
        RECT 94.705 124.355 97.455 125.165 ;
        RECT 100.665 125.035 101.595 125.265 ;
        RECT 97.695 124.355 101.595 125.035 ;
        RECT 101.615 124.440 102.045 125.225 ;
        RECT 102.265 125.175 103.215 125.265 ;
        RECT 102.265 124.355 104.195 125.175 ;
        RECT 104.375 124.355 105.725 125.265 ;
        RECT 109.405 125.035 110.335 125.265 ;
        RECT 114.005 125.035 114.935 125.265 ;
        RECT 106.435 124.355 110.335 125.035 ;
        RECT 111.035 124.355 114.935 125.035 ;
        RECT 115.315 125.155 116.235 125.265 ;
        RECT 115.315 125.035 117.650 125.155 ;
        RECT 122.315 125.035 123.235 125.255 ;
        RECT 115.315 124.355 124.595 125.035 ;
        RECT 124.605 124.355 125.975 125.135 ;
        RECT 126.445 124.355 127.815 125.165 ;
        RECT 20.785 124.145 20.955 124.355 ;
        RECT 22.220 124.195 22.340 124.305 ;
        RECT 22.625 124.200 22.785 124.310 ;
        RECT 24.005 124.165 24.175 124.355 ;
        RECT 24.925 124.165 25.095 124.355 ;
        RECT 26.305 124.165 26.475 124.355 ;
        RECT 27.960 124.165 28.130 124.355 ;
        RECT 31.825 124.145 31.995 124.335 ;
        RECT 32.285 124.200 32.445 124.310 ;
        RECT 32.745 124.190 32.905 124.300 ;
        RECT 36.610 124.145 36.780 124.335 ;
        RECT 37.805 124.145 37.975 124.335 ;
        RECT 41.945 124.165 42.115 124.355 ;
        RECT 42.460 124.195 42.580 124.305 ;
        RECT 46.270 124.165 46.440 124.355 ;
        RECT 47.060 124.195 47.180 124.305 ;
        RECT 48.385 124.145 48.555 124.335 ;
        RECT 49.765 124.165 49.935 124.355 ;
        RECT 54.090 124.165 54.260 124.355 ;
        RECT 55.285 124.200 55.445 124.310 ;
        RECT 58.045 124.145 58.215 124.335 ;
        RECT 58.560 124.195 58.680 124.305 ;
        RECT 60.805 124.165 60.975 124.355 ;
        RECT 61.265 124.145 61.435 124.335 ;
        RECT 61.725 124.145 61.895 124.335 ;
        RECT 64.025 124.190 64.185 124.300 ;
        RECT 64.670 124.165 64.840 124.355 ;
        RECT 65.405 124.145 65.575 124.335 ;
        RECT 66.325 124.165 66.495 124.355 ;
        RECT 70.190 124.165 70.360 124.355 ;
        RECT 71.845 124.165 72.015 124.355 ;
        RECT 72.360 124.195 72.480 124.305 ;
        RECT 72.765 124.165 72.935 124.355 ;
        RECT 74.200 124.195 74.320 124.305 ;
        RECT 74.605 124.165 74.775 124.355 ;
        RECT 75.065 124.145 75.235 124.335 ;
        RECT 75.580 124.195 75.700 124.305 ;
        RECT 75.985 124.145 76.155 124.335 ;
        RECT 76.905 124.200 77.065 124.310 ;
        RECT 77.365 124.165 77.535 124.355 ;
        RECT 86.565 124.145 86.735 124.335 ;
        RECT 87.945 124.145 88.115 124.355 ;
        RECT 88.460 124.195 88.580 124.305 ;
        RECT 88.865 124.200 89.025 124.310 ;
        RECT 89.325 124.145 89.495 124.355 ;
        RECT 90.705 124.145 90.875 124.335 ;
        RECT 90.980 124.165 91.150 124.355 ;
        RECT 97.145 124.165 97.315 124.355 ;
        RECT 101.010 124.165 101.180 124.355 ;
        RECT 104.045 124.335 104.195 124.355 ;
        RECT 101.285 124.145 101.455 124.335 ;
        RECT 104.045 124.165 104.215 124.335 ;
        RECT 104.505 124.165 104.675 124.355 ;
        RECT 105.940 124.195 106.060 124.305 ;
        RECT 109.750 124.165 109.920 124.355 ;
        RECT 110.540 124.195 110.660 124.305 ;
        RECT 110.945 124.145 111.115 124.335 ;
        RECT 112.325 124.145 112.495 124.335 ;
        RECT 113.705 124.145 113.875 124.335 ;
        RECT 114.220 124.195 114.340 124.305 ;
        RECT 114.350 124.165 114.520 124.355 ;
        RECT 115.360 124.145 115.530 124.335 ;
        RECT 119.225 124.145 119.395 124.335 ;
        RECT 120.660 124.195 120.780 124.305 ;
        RECT 124.285 124.165 124.455 124.355 ;
        RECT 125.665 124.165 125.835 124.355 ;
        RECT 126.125 124.305 126.295 124.335 ;
        RECT 126.125 124.195 126.300 124.305 ;
        RECT 126.125 124.145 126.295 124.195 ;
        RECT 127.505 124.145 127.675 124.355 ;
        RECT 20.645 123.335 22.015 124.145 ;
        RECT 22.855 123.465 32.135 124.145 ;
        RECT 33.295 123.465 37.195 124.145 ;
        RECT 22.855 123.345 25.190 123.465 ;
        RECT 22.855 123.235 23.775 123.345 ;
        RECT 29.855 123.245 30.775 123.465 ;
        RECT 36.265 123.235 37.195 123.465 ;
        RECT 37.215 123.275 37.645 124.060 ;
        RECT 37.665 123.365 39.035 124.145 ;
        RECT 39.415 123.465 48.695 124.145 ;
        RECT 49.075 123.465 58.355 124.145 ;
        RECT 39.415 123.345 41.750 123.465 ;
        RECT 39.415 123.235 40.335 123.345 ;
        RECT 46.415 123.245 47.335 123.465 ;
        RECT 49.075 123.345 51.410 123.465 ;
        RECT 49.075 123.235 49.995 123.345 ;
        RECT 56.075 123.245 56.995 123.465 ;
        RECT 58.825 123.335 61.575 124.145 ;
        RECT 61.595 123.235 62.945 124.145 ;
        RECT 62.975 123.275 63.405 124.060 ;
        RECT 64.345 123.365 65.715 124.145 ;
        RECT 66.095 123.465 75.375 124.145 ;
        RECT 75.845 123.465 85.125 124.145 ;
        RECT 66.095 123.345 68.430 123.465 ;
        RECT 66.095 123.235 67.015 123.345 ;
        RECT 73.095 123.245 74.015 123.465 ;
        RECT 77.205 123.245 78.125 123.465 ;
        RECT 82.790 123.345 85.125 123.465 ;
        RECT 84.205 123.235 85.125 123.345 ;
        RECT 85.515 123.235 86.865 124.145 ;
        RECT 86.885 123.365 88.255 124.145 ;
        RECT 88.735 123.275 89.165 124.060 ;
        RECT 89.195 123.235 90.545 124.145 ;
        RECT 90.565 123.365 91.935 124.145 ;
        RECT 92.315 123.465 101.595 124.145 ;
        RECT 101.975 123.465 111.255 124.145 ;
        RECT 92.315 123.345 94.650 123.465 ;
        RECT 92.315 123.235 93.235 123.345 ;
        RECT 99.315 123.245 100.235 123.465 ;
        RECT 101.975 123.345 104.310 123.465 ;
        RECT 101.975 123.235 102.895 123.345 ;
        RECT 108.975 123.245 109.895 123.465 ;
        RECT 111.265 123.365 112.635 124.145 ;
        RECT 112.655 123.235 114.005 124.145 ;
        RECT 114.495 123.275 114.925 124.060 ;
        RECT 114.945 123.465 118.845 124.145 ;
        RECT 114.945 123.235 115.875 123.465 ;
        RECT 119.095 123.235 120.445 124.145 ;
        RECT 120.925 123.335 126.435 124.145 ;
        RECT 126.445 123.335 127.815 124.145 ;
      LAYER nwell ;
        RECT 20.450 120.115 128.010 122.945 ;
      LAYER pwell ;
        RECT 20.645 118.915 22.015 119.725 ;
        RECT 22.485 118.915 24.315 119.725 ;
        RECT 24.335 119.000 24.765 119.785 ;
        RECT 25.155 119.715 26.075 119.825 ;
        RECT 25.155 119.595 27.490 119.715 ;
        RECT 32.155 119.595 33.075 119.815 ;
        RECT 25.155 118.915 34.435 119.595 ;
        RECT 34.445 118.915 35.815 119.725 ;
        RECT 35.835 118.915 37.185 119.825 ;
        RECT 37.205 118.915 42.715 119.725 ;
        RECT 42.735 118.915 44.085 119.825 ;
        RECT 44.105 118.915 45.935 119.725 ;
        RECT 45.945 118.915 47.315 119.695 ;
        RECT 47.325 118.915 50.075 119.725 ;
        RECT 50.095 119.000 50.525 119.785 ;
        RECT 50.545 118.915 52.375 119.725 ;
        RECT 52.395 118.915 53.745 119.825 ;
        RECT 54.685 118.915 56.055 119.695 ;
        RECT 56.665 118.915 59.275 119.825 ;
        RECT 61.105 119.595 62.025 119.815 ;
        RECT 68.105 119.715 69.025 119.825 ;
        RECT 66.690 119.595 69.025 119.715 ;
        RECT 59.745 118.915 69.025 119.595 ;
        RECT 69.415 118.915 70.765 119.825 ;
        RECT 71.245 118.915 72.615 119.695 ;
        RECT 73.085 118.915 75.835 119.725 ;
        RECT 75.855 119.000 76.285 119.785 ;
        RECT 76.305 118.915 81.815 119.725 ;
        RECT 85.025 119.595 85.955 119.825 ;
        RECT 82.055 118.915 85.955 119.595 ;
        RECT 86.335 119.715 87.255 119.825 ;
        RECT 86.335 119.595 88.670 119.715 ;
        RECT 93.335 119.595 94.255 119.815 ;
        RECT 86.335 118.915 95.615 119.595 ;
        RECT 96.545 118.915 100.215 119.725 ;
        RECT 100.225 118.915 101.595 119.695 ;
        RECT 101.615 119.000 102.045 119.785 ;
        RECT 102.525 118.915 108.035 119.725 ;
        RECT 108.415 119.715 109.335 119.825 ;
        RECT 108.415 119.595 110.750 119.715 ;
        RECT 115.415 119.595 116.335 119.815 ;
        RECT 108.415 118.915 117.695 119.595 ;
        RECT 118.165 118.915 120.915 119.725 ;
        RECT 120.925 118.915 126.435 119.725 ;
        RECT 126.445 118.915 127.815 119.725 ;
        RECT 20.785 118.705 20.955 118.915 ;
        RECT 22.220 118.755 22.340 118.865 ;
        RECT 24.005 118.725 24.175 118.915 ;
        RECT 25.385 118.705 25.555 118.895 ;
        RECT 30.905 118.705 31.075 118.895 ;
        RECT 31.365 118.705 31.535 118.895 ;
        RECT 33.205 118.750 33.365 118.860 ;
        RECT 34.125 118.725 34.295 118.915 ;
        RECT 35.505 118.725 35.675 118.915 ;
        RECT 35.965 118.725 36.135 118.915 ;
        RECT 36.885 118.705 37.055 118.895 ;
        RECT 37.860 118.755 37.980 118.865 ;
        RECT 40.565 118.705 40.735 118.895 ;
        RECT 42.405 118.725 42.575 118.915 ;
        RECT 43.785 118.725 43.955 118.915 ;
        RECT 45.625 118.725 45.795 118.915 ;
        RECT 46.085 118.705 46.255 118.915 ;
        RECT 49.765 118.725 49.935 118.915 ;
        RECT 51.605 118.705 51.775 118.895 ;
        RECT 52.065 118.725 52.235 118.915 ;
        RECT 53.445 118.725 53.615 118.915 ;
        RECT 54.365 118.760 54.525 118.870 ;
        RECT 54.825 118.725 54.995 118.915 ;
        RECT 56.260 118.755 56.380 118.865 ;
        RECT 57.125 118.705 57.295 118.895 ;
        RECT 58.960 118.725 59.130 118.915 ;
        RECT 59.480 118.755 59.600 118.865 ;
        RECT 59.885 118.725 60.055 118.915 ;
        RECT 62.645 118.705 62.815 118.895 ;
        RECT 63.620 118.755 63.740 118.865 ;
        RECT 66.325 118.705 66.495 118.895 ;
        RECT 70.465 118.725 70.635 118.915 ;
        RECT 70.980 118.755 71.100 118.865 ;
        RECT 71.385 118.725 71.555 118.915 ;
        RECT 71.845 118.705 72.015 118.895 ;
        RECT 72.820 118.755 72.940 118.865 ;
        RECT 75.525 118.725 75.695 118.915 ;
        RECT 77.365 118.705 77.535 118.895 ;
        RECT 81.505 118.725 81.675 118.915 ;
        RECT 82.885 118.705 83.055 118.895 ;
        RECT 85.370 118.725 85.540 118.915 ;
        RECT 88.405 118.705 88.575 118.895 ;
        RECT 89.380 118.755 89.500 118.865 ;
        RECT 92.085 118.705 92.255 118.895 ;
        RECT 95.305 118.725 95.475 118.915 ;
        RECT 96.225 118.760 96.385 118.870 ;
        RECT 97.605 118.705 97.775 118.895 ;
        RECT 99.905 118.725 100.075 118.915 ;
        RECT 101.285 118.725 101.455 118.915 ;
        RECT 102.260 118.755 102.380 118.865 ;
        RECT 103.125 118.705 103.295 118.895 ;
        RECT 107.725 118.725 107.895 118.915 ;
        RECT 108.645 118.705 108.815 118.895 ;
        RECT 114.165 118.705 114.335 118.895 ;
        RECT 115.085 118.705 115.255 118.895 ;
        RECT 116.520 118.755 116.640 118.865 ;
        RECT 117.385 118.725 117.555 118.915 ;
        RECT 117.900 118.755 118.020 118.865 ;
        RECT 119.225 118.705 119.395 118.895 ;
        RECT 119.685 118.705 119.855 118.895 ;
        RECT 120.605 118.725 120.775 118.915 ;
        RECT 121.065 118.705 121.235 118.895 ;
        RECT 123.365 118.705 123.535 118.895 ;
        RECT 126.125 118.705 126.295 118.915 ;
        RECT 127.505 118.705 127.675 118.915 ;
        RECT 20.645 117.895 22.015 118.705 ;
        RECT 22.025 117.895 25.695 118.705 ;
        RECT 25.705 117.895 31.215 118.705 ;
        RECT 31.225 117.925 32.595 118.705 ;
        RECT 33.525 117.895 37.195 118.705 ;
        RECT 37.215 117.835 37.645 118.620 ;
        RECT 38.125 117.895 40.875 118.705 ;
        RECT 40.885 117.895 46.395 118.705 ;
        RECT 46.405 117.895 51.915 118.705 ;
        RECT 51.925 117.895 57.435 118.705 ;
        RECT 57.445 117.895 62.955 118.705 ;
        RECT 62.975 117.835 63.405 118.620 ;
        RECT 63.885 117.895 66.635 118.705 ;
        RECT 66.645 117.895 72.155 118.705 ;
        RECT 72.165 117.895 77.675 118.705 ;
        RECT 77.685 117.895 83.195 118.705 ;
        RECT 83.205 117.895 88.715 118.705 ;
        RECT 88.735 117.835 89.165 118.620 ;
        RECT 89.645 117.895 92.395 118.705 ;
        RECT 92.405 117.895 97.915 118.705 ;
        RECT 97.925 117.895 103.435 118.705 ;
        RECT 103.445 117.895 108.955 118.705 ;
        RECT 108.965 117.895 114.475 118.705 ;
        RECT 114.495 117.835 114.925 118.620 ;
        RECT 114.945 117.925 116.315 118.705 ;
        RECT 116.785 117.895 119.535 118.705 ;
        RECT 119.555 117.795 120.905 118.705 ;
        RECT 120.925 117.925 122.295 118.705 ;
        RECT 122.305 117.925 123.675 118.705 ;
        RECT 123.685 117.895 126.435 118.705 ;
        RECT 126.445 117.895 127.815 118.705 ;
      LAYER nwell ;
        RECT 20.450 114.675 128.010 117.505 ;
      LAYER pwell ;
        RECT 20.645 113.475 22.015 114.285 ;
        RECT 22.485 113.475 24.315 114.285 ;
        RECT 24.335 113.560 24.765 114.345 ;
        RECT 24.785 113.475 26.615 114.285 ;
        RECT 26.625 114.155 27.545 114.385 ;
        RECT 30.375 114.155 31.305 114.375 ;
        RECT 26.625 113.475 35.815 114.155 ;
        RECT 35.825 113.475 37.195 114.255 ;
        RECT 37.205 113.475 38.575 114.255 ;
        RECT 38.595 113.475 39.945 114.385 ;
        RECT 39.965 113.475 45.475 114.285 ;
        RECT 45.485 113.475 46.855 114.255 ;
        RECT 46.865 113.475 48.235 114.285 ;
        RECT 48.255 113.475 49.605 114.385 ;
        RECT 50.095 113.560 50.525 114.345 ;
        RECT 51.005 113.475 53.755 114.285 ;
        RECT 53.765 113.475 55.135 114.255 ;
        RECT 55.145 113.475 56.975 114.285 ;
        RECT 56.985 113.475 62.495 114.285 ;
        RECT 62.505 113.475 65.115 114.385 ;
        RECT 65.265 113.475 70.775 114.285 ;
        RECT 70.785 113.475 72.155 114.255 ;
        RECT 72.165 113.475 75.835 114.285 ;
        RECT 75.855 113.560 76.285 114.345 ;
        RECT 76.765 113.475 78.595 114.285 ;
        RECT 78.615 113.475 79.965 114.385 ;
        RECT 79.995 113.475 81.345 114.385 ;
        RECT 81.365 113.475 82.735 114.255 ;
        RECT 83.205 113.475 85.815 114.385 ;
        RECT 85.965 113.475 87.335 114.255 ;
        RECT 87.805 113.475 93.315 114.285 ;
        RECT 93.335 113.475 94.685 114.385 ;
        RECT 94.705 113.475 96.075 114.255 ;
        RECT 96.085 113.475 97.455 114.285 ;
        RECT 97.475 113.475 98.825 114.385 ;
        RECT 98.845 113.475 101.595 114.285 ;
        RECT 101.615 113.560 102.045 114.345 ;
        RECT 102.525 113.475 104.355 114.285 ;
        RECT 104.375 113.475 105.725 114.385 ;
        RECT 106.665 113.475 108.035 114.255 ;
        RECT 108.055 113.475 109.405 114.385 ;
        RECT 110.345 113.475 115.855 114.285 ;
        RECT 115.875 113.475 117.225 114.385 ;
        RECT 121.755 114.155 122.685 114.375 ;
        RECT 125.515 114.155 126.435 114.385 ;
        RECT 117.245 113.475 126.435 114.155 ;
        RECT 126.445 113.475 127.815 114.285 ;
        RECT 20.785 113.265 20.955 113.475 ;
        RECT 22.220 113.315 22.340 113.425 ;
        RECT 23.545 113.265 23.715 113.455 ;
        RECT 24.005 113.285 24.175 113.475 ;
        RECT 24.925 113.265 25.095 113.455 ;
        RECT 25.385 113.265 25.555 113.455 ;
        RECT 26.305 113.285 26.475 113.475 ;
        RECT 26.765 113.265 26.935 113.455 ;
        RECT 35.505 113.285 35.675 113.475 ;
        RECT 36.885 113.265 37.055 113.475 ;
        RECT 37.805 113.265 37.975 113.455 ;
        RECT 38.265 113.285 38.435 113.475 ;
        RECT 39.185 113.265 39.355 113.455 ;
        RECT 39.645 113.285 39.815 113.475 ;
        RECT 45.165 113.285 45.335 113.475 ;
        RECT 45.625 113.285 45.795 113.475 ;
        RECT 47.925 113.285 48.095 113.475 ;
        RECT 49.305 113.265 49.475 113.475 ;
        RECT 50.685 113.425 50.855 113.455 ;
        RECT 49.820 113.315 49.940 113.425 ;
        RECT 50.685 113.315 50.860 113.425 ;
        RECT 51.200 113.315 51.320 113.425 ;
        RECT 50.685 113.265 50.855 113.315 ;
        RECT 53.445 113.285 53.615 113.475 ;
        RECT 53.905 113.285 54.075 113.475 ;
        RECT 56.665 113.285 56.835 113.475 ;
        RECT 60.345 113.265 60.515 113.455 ;
        RECT 60.805 113.265 60.975 113.455 ;
        RECT 62.185 113.285 62.355 113.475 ;
        RECT 62.650 113.420 62.820 113.475 ;
        RECT 62.645 113.310 62.820 113.420 ;
        RECT 62.650 113.285 62.820 113.310 ;
        RECT 64.485 113.265 64.655 113.455 ;
        RECT 64.945 113.265 65.115 113.455 ;
        RECT 70.465 113.285 70.635 113.475 ;
        RECT 70.925 113.285 71.095 113.475 ;
        RECT 75.065 113.265 75.235 113.455 ;
        RECT 75.525 113.285 75.695 113.475 ;
        RECT 76.445 113.425 76.615 113.455 ;
        RECT 76.445 113.315 76.620 113.425 ;
        RECT 76.445 113.265 76.615 113.315 ;
        RECT 77.825 113.265 77.995 113.455 ;
        RECT 78.285 113.285 78.455 113.475 ;
        RECT 79.665 113.285 79.835 113.475 ;
        RECT 80.125 113.285 80.295 113.475 ;
        RECT 81.505 113.285 81.675 113.475 ;
        RECT 82.940 113.315 83.060 113.425 ;
        RECT 83.350 113.285 83.520 113.475 ;
        RECT 86.105 113.285 86.275 113.475 ;
        RECT 87.025 113.265 87.195 113.455 ;
        RECT 87.540 113.315 87.660 113.425 ;
        RECT 88.405 113.265 88.575 113.455 ;
        RECT 90.245 113.265 90.415 113.455 ;
        RECT 93.005 113.285 93.175 113.475 ;
        RECT 94.385 113.285 94.555 113.475 ;
        RECT 94.845 113.285 95.015 113.475 ;
        RECT 97.145 113.285 97.315 113.475 ;
        RECT 97.605 113.285 97.775 113.475 ;
        RECT 99.445 113.265 99.615 113.455 ;
        RECT 100.825 113.265 100.995 113.455 ;
        RECT 101.285 113.425 101.455 113.475 ;
        RECT 101.285 113.315 101.460 113.425 ;
        RECT 102.260 113.315 102.380 113.425 ;
        RECT 101.285 113.285 101.455 113.315 ;
        RECT 104.045 113.285 104.215 113.475 ;
        RECT 105.425 113.285 105.595 113.475 ;
        RECT 106.345 113.320 106.505 113.430 ;
        RECT 106.805 113.285 106.975 113.475 ;
        RECT 109.105 113.285 109.275 113.475 ;
        RECT 110.025 113.320 110.185 113.430 ;
        RECT 110.485 113.265 110.655 113.455 ;
        RECT 110.945 113.265 111.115 113.455 ;
        RECT 112.785 113.310 112.945 113.420 ;
        RECT 113.245 113.265 113.415 113.455 ;
        RECT 115.140 113.315 115.260 113.425 ;
        RECT 115.545 113.265 115.715 113.475 ;
        RECT 116.005 113.285 116.175 113.475 ;
        RECT 116.980 113.315 117.100 113.425 ;
        RECT 117.385 113.285 117.555 113.475 ;
        RECT 126.125 113.265 126.295 113.455 ;
        RECT 127.505 113.265 127.675 113.475 ;
        RECT 20.645 112.455 22.015 113.265 ;
        RECT 22.025 112.455 23.855 113.265 ;
        RECT 23.875 112.355 25.225 113.265 ;
        RECT 25.255 112.355 26.605 113.265 ;
        RECT 26.635 112.355 27.985 113.265 ;
        RECT 28.005 112.585 37.195 113.265 ;
        RECT 28.005 112.355 28.925 112.585 ;
        RECT 31.755 112.365 32.685 112.585 ;
        RECT 37.215 112.395 37.645 113.180 ;
        RECT 37.665 112.485 39.035 113.265 ;
        RECT 39.055 112.355 40.405 113.265 ;
        RECT 40.425 112.585 49.615 113.265 ;
        RECT 40.425 112.355 41.345 112.585 ;
        RECT 44.175 112.365 45.105 112.585 ;
        RECT 49.625 112.485 50.995 113.265 ;
        RECT 51.465 112.585 60.655 113.265 ;
        RECT 51.465 112.355 52.385 112.585 ;
        RECT 55.215 112.365 56.145 112.585 ;
        RECT 60.665 112.485 62.035 113.265 ;
        RECT 62.975 112.395 63.405 113.180 ;
        RECT 63.425 112.455 64.795 113.265 ;
        RECT 64.805 112.485 66.175 113.265 ;
        RECT 66.185 112.585 75.375 113.265 ;
        RECT 66.185 112.355 67.105 112.585 ;
        RECT 69.935 112.365 70.865 112.585 ;
        RECT 75.385 112.455 76.755 113.265 ;
        RECT 76.775 112.355 78.125 113.265 ;
        RECT 78.145 112.585 87.335 113.265 ;
        RECT 78.145 112.355 79.065 112.585 ;
        RECT 81.895 112.365 82.825 112.585 ;
        RECT 87.345 112.485 88.715 113.265 ;
        RECT 88.735 112.395 89.165 113.180 ;
        RECT 89.195 112.355 90.545 113.265 ;
        RECT 90.565 112.585 99.755 113.265 ;
        RECT 90.565 112.355 91.485 112.585 ;
        RECT 94.315 112.365 95.245 112.585 ;
        RECT 99.765 112.485 101.135 113.265 ;
        RECT 101.605 112.585 110.795 113.265 ;
        RECT 101.605 112.355 102.525 112.585 ;
        RECT 105.355 112.365 106.285 112.585 ;
        RECT 110.805 112.485 112.175 113.265 ;
        RECT 113.105 112.485 114.475 113.265 ;
        RECT 114.495 112.395 114.925 113.180 ;
        RECT 115.415 112.355 116.765 113.265 ;
        RECT 117.245 112.585 126.435 113.265 ;
        RECT 117.245 112.355 118.165 112.585 ;
        RECT 120.995 112.365 121.925 112.585 ;
        RECT 126.445 112.455 127.815 113.265 ;
      LAYER nwell ;
        RECT 20.450 109.235 128.010 112.065 ;
      LAYER pwell ;
        RECT 20.645 108.035 22.015 108.845 ;
        RECT 22.485 108.035 24.315 108.845 ;
        RECT 24.335 108.120 24.765 108.905 ;
        RECT 24.785 108.035 30.295 108.845 ;
        RECT 30.305 108.035 31.675 108.815 ;
        RECT 36.195 108.715 37.125 108.935 ;
        RECT 39.955 108.715 40.875 108.945 ;
        RECT 45.395 108.715 46.325 108.935 ;
        RECT 49.155 108.715 50.075 108.945 ;
        RECT 31.685 108.035 40.875 108.715 ;
        RECT 40.885 108.035 50.075 108.715 ;
        RECT 50.095 108.120 50.525 108.905 ;
        RECT 51.005 108.035 53.755 108.845 ;
        RECT 53.775 108.035 55.125 108.945 ;
        RECT 55.155 108.035 56.505 108.945 ;
        RECT 56.525 108.715 57.445 108.945 ;
        RECT 60.275 108.715 61.205 108.935 ;
        RECT 65.725 108.715 66.645 108.945 ;
        RECT 69.475 108.715 70.405 108.935 ;
        RECT 56.525 108.035 65.715 108.715 ;
        RECT 65.725 108.035 74.915 108.715 ;
        RECT 75.855 108.120 76.285 108.905 ;
        RECT 76.305 108.715 77.225 108.945 ;
        RECT 80.055 108.715 80.985 108.935 ;
        RECT 90.015 108.715 90.945 108.935 ;
        RECT 93.775 108.715 94.695 108.945 ;
        RECT 76.305 108.035 85.495 108.715 ;
        RECT 85.505 108.035 94.695 108.715 ;
        RECT 94.705 108.035 96.075 108.845 ;
        RECT 96.085 108.035 101.595 108.845 ;
        RECT 101.615 108.120 102.045 108.905 ;
        RECT 102.525 108.035 105.275 108.845 ;
        RECT 105.285 108.715 106.205 108.945 ;
        RECT 109.035 108.715 109.965 108.935 ;
        RECT 114.485 108.715 115.405 108.945 ;
        RECT 118.235 108.715 119.165 108.935 ;
        RECT 105.285 108.035 114.475 108.715 ;
        RECT 114.485 108.035 123.675 108.715 ;
        RECT 123.685 108.035 125.055 108.845 ;
        RECT 125.065 108.035 126.435 108.815 ;
        RECT 126.445 108.035 127.815 108.845 ;
        RECT 20.785 107.825 20.955 108.035 ;
        RECT 22.220 107.875 22.340 107.985 ;
        RECT 24.005 107.825 24.175 108.035 ;
        RECT 29.985 107.845 30.155 108.035 ;
        RECT 30.445 107.845 30.615 108.035 ;
        RECT 31.825 107.845 31.995 108.035 ;
        RECT 33.665 107.825 33.835 108.015 ;
        RECT 34.180 107.875 34.300 107.985 ;
        RECT 36.885 107.825 37.055 108.015 ;
        RECT 38.725 107.825 38.895 108.015 ;
        RECT 41.025 107.845 41.195 108.035 ;
        RECT 44.245 107.825 44.415 108.015 ;
        RECT 49.765 107.825 49.935 108.015 ;
        RECT 50.740 107.875 50.860 107.985 ;
        RECT 51.605 107.825 51.775 108.015 ;
        RECT 53.445 107.845 53.615 108.035 ;
        RECT 53.905 107.845 54.075 108.035 ;
        RECT 55.285 107.845 55.455 108.035 ;
        RECT 57.125 107.825 57.295 108.015 ;
        RECT 62.645 107.825 62.815 108.015 ;
        RECT 64.945 107.825 65.115 108.015 ;
        RECT 65.405 107.825 65.575 108.035 ;
        RECT 66.840 107.875 66.960 107.985 ;
        RECT 67.245 107.825 67.415 108.015 ;
        RECT 70.005 107.825 70.175 108.015 ;
        RECT 74.605 107.845 74.775 108.035 ;
        RECT 75.525 107.825 75.695 108.015 ;
        RECT 77.365 107.825 77.535 108.015 ;
        RECT 82.885 107.825 83.055 108.015 ;
        RECT 85.185 107.845 85.355 108.035 ;
        RECT 85.645 107.845 85.815 108.035 ;
        RECT 88.405 107.825 88.575 108.015 ;
        RECT 89.380 107.875 89.500 107.985 ;
        RECT 92.085 107.825 92.255 108.015 ;
        RECT 92.545 107.825 92.715 108.015 ;
        RECT 95.765 107.845 95.935 108.035 ;
        RECT 101.285 107.845 101.455 108.035 ;
        RECT 102.260 107.875 102.380 107.985 ;
        RECT 103.125 107.825 103.295 108.015 ;
        RECT 104.965 107.845 105.135 108.035 ;
        RECT 108.645 107.825 108.815 108.015 ;
        RECT 114.165 107.825 114.335 108.035 ;
        RECT 115.140 107.875 115.260 107.985 ;
        RECT 120.605 107.825 120.775 108.015 ;
        RECT 123.365 107.845 123.535 108.035 ;
        RECT 124.745 107.845 124.915 108.035 ;
        RECT 126.115 108.015 126.285 108.035 ;
        RECT 126.115 107.845 126.295 108.015 ;
        RECT 126.125 107.825 126.295 107.845 ;
        RECT 127.505 107.825 127.675 108.035 ;
        RECT 20.645 107.015 22.015 107.825 ;
        RECT 22.485 107.015 24.315 107.825 ;
        RECT 24.335 106.955 24.765 107.740 ;
        RECT 24.785 107.145 33.975 107.825 ;
        RECT 24.785 106.915 25.705 107.145 ;
        RECT 28.535 106.925 29.465 107.145 ;
        RECT 34.445 107.015 37.195 107.825 ;
        RECT 37.215 106.955 37.645 107.740 ;
        RECT 37.665 107.015 39.035 107.825 ;
        RECT 39.045 107.015 44.555 107.825 ;
        RECT 44.565 107.015 50.075 107.825 ;
        RECT 50.095 106.955 50.525 107.740 ;
        RECT 50.545 107.015 51.915 107.825 ;
        RECT 51.925 107.015 57.435 107.825 ;
        RECT 57.445 107.015 62.955 107.825 ;
        RECT 62.975 106.955 63.405 107.740 ;
        RECT 63.425 107.015 65.255 107.825 ;
        RECT 65.275 106.915 66.625 107.825 ;
        RECT 67.115 106.915 68.465 107.825 ;
        RECT 68.485 107.015 70.315 107.825 ;
        RECT 70.325 107.015 75.835 107.825 ;
        RECT 75.855 106.955 76.285 107.740 ;
        RECT 76.305 107.015 77.675 107.825 ;
        RECT 77.685 107.015 83.195 107.825 ;
        RECT 83.205 107.015 88.715 107.825 ;
        RECT 88.735 106.955 89.165 107.740 ;
        RECT 89.645 107.015 92.395 107.825 ;
        RECT 92.405 107.145 101.595 107.825 ;
        RECT 96.915 106.925 97.845 107.145 ;
        RECT 100.675 106.915 101.595 107.145 ;
        RECT 101.615 106.955 102.045 107.740 ;
        RECT 102.065 107.015 103.435 107.825 ;
        RECT 103.445 107.015 108.955 107.825 ;
        RECT 108.965 107.015 114.475 107.825 ;
        RECT 114.495 106.955 114.925 107.740 ;
        RECT 115.405 107.015 120.915 107.825 ;
        RECT 120.925 107.015 126.435 107.825 ;
        RECT 126.445 107.015 127.815 107.825 ;
      LAYER nwell ;
        RECT 20.450 105.020 128.010 106.625 ;
        RECT 20.485 54.580 29.875 66.420 ;
        RECT 31.685 54.590 41.075 66.430 ;
        RECT 42.905 54.560 52.295 66.400 ;
        RECT 54.155 54.540 63.545 66.380 ;
        RECT 65.375 54.530 74.765 66.370 ;
        RECT 76.615 54.520 86.005 66.360 ;
        RECT 87.865 54.530 97.255 66.370 ;
        RECT 99.145 54.520 108.535 66.360 ;
        RECT 110.415 54.520 119.805 66.360 ;
        RECT 121.665 54.520 131.055 66.360 ;
        RECT 132.415 54.490 139.375 66.330 ;
        RECT 20.655 49.020 23.115 53.210 ;
      LAYER pwell ;
        RECT 20.555 45.340 22.915 48.340 ;
      LAYER nwell ;
        RECT 24.735 45.940 29.125 53.130 ;
        RECT 31.855 49.030 34.315 53.220 ;
      LAYER pwell ;
        RECT 31.755 45.350 34.115 48.350 ;
      LAYER nwell ;
        RECT 35.935 45.950 40.325 53.140 ;
        RECT 43.075 49.000 45.535 53.190 ;
      LAYER pwell ;
        RECT 42.975 45.320 45.335 48.320 ;
      LAYER nwell ;
        RECT 47.155 45.920 51.545 53.110 ;
        RECT 54.325 48.980 56.785 53.170 ;
      LAYER pwell ;
        RECT 54.225 45.300 56.585 48.300 ;
      LAYER nwell ;
        RECT 58.405 45.900 62.795 53.090 ;
        RECT 65.545 48.970 68.005 53.160 ;
      LAYER pwell ;
        RECT 65.445 45.290 67.805 48.290 ;
      LAYER nwell ;
        RECT 69.625 45.890 74.015 53.080 ;
        RECT 76.785 48.960 79.245 53.150 ;
      LAYER pwell ;
        RECT 76.685 45.280 79.045 48.280 ;
      LAYER nwell ;
        RECT 80.865 45.880 85.255 53.070 ;
        RECT 88.035 48.970 90.495 53.160 ;
      LAYER pwell ;
        RECT 87.935 45.290 90.295 48.290 ;
      LAYER nwell ;
        RECT 92.115 45.890 96.505 53.080 ;
        RECT 99.315 48.960 101.775 53.150 ;
      LAYER pwell ;
        RECT 99.215 45.280 101.575 48.280 ;
      LAYER nwell ;
        RECT 103.395 45.880 107.785 53.070 ;
        RECT 110.585 48.960 113.045 53.150 ;
      LAYER pwell ;
        RECT 110.485 45.280 112.845 48.280 ;
      LAYER nwell ;
        RECT 114.665 45.880 119.055 53.070 ;
        RECT 121.835 48.960 124.295 53.150 ;
      LAYER pwell ;
        RECT 121.735 45.280 124.095 48.280 ;
      LAYER nwell ;
        RECT 125.915 45.880 130.305 53.070 ;
        RECT 19.615 32.280 24.005 39.470 ;
      LAYER pwell ;
        RECT 25.825 37.070 28.185 40.070 ;
      LAYER nwell ;
        RECT 25.625 32.200 28.085 36.390 ;
        RECT 30.895 32.280 35.285 39.470 ;
      LAYER pwell ;
        RECT 37.105 37.070 39.465 40.070 ;
      LAYER nwell ;
        RECT 36.905 32.200 39.365 36.390 ;
        RECT 42.185 32.260 46.575 39.450 ;
      LAYER pwell ;
        RECT 48.395 37.050 50.755 40.050 ;
      LAYER nwell ;
        RECT 48.195 32.180 50.655 36.370 ;
        RECT 53.405 32.260 57.795 39.450 ;
      LAYER pwell ;
        RECT 59.615 37.050 61.975 40.050 ;
      LAYER nwell ;
        RECT 59.415 32.180 61.875 36.370 ;
        RECT 64.605 32.260 68.995 39.450 ;
      LAYER pwell ;
        RECT 70.815 37.050 73.175 40.050 ;
      LAYER nwell ;
        RECT 70.615 32.180 73.075 36.370 ;
        RECT 75.895 32.250 80.285 39.440 ;
      LAYER pwell ;
        RECT 82.105 37.040 84.465 40.040 ;
      LAYER nwell ;
        RECT 81.905 32.170 84.365 36.360 ;
        RECT 87.135 32.270 91.525 39.460 ;
      LAYER pwell ;
        RECT 93.345 37.060 95.705 40.060 ;
      LAYER nwell ;
        RECT 93.145 32.190 95.605 36.380 ;
        RECT 98.345 32.290 102.735 39.480 ;
      LAYER pwell ;
        RECT 104.555 37.080 106.915 40.080 ;
      LAYER nwell ;
        RECT 104.355 32.210 106.815 36.400 ;
        RECT 109.545 32.330 113.935 39.520 ;
      LAYER pwell ;
        RECT 115.755 37.120 118.115 40.120 ;
      LAYER nwell ;
        RECT 115.555 32.250 118.015 36.440 ;
        RECT 120.755 32.350 125.145 39.540 ;
      LAYER pwell ;
        RECT 126.965 37.140 129.325 40.140 ;
      LAYER nwell ;
        RECT 126.765 32.270 129.225 36.460 ;
        RECT 18.865 18.990 28.255 30.830 ;
        RECT 30.145 18.990 39.535 30.830 ;
        RECT 41.435 18.970 50.825 30.810 ;
        RECT 52.655 18.970 62.045 30.810 ;
        RECT 63.855 18.970 73.245 30.810 ;
        RECT 75.145 18.960 84.535 30.800 ;
        RECT 86.385 18.980 95.775 30.820 ;
        RECT 97.595 19.000 106.985 30.840 ;
        RECT 108.795 19.040 118.185 30.880 ;
        RECT 120.005 19.060 129.395 30.900 ;
        RECT 131.725 19.030 138.685 30.870 ;
      LAYER li1 ;
        RECT 20.640 211.205 127.820 211.375 ;
        RECT 20.725 210.455 21.935 211.205 ;
        RECT 20.725 209.915 21.245 210.455 ;
        RECT 22.565 210.435 24.235 211.205 ;
        RECT 24.405 210.480 24.695 211.205 ;
        RECT 24.865 210.455 26.075 211.205 ;
        RECT 26.250 210.660 31.595 211.205 ;
        RECT 31.770 210.660 37.115 211.205 ;
        RECT 21.415 209.745 21.935 210.285 ;
        RECT 20.725 208.655 21.935 209.745 ;
        RECT 22.565 209.745 23.315 210.265 ;
        RECT 23.485 209.915 24.235 210.435 ;
        RECT 22.565 208.655 24.235 209.745 ;
        RECT 24.405 208.655 24.695 209.820 ;
        RECT 24.865 209.745 25.385 210.285 ;
        RECT 25.555 209.915 26.075 210.455 ;
        RECT 24.865 208.655 26.075 209.745 ;
        RECT 27.840 209.090 28.190 210.340 ;
        RECT 29.670 209.830 30.010 210.660 ;
        RECT 33.360 209.090 33.710 210.340 ;
        RECT 35.190 209.830 35.530 210.660 ;
        RECT 37.285 210.480 37.575 211.205 ;
        RECT 37.745 210.455 38.955 211.205 ;
        RECT 39.130 210.660 44.475 211.205 ;
        RECT 44.650 210.660 49.995 211.205 ;
        RECT 26.250 208.655 31.595 209.090 ;
        RECT 31.770 208.655 37.115 209.090 ;
        RECT 37.285 208.655 37.575 209.820 ;
        RECT 37.745 209.745 38.265 210.285 ;
        RECT 38.435 209.915 38.955 210.455 ;
        RECT 37.745 208.655 38.955 209.745 ;
        RECT 40.720 209.090 41.070 210.340 ;
        RECT 42.550 209.830 42.890 210.660 ;
        RECT 46.240 209.090 46.590 210.340 ;
        RECT 48.070 209.830 48.410 210.660 ;
        RECT 50.165 210.480 50.455 211.205 ;
        RECT 50.625 210.455 51.835 211.205 ;
        RECT 52.010 210.660 57.355 211.205 ;
        RECT 57.530 210.660 62.875 211.205 ;
        RECT 39.130 208.655 44.475 209.090 ;
        RECT 44.650 208.655 49.995 209.090 ;
        RECT 50.165 208.655 50.455 209.820 ;
        RECT 50.625 209.745 51.145 210.285 ;
        RECT 51.315 209.915 51.835 210.455 ;
        RECT 50.625 208.655 51.835 209.745 ;
        RECT 53.600 209.090 53.950 210.340 ;
        RECT 55.430 209.830 55.770 210.660 ;
        RECT 59.120 209.090 59.470 210.340 ;
        RECT 60.950 209.830 61.290 210.660 ;
        RECT 63.045 210.480 63.335 211.205 ;
        RECT 63.505 210.455 64.715 211.205 ;
        RECT 64.890 210.660 70.235 211.205 ;
        RECT 70.410 210.660 75.755 211.205 ;
        RECT 52.010 208.655 57.355 209.090 ;
        RECT 57.530 208.655 62.875 209.090 ;
        RECT 63.045 208.655 63.335 209.820 ;
        RECT 63.505 209.745 64.025 210.285 ;
        RECT 64.195 209.915 64.715 210.455 ;
        RECT 63.505 208.655 64.715 209.745 ;
        RECT 66.480 209.090 66.830 210.340 ;
        RECT 68.310 209.830 68.650 210.660 ;
        RECT 72.000 209.090 72.350 210.340 ;
        RECT 73.830 209.830 74.170 210.660 ;
        RECT 75.925 210.480 76.215 211.205 ;
        RECT 76.385 210.455 77.595 211.205 ;
        RECT 77.770 210.660 83.115 211.205 ;
        RECT 83.290 210.660 88.635 211.205 ;
        RECT 64.890 208.655 70.235 209.090 ;
        RECT 70.410 208.655 75.755 209.090 ;
        RECT 75.925 208.655 76.215 209.820 ;
        RECT 76.385 209.745 76.905 210.285 ;
        RECT 77.075 209.915 77.595 210.455 ;
        RECT 76.385 208.655 77.595 209.745 ;
        RECT 79.360 209.090 79.710 210.340 ;
        RECT 81.190 209.830 81.530 210.660 ;
        RECT 84.880 209.090 85.230 210.340 ;
        RECT 86.710 209.830 87.050 210.660 ;
        RECT 88.805 210.480 89.095 211.205 ;
        RECT 89.265 210.455 90.475 211.205 ;
        RECT 90.650 210.660 95.995 211.205 ;
        RECT 96.170 210.660 101.515 211.205 ;
        RECT 77.770 208.655 83.115 209.090 ;
        RECT 83.290 208.655 88.635 209.090 ;
        RECT 88.805 208.655 89.095 209.820 ;
        RECT 89.265 209.745 89.785 210.285 ;
        RECT 89.955 209.915 90.475 210.455 ;
        RECT 89.265 208.655 90.475 209.745 ;
        RECT 92.240 209.090 92.590 210.340 ;
        RECT 94.070 209.830 94.410 210.660 ;
        RECT 97.760 209.090 98.110 210.340 ;
        RECT 99.590 209.830 99.930 210.660 ;
        RECT 101.685 210.480 101.975 211.205 ;
        RECT 102.145 210.455 103.355 211.205 ;
        RECT 103.530 210.660 108.875 211.205 ;
        RECT 109.050 210.660 114.395 211.205 ;
        RECT 90.650 208.655 95.995 209.090 ;
        RECT 96.170 208.655 101.515 209.090 ;
        RECT 101.685 208.655 101.975 209.820 ;
        RECT 102.145 209.745 102.665 210.285 ;
        RECT 102.835 209.915 103.355 210.455 ;
        RECT 102.145 208.655 103.355 209.745 ;
        RECT 105.120 209.090 105.470 210.340 ;
        RECT 106.950 209.830 107.290 210.660 ;
        RECT 110.640 209.090 110.990 210.340 ;
        RECT 112.470 209.830 112.810 210.660 ;
        RECT 114.565 210.480 114.855 211.205 ;
        RECT 115.490 210.660 120.835 211.205 ;
        RECT 121.010 210.660 126.355 211.205 ;
        RECT 103.530 208.655 108.875 209.090 ;
        RECT 109.050 208.655 114.395 209.090 ;
        RECT 114.565 208.655 114.855 209.820 ;
        RECT 117.080 209.090 117.430 210.340 ;
        RECT 118.910 209.830 119.250 210.660 ;
        RECT 122.600 209.090 122.950 210.340 ;
        RECT 124.430 209.830 124.770 210.660 ;
        RECT 126.525 210.455 127.735 211.205 ;
        RECT 126.525 209.745 127.045 210.285 ;
        RECT 127.215 209.915 127.735 210.455 ;
        RECT 115.490 208.655 120.835 209.090 ;
        RECT 121.010 208.655 126.355 209.090 ;
        RECT 126.525 208.655 127.735 209.745 ;
        RECT 20.640 208.485 127.820 208.655 ;
        RECT 20.725 207.395 21.935 208.485 ;
        RECT 20.725 206.685 21.245 207.225 ;
        RECT 21.415 206.855 21.935 207.395 ;
        RECT 22.565 207.395 24.235 208.485 ;
        RECT 22.565 206.875 23.315 207.395 ;
        RECT 24.405 207.320 24.695 208.485 ;
        RECT 25.325 207.395 27.915 208.485 ;
        RECT 28.090 208.050 33.435 208.485 ;
        RECT 33.610 208.050 38.955 208.485 ;
        RECT 39.130 208.050 44.475 208.485 ;
        RECT 44.650 208.050 49.995 208.485 ;
        RECT 23.485 206.705 24.235 207.225 ;
        RECT 25.325 206.875 26.535 207.395 ;
        RECT 26.705 206.705 27.915 207.225 ;
        RECT 29.680 206.800 30.030 208.050 ;
        RECT 20.725 205.935 21.935 206.685 ;
        RECT 22.565 205.935 24.235 206.705 ;
        RECT 24.405 205.935 24.695 206.660 ;
        RECT 25.325 205.935 27.915 206.705 ;
        RECT 31.510 206.480 31.850 207.310 ;
        RECT 35.200 206.800 35.550 208.050 ;
        RECT 37.030 206.480 37.370 207.310 ;
        RECT 40.720 206.800 41.070 208.050 ;
        RECT 42.550 206.480 42.890 207.310 ;
        RECT 46.240 206.800 46.590 208.050 ;
        RECT 50.165 207.320 50.455 208.485 ;
        RECT 51.085 207.395 53.675 208.485 ;
        RECT 53.850 208.050 59.195 208.485 ;
        RECT 59.370 208.050 64.715 208.485 ;
        RECT 64.890 208.050 70.235 208.485 ;
        RECT 70.410 208.050 75.755 208.485 ;
        RECT 48.070 206.480 48.410 207.310 ;
        RECT 51.085 206.875 52.295 207.395 ;
        RECT 52.465 206.705 53.675 207.225 ;
        RECT 55.440 206.800 55.790 208.050 ;
        RECT 28.090 205.935 33.435 206.480 ;
        RECT 33.610 205.935 38.955 206.480 ;
        RECT 39.130 205.935 44.475 206.480 ;
        RECT 44.650 205.935 49.995 206.480 ;
        RECT 50.165 205.935 50.455 206.660 ;
        RECT 51.085 205.935 53.675 206.705 ;
        RECT 57.270 206.480 57.610 207.310 ;
        RECT 60.960 206.800 61.310 208.050 ;
        RECT 62.790 206.480 63.130 207.310 ;
        RECT 66.480 206.800 66.830 208.050 ;
        RECT 68.310 206.480 68.650 207.310 ;
        RECT 72.000 206.800 72.350 208.050 ;
        RECT 75.925 207.320 76.215 208.485 ;
        RECT 76.845 207.395 79.435 208.485 ;
        RECT 79.610 208.050 84.955 208.485 ;
        RECT 85.130 208.050 90.475 208.485 ;
        RECT 90.650 208.050 95.995 208.485 ;
        RECT 96.170 208.050 101.515 208.485 ;
        RECT 73.830 206.480 74.170 207.310 ;
        RECT 76.845 206.875 78.055 207.395 ;
        RECT 78.225 206.705 79.435 207.225 ;
        RECT 81.200 206.800 81.550 208.050 ;
        RECT 53.850 205.935 59.195 206.480 ;
        RECT 59.370 205.935 64.715 206.480 ;
        RECT 64.890 205.935 70.235 206.480 ;
        RECT 70.410 205.935 75.755 206.480 ;
        RECT 75.925 205.935 76.215 206.660 ;
        RECT 76.845 205.935 79.435 206.705 ;
        RECT 83.030 206.480 83.370 207.310 ;
        RECT 86.720 206.800 87.070 208.050 ;
        RECT 88.550 206.480 88.890 207.310 ;
        RECT 92.240 206.800 92.590 208.050 ;
        RECT 94.070 206.480 94.410 207.310 ;
        RECT 97.760 206.800 98.110 208.050 ;
        RECT 101.685 207.320 101.975 208.485 ;
        RECT 102.605 207.395 104.275 208.485 ;
        RECT 104.450 208.050 109.795 208.485 ;
        RECT 109.970 208.050 115.315 208.485 ;
        RECT 115.490 208.050 120.835 208.485 ;
        RECT 121.010 208.050 126.355 208.485 ;
        RECT 99.590 206.480 99.930 207.310 ;
        RECT 102.605 206.875 103.355 207.395 ;
        RECT 103.525 206.705 104.275 207.225 ;
        RECT 106.040 206.800 106.390 208.050 ;
        RECT 79.610 205.935 84.955 206.480 ;
        RECT 85.130 205.935 90.475 206.480 ;
        RECT 90.650 205.935 95.995 206.480 ;
        RECT 96.170 205.935 101.515 206.480 ;
        RECT 101.685 205.935 101.975 206.660 ;
        RECT 102.605 205.935 104.275 206.705 ;
        RECT 107.870 206.480 108.210 207.310 ;
        RECT 111.560 206.800 111.910 208.050 ;
        RECT 113.390 206.480 113.730 207.310 ;
        RECT 117.080 206.800 117.430 208.050 ;
        RECT 118.910 206.480 119.250 207.310 ;
        RECT 122.600 206.800 122.950 208.050 ;
        RECT 126.525 207.395 127.735 208.485 ;
        RECT 124.430 206.480 124.770 207.310 ;
        RECT 126.525 206.855 127.045 207.395 ;
        RECT 127.215 206.685 127.735 207.225 ;
        RECT 104.450 205.935 109.795 206.480 ;
        RECT 109.970 205.935 115.315 206.480 ;
        RECT 115.490 205.935 120.835 206.480 ;
        RECT 121.010 205.935 126.355 206.480 ;
        RECT 126.525 205.935 127.735 206.685 ;
        RECT 20.640 205.765 127.820 205.935 ;
        RECT 20.725 205.015 21.935 205.765 ;
        RECT 20.725 204.475 21.245 205.015 ;
        RECT 22.565 204.995 26.075 205.765 ;
        RECT 26.250 205.220 31.595 205.765 ;
        RECT 31.770 205.220 37.115 205.765 ;
        RECT 21.415 204.305 21.935 204.845 ;
        RECT 20.725 203.215 21.935 204.305 ;
        RECT 22.565 204.305 24.255 204.825 ;
        RECT 24.425 204.475 26.075 204.995 ;
        RECT 22.565 203.215 26.075 204.305 ;
        RECT 27.840 203.650 28.190 204.900 ;
        RECT 29.670 204.390 30.010 205.220 ;
        RECT 33.360 203.650 33.710 204.900 ;
        RECT 35.190 204.390 35.530 205.220 ;
        RECT 37.285 205.040 37.575 205.765 ;
        RECT 38.205 204.995 40.795 205.765 ;
        RECT 40.970 205.220 46.315 205.765 ;
        RECT 46.490 205.220 51.835 205.765 ;
        RECT 52.010 205.220 57.355 205.765 ;
        RECT 57.530 205.220 62.875 205.765 ;
        RECT 26.250 203.215 31.595 203.650 ;
        RECT 31.770 203.215 37.115 203.650 ;
        RECT 37.285 203.215 37.575 204.380 ;
        RECT 38.205 204.305 39.415 204.825 ;
        RECT 39.585 204.475 40.795 204.995 ;
        RECT 38.205 203.215 40.795 204.305 ;
        RECT 42.560 203.650 42.910 204.900 ;
        RECT 44.390 204.390 44.730 205.220 ;
        RECT 48.080 203.650 48.430 204.900 ;
        RECT 49.910 204.390 50.250 205.220 ;
        RECT 53.600 203.650 53.950 204.900 ;
        RECT 55.430 204.390 55.770 205.220 ;
        RECT 59.120 203.650 59.470 204.900 ;
        RECT 60.950 204.390 61.290 205.220 ;
        RECT 63.045 205.040 63.335 205.765 ;
        RECT 63.965 204.995 66.555 205.765 ;
        RECT 66.730 205.220 72.075 205.765 ;
        RECT 72.250 205.220 77.595 205.765 ;
        RECT 77.770 205.220 83.115 205.765 ;
        RECT 83.290 205.220 88.635 205.765 ;
        RECT 40.970 203.215 46.315 203.650 ;
        RECT 46.490 203.215 51.835 203.650 ;
        RECT 52.010 203.215 57.355 203.650 ;
        RECT 57.530 203.215 62.875 203.650 ;
        RECT 63.045 203.215 63.335 204.380 ;
        RECT 63.965 204.305 65.175 204.825 ;
        RECT 65.345 204.475 66.555 204.995 ;
        RECT 63.965 203.215 66.555 204.305 ;
        RECT 68.320 203.650 68.670 204.900 ;
        RECT 70.150 204.390 70.490 205.220 ;
        RECT 73.840 203.650 74.190 204.900 ;
        RECT 75.670 204.390 76.010 205.220 ;
        RECT 79.360 203.650 79.710 204.900 ;
        RECT 81.190 204.390 81.530 205.220 ;
        RECT 84.880 203.650 85.230 204.900 ;
        RECT 86.710 204.390 87.050 205.220 ;
        RECT 88.805 205.040 89.095 205.765 ;
        RECT 89.725 204.995 92.315 205.765 ;
        RECT 92.490 205.220 97.835 205.765 ;
        RECT 98.010 205.220 103.355 205.765 ;
        RECT 103.530 205.220 108.875 205.765 ;
        RECT 109.050 205.220 114.395 205.765 ;
        RECT 66.730 203.215 72.075 203.650 ;
        RECT 72.250 203.215 77.595 203.650 ;
        RECT 77.770 203.215 83.115 203.650 ;
        RECT 83.290 203.215 88.635 203.650 ;
        RECT 88.805 203.215 89.095 204.380 ;
        RECT 89.725 204.305 90.935 204.825 ;
        RECT 91.105 204.475 92.315 204.995 ;
        RECT 89.725 203.215 92.315 204.305 ;
        RECT 94.080 203.650 94.430 204.900 ;
        RECT 95.910 204.390 96.250 205.220 ;
        RECT 99.600 203.650 99.950 204.900 ;
        RECT 101.430 204.390 101.770 205.220 ;
        RECT 105.120 203.650 105.470 204.900 ;
        RECT 106.950 204.390 107.290 205.220 ;
        RECT 110.640 203.650 110.990 204.900 ;
        RECT 112.470 204.390 112.810 205.220 ;
        RECT 114.565 205.040 114.855 205.765 ;
        RECT 115.490 205.220 120.835 205.765 ;
        RECT 121.010 205.220 126.355 205.765 ;
        RECT 92.490 203.215 97.835 203.650 ;
        RECT 98.010 203.215 103.355 203.650 ;
        RECT 103.530 203.215 108.875 203.650 ;
        RECT 109.050 203.215 114.395 203.650 ;
        RECT 114.565 203.215 114.855 204.380 ;
        RECT 117.080 203.650 117.430 204.900 ;
        RECT 118.910 204.390 119.250 205.220 ;
        RECT 122.600 203.650 122.950 204.900 ;
        RECT 124.430 204.390 124.770 205.220 ;
        RECT 126.525 205.015 127.735 205.765 ;
        RECT 126.525 204.305 127.045 204.845 ;
        RECT 127.215 204.475 127.735 205.015 ;
        RECT 115.490 203.215 120.835 203.650 ;
        RECT 121.010 203.215 126.355 203.650 ;
        RECT 126.525 203.215 127.735 204.305 ;
        RECT 20.640 203.045 127.820 203.215 ;
        RECT 20.725 201.955 21.935 203.045 ;
        RECT 20.725 201.245 21.245 201.785 ;
        RECT 21.415 201.415 21.935 201.955 ;
        RECT 22.565 201.955 24.235 203.045 ;
        RECT 22.565 201.435 23.315 201.955 ;
        RECT 24.405 201.880 24.695 203.045 ;
        RECT 25.325 201.955 27.915 203.045 ;
        RECT 28.090 202.610 33.435 203.045 ;
        RECT 33.610 202.610 38.955 203.045 ;
        RECT 39.130 202.610 44.475 203.045 ;
        RECT 44.650 202.610 49.995 203.045 ;
        RECT 23.485 201.265 24.235 201.785 ;
        RECT 25.325 201.435 26.535 201.955 ;
        RECT 26.705 201.265 27.915 201.785 ;
        RECT 29.680 201.360 30.030 202.610 ;
        RECT 20.725 200.495 21.935 201.245 ;
        RECT 22.565 200.495 24.235 201.265 ;
        RECT 24.405 200.495 24.695 201.220 ;
        RECT 25.325 200.495 27.915 201.265 ;
        RECT 31.510 201.040 31.850 201.870 ;
        RECT 35.200 201.360 35.550 202.610 ;
        RECT 37.030 201.040 37.370 201.870 ;
        RECT 40.720 201.360 41.070 202.610 ;
        RECT 42.550 201.040 42.890 201.870 ;
        RECT 46.240 201.360 46.590 202.610 ;
        RECT 50.165 201.880 50.455 203.045 ;
        RECT 51.085 201.955 53.675 203.045 ;
        RECT 53.850 202.610 59.195 203.045 ;
        RECT 59.370 202.610 64.715 203.045 ;
        RECT 64.890 202.610 70.235 203.045 ;
        RECT 48.070 201.040 48.410 201.870 ;
        RECT 51.085 201.435 52.295 201.955 ;
        RECT 52.465 201.265 53.675 201.785 ;
        RECT 55.440 201.360 55.790 202.610 ;
        RECT 28.090 200.495 33.435 201.040 ;
        RECT 33.610 200.495 38.955 201.040 ;
        RECT 39.130 200.495 44.475 201.040 ;
        RECT 44.650 200.495 49.995 201.040 ;
        RECT 50.165 200.495 50.455 201.220 ;
        RECT 51.085 200.495 53.675 201.265 ;
        RECT 57.270 201.040 57.610 201.870 ;
        RECT 60.960 201.360 61.310 202.610 ;
        RECT 62.790 201.040 63.130 201.870 ;
        RECT 66.480 201.360 66.830 202.610 ;
        RECT 70.425 202.535 70.725 203.045 ;
        RECT 70.895 202.535 71.275 202.705 ;
        RECT 71.855 202.535 72.485 203.045 ;
        RECT 70.895 202.365 71.065 202.535 ;
        RECT 72.655 202.365 72.985 202.875 ;
        RECT 73.155 202.535 73.455 203.045 ;
        RECT 70.405 202.165 71.065 202.365 ;
        RECT 71.235 202.195 73.455 202.365 ;
        RECT 68.310 201.040 68.650 201.870 ;
        RECT 70.405 201.235 70.575 202.165 ;
        RECT 71.235 201.995 71.405 202.195 ;
        RECT 70.745 201.825 71.405 201.995 ;
        RECT 71.575 201.855 73.115 202.025 ;
        RECT 70.745 201.405 70.915 201.825 ;
        RECT 71.575 201.655 71.745 201.855 ;
        RECT 71.145 201.485 71.745 201.655 ;
        RECT 71.915 201.485 72.610 201.685 ;
        RECT 72.870 201.405 73.115 201.855 ;
        RECT 71.235 201.235 72.145 201.315 ;
        RECT 53.850 200.495 59.195 201.040 ;
        RECT 59.370 200.495 64.715 201.040 ;
        RECT 64.890 200.495 70.235 201.040 ;
        RECT 70.405 200.755 70.725 201.235 ;
        RECT 70.895 201.145 72.145 201.235 ;
        RECT 70.895 201.065 71.405 201.145 ;
        RECT 70.895 200.665 71.125 201.065 ;
        RECT 71.295 200.495 71.645 200.885 ;
        RECT 71.815 200.665 72.145 201.145 ;
        RECT 72.315 200.495 72.485 201.315 ;
        RECT 73.285 201.235 73.455 202.195 ;
        RECT 74.085 201.955 75.755 203.045 ;
        RECT 74.085 201.435 74.835 201.955 ;
        RECT 75.925 201.880 76.215 203.045 ;
        RECT 76.845 201.955 79.435 203.045 ;
        RECT 79.610 202.610 84.955 203.045 ;
        RECT 85.130 202.610 90.475 203.045 ;
        RECT 90.650 202.610 95.995 203.045 ;
        RECT 96.170 202.610 101.515 203.045 ;
        RECT 75.005 201.265 75.755 201.785 ;
        RECT 76.845 201.435 78.055 201.955 ;
        RECT 78.225 201.265 79.435 201.785 ;
        RECT 81.200 201.360 81.550 202.610 ;
        RECT 72.990 200.690 73.455 201.235 ;
        RECT 74.085 200.495 75.755 201.265 ;
        RECT 75.925 200.495 76.215 201.220 ;
        RECT 76.845 200.495 79.435 201.265 ;
        RECT 83.030 201.040 83.370 201.870 ;
        RECT 86.720 201.360 87.070 202.610 ;
        RECT 88.550 201.040 88.890 201.870 ;
        RECT 92.240 201.360 92.590 202.610 ;
        RECT 94.070 201.040 94.410 201.870 ;
        RECT 97.760 201.360 98.110 202.610 ;
        RECT 101.685 201.880 101.975 203.045 ;
        RECT 102.605 201.955 104.275 203.045 ;
        RECT 104.450 202.610 109.795 203.045 ;
        RECT 109.970 202.610 115.315 203.045 ;
        RECT 115.490 202.610 120.835 203.045 ;
        RECT 121.010 202.610 126.355 203.045 ;
        RECT 99.590 201.040 99.930 201.870 ;
        RECT 102.605 201.435 103.355 201.955 ;
        RECT 103.525 201.265 104.275 201.785 ;
        RECT 106.040 201.360 106.390 202.610 ;
        RECT 79.610 200.495 84.955 201.040 ;
        RECT 85.130 200.495 90.475 201.040 ;
        RECT 90.650 200.495 95.995 201.040 ;
        RECT 96.170 200.495 101.515 201.040 ;
        RECT 101.685 200.495 101.975 201.220 ;
        RECT 102.605 200.495 104.275 201.265 ;
        RECT 107.870 201.040 108.210 201.870 ;
        RECT 111.560 201.360 111.910 202.610 ;
        RECT 113.390 201.040 113.730 201.870 ;
        RECT 117.080 201.360 117.430 202.610 ;
        RECT 118.910 201.040 119.250 201.870 ;
        RECT 122.600 201.360 122.950 202.610 ;
        RECT 126.525 201.955 127.735 203.045 ;
        RECT 124.430 201.040 124.770 201.870 ;
        RECT 126.525 201.415 127.045 201.955 ;
        RECT 127.215 201.245 127.735 201.785 ;
        RECT 104.450 200.495 109.795 201.040 ;
        RECT 109.970 200.495 115.315 201.040 ;
        RECT 115.490 200.495 120.835 201.040 ;
        RECT 121.010 200.495 126.355 201.040 ;
        RECT 126.525 200.495 127.735 201.245 ;
        RECT 20.640 200.325 127.820 200.495 ;
        RECT 20.725 199.575 21.935 200.325 ;
        RECT 20.725 199.035 21.245 199.575 ;
        RECT 22.565 199.555 26.075 200.325 ;
        RECT 26.250 199.780 31.595 200.325 ;
        RECT 31.770 199.780 37.115 200.325 ;
        RECT 21.415 198.865 21.935 199.405 ;
        RECT 20.725 197.775 21.935 198.865 ;
        RECT 22.565 198.865 24.255 199.385 ;
        RECT 24.425 199.035 26.075 199.555 ;
        RECT 22.565 197.775 26.075 198.865 ;
        RECT 27.840 198.210 28.190 199.460 ;
        RECT 29.670 198.950 30.010 199.780 ;
        RECT 33.360 198.210 33.710 199.460 ;
        RECT 35.190 198.950 35.530 199.780 ;
        RECT 37.285 199.600 37.575 200.325 ;
        RECT 37.745 199.555 40.335 200.325 ;
        RECT 40.510 199.780 45.855 200.325 ;
        RECT 26.250 197.775 31.595 198.210 ;
        RECT 31.770 197.775 37.115 198.210 ;
        RECT 37.285 197.775 37.575 198.940 ;
        RECT 37.745 198.865 38.955 199.385 ;
        RECT 39.125 199.035 40.335 199.555 ;
        RECT 37.745 197.775 40.335 198.865 ;
        RECT 42.100 198.210 42.450 199.460 ;
        RECT 43.930 198.950 44.270 199.780 ;
        RECT 46.030 199.775 46.285 200.065 ;
        RECT 46.455 199.945 46.785 200.325 ;
        RECT 46.030 199.605 46.780 199.775 ;
        RECT 46.030 198.785 46.380 199.435 ;
        RECT 46.550 198.615 46.780 199.605 ;
        RECT 46.030 198.445 46.780 198.615 ;
        RECT 40.510 197.775 45.855 198.210 ;
        RECT 46.030 197.945 46.285 198.445 ;
        RECT 46.455 197.775 46.785 198.275 ;
        RECT 46.955 197.945 47.125 200.065 ;
        RECT 47.485 199.965 47.815 200.325 ;
        RECT 47.985 199.935 48.480 200.105 ;
        RECT 48.685 199.935 49.540 200.105 ;
        RECT 47.355 198.745 47.815 199.795 ;
        RECT 47.295 197.960 47.620 198.745 ;
        RECT 47.985 198.575 48.155 199.935 ;
        RECT 48.325 199.025 48.675 199.645 ;
        RECT 48.845 199.425 49.200 199.645 ;
        RECT 48.845 198.835 49.015 199.425 ;
        RECT 49.370 199.225 49.540 199.935 ;
        RECT 50.415 199.865 50.745 200.325 ;
        RECT 50.955 199.965 51.305 200.135 ;
        RECT 49.745 199.395 50.535 199.645 ;
        RECT 50.955 199.575 51.215 199.965 ;
        RECT 51.525 199.875 52.475 200.155 ;
        RECT 52.645 199.885 52.835 200.325 ;
        RECT 53.005 199.945 54.075 200.115 ;
        RECT 50.705 199.225 50.875 199.405 ;
        RECT 47.985 198.405 48.380 198.575 ;
        RECT 48.550 198.445 49.015 198.835 ;
        RECT 49.185 199.055 50.875 199.225 ;
        RECT 48.210 198.275 48.380 198.405 ;
        RECT 49.185 198.275 49.355 199.055 ;
        RECT 51.045 198.885 51.215 199.575 ;
        RECT 49.715 198.715 51.215 198.885 ;
        RECT 51.405 198.915 51.615 199.705 ;
        RECT 51.785 199.085 52.135 199.705 ;
        RECT 52.305 199.095 52.475 199.875 ;
        RECT 53.005 199.715 53.175 199.945 ;
        RECT 52.645 199.545 53.175 199.715 ;
        RECT 52.645 199.265 52.865 199.545 ;
        RECT 53.345 199.375 53.585 199.775 ;
        RECT 52.305 198.925 52.710 199.095 ;
        RECT 53.045 199.005 53.585 199.375 ;
        RECT 53.755 199.590 54.075 199.945 ;
        RECT 54.320 199.865 54.625 200.325 ;
        RECT 54.795 199.615 55.050 200.145 ;
        RECT 56.150 199.780 61.495 200.325 ;
        RECT 53.755 199.415 54.080 199.590 ;
        RECT 53.755 199.115 54.670 199.415 ;
        RECT 53.930 199.085 54.670 199.115 ;
        RECT 51.405 198.755 52.080 198.915 ;
        RECT 52.540 198.835 52.710 198.925 ;
        RECT 51.405 198.745 52.370 198.755 ;
        RECT 51.045 198.575 51.215 198.715 ;
        RECT 47.790 197.775 48.040 198.235 ;
        RECT 48.210 197.945 48.460 198.275 ;
        RECT 48.675 197.945 49.355 198.275 ;
        RECT 49.525 198.375 50.600 198.545 ;
        RECT 51.045 198.405 51.605 198.575 ;
        RECT 51.910 198.455 52.370 198.745 ;
        RECT 52.540 198.665 53.760 198.835 ;
        RECT 49.525 198.035 49.695 198.375 ;
        RECT 49.930 197.775 50.260 198.205 ;
        RECT 50.430 198.035 50.600 198.375 ;
        RECT 50.895 197.775 51.265 198.235 ;
        RECT 51.435 197.945 51.605 198.405 ;
        RECT 52.540 198.285 52.710 198.665 ;
        RECT 53.930 198.495 54.100 199.085 ;
        RECT 54.840 198.965 55.050 199.615 ;
        RECT 51.840 197.945 52.710 198.285 ;
        RECT 53.300 198.325 54.100 198.495 ;
        RECT 52.880 197.775 53.130 198.235 ;
        RECT 53.300 198.035 53.470 198.325 ;
        RECT 53.650 197.775 53.980 198.155 ;
        RECT 54.320 197.775 54.625 198.915 ;
        RECT 54.795 198.085 55.050 198.965 ;
        RECT 57.740 198.210 58.090 199.460 ;
        RECT 59.570 198.950 59.910 199.780 ;
        RECT 61.725 199.505 61.935 200.325 ;
        RECT 62.105 199.525 62.435 200.155 ;
        RECT 62.105 198.925 62.355 199.525 ;
        RECT 62.605 199.505 62.835 200.325 ;
        RECT 63.045 199.600 63.335 200.325 ;
        RECT 63.510 199.775 63.765 200.065 ;
        RECT 63.935 199.945 64.265 200.325 ;
        RECT 63.510 199.605 64.260 199.775 ;
        RECT 62.525 199.085 62.855 199.335 ;
        RECT 56.150 197.775 61.495 198.210 ;
        RECT 61.725 197.775 61.935 198.915 ;
        RECT 62.105 197.945 62.435 198.925 ;
        RECT 62.605 197.775 62.835 198.915 ;
        RECT 63.045 197.775 63.335 198.940 ;
        RECT 63.510 198.785 63.860 199.435 ;
        RECT 64.030 198.615 64.260 199.605 ;
        RECT 63.510 198.445 64.260 198.615 ;
        RECT 63.510 197.945 63.765 198.445 ;
        RECT 63.935 197.775 64.265 198.275 ;
        RECT 64.435 197.945 64.605 200.065 ;
        RECT 64.965 199.965 65.295 200.325 ;
        RECT 65.465 199.935 65.960 200.105 ;
        RECT 66.165 199.935 67.020 200.105 ;
        RECT 64.835 198.745 65.295 199.795 ;
        RECT 64.775 197.960 65.100 198.745 ;
        RECT 65.465 198.575 65.635 199.935 ;
        RECT 65.805 199.025 66.155 199.645 ;
        RECT 66.325 199.425 66.680 199.645 ;
        RECT 66.325 198.835 66.495 199.425 ;
        RECT 66.850 199.225 67.020 199.935 ;
        RECT 67.895 199.865 68.225 200.325 ;
        RECT 68.435 199.965 68.785 200.135 ;
        RECT 67.225 199.395 68.015 199.645 ;
        RECT 68.435 199.575 68.695 199.965 ;
        RECT 69.005 199.875 69.955 200.155 ;
        RECT 70.125 199.885 70.315 200.325 ;
        RECT 70.485 199.945 71.555 200.115 ;
        RECT 68.185 199.225 68.355 199.405 ;
        RECT 65.465 198.405 65.860 198.575 ;
        RECT 66.030 198.445 66.495 198.835 ;
        RECT 66.665 199.055 68.355 199.225 ;
        RECT 65.690 198.275 65.860 198.405 ;
        RECT 66.665 198.275 66.835 199.055 ;
        RECT 68.525 198.885 68.695 199.575 ;
        RECT 67.195 198.715 68.695 198.885 ;
        RECT 68.885 198.915 69.095 199.705 ;
        RECT 69.265 199.085 69.615 199.705 ;
        RECT 69.785 199.095 69.955 199.875 ;
        RECT 70.485 199.715 70.655 199.945 ;
        RECT 70.125 199.545 70.655 199.715 ;
        RECT 70.125 199.265 70.345 199.545 ;
        RECT 70.825 199.375 71.065 199.775 ;
        RECT 69.785 198.925 70.190 199.095 ;
        RECT 70.525 199.005 71.065 199.375 ;
        RECT 71.235 199.590 71.555 199.945 ;
        RECT 71.800 199.865 72.105 200.325 ;
        RECT 72.275 199.615 72.525 200.145 ;
        RECT 71.235 199.415 71.560 199.590 ;
        RECT 71.235 199.115 72.150 199.415 ;
        RECT 71.410 199.085 72.150 199.115 ;
        RECT 68.885 198.755 69.560 198.915 ;
        RECT 70.020 198.835 70.190 198.925 ;
        RECT 68.885 198.745 69.850 198.755 ;
        RECT 68.525 198.575 68.695 198.715 ;
        RECT 65.270 197.775 65.520 198.235 ;
        RECT 65.690 197.945 65.940 198.275 ;
        RECT 66.155 197.945 66.835 198.275 ;
        RECT 67.005 198.375 68.080 198.545 ;
        RECT 68.525 198.405 69.085 198.575 ;
        RECT 69.390 198.455 69.850 198.745 ;
        RECT 70.020 198.665 71.240 198.835 ;
        RECT 67.005 198.035 67.175 198.375 ;
        RECT 67.410 197.775 67.740 198.205 ;
        RECT 67.910 198.035 68.080 198.375 ;
        RECT 68.375 197.775 68.745 198.235 ;
        RECT 68.915 197.945 69.085 198.405 ;
        RECT 70.020 198.285 70.190 198.665 ;
        RECT 71.410 198.495 71.580 199.085 ;
        RECT 72.320 198.965 72.525 199.615 ;
        RECT 72.695 199.570 72.945 200.325 ;
        RECT 73.165 199.650 73.440 199.995 ;
        RECT 73.630 199.925 74.005 200.325 ;
        RECT 74.175 199.755 74.345 200.105 ;
        RECT 74.515 199.925 74.845 200.325 ;
        RECT 75.015 199.755 75.275 200.155 ;
        RECT 69.320 197.945 70.190 198.285 ;
        RECT 70.780 198.325 71.580 198.495 ;
        RECT 70.360 197.775 70.610 198.235 ;
        RECT 70.780 198.035 70.950 198.325 ;
        RECT 71.130 197.775 71.460 198.155 ;
        RECT 71.800 197.775 72.105 198.915 ;
        RECT 72.275 198.085 72.525 198.965 ;
        RECT 73.165 198.915 73.335 199.650 ;
        RECT 73.610 199.585 75.275 199.755 ;
        RECT 73.610 199.415 73.780 199.585 ;
        RECT 75.455 199.505 75.785 199.925 ;
        RECT 75.955 199.505 76.215 200.325 ;
        RECT 76.845 199.555 78.515 200.325 ;
        RECT 75.455 199.415 75.705 199.505 ;
        RECT 73.505 199.085 73.780 199.415 ;
        RECT 73.950 199.085 74.775 199.415 ;
        RECT 74.990 199.085 75.705 199.415 ;
        RECT 75.875 199.085 76.210 199.335 ;
        RECT 73.610 198.915 73.780 199.085 ;
        RECT 72.695 197.775 72.945 198.915 ;
        RECT 73.165 197.945 73.440 198.915 ;
        RECT 73.610 198.745 74.270 198.915 ;
        RECT 74.530 198.795 74.775 199.085 ;
        RECT 74.100 198.625 74.270 198.745 ;
        RECT 74.945 198.625 75.275 198.915 ;
        RECT 73.650 197.775 73.930 198.575 ;
        RECT 74.100 198.455 75.275 198.625 ;
        RECT 75.535 198.525 75.705 199.085 ;
        RECT 74.100 197.955 75.715 198.285 ;
        RECT 75.955 197.775 76.215 198.915 ;
        RECT 76.845 198.865 77.595 199.385 ;
        RECT 77.765 199.035 78.515 199.555 ;
        RECT 78.725 199.505 78.955 200.325 ;
        RECT 79.125 199.525 79.455 200.155 ;
        RECT 78.705 199.085 79.035 199.335 ;
        RECT 79.205 198.925 79.455 199.525 ;
        RECT 79.625 199.505 79.835 200.325 ;
        RECT 80.065 199.585 80.530 200.130 ;
        RECT 76.845 197.775 78.515 198.865 ;
        RECT 78.725 197.775 78.955 198.915 ;
        RECT 79.125 197.945 79.455 198.925 ;
        RECT 79.625 197.775 79.835 198.915 ;
        RECT 80.065 198.625 80.235 199.585 ;
        RECT 81.035 199.505 81.205 200.325 ;
        RECT 81.375 199.675 81.705 200.155 ;
        RECT 81.875 199.935 82.225 200.325 ;
        RECT 82.395 199.755 82.625 200.155 ;
        RECT 82.115 199.675 82.625 199.755 ;
        RECT 81.375 199.585 82.625 199.675 ;
        RECT 82.795 199.585 83.115 200.065 ;
        RECT 83.290 199.780 88.635 200.325 ;
        RECT 81.375 199.505 82.285 199.585 ;
        RECT 80.405 198.965 80.650 199.415 ;
        RECT 80.910 199.135 81.605 199.335 ;
        RECT 81.775 199.165 82.375 199.335 ;
        RECT 81.775 198.965 81.945 199.165 ;
        RECT 82.605 198.995 82.775 199.415 ;
        RECT 80.405 198.795 81.945 198.965 ;
        RECT 82.115 198.825 82.775 198.995 ;
        RECT 82.115 198.625 82.285 198.825 ;
        RECT 82.945 198.655 83.115 199.585 ;
        RECT 80.065 198.455 82.285 198.625 ;
        RECT 82.455 198.455 83.115 198.655 ;
        RECT 80.065 197.775 80.365 198.285 ;
        RECT 80.535 197.945 80.865 198.455 ;
        RECT 82.455 198.285 82.625 198.455 ;
        RECT 81.035 197.775 81.665 198.285 ;
        RECT 82.245 198.115 82.625 198.285 ;
        RECT 82.795 197.775 83.095 198.285 ;
        RECT 84.880 198.210 85.230 199.460 ;
        RECT 86.710 198.950 87.050 199.780 ;
        RECT 88.805 199.600 89.095 200.325 ;
        RECT 89.265 199.555 92.775 200.325 ;
        RECT 92.950 199.780 98.295 200.325 ;
        RECT 83.290 197.775 88.635 198.210 ;
        RECT 88.805 197.775 89.095 198.940 ;
        RECT 89.265 198.865 90.955 199.385 ;
        RECT 91.125 199.035 92.775 199.555 ;
        RECT 89.265 197.775 92.775 198.865 ;
        RECT 94.540 198.210 94.890 199.460 ;
        RECT 96.370 198.950 96.710 199.780 ;
        RECT 98.470 199.615 98.725 200.145 ;
        RECT 98.895 199.865 99.200 200.325 ;
        RECT 99.445 199.945 100.515 200.115 ;
        RECT 98.470 198.965 98.680 199.615 ;
        RECT 99.445 199.590 99.765 199.945 ;
        RECT 99.440 199.415 99.765 199.590 ;
        RECT 98.850 199.115 99.765 199.415 ;
        RECT 99.935 199.375 100.175 199.775 ;
        RECT 100.345 199.715 100.515 199.945 ;
        RECT 100.685 199.885 100.875 200.325 ;
        RECT 101.045 199.875 101.995 200.155 ;
        RECT 102.215 199.965 102.565 200.135 ;
        RECT 100.345 199.545 100.875 199.715 ;
        RECT 98.850 199.085 99.590 199.115 ;
        RECT 92.950 197.775 98.295 198.210 ;
        RECT 98.470 198.085 98.725 198.965 ;
        RECT 98.895 197.775 99.200 198.915 ;
        RECT 99.420 198.495 99.590 199.085 ;
        RECT 99.935 199.005 100.475 199.375 ;
        RECT 100.655 199.265 100.875 199.545 ;
        RECT 101.045 199.095 101.215 199.875 ;
        RECT 100.810 198.925 101.215 199.095 ;
        RECT 101.385 199.085 101.735 199.705 ;
        RECT 100.810 198.835 100.980 198.925 ;
        RECT 101.905 198.915 102.115 199.705 ;
        RECT 99.760 198.665 100.980 198.835 ;
        RECT 101.440 198.755 102.115 198.915 ;
        RECT 99.420 198.325 100.220 198.495 ;
        RECT 99.540 197.775 99.870 198.155 ;
        RECT 100.050 198.035 100.220 198.325 ;
        RECT 100.810 198.285 100.980 198.665 ;
        RECT 101.150 198.745 102.115 198.755 ;
        RECT 102.305 199.575 102.565 199.965 ;
        RECT 102.775 199.865 103.105 200.325 ;
        RECT 103.980 199.935 104.835 200.105 ;
        RECT 105.040 199.935 105.535 200.105 ;
        RECT 105.705 199.965 106.035 200.325 ;
        RECT 102.305 198.885 102.475 199.575 ;
        RECT 102.645 199.225 102.815 199.405 ;
        RECT 102.985 199.395 103.775 199.645 ;
        RECT 103.980 199.225 104.150 199.935 ;
        RECT 104.320 199.425 104.675 199.645 ;
        RECT 102.645 199.055 104.335 199.225 ;
        RECT 101.150 198.455 101.610 198.745 ;
        RECT 102.305 198.715 103.805 198.885 ;
        RECT 102.305 198.575 102.475 198.715 ;
        RECT 101.915 198.405 102.475 198.575 ;
        RECT 100.390 197.775 100.640 198.235 ;
        RECT 100.810 197.945 101.680 198.285 ;
        RECT 101.915 197.945 102.085 198.405 ;
        RECT 102.920 198.375 103.995 198.545 ;
        RECT 102.255 197.775 102.625 198.235 ;
        RECT 102.920 198.035 103.090 198.375 ;
        RECT 103.260 197.775 103.590 198.205 ;
        RECT 103.825 198.035 103.995 198.375 ;
        RECT 104.165 198.275 104.335 199.055 ;
        RECT 104.505 198.835 104.675 199.425 ;
        RECT 104.845 199.025 105.195 199.645 ;
        RECT 104.505 198.445 104.970 198.835 ;
        RECT 105.365 198.575 105.535 199.935 ;
        RECT 105.705 198.745 106.165 199.795 ;
        RECT 105.140 198.405 105.535 198.575 ;
        RECT 105.140 198.275 105.310 198.405 ;
        RECT 104.165 197.945 104.845 198.275 ;
        RECT 105.060 197.945 105.310 198.275 ;
        RECT 105.480 197.775 105.730 198.235 ;
        RECT 105.900 197.960 106.225 198.745 ;
        RECT 106.395 197.945 106.565 200.065 ;
        RECT 106.735 199.945 107.065 200.325 ;
        RECT 107.235 199.775 107.490 200.065 ;
        RECT 106.740 199.605 107.490 199.775 ;
        RECT 106.740 198.615 106.970 199.605 ;
        RECT 107.665 199.555 110.255 200.325 ;
        RECT 107.140 198.785 107.490 199.435 ;
        RECT 107.665 198.865 108.875 199.385 ;
        RECT 109.045 199.035 110.255 199.555 ;
        RECT 110.700 199.515 110.945 200.120 ;
        RECT 111.165 199.790 111.675 200.325 ;
        RECT 110.425 199.345 111.655 199.515 ;
        RECT 106.740 198.445 107.490 198.615 ;
        RECT 106.735 197.775 107.065 198.275 ;
        RECT 107.235 197.945 107.490 198.445 ;
        RECT 107.665 197.775 110.255 198.865 ;
        RECT 110.425 198.535 110.765 199.345 ;
        RECT 110.935 198.780 111.685 198.970 ;
        RECT 110.425 198.125 110.940 198.535 ;
        RECT 111.175 197.775 111.345 198.535 ;
        RECT 111.515 198.115 111.685 198.780 ;
        RECT 111.855 198.795 112.045 200.155 ;
        RECT 112.215 199.645 112.490 200.155 ;
        RECT 112.680 199.790 113.210 200.155 ;
        RECT 113.635 199.925 113.965 200.325 ;
        RECT 113.035 199.755 113.210 199.790 ;
        RECT 112.215 199.475 112.495 199.645 ;
        RECT 112.215 198.995 112.490 199.475 ;
        RECT 112.695 198.795 112.865 199.595 ;
        RECT 111.855 198.625 112.865 198.795 ;
        RECT 113.035 199.585 113.965 199.755 ;
        RECT 114.135 199.585 114.390 200.155 ;
        RECT 114.565 199.600 114.855 200.325 ;
        RECT 115.030 199.615 115.285 200.145 ;
        RECT 115.455 199.865 115.760 200.325 ;
        RECT 116.005 199.945 117.075 200.115 ;
        RECT 113.035 198.455 113.205 199.585 ;
        RECT 113.795 199.415 113.965 199.585 ;
        RECT 112.080 198.285 113.205 198.455 ;
        RECT 113.375 199.085 113.570 199.415 ;
        RECT 113.795 199.085 114.050 199.415 ;
        RECT 113.375 198.115 113.545 199.085 ;
        RECT 114.220 198.915 114.390 199.585 ;
        RECT 115.030 198.965 115.240 199.615 ;
        RECT 116.005 199.590 116.325 199.945 ;
        RECT 116.000 199.415 116.325 199.590 ;
        RECT 115.410 199.115 116.325 199.415 ;
        RECT 116.495 199.375 116.735 199.775 ;
        RECT 116.905 199.715 117.075 199.945 ;
        RECT 117.245 199.885 117.435 200.325 ;
        RECT 117.605 199.875 118.555 200.155 ;
        RECT 118.775 199.965 119.125 200.135 ;
        RECT 116.905 199.545 117.435 199.715 ;
        RECT 115.410 199.085 116.150 199.115 ;
        RECT 111.515 197.945 113.545 198.115 ;
        RECT 113.715 197.775 113.885 198.915 ;
        RECT 114.055 197.945 114.390 198.915 ;
        RECT 114.565 197.775 114.855 198.940 ;
        RECT 115.030 198.085 115.285 198.965 ;
        RECT 115.455 197.775 115.760 198.915 ;
        RECT 115.980 198.495 116.150 199.085 ;
        RECT 116.495 199.005 117.035 199.375 ;
        RECT 117.215 199.265 117.435 199.545 ;
        RECT 117.605 199.095 117.775 199.875 ;
        RECT 117.370 198.925 117.775 199.095 ;
        RECT 117.945 199.085 118.295 199.705 ;
        RECT 117.370 198.835 117.540 198.925 ;
        RECT 118.465 198.915 118.675 199.705 ;
        RECT 116.320 198.665 117.540 198.835 ;
        RECT 118.000 198.755 118.675 198.915 ;
        RECT 115.980 198.325 116.780 198.495 ;
        RECT 116.100 197.775 116.430 198.155 ;
        RECT 116.610 198.035 116.780 198.325 ;
        RECT 117.370 198.285 117.540 198.665 ;
        RECT 117.710 198.745 118.675 198.755 ;
        RECT 118.865 199.575 119.125 199.965 ;
        RECT 119.335 199.865 119.665 200.325 ;
        RECT 120.540 199.935 121.395 200.105 ;
        RECT 121.600 199.935 122.095 200.105 ;
        RECT 122.265 199.965 122.595 200.325 ;
        RECT 118.865 198.885 119.035 199.575 ;
        RECT 119.205 199.225 119.375 199.405 ;
        RECT 119.545 199.395 120.335 199.645 ;
        RECT 120.540 199.225 120.710 199.935 ;
        RECT 120.880 199.425 121.235 199.645 ;
        RECT 119.205 199.055 120.895 199.225 ;
        RECT 117.710 198.455 118.170 198.745 ;
        RECT 118.865 198.715 120.365 198.885 ;
        RECT 118.865 198.575 119.035 198.715 ;
        RECT 118.475 198.405 119.035 198.575 ;
        RECT 116.950 197.775 117.200 198.235 ;
        RECT 117.370 197.945 118.240 198.285 ;
        RECT 118.475 197.945 118.645 198.405 ;
        RECT 119.480 198.375 120.555 198.545 ;
        RECT 118.815 197.775 119.185 198.235 ;
        RECT 119.480 198.035 119.650 198.375 ;
        RECT 119.820 197.775 120.150 198.205 ;
        RECT 120.385 198.035 120.555 198.375 ;
        RECT 120.725 198.275 120.895 199.055 ;
        RECT 121.065 198.835 121.235 199.425 ;
        RECT 121.405 199.025 121.755 199.645 ;
        RECT 121.065 198.445 121.530 198.835 ;
        RECT 121.925 198.575 122.095 199.935 ;
        RECT 122.265 198.745 122.725 199.795 ;
        RECT 121.700 198.405 122.095 198.575 ;
        RECT 121.700 198.275 121.870 198.405 ;
        RECT 120.725 197.945 121.405 198.275 ;
        RECT 121.620 197.945 121.870 198.275 ;
        RECT 122.040 197.775 122.290 198.235 ;
        RECT 122.460 197.960 122.785 198.745 ;
        RECT 122.955 197.945 123.125 200.065 ;
        RECT 123.295 199.945 123.625 200.325 ;
        RECT 123.795 199.775 124.050 200.065 ;
        RECT 123.300 199.605 124.050 199.775 ;
        RECT 123.300 198.615 123.530 199.605 ;
        RECT 124.685 199.555 126.355 200.325 ;
        RECT 126.525 199.575 127.735 200.325 ;
        RECT 123.700 198.785 124.050 199.435 ;
        RECT 124.685 198.865 125.435 199.385 ;
        RECT 125.605 199.035 126.355 199.555 ;
        RECT 126.525 198.865 127.045 199.405 ;
        RECT 127.215 199.035 127.735 199.575 ;
        RECT 123.300 198.445 124.050 198.615 ;
        RECT 123.295 197.775 123.625 198.275 ;
        RECT 123.795 197.945 124.050 198.445 ;
        RECT 124.685 197.775 126.355 198.865 ;
        RECT 126.525 197.775 127.735 198.865 ;
        RECT 20.640 197.605 127.820 197.775 ;
        RECT 20.725 196.515 21.935 197.605 ;
        RECT 20.725 195.805 21.245 196.345 ;
        RECT 21.415 195.975 21.935 196.515 ;
        RECT 22.565 196.515 24.235 197.605 ;
        RECT 22.565 195.995 23.315 196.515 ;
        RECT 24.405 196.440 24.695 197.605 ;
        RECT 25.325 196.515 27.915 197.605 ;
        RECT 28.090 197.170 33.435 197.605 ;
        RECT 23.485 195.825 24.235 196.345 ;
        RECT 25.325 195.995 26.535 196.515 ;
        RECT 26.705 195.825 27.915 196.345 ;
        RECT 29.680 195.920 30.030 197.170 ;
        RECT 33.665 196.465 33.875 197.605 ;
        RECT 34.045 196.455 34.375 197.435 ;
        RECT 34.545 196.465 34.775 197.605 ;
        RECT 34.985 196.515 36.655 197.605 ;
        RECT 36.830 197.170 42.175 197.605 ;
        RECT 20.725 195.055 21.935 195.805 ;
        RECT 22.565 195.055 24.235 195.825 ;
        RECT 24.405 195.055 24.695 195.780 ;
        RECT 25.325 195.055 27.915 195.825 ;
        RECT 31.510 195.600 31.850 196.430 ;
        RECT 28.090 195.055 33.435 195.600 ;
        RECT 33.665 195.055 33.875 195.875 ;
        RECT 34.045 195.855 34.295 196.455 ;
        RECT 34.465 196.045 34.795 196.295 ;
        RECT 34.985 195.995 35.735 196.515 ;
        RECT 34.045 195.225 34.375 195.855 ;
        RECT 34.545 195.055 34.775 195.875 ;
        RECT 35.905 195.825 36.655 196.345 ;
        RECT 38.420 195.920 38.770 197.170 ;
        RECT 42.385 196.465 42.615 197.605 ;
        RECT 42.785 196.455 43.115 197.435 ;
        RECT 43.285 196.465 43.495 197.605 ;
        RECT 43.725 196.515 45.395 197.605 ;
        RECT 45.565 196.845 46.080 197.255 ;
        RECT 46.315 196.845 46.485 197.605 ;
        RECT 46.655 197.265 48.685 197.435 ;
        RECT 34.985 195.055 36.655 195.825 ;
        RECT 40.250 195.600 40.590 196.430 ;
        RECT 42.365 196.045 42.695 196.295 ;
        RECT 36.830 195.055 42.175 195.600 ;
        RECT 42.385 195.055 42.615 195.875 ;
        RECT 42.865 195.855 43.115 196.455 ;
        RECT 43.725 195.995 44.475 196.515 ;
        RECT 42.785 195.225 43.115 195.855 ;
        RECT 43.285 195.055 43.495 195.875 ;
        RECT 44.645 195.825 45.395 196.345 ;
        RECT 45.565 196.035 45.905 196.845 ;
        RECT 46.655 196.600 46.825 197.265 ;
        RECT 47.220 196.925 48.345 197.095 ;
        RECT 46.075 196.410 46.825 196.600 ;
        RECT 46.995 196.585 48.005 196.755 ;
        RECT 45.565 195.865 46.795 196.035 ;
        RECT 43.725 195.055 45.395 195.825 ;
        RECT 45.840 195.260 46.085 195.865 ;
        RECT 46.305 195.055 46.815 195.590 ;
        RECT 46.995 195.225 47.185 196.585 ;
        RECT 47.355 195.565 47.630 196.385 ;
        RECT 47.835 195.785 48.005 196.585 ;
        RECT 48.175 195.795 48.345 196.925 ;
        RECT 48.515 196.295 48.685 197.265 ;
        RECT 48.855 196.465 49.025 197.605 ;
        RECT 49.195 196.465 49.530 197.435 ;
        RECT 48.515 195.965 48.710 196.295 ;
        RECT 48.935 195.965 49.190 196.295 ;
        RECT 48.935 195.795 49.105 195.965 ;
        RECT 49.360 195.795 49.530 196.465 ;
        RECT 50.165 196.440 50.455 197.605 ;
        RECT 51.545 196.515 55.055 197.605 ;
        RECT 55.225 196.845 55.740 197.255 ;
        RECT 55.975 196.845 56.145 197.605 ;
        RECT 56.315 197.265 58.345 197.435 ;
        RECT 51.545 195.995 53.235 196.515 ;
        RECT 53.405 195.825 55.055 196.345 ;
        RECT 55.225 196.035 55.565 196.845 ;
        RECT 56.315 196.600 56.485 197.265 ;
        RECT 56.880 196.925 58.005 197.095 ;
        RECT 55.735 196.410 56.485 196.600 ;
        RECT 56.655 196.585 57.665 196.755 ;
        RECT 55.225 195.865 56.455 196.035 ;
        RECT 48.175 195.625 49.105 195.795 ;
        RECT 48.175 195.590 48.350 195.625 ;
        RECT 47.355 195.395 47.635 195.565 ;
        RECT 47.355 195.225 47.630 195.395 ;
        RECT 47.820 195.225 48.350 195.590 ;
        RECT 48.775 195.055 49.105 195.455 ;
        RECT 49.275 195.225 49.530 195.795 ;
        RECT 50.165 195.055 50.455 195.780 ;
        RECT 51.545 195.055 55.055 195.825 ;
        RECT 55.500 195.260 55.745 195.865 ;
        RECT 55.965 195.055 56.475 195.590 ;
        RECT 56.655 195.225 56.845 196.585 ;
        RECT 57.015 195.905 57.290 196.385 ;
        RECT 57.015 195.735 57.295 195.905 ;
        RECT 57.495 195.785 57.665 196.585 ;
        RECT 57.835 195.795 58.005 196.925 ;
        RECT 58.175 196.295 58.345 197.265 ;
        RECT 58.515 196.465 58.685 197.605 ;
        RECT 58.855 196.465 59.190 197.435 ;
        RECT 59.915 196.675 60.085 197.435 ;
        RECT 60.265 196.845 60.595 197.605 ;
        RECT 59.915 196.505 60.580 196.675 ;
        RECT 60.765 196.530 61.035 197.435 ;
        RECT 61.210 197.170 66.555 197.605 ;
        RECT 58.175 195.965 58.370 196.295 ;
        RECT 58.595 195.965 58.850 196.295 ;
        RECT 58.595 195.795 58.765 195.965 ;
        RECT 59.020 195.795 59.190 196.465 ;
        RECT 60.410 196.360 60.580 196.505 ;
        RECT 59.845 195.955 60.175 196.325 ;
        RECT 60.410 196.030 60.695 196.360 ;
        RECT 57.015 195.225 57.290 195.735 ;
        RECT 57.835 195.625 58.765 195.795 ;
        RECT 57.835 195.590 58.010 195.625 ;
        RECT 57.480 195.225 58.010 195.590 ;
        RECT 58.435 195.055 58.765 195.455 ;
        RECT 58.935 195.225 59.190 195.795 ;
        RECT 60.410 195.775 60.580 196.030 ;
        RECT 59.915 195.605 60.580 195.775 ;
        RECT 60.865 195.730 61.035 196.530 ;
        RECT 62.800 195.920 63.150 197.170 ;
        RECT 66.765 196.465 66.995 197.605 ;
        RECT 67.165 196.455 67.495 197.435 ;
        RECT 67.665 196.465 67.875 197.605 ;
        RECT 69.025 197.050 69.630 197.605 ;
        RECT 69.805 197.095 70.285 197.435 ;
        RECT 70.455 197.060 70.710 197.605 ;
        RECT 69.025 196.950 69.640 197.050 ;
        RECT 69.455 196.925 69.640 196.950 ;
        RECT 59.915 195.225 60.085 195.605 ;
        RECT 60.265 195.055 60.595 195.435 ;
        RECT 60.775 195.225 61.035 195.730 ;
        RECT 64.630 195.600 64.970 196.430 ;
        RECT 66.745 196.045 67.075 196.295 ;
        RECT 61.210 195.055 66.555 195.600 ;
        RECT 66.765 195.055 66.995 195.875 ;
        RECT 67.245 195.855 67.495 196.455 ;
        RECT 69.025 196.330 69.285 196.780 ;
        RECT 69.455 196.680 69.785 196.925 ;
        RECT 69.955 196.605 70.710 196.855 ;
        RECT 70.880 196.735 71.155 197.435 ;
        RECT 69.940 196.570 70.710 196.605 ;
        RECT 69.925 196.560 70.710 196.570 ;
        RECT 69.920 196.545 70.815 196.560 ;
        RECT 69.900 196.530 70.815 196.545 ;
        RECT 69.880 196.520 70.815 196.530 ;
        RECT 69.855 196.510 70.815 196.520 ;
        RECT 69.785 196.480 70.815 196.510 ;
        RECT 69.765 196.450 70.815 196.480 ;
        RECT 69.745 196.420 70.815 196.450 ;
        RECT 69.715 196.395 70.815 196.420 ;
        RECT 69.680 196.360 70.815 196.395 ;
        RECT 69.650 196.355 70.815 196.360 ;
        RECT 69.650 196.350 70.040 196.355 ;
        RECT 69.650 196.340 70.015 196.350 ;
        RECT 69.650 196.335 70.000 196.340 ;
        RECT 69.650 196.330 69.985 196.335 ;
        RECT 69.025 196.325 69.985 196.330 ;
        RECT 69.025 196.315 69.975 196.325 ;
        RECT 69.025 196.310 69.965 196.315 ;
        RECT 69.025 196.300 69.955 196.310 ;
        RECT 69.025 196.290 69.950 196.300 ;
        RECT 69.025 196.285 69.945 196.290 ;
        RECT 69.025 196.270 69.935 196.285 ;
        RECT 69.025 196.255 69.930 196.270 ;
        RECT 69.025 196.230 69.920 196.255 ;
        RECT 69.025 196.160 69.915 196.230 ;
        RECT 67.165 195.225 67.495 195.855 ;
        RECT 67.665 195.055 67.875 195.875 ;
        RECT 69.025 195.605 69.575 195.990 ;
        RECT 69.745 195.435 69.915 196.160 ;
        RECT 69.025 195.265 69.915 195.435 ;
        RECT 70.085 195.760 70.415 196.185 ;
        RECT 70.585 195.960 70.815 196.355 ;
        RECT 70.085 195.735 70.335 195.760 ;
        RECT 70.085 195.275 70.305 195.735 ;
        RECT 70.985 195.705 71.155 196.735 ;
        RECT 70.475 195.055 70.725 195.595 ;
        RECT 70.895 195.225 71.155 195.705 ;
        RECT 71.335 196.545 71.665 197.395 ;
        RECT 71.335 195.780 71.525 196.545 ;
        RECT 71.835 196.465 72.085 197.605 ;
        RECT 72.275 196.965 72.525 197.385 ;
        RECT 72.755 197.135 73.085 197.605 ;
        RECT 73.315 196.965 73.565 197.385 ;
        RECT 72.275 196.795 73.565 196.965 ;
        RECT 73.745 196.965 74.075 197.395 ;
        RECT 73.745 196.795 74.200 196.965 ;
        RECT 72.265 196.295 72.480 196.625 ;
        RECT 71.695 195.965 72.005 196.295 ;
        RECT 72.175 195.965 72.480 196.295 ;
        RECT 72.655 195.965 72.940 196.625 ;
        RECT 73.135 195.965 73.400 196.625 ;
        RECT 73.615 195.965 73.860 196.625 ;
        RECT 71.835 195.795 72.005 195.965 ;
        RECT 74.030 195.795 74.200 196.795 ;
        RECT 74.545 196.515 75.755 197.605 ;
        RECT 74.545 195.975 75.065 196.515 ;
        RECT 75.925 196.440 76.215 197.605 ;
        RECT 77.310 196.415 77.565 197.295 ;
        RECT 77.735 196.465 78.040 197.605 ;
        RECT 78.380 197.225 78.710 197.605 ;
        RECT 78.890 197.055 79.060 197.345 ;
        RECT 79.230 197.145 79.480 197.605 ;
        RECT 78.260 196.885 79.060 197.055 ;
        RECT 79.650 197.095 80.520 197.435 ;
        RECT 75.235 195.805 75.755 196.345 ;
        RECT 71.335 195.270 71.665 195.780 ;
        RECT 71.835 195.625 74.200 195.795 ;
        RECT 71.835 195.055 72.165 195.455 ;
        RECT 73.215 195.285 73.545 195.625 ;
        RECT 73.715 195.055 74.045 195.455 ;
        RECT 74.545 195.055 75.755 195.805 ;
        RECT 75.925 195.055 76.215 195.780 ;
        RECT 77.310 195.765 77.520 196.415 ;
        RECT 78.260 196.295 78.430 196.885 ;
        RECT 79.650 196.715 79.820 197.095 ;
        RECT 80.755 196.975 80.925 197.435 ;
        RECT 81.095 197.145 81.465 197.605 ;
        RECT 81.760 197.005 81.930 197.345 ;
        RECT 82.100 197.175 82.430 197.605 ;
        RECT 82.665 197.005 82.835 197.345 ;
        RECT 78.600 196.545 79.820 196.715 ;
        RECT 79.990 196.635 80.450 196.925 ;
        RECT 80.755 196.805 81.315 196.975 ;
        RECT 81.760 196.835 82.835 197.005 ;
        RECT 83.005 197.105 83.685 197.435 ;
        RECT 83.900 197.105 84.150 197.435 ;
        RECT 84.320 197.145 84.570 197.605 ;
        RECT 81.145 196.665 81.315 196.805 ;
        RECT 79.990 196.625 80.955 196.635 ;
        RECT 79.650 196.455 79.820 196.545 ;
        RECT 80.280 196.465 80.955 196.625 ;
        RECT 77.690 196.265 78.430 196.295 ;
        RECT 77.690 195.965 78.605 196.265 ;
        RECT 78.280 195.790 78.605 195.965 ;
        RECT 77.310 195.235 77.565 195.765 ;
        RECT 77.735 195.055 78.040 195.515 ;
        RECT 78.285 195.435 78.605 195.790 ;
        RECT 78.775 196.005 79.315 196.375 ;
        RECT 79.650 196.285 80.055 196.455 ;
        RECT 78.775 195.605 79.015 196.005 ;
        RECT 79.495 195.835 79.715 196.115 ;
        RECT 79.185 195.665 79.715 195.835 ;
        RECT 79.185 195.435 79.355 195.665 ;
        RECT 79.885 195.505 80.055 196.285 ;
        RECT 80.225 195.675 80.575 196.295 ;
        RECT 80.745 195.675 80.955 196.465 ;
        RECT 81.145 196.495 82.645 196.665 ;
        RECT 81.145 195.805 81.315 196.495 ;
        RECT 83.005 196.325 83.175 197.105 ;
        RECT 83.980 196.975 84.150 197.105 ;
        RECT 81.485 196.155 83.175 196.325 ;
        RECT 83.345 196.545 83.810 196.935 ;
        RECT 83.980 196.805 84.375 196.975 ;
        RECT 81.485 195.975 81.655 196.155 ;
        RECT 78.285 195.265 79.355 195.435 ;
        RECT 79.525 195.055 79.715 195.495 ;
        RECT 79.885 195.225 80.835 195.505 ;
        RECT 81.145 195.415 81.405 195.805 ;
        RECT 81.825 195.735 82.615 195.985 ;
        RECT 81.055 195.245 81.405 195.415 ;
        RECT 81.615 195.055 81.945 195.515 ;
        RECT 82.820 195.445 82.990 196.155 ;
        RECT 83.345 195.955 83.515 196.545 ;
        RECT 83.160 195.735 83.515 195.955 ;
        RECT 83.685 195.735 84.035 196.355 ;
        RECT 84.205 195.445 84.375 196.805 ;
        RECT 84.740 196.635 85.065 197.420 ;
        RECT 84.545 195.585 85.005 196.635 ;
        RECT 82.820 195.275 83.675 195.445 ;
        RECT 83.880 195.275 84.375 195.445 ;
        RECT 84.545 195.055 84.875 195.415 ;
        RECT 85.235 195.315 85.405 197.435 ;
        RECT 85.575 197.105 85.905 197.605 ;
        RECT 86.075 196.935 86.330 197.435 ;
        RECT 85.580 196.765 86.330 196.935 ;
        RECT 87.055 196.935 87.225 197.435 ;
        RECT 87.395 197.105 87.725 197.605 ;
        RECT 87.055 196.765 87.720 196.935 ;
        RECT 85.580 195.775 85.810 196.765 ;
        RECT 85.980 195.945 86.330 196.595 ;
        RECT 86.970 195.945 87.320 196.595 ;
        RECT 87.490 195.775 87.720 196.765 ;
        RECT 85.580 195.605 86.330 195.775 ;
        RECT 85.575 195.055 85.905 195.435 ;
        RECT 86.075 195.315 86.330 195.605 ;
        RECT 87.055 195.605 87.720 195.775 ;
        RECT 87.055 195.315 87.225 195.605 ;
        RECT 87.395 195.055 87.725 195.435 ;
        RECT 87.895 195.315 88.120 197.435 ;
        RECT 88.335 197.105 88.665 197.605 ;
        RECT 88.835 196.935 89.005 197.435 ;
        RECT 89.240 197.220 90.070 197.390 ;
        RECT 90.310 197.225 90.690 197.605 ;
        RECT 88.310 196.765 89.005 196.935 ;
        RECT 88.310 195.795 88.480 196.765 ;
        RECT 88.650 195.975 89.060 196.595 ;
        RECT 89.230 196.545 89.730 196.925 ;
        RECT 88.310 195.605 89.005 195.795 ;
        RECT 89.230 195.675 89.450 196.545 ;
        RECT 89.900 196.375 90.070 197.220 ;
        RECT 90.870 197.055 91.040 197.345 ;
        RECT 91.210 197.225 91.540 197.605 ;
        RECT 92.010 197.135 92.640 197.385 ;
        RECT 92.820 197.225 93.240 197.605 ;
        RECT 92.470 197.055 92.640 197.135 ;
        RECT 93.440 197.055 93.680 197.345 ;
        RECT 90.240 196.805 91.610 197.055 ;
        RECT 90.240 196.545 90.490 196.805 ;
        RECT 91.000 196.375 91.250 196.535 ;
        RECT 89.900 196.205 91.250 196.375 ;
        RECT 89.900 196.165 90.320 196.205 ;
        RECT 89.630 195.615 89.980 195.985 ;
        RECT 88.335 195.055 88.665 195.435 ;
        RECT 88.835 195.275 89.005 195.605 ;
        RECT 90.150 195.435 90.320 196.165 ;
        RECT 91.420 196.035 91.610 196.805 ;
        RECT 90.490 195.705 90.900 196.035 ;
        RECT 91.190 195.695 91.610 196.035 ;
        RECT 91.780 196.625 92.300 196.935 ;
        RECT 92.470 196.885 93.680 197.055 ;
        RECT 93.910 196.915 94.240 197.605 ;
        RECT 91.780 195.865 91.950 196.625 ;
        RECT 92.120 196.035 92.300 196.445 ;
        RECT 92.470 196.375 92.640 196.885 ;
        RECT 94.410 196.735 94.580 197.345 ;
        RECT 94.850 196.885 95.180 197.395 ;
        RECT 94.410 196.715 94.730 196.735 ;
        RECT 92.810 196.545 94.730 196.715 ;
        RECT 92.470 196.205 94.370 196.375 ;
        RECT 92.700 195.865 93.030 195.985 ;
        RECT 91.780 195.695 93.030 195.865 ;
        RECT 89.305 195.235 90.320 195.435 ;
        RECT 90.490 195.055 90.900 195.495 ;
        RECT 91.190 195.265 91.440 195.695 ;
        RECT 91.640 195.055 91.960 195.515 ;
        RECT 93.200 195.445 93.370 196.205 ;
        RECT 94.040 196.145 94.370 196.205 ;
        RECT 93.560 195.975 93.890 196.035 ;
        RECT 93.560 195.705 94.220 195.975 ;
        RECT 94.540 195.650 94.730 196.545 ;
        RECT 92.520 195.275 93.370 195.445 ;
        RECT 93.570 195.055 94.230 195.535 ;
        RECT 94.410 195.320 94.730 195.650 ;
        RECT 94.930 196.295 95.180 196.885 ;
        RECT 95.360 196.805 95.645 197.605 ;
        RECT 95.825 196.625 96.080 197.295 ;
        RECT 94.930 195.965 95.730 196.295 ;
        RECT 94.930 195.315 95.180 195.965 ;
        RECT 95.900 195.765 96.080 196.625 ;
        RECT 96.625 196.515 100.135 197.605 ;
        RECT 96.625 195.995 98.315 196.515 ;
        RECT 100.345 196.465 100.575 197.605 ;
        RECT 100.745 196.455 101.075 197.435 ;
        RECT 101.245 196.465 101.455 197.605 ;
        RECT 98.485 195.825 100.135 196.345 ;
        RECT 100.325 196.045 100.655 196.295 ;
        RECT 95.825 195.565 96.080 195.765 ;
        RECT 95.360 195.055 95.645 195.515 ;
        RECT 95.825 195.395 96.165 195.565 ;
        RECT 95.825 195.235 96.080 195.395 ;
        RECT 96.625 195.055 100.135 195.825 ;
        RECT 100.345 195.055 100.575 195.875 ;
        RECT 100.825 195.855 101.075 196.455 ;
        RECT 101.685 196.440 101.975 197.605 ;
        RECT 103.155 196.675 103.325 197.435 ;
        RECT 103.505 196.845 103.835 197.605 ;
        RECT 103.155 196.505 103.820 196.675 ;
        RECT 104.005 196.530 104.275 197.435 ;
        RECT 103.650 196.360 103.820 196.505 ;
        RECT 103.085 195.955 103.415 196.325 ;
        RECT 103.650 196.030 103.935 196.360 ;
        RECT 100.745 195.225 101.075 195.855 ;
        RECT 101.245 195.055 101.455 195.875 ;
        RECT 101.685 195.055 101.975 195.780 ;
        RECT 103.650 195.775 103.820 196.030 ;
        RECT 103.155 195.605 103.820 195.775 ;
        RECT 104.105 195.730 104.275 196.530 ;
        RECT 104.445 196.515 107.955 197.605 ;
        RECT 104.445 195.995 106.135 196.515 ;
        RECT 108.165 196.465 108.395 197.605 ;
        RECT 108.565 196.455 108.895 197.435 ;
        RECT 109.065 196.465 109.275 197.605 ;
        RECT 106.305 195.825 107.955 196.345 ;
        RECT 108.145 196.045 108.475 196.295 ;
        RECT 103.155 195.225 103.325 195.605 ;
        RECT 103.505 195.055 103.835 195.435 ;
        RECT 104.015 195.225 104.275 195.730 ;
        RECT 104.445 195.055 107.955 195.825 ;
        RECT 108.165 195.055 108.395 195.875 ;
        RECT 108.645 195.855 108.895 196.455 ;
        RECT 109.510 196.415 109.765 197.295 ;
        RECT 109.935 196.465 110.240 197.605 ;
        RECT 110.580 197.225 110.910 197.605 ;
        RECT 111.090 197.055 111.260 197.345 ;
        RECT 111.430 197.145 111.680 197.605 ;
        RECT 110.460 196.885 111.260 197.055 ;
        RECT 111.850 197.095 112.720 197.435 ;
        RECT 108.565 195.225 108.895 195.855 ;
        RECT 109.065 195.055 109.275 195.875 ;
        RECT 109.510 195.765 109.720 196.415 ;
        RECT 110.460 196.295 110.630 196.885 ;
        RECT 111.850 196.715 112.020 197.095 ;
        RECT 112.955 196.975 113.125 197.435 ;
        RECT 113.295 197.145 113.665 197.605 ;
        RECT 113.960 197.005 114.130 197.345 ;
        RECT 114.300 197.175 114.630 197.605 ;
        RECT 114.865 197.005 115.035 197.345 ;
        RECT 110.800 196.545 112.020 196.715 ;
        RECT 112.190 196.635 112.650 196.925 ;
        RECT 112.955 196.805 113.515 196.975 ;
        RECT 113.960 196.835 115.035 197.005 ;
        RECT 115.205 197.105 115.885 197.435 ;
        RECT 116.100 197.105 116.350 197.435 ;
        RECT 116.520 197.145 116.770 197.605 ;
        RECT 113.345 196.665 113.515 196.805 ;
        RECT 112.190 196.625 113.155 196.635 ;
        RECT 111.850 196.455 112.020 196.545 ;
        RECT 112.480 196.465 113.155 196.625 ;
        RECT 109.890 196.265 110.630 196.295 ;
        RECT 109.890 195.965 110.805 196.265 ;
        RECT 110.480 195.790 110.805 195.965 ;
        RECT 109.510 195.235 109.765 195.765 ;
        RECT 109.935 195.055 110.240 195.515 ;
        RECT 110.485 195.435 110.805 195.790 ;
        RECT 110.975 196.005 111.515 196.375 ;
        RECT 111.850 196.285 112.255 196.455 ;
        RECT 110.975 195.605 111.215 196.005 ;
        RECT 111.695 195.835 111.915 196.115 ;
        RECT 111.385 195.665 111.915 195.835 ;
        RECT 111.385 195.435 111.555 195.665 ;
        RECT 112.085 195.505 112.255 196.285 ;
        RECT 112.425 195.675 112.775 196.295 ;
        RECT 112.945 195.675 113.155 196.465 ;
        RECT 113.345 196.495 114.845 196.665 ;
        RECT 113.345 195.805 113.515 196.495 ;
        RECT 115.205 196.325 115.375 197.105 ;
        RECT 116.180 196.975 116.350 197.105 ;
        RECT 113.685 196.155 115.375 196.325 ;
        RECT 115.545 196.545 116.010 196.935 ;
        RECT 116.180 196.805 116.575 196.975 ;
        RECT 113.685 195.975 113.855 196.155 ;
        RECT 110.485 195.265 111.555 195.435 ;
        RECT 111.725 195.055 111.915 195.495 ;
        RECT 112.085 195.225 113.035 195.505 ;
        RECT 113.345 195.415 113.605 195.805 ;
        RECT 114.025 195.735 114.815 195.985 ;
        RECT 113.255 195.245 113.605 195.415 ;
        RECT 113.815 195.055 114.145 195.515 ;
        RECT 115.020 195.445 115.190 196.155 ;
        RECT 115.545 195.955 115.715 196.545 ;
        RECT 115.360 195.735 115.715 195.955 ;
        RECT 115.885 195.735 116.235 196.355 ;
        RECT 116.405 195.445 116.575 196.805 ;
        RECT 116.940 196.635 117.265 197.420 ;
        RECT 116.745 195.585 117.205 196.635 ;
        RECT 115.020 195.275 115.875 195.445 ;
        RECT 116.080 195.275 116.575 195.445 ;
        RECT 116.745 195.055 117.075 195.415 ;
        RECT 117.435 195.315 117.605 197.435 ;
        RECT 117.775 197.105 118.105 197.605 ;
        RECT 118.275 196.935 118.530 197.435 ;
        RECT 117.780 196.765 118.530 196.935 ;
        RECT 117.780 195.775 118.010 196.765 ;
        RECT 118.180 195.945 118.530 196.595 ;
        RECT 118.705 196.530 118.975 197.435 ;
        RECT 119.145 196.845 119.475 197.605 ;
        RECT 119.655 196.675 119.825 197.435 ;
        RECT 121.010 197.170 126.355 197.605 ;
        RECT 117.780 195.605 118.530 195.775 ;
        RECT 117.775 195.055 118.105 195.435 ;
        RECT 118.275 195.315 118.530 195.605 ;
        RECT 118.705 195.730 118.875 196.530 ;
        RECT 119.160 196.505 119.825 196.675 ;
        RECT 119.160 196.360 119.330 196.505 ;
        RECT 119.045 196.030 119.330 196.360 ;
        RECT 119.160 195.775 119.330 196.030 ;
        RECT 119.565 195.955 119.895 196.325 ;
        RECT 122.600 195.920 122.950 197.170 ;
        RECT 126.525 196.515 127.735 197.605 ;
        RECT 118.705 195.225 118.965 195.730 ;
        RECT 119.160 195.605 119.825 195.775 ;
        RECT 119.145 195.055 119.475 195.435 ;
        RECT 119.655 195.225 119.825 195.605 ;
        RECT 124.430 195.600 124.770 196.430 ;
        RECT 126.525 195.975 127.045 196.515 ;
        RECT 127.215 195.805 127.735 196.345 ;
        RECT 121.010 195.055 126.355 195.600 ;
        RECT 126.525 195.055 127.735 195.805 ;
        RECT 20.640 194.885 127.820 195.055 ;
        RECT 20.725 194.135 21.935 194.885 ;
        RECT 22.570 194.340 27.915 194.885 ;
        RECT 20.725 193.595 21.245 194.135 ;
        RECT 21.415 193.425 21.935 193.965 ;
        RECT 20.725 192.335 21.935 193.425 ;
        RECT 24.160 192.770 24.510 194.020 ;
        RECT 25.990 193.510 26.330 194.340 ;
        RECT 28.090 194.335 28.345 194.625 ;
        RECT 28.515 194.505 28.845 194.885 ;
        RECT 28.090 194.165 28.840 194.335 ;
        RECT 28.090 193.345 28.440 193.995 ;
        RECT 28.610 193.175 28.840 194.165 ;
        RECT 28.090 193.005 28.840 193.175 ;
        RECT 22.570 192.335 27.915 192.770 ;
        RECT 28.090 192.505 28.345 193.005 ;
        RECT 28.515 192.335 28.845 192.835 ;
        RECT 29.015 192.505 29.185 194.625 ;
        RECT 29.545 194.525 29.875 194.885 ;
        RECT 30.045 194.495 30.540 194.665 ;
        RECT 30.745 194.495 31.600 194.665 ;
        RECT 29.415 193.305 29.875 194.355 ;
        RECT 29.355 192.520 29.680 193.305 ;
        RECT 30.045 193.135 30.215 194.495 ;
        RECT 30.385 193.585 30.735 194.205 ;
        RECT 30.905 193.985 31.260 194.205 ;
        RECT 30.905 193.395 31.075 193.985 ;
        RECT 31.430 193.785 31.600 194.495 ;
        RECT 32.475 194.425 32.805 194.885 ;
        RECT 33.015 194.525 33.365 194.695 ;
        RECT 31.805 193.955 32.595 194.205 ;
        RECT 33.015 194.135 33.275 194.525 ;
        RECT 33.585 194.435 34.535 194.715 ;
        RECT 34.705 194.445 34.895 194.885 ;
        RECT 35.065 194.505 36.135 194.675 ;
        RECT 32.765 193.785 32.935 193.965 ;
        RECT 30.045 192.965 30.440 193.135 ;
        RECT 30.610 193.005 31.075 193.395 ;
        RECT 31.245 193.615 32.935 193.785 ;
        RECT 30.270 192.835 30.440 192.965 ;
        RECT 31.245 192.835 31.415 193.615 ;
        RECT 33.105 193.445 33.275 194.135 ;
        RECT 31.775 193.275 33.275 193.445 ;
        RECT 33.465 193.475 33.675 194.265 ;
        RECT 33.845 193.645 34.195 194.265 ;
        RECT 34.365 193.655 34.535 194.435 ;
        RECT 35.065 194.275 35.235 194.505 ;
        RECT 34.705 194.105 35.235 194.275 ;
        RECT 34.705 193.825 34.925 194.105 ;
        RECT 35.405 193.935 35.645 194.335 ;
        RECT 34.365 193.485 34.770 193.655 ;
        RECT 35.105 193.565 35.645 193.935 ;
        RECT 35.815 194.150 36.135 194.505 ;
        RECT 36.380 194.425 36.685 194.885 ;
        RECT 36.855 194.175 37.110 194.705 ;
        RECT 35.815 193.975 36.140 194.150 ;
        RECT 35.815 193.675 36.730 193.975 ;
        RECT 35.990 193.645 36.730 193.675 ;
        RECT 33.465 193.315 34.140 193.475 ;
        RECT 34.600 193.395 34.770 193.485 ;
        RECT 33.465 193.305 34.430 193.315 ;
        RECT 33.105 193.135 33.275 193.275 ;
        RECT 29.850 192.335 30.100 192.795 ;
        RECT 30.270 192.505 30.520 192.835 ;
        RECT 30.735 192.505 31.415 192.835 ;
        RECT 31.585 192.935 32.660 193.105 ;
        RECT 33.105 192.965 33.665 193.135 ;
        RECT 33.970 193.015 34.430 193.305 ;
        RECT 34.600 193.225 35.820 193.395 ;
        RECT 31.585 192.595 31.755 192.935 ;
        RECT 31.990 192.335 32.320 192.765 ;
        RECT 32.490 192.595 32.660 192.935 ;
        RECT 32.955 192.335 33.325 192.795 ;
        RECT 33.495 192.505 33.665 192.965 ;
        RECT 34.600 192.845 34.770 193.225 ;
        RECT 35.990 193.055 36.160 193.645 ;
        RECT 36.900 193.525 37.110 194.175 ;
        RECT 37.285 194.160 37.575 194.885 ;
        RECT 37.745 194.135 38.955 194.885 ;
        RECT 33.900 192.505 34.770 192.845 ;
        RECT 35.360 192.885 36.160 193.055 ;
        RECT 34.940 192.335 35.190 192.795 ;
        RECT 35.360 192.595 35.530 192.885 ;
        RECT 35.710 192.335 36.040 192.715 ;
        RECT 36.380 192.335 36.685 193.475 ;
        RECT 36.855 192.645 37.110 193.525 ;
        RECT 37.285 192.335 37.575 193.500 ;
        RECT 37.745 193.425 38.265 193.965 ;
        RECT 38.435 193.595 38.955 194.135 ;
        RECT 39.500 194.175 39.755 194.705 ;
        RECT 39.935 194.425 40.220 194.885 ;
        RECT 37.745 192.335 38.955 193.425 ;
        RECT 39.500 193.315 39.680 194.175 ;
        RECT 40.400 193.975 40.650 194.625 ;
        RECT 39.850 193.645 40.650 193.975 ;
        RECT 39.500 192.845 39.755 193.315 ;
        RECT 39.415 192.675 39.755 192.845 ;
        RECT 39.500 192.645 39.755 192.675 ;
        RECT 39.935 192.335 40.220 193.135 ;
        RECT 40.400 193.055 40.650 193.645 ;
        RECT 40.850 194.290 41.170 194.620 ;
        RECT 41.350 194.405 42.010 194.885 ;
        RECT 42.210 194.495 43.060 194.665 ;
        RECT 40.850 193.395 41.040 194.290 ;
        RECT 41.360 193.965 42.020 194.235 ;
        RECT 41.690 193.905 42.020 193.965 ;
        RECT 41.210 193.735 41.540 193.795 ;
        RECT 42.210 193.735 42.380 194.495 ;
        RECT 43.620 194.425 43.940 194.885 ;
        RECT 44.140 194.245 44.390 194.675 ;
        RECT 44.680 194.445 45.090 194.885 ;
        RECT 45.260 194.505 46.275 194.705 ;
        RECT 42.550 194.075 43.800 194.245 ;
        RECT 42.550 193.955 42.880 194.075 ;
        RECT 41.210 193.565 43.110 193.735 ;
        RECT 40.850 193.225 42.770 193.395 ;
        RECT 40.850 193.205 41.170 193.225 ;
        RECT 40.400 192.545 40.730 193.055 ;
        RECT 41.000 192.595 41.170 193.205 ;
        RECT 42.940 193.055 43.110 193.565 ;
        RECT 43.280 193.495 43.460 193.905 ;
        RECT 43.630 193.315 43.800 194.075 ;
        RECT 41.340 192.335 41.670 193.025 ;
        RECT 41.900 192.885 43.110 193.055 ;
        RECT 43.280 193.005 43.800 193.315 ;
        RECT 43.970 193.905 44.390 194.245 ;
        RECT 44.680 193.905 45.090 194.235 ;
        RECT 43.970 193.135 44.160 193.905 ;
        RECT 45.260 193.775 45.430 194.505 ;
        RECT 46.575 194.335 46.745 194.665 ;
        RECT 46.915 194.505 47.245 194.885 ;
        RECT 45.600 193.955 45.950 194.325 ;
        RECT 45.260 193.735 45.680 193.775 ;
        RECT 44.330 193.565 45.680 193.735 ;
        RECT 44.330 193.405 44.580 193.565 ;
        RECT 45.090 193.135 45.340 193.395 ;
        RECT 43.970 192.885 45.340 193.135 ;
        RECT 41.900 192.595 42.140 192.885 ;
        RECT 42.940 192.805 43.110 192.885 ;
        RECT 42.340 192.335 42.760 192.715 ;
        RECT 42.940 192.555 43.570 192.805 ;
        RECT 44.040 192.335 44.370 192.715 ;
        RECT 44.540 192.595 44.710 192.885 ;
        RECT 45.510 192.720 45.680 193.565 ;
        RECT 46.130 193.395 46.350 194.265 ;
        RECT 46.575 194.145 47.270 194.335 ;
        RECT 45.850 193.015 46.350 193.395 ;
        RECT 46.520 193.345 46.930 193.965 ;
        RECT 47.100 193.175 47.270 194.145 ;
        RECT 46.575 193.005 47.270 193.175 ;
        RECT 44.890 192.335 45.270 192.715 ;
        RECT 45.510 192.550 46.340 192.720 ;
        RECT 46.575 192.505 46.745 193.005 ;
        RECT 46.915 192.335 47.245 192.835 ;
        RECT 47.460 192.505 47.685 194.625 ;
        RECT 47.855 194.505 48.185 194.885 ;
        RECT 48.355 194.335 48.525 194.625 ;
        RECT 47.860 194.165 48.525 194.335 ;
        RECT 48.785 194.210 49.045 194.715 ;
        RECT 49.225 194.505 49.555 194.885 ;
        RECT 49.735 194.335 49.905 194.715 ;
        RECT 47.860 193.175 48.090 194.165 ;
        RECT 48.260 193.345 48.610 193.995 ;
        RECT 48.785 193.410 48.955 194.210 ;
        RECT 49.240 194.165 49.905 194.335 ;
        RECT 50.165 194.210 50.425 194.715 ;
        RECT 50.605 194.505 50.935 194.885 ;
        RECT 51.115 194.335 51.285 194.715 ;
        RECT 49.240 193.910 49.410 194.165 ;
        RECT 49.125 193.580 49.410 193.910 ;
        RECT 49.645 193.615 49.975 193.985 ;
        RECT 49.240 193.435 49.410 193.580 ;
        RECT 47.860 193.005 48.525 193.175 ;
        RECT 47.855 192.335 48.185 192.835 ;
        RECT 48.355 192.505 48.525 193.005 ;
        RECT 48.785 192.505 49.055 193.410 ;
        RECT 49.240 193.265 49.905 193.435 ;
        RECT 49.225 192.335 49.555 193.095 ;
        RECT 49.735 192.505 49.905 193.265 ;
        RECT 50.165 193.410 50.335 194.210 ;
        RECT 50.620 194.165 51.285 194.335 ;
        RECT 50.620 193.910 50.790 194.165 ;
        RECT 51.605 194.065 51.815 194.885 ;
        RECT 51.985 194.085 52.315 194.715 ;
        RECT 50.505 193.580 50.790 193.910 ;
        RECT 51.025 193.615 51.355 193.985 ;
        RECT 50.620 193.435 50.790 193.580 ;
        RECT 51.985 193.485 52.235 194.085 ;
        RECT 52.485 194.065 52.715 194.885 ;
        RECT 53.850 194.175 54.105 194.705 ;
        RECT 54.275 194.425 54.580 194.885 ;
        RECT 54.825 194.505 55.895 194.675 ;
        RECT 52.405 193.645 52.735 193.895 ;
        RECT 53.850 193.525 54.060 194.175 ;
        RECT 54.825 194.150 55.145 194.505 ;
        RECT 54.820 193.975 55.145 194.150 ;
        RECT 54.230 193.675 55.145 193.975 ;
        RECT 55.315 193.935 55.555 194.335 ;
        RECT 55.725 194.275 55.895 194.505 ;
        RECT 56.065 194.445 56.255 194.885 ;
        RECT 56.425 194.435 57.375 194.715 ;
        RECT 57.595 194.525 57.945 194.695 ;
        RECT 55.725 194.105 56.255 194.275 ;
        RECT 54.230 193.645 54.970 193.675 ;
        RECT 50.165 192.505 50.435 193.410 ;
        RECT 50.620 193.265 51.285 193.435 ;
        RECT 50.605 192.335 50.935 193.095 ;
        RECT 51.115 192.505 51.285 193.265 ;
        RECT 51.605 192.335 51.815 193.475 ;
        RECT 51.985 192.505 52.315 193.485 ;
        RECT 52.485 192.335 52.715 193.475 ;
        RECT 53.850 192.645 54.105 193.525 ;
        RECT 54.275 192.335 54.580 193.475 ;
        RECT 54.800 193.055 54.970 193.645 ;
        RECT 55.315 193.565 55.855 193.935 ;
        RECT 56.035 193.825 56.255 194.105 ;
        RECT 56.425 193.655 56.595 194.435 ;
        RECT 56.190 193.485 56.595 193.655 ;
        RECT 56.765 193.645 57.115 194.265 ;
        RECT 56.190 193.395 56.360 193.485 ;
        RECT 57.285 193.475 57.495 194.265 ;
        RECT 55.140 193.225 56.360 193.395 ;
        RECT 56.820 193.315 57.495 193.475 ;
        RECT 54.800 192.885 55.600 193.055 ;
        RECT 54.920 192.335 55.250 192.715 ;
        RECT 55.430 192.595 55.600 192.885 ;
        RECT 56.190 192.845 56.360 193.225 ;
        RECT 56.530 193.305 57.495 193.315 ;
        RECT 57.685 194.135 57.945 194.525 ;
        RECT 58.155 194.425 58.485 194.885 ;
        RECT 59.360 194.495 60.215 194.665 ;
        RECT 60.420 194.495 60.915 194.665 ;
        RECT 61.085 194.525 61.415 194.885 ;
        RECT 57.685 193.445 57.855 194.135 ;
        RECT 58.025 193.785 58.195 193.965 ;
        RECT 58.365 193.955 59.155 194.205 ;
        RECT 59.360 193.785 59.530 194.495 ;
        RECT 59.700 193.985 60.055 194.205 ;
        RECT 58.025 193.615 59.715 193.785 ;
        RECT 56.530 193.015 56.990 193.305 ;
        RECT 57.685 193.275 59.185 193.445 ;
        RECT 57.685 193.135 57.855 193.275 ;
        RECT 57.295 192.965 57.855 193.135 ;
        RECT 55.770 192.335 56.020 192.795 ;
        RECT 56.190 192.505 57.060 192.845 ;
        RECT 57.295 192.505 57.465 192.965 ;
        RECT 58.300 192.935 59.375 193.105 ;
        RECT 57.635 192.335 58.005 192.795 ;
        RECT 58.300 192.595 58.470 192.935 ;
        RECT 58.640 192.335 58.970 192.765 ;
        RECT 59.205 192.595 59.375 192.935 ;
        RECT 59.545 192.835 59.715 193.615 ;
        RECT 59.885 193.395 60.055 193.985 ;
        RECT 60.225 193.585 60.575 194.205 ;
        RECT 59.885 193.005 60.350 193.395 ;
        RECT 60.745 193.135 60.915 194.495 ;
        RECT 61.085 193.305 61.545 194.355 ;
        RECT 60.520 192.965 60.915 193.135 ;
        RECT 60.520 192.835 60.690 192.965 ;
        RECT 59.545 192.505 60.225 192.835 ;
        RECT 60.440 192.505 60.690 192.835 ;
        RECT 60.860 192.335 61.110 192.795 ;
        RECT 61.280 192.520 61.605 193.305 ;
        RECT 61.775 192.505 61.945 194.625 ;
        RECT 62.115 194.505 62.445 194.885 ;
        RECT 62.615 194.335 62.870 194.625 ;
        RECT 62.120 194.165 62.870 194.335 ;
        RECT 62.120 193.175 62.350 194.165 ;
        RECT 63.045 194.160 63.335 194.885 ;
        RECT 63.815 194.415 63.985 194.885 ;
        RECT 64.155 194.235 64.485 194.715 ;
        RECT 64.655 194.415 64.825 194.885 ;
        RECT 64.995 194.235 65.325 194.715 ;
        RECT 63.560 194.065 65.325 194.235 ;
        RECT 65.495 194.075 65.665 194.885 ;
        RECT 65.865 194.505 66.935 194.675 ;
        RECT 65.865 194.150 66.185 194.505 ;
        RECT 62.520 193.345 62.870 193.995 ;
        RECT 63.560 193.515 63.970 194.065 ;
        RECT 65.860 193.895 66.185 194.150 ;
        RECT 64.155 193.685 66.185 193.895 ;
        RECT 65.840 193.675 66.185 193.685 ;
        RECT 66.355 193.935 66.595 194.335 ;
        RECT 66.765 194.275 66.935 194.505 ;
        RECT 67.105 194.445 67.295 194.885 ;
        RECT 67.465 194.435 68.415 194.715 ;
        RECT 68.635 194.525 68.985 194.695 ;
        RECT 66.765 194.105 67.295 194.275 ;
        RECT 62.120 193.005 62.870 193.175 ;
        RECT 62.115 192.335 62.445 192.835 ;
        RECT 62.615 192.505 62.870 193.005 ;
        RECT 63.045 192.335 63.335 193.500 ;
        RECT 63.560 193.345 65.285 193.515 ;
        RECT 63.815 192.335 63.985 193.175 ;
        RECT 64.195 192.505 64.445 193.345 ;
        RECT 64.655 192.335 64.825 193.175 ;
        RECT 64.995 192.505 65.285 193.345 ;
        RECT 65.495 192.335 65.665 193.395 ;
        RECT 65.840 193.055 66.010 193.675 ;
        RECT 66.355 193.565 66.895 193.935 ;
        RECT 67.075 193.825 67.295 194.105 ;
        RECT 67.465 193.655 67.635 194.435 ;
        RECT 67.230 193.485 67.635 193.655 ;
        RECT 67.805 193.645 68.155 194.265 ;
        RECT 67.230 193.395 67.400 193.485 ;
        RECT 68.325 193.475 68.535 194.265 ;
        RECT 66.180 193.225 67.400 193.395 ;
        RECT 67.860 193.315 68.535 193.475 ;
        RECT 65.840 192.885 66.640 193.055 ;
        RECT 65.960 192.335 66.290 192.715 ;
        RECT 66.470 192.595 66.640 192.885 ;
        RECT 67.230 192.845 67.400 193.225 ;
        RECT 67.570 193.305 68.535 193.315 ;
        RECT 68.725 194.135 68.985 194.525 ;
        RECT 69.195 194.425 69.525 194.885 ;
        RECT 70.400 194.495 71.255 194.665 ;
        RECT 71.460 194.495 71.955 194.665 ;
        RECT 72.125 194.525 72.455 194.885 ;
        RECT 68.725 193.445 68.895 194.135 ;
        RECT 69.065 193.785 69.235 193.965 ;
        RECT 69.405 193.955 70.195 194.205 ;
        RECT 70.400 193.785 70.570 194.495 ;
        RECT 70.740 193.985 71.095 194.205 ;
        RECT 69.065 193.615 70.755 193.785 ;
        RECT 67.570 193.015 68.030 193.305 ;
        RECT 68.725 193.275 70.225 193.445 ;
        RECT 68.725 193.135 68.895 193.275 ;
        RECT 68.335 192.965 68.895 193.135 ;
        RECT 66.810 192.335 67.060 192.795 ;
        RECT 67.230 192.505 68.100 192.845 ;
        RECT 68.335 192.505 68.505 192.965 ;
        RECT 69.340 192.935 70.415 193.105 ;
        RECT 68.675 192.335 69.045 192.795 ;
        RECT 69.340 192.595 69.510 192.935 ;
        RECT 69.680 192.335 70.010 192.765 ;
        RECT 70.245 192.595 70.415 192.935 ;
        RECT 70.585 192.835 70.755 193.615 ;
        RECT 70.925 193.395 71.095 193.985 ;
        RECT 71.265 193.585 71.615 194.205 ;
        RECT 70.925 193.005 71.390 193.395 ;
        RECT 71.785 193.135 71.955 194.495 ;
        RECT 72.125 193.305 72.585 194.355 ;
        RECT 71.560 192.965 71.955 193.135 ;
        RECT 71.560 192.835 71.730 192.965 ;
        RECT 70.585 192.505 71.265 192.835 ;
        RECT 71.480 192.505 71.730 192.835 ;
        RECT 71.900 192.335 72.150 192.795 ;
        RECT 72.320 192.520 72.645 193.305 ;
        RECT 72.815 192.505 72.985 194.625 ;
        RECT 73.155 194.505 73.485 194.885 ;
        RECT 73.655 194.335 73.910 194.625 ;
        RECT 73.160 194.165 73.910 194.335 ;
        RECT 74.085 194.210 74.360 194.555 ;
        RECT 74.550 194.485 74.925 194.885 ;
        RECT 75.095 194.315 75.265 194.665 ;
        RECT 75.435 194.485 75.765 194.885 ;
        RECT 75.935 194.315 76.195 194.715 ;
        RECT 73.160 193.175 73.390 194.165 ;
        RECT 73.560 193.345 73.910 193.995 ;
        RECT 74.085 193.475 74.255 194.210 ;
        RECT 74.530 194.145 76.195 194.315 ;
        RECT 74.530 193.975 74.700 194.145 ;
        RECT 76.375 194.065 76.705 194.485 ;
        RECT 76.875 194.065 77.135 194.885 ;
        RECT 77.340 194.145 77.955 194.715 ;
        RECT 78.125 194.375 78.340 194.885 ;
        RECT 78.570 194.375 78.850 194.705 ;
        RECT 79.030 194.375 79.270 194.885 ;
        RECT 76.375 193.975 76.625 194.065 ;
        RECT 74.425 193.645 74.700 193.975 ;
        RECT 74.870 193.645 75.695 193.975 ;
        RECT 75.910 193.645 76.625 193.975 ;
        RECT 76.795 193.645 77.130 193.895 ;
        RECT 74.530 193.475 74.700 193.645 ;
        RECT 73.160 193.005 73.910 193.175 ;
        RECT 73.155 192.335 73.485 192.835 ;
        RECT 73.655 192.505 73.910 193.005 ;
        RECT 74.085 192.505 74.360 193.475 ;
        RECT 74.530 193.305 75.190 193.475 ;
        RECT 75.450 193.355 75.695 193.645 ;
        RECT 75.020 193.185 75.190 193.305 ;
        RECT 75.865 193.185 76.195 193.475 ;
        RECT 74.570 192.335 74.850 193.135 ;
        RECT 75.020 193.015 76.195 193.185 ;
        RECT 76.455 193.085 76.625 193.645 ;
        RECT 75.020 192.515 76.635 192.845 ;
        RECT 76.875 192.335 77.135 193.475 ;
        RECT 77.340 193.125 77.655 194.145 ;
        RECT 77.825 193.475 77.995 193.975 ;
        RECT 78.245 193.645 78.510 194.205 ;
        RECT 78.680 193.475 78.850 194.375 ;
        RECT 79.695 194.335 79.865 194.715 ;
        RECT 80.080 194.505 80.410 194.885 ;
        RECT 79.020 193.645 79.375 194.205 ;
        RECT 79.695 194.165 80.410 194.335 ;
        RECT 79.605 193.615 79.960 193.985 ;
        RECT 80.240 193.975 80.410 194.165 ;
        RECT 80.580 194.140 80.835 194.715 ;
        RECT 80.240 193.645 80.495 193.975 ;
        RECT 77.825 193.305 79.250 193.475 ;
        RECT 80.240 193.435 80.410 193.645 ;
        RECT 77.340 192.505 77.875 193.125 ;
        RECT 78.045 192.335 78.375 193.135 ;
        RECT 78.860 193.130 79.250 193.305 ;
        RECT 79.695 193.265 80.410 193.435 ;
        RECT 80.665 193.410 80.835 194.140 ;
        RECT 81.010 194.045 81.270 194.885 ;
        RECT 81.445 194.085 82.140 194.715 ;
        RECT 82.345 194.085 82.655 194.885 ;
        RECT 82.825 194.115 84.495 194.885 ;
        RECT 84.755 194.335 84.925 194.715 ;
        RECT 85.105 194.505 85.435 194.885 ;
        RECT 84.755 194.165 85.420 194.335 ;
        RECT 85.615 194.210 85.875 194.715 ;
        RECT 81.465 193.645 81.800 193.895 ;
        RECT 81.970 193.485 82.140 194.085 ;
        RECT 82.310 193.645 82.645 193.915 ;
        RECT 79.695 192.505 79.865 193.265 ;
        RECT 80.080 192.335 80.410 193.095 ;
        RECT 80.580 192.505 80.835 193.410 ;
        RECT 81.010 192.335 81.270 193.485 ;
        RECT 81.445 192.335 81.705 193.475 ;
        RECT 81.875 192.505 82.205 193.485 ;
        RECT 82.375 192.335 82.655 193.475 ;
        RECT 82.825 193.425 83.575 193.945 ;
        RECT 83.745 193.595 84.495 194.115 ;
        RECT 84.685 193.615 85.015 193.985 ;
        RECT 85.250 193.910 85.420 194.165 ;
        RECT 85.250 193.580 85.535 193.910 ;
        RECT 85.250 193.435 85.420 193.580 ;
        RECT 82.825 192.335 84.495 193.425 ;
        RECT 84.755 193.265 85.420 193.435 ;
        RECT 85.705 193.410 85.875 194.210 ;
        RECT 86.105 194.065 86.315 194.885 ;
        RECT 86.485 194.085 86.815 194.715 ;
        RECT 86.485 193.485 86.735 194.085 ;
        RECT 86.985 194.065 87.215 194.885 ;
        RECT 87.465 194.065 87.695 194.885 ;
        RECT 87.865 194.085 88.195 194.715 ;
        RECT 86.905 193.645 87.235 193.895 ;
        RECT 87.445 193.645 87.775 193.895 ;
        RECT 87.945 193.485 88.195 194.085 ;
        RECT 88.365 194.065 88.575 194.885 ;
        RECT 88.805 194.160 89.095 194.885 ;
        RECT 89.640 194.175 89.895 194.705 ;
        RECT 90.075 194.425 90.360 194.885 ;
        RECT 84.755 192.505 84.925 193.265 ;
        RECT 85.105 192.335 85.435 193.095 ;
        RECT 85.605 192.505 85.875 193.410 ;
        RECT 86.105 192.335 86.315 193.475 ;
        RECT 86.485 192.505 86.815 193.485 ;
        RECT 86.985 192.335 87.215 193.475 ;
        RECT 87.465 192.335 87.695 193.475 ;
        RECT 87.865 192.505 88.195 193.485 ;
        RECT 88.365 192.335 88.575 193.475 ;
        RECT 88.805 192.335 89.095 193.500 ;
        RECT 89.640 193.315 89.820 194.175 ;
        RECT 90.540 193.975 90.790 194.625 ;
        RECT 89.990 193.645 90.790 193.975 ;
        RECT 89.640 192.845 89.895 193.315 ;
        RECT 89.555 192.675 89.895 192.845 ;
        RECT 89.640 192.645 89.895 192.675 ;
        RECT 90.075 192.335 90.360 193.135 ;
        RECT 90.540 193.055 90.790 193.645 ;
        RECT 90.990 194.290 91.310 194.620 ;
        RECT 91.490 194.405 92.150 194.885 ;
        RECT 92.350 194.495 93.200 194.665 ;
        RECT 90.990 193.395 91.180 194.290 ;
        RECT 91.500 193.965 92.160 194.235 ;
        RECT 91.830 193.905 92.160 193.965 ;
        RECT 91.350 193.735 91.680 193.795 ;
        RECT 92.350 193.735 92.520 194.495 ;
        RECT 93.760 194.425 94.080 194.885 ;
        RECT 94.280 194.245 94.530 194.675 ;
        RECT 94.820 194.445 95.230 194.885 ;
        RECT 95.400 194.505 96.415 194.705 ;
        RECT 92.690 194.075 93.940 194.245 ;
        RECT 92.690 193.955 93.020 194.075 ;
        RECT 91.350 193.565 93.250 193.735 ;
        RECT 90.990 193.225 92.910 193.395 ;
        RECT 90.990 193.205 91.310 193.225 ;
        RECT 90.540 192.545 90.870 193.055 ;
        RECT 91.140 192.595 91.310 193.205 ;
        RECT 93.080 193.055 93.250 193.565 ;
        RECT 93.420 193.495 93.600 193.905 ;
        RECT 93.770 193.315 93.940 194.075 ;
        RECT 91.480 192.335 91.810 193.025 ;
        RECT 92.040 192.885 93.250 193.055 ;
        RECT 93.420 193.005 93.940 193.315 ;
        RECT 94.110 193.905 94.530 194.245 ;
        RECT 94.820 193.905 95.230 194.235 ;
        RECT 94.110 193.135 94.300 193.905 ;
        RECT 95.400 193.775 95.570 194.505 ;
        RECT 96.715 194.335 96.885 194.665 ;
        RECT 97.055 194.505 97.385 194.885 ;
        RECT 95.740 193.955 96.090 194.325 ;
        RECT 95.400 193.735 95.820 193.775 ;
        RECT 94.470 193.565 95.820 193.735 ;
        RECT 94.470 193.405 94.720 193.565 ;
        RECT 95.230 193.135 95.480 193.395 ;
        RECT 94.110 192.885 95.480 193.135 ;
        RECT 92.040 192.595 92.280 192.885 ;
        RECT 93.080 192.805 93.250 192.885 ;
        RECT 92.480 192.335 92.900 192.715 ;
        RECT 93.080 192.555 93.710 192.805 ;
        RECT 94.180 192.335 94.510 192.715 ;
        RECT 94.680 192.595 94.850 192.885 ;
        RECT 95.650 192.720 95.820 193.565 ;
        RECT 96.270 193.395 96.490 194.265 ;
        RECT 96.715 194.145 97.410 194.335 ;
        RECT 95.990 193.015 96.490 193.395 ;
        RECT 96.660 193.345 97.070 193.965 ;
        RECT 97.240 193.175 97.410 194.145 ;
        RECT 96.715 193.005 97.410 193.175 ;
        RECT 95.030 192.335 95.410 192.715 ;
        RECT 95.650 192.550 96.480 192.720 ;
        RECT 96.715 192.505 96.885 193.005 ;
        RECT 97.055 192.335 97.385 192.835 ;
        RECT 97.600 192.505 97.825 194.625 ;
        RECT 97.995 194.505 98.325 194.885 ;
        RECT 98.495 194.335 98.665 194.625 ;
        RECT 98.000 194.165 98.665 194.335 ;
        RECT 98.000 193.175 98.230 194.165 ;
        RECT 99.200 194.075 99.445 194.680 ;
        RECT 99.665 194.350 100.175 194.885 ;
        RECT 98.400 193.345 98.750 193.995 ;
        RECT 98.925 193.905 100.155 194.075 ;
        RECT 98.000 193.005 98.665 193.175 ;
        RECT 97.995 192.335 98.325 192.835 ;
        RECT 98.495 192.505 98.665 193.005 ;
        RECT 98.925 193.095 99.265 193.905 ;
        RECT 99.435 193.340 100.185 193.530 ;
        RECT 98.925 192.685 99.440 193.095 ;
        RECT 99.675 192.335 99.845 193.095 ;
        RECT 100.015 192.675 100.185 193.340 ;
        RECT 100.355 193.355 100.545 194.715 ;
        RECT 100.715 193.865 100.990 194.715 ;
        RECT 101.180 194.350 101.710 194.715 ;
        RECT 102.135 194.485 102.465 194.885 ;
        RECT 101.535 194.315 101.710 194.350 ;
        RECT 100.715 193.695 100.995 193.865 ;
        RECT 100.715 193.555 100.990 193.695 ;
        RECT 101.195 193.355 101.365 194.155 ;
        RECT 100.355 193.185 101.365 193.355 ;
        RECT 101.535 194.145 102.465 194.315 ;
        RECT 102.635 194.145 102.890 194.715 ;
        RECT 101.535 193.015 101.705 194.145 ;
        RECT 102.295 193.975 102.465 194.145 ;
        RECT 100.580 192.845 101.705 193.015 ;
        RECT 101.875 193.645 102.070 193.975 ;
        RECT 102.295 193.645 102.550 193.975 ;
        RECT 101.875 192.675 102.045 193.645 ;
        RECT 102.720 193.475 102.890 194.145 ;
        RECT 103.065 194.115 104.735 194.885 ;
        RECT 104.910 194.340 110.255 194.885 ;
        RECT 100.015 192.505 102.045 192.675 ;
        RECT 102.215 192.335 102.385 193.475 ;
        RECT 102.555 192.505 102.890 193.475 ;
        RECT 103.065 193.425 103.815 193.945 ;
        RECT 103.985 193.595 104.735 194.115 ;
        RECT 103.065 192.335 104.735 193.425 ;
        RECT 106.500 192.770 106.850 194.020 ;
        RECT 108.330 193.510 108.670 194.340 ;
        RECT 110.700 194.075 110.945 194.680 ;
        RECT 111.165 194.350 111.675 194.885 ;
        RECT 110.425 193.905 111.655 194.075 ;
        RECT 110.425 193.095 110.765 193.905 ;
        RECT 110.935 193.340 111.685 193.530 ;
        RECT 104.910 192.335 110.255 192.770 ;
        RECT 110.425 192.685 110.940 193.095 ;
        RECT 111.175 192.335 111.345 193.095 ;
        RECT 111.515 192.675 111.685 193.340 ;
        RECT 111.855 193.355 112.045 194.715 ;
        RECT 112.215 193.865 112.490 194.715 ;
        RECT 112.680 194.350 113.210 194.715 ;
        RECT 113.635 194.485 113.965 194.885 ;
        RECT 113.035 194.315 113.210 194.350 ;
        RECT 112.215 193.695 112.495 193.865 ;
        RECT 112.215 193.555 112.490 193.695 ;
        RECT 112.695 193.355 112.865 194.155 ;
        RECT 111.855 193.185 112.865 193.355 ;
        RECT 113.035 194.145 113.965 194.315 ;
        RECT 114.135 194.145 114.390 194.715 ;
        RECT 114.565 194.160 114.855 194.885 ;
        RECT 113.035 193.015 113.205 194.145 ;
        RECT 113.795 193.975 113.965 194.145 ;
        RECT 112.080 192.845 113.205 193.015 ;
        RECT 113.375 193.645 113.570 193.975 ;
        RECT 113.795 193.645 114.050 193.975 ;
        RECT 113.375 192.675 113.545 193.645 ;
        RECT 114.220 193.475 114.390 194.145 ;
        RECT 115.985 194.065 116.215 194.885 ;
        RECT 116.385 194.085 116.715 194.715 ;
        RECT 115.965 193.645 116.295 193.895 ;
        RECT 111.515 192.505 113.545 192.675 ;
        RECT 113.715 192.335 113.885 193.475 ;
        RECT 114.055 192.505 114.390 193.475 ;
        RECT 114.565 192.335 114.855 193.500 ;
        RECT 116.465 193.485 116.715 194.085 ;
        RECT 116.885 194.065 117.095 194.885 ;
        RECT 117.325 194.115 118.995 194.885 ;
        RECT 119.255 194.335 119.425 194.715 ;
        RECT 119.605 194.505 119.935 194.885 ;
        RECT 119.255 194.165 119.920 194.335 ;
        RECT 120.115 194.210 120.375 194.715 ;
        RECT 121.010 194.340 126.355 194.885 ;
        RECT 115.985 192.335 116.215 193.475 ;
        RECT 116.385 192.505 116.715 193.485 ;
        RECT 116.885 192.335 117.095 193.475 ;
        RECT 117.325 193.425 118.075 193.945 ;
        RECT 118.245 193.595 118.995 194.115 ;
        RECT 119.185 193.615 119.515 193.985 ;
        RECT 119.750 193.910 119.920 194.165 ;
        RECT 119.750 193.580 120.035 193.910 ;
        RECT 119.750 193.435 119.920 193.580 ;
        RECT 117.325 192.335 118.995 193.425 ;
        RECT 119.255 193.265 119.920 193.435 ;
        RECT 120.205 193.410 120.375 194.210 ;
        RECT 119.255 192.505 119.425 193.265 ;
        RECT 119.605 192.335 119.935 193.095 ;
        RECT 120.105 192.505 120.375 193.410 ;
        RECT 122.600 192.770 122.950 194.020 ;
        RECT 124.430 193.510 124.770 194.340 ;
        RECT 126.525 194.135 127.735 194.885 ;
        RECT 126.525 193.425 127.045 193.965 ;
        RECT 127.215 193.595 127.735 194.135 ;
        RECT 121.010 192.335 126.355 192.770 ;
        RECT 126.525 192.335 127.735 193.425 ;
        RECT 20.640 192.165 127.820 192.335 ;
        RECT 20.725 191.075 21.935 192.165 ;
        RECT 20.725 190.365 21.245 190.905 ;
        RECT 21.415 190.535 21.935 191.075 ;
        RECT 22.565 191.075 24.235 192.165 ;
        RECT 22.565 190.555 23.315 191.075 ;
        RECT 24.405 191.000 24.695 192.165 ;
        RECT 24.865 191.075 26.075 192.165 ;
        RECT 26.250 191.730 31.595 192.165 ;
        RECT 23.485 190.385 24.235 190.905 ;
        RECT 24.865 190.535 25.385 191.075 ;
        RECT 20.725 189.615 21.935 190.365 ;
        RECT 22.565 189.615 24.235 190.385 ;
        RECT 25.555 190.365 26.075 190.905 ;
        RECT 27.840 190.480 28.190 191.730 ;
        RECT 31.805 191.025 32.035 192.165 ;
        RECT 32.205 191.015 32.535 191.995 ;
        RECT 32.705 191.025 32.915 192.165 ;
        RECT 34.065 191.090 34.335 191.995 ;
        RECT 34.505 191.405 34.835 192.165 ;
        RECT 35.015 191.235 35.185 191.995 ;
        RECT 24.405 189.615 24.695 190.340 ;
        RECT 24.865 189.615 26.075 190.365 ;
        RECT 29.670 190.160 30.010 190.990 ;
        RECT 31.785 190.605 32.115 190.855 ;
        RECT 26.250 189.615 31.595 190.160 ;
        RECT 31.805 189.615 32.035 190.435 ;
        RECT 32.285 190.415 32.535 191.015 ;
        RECT 32.205 189.785 32.535 190.415 ;
        RECT 32.705 189.615 32.915 190.435 ;
        RECT 34.065 190.290 34.235 191.090 ;
        RECT 34.520 191.065 35.185 191.235 ;
        RECT 34.520 190.920 34.690 191.065 ;
        RECT 34.405 190.590 34.690 190.920 ;
        RECT 35.450 191.025 35.785 191.995 ;
        RECT 35.955 191.025 36.125 192.165 ;
        RECT 36.295 191.825 38.325 191.995 ;
        RECT 34.520 190.335 34.690 190.590 ;
        RECT 34.925 190.515 35.255 190.885 ;
        RECT 35.450 190.355 35.620 191.025 ;
        RECT 36.295 190.855 36.465 191.825 ;
        RECT 35.790 190.525 36.045 190.855 ;
        RECT 36.270 190.525 36.465 190.855 ;
        RECT 36.635 191.485 37.760 191.655 ;
        RECT 35.875 190.355 36.045 190.525 ;
        RECT 36.635 190.355 36.805 191.485 ;
        RECT 34.065 189.785 34.325 190.290 ;
        RECT 34.520 190.165 35.185 190.335 ;
        RECT 34.505 189.615 34.835 189.995 ;
        RECT 35.015 189.785 35.185 190.165 ;
        RECT 35.450 189.785 35.705 190.355 ;
        RECT 35.875 190.185 36.805 190.355 ;
        RECT 36.975 191.145 37.985 191.315 ;
        RECT 36.975 190.345 37.145 191.145 ;
        RECT 36.630 190.150 36.805 190.185 ;
        RECT 35.875 189.615 36.205 190.015 ;
        RECT 36.630 189.785 37.160 190.150 ;
        RECT 37.350 190.125 37.625 190.945 ;
        RECT 37.345 189.955 37.625 190.125 ;
        RECT 37.350 189.785 37.625 189.955 ;
        RECT 37.795 189.785 37.985 191.145 ;
        RECT 38.155 191.160 38.325 191.825 ;
        RECT 38.495 191.405 38.665 192.165 ;
        RECT 38.900 191.405 39.415 191.815 ;
        RECT 38.155 190.970 38.905 191.160 ;
        RECT 39.075 190.595 39.415 191.405 ;
        RECT 38.185 190.425 39.415 190.595 ;
        RECT 39.585 191.075 42.175 192.165 ;
        RECT 42.345 191.405 42.860 191.815 ;
        RECT 43.095 191.405 43.265 192.165 ;
        RECT 43.435 191.825 45.465 191.995 ;
        RECT 39.585 190.555 40.795 191.075 ;
        RECT 38.165 189.615 38.675 190.150 ;
        RECT 38.895 189.820 39.140 190.425 ;
        RECT 40.965 190.385 42.175 190.905 ;
        RECT 42.345 190.595 42.685 191.405 ;
        RECT 43.435 191.160 43.605 191.825 ;
        RECT 44.000 191.485 45.125 191.655 ;
        RECT 42.855 190.970 43.605 191.160 ;
        RECT 43.775 191.145 44.785 191.315 ;
        RECT 42.345 190.425 43.575 190.595 ;
        RECT 39.585 189.615 42.175 190.385 ;
        RECT 42.620 189.820 42.865 190.425 ;
        RECT 43.085 189.615 43.595 190.150 ;
        RECT 43.775 189.785 43.965 191.145 ;
        RECT 44.135 190.125 44.410 190.945 ;
        RECT 44.615 190.345 44.785 191.145 ;
        RECT 44.955 190.355 45.125 191.485 ;
        RECT 45.295 190.855 45.465 191.825 ;
        RECT 45.635 191.025 45.805 192.165 ;
        RECT 45.975 191.025 46.310 191.995 ;
        RECT 45.295 190.525 45.490 190.855 ;
        RECT 45.715 190.525 45.970 190.855 ;
        RECT 45.715 190.355 45.885 190.525 ;
        RECT 46.140 190.355 46.310 191.025 ;
        RECT 46.485 191.075 49.995 192.165 ;
        RECT 46.485 190.555 48.175 191.075 ;
        RECT 50.165 191.000 50.455 192.165 ;
        RECT 51.085 191.075 52.755 192.165 ;
        RECT 48.345 190.385 49.995 190.905 ;
        RECT 51.085 190.555 51.835 191.075 ;
        RECT 52.985 191.025 53.195 192.165 ;
        RECT 53.365 191.015 53.695 191.995 ;
        RECT 53.865 191.025 54.095 192.165 ;
        RECT 54.305 191.075 55.515 192.165 ;
        RECT 55.775 191.235 55.945 191.995 ;
        RECT 56.125 191.405 56.455 192.165 ;
        RECT 52.005 190.385 52.755 190.905 ;
        RECT 44.955 190.185 45.885 190.355 ;
        RECT 44.955 190.150 45.130 190.185 ;
        RECT 44.135 189.955 44.415 190.125 ;
        RECT 44.135 189.785 44.410 189.955 ;
        RECT 44.600 189.785 45.130 190.150 ;
        RECT 45.555 189.615 45.885 190.015 ;
        RECT 46.055 189.785 46.310 190.355 ;
        RECT 46.485 189.615 49.995 190.385 ;
        RECT 50.165 189.615 50.455 190.340 ;
        RECT 51.085 189.615 52.755 190.385 ;
        RECT 52.985 189.615 53.195 190.435 ;
        RECT 53.365 190.415 53.615 191.015 ;
        RECT 53.785 190.605 54.115 190.855 ;
        RECT 54.305 190.535 54.825 191.075 ;
        RECT 55.775 191.065 56.440 191.235 ;
        RECT 56.625 191.090 56.895 191.995 ;
        RECT 56.270 190.920 56.440 191.065 ;
        RECT 53.365 189.785 53.695 190.415 ;
        RECT 53.865 189.615 54.095 190.435 ;
        RECT 54.995 190.365 55.515 190.905 ;
        RECT 55.705 190.515 56.035 190.885 ;
        RECT 56.270 190.590 56.555 190.920 ;
        RECT 54.305 189.615 55.515 190.365 ;
        RECT 56.270 190.335 56.440 190.590 ;
        RECT 55.775 190.165 56.440 190.335 ;
        RECT 56.725 190.290 56.895 191.090 ;
        RECT 57.125 191.025 57.335 192.165 ;
        RECT 57.505 191.015 57.835 191.995 ;
        RECT 58.005 191.025 58.235 192.165 ;
        RECT 58.445 191.075 59.655 192.165 ;
        RECT 59.830 191.730 65.175 192.165 ;
        RECT 65.350 191.730 70.695 192.165 ;
        RECT 55.775 189.785 55.945 190.165 ;
        RECT 56.125 189.615 56.455 189.995 ;
        RECT 56.635 189.785 56.895 190.290 ;
        RECT 57.125 189.615 57.335 190.435 ;
        RECT 57.505 190.415 57.755 191.015 ;
        RECT 57.925 190.605 58.255 190.855 ;
        RECT 58.445 190.535 58.965 191.075 ;
        RECT 57.505 189.785 57.835 190.415 ;
        RECT 58.005 189.615 58.235 190.435 ;
        RECT 59.135 190.365 59.655 190.905 ;
        RECT 61.420 190.480 61.770 191.730 ;
        RECT 58.445 189.615 59.655 190.365 ;
        RECT 63.250 190.160 63.590 190.990 ;
        RECT 66.940 190.480 67.290 191.730 ;
        RECT 70.955 191.235 71.125 191.995 ;
        RECT 71.305 191.405 71.635 192.165 ;
        RECT 70.955 191.065 71.620 191.235 ;
        RECT 71.805 191.090 72.075 191.995 ;
        RECT 68.770 190.160 69.110 190.990 ;
        RECT 71.450 190.920 71.620 191.065 ;
        RECT 70.885 190.515 71.215 190.885 ;
        RECT 71.450 190.590 71.735 190.920 ;
        RECT 71.450 190.335 71.620 190.590 ;
        RECT 70.955 190.165 71.620 190.335 ;
        RECT 71.905 190.290 72.075 191.090 ;
        RECT 72.245 191.075 73.455 192.165 ;
        RECT 73.645 191.365 73.925 192.165 ;
        RECT 74.125 191.195 74.455 191.995 ;
        RECT 74.655 191.365 74.825 192.165 ;
        RECT 74.995 191.195 75.325 191.995 ;
        RECT 72.245 190.535 72.765 191.075 ;
        RECT 72.935 190.365 73.455 190.905 ;
        RECT 73.625 190.525 73.865 191.195 ;
        RECT 74.045 191.025 75.325 191.195 ;
        RECT 75.495 191.025 75.755 192.165 ;
        RECT 59.830 189.615 65.175 190.160 ;
        RECT 65.350 189.615 70.695 190.160 ;
        RECT 70.955 189.785 71.125 190.165 ;
        RECT 71.305 189.615 71.635 189.995 ;
        RECT 71.815 189.785 72.075 190.290 ;
        RECT 72.245 189.615 73.455 190.365 ;
        RECT 74.045 190.355 74.215 191.025 ;
        RECT 75.925 191.000 76.215 192.165 ;
        RECT 76.845 191.610 77.450 192.165 ;
        RECT 77.625 191.655 78.105 191.995 ;
        RECT 78.275 191.620 78.530 192.165 ;
        RECT 76.845 191.510 77.460 191.610 ;
        RECT 77.275 191.485 77.460 191.510 ;
        RECT 76.845 190.890 77.105 191.340 ;
        RECT 77.275 191.240 77.605 191.485 ;
        RECT 77.775 191.165 78.530 191.415 ;
        RECT 78.700 191.295 78.975 191.995 ;
        RECT 77.760 191.130 78.530 191.165 ;
        RECT 77.745 191.120 78.530 191.130 ;
        RECT 77.740 191.105 78.635 191.120 ;
        RECT 77.720 191.090 78.635 191.105 ;
        RECT 77.700 191.080 78.635 191.090 ;
        RECT 77.675 191.070 78.635 191.080 ;
        RECT 77.605 191.040 78.635 191.070 ;
        RECT 77.585 191.010 78.635 191.040 ;
        RECT 77.565 190.980 78.635 191.010 ;
        RECT 77.535 190.955 78.635 190.980 ;
        RECT 77.500 190.920 78.635 190.955 ;
        RECT 77.470 190.915 78.635 190.920 ;
        RECT 77.470 190.910 77.860 190.915 ;
        RECT 77.470 190.900 77.835 190.910 ;
        RECT 77.470 190.895 77.820 190.900 ;
        RECT 77.470 190.890 77.805 190.895 ;
        RECT 76.845 190.885 77.805 190.890 ;
        RECT 76.845 190.875 77.795 190.885 ;
        RECT 76.845 190.870 77.785 190.875 ;
        RECT 76.845 190.860 77.775 190.870 ;
        RECT 74.385 190.525 74.695 190.855 ;
        RECT 74.865 190.525 75.245 190.855 ;
        RECT 75.445 190.525 75.730 190.855 ;
        RECT 76.845 190.850 77.770 190.860 ;
        RECT 76.845 190.845 77.765 190.850 ;
        RECT 76.845 190.830 77.755 190.845 ;
        RECT 76.845 190.815 77.750 190.830 ;
        RECT 76.845 190.790 77.740 190.815 ;
        RECT 76.845 190.720 77.735 190.790 ;
        RECT 74.490 190.355 74.695 190.525 ;
        RECT 73.625 189.785 74.320 190.355 ;
        RECT 74.490 189.830 74.840 190.355 ;
        RECT 75.030 189.830 75.245 190.525 ;
        RECT 75.415 189.615 75.750 190.355 ;
        RECT 75.925 189.615 76.215 190.340 ;
        RECT 76.845 190.165 77.395 190.550 ;
        RECT 77.565 189.995 77.735 190.720 ;
        RECT 76.845 189.825 77.735 189.995 ;
        RECT 77.905 190.320 78.235 190.745 ;
        RECT 78.405 190.520 78.635 190.915 ;
        RECT 77.905 189.835 78.125 190.320 ;
        RECT 78.805 190.265 78.975 191.295 ;
        RECT 79.235 191.235 79.405 191.995 ;
        RECT 79.585 191.405 79.915 192.165 ;
        RECT 79.235 191.065 79.900 191.235 ;
        RECT 80.085 191.090 80.355 191.995 ;
        RECT 79.730 190.920 79.900 191.065 ;
        RECT 79.165 190.515 79.495 190.885 ;
        RECT 79.730 190.590 80.015 190.920 ;
        RECT 79.730 190.335 79.900 190.590 ;
        RECT 78.295 189.615 78.545 190.155 ;
        RECT 78.715 189.785 78.975 190.265 ;
        RECT 79.235 190.165 79.900 190.335 ;
        RECT 80.185 190.290 80.355 191.090 ;
        RECT 80.985 191.075 83.575 192.165 ;
        RECT 83.750 191.730 89.095 192.165 ;
        RECT 80.985 190.555 82.195 191.075 ;
        RECT 82.365 190.385 83.575 190.905 ;
        RECT 85.340 190.480 85.690 191.730 ;
        RECT 89.270 191.025 89.605 191.995 ;
        RECT 89.775 191.025 89.945 192.165 ;
        RECT 90.115 191.825 92.145 191.995 ;
        RECT 79.235 189.785 79.405 190.165 ;
        RECT 79.585 189.615 79.915 189.995 ;
        RECT 80.095 189.785 80.355 190.290 ;
        RECT 80.985 189.615 83.575 190.385 ;
        RECT 87.170 190.160 87.510 190.990 ;
        RECT 89.270 190.355 89.440 191.025 ;
        RECT 90.115 190.855 90.285 191.825 ;
        RECT 89.610 190.525 89.865 190.855 ;
        RECT 90.090 190.525 90.285 190.855 ;
        RECT 90.455 191.485 91.580 191.655 ;
        RECT 89.695 190.355 89.865 190.525 ;
        RECT 90.455 190.355 90.625 191.485 ;
        RECT 83.750 189.615 89.095 190.160 ;
        RECT 89.270 189.785 89.525 190.355 ;
        RECT 89.695 190.185 90.625 190.355 ;
        RECT 90.795 191.145 91.805 191.315 ;
        RECT 90.795 190.345 90.965 191.145 ;
        RECT 90.450 190.150 90.625 190.185 ;
        RECT 89.695 189.615 90.025 190.015 ;
        RECT 90.450 189.785 90.980 190.150 ;
        RECT 91.170 190.125 91.445 190.945 ;
        RECT 91.165 189.955 91.445 190.125 ;
        RECT 91.170 189.785 91.445 189.955 ;
        RECT 91.615 189.785 91.805 191.145 ;
        RECT 91.975 191.160 92.145 191.825 ;
        RECT 92.315 191.405 92.485 192.165 ;
        RECT 92.720 191.405 93.235 191.815 ;
        RECT 91.975 190.970 92.725 191.160 ;
        RECT 92.895 190.595 93.235 191.405 ;
        RECT 93.495 191.235 93.665 191.995 ;
        RECT 93.845 191.405 94.175 192.165 ;
        RECT 93.495 191.065 94.160 191.235 ;
        RECT 94.345 191.090 94.615 191.995 ;
        RECT 93.990 190.920 94.160 191.065 ;
        RECT 92.005 190.425 93.235 190.595 ;
        RECT 93.425 190.515 93.755 190.885 ;
        RECT 93.990 190.590 94.275 190.920 ;
        RECT 91.985 189.615 92.495 190.150 ;
        RECT 92.715 189.820 92.960 190.425 ;
        RECT 93.990 190.335 94.160 190.590 ;
        RECT 93.495 190.165 94.160 190.335 ;
        RECT 94.445 190.290 94.615 191.090 ;
        RECT 94.785 191.075 95.995 192.165 ;
        RECT 96.170 191.730 101.515 192.165 ;
        RECT 94.785 190.535 95.305 191.075 ;
        RECT 95.475 190.365 95.995 190.905 ;
        RECT 97.760 190.480 98.110 191.730 ;
        RECT 101.685 191.000 101.975 192.165 ;
        RECT 103.070 191.730 108.415 192.165 ;
        RECT 93.495 189.785 93.665 190.165 ;
        RECT 93.845 189.615 94.175 189.995 ;
        RECT 94.355 189.785 94.615 190.290 ;
        RECT 94.785 189.615 95.995 190.365 ;
        RECT 99.590 190.160 99.930 190.990 ;
        RECT 104.660 190.480 105.010 191.730 ;
        RECT 96.170 189.615 101.515 190.160 ;
        RECT 101.685 189.615 101.975 190.340 ;
        RECT 106.490 190.160 106.830 190.990 ;
        RECT 108.590 190.975 108.845 191.855 ;
        RECT 109.015 191.025 109.320 192.165 ;
        RECT 109.660 191.785 109.990 192.165 ;
        RECT 110.170 191.615 110.340 191.905 ;
        RECT 110.510 191.705 110.760 192.165 ;
        RECT 109.540 191.445 110.340 191.615 ;
        RECT 110.930 191.655 111.800 191.995 ;
        RECT 108.590 190.325 108.800 190.975 ;
        RECT 109.540 190.855 109.710 191.445 ;
        RECT 110.930 191.275 111.100 191.655 ;
        RECT 112.035 191.535 112.205 191.995 ;
        RECT 112.375 191.705 112.745 192.165 ;
        RECT 113.040 191.565 113.210 191.905 ;
        RECT 113.380 191.735 113.710 192.165 ;
        RECT 113.945 191.565 114.115 191.905 ;
        RECT 109.880 191.105 111.100 191.275 ;
        RECT 111.270 191.195 111.730 191.485 ;
        RECT 112.035 191.365 112.595 191.535 ;
        RECT 113.040 191.395 114.115 191.565 ;
        RECT 114.285 191.665 114.965 191.995 ;
        RECT 115.180 191.665 115.430 191.995 ;
        RECT 115.600 191.705 115.850 192.165 ;
        RECT 112.425 191.225 112.595 191.365 ;
        RECT 111.270 191.185 112.235 191.195 ;
        RECT 110.930 191.015 111.100 191.105 ;
        RECT 111.560 191.025 112.235 191.185 ;
        RECT 108.970 190.825 109.710 190.855 ;
        RECT 108.970 190.525 109.885 190.825 ;
        RECT 109.560 190.350 109.885 190.525 ;
        RECT 103.070 189.615 108.415 190.160 ;
        RECT 108.590 189.795 108.845 190.325 ;
        RECT 109.015 189.615 109.320 190.075 ;
        RECT 109.565 189.995 109.885 190.350 ;
        RECT 110.055 190.565 110.595 190.935 ;
        RECT 110.930 190.845 111.335 191.015 ;
        RECT 110.055 190.165 110.295 190.565 ;
        RECT 110.775 190.395 110.995 190.675 ;
        RECT 110.465 190.225 110.995 190.395 ;
        RECT 110.465 189.995 110.635 190.225 ;
        RECT 111.165 190.065 111.335 190.845 ;
        RECT 111.505 190.235 111.855 190.855 ;
        RECT 112.025 190.235 112.235 191.025 ;
        RECT 112.425 191.055 113.925 191.225 ;
        RECT 112.425 190.365 112.595 191.055 ;
        RECT 114.285 190.885 114.455 191.665 ;
        RECT 115.260 191.535 115.430 191.665 ;
        RECT 112.765 190.715 114.455 190.885 ;
        RECT 114.625 191.105 115.090 191.495 ;
        RECT 115.260 191.365 115.655 191.535 ;
        RECT 112.765 190.535 112.935 190.715 ;
        RECT 109.565 189.825 110.635 189.995 ;
        RECT 110.805 189.615 110.995 190.055 ;
        RECT 111.165 189.785 112.115 190.065 ;
        RECT 112.425 189.975 112.685 190.365 ;
        RECT 113.105 190.295 113.895 190.545 ;
        RECT 112.335 189.805 112.685 189.975 ;
        RECT 112.895 189.615 113.225 190.075 ;
        RECT 114.100 190.005 114.270 190.715 ;
        RECT 114.625 190.515 114.795 191.105 ;
        RECT 114.440 190.295 114.795 190.515 ;
        RECT 114.965 190.295 115.315 190.915 ;
        RECT 115.485 190.005 115.655 191.365 ;
        RECT 116.020 191.195 116.345 191.980 ;
        RECT 115.825 190.145 116.285 191.195 ;
        RECT 114.100 189.835 114.955 190.005 ;
        RECT 115.160 189.835 115.655 190.005 ;
        RECT 115.825 189.615 116.155 189.975 ;
        RECT 116.515 189.875 116.685 191.995 ;
        RECT 116.855 191.665 117.185 192.165 ;
        RECT 117.355 191.495 117.610 191.995 ;
        RECT 116.860 191.325 117.610 191.495 ;
        RECT 116.860 190.335 117.090 191.325 ;
        RECT 117.260 190.505 117.610 191.155 ;
        RECT 117.785 191.075 120.375 192.165 ;
        RECT 120.635 191.235 120.805 191.995 ;
        RECT 120.985 191.405 121.315 192.165 ;
        RECT 117.785 190.555 118.995 191.075 ;
        RECT 120.635 191.065 121.300 191.235 ;
        RECT 121.485 191.090 121.755 191.995 ;
        RECT 121.130 190.920 121.300 191.065 ;
        RECT 119.165 190.385 120.375 190.905 ;
        RECT 120.565 190.515 120.895 190.885 ;
        RECT 121.130 190.590 121.415 190.920 ;
        RECT 116.860 190.165 117.610 190.335 ;
        RECT 116.855 189.615 117.185 189.995 ;
        RECT 117.355 189.875 117.610 190.165 ;
        RECT 117.785 189.615 120.375 190.385 ;
        RECT 121.130 190.335 121.300 190.590 ;
        RECT 120.635 190.165 121.300 190.335 ;
        RECT 121.585 190.290 121.755 191.090 ;
        RECT 122.845 191.075 126.355 192.165 ;
        RECT 126.525 191.075 127.735 192.165 ;
        RECT 122.845 190.555 124.535 191.075 ;
        RECT 124.705 190.385 126.355 190.905 ;
        RECT 126.525 190.535 127.045 191.075 ;
        RECT 120.635 189.785 120.805 190.165 ;
        RECT 120.985 189.615 121.315 189.995 ;
        RECT 121.495 189.785 121.755 190.290 ;
        RECT 122.845 189.615 126.355 190.385 ;
        RECT 127.215 190.365 127.735 190.905 ;
        RECT 126.525 189.615 127.735 190.365 ;
        RECT 20.640 189.445 127.820 189.615 ;
        RECT 20.725 188.695 21.935 189.445 ;
        RECT 22.570 188.900 27.915 189.445 ;
        RECT 20.725 188.155 21.245 188.695 ;
        RECT 21.415 187.985 21.935 188.525 ;
        RECT 20.725 186.895 21.935 187.985 ;
        RECT 24.160 187.330 24.510 188.580 ;
        RECT 25.990 188.070 26.330 188.900 ;
        RECT 28.090 188.895 28.345 189.185 ;
        RECT 28.515 189.065 28.845 189.445 ;
        RECT 28.090 188.725 28.840 188.895 ;
        RECT 28.090 187.905 28.440 188.555 ;
        RECT 28.610 187.735 28.840 188.725 ;
        RECT 28.090 187.565 28.840 187.735 ;
        RECT 22.570 186.895 27.915 187.330 ;
        RECT 28.090 187.065 28.345 187.565 ;
        RECT 28.515 186.895 28.845 187.395 ;
        RECT 29.015 187.065 29.185 189.185 ;
        RECT 29.545 189.085 29.875 189.445 ;
        RECT 30.045 189.055 30.540 189.225 ;
        RECT 30.745 189.055 31.600 189.225 ;
        RECT 29.415 187.865 29.875 188.915 ;
        RECT 29.355 187.080 29.680 187.865 ;
        RECT 30.045 187.695 30.215 189.055 ;
        RECT 30.385 188.145 30.735 188.765 ;
        RECT 30.905 188.545 31.260 188.765 ;
        RECT 30.905 187.955 31.075 188.545 ;
        RECT 31.430 188.345 31.600 189.055 ;
        RECT 32.475 188.985 32.805 189.445 ;
        RECT 33.015 189.085 33.365 189.255 ;
        RECT 31.805 188.515 32.595 188.765 ;
        RECT 33.015 188.695 33.275 189.085 ;
        RECT 33.585 188.995 34.535 189.275 ;
        RECT 34.705 189.005 34.895 189.445 ;
        RECT 35.065 189.065 36.135 189.235 ;
        RECT 32.765 188.345 32.935 188.525 ;
        RECT 30.045 187.525 30.440 187.695 ;
        RECT 30.610 187.565 31.075 187.955 ;
        RECT 31.245 188.175 32.935 188.345 ;
        RECT 30.270 187.395 30.440 187.525 ;
        RECT 31.245 187.395 31.415 188.175 ;
        RECT 33.105 188.005 33.275 188.695 ;
        RECT 31.775 187.835 33.275 188.005 ;
        RECT 33.465 188.035 33.675 188.825 ;
        RECT 33.845 188.205 34.195 188.825 ;
        RECT 34.365 188.215 34.535 188.995 ;
        RECT 35.065 188.835 35.235 189.065 ;
        RECT 34.705 188.665 35.235 188.835 ;
        RECT 34.705 188.385 34.925 188.665 ;
        RECT 35.405 188.495 35.645 188.895 ;
        RECT 34.365 188.045 34.770 188.215 ;
        RECT 35.105 188.125 35.645 188.495 ;
        RECT 35.815 188.710 36.135 189.065 ;
        RECT 36.380 188.985 36.685 189.445 ;
        RECT 36.855 188.735 37.110 189.265 ;
        RECT 35.815 188.535 36.140 188.710 ;
        RECT 35.815 188.235 36.730 188.535 ;
        RECT 35.990 188.205 36.730 188.235 ;
        RECT 33.465 187.875 34.140 188.035 ;
        RECT 34.600 187.955 34.770 188.045 ;
        RECT 33.465 187.865 34.430 187.875 ;
        RECT 33.105 187.695 33.275 187.835 ;
        RECT 29.850 186.895 30.100 187.355 ;
        RECT 30.270 187.065 30.520 187.395 ;
        RECT 30.735 187.065 31.415 187.395 ;
        RECT 31.585 187.495 32.660 187.665 ;
        RECT 33.105 187.525 33.665 187.695 ;
        RECT 33.970 187.575 34.430 187.865 ;
        RECT 34.600 187.785 35.820 187.955 ;
        RECT 31.585 187.155 31.755 187.495 ;
        RECT 31.990 186.895 32.320 187.325 ;
        RECT 32.490 187.155 32.660 187.495 ;
        RECT 32.955 186.895 33.325 187.355 ;
        RECT 33.495 187.065 33.665 187.525 ;
        RECT 34.600 187.405 34.770 187.785 ;
        RECT 35.990 187.615 36.160 188.205 ;
        RECT 36.900 188.085 37.110 188.735 ;
        RECT 37.285 188.720 37.575 189.445 ;
        RECT 38.210 188.900 43.555 189.445 ;
        RECT 43.730 188.900 49.075 189.445 ;
        RECT 33.900 187.065 34.770 187.405 ;
        RECT 35.360 187.445 36.160 187.615 ;
        RECT 34.940 186.895 35.190 187.355 ;
        RECT 35.360 187.155 35.530 187.445 ;
        RECT 35.710 186.895 36.040 187.275 ;
        RECT 36.380 186.895 36.685 188.035 ;
        RECT 36.855 187.205 37.110 188.085 ;
        RECT 37.285 186.895 37.575 188.060 ;
        RECT 39.800 187.330 40.150 188.580 ;
        RECT 41.630 188.070 41.970 188.900 ;
        RECT 45.320 187.330 45.670 188.580 ;
        RECT 47.150 188.070 47.490 188.900 ;
        RECT 49.250 188.735 49.505 189.265 ;
        RECT 49.675 188.985 49.980 189.445 ;
        RECT 50.225 189.065 51.295 189.235 ;
        RECT 49.250 188.085 49.460 188.735 ;
        RECT 50.225 188.710 50.545 189.065 ;
        RECT 50.220 188.535 50.545 188.710 ;
        RECT 49.630 188.235 50.545 188.535 ;
        RECT 50.715 188.495 50.955 188.895 ;
        RECT 51.125 188.835 51.295 189.065 ;
        RECT 51.465 189.005 51.655 189.445 ;
        RECT 51.825 188.995 52.775 189.275 ;
        RECT 52.995 189.085 53.345 189.255 ;
        RECT 51.125 188.665 51.655 188.835 ;
        RECT 49.630 188.205 50.370 188.235 ;
        RECT 38.210 186.895 43.555 187.330 ;
        RECT 43.730 186.895 49.075 187.330 ;
        RECT 49.250 187.205 49.505 188.085 ;
        RECT 49.675 186.895 49.980 188.035 ;
        RECT 50.200 187.615 50.370 188.205 ;
        RECT 50.715 188.125 51.255 188.495 ;
        RECT 51.435 188.385 51.655 188.665 ;
        RECT 51.825 188.215 51.995 188.995 ;
        RECT 51.590 188.045 51.995 188.215 ;
        RECT 52.165 188.205 52.515 188.825 ;
        RECT 51.590 187.955 51.760 188.045 ;
        RECT 52.685 188.035 52.895 188.825 ;
        RECT 50.540 187.785 51.760 187.955 ;
        RECT 52.220 187.875 52.895 188.035 ;
        RECT 50.200 187.445 51.000 187.615 ;
        RECT 50.320 186.895 50.650 187.275 ;
        RECT 50.830 187.155 51.000 187.445 ;
        RECT 51.590 187.405 51.760 187.785 ;
        RECT 51.930 187.865 52.895 187.875 ;
        RECT 53.085 188.695 53.345 189.085 ;
        RECT 53.555 188.985 53.885 189.445 ;
        RECT 54.760 189.055 55.615 189.225 ;
        RECT 55.820 189.055 56.315 189.225 ;
        RECT 56.485 189.085 56.815 189.445 ;
        RECT 53.085 188.005 53.255 188.695 ;
        RECT 53.425 188.345 53.595 188.525 ;
        RECT 53.765 188.515 54.555 188.765 ;
        RECT 54.760 188.345 54.930 189.055 ;
        RECT 55.100 188.545 55.455 188.765 ;
        RECT 53.425 188.175 55.115 188.345 ;
        RECT 51.930 187.575 52.390 187.865 ;
        RECT 53.085 187.835 54.585 188.005 ;
        RECT 53.085 187.695 53.255 187.835 ;
        RECT 52.695 187.525 53.255 187.695 ;
        RECT 51.170 186.895 51.420 187.355 ;
        RECT 51.590 187.065 52.460 187.405 ;
        RECT 52.695 187.065 52.865 187.525 ;
        RECT 53.700 187.495 54.775 187.665 ;
        RECT 53.035 186.895 53.405 187.355 ;
        RECT 53.700 187.155 53.870 187.495 ;
        RECT 54.040 186.895 54.370 187.325 ;
        RECT 54.605 187.155 54.775 187.495 ;
        RECT 54.945 187.395 55.115 188.175 ;
        RECT 55.285 187.955 55.455 188.545 ;
        RECT 55.625 188.145 55.975 188.765 ;
        RECT 55.285 187.565 55.750 187.955 ;
        RECT 56.145 187.695 56.315 189.055 ;
        RECT 56.485 187.865 56.945 188.915 ;
        RECT 55.920 187.525 56.315 187.695 ;
        RECT 55.920 187.395 56.090 187.525 ;
        RECT 54.945 187.065 55.625 187.395 ;
        RECT 55.840 187.065 56.090 187.395 ;
        RECT 56.260 186.895 56.510 187.355 ;
        RECT 56.680 187.080 57.005 187.865 ;
        RECT 57.175 187.065 57.345 189.185 ;
        RECT 57.515 189.065 57.845 189.445 ;
        RECT 58.015 188.895 58.270 189.185 ;
        RECT 57.520 188.725 58.270 188.895 ;
        RECT 57.520 187.735 57.750 188.725 ;
        RECT 58.505 188.625 58.715 189.445 ;
        RECT 58.885 188.645 59.215 189.275 ;
        RECT 57.920 187.905 58.270 188.555 ;
        RECT 58.885 188.045 59.135 188.645 ;
        RECT 59.385 188.625 59.615 189.445 ;
        RECT 60.285 188.675 62.875 189.445 ;
        RECT 63.045 188.720 63.335 189.445 ;
        RECT 63.965 188.675 66.555 189.445 ;
        RECT 66.730 188.900 72.075 189.445 ;
        RECT 59.305 188.205 59.635 188.455 ;
        RECT 57.520 187.565 58.270 187.735 ;
        RECT 57.515 186.895 57.845 187.395 ;
        RECT 58.015 187.065 58.270 187.565 ;
        RECT 58.505 186.895 58.715 188.035 ;
        RECT 58.885 187.065 59.215 188.045 ;
        RECT 59.385 186.895 59.615 188.035 ;
        RECT 60.285 187.985 61.495 188.505 ;
        RECT 61.665 188.155 62.875 188.675 ;
        RECT 60.285 186.895 62.875 187.985 ;
        RECT 63.045 186.895 63.335 188.060 ;
        RECT 63.965 187.985 65.175 188.505 ;
        RECT 65.345 188.155 66.555 188.675 ;
        RECT 63.965 186.895 66.555 187.985 ;
        RECT 68.320 187.330 68.670 188.580 ;
        RECT 70.150 188.070 70.490 188.900 ;
        RECT 72.285 188.625 72.515 189.445 ;
        RECT 72.685 188.645 73.015 189.275 ;
        RECT 72.265 188.205 72.595 188.455 ;
        RECT 72.765 188.045 73.015 188.645 ;
        RECT 73.185 188.625 73.395 189.445 ;
        RECT 73.630 188.735 73.885 189.265 ;
        RECT 74.055 188.985 74.360 189.445 ;
        RECT 74.605 189.065 75.675 189.235 ;
        RECT 66.730 186.895 72.075 187.330 ;
        RECT 72.285 186.895 72.515 188.035 ;
        RECT 72.685 187.065 73.015 188.045 ;
        RECT 73.630 188.085 73.840 188.735 ;
        RECT 74.605 188.710 74.925 189.065 ;
        RECT 74.600 188.535 74.925 188.710 ;
        RECT 74.010 188.235 74.925 188.535 ;
        RECT 75.095 188.495 75.335 188.895 ;
        RECT 75.505 188.835 75.675 189.065 ;
        RECT 75.845 189.005 76.035 189.445 ;
        RECT 76.205 188.995 77.155 189.275 ;
        RECT 77.375 189.085 77.725 189.255 ;
        RECT 75.505 188.665 76.035 188.835 ;
        RECT 74.010 188.205 74.750 188.235 ;
        RECT 73.185 186.895 73.395 188.035 ;
        RECT 73.630 187.205 73.885 188.085 ;
        RECT 74.055 186.895 74.360 188.035 ;
        RECT 74.580 187.615 74.750 188.205 ;
        RECT 75.095 188.125 75.635 188.495 ;
        RECT 75.815 188.385 76.035 188.665 ;
        RECT 76.205 188.215 76.375 188.995 ;
        RECT 75.970 188.045 76.375 188.215 ;
        RECT 76.545 188.205 76.895 188.825 ;
        RECT 75.970 187.955 76.140 188.045 ;
        RECT 77.065 188.035 77.275 188.825 ;
        RECT 74.920 187.785 76.140 187.955 ;
        RECT 76.600 187.875 77.275 188.035 ;
        RECT 74.580 187.445 75.380 187.615 ;
        RECT 74.700 186.895 75.030 187.275 ;
        RECT 75.210 187.155 75.380 187.445 ;
        RECT 75.970 187.405 76.140 187.785 ;
        RECT 76.310 187.865 77.275 187.875 ;
        RECT 77.465 188.695 77.725 189.085 ;
        RECT 77.935 188.985 78.265 189.445 ;
        RECT 79.140 189.055 79.995 189.225 ;
        RECT 80.200 189.055 80.695 189.225 ;
        RECT 80.865 189.085 81.195 189.445 ;
        RECT 77.465 188.005 77.635 188.695 ;
        RECT 77.805 188.345 77.975 188.525 ;
        RECT 78.145 188.515 78.935 188.765 ;
        RECT 79.140 188.345 79.310 189.055 ;
        RECT 79.480 188.545 79.835 188.765 ;
        RECT 77.805 188.175 79.495 188.345 ;
        RECT 76.310 187.575 76.770 187.865 ;
        RECT 77.465 187.835 78.965 188.005 ;
        RECT 77.465 187.695 77.635 187.835 ;
        RECT 77.075 187.525 77.635 187.695 ;
        RECT 75.550 186.895 75.800 187.355 ;
        RECT 75.970 187.065 76.840 187.405 ;
        RECT 77.075 187.065 77.245 187.525 ;
        RECT 78.080 187.495 79.155 187.665 ;
        RECT 77.415 186.895 77.785 187.355 ;
        RECT 78.080 187.155 78.250 187.495 ;
        RECT 78.420 186.895 78.750 187.325 ;
        RECT 78.985 187.155 79.155 187.495 ;
        RECT 79.325 187.395 79.495 188.175 ;
        RECT 79.665 187.955 79.835 188.545 ;
        RECT 80.005 188.145 80.355 188.765 ;
        RECT 79.665 187.565 80.130 187.955 ;
        RECT 80.525 187.695 80.695 189.055 ;
        RECT 80.865 187.865 81.325 188.915 ;
        RECT 80.300 187.525 80.695 187.695 ;
        RECT 80.300 187.395 80.470 187.525 ;
        RECT 79.325 187.065 80.005 187.395 ;
        RECT 80.220 187.065 80.470 187.395 ;
        RECT 80.640 186.895 80.890 187.355 ;
        RECT 81.060 187.080 81.385 187.865 ;
        RECT 81.555 187.065 81.725 189.185 ;
        RECT 81.895 189.065 82.225 189.445 ;
        RECT 82.395 188.895 82.650 189.185 ;
        RECT 81.900 188.725 82.650 188.895 ;
        RECT 81.900 187.735 82.130 188.725 ;
        RECT 82.825 188.675 84.495 189.445 ;
        RECT 82.300 187.905 82.650 188.555 ;
        RECT 82.825 187.985 83.575 188.505 ;
        RECT 83.745 188.155 84.495 188.675 ;
        RECT 84.940 188.635 85.185 189.240 ;
        RECT 85.405 188.910 85.915 189.445 ;
        RECT 84.665 188.465 85.895 188.635 ;
        RECT 81.900 187.565 82.650 187.735 ;
        RECT 81.895 186.895 82.225 187.395 ;
        RECT 82.395 187.065 82.650 187.565 ;
        RECT 82.825 186.895 84.495 187.985 ;
        RECT 84.665 187.655 85.005 188.465 ;
        RECT 85.175 187.900 85.925 188.090 ;
        RECT 84.665 187.245 85.180 187.655 ;
        RECT 85.415 186.895 85.585 187.655 ;
        RECT 85.755 187.235 85.925 187.900 ;
        RECT 86.095 187.915 86.285 189.275 ;
        RECT 86.455 188.765 86.730 189.275 ;
        RECT 86.920 188.910 87.450 189.275 ;
        RECT 87.875 189.045 88.205 189.445 ;
        RECT 87.275 188.875 87.450 188.910 ;
        RECT 86.455 188.595 86.735 188.765 ;
        RECT 86.455 188.115 86.730 188.595 ;
        RECT 86.935 187.915 87.105 188.715 ;
        RECT 86.095 187.745 87.105 187.915 ;
        RECT 87.275 188.705 88.205 188.875 ;
        RECT 88.375 188.705 88.630 189.275 ;
        RECT 88.805 188.720 89.095 189.445 ;
        RECT 87.275 187.575 87.445 188.705 ;
        RECT 88.035 188.535 88.205 188.705 ;
        RECT 86.320 187.405 87.445 187.575 ;
        RECT 87.615 188.205 87.810 188.535 ;
        RECT 88.035 188.205 88.290 188.535 ;
        RECT 87.615 187.235 87.785 188.205 ;
        RECT 88.460 188.035 88.630 188.705 ;
        RECT 89.265 188.695 90.475 189.445 ;
        RECT 85.755 187.065 87.785 187.235 ;
        RECT 87.955 186.895 88.125 188.035 ;
        RECT 88.295 187.065 88.630 188.035 ;
        RECT 88.805 186.895 89.095 188.060 ;
        RECT 89.265 187.985 89.785 188.525 ;
        RECT 89.955 188.155 90.475 188.695 ;
        RECT 90.705 188.625 90.915 189.445 ;
        RECT 91.085 188.645 91.415 189.275 ;
        RECT 91.085 188.045 91.335 188.645 ;
        RECT 91.585 188.625 91.815 189.445 ;
        RECT 92.950 188.900 98.295 189.445 ;
        RECT 91.505 188.205 91.835 188.455 ;
        RECT 89.265 186.895 90.475 187.985 ;
        RECT 90.705 186.895 90.915 188.035 ;
        RECT 91.085 187.065 91.415 188.045 ;
        RECT 91.585 186.895 91.815 188.035 ;
        RECT 94.540 187.330 94.890 188.580 ;
        RECT 96.370 188.070 96.710 188.900 ;
        RECT 98.505 188.625 98.735 189.445 ;
        RECT 98.905 188.645 99.235 189.275 ;
        RECT 98.485 188.205 98.815 188.455 ;
        RECT 98.985 188.045 99.235 188.645 ;
        RECT 99.405 188.625 99.615 189.445 ;
        RECT 99.850 188.735 100.105 189.265 ;
        RECT 100.275 188.985 100.580 189.445 ;
        RECT 100.825 189.065 101.895 189.235 ;
        RECT 92.950 186.895 98.295 187.330 ;
        RECT 98.505 186.895 98.735 188.035 ;
        RECT 98.905 187.065 99.235 188.045 ;
        RECT 99.850 188.085 100.060 188.735 ;
        RECT 100.825 188.710 101.145 189.065 ;
        RECT 100.820 188.535 101.145 188.710 ;
        RECT 100.230 188.235 101.145 188.535 ;
        RECT 101.315 188.495 101.555 188.895 ;
        RECT 101.725 188.835 101.895 189.065 ;
        RECT 102.065 189.005 102.255 189.445 ;
        RECT 102.425 188.995 103.375 189.275 ;
        RECT 103.595 189.085 103.945 189.255 ;
        RECT 101.725 188.665 102.255 188.835 ;
        RECT 100.230 188.205 100.970 188.235 ;
        RECT 99.405 186.895 99.615 188.035 ;
        RECT 99.850 187.205 100.105 188.085 ;
        RECT 100.275 186.895 100.580 188.035 ;
        RECT 100.800 187.615 100.970 188.205 ;
        RECT 101.315 188.125 101.855 188.495 ;
        RECT 102.035 188.385 102.255 188.665 ;
        RECT 102.425 188.215 102.595 188.995 ;
        RECT 102.190 188.045 102.595 188.215 ;
        RECT 102.765 188.205 103.115 188.825 ;
        RECT 102.190 187.955 102.360 188.045 ;
        RECT 103.285 188.035 103.495 188.825 ;
        RECT 101.140 187.785 102.360 187.955 ;
        RECT 102.820 187.875 103.495 188.035 ;
        RECT 100.800 187.445 101.600 187.615 ;
        RECT 100.920 186.895 101.250 187.275 ;
        RECT 101.430 187.155 101.600 187.445 ;
        RECT 102.190 187.405 102.360 187.785 ;
        RECT 102.530 187.865 103.495 187.875 ;
        RECT 103.685 188.695 103.945 189.085 ;
        RECT 104.155 188.985 104.485 189.445 ;
        RECT 105.360 189.055 106.215 189.225 ;
        RECT 106.420 189.055 106.915 189.225 ;
        RECT 107.085 189.085 107.415 189.445 ;
        RECT 103.685 188.005 103.855 188.695 ;
        RECT 104.025 188.345 104.195 188.525 ;
        RECT 104.365 188.515 105.155 188.765 ;
        RECT 105.360 188.345 105.530 189.055 ;
        RECT 105.700 188.545 106.055 188.765 ;
        RECT 104.025 188.175 105.715 188.345 ;
        RECT 102.530 187.575 102.990 187.865 ;
        RECT 103.685 187.835 105.185 188.005 ;
        RECT 103.685 187.695 103.855 187.835 ;
        RECT 103.295 187.525 103.855 187.695 ;
        RECT 101.770 186.895 102.020 187.355 ;
        RECT 102.190 187.065 103.060 187.405 ;
        RECT 103.295 187.065 103.465 187.525 ;
        RECT 104.300 187.495 105.375 187.665 ;
        RECT 103.635 186.895 104.005 187.355 ;
        RECT 104.300 187.155 104.470 187.495 ;
        RECT 104.640 186.895 104.970 187.325 ;
        RECT 105.205 187.155 105.375 187.495 ;
        RECT 105.545 187.395 105.715 188.175 ;
        RECT 105.885 187.955 106.055 188.545 ;
        RECT 106.225 188.145 106.575 188.765 ;
        RECT 105.885 187.565 106.350 187.955 ;
        RECT 106.745 187.695 106.915 189.055 ;
        RECT 107.085 187.865 107.545 188.915 ;
        RECT 106.520 187.525 106.915 187.695 ;
        RECT 106.520 187.395 106.690 187.525 ;
        RECT 105.545 187.065 106.225 187.395 ;
        RECT 106.440 187.065 106.690 187.395 ;
        RECT 106.860 186.895 107.110 187.355 ;
        RECT 107.280 187.080 107.605 187.865 ;
        RECT 107.775 187.065 107.945 189.185 ;
        RECT 108.115 189.065 108.445 189.445 ;
        RECT 108.615 188.895 108.870 189.185 ;
        RECT 108.120 188.725 108.870 188.895 ;
        RECT 109.045 188.770 109.305 189.275 ;
        RECT 109.485 189.065 109.815 189.445 ;
        RECT 109.995 188.895 110.165 189.275 ;
        RECT 108.120 187.735 108.350 188.725 ;
        RECT 108.520 187.905 108.870 188.555 ;
        RECT 109.045 187.970 109.215 188.770 ;
        RECT 109.500 188.725 110.165 188.895 ;
        RECT 109.500 188.470 109.670 188.725 ;
        RECT 111.405 188.625 111.615 189.445 ;
        RECT 111.785 188.645 112.115 189.275 ;
        RECT 109.385 188.140 109.670 188.470 ;
        RECT 109.905 188.175 110.235 188.545 ;
        RECT 109.500 187.995 109.670 188.140 ;
        RECT 111.785 188.045 112.035 188.645 ;
        RECT 112.285 188.625 112.515 189.445 ;
        RECT 113.225 188.625 113.455 189.445 ;
        RECT 113.625 188.645 113.955 189.275 ;
        RECT 112.205 188.205 112.535 188.455 ;
        RECT 113.205 188.205 113.535 188.455 ;
        RECT 113.705 188.045 113.955 188.645 ;
        RECT 114.125 188.625 114.335 189.445 ;
        RECT 114.565 188.720 114.855 189.445 ;
        RECT 115.950 188.735 116.205 189.265 ;
        RECT 116.375 188.985 116.680 189.445 ;
        RECT 116.925 189.065 117.995 189.235 ;
        RECT 115.950 188.085 116.160 188.735 ;
        RECT 116.925 188.710 117.245 189.065 ;
        RECT 116.920 188.535 117.245 188.710 ;
        RECT 116.330 188.235 117.245 188.535 ;
        RECT 117.415 188.495 117.655 188.895 ;
        RECT 117.825 188.835 117.995 189.065 ;
        RECT 118.165 189.005 118.355 189.445 ;
        RECT 118.525 188.995 119.475 189.275 ;
        RECT 119.695 189.085 120.045 189.255 ;
        RECT 117.825 188.665 118.355 188.835 ;
        RECT 116.330 188.205 117.070 188.235 ;
        RECT 108.120 187.565 108.870 187.735 ;
        RECT 108.115 186.895 108.445 187.395 ;
        RECT 108.615 187.065 108.870 187.565 ;
        RECT 109.045 187.065 109.315 187.970 ;
        RECT 109.500 187.825 110.165 187.995 ;
        RECT 109.485 186.895 109.815 187.655 ;
        RECT 109.995 187.065 110.165 187.825 ;
        RECT 111.405 186.895 111.615 188.035 ;
        RECT 111.785 187.065 112.115 188.045 ;
        RECT 112.285 186.895 112.515 188.035 ;
        RECT 113.225 186.895 113.455 188.035 ;
        RECT 113.625 187.065 113.955 188.045 ;
        RECT 114.125 186.895 114.335 188.035 ;
        RECT 114.565 186.895 114.855 188.060 ;
        RECT 115.950 187.205 116.205 188.085 ;
        RECT 116.375 186.895 116.680 188.035 ;
        RECT 116.900 187.615 117.070 188.205 ;
        RECT 117.415 188.125 117.955 188.495 ;
        RECT 118.135 188.385 118.355 188.665 ;
        RECT 118.525 188.215 118.695 188.995 ;
        RECT 118.290 188.045 118.695 188.215 ;
        RECT 118.865 188.205 119.215 188.825 ;
        RECT 118.290 187.955 118.460 188.045 ;
        RECT 119.385 188.035 119.595 188.825 ;
        RECT 117.240 187.785 118.460 187.955 ;
        RECT 118.920 187.875 119.595 188.035 ;
        RECT 116.900 187.445 117.700 187.615 ;
        RECT 117.020 186.895 117.350 187.275 ;
        RECT 117.530 187.155 117.700 187.445 ;
        RECT 118.290 187.405 118.460 187.785 ;
        RECT 118.630 187.865 119.595 187.875 ;
        RECT 119.785 188.695 120.045 189.085 ;
        RECT 120.255 188.985 120.585 189.445 ;
        RECT 121.460 189.055 122.315 189.225 ;
        RECT 122.520 189.055 123.015 189.225 ;
        RECT 123.185 189.085 123.515 189.445 ;
        RECT 119.785 188.005 119.955 188.695 ;
        RECT 120.125 188.345 120.295 188.525 ;
        RECT 120.465 188.515 121.255 188.765 ;
        RECT 121.460 188.345 121.630 189.055 ;
        RECT 121.800 188.545 122.155 188.765 ;
        RECT 120.125 188.175 121.815 188.345 ;
        RECT 118.630 187.575 119.090 187.865 ;
        RECT 119.785 187.835 121.285 188.005 ;
        RECT 119.785 187.695 119.955 187.835 ;
        RECT 119.395 187.525 119.955 187.695 ;
        RECT 117.870 186.895 118.120 187.355 ;
        RECT 118.290 187.065 119.160 187.405 ;
        RECT 119.395 187.065 119.565 187.525 ;
        RECT 120.400 187.495 121.475 187.665 ;
        RECT 119.735 186.895 120.105 187.355 ;
        RECT 120.400 187.155 120.570 187.495 ;
        RECT 120.740 186.895 121.070 187.325 ;
        RECT 121.305 187.155 121.475 187.495 ;
        RECT 121.645 187.395 121.815 188.175 ;
        RECT 121.985 187.955 122.155 188.545 ;
        RECT 122.325 188.145 122.675 188.765 ;
        RECT 121.985 187.565 122.450 187.955 ;
        RECT 122.845 187.695 123.015 189.055 ;
        RECT 123.185 187.865 123.645 188.915 ;
        RECT 122.620 187.525 123.015 187.695 ;
        RECT 122.620 187.395 122.790 187.525 ;
        RECT 121.645 187.065 122.325 187.395 ;
        RECT 122.540 187.065 122.790 187.395 ;
        RECT 122.960 186.895 123.210 187.355 ;
        RECT 123.380 187.080 123.705 187.865 ;
        RECT 123.875 187.065 124.045 189.185 ;
        RECT 124.215 189.065 124.545 189.445 ;
        RECT 124.715 188.895 124.970 189.185 ;
        RECT 124.220 188.725 124.970 188.895 ;
        RECT 124.220 187.735 124.450 188.725 ;
        RECT 125.145 188.695 126.355 189.445 ;
        RECT 126.525 188.695 127.735 189.445 ;
        RECT 124.620 187.905 124.970 188.555 ;
        RECT 125.145 187.985 125.665 188.525 ;
        RECT 125.835 188.155 126.355 188.695 ;
        RECT 126.525 187.985 127.045 188.525 ;
        RECT 127.215 188.155 127.735 188.695 ;
        RECT 124.220 187.565 124.970 187.735 ;
        RECT 124.215 186.895 124.545 187.395 ;
        RECT 124.715 187.065 124.970 187.565 ;
        RECT 125.145 186.895 126.355 187.985 ;
        RECT 126.525 186.895 127.735 187.985 ;
        RECT 20.640 186.725 127.820 186.895 ;
        RECT 20.725 185.635 21.935 186.725 ;
        RECT 20.725 184.925 21.245 185.465 ;
        RECT 21.415 185.095 21.935 185.635 ;
        RECT 22.565 185.635 24.235 186.725 ;
        RECT 22.565 185.115 23.315 185.635 ;
        RECT 24.405 185.560 24.695 186.725 ;
        RECT 25.790 186.290 31.135 186.725 ;
        RECT 23.485 184.945 24.235 185.465 ;
        RECT 27.380 185.040 27.730 186.290 ;
        RECT 31.345 185.585 31.575 186.725 ;
        RECT 31.745 185.575 32.075 186.555 ;
        RECT 32.245 185.585 32.455 186.725 ;
        RECT 33.145 185.650 33.415 186.555 ;
        RECT 33.585 185.965 33.915 186.725 ;
        RECT 34.095 185.795 34.265 186.555 ;
        RECT 20.725 184.175 21.935 184.925 ;
        RECT 22.565 184.175 24.235 184.945 ;
        RECT 24.405 184.175 24.695 184.900 ;
        RECT 29.210 184.720 29.550 185.550 ;
        RECT 31.325 185.165 31.655 185.415 ;
        RECT 25.790 184.175 31.135 184.720 ;
        RECT 31.345 184.175 31.575 184.995 ;
        RECT 31.825 184.975 32.075 185.575 ;
        RECT 31.745 184.345 32.075 184.975 ;
        RECT 32.245 184.175 32.455 184.995 ;
        RECT 33.145 184.850 33.315 185.650 ;
        RECT 33.600 185.625 34.265 185.795 ;
        RECT 33.600 185.480 33.770 185.625 ;
        RECT 33.485 185.150 33.770 185.480 ;
        RECT 34.530 185.585 34.865 186.555 ;
        RECT 35.035 185.585 35.205 186.725 ;
        RECT 35.375 186.385 37.405 186.555 ;
        RECT 33.600 184.895 33.770 185.150 ;
        RECT 34.005 185.075 34.335 185.445 ;
        RECT 34.530 184.915 34.700 185.585 ;
        RECT 35.375 185.415 35.545 186.385 ;
        RECT 34.870 185.085 35.125 185.415 ;
        RECT 35.350 185.085 35.545 185.415 ;
        RECT 35.715 186.045 36.840 186.215 ;
        RECT 34.955 184.915 35.125 185.085 ;
        RECT 35.715 184.915 35.885 186.045 ;
        RECT 33.145 184.345 33.405 184.850 ;
        RECT 33.600 184.725 34.265 184.895 ;
        RECT 33.585 184.175 33.915 184.555 ;
        RECT 34.095 184.345 34.265 184.725 ;
        RECT 34.530 184.345 34.785 184.915 ;
        RECT 34.955 184.745 35.885 184.915 ;
        RECT 36.055 185.705 37.065 185.875 ;
        RECT 36.055 184.905 36.225 185.705 ;
        RECT 36.430 185.025 36.705 185.505 ;
        RECT 36.425 184.855 36.705 185.025 ;
        RECT 35.710 184.710 35.885 184.745 ;
        RECT 34.955 184.175 35.285 184.575 ;
        RECT 35.710 184.345 36.240 184.710 ;
        RECT 36.430 184.345 36.705 184.855 ;
        RECT 36.875 184.345 37.065 185.705 ;
        RECT 37.235 185.720 37.405 186.385 ;
        RECT 37.575 185.965 37.745 186.725 ;
        RECT 37.980 185.965 38.495 186.375 ;
        RECT 37.235 185.530 37.985 185.720 ;
        RECT 38.155 185.155 38.495 185.965 ;
        RECT 37.265 184.985 38.495 185.155 ;
        RECT 38.665 185.635 39.875 186.725 ;
        RECT 40.045 185.635 43.555 186.725 ;
        RECT 38.665 185.095 39.185 185.635 ;
        RECT 37.245 184.175 37.755 184.710 ;
        RECT 37.975 184.380 38.220 184.985 ;
        RECT 39.355 184.925 39.875 185.465 ;
        RECT 40.045 185.115 41.735 185.635 ;
        RECT 43.785 185.585 43.995 186.725 ;
        RECT 44.165 185.575 44.495 186.555 ;
        RECT 44.665 185.585 44.895 186.725 ;
        RECT 46.025 185.965 46.540 186.375 ;
        RECT 46.775 185.965 46.945 186.725 ;
        RECT 47.115 186.385 49.145 186.555 ;
        RECT 41.905 184.945 43.555 185.465 ;
        RECT 38.665 184.175 39.875 184.925 ;
        RECT 40.045 184.175 43.555 184.945 ;
        RECT 43.785 184.175 43.995 184.995 ;
        RECT 44.165 184.975 44.415 185.575 ;
        RECT 44.585 185.165 44.915 185.415 ;
        RECT 46.025 185.155 46.365 185.965 ;
        RECT 47.115 185.720 47.285 186.385 ;
        RECT 47.680 186.045 48.805 186.215 ;
        RECT 46.535 185.530 47.285 185.720 ;
        RECT 47.455 185.705 48.465 185.875 ;
        RECT 44.165 184.345 44.495 184.975 ;
        RECT 44.665 184.175 44.895 184.995 ;
        RECT 46.025 184.985 47.255 185.155 ;
        RECT 46.300 184.380 46.545 184.985 ;
        RECT 46.765 184.175 47.275 184.710 ;
        RECT 47.455 184.345 47.645 185.705 ;
        RECT 47.815 184.685 48.090 185.505 ;
        RECT 48.295 184.905 48.465 185.705 ;
        RECT 48.635 184.915 48.805 186.045 ;
        RECT 48.975 185.415 49.145 186.385 ;
        RECT 49.315 185.585 49.485 186.725 ;
        RECT 49.655 185.585 49.990 186.555 ;
        RECT 48.975 185.085 49.170 185.415 ;
        RECT 49.395 185.085 49.650 185.415 ;
        RECT 49.395 184.915 49.565 185.085 ;
        RECT 49.820 184.915 49.990 185.585 ;
        RECT 50.165 185.560 50.455 186.725 ;
        RECT 51.085 185.965 51.600 186.375 ;
        RECT 51.835 185.965 52.005 186.725 ;
        RECT 52.175 186.385 54.205 186.555 ;
        RECT 51.085 185.155 51.425 185.965 ;
        RECT 52.175 185.720 52.345 186.385 ;
        RECT 52.740 186.045 53.865 186.215 ;
        RECT 51.595 185.530 52.345 185.720 ;
        RECT 52.515 185.705 53.525 185.875 ;
        RECT 51.085 184.985 52.315 185.155 ;
        RECT 48.635 184.745 49.565 184.915 ;
        RECT 48.635 184.710 48.810 184.745 ;
        RECT 47.815 184.515 48.095 184.685 ;
        RECT 47.815 184.345 48.090 184.515 ;
        RECT 48.280 184.345 48.810 184.710 ;
        RECT 49.235 184.175 49.565 184.575 ;
        RECT 49.735 184.345 49.990 184.915 ;
        RECT 50.165 184.175 50.455 184.900 ;
        RECT 51.360 184.380 51.605 184.985 ;
        RECT 51.825 184.175 52.335 184.710 ;
        RECT 52.515 184.345 52.705 185.705 ;
        RECT 52.875 184.685 53.150 185.505 ;
        RECT 53.355 184.905 53.525 185.705 ;
        RECT 53.695 184.915 53.865 186.045 ;
        RECT 54.035 185.415 54.205 186.385 ;
        RECT 54.375 185.585 54.545 186.725 ;
        RECT 54.715 185.585 55.050 186.555 ;
        RECT 54.035 185.085 54.230 185.415 ;
        RECT 54.455 185.085 54.710 185.415 ;
        RECT 54.455 184.915 54.625 185.085 ;
        RECT 54.880 184.915 55.050 185.585 ;
        RECT 53.695 184.745 54.625 184.915 ;
        RECT 53.695 184.710 53.870 184.745 ;
        RECT 52.875 184.515 53.155 184.685 ;
        RECT 52.875 184.345 53.150 184.515 ;
        RECT 53.340 184.345 53.870 184.710 ;
        RECT 54.295 184.175 54.625 184.575 ;
        RECT 54.795 184.345 55.050 184.915 ;
        RECT 55.230 185.535 55.485 186.415 ;
        RECT 55.655 185.585 55.960 186.725 ;
        RECT 56.300 186.345 56.630 186.725 ;
        RECT 56.810 186.175 56.980 186.465 ;
        RECT 57.150 186.265 57.400 186.725 ;
        RECT 56.180 186.005 56.980 186.175 ;
        RECT 57.570 186.215 58.440 186.555 ;
        RECT 55.230 184.885 55.440 185.535 ;
        RECT 56.180 185.415 56.350 186.005 ;
        RECT 57.570 185.835 57.740 186.215 ;
        RECT 58.675 186.095 58.845 186.555 ;
        RECT 59.015 186.265 59.385 186.725 ;
        RECT 59.680 186.125 59.850 186.465 ;
        RECT 60.020 186.295 60.350 186.725 ;
        RECT 60.585 186.125 60.755 186.465 ;
        RECT 56.520 185.665 57.740 185.835 ;
        RECT 57.910 185.755 58.370 186.045 ;
        RECT 58.675 185.925 59.235 186.095 ;
        RECT 59.680 185.955 60.755 186.125 ;
        RECT 60.925 186.225 61.605 186.555 ;
        RECT 61.820 186.225 62.070 186.555 ;
        RECT 62.240 186.265 62.490 186.725 ;
        RECT 59.065 185.785 59.235 185.925 ;
        RECT 57.910 185.745 58.875 185.755 ;
        RECT 57.570 185.575 57.740 185.665 ;
        RECT 58.200 185.585 58.875 185.745 ;
        RECT 55.610 185.385 56.350 185.415 ;
        RECT 55.610 185.085 56.525 185.385 ;
        RECT 56.200 184.910 56.525 185.085 ;
        RECT 55.230 184.355 55.485 184.885 ;
        RECT 55.655 184.175 55.960 184.635 ;
        RECT 56.205 184.555 56.525 184.910 ;
        RECT 56.695 185.125 57.235 185.495 ;
        RECT 57.570 185.405 57.975 185.575 ;
        RECT 56.695 184.725 56.935 185.125 ;
        RECT 57.415 184.955 57.635 185.235 ;
        RECT 57.105 184.785 57.635 184.955 ;
        RECT 57.105 184.555 57.275 184.785 ;
        RECT 57.805 184.625 57.975 185.405 ;
        RECT 58.145 184.795 58.495 185.415 ;
        RECT 58.665 184.795 58.875 185.585 ;
        RECT 59.065 185.615 60.565 185.785 ;
        RECT 59.065 184.925 59.235 185.615 ;
        RECT 60.925 185.445 61.095 186.225 ;
        RECT 61.900 186.095 62.070 186.225 ;
        RECT 59.405 185.275 61.095 185.445 ;
        RECT 61.265 185.665 61.730 186.055 ;
        RECT 61.900 185.925 62.295 186.095 ;
        RECT 59.405 185.095 59.575 185.275 ;
        RECT 56.205 184.385 57.275 184.555 ;
        RECT 57.445 184.175 57.635 184.615 ;
        RECT 57.805 184.345 58.755 184.625 ;
        RECT 59.065 184.535 59.325 184.925 ;
        RECT 59.745 184.855 60.535 185.105 ;
        RECT 58.975 184.365 59.325 184.535 ;
        RECT 59.535 184.175 59.865 184.635 ;
        RECT 60.740 184.565 60.910 185.275 ;
        RECT 61.265 185.075 61.435 185.665 ;
        RECT 61.080 184.855 61.435 185.075 ;
        RECT 61.605 184.855 61.955 185.475 ;
        RECT 62.125 184.565 62.295 185.925 ;
        RECT 62.660 185.755 62.985 186.540 ;
        RECT 62.465 184.705 62.925 185.755 ;
        RECT 60.740 184.395 61.595 184.565 ;
        RECT 61.800 184.395 62.295 184.565 ;
        RECT 62.465 184.175 62.795 184.535 ;
        RECT 63.155 184.435 63.325 186.555 ;
        RECT 63.495 186.225 63.825 186.725 ;
        RECT 63.995 186.055 64.250 186.555 ;
        RECT 63.500 185.885 64.250 186.055 ;
        RECT 63.500 184.895 63.730 185.885 ;
        RECT 63.900 185.065 64.250 185.715 ;
        RECT 64.885 185.635 68.395 186.725 ;
        RECT 68.565 185.755 68.835 186.525 ;
        RECT 69.005 185.945 69.335 186.725 ;
        RECT 69.540 186.120 69.725 186.525 ;
        RECT 69.895 186.300 70.230 186.725 ;
        RECT 69.540 185.945 70.205 186.120 ;
        RECT 64.885 185.115 66.575 185.635 ;
        RECT 68.565 185.585 69.695 185.755 ;
        RECT 66.745 184.945 68.395 185.465 ;
        RECT 63.500 184.725 64.250 184.895 ;
        RECT 63.495 184.175 63.825 184.555 ;
        RECT 63.995 184.435 64.250 184.725 ;
        RECT 64.885 184.175 68.395 184.945 ;
        RECT 68.565 184.675 68.735 185.585 ;
        RECT 68.905 184.835 69.265 185.415 ;
        RECT 69.445 185.085 69.695 185.585 ;
        RECT 69.865 184.915 70.205 185.945 ;
        RECT 70.410 185.575 70.670 186.725 ;
        RECT 70.845 185.650 71.100 186.555 ;
        RECT 71.270 185.965 71.600 186.725 ;
        RECT 71.815 185.795 71.985 186.555 ;
        RECT 69.520 184.745 70.205 184.915 ;
        RECT 68.565 184.345 68.825 184.675 ;
        RECT 69.035 184.175 69.310 184.655 ;
        RECT 69.520 184.345 69.725 184.745 ;
        RECT 69.895 184.175 70.230 184.575 ;
        RECT 70.410 184.175 70.670 185.015 ;
        RECT 70.845 184.920 71.015 185.650 ;
        RECT 71.270 185.625 71.985 185.795 ;
        RECT 71.270 185.415 71.440 185.625 ;
        RECT 72.245 185.585 72.505 186.555 ;
        RECT 72.700 186.315 73.030 186.725 ;
        RECT 73.230 186.135 73.400 186.555 ;
        RECT 73.615 186.315 74.285 186.725 ;
        RECT 74.520 186.135 74.690 186.555 ;
        RECT 74.995 186.285 75.325 186.725 ;
        RECT 72.675 185.965 74.690 186.135 ;
        RECT 75.495 186.105 75.670 186.555 ;
        RECT 71.185 185.085 71.440 185.415 ;
        RECT 70.845 184.345 71.100 184.920 ;
        RECT 71.270 184.895 71.440 185.085 ;
        RECT 71.720 185.075 72.075 185.445 ;
        RECT 72.245 184.895 72.415 185.585 ;
        RECT 72.675 185.415 72.845 185.965 ;
        RECT 72.585 185.085 72.845 185.415 ;
        RECT 71.270 184.725 71.985 184.895 ;
        RECT 71.270 184.175 71.600 184.555 ;
        RECT 71.815 184.345 71.985 184.725 ;
        RECT 72.245 184.430 72.585 184.895 ;
        RECT 73.015 184.755 73.355 185.785 ;
        RECT 73.545 185.705 73.815 185.785 ;
        RECT 73.545 185.535 73.855 185.705 ;
        RECT 72.250 184.385 72.585 184.430 ;
        RECT 72.755 184.175 73.085 184.555 ;
        RECT 73.545 184.510 73.815 185.535 ;
        RECT 74.040 184.510 74.320 185.785 ;
        RECT 74.520 184.675 74.690 185.965 ;
        RECT 75.040 185.935 75.670 186.105 ;
        RECT 75.040 185.415 75.210 185.935 ;
        RECT 74.860 185.085 75.210 185.415 ;
        RECT 75.390 185.085 75.755 185.765 ;
        RECT 75.925 185.560 76.215 186.725 ;
        RECT 76.390 185.535 76.645 186.415 ;
        RECT 76.815 185.585 77.120 186.725 ;
        RECT 77.460 186.345 77.790 186.725 ;
        RECT 77.970 186.175 78.140 186.465 ;
        RECT 78.310 186.265 78.560 186.725 ;
        RECT 77.340 186.005 78.140 186.175 ;
        RECT 78.730 186.215 79.600 186.555 ;
        RECT 75.040 184.915 75.210 185.085 ;
        RECT 75.040 184.745 75.670 184.915 ;
        RECT 74.520 184.345 74.750 184.675 ;
        RECT 74.995 184.175 75.325 184.555 ;
        RECT 75.495 184.345 75.670 184.745 ;
        RECT 75.925 184.175 76.215 184.900 ;
        RECT 76.390 184.885 76.600 185.535 ;
        RECT 77.340 185.415 77.510 186.005 ;
        RECT 78.730 185.835 78.900 186.215 ;
        RECT 79.835 186.095 80.005 186.555 ;
        RECT 80.175 186.265 80.545 186.725 ;
        RECT 80.840 186.125 81.010 186.465 ;
        RECT 81.180 186.295 81.510 186.725 ;
        RECT 81.745 186.125 81.915 186.465 ;
        RECT 77.680 185.665 78.900 185.835 ;
        RECT 79.070 185.755 79.530 186.045 ;
        RECT 79.835 185.925 80.395 186.095 ;
        RECT 80.840 185.955 81.915 186.125 ;
        RECT 82.085 186.225 82.765 186.555 ;
        RECT 82.980 186.225 83.230 186.555 ;
        RECT 83.400 186.265 83.650 186.725 ;
        RECT 80.225 185.785 80.395 185.925 ;
        RECT 79.070 185.745 80.035 185.755 ;
        RECT 78.730 185.575 78.900 185.665 ;
        RECT 79.360 185.585 80.035 185.745 ;
        RECT 76.770 185.385 77.510 185.415 ;
        RECT 76.770 185.085 77.685 185.385 ;
        RECT 77.360 184.910 77.685 185.085 ;
        RECT 76.390 184.355 76.645 184.885 ;
        RECT 76.815 184.175 77.120 184.635 ;
        RECT 77.365 184.555 77.685 184.910 ;
        RECT 77.855 185.125 78.395 185.495 ;
        RECT 78.730 185.405 79.135 185.575 ;
        RECT 77.855 184.725 78.095 185.125 ;
        RECT 78.575 184.955 78.795 185.235 ;
        RECT 78.265 184.785 78.795 184.955 ;
        RECT 78.265 184.555 78.435 184.785 ;
        RECT 78.965 184.625 79.135 185.405 ;
        RECT 79.305 184.795 79.655 185.415 ;
        RECT 79.825 184.795 80.035 185.585 ;
        RECT 80.225 185.615 81.725 185.785 ;
        RECT 80.225 184.925 80.395 185.615 ;
        RECT 82.085 185.445 82.255 186.225 ;
        RECT 83.060 186.095 83.230 186.225 ;
        RECT 80.565 185.275 82.255 185.445 ;
        RECT 82.425 185.665 82.890 186.055 ;
        RECT 83.060 185.925 83.455 186.095 ;
        RECT 80.565 185.095 80.735 185.275 ;
        RECT 77.365 184.385 78.435 184.555 ;
        RECT 78.605 184.175 78.795 184.615 ;
        RECT 78.965 184.345 79.915 184.625 ;
        RECT 80.225 184.535 80.485 184.925 ;
        RECT 80.905 184.855 81.695 185.105 ;
        RECT 80.135 184.365 80.485 184.535 ;
        RECT 80.695 184.175 81.025 184.635 ;
        RECT 81.900 184.565 82.070 185.275 ;
        RECT 82.425 185.075 82.595 185.665 ;
        RECT 82.240 184.855 82.595 185.075 ;
        RECT 82.765 184.855 83.115 185.475 ;
        RECT 83.285 184.565 83.455 185.925 ;
        RECT 83.820 185.755 84.145 186.540 ;
        RECT 83.625 184.705 84.085 185.755 ;
        RECT 81.900 184.395 82.755 184.565 ;
        RECT 82.960 184.395 83.455 184.565 ;
        RECT 83.625 184.175 83.955 184.535 ;
        RECT 84.315 184.435 84.485 186.555 ;
        RECT 84.655 186.225 84.985 186.725 ;
        RECT 85.155 186.055 85.410 186.555 ;
        RECT 84.660 185.885 85.410 186.055 ;
        RECT 84.660 184.895 84.890 185.885 ;
        RECT 85.060 185.065 85.410 185.715 ;
        RECT 85.585 185.635 87.255 186.725 ;
        RECT 85.585 185.115 86.335 185.635 ;
        RECT 87.430 185.535 87.685 186.415 ;
        RECT 87.855 185.585 88.160 186.725 ;
        RECT 88.500 186.345 88.830 186.725 ;
        RECT 89.010 186.175 89.180 186.465 ;
        RECT 89.350 186.265 89.600 186.725 ;
        RECT 88.380 186.005 89.180 186.175 ;
        RECT 89.770 186.215 90.640 186.555 ;
        RECT 86.505 184.945 87.255 185.465 ;
        RECT 84.660 184.725 85.410 184.895 ;
        RECT 84.655 184.175 84.985 184.555 ;
        RECT 85.155 184.435 85.410 184.725 ;
        RECT 85.585 184.175 87.255 184.945 ;
        RECT 87.430 184.885 87.640 185.535 ;
        RECT 88.380 185.415 88.550 186.005 ;
        RECT 89.770 185.835 89.940 186.215 ;
        RECT 90.875 186.095 91.045 186.555 ;
        RECT 91.215 186.265 91.585 186.725 ;
        RECT 91.880 186.125 92.050 186.465 ;
        RECT 92.220 186.295 92.550 186.725 ;
        RECT 92.785 186.125 92.955 186.465 ;
        RECT 88.720 185.665 89.940 185.835 ;
        RECT 90.110 185.755 90.570 186.045 ;
        RECT 90.875 185.925 91.435 186.095 ;
        RECT 91.880 185.955 92.955 186.125 ;
        RECT 93.125 186.225 93.805 186.555 ;
        RECT 94.020 186.225 94.270 186.555 ;
        RECT 94.440 186.265 94.690 186.725 ;
        RECT 91.265 185.785 91.435 185.925 ;
        RECT 90.110 185.745 91.075 185.755 ;
        RECT 89.770 185.575 89.940 185.665 ;
        RECT 90.400 185.585 91.075 185.745 ;
        RECT 87.810 185.385 88.550 185.415 ;
        RECT 87.810 185.085 88.725 185.385 ;
        RECT 88.400 184.910 88.725 185.085 ;
        RECT 87.430 184.355 87.685 184.885 ;
        RECT 87.855 184.175 88.160 184.635 ;
        RECT 88.405 184.555 88.725 184.910 ;
        RECT 88.895 185.125 89.435 185.495 ;
        RECT 89.770 185.405 90.175 185.575 ;
        RECT 88.895 184.725 89.135 185.125 ;
        RECT 89.615 184.955 89.835 185.235 ;
        RECT 89.305 184.785 89.835 184.955 ;
        RECT 89.305 184.555 89.475 184.785 ;
        RECT 90.005 184.625 90.175 185.405 ;
        RECT 90.345 184.795 90.695 185.415 ;
        RECT 90.865 184.795 91.075 185.585 ;
        RECT 91.265 185.615 92.765 185.785 ;
        RECT 91.265 184.925 91.435 185.615 ;
        RECT 93.125 185.445 93.295 186.225 ;
        RECT 94.100 186.095 94.270 186.225 ;
        RECT 91.605 185.275 93.295 185.445 ;
        RECT 93.465 185.665 93.930 186.055 ;
        RECT 94.100 185.925 94.495 186.095 ;
        RECT 91.605 185.095 91.775 185.275 ;
        RECT 88.405 184.385 89.475 184.555 ;
        RECT 89.645 184.175 89.835 184.615 ;
        RECT 90.005 184.345 90.955 184.625 ;
        RECT 91.265 184.535 91.525 184.925 ;
        RECT 91.945 184.855 92.735 185.105 ;
        RECT 91.175 184.365 91.525 184.535 ;
        RECT 91.735 184.175 92.065 184.635 ;
        RECT 92.940 184.565 93.110 185.275 ;
        RECT 93.465 185.075 93.635 185.665 ;
        RECT 93.280 184.855 93.635 185.075 ;
        RECT 93.805 184.855 94.155 185.475 ;
        RECT 94.325 184.565 94.495 185.925 ;
        RECT 94.860 185.755 95.185 186.540 ;
        RECT 94.665 184.705 95.125 185.755 ;
        RECT 92.940 184.395 93.795 184.565 ;
        RECT 94.000 184.395 94.495 184.565 ;
        RECT 94.665 184.175 94.995 184.535 ;
        RECT 95.355 184.435 95.525 186.555 ;
        RECT 95.695 186.225 96.025 186.725 ;
        RECT 96.195 186.055 96.450 186.555 ;
        RECT 95.700 185.885 96.450 186.055 ;
        RECT 97.085 185.965 97.600 186.375 ;
        RECT 97.835 185.965 98.005 186.725 ;
        RECT 98.175 186.385 100.205 186.555 ;
        RECT 95.700 184.895 95.930 185.885 ;
        RECT 96.100 185.065 96.450 185.715 ;
        RECT 97.085 185.155 97.425 185.965 ;
        RECT 98.175 185.720 98.345 186.385 ;
        RECT 98.740 186.045 99.865 186.215 ;
        RECT 97.595 185.530 98.345 185.720 ;
        RECT 98.515 185.705 99.525 185.875 ;
        RECT 97.085 184.985 98.315 185.155 ;
        RECT 95.700 184.725 96.450 184.895 ;
        RECT 95.695 184.175 96.025 184.555 ;
        RECT 96.195 184.435 96.450 184.725 ;
        RECT 97.360 184.380 97.605 184.985 ;
        RECT 97.825 184.175 98.335 184.710 ;
        RECT 98.515 184.345 98.705 185.705 ;
        RECT 98.875 184.685 99.150 185.505 ;
        RECT 99.355 184.905 99.525 185.705 ;
        RECT 99.695 184.915 99.865 186.045 ;
        RECT 100.035 185.415 100.205 186.385 ;
        RECT 100.375 185.585 100.545 186.725 ;
        RECT 100.715 185.585 101.050 186.555 ;
        RECT 100.035 185.085 100.230 185.415 ;
        RECT 100.455 185.085 100.710 185.415 ;
        RECT 100.455 184.915 100.625 185.085 ;
        RECT 100.880 184.915 101.050 185.585 ;
        RECT 101.685 185.560 101.975 186.725 ;
        RECT 102.145 185.635 103.815 186.725 ;
        RECT 103.985 185.965 104.500 186.375 ;
        RECT 104.735 185.965 104.905 186.725 ;
        RECT 105.075 186.385 107.105 186.555 ;
        RECT 102.145 185.115 102.895 185.635 ;
        RECT 103.065 184.945 103.815 185.465 ;
        RECT 103.985 185.155 104.325 185.965 ;
        RECT 105.075 185.720 105.245 186.385 ;
        RECT 105.640 186.045 106.765 186.215 ;
        RECT 104.495 185.530 105.245 185.720 ;
        RECT 105.415 185.705 106.425 185.875 ;
        RECT 103.985 184.985 105.215 185.155 ;
        RECT 99.695 184.745 100.625 184.915 ;
        RECT 99.695 184.710 99.870 184.745 ;
        RECT 98.875 184.515 99.155 184.685 ;
        RECT 98.875 184.345 99.150 184.515 ;
        RECT 99.340 184.345 99.870 184.710 ;
        RECT 100.295 184.175 100.625 184.575 ;
        RECT 100.795 184.345 101.050 184.915 ;
        RECT 101.685 184.175 101.975 184.900 ;
        RECT 102.145 184.175 103.815 184.945 ;
        RECT 104.260 184.380 104.505 184.985 ;
        RECT 104.725 184.175 105.235 184.710 ;
        RECT 105.415 184.345 105.605 185.705 ;
        RECT 105.775 185.365 106.050 185.505 ;
        RECT 105.775 185.195 106.055 185.365 ;
        RECT 105.775 184.345 106.050 185.195 ;
        RECT 106.255 184.905 106.425 185.705 ;
        RECT 106.595 184.915 106.765 186.045 ;
        RECT 106.935 185.415 107.105 186.385 ;
        RECT 107.275 185.585 107.445 186.725 ;
        RECT 107.615 185.585 107.950 186.555 ;
        RECT 106.935 185.085 107.130 185.415 ;
        RECT 107.355 185.085 107.610 185.415 ;
        RECT 107.355 184.915 107.525 185.085 ;
        RECT 107.780 184.915 107.950 185.585 ;
        RECT 108.585 185.635 111.175 186.725 ;
        RECT 111.345 185.965 111.860 186.375 ;
        RECT 112.095 185.965 112.265 186.725 ;
        RECT 112.435 186.385 114.465 186.555 ;
        RECT 108.585 185.115 109.795 185.635 ;
        RECT 109.965 184.945 111.175 185.465 ;
        RECT 111.345 185.155 111.685 185.965 ;
        RECT 112.435 185.720 112.605 186.385 ;
        RECT 113.000 186.045 114.125 186.215 ;
        RECT 111.855 185.530 112.605 185.720 ;
        RECT 112.775 185.705 113.785 185.875 ;
        RECT 111.345 184.985 112.575 185.155 ;
        RECT 106.595 184.745 107.525 184.915 ;
        RECT 106.595 184.710 106.770 184.745 ;
        RECT 106.240 184.345 106.770 184.710 ;
        RECT 107.195 184.175 107.525 184.575 ;
        RECT 107.695 184.345 107.950 184.915 ;
        RECT 108.585 184.175 111.175 184.945 ;
        RECT 111.620 184.380 111.865 184.985 ;
        RECT 112.085 184.175 112.595 184.710 ;
        RECT 112.775 184.345 112.965 185.705 ;
        RECT 113.135 184.685 113.410 185.505 ;
        RECT 113.615 184.905 113.785 185.705 ;
        RECT 113.955 184.915 114.125 186.045 ;
        RECT 114.295 185.415 114.465 186.385 ;
        RECT 114.635 185.585 114.805 186.725 ;
        RECT 114.975 185.585 115.310 186.555 ;
        RECT 114.295 185.085 114.490 185.415 ;
        RECT 114.715 185.085 114.970 185.415 ;
        RECT 114.715 184.915 114.885 185.085 ;
        RECT 115.140 184.915 115.310 185.585 ;
        RECT 115.485 185.965 116.000 186.375 ;
        RECT 116.235 185.965 116.405 186.725 ;
        RECT 116.575 186.385 118.605 186.555 ;
        RECT 115.485 185.155 115.825 185.965 ;
        RECT 116.575 185.720 116.745 186.385 ;
        RECT 117.140 186.045 118.265 186.215 ;
        RECT 115.995 185.530 116.745 185.720 ;
        RECT 116.915 185.705 117.925 185.875 ;
        RECT 115.485 184.985 116.715 185.155 ;
        RECT 113.955 184.745 114.885 184.915 ;
        RECT 113.955 184.710 114.130 184.745 ;
        RECT 113.135 184.515 113.415 184.685 ;
        RECT 113.135 184.345 113.410 184.515 ;
        RECT 113.600 184.345 114.130 184.710 ;
        RECT 114.555 184.175 114.885 184.575 ;
        RECT 115.055 184.345 115.310 184.915 ;
        RECT 115.760 184.380 116.005 184.985 ;
        RECT 116.225 184.175 116.735 184.710 ;
        RECT 116.915 184.345 117.105 185.705 ;
        RECT 117.275 185.365 117.550 185.505 ;
        RECT 117.275 185.195 117.555 185.365 ;
        RECT 117.275 184.345 117.550 185.195 ;
        RECT 117.755 184.905 117.925 185.705 ;
        RECT 118.095 184.915 118.265 186.045 ;
        RECT 118.435 185.415 118.605 186.385 ;
        RECT 118.775 185.585 118.945 186.725 ;
        RECT 119.115 185.585 119.450 186.555 ;
        RECT 118.435 185.085 118.630 185.415 ;
        RECT 118.855 185.085 119.110 185.415 ;
        RECT 118.855 184.915 119.025 185.085 ;
        RECT 119.280 184.915 119.450 185.585 ;
        RECT 119.625 185.635 120.835 186.725 ;
        RECT 121.010 186.290 126.355 186.725 ;
        RECT 119.625 185.095 120.145 185.635 ;
        RECT 120.315 184.925 120.835 185.465 ;
        RECT 122.600 185.040 122.950 186.290 ;
        RECT 126.525 185.635 127.735 186.725 ;
        RECT 118.095 184.745 119.025 184.915 ;
        RECT 118.095 184.710 118.270 184.745 ;
        RECT 117.740 184.345 118.270 184.710 ;
        RECT 118.695 184.175 119.025 184.575 ;
        RECT 119.195 184.345 119.450 184.915 ;
        RECT 119.625 184.175 120.835 184.925 ;
        RECT 124.430 184.720 124.770 185.550 ;
        RECT 126.525 185.095 127.045 185.635 ;
        RECT 127.215 184.925 127.735 185.465 ;
        RECT 121.010 184.175 126.355 184.720 ;
        RECT 126.525 184.175 127.735 184.925 ;
        RECT 20.640 184.005 127.820 184.175 ;
        RECT 20.725 183.255 21.935 184.005 ;
        RECT 22.570 183.460 27.915 184.005 ;
        RECT 20.725 182.715 21.245 183.255 ;
        RECT 21.415 182.545 21.935 183.085 ;
        RECT 20.725 181.455 21.935 182.545 ;
        RECT 24.160 181.890 24.510 183.140 ;
        RECT 25.990 182.630 26.330 183.460 ;
        RECT 28.090 183.455 28.345 183.745 ;
        RECT 28.515 183.625 28.845 184.005 ;
        RECT 28.090 183.285 28.840 183.455 ;
        RECT 28.090 182.465 28.440 183.115 ;
        RECT 28.610 182.295 28.840 183.285 ;
        RECT 28.090 182.125 28.840 182.295 ;
        RECT 22.570 181.455 27.915 181.890 ;
        RECT 28.090 181.625 28.345 182.125 ;
        RECT 28.515 181.455 28.845 181.955 ;
        RECT 29.015 181.625 29.185 183.745 ;
        RECT 29.545 183.645 29.875 184.005 ;
        RECT 30.045 183.615 30.540 183.785 ;
        RECT 30.745 183.615 31.600 183.785 ;
        RECT 29.415 182.425 29.875 183.475 ;
        RECT 29.355 181.640 29.680 182.425 ;
        RECT 30.045 182.255 30.215 183.615 ;
        RECT 30.385 182.705 30.735 183.325 ;
        RECT 30.905 183.105 31.260 183.325 ;
        RECT 30.905 182.515 31.075 183.105 ;
        RECT 31.430 182.905 31.600 183.615 ;
        RECT 32.475 183.545 32.805 184.005 ;
        RECT 33.015 183.645 33.365 183.815 ;
        RECT 31.805 183.075 32.595 183.325 ;
        RECT 33.015 183.255 33.275 183.645 ;
        RECT 33.585 183.555 34.535 183.835 ;
        RECT 34.705 183.565 34.895 184.005 ;
        RECT 35.065 183.625 36.135 183.795 ;
        RECT 32.765 182.905 32.935 183.085 ;
        RECT 30.045 182.085 30.440 182.255 ;
        RECT 30.610 182.125 31.075 182.515 ;
        RECT 31.245 182.735 32.935 182.905 ;
        RECT 30.270 181.955 30.440 182.085 ;
        RECT 31.245 181.955 31.415 182.735 ;
        RECT 33.105 182.565 33.275 183.255 ;
        RECT 31.775 182.395 33.275 182.565 ;
        RECT 33.465 182.595 33.675 183.385 ;
        RECT 33.845 182.765 34.195 183.385 ;
        RECT 34.365 182.775 34.535 183.555 ;
        RECT 35.065 183.395 35.235 183.625 ;
        RECT 34.705 183.225 35.235 183.395 ;
        RECT 34.705 182.945 34.925 183.225 ;
        RECT 35.405 183.055 35.645 183.455 ;
        RECT 34.365 182.605 34.770 182.775 ;
        RECT 35.105 182.685 35.645 183.055 ;
        RECT 35.815 183.270 36.135 183.625 ;
        RECT 36.380 183.545 36.685 184.005 ;
        RECT 36.855 183.295 37.110 183.825 ;
        RECT 35.815 183.095 36.140 183.270 ;
        RECT 35.815 182.795 36.730 183.095 ;
        RECT 35.990 182.765 36.730 182.795 ;
        RECT 33.465 182.435 34.140 182.595 ;
        RECT 34.600 182.515 34.770 182.605 ;
        RECT 33.465 182.425 34.430 182.435 ;
        RECT 33.105 182.255 33.275 182.395 ;
        RECT 29.850 181.455 30.100 181.915 ;
        RECT 30.270 181.625 30.520 181.955 ;
        RECT 30.735 181.625 31.415 181.955 ;
        RECT 31.585 182.055 32.660 182.225 ;
        RECT 33.105 182.085 33.665 182.255 ;
        RECT 33.970 182.135 34.430 182.425 ;
        RECT 34.600 182.345 35.820 182.515 ;
        RECT 31.585 181.715 31.755 182.055 ;
        RECT 31.990 181.455 32.320 181.885 ;
        RECT 32.490 181.715 32.660 182.055 ;
        RECT 32.955 181.455 33.325 181.915 ;
        RECT 33.495 181.625 33.665 182.085 ;
        RECT 34.600 181.965 34.770 182.345 ;
        RECT 35.990 182.175 36.160 182.765 ;
        RECT 36.900 182.645 37.110 183.295 ;
        RECT 37.285 183.280 37.575 184.005 ;
        RECT 37.745 183.235 40.335 184.005 ;
        RECT 33.900 181.625 34.770 181.965 ;
        RECT 35.360 182.005 36.160 182.175 ;
        RECT 34.940 181.455 35.190 181.915 ;
        RECT 35.360 181.715 35.530 182.005 ;
        RECT 35.710 181.455 36.040 181.835 ;
        RECT 36.380 181.455 36.685 182.595 ;
        RECT 36.855 181.765 37.110 182.645 ;
        RECT 37.285 181.455 37.575 182.620 ;
        RECT 37.745 182.545 38.955 183.065 ;
        RECT 39.125 182.715 40.335 183.235 ;
        RECT 40.510 183.295 40.765 183.825 ;
        RECT 40.935 183.545 41.240 184.005 ;
        RECT 41.485 183.625 42.555 183.795 ;
        RECT 40.510 182.645 40.720 183.295 ;
        RECT 41.485 183.270 41.805 183.625 ;
        RECT 41.480 183.095 41.805 183.270 ;
        RECT 40.890 182.795 41.805 183.095 ;
        RECT 41.975 183.055 42.215 183.455 ;
        RECT 42.385 183.395 42.555 183.625 ;
        RECT 42.725 183.565 42.915 184.005 ;
        RECT 43.085 183.555 44.035 183.835 ;
        RECT 44.255 183.645 44.605 183.815 ;
        RECT 42.385 183.225 42.915 183.395 ;
        RECT 40.890 182.765 41.630 182.795 ;
        RECT 37.745 181.455 40.335 182.545 ;
        RECT 40.510 181.765 40.765 182.645 ;
        RECT 40.935 181.455 41.240 182.595 ;
        RECT 41.460 182.175 41.630 182.765 ;
        RECT 41.975 182.685 42.515 183.055 ;
        RECT 42.695 182.945 42.915 183.225 ;
        RECT 43.085 182.775 43.255 183.555 ;
        RECT 42.850 182.605 43.255 182.775 ;
        RECT 43.425 182.765 43.775 183.385 ;
        RECT 42.850 182.515 43.020 182.605 ;
        RECT 43.945 182.595 44.155 183.385 ;
        RECT 41.800 182.345 43.020 182.515 ;
        RECT 43.480 182.435 44.155 182.595 ;
        RECT 41.460 182.005 42.260 182.175 ;
        RECT 41.580 181.455 41.910 181.835 ;
        RECT 42.090 181.715 42.260 182.005 ;
        RECT 42.850 181.965 43.020 182.345 ;
        RECT 43.190 182.425 44.155 182.435 ;
        RECT 44.345 183.255 44.605 183.645 ;
        RECT 44.815 183.545 45.145 184.005 ;
        RECT 46.020 183.615 46.875 183.785 ;
        RECT 47.080 183.615 47.575 183.785 ;
        RECT 47.745 183.645 48.075 184.005 ;
        RECT 44.345 182.565 44.515 183.255 ;
        RECT 44.685 182.905 44.855 183.085 ;
        RECT 45.025 183.075 45.815 183.325 ;
        RECT 46.020 182.905 46.190 183.615 ;
        RECT 46.360 183.105 46.715 183.325 ;
        RECT 44.685 182.735 46.375 182.905 ;
        RECT 43.190 182.135 43.650 182.425 ;
        RECT 44.345 182.395 45.845 182.565 ;
        RECT 44.345 182.255 44.515 182.395 ;
        RECT 43.955 182.085 44.515 182.255 ;
        RECT 42.430 181.455 42.680 181.915 ;
        RECT 42.850 181.625 43.720 181.965 ;
        RECT 43.955 181.625 44.125 182.085 ;
        RECT 44.960 182.055 46.035 182.225 ;
        RECT 44.295 181.455 44.665 181.915 ;
        RECT 44.960 181.715 45.130 182.055 ;
        RECT 45.300 181.455 45.630 181.885 ;
        RECT 45.865 181.715 46.035 182.055 ;
        RECT 46.205 181.955 46.375 182.735 ;
        RECT 46.545 182.515 46.715 183.105 ;
        RECT 46.885 182.705 47.235 183.325 ;
        RECT 46.545 182.125 47.010 182.515 ;
        RECT 47.405 182.255 47.575 183.615 ;
        RECT 47.745 182.425 48.205 183.475 ;
        RECT 47.180 182.085 47.575 182.255 ;
        RECT 47.180 181.955 47.350 182.085 ;
        RECT 46.205 181.625 46.885 181.955 ;
        RECT 47.100 181.625 47.350 181.955 ;
        RECT 47.520 181.455 47.770 181.915 ;
        RECT 47.940 181.640 48.265 182.425 ;
        RECT 48.435 181.625 48.605 183.745 ;
        RECT 48.775 183.625 49.105 184.005 ;
        RECT 49.275 183.455 49.530 183.745 ;
        RECT 48.780 183.285 49.530 183.455 ;
        RECT 49.705 183.330 49.965 183.835 ;
        RECT 50.145 183.625 50.475 184.005 ;
        RECT 50.655 183.455 50.825 183.835 ;
        RECT 48.780 182.295 49.010 183.285 ;
        RECT 49.180 182.465 49.530 183.115 ;
        RECT 49.705 182.530 49.875 183.330 ;
        RECT 50.160 183.285 50.825 183.455 ;
        RECT 50.160 183.030 50.330 183.285 ;
        RECT 51.545 183.235 55.055 184.005 ;
        RECT 55.230 183.460 60.575 184.005 ;
        RECT 50.045 182.700 50.330 183.030 ;
        RECT 50.565 182.735 50.895 183.105 ;
        RECT 50.160 182.555 50.330 182.700 ;
        RECT 48.780 182.125 49.530 182.295 ;
        RECT 48.775 181.455 49.105 181.955 ;
        RECT 49.275 181.625 49.530 182.125 ;
        RECT 49.705 181.625 49.975 182.530 ;
        RECT 50.160 182.385 50.825 182.555 ;
        RECT 50.145 181.455 50.475 182.215 ;
        RECT 50.655 181.625 50.825 182.385 ;
        RECT 51.545 182.545 53.235 183.065 ;
        RECT 53.405 182.715 55.055 183.235 ;
        RECT 51.545 181.455 55.055 182.545 ;
        RECT 56.820 181.890 57.170 183.140 ;
        RECT 58.650 182.630 58.990 183.460 ;
        RECT 60.835 183.455 61.005 183.835 ;
        RECT 61.185 183.625 61.515 184.005 ;
        RECT 60.835 183.285 61.500 183.455 ;
        RECT 61.695 183.330 61.955 183.835 ;
        RECT 60.765 182.735 61.095 183.105 ;
        RECT 61.330 183.030 61.500 183.285 ;
        RECT 61.330 182.700 61.615 183.030 ;
        RECT 61.330 182.555 61.500 182.700 ;
        RECT 60.835 182.385 61.500 182.555 ;
        RECT 61.785 182.530 61.955 183.330 ;
        RECT 63.045 183.280 63.335 184.005 ;
        RECT 63.505 183.235 66.095 184.005 ;
        RECT 66.270 183.460 71.615 184.005 ;
        RECT 55.230 181.455 60.575 181.890 ;
        RECT 60.835 181.625 61.005 182.385 ;
        RECT 61.185 181.455 61.515 182.215 ;
        RECT 61.685 181.625 61.955 182.530 ;
        RECT 63.045 181.455 63.335 182.620 ;
        RECT 63.505 182.545 64.715 183.065 ;
        RECT 64.885 182.715 66.095 183.235 ;
        RECT 63.505 181.455 66.095 182.545 ;
        RECT 67.860 181.890 68.210 183.140 ;
        RECT 69.690 182.630 70.030 183.460 ;
        RECT 66.270 181.455 71.615 181.890 ;
        RECT 71.785 181.625 72.045 183.835 ;
        RECT 72.215 183.625 72.545 184.005 ;
        RECT 72.755 183.095 72.950 183.670 ;
        RECT 73.220 183.095 73.405 183.675 ;
        RECT 72.215 182.175 72.385 183.095 ;
        RECT 72.695 182.765 72.950 183.095 ;
        RECT 73.175 182.765 73.405 183.095 ;
        RECT 73.655 183.665 75.135 183.835 ;
        RECT 73.655 182.765 73.825 183.665 ;
        RECT 73.995 183.165 74.545 183.495 ;
        RECT 74.735 183.335 75.135 183.665 ;
        RECT 75.315 183.625 75.645 184.005 ;
        RECT 75.955 183.505 76.215 183.835 ;
        RECT 72.755 182.455 72.950 182.765 ;
        RECT 73.220 182.455 73.405 182.765 ;
        RECT 73.995 182.175 74.165 183.165 ;
        RECT 74.735 182.855 74.905 183.335 ;
        RECT 75.485 183.145 75.695 183.325 ;
        RECT 75.075 182.975 75.695 183.145 ;
        RECT 72.215 182.005 74.165 182.175 ;
        RECT 74.335 182.685 74.905 182.855 ;
        RECT 76.045 182.805 76.215 183.505 ;
        RECT 76.885 183.185 77.115 184.005 ;
        RECT 77.285 183.205 77.615 183.835 ;
        RECT 74.335 182.175 74.505 182.685 ;
        RECT 75.085 182.635 76.215 182.805 ;
        RECT 76.865 182.765 77.195 183.015 ;
        RECT 75.085 182.515 75.255 182.635 ;
        RECT 74.675 182.345 75.255 182.515 ;
        RECT 74.335 182.005 75.075 182.175 ;
        RECT 75.525 182.135 75.875 182.465 ;
        RECT 72.215 181.455 72.545 181.835 ;
        RECT 72.970 181.625 73.140 182.005 ;
        RECT 73.400 181.455 73.730 181.835 ;
        RECT 73.925 181.625 74.095 182.005 ;
        RECT 74.305 181.455 74.635 181.835 ;
        RECT 74.885 181.625 75.075 182.005 ;
        RECT 76.045 181.955 76.215 182.635 ;
        RECT 77.365 182.605 77.615 183.205 ;
        RECT 77.785 183.185 77.995 184.005 ;
        RECT 79.185 183.185 79.415 184.005 ;
        RECT 79.585 183.205 79.915 183.835 ;
        RECT 79.165 182.765 79.495 183.015 ;
        RECT 79.665 182.605 79.915 183.205 ;
        RECT 80.085 183.185 80.295 184.005 ;
        RECT 80.525 183.235 84.035 184.005 ;
        RECT 75.315 181.455 75.645 181.835 ;
        RECT 75.955 181.625 76.215 181.955 ;
        RECT 76.885 181.455 77.115 182.595 ;
        RECT 77.285 181.625 77.615 182.605 ;
        RECT 77.785 181.455 77.995 182.595 ;
        RECT 79.185 181.455 79.415 182.595 ;
        RECT 79.585 181.625 79.915 182.605 ;
        RECT 80.085 181.455 80.295 182.595 ;
        RECT 80.525 182.545 82.215 183.065 ;
        RECT 82.385 182.715 84.035 183.235 ;
        RECT 84.295 183.355 84.465 183.835 ;
        RECT 84.645 183.525 84.885 184.005 ;
        RECT 85.135 183.355 85.305 183.835 ;
        RECT 85.475 183.525 85.805 184.005 ;
        RECT 85.975 183.355 86.145 183.835 ;
        RECT 84.295 183.185 84.930 183.355 ;
        RECT 85.135 183.185 86.145 183.355 ;
        RECT 86.315 183.205 86.645 184.005 ;
        RECT 86.965 183.235 88.635 184.005 ;
        RECT 88.805 183.280 89.095 184.005 ;
        RECT 84.760 183.015 84.930 183.185 ;
        RECT 85.645 183.155 86.145 183.185 ;
        RECT 84.210 182.775 84.590 183.015 ;
        RECT 84.760 182.845 85.260 183.015 ;
        RECT 84.760 182.605 84.930 182.845 ;
        RECT 85.650 182.645 86.145 183.155 ;
        RECT 80.525 181.455 84.035 182.545 ;
        RECT 84.215 182.435 84.930 182.605 ;
        RECT 85.135 182.475 86.145 182.645 ;
        RECT 84.215 181.625 84.545 182.435 ;
        RECT 84.715 181.455 84.955 182.255 ;
        RECT 85.135 181.625 85.305 182.475 ;
        RECT 85.475 181.455 85.805 182.255 ;
        RECT 85.975 181.625 86.145 182.475 ;
        RECT 86.315 181.455 86.645 182.605 ;
        RECT 86.965 182.545 87.715 183.065 ;
        RECT 87.885 182.715 88.635 183.235 ;
        RECT 90.000 183.195 90.245 183.800 ;
        RECT 90.465 183.470 90.975 184.005 ;
        RECT 89.725 183.025 90.955 183.195 ;
        RECT 86.965 181.455 88.635 182.545 ;
        RECT 88.805 181.455 89.095 182.620 ;
        RECT 89.725 182.215 90.065 183.025 ;
        RECT 90.235 182.460 90.985 182.650 ;
        RECT 89.725 181.805 90.240 182.215 ;
        RECT 90.475 181.455 90.645 182.215 ;
        RECT 90.815 181.795 90.985 182.460 ;
        RECT 91.155 182.475 91.345 183.835 ;
        RECT 91.515 183.665 91.790 183.835 ;
        RECT 91.515 183.495 91.795 183.665 ;
        RECT 91.515 182.675 91.790 183.495 ;
        RECT 91.980 183.470 92.510 183.835 ;
        RECT 92.935 183.605 93.265 184.005 ;
        RECT 92.335 183.435 92.510 183.470 ;
        RECT 91.995 182.475 92.165 183.275 ;
        RECT 91.155 182.305 92.165 182.475 ;
        RECT 92.335 183.265 93.265 183.435 ;
        RECT 93.435 183.265 93.690 183.835 ;
        RECT 92.335 182.135 92.505 183.265 ;
        RECT 93.095 183.095 93.265 183.265 ;
        RECT 91.380 181.965 92.505 182.135 ;
        RECT 92.675 182.765 92.870 183.095 ;
        RECT 93.095 182.765 93.350 183.095 ;
        RECT 92.675 181.795 92.845 182.765 ;
        RECT 93.520 182.595 93.690 183.265 ;
        RECT 90.815 181.625 92.845 181.795 ;
        RECT 93.015 181.455 93.185 182.595 ;
        RECT 93.355 181.625 93.690 182.595 ;
        RECT 93.870 183.295 94.125 183.825 ;
        RECT 94.295 183.545 94.600 184.005 ;
        RECT 94.845 183.625 95.915 183.795 ;
        RECT 93.870 182.645 94.080 183.295 ;
        RECT 94.845 183.270 95.165 183.625 ;
        RECT 94.840 183.095 95.165 183.270 ;
        RECT 94.250 182.795 95.165 183.095 ;
        RECT 95.335 183.055 95.575 183.455 ;
        RECT 95.745 183.395 95.915 183.625 ;
        RECT 96.085 183.565 96.275 184.005 ;
        RECT 96.445 183.555 97.395 183.835 ;
        RECT 97.615 183.645 97.965 183.815 ;
        RECT 95.745 183.225 96.275 183.395 ;
        RECT 94.250 182.765 94.990 182.795 ;
        RECT 93.870 181.765 94.125 182.645 ;
        RECT 94.295 181.455 94.600 182.595 ;
        RECT 94.820 182.175 94.990 182.765 ;
        RECT 95.335 182.685 95.875 183.055 ;
        RECT 96.055 182.945 96.275 183.225 ;
        RECT 96.445 182.775 96.615 183.555 ;
        RECT 96.210 182.605 96.615 182.775 ;
        RECT 96.785 182.765 97.135 183.385 ;
        RECT 96.210 182.515 96.380 182.605 ;
        RECT 97.305 182.595 97.515 183.385 ;
        RECT 95.160 182.345 96.380 182.515 ;
        RECT 96.840 182.435 97.515 182.595 ;
        RECT 94.820 182.005 95.620 182.175 ;
        RECT 94.940 181.455 95.270 181.835 ;
        RECT 95.450 181.715 95.620 182.005 ;
        RECT 96.210 181.965 96.380 182.345 ;
        RECT 96.550 182.425 97.515 182.435 ;
        RECT 97.705 183.255 97.965 183.645 ;
        RECT 98.175 183.545 98.505 184.005 ;
        RECT 99.380 183.615 100.235 183.785 ;
        RECT 100.440 183.615 100.935 183.785 ;
        RECT 101.105 183.645 101.435 184.005 ;
        RECT 97.705 182.565 97.875 183.255 ;
        RECT 98.045 182.905 98.215 183.085 ;
        RECT 98.385 183.075 99.175 183.325 ;
        RECT 99.380 182.905 99.550 183.615 ;
        RECT 99.720 183.105 100.075 183.325 ;
        RECT 98.045 182.735 99.735 182.905 ;
        RECT 96.550 182.135 97.010 182.425 ;
        RECT 97.705 182.395 99.205 182.565 ;
        RECT 97.705 182.255 97.875 182.395 ;
        RECT 97.315 182.085 97.875 182.255 ;
        RECT 95.790 181.455 96.040 181.915 ;
        RECT 96.210 181.625 97.080 181.965 ;
        RECT 97.315 181.625 97.485 182.085 ;
        RECT 98.320 182.055 99.395 182.225 ;
        RECT 97.655 181.455 98.025 181.915 ;
        RECT 98.320 181.715 98.490 182.055 ;
        RECT 98.660 181.455 98.990 181.885 ;
        RECT 99.225 181.715 99.395 182.055 ;
        RECT 99.565 181.955 99.735 182.735 ;
        RECT 99.905 182.515 100.075 183.105 ;
        RECT 100.245 182.705 100.595 183.325 ;
        RECT 99.905 182.125 100.370 182.515 ;
        RECT 100.765 182.255 100.935 183.615 ;
        RECT 101.105 182.425 101.565 183.475 ;
        RECT 100.540 182.085 100.935 182.255 ;
        RECT 100.540 181.955 100.710 182.085 ;
        RECT 99.565 181.625 100.245 181.955 ;
        RECT 100.460 181.625 100.710 181.955 ;
        RECT 100.880 181.455 101.130 181.915 ;
        RECT 101.300 181.640 101.625 182.425 ;
        RECT 101.795 181.625 101.965 183.745 ;
        RECT 102.135 183.625 102.465 184.005 ;
        RECT 102.635 183.455 102.890 183.745 ;
        RECT 102.140 183.285 102.890 183.455 ;
        RECT 102.140 182.295 102.370 183.285 ;
        RECT 103.065 183.255 104.275 184.005 ;
        RECT 104.450 183.460 109.795 184.005 ;
        RECT 102.540 182.465 102.890 183.115 ;
        RECT 103.065 182.545 103.585 183.085 ;
        RECT 103.755 182.715 104.275 183.255 ;
        RECT 102.140 182.125 102.890 182.295 ;
        RECT 102.135 181.455 102.465 181.955 ;
        RECT 102.635 181.625 102.890 182.125 ;
        RECT 103.065 181.455 104.275 182.545 ;
        RECT 106.040 181.890 106.390 183.140 ;
        RECT 107.870 182.630 108.210 183.460 ;
        RECT 109.965 183.205 110.305 183.835 ;
        RECT 110.475 183.205 110.725 184.005 ;
        RECT 110.915 183.355 111.245 183.835 ;
        RECT 111.415 183.545 111.640 184.005 ;
        RECT 111.810 183.355 112.140 183.835 ;
        RECT 109.965 182.595 110.140 183.205 ;
        RECT 110.915 183.185 112.140 183.355 ;
        RECT 112.770 183.225 113.270 183.835 ;
        RECT 114.565 183.280 114.855 184.005 ;
        RECT 115.115 183.455 115.285 183.835 ;
        RECT 115.465 183.625 115.795 184.005 ;
        RECT 115.115 183.285 115.780 183.455 ;
        RECT 115.975 183.330 116.235 183.835 ;
        RECT 110.310 182.845 111.005 183.015 ;
        RECT 110.835 182.595 111.005 182.845 ;
        RECT 111.180 182.815 111.600 183.015 ;
        RECT 111.770 182.815 112.100 183.015 ;
        RECT 112.270 182.815 112.600 183.015 ;
        RECT 112.770 182.595 112.940 183.225 ;
        RECT 113.125 182.765 113.475 183.015 ;
        RECT 115.045 182.735 115.375 183.105 ;
        RECT 115.610 183.030 115.780 183.285 ;
        RECT 115.610 182.700 115.895 183.030 ;
        RECT 104.450 181.455 109.795 181.890 ;
        RECT 109.965 181.625 110.305 182.595 ;
        RECT 110.475 181.455 110.645 182.595 ;
        RECT 110.835 182.425 113.270 182.595 ;
        RECT 110.915 181.455 111.165 182.255 ;
        RECT 111.810 181.625 112.140 182.425 ;
        RECT 112.440 181.455 112.770 182.255 ;
        RECT 112.940 181.625 113.270 182.425 ;
        RECT 114.565 181.455 114.855 182.620 ;
        RECT 115.610 182.555 115.780 182.700 ;
        RECT 115.115 182.385 115.780 182.555 ;
        RECT 116.065 182.530 116.235 183.330 ;
        RECT 117.325 183.235 120.835 184.005 ;
        RECT 121.010 183.460 126.355 184.005 ;
        RECT 115.115 181.625 115.285 182.385 ;
        RECT 115.465 181.455 115.795 182.215 ;
        RECT 115.965 181.625 116.235 182.530 ;
        RECT 117.325 182.545 119.015 183.065 ;
        RECT 119.185 182.715 120.835 183.235 ;
        RECT 117.325 181.455 120.835 182.545 ;
        RECT 122.600 181.890 122.950 183.140 ;
        RECT 124.430 182.630 124.770 183.460 ;
        RECT 126.525 183.255 127.735 184.005 ;
        RECT 126.525 182.545 127.045 183.085 ;
        RECT 127.215 182.715 127.735 183.255 ;
        RECT 121.010 181.455 126.355 181.890 ;
        RECT 126.525 181.455 127.735 182.545 ;
        RECT 20.640 181.285 127.820 181.455 ;
        RECT 20.725 180.195 21.935 181.285 ;
        RECT 20.725 179.485 21.245 180.025 ;
        RECT 21.415 179.655 21.935 180.195 ;
        RECT 22.565 180.195 24.235 181.285 ;
        RECT 22.565 179.675 23.315 180.195 ;
        RECT 24.405 180.120 24.695 181.285 ;
        RECT 24.865 180.195 26.075 181.285 ;
        RECT 26.245 180.195 29.755 181.285 ;
        RECT 29.930 180.850 35.275 181.285 ;
        RECT 23.485 179.505 24.235 180.025 ;
        RECT 24.865 179.655 25.385 180.195 ;
        RECT 20.725 178.735 21.935 179.485 ;
        RECT 22.565 178.735 24.235 179.505 ;
        RECT 25.555 179.485 26.075 180.025 ;
        RECT 26.245 179.675 27.935 180.195 ;
        RECT 28.105 179.505 29.755 180.025 ;
        RECT 31.520 179.600 31.870 180.850 ;
        RECT 35.445 180.210 35.715 181.115 ;
        RECT 35.885 180.525 36.215 181.285 ;
        RECT 36.395 180.355 36.565 181.115 ;
        RECT 24.405 178.735 24.695 179.460 ;
        RECT 24.865 178.735 26.075 179.485 ;
        RECT 26.245 178.735 29.755 179.505 ;
        RECT 33.350 179.280 33.690 180.110 ;
        RECT 35.445 179.410 35.615 180.210 ;
        RECT 35.900 180.185 36.565 180.355 ;
        RECT 35.900 180.040 36.070 180.185 ;
        RECT 35.785 179.710 36.070 180.040 ;
        RECT 36.830 180.145 37.165 181.115 ;
        RECT 37.335 180.145 37.505 181.285 ;
        RECT 37.675 180.945 39.705 181.115 ;
        RECT 35.900 179.455 36.070 179.710 ;
        RECT 36.305 179.635 36.635 180.005 ;
        RECT 36.830 179.475 37.000 180.145 ;
        RECT 37.675 179.975 37.845 180.945 ;
        RECT 37.170 179.645 37.425 179.975 ;
        RECT 37.650 179.645 37.845 179.975 ;
        RECT 38.015 180.605 39.140 180.775 ;
        RECT 37.255 179.475 37.425 179.645 ;
        RECT 38.015 179.475 38.185 180.605 ;
        RECT 29.930 178.735 35.275 179.280 ;
        RECT 35.445 178.905 35.705 179.410 ;
        RECT 35.900 179.285 36.565 179.455 ;
        RECT 35.885 178.735 36.215 179.115 ;
        RECT 36.395 178.905 36.565 179.285 ;
        RECT 36.830 178.905 37.085 179.475 ;
        RECT 37.255 179.305 38.185 179.475 ;
        RECT 38.355 180.265 39.365 180.435 ;
        RECT 38.355 179.465 38.525 180.265 ;
        RECT 38.730 179.925 39.005 180.065 ;
        RECT 38.725 179.755 39.005 179.925 ;
        RECT 38.010 179.270 38.185 179.305 ;
        RECT 37.255 178.735 37.585 179.135 ;
        RECT 38.010 178.905 38.540 179.270 ;
        RECT 38.730 178.905 39.005 179.755 ;
        RECT 39.175 178.905 39.365 180.265 ;
        RECT 39.535 180.280 39.705 180.945 ;
        RECT 39.875 180.525 40.045 181.285 ;
        RECT 40.280 180.525 40.795 180.935 ;
        RECT 40.970 180.850 46.315 181.285 ;
        RECT 39.535 180.090 40.285 180.280 ;
        RECT 40.455 179.715 40.795 180.525 ;
        RECT 39.565 179.545 40.795 179.715 ;
        RECT 42.560 179.600 42.910 180.850 ;
        RECT 46.485 180.145 46.825 181.115 ;
        RECT 46.995 180.145 47.165 181.285 ;
        RECT 47.435 180.485 47.685 181.285 ;
        RECT 48.330 180.315 48.660 181.115 ;
        RECT 48.960 180.485 49.290 181.285 ;
        RECT 49.460 180.315 49.790 181.115 ;
        RECT 47.355 180.145 49.790 180.315 ;
        RECT 39.545 178.735 40.055 179.270 ;
        RECT 40.275 178.940 40.520 179.545 ;
        RECT 44.390 179.280 44.730 180.110 ;
        RECT 46.485 179.535 46.660 180.145 ;
        RECT 47.355 179.895 47.525 180.145 ;
        RECT 46.830 179.725 47.525 179.895 ;
        RECT 47.700 179.725 48.120 179.925 ;
        RECT 48.290 179.725 48.620 179.925 ;
        RECT 48.790 179.725 49.120 179.925 ;
        RECT 40.970 178.735 46.315 179.280 ;
        RECT 46.485 178.905 46.825 179.535 ;
        RECT 46.995 178.735 47.245 179.535 ;
        RECT 47.435 179.385 48.660 179.555 ;
        RECT 47.435 178.905 47.765 179.385 ;
        RECT 47.935 178.735 48.160 179.195 ;
        RECT 48.330 178.905 48.660 179.385 ;
        RECT 49.290 179.515 49.460 180.145 ;
        RECT 50.165 180.120 50.455 181.285 ;
        RECT 51.085 180.195 52.755 181.285 ;
        RECT 52.925 180.525 53.440 180.935 ;
        RECT 53.675 180.525 53.845 181.285 ;
        RECT 54.015 180.945 56.045 181.115 ;
        RECT 49.645 179.725 49.995 179.975 ;
        RECT 51.085 179.675 51.835 180.195 ;
        RECT 49.290 178.905 49.790 179.515 ;
        RECT 52.005 179.505 52.755 180.025 ;
        RECT 52.925 179.715 53.265 180.525 ;
        RECT 54.015 180.280 54.185 180.945 ;
        RECT 54.580 180.605 55.705 180.775 ;
        RECT 53.435 180.090 54.185 180.280 ;
        RECT 54.355 180.265 55.365 180.435 ;
        RECT 52.925 179.545 54.155 179.715 ;
        RECT 50.165 178.735 50.455 179.460 ;
        RECT 51.085 178.735 52.755 179.505 ;
        RECT 53.200 178.940 53.445 179.545 ;
        RECT 53.665 178.735 54.175 179.270 ;
        RECT 54.355 178.905 54.545 180.265 ;
        RECT 54.715 179.245 54.990 180.065 ;
        RECT 55.195 179.465 55.365 180.265 ;
        RECT 55.535 179.475 55.705 180.605 ;
        RECT 55.875 179.975 56.045 180.945 ;
        RECT 56.215 180.145 56.385 181.285 ;
        RECT 56.555 180.145 56.890 181.115 ;
        RECT 55.875 179.645 56.070 179.975 ;
        RECT 56.295 179.645 56.550 179.975 ;
        RECT 56.295 179.475 56.465 179.645 ;
        RECT 56.720 179.475 56.890 180.145 ;
        RECT 57.065 180.525 57.580 180.935 ;
        RECT 57.815 180.525 57.985 181.285 ;
        RECT 58.155 180.945 60.185 181.115 ;
        RECT 57.065 179.715 57.405 180.525 ;
        RECT 58.155 180.280 58.325 180.945 ;
        RECT 58.720 180.605 59.845 180.775 ;
        RECT 57.575 180.090 58.325 180.280 ;
        RECT 58.495 180.265 59.505 180.435 ;
        RECT 57.065 179.545 58.295 179.715 ;
        RECT 55.535 179.305 56.465 179.475 ;
        RECT 55.535 179.270 55.710 179.305 ;
        RECT 54.715 179.075 54.995 179.245 ;
        RECT 54.715 178.905 54.990 179.075 ;
        RECT 55.180 178.905 55.710 179.270 ;
        RECT 56.135 178.735 56.465 179.135 ;
        RECT 56.635 178.905 56.890 179.475 ;
        RECT 57.340 178.940 57.585 179.545 ;
        RECT 57.805 178.735 58.315 179.270 ;
        RECT 58.495 178.905 58.685 180.265 ;
        RECT 58.855 179.585 59.130 180.065 ;
        RECT 58.855 179.415 59.135 179.585 ;
        RECT 59.335 179.465 59.505 180.265 ;
        RECT 59.675 179.475 59.845 180.605 ;
        RECT 60.015 179.975 60.185 180.945 ;
        RECT 60.355 180.145 60.525 181.285 ;
        RECT 60.695 180.145 61.030 181.115 ;
        RECT 61.260 180.415 61.545 181.285 ;
        RECT 61.715 180.655 61.975 181.115 ;
        RECT 62.150 180.825 62.405 181.285 ;
        RECT 62.575 180.655 62.835 181.115 ;
        RECT 61.715 180.485 62.835 180.655 ;
        RECT 63.005 180.485 63.315 181.285 ;
        RECT 61.715 180.235 61.975 180.485 ;
        RECT 63.485 180.315 63.795 181.115 ;
        RECT 60.015 179.645 60.210 179.975 ;
        RECT 60.435 179.645 60.690 179.975 ;
        RECT 60.435 179.475 60.605 179.645 ;
        RECT 60.860 179.475 61.030 180.145 ;
        RECT 58.855 178.905 59.130 179.415 ;
        RECT 59.675 179.305 60.605 179.475 ;
        RECT 59.675 179.270 59.850 179.305 ;
        RECT 59.320 178.905 59.850 179.270 ;
        RECT 60.275 178.735 60.605 179.135 ;
        RECT 60.775 178.905 61.030 179.475 ;
        RECT 61.220 180.065 61.975 180.235 ;
        RECT 62.765 180.145 63.795 180.315 ;
        RECT 61.220 179.555 61.625 180.065 ;
        RECT 62.765 179.895 62.935 180.145 ;
        RECT 61.795 179.725 62.935 179.895 ;
        RECT 61.220 179.385 62.870 179.555 ;
        RECT 63.105 179.405 63.455 179.975 ;
        RECT 61.265 178.735 61.545 179.215 ;
        RECT 61.715 178.995 61.975 179.385 ;
        RECT 62.150 178.735 62.405 179.215 ;
        RECT 62.575 178.995 62.870 179.385 ;
        RECT 63.625 179.235 63.795 180.145 ;
        RECT 63.965 180.195 67.475 181.285 ;
        RECT 63.965 179.675 65.655 180.195 ;
        RECT 67.650 180.135 67.910 181.285 ;
        RECT 68.085 180.210 68.340 181.115 ;
        RECT 68.510 180.525 68.840 181.285 ;
        RECT 69.055 180.355 69.225 181.115 ;
        RECT 65.825 179.505 67.475 180.025 ;
        RECT 63.050 178.735 63.325 179.215 ;
        RECT 63.495 178.905 63.795 179.235 ;
        RECT 63.965 178.735 67.475 179.505 ;
        RECT 67.650 178.735 67.910 179.575 ;
        RECT 68.085 179.480 68.255 180.210 ;
        RECT 68.510 180.185 69.225 180.355 ;
        RECT 69.575 180.355 69.745 181.115 ;
        RECT 69.960 180.525 70.290 181.285 ;
        RECT 69.575 180.185 70.290 180.355 ;
        RECT 70.460 180.210 70.715 181.115 ;
        RECT 68.510 179.975 68.680 180.185 ;
        RECT 68.425 179.645 68.680 179.975 ;
        RECT 68.085 178.905 68.340 179.480 ;
        RECT 68.510 179.455 68.680 179.645 ;
        RECT 68.960 179.635 69.315 180.005 ;
        RECT 69.485 179.635 69.840 180.005 ;
        RECT 70.120 179.975 70.290 180.185 ;
        RECT 70.120 179.645 70.375 179.975 ;
        RECT 70.120 179.455 70.290 179.645 ;
        RECT 70.545 179.480 70.715 180.210 ;
        RECT 70.890 180.135 71.150 181.285 ;
        RECT 72.245 180.195 75.755 181.285 ;
        RECT 72.245 179.675 73.935 180.195 ;
        RECT 75.925 180.120 76.215 181.285 ;
        RECT 76.845 180.195 80.355 181.285 ;
        RECT 80.525 180.315 80.835 181.115 ;
        RECT 81.005 180.485 81.315 181.285 ;
        RECT 81.485 180.655 81.745 181.115 ;
        RECT 81.915 180.825 82.170 181.285 ;
        RECT 82.345 180.655 82.605 181.115 ;
        RECT 81.485 180.485 82.605 180.655 ;
        RECT 68.510 179.285 69.225 179.455 ;
        RECT 68.510 178.735 68.840 179.115 ;
        RECT 69.055 178.905 69.225 179.285 ;
        RECT 69.575 179.285 70.290 179.455 ;
        RECT 69.575 178.905 69.745 179.285 ;
        RECT 69.960 178.735 70.290 179.115 ;
        RECT 70.460 178.905 70.715 179.480 ;
        RECT 70.890 178.735 71.150 179.575 ;
        RECT 74.105 179.505 75.755 180.025 ;
        RECT 76.845 179.675 78.535 180.195 ;
        RECT 80.525 180.145 81.555 180.315 ;
        RECT 78.705 179.505 80.355 180.025 ;
        RECT 72.245 178.735 75.755 179.505 ;
        RECT 75.925 178.735 76.215 179.460 ;
        RECT 76.845 178.735 80.355 179.505 ;
        RECT 80.525 179.235 80.695 180.145 ;
        RECT 80.865 179.405 81.215 179.975 ;
        RECT 81.385 179.895 81.555 180.145 ;
        RECT 82.345 180.235 82.605 180.485 ;
        RECT 82.775 180.415 83.060 181.285 ;
        RECT 82.345 180.065 83.100 180.235 ;
        RECT 81.385 179.725 82.525 179.895 ;
        RECT 82.695 179.555 83.100 180.065 ;
        RECT 81.450 179.385 83.100 179.555 ;
        RECT 83.285 180.145 83.625 181.115 ;
        RECT 83.795 180.145 83.965 181.285 ;
        RECT 84.235 180.485 84.485 181.285 ;
        RECT 85.130 180.315 85.460 181.115 ;
        RECT 85.760 180.485 86.090 181.285 ;
        RECT 86.260 180.315 86.590 181.115 ;
        RECT 87.890 180.850 93.235 181.285 ;
        RECT 84.155 180.145 86.590 180.315 ;
        RECT 83.285 179.535 83.460 180.145 ;
        RECT 84.155 179.895 84.325 180.145 ;
        RECT 83.630 179.725 84.325 179.895 ;
        RECT 84.500 179.725 84.920 179.925 ;
        RECT 85.090 179.725 85.420 179.925 ;
        RECT 85.590 179.725 85.920 179.925 ;
        RECT 80.525 178.905 80.825 179.235 ;
        RECT 80.995 178.735 81.270 179.215 ;
        RECT 81.450 178.995 81.745 179.385 ;
        RECT 81.915 178.735 82.170 179.215 ;
        RECT 82.345 178.995 82.605 179.385 ;
        RECT 82.775 178.735 83.055 179.215 ;
        RECT 83.285 178.905 83.625 179.535 ;
        RECT 83.795 178.735 84.045 179.535 ;
        RECT 84.235 179.385 85.460 179.555 ;
        RECT 84.235 178.905 84.565 179.385 ;
        RECT 84.735 178.735 84.960 179.195 ;
        RECT 85.130 178.905 85.460 179.385 ;
        RECT 86.090 179.515 86.260 180.145 ;
        RECT 86.445 179.725 86.795 179.975 ;
        RECT 89.480 179.600 89.830 180.850 ;
        RECT 93.495 180.355 93.665 181.115 ;
        RECT 93.845 180.525 94.175 181.285 ;
        RECT 93.495 180.185 94.160 180.355 ;
        RECT 94.345 180.210 94.615 181.115 ;
        RECT 86.090 178.905 86.590 179.515 ;
        RECT 91.310 179.280 91.650 180.110 ;
        RECT 93.990 180.040 94.160 180.185 ;
        RECT 93.425 179.635 93.755 180.005 ;
        RECT 93.990 179.710 94.275 180.040 ;
        RECT 93.990 179.455 94.160 179.710 ;
        RECT 93.495 179.285 94.160 179.455 ;
        RECT 94.445 179.410 94.615 180.210 ;
        RECT 94.785 180.195 96.455 181.285 ;
        RECT 94.785 179.675 95.535 180.195 ;
        RECT 96.685 180.145 96.895 181.285 ;
        RECT 97.065 180.135 97.395 181.115 ;
        RECT 97.565 180.145 97.795 181.285 ;
        RECT 98.465 180.195 100.135 181.285 ;
        RECT 100.395 180.355 100.565 181.115 ;
        RECT 100.745 180.525 101.075 181.285 ;
        RECT 95.705 179.505 96.455 180.025 ;
        RECT 87.890 178.735 93.235 179.280 ;
        RECT 93.495 178.905 93.665 179.285 ;
        RECT 93.845 178.735 94.175 179.115 ;
        RECT 94.355 178.905 94.615 179.410 ;
        RECT 94.785 178.735 96.455 179.505 ;
        RECT 96.685 178.735 96.895 179.555 ;
        RECT 97.065 179.535 97.315 180.135 ;
        RECT 97.485 179.725 97.815 179.975 ;
        RECT 98.465 179.675 99.215 180.195 ;
        RECT 100.395 180.185 101.060 180.355 ;
        RECT 101.245 180.210 101.515 181.115 ;
        RECT 100.890 180.040 101.060 180.185 ;
        RECT 97.065 178.905 97.395 179.535 ;
        RECT 97.565 178.735 97.795 179.555 ;
        RECT 99.385 179.505 100.135 180.025 ;
        RECT 100.325 179.635 100.655 180.005 ;
        RECT 100.890 179.710 101.175 180.040 ;
        RECT 98.465 178.735 100.135 179.505 ;
        RECT 100.890 179.455 101.060 179.710 ;
        RECT 100.395 179.285 101.060 179.455 ;
        RECT 101.345 179.410 101.515 180.210 ;
        RECT 101.685 180.120 101.975 181.285 ;
        RECT 102.205 180.145 102.415 181.285 ;
        RECT 102.585 180.135 102.915 181.115 ;
        RECT 103.085 180.145 103.315 181.285 ;
        RECT 103.985 180.195 106.575 181.285 ;
        RECT 100.395 178.905 100.565 179.285 ;
        RECT 100.745 178.735 101.075 179.115 ;
        RECT 101.255 178.905 101.515 179.410 ;
        RECT 101.685 178.735 101.975 179.460 ;
        RECT 102.205 178.735 102.415 179.555 ;
        RECT 102.585 179.535 102.835 180.135 ;
        RECT 103.005 179.725 103.335 179.975 ;
        RECT 103.985 179.675 105.195 180.195 ;
        RECT 106.745 180.145 107.085 181.115 ;
        RECT 107.255 180.145 107.425 181.285 ;
        RECT 107.695 180.485 107.945 181.285 ;
        RECT 108.590 180.315 108.920 181.115 ;
        RECT 109.220 180.485 109.550 181.285 ;
        RECT 109.720 180.315 110.050 181.115 ;
        RECT 107.615 180.145 110.050 180.315 ;
        RECT 110.630 180.315 110.960 181.115 ;
        RECT 111.130 180.485 111.460 181.285 ;
        RECT 111.760 180.315 112.090 181.115 ;
        RECT 112.735 180.485 112.985 181.285 ;
        RECT 110.630 180.145 113.065 180.315 ;
        RECT 113.255 180.145 113.425 181.285 ;
        RECT 113.595 180.145 113.935 181.115 ;
        RECT 102.585 178.905 102.915 179.535 ;
        RECT 103.085 178.735 103.315 179.555 ;
        RECT 105.365 179.505 106.575 180.025 ;
        RECT 103.985 178.735 106.575 179.505 ;
        RECT 106.745 179.535 106.920 180.145 ;
        RECT 107.615 179.895 107.785 180.145 ;
        RECT 107.090 179.725 107.785 179.895 ;
        RECT 107.960 179.725 108.380 179.925 ;
        RECT 108.550 179.725 108.880 179.925 ;
        RECT 109.050 179.725 109.380 179.925 ;
        RECT 106.745 178.905 107.085 179.535 ;
        RECT 107.255 178.735 107.505 179.535 ;
        RECT 107.695 179.385 108.920 179.555 ;
        RECT 107.695 178.905 108.025 179.385 ;
        RECT 108.195 178.735 108.420 179.195 ;
        RECT 108.590 178.905 108.920 179.385 ;
        RECT 109.550 179.515 109.720 180.145 ;
        RECT 109.905 179.725 110.255 179.975 ;
        RECT 110.425 179.725 110.775 179.975 ;
        RECT 110.960 179.515 111.130 180.145 ;
        RECT 111.300 179.725 111.630 179.925 ;
        RECT 111.800 179.725 112.130 179.925 ;
        RECT 112.300 179.725 112.720 179.925 ;
        RECT 112.895 179.895 113.065 180.145 ;
        RECT 112.895 179.725 113.590 179.895 ;
        RECT 109.550 178.905 110.050 179.515 ;
        RECT 110.630 178.905 111.130 179.515 ;
        RECT 111.760 179.385 112.985 179.555 ;
        RECT 113.760 179.535 113.935 180.145 ;
        RECT 114.105 180.195 115.775 181.285 ;
        RECT 114.105 179.675 114.855 180.195 ;
        RECT 115.985 180.145 116.215 181.285 ;
        RECT 116.385 180.135 116.715 181.115 ;
        RECT 116.885 180.145 117.095 181.285 ;
        RECT 111.760 178.905 112.090 179.385 ;
        RECT 112.260 178.735 112.485 179.195 ;
        RECT 112.655 178.905 112.985 179.385 ;
        RECT 113.175 178.735 113.425 179.535 ;
        RECT 113.595 178.905 113.935 179.535 ;
        RECT 115.025 179.505 115.775 180.025 ;
        RECT 115.965 179.725 116.295 179.975 ;
        RECT 114.105 178.735 115.775 179.505 ;
        RECT 115.985 178.735 116.215 179.555 ;
        RECT 116.465 179.535 116.715 180.135 ;
        RECT 117.330 180.095 117.585 180.975 ;
        RECT 117.755 180.145 118.060 181.285 ;
        RECT 118.400 180.905 118.730 181.285 ;
        RECT 118.910 180.735 119.080 181.025 ;
        RECT 119.250 180.825 119.500 181.285 ;
        RECT 118.280 180.565 119.080 180.735 ;
        RECT 119.670 180.775 120.540 181.115 ;
        RECT 116.385 178.905 116.715 179.535 ;
        RECT 116.885 178.735 117.095 179.555 ;
        RECT 117.330 179.445 117.540 180.095 ;
        RECT 118.280 179.975 118.450 180.565 ;
        RECT 119.670 180.395 119.840 180.775 ;
        RECT 120.775 180.655 120.945 181.115 ;
        RECT 121.115 180.825 121.485 181.285 ;
        RECT 121.780 180.685 121.950 181.025 ;
        RECT 122.120 180.855 122.450 181.285 ;
        RECT 122.685 180.685 122.855 181.025 ;
        RECT 118.620 180.225 119.840 180.395 ;
        RECT 120.010 180.315 120.470 180.605 ;
        RECT 120.775 180.485 121.335 180.655 ;
        RECT 121.780 180.515 122.855 180.685 ;
        RECT 123.025 180.785 123.705 181.115 ;
        RECT 123.920 180.785 124.170 181.115 ;
        RECT 124.340 180.825 124.590 181.285 ;
        RECT 121.165 180.345 121.335 180.485 ;
        RECT 120.010 180.305 120.975 180.315 ;
        RECT 119.670 180.135 119.840 180.225 ;
        RECT 120.300 180.145 120.975 180.305 ;
        RECT 117.710 179.945 118.450 179.975 ;
        RECT 117.710 179.645 118.625 179.945 ;
        RECT 118.300 179.470 118.625 179.645 ;
        RECT 117.330 178.915 117.585 179.445 ;
        RECT 117.755 178.735 118.060 179.195 ;
        RECT 118.305 179.115 118.625 179.470 ;
        RECT 118.795 179.685 119.335 180.055 ;
        RECT 119.670 179.965 120.075 180.135 ;
        RECT 118.795 179.285 119.035 179.685 ;
        RECT 119.515 179.515 119.735 179.795 ;
        RECT 119.205 179.345 119.735 179.515 ;
        RECT 119.205 179.115 119.375 179.345 ;
        RECT 119.905 179.185 120.075 179.965 ;
        RECT 120.245 179.355 120.595 179.975 ;
        RECT 120.765 179.355 120.975 180.145 ;
        RECT 121.165 180.175 122.665 180.345 ;
        RECT 121.165 179.485 121.335 180.175 ;
        RECT 123.025 180.005 123.195 180.785 ;
        RECT 124.000 180.655 124.170 180.785 ;
        RECT 121.505 179.835 123.195 180.005 ;
        RECT 123.365 180.225 123.830 180.615 ;
        RECT 124.000 180.485 124.395 180.655 ;
        RECT 121.505 179.655 121.675 179.835 ;
        RECT 118.305 178.945 119.375 179.115 ;
        RECT 119.545 178.735 119.735 179.175 ;
        RECT 119.905 178.905 120.855 179.185 ;
        RECT 121.165 179.095 121.425 179.485 ;
        RECT 121.845 179.415 122.635 179.665 ;
        RECT 121.075 178.925 121.425 179.095 ;
        RECT 121.635 178.735 121.965 179.195 ;
        RECT 122.840 179.125 123.010 179.835 ;
        RECT 123.365 179.635 123.535 180.225 ;
        RECT 123.180 179.415 123.535 179.635 ;
        RECT 123.705 179.415 124.055 180.035 ;
        RECT 124.225 179.125 124.395 180.485 ;
        RECT 124.760 180.315 125.085 181.100 ;
        RECT 124.565 179.265 125.025 180.315 ;
        RECT 122.840 178.955 123.695 179.125 ;
        RECT 123.900 178.955 124.395 179.125 ;
        RECT 124.565 178.735 124.895 179.095 ;
        RECT 125.255 178.995 125.425 181.115 ;
        RECT 125.595 180.785 125.925 181.285 ;
        RECT 126.095 180.615 126.350 181.115 ;
        RECT 125.600 180.445 126.350 180.615 ;
        RECT 125.600 179.455 125.830 180.445 ;
        RECT 126.000 179.625 126.350 180.275 ;
        RECT 126.525 180.195 127.735 181.285 ;
        RECT 126.525 179.655 127.045 180.195 ;
        RECT 127.215 179.485 127.735 180.025 ;
        RECT 125.600 179.285 126.350 179.455 ;
        RECT 125.595 178.735 125.925 179.115 ;
        RECT 126.095 178.995 126.350 179.285 ;
        RECT 126.525 178.735 127.735 179.485 ;
        RECT 20.640 178.565 127.820 178.735 ;
        RECT 20.725 177.815 21.935 178.565 ;
        RECT 20.725 177.275 21.245 177.815 ;
        RECT 22.565 177.795 26.075 178.565 ;
        RECT 26.250 178.020 31.595 178.565 ;
        RECT 31.770 178.020 37.115 178.565 ;
        RECT 21.415 177.105 21.935 177.645 ;
        RECT 20.725 176.015 21.935 177.105 ;
        RECT 22.565 177.105 24.255 177.625 ;
        RECT 24.425 177.275 26.075 177.795 ;
        RECT 22.565 176.015 26.075 177.105 ;
        RECT 27.840 176.450 28.190 177.700 ;
        RECT 29.670 177.190 30.010 178.020 ;
        RECT 33.360 176.450 33.710 177.700 ;
        RECT 35.190 177.190 35.530 178.020 ;
        RECT 37.285 177.840 37.575 178.565 ;
        RECT 37.745 177.815 38.955 178.565 ;
        RECT 26.250 176.015 31.595 176.450 ;
        RECT 31.770 176.015 37.115 176.450 ;
        RECT 37.285 176.015 37.575 177.180 ;
        RECT 37.745 177.105 38.265 177.645 ;
        RECT 38.435 177.275 38.955 177.815 ;
        RECT 39.330 177.785 39.830 178.395 ;
        RECT 39.125 177.325 39.475 177.575 ;
        RECT 39.660 177.155 39.830 177.785 ;
        RECT 40.460 177.915 40.790 178.395 ;
        RECT 40.960 178.105 41.185 178.565 ;
        RECT 41.355 177.915 41.685 178.395 ;
        RECT 40.460 177.745 41.685 177.915 ;
        RECT 41.875 177.765 42.125 178.565 ;
        RECT 42.295 177.765 42.635 178.395 ;
        RECT 40.000 177.375 40.330 177.575 ;
        RECT 40.500 177.375 40.830 177.575 ;
        RECT 41.000 177.375 41.420 177.575 ;
        RECT 41.595 177.405 42.290 177.575 ;
        RECT 41.595 177.155 41.765 177.405 ;
        RECT 42.460 177.205 42.635 177.765 ;
        RECT 42.405 177.155 42.635 177.205 ;
        RECT 37.745 176.015 38.955 177.105 ;
        RECT 39.330 176.985 41.765 177.155 ;
        RECT 39.330 176.185 39.660 176.985 ;
        RECT 39.830 176.015 40.160 176.815 ;
        RECT 40.460 176.185 40.790 176.985 ;
        RECT 41.435 176.015 41.685 176.815 ;
        RECT 41.955 176.015 42.125 177.155 ;
        RECT 42.295 176.185 42.635 177.155 ;
        RECT 42.805 177.765 43.145 178.395 ;
        RECT 43.315 177.765 43.565 178.565 ;
        RECT 43.755 177.915 44.085 178.395 ;
        RECT 44.255 178.105 44.480 178.565 ;
        RECT 44.650 177.915 44.980 178.395 ;
        RECT 42.805 177.155 42.980 177.765 ;
        RECT 43.755 177.745 44.980 177.915 ;
        RECT 45.610 177.785 46.110 178.395 ;
        RECT 46.690 177.785 47.190 178.395 ;
        RECT 43.150 177.405 43.845 177.575 ;
        RECT 43.675 177.155 43.845 177.405 ;
        RECT 44.020 177.375 44.440 177.575 ;
        RECT 44.610 177.375 44.940 177.575 ;
        RECT 45.110 177.375 45.440 177.575 ;
        RECT 45.610 177.155 45.780 177.785 ;
        RECT 45.965 177.325 46.315 177.575 ;
        RECT 46.485 177.325 46.835 177.575 ;
        RECT 47.020 177.155 47.190 177.785 ;
        RECT 47.820 177.915 48.150 178.395 ;
        RECT 48.320 178.105 48.545 178.565 ;
        RECT 48.715 177.915 49.045 178.395 ;
        RECT 47.820 177.745 49.045 177.915 ;
        RECT 49.235 177.765 49.485 178.565 ;
        RECT 49.655 177.765 49.995 178.395 ;
        RECT 50.370 177.785 50.870 178.395 ;
        RECT 47.360 177.375 47.690 177.575 ;
        RECT 47.860 177.375 48.190 177.575 ;
        RECT 48.360 177.375 48.780 177.575 ;
        RECT 48.955 177.405 49.650 177.575 ;
        RECT 48.955 177.155 49.125 177.405 ;
        RECT 49.820 177.155 49.995 177.765 ;
        RECT 50.165 177.325 50.515 177.575 ;
        RECT 50.700 177.155 50.870 177.785 ;
        RECT 51.500 177.915 51.830 178.395 ;
        RECT 52.000 178.105 52.225 178.565 ;
        RECT 52.395 177.915 52.725 178.395 ;
        RECT 51.500 177.745 52.725 177.915 ;
        RECT 52.915 177.765 53.165 178.565 ;
        RECT 53.335 177.765 53.675 178.395 ;
        RECT 51.040 177.375 51.370 177.575 ;
        RECT 51.540 177.375 51.870 177.575 ;
        RECT 52.040 177.375 52.460 177.575 ;
        RECT 52.635 177.405 53.330 177.575 ;
        RECT 52.635 177.155 52.805 177.405 ;
        RECT 53.500 177.155 53.675 177.765 ;
        RECT 42.805 176.185 43.145 177.155 ;
        RECT 43.315 176.015 43.485 177.155 ;
        RECT 43.675 176.985 46.110 177.155 ;
        RECT 43.755 176.015 44.005 176.815 ;
        RECT 44.650 176.185 44.980 176.985 ;
        RECT 45.280 176.015 45.610 176.815 ;
        RECT 45.780 176.185 46.110 176.985 ;
        RECT 46.690 176.985 49.125 177.155 ;
        RECT 46.690 176.185 47.020 176.985 ;
        RECT 47.190 176.015 47.520 176.815 ;
        RECT 47.820 176.185 48.150 176.985 ;
        RECT 48.795 176.015 49.045 176.815 ;
        RECT 49.315 176.015 49.485 177.155 ;
        RECT 49.655 176.185 49.995 177.155 ;
        RECT 50.370 176.985 52.805 177.155 ;
        RECT 50.370 176.185 50.700 176.985 ;
        RECT 50.870 176.015 51.200 176.815 ;
        RECT 51.500 176.185 51.830 176.985 ;
        RECT 52.475 176.015 52.725 176.815 ;
        RECT 52.995 176.015 53.165 177.155 ;
        RECT 53.335 176.185 53.675 177.155 ;
        RECT 53.850 177.855 54.105 178.385 ;
        RECT 54.275 178.105 54.580 178.565 ;
        RECT 54.825 178.185 55.895 178.355 ;
        RECT 53.850 177.205 54.060 177.855 ;
        RECT 54.825 177.830 55.145 178.185 ;
        RECT 54.820 177.655 55.145 177.830 ;
        RECT 54.230 177.355 55.145 177.655 ;
        RECT 55.315 177.615 55.555 178.015 ;
        RECT 55.725 177.955 55.895 178.185 ;
        RECT 56.065 178.125 56.255 178.565 ;
        RECT 56.425 178.115 57.375 178.395 ;
        RECT 57.595 178.205 57.945 178.375 ;
        RECT 55.725 177.785 56.255 177.955 ;
        RECT 54.230 177.325 54.970 177.355 ;
        RECT 53.850 176.325 54.105 177.205 ;
        RECT 54.275 176.015 54.580 177.155 ;
        RECT 54.800 176.735 54.970 177.325 ;
        RECT 55.315 177.245 55.855 177.615 ;
        RECT 56.035 177.505 56.255 177.785 ;
        RECT 56.425 177.335 56.595 178.115 ;
        RECT 56.190 177.165 56.595 177.335 ;
        RECT 56.765 177.325 57.115 177.945 ;
        RECT 56.190 177.075 56.360 177.165 ;
        RECT 57.285 177.155 57.495 177.945 ;
        RECT 55.140 176.905 56.360 177.075 ;
        RECT 56.820 176.995 57.495 177.155 ;
        RECT 54.800 176.565 55.600 176.735 ;
        RECT 54.920 176.015 55.250 176.395 ;
        RECT 55.430 176.275 55.600 176.565 ;
        RECT 56.190 176.525 56.360 176.905 ;
        RECT 56.530 176.985 57.495 176.995 ;
        RECT 57.685 177.815 57.945 178.205 ;
        RECT 58.155 178.105 58.485 178.565 ;
        RECT 59.360 178.175 60.215 178.345 ;
        RECT 60.420 178.175 60.915 178.345 ;
        RECT 61.085 178.205 61.415 178.565 ;
        RECT 57.685 177.125 57.855 177.815 ;
        RECT 58.025 177.465 58.195 177.645 ;
        RECT 58.365 177.635 59.155 177.885 ;
        RECT 59.360 177.465 59.530 178.175 ;
        RECT 59.700 177.665 60.055 177.885 ;
        RECT 58.025 177.295 59.715 177.465 ;
        RECT 56.530 176.695 56.990 176.985 ;
        RECT 57.685 176.955 59.185 177.125 ;
        RECT 57.685 176.815 57.855 176.955 ;
        RECT 57.295 176.645 57.855 176.815 ;
        RECT 55.770 176.015 56.020 176.475 ;
        RECT 56.190 176.185 57.060 176.525 ;
        RECT 57.295 176.185 57.465 176.645 ;
        RECT 58.300 176.615 59.375 176.785 ;
        RECT 57.635 176.015 58.005 176.475 ;
        RECT 58.300 176.275 58.470 176.615 ;
        RECT 58.640 176.015 58.970 176.445 ;
        RECT 59.205 176.275 59.375 176.615 ;
        RECT 59.545 176.515 59.715 177.295 ;
        RECT 59.885 177.075 60.055 177.665 ;
        RECT 60.225 177.265 60.575 177.885 ;
        RECT 59.885 176.685 60.350 177.075 ;
        RECT 60.745 176.815 60.915 178.175 ;
        RECT 61.085 176.985 61.545 178.035 ;
        RECT 60.520 176.645 60.915 176.815 ;
        RECT 60.520 176.515 60.690 176.645 ;
        RECT 59.545 176.185 60.225 176.515 ;
        RECT 60.440 176.185 60.690 176.515 ;
        RECT 60.860 176.015 61.110 176.475 ;
        RECT 61.280 176.200 61.605 176.985 ;
        RECT 61.775 176.185 61.945 178.305 ;
        RECT 62.115 178.185 62.445 178.565 ;
        RECT 62.615 178.015 62.870 178.305 ;
        RECT 62.120 177.845 62.870 178.015 ;
        RECT 62.120 176.855 62.350 177.845 ;
        RECT 63.045 177.840 63.335 178.565 ;
        RECT 63.505 177.890 63.765 178.395 ;
        RECT 63.945 178.185 64.275 178.565 ;
        RECT 64.455 178.015 64.625 178.395 ;
        RECT 62.520 177.025 62.870 177.675 ;
        RECT 62.120 176.685 62.870 176.855 ;
        RECT 62.115 176.015 62.445 176.515 ;
        RECT 62.615 176.185 62.870 176.685 ;
        RECT 63.045 176.015 63.335 177.180 ;
        RECT 63.505 177.090 63.675 177.890 ;
        RECT 63.960 177.845 64.625 178.015 ;
        RECT 63.960 177.590 64.130 177.845 ;
        RECT 65.810 177.725 66.070 178.565 ;
        RECT 66.245 177.820 66.500 178.395 ;
        RECT 66.670 178.185 67.000 178.565 ;
        RECT 67.215 178.015 67.385 178.395 ;
        RECT 67.915 178.170 68.245 178.565 ;
        RECT 66.670 177.845 67.385 178.015 ;
        RECT 68.415 177.995 68.615 178.350 ;
        RECT 68.785 178.165 69.115 178.565 ;
        RECT 69.285 177.995 69.485 178.340 ;
        RECT 63.845 177.260 64.130 177.590 ;
        RECT 64.365 177.295 64.695 177.665 ;
        RECT 63.960 177.115 64.130 177.260 ;
        RECT 63.505 176.185 63.775 177.090 ;
        RECT 63.960 176.945 64.625 177.115 ;
        RECT 63.945 176.015 64.275 176.775 ;
        RECT 64.455 176.185 64.625 176.945 ;
        RECT 65.810 176.015 66.070 177.165 ;
        RECT 66.245 177.090 66.415 177.820 ;
        RECT 66.670 177.655 66.840 177.845 ;
        RECT 67.645 177.825 69.485 177.995 ;
        RECT 69.655 177.825 69.985 178.565 ;
        RECT 70.220 177.995 70.390 178.245 ;
        RECT 71.135 178.170 71.465 178.565 ;
        RECT 71.635 177.995 71.835 178.350 ;
        RECT 72.005 178.165 72.335 178.565 ;
        RECT 72.505 177.995 72.705 178.340 ;
        RECT 70.220 177.825 70.695 177.995 ;
        RECT 66.585 177.325 66.840 177.655 ;
        RECT 66.670 177.115 66.840 177.325 ;
        RECT 67.120 177.295 67.475 177.665 ;
        RECT 66.245 176.185 66.500 177.090 ;
        RECT 66.670 176.945 67.385 177.115 ;
        RECT 66.670 176.015 67.000 176.775 ;
        RECT 67.215 176.185 67.385 176.945 ;
        RECT 67.645 176.200 67.905 177.825 ;
        RECT 68.085 176.855 68.305 177.655 ;
        RECT 68.545 177.035 68.845 177.655 ;
        RECT 69.015 177.035 69.345 177.655 ;
        RECT 69.515 177.035 69.835 177.655 ;
        RECT 70.005 177.035 70.355 177.655 ;
        RECT 70.525 176.855 70.695 177.825 ;
        RECT 68.085 176.645 70.695 176.855 ;
        RECT 70.865 177.825 72.705 177.995 ;
        RECT 72.875 177.825 73.205 178.565 ;
        RECT 73.440 177.995 73.610 178.245 ;
        RECT 74.175 178.015 74.345 178.395 ;
        RECT 74.560 178.185 74.890 178.565 ;
        RECT 73.440 177.825 73.915 177.995 ;
        RECT 74.175 177.845 74.890 178.015 ;
        RECT 69.655 176.015 69.985 176.465 ;
        RECT 70.865 176.200 71.125 177.825 ;
        RECT 71.305 176.855 71.525 177.655 ;
        RECT 71.765 177.035 72.065 177.655 ;
        RECT 72.235 177.035 72.565 177.655 ;
        RECT 72.735 177.035 73.055 177.655 ;
        RECT 73.225 177.035 73.575 177.655 ;
        RECT 73.745 176.855 73.915 177.825 ;
        RECT 74.085 177.295 74.440 177.665 ;
        RECT 74.720 177.655 74.890 177.845 ;
        RECT 75.060 177.820 75.315 178.395 ;
        RECT 74.720 177.325 74.975 177.655 ;
        RECT 74.720 177.115 74.890 177.325 ;
        RECT 71.305 176.645 73.915 176.855 ;
        RECT 74.175 176.945 74.890 177.115 ;
        RECT 75.145 177.090 75.315 177.820 ;
        RECT 75.490 177.725 75.750 178.565 ;
        RECT 75.925 177.795 79.435 178.565 ;
        RECT 72.875 176.015 73.205 176.465 ;
        RECT 74.175 176.185 74.345 176.945 ;
        RECT 74.560 176.015 74.890 176.775 ;
        RECT 75.060 176.185 75.315 177.090 ;
        RECT 75.490 176.015 75.750 177.165 ;
        RECT 75.925 177.105 77.615 177.625 ;
        RECT 77.785 177.275 79.435 177.795 ;
        RECT 79.605 177.765 79.945 178.395 ;
        RECT 80.115 177.765 80.365 178.565 ;
        RECT 80.555 177.915 80.885 178.395 ;
        RECT 81.055 178.105 81.280 178.565 ;
        RECT 81.450 177.915 81.780 178.395 ;
        RECT 79.605 177.155 79.780 177.765 ;
        RECT 80.555 177.745 81.780 177.915 ;
        RECT 82.410 177.785 82.910 178.395 ;
        RECT 79.950 177.405 80.645 177.575 ;
        RECT 80.475 177.155 80.645 177.405 ;
        RECT 80.820 177.375 81.240 177.575 ;
        RECT 81.410 177.375 81.740 177.575 ;
        RECT 81.910 177.375 82.240 177.575 ;
        RECT 82.410 177.155 82.580 177.785 ;
        RECT 83.285 177.765 83.625 178.395 ;
        RECT 83.795 177.765 84.045 178.565 ;
        RECT 84.235 177.915 84.565 178.395 ;
        RECT 84.735 178.105 84.960 178.565 ;
        RECT 85.130 177.915 85.460 178.395 ;
        RECT 82.765 177.325 83.115 177.575 ;
        RECT 83.285 177.155 83.460 177.765 ;
        RECT 84.235 177.745 85.460 177.915 ;
        RECT 86.090 177.785 86.590 178.395 ;
        RECT 86.965 177.795 88.635 178.565 ;
        RECT 88.805 177.840 89.095 178.565 ;
        RECT 89.355 177.915 89.525 178.395 ;
        RECT 89.705 178.085 89.945 178.565 ;
        RECT 90.195 177.915 90.365 178.395 ;
        RECT 90.535 178.085 90.865 178.565 ;
        RECT 91.035 177.915 91.205 178.395 ;
        RECT 83.630 177.405 84.325 177.575 ;
        RECT 84.155 177.155 84.325 177.405 ;
        RECT 84.500 177.375 84.920 177.575 ;
        RECT 85.090 177.375 85.420 177.575 ;
        RECT 85.590 177.375 85.920 177.575 ;
        RECT 86.090 177.155 86.260 177.785 ;
        RECT 86.445 177.325 86.795 177.575 ;
        RECT 75.925 176.015 79.435 177.105 ;
        RECT 79.605 176.185 79.945 177.155 ;
        RECT 80.115 176.015 80.285 177.155 ;
        RECT 80.475 176.985 82.910 177.155 ;
        RECT 80.555 176.015 80.805 176.815 ;
        RECT 81.450 176.185 81.780 176.985 ;
        RECT 82.080 176.015 82.410 176.815 ;
        RECT 82.580 176.185 82.910 176.985 ;
        RECT 83.285 176.185 83.625 177.155 ;
        RECT 83.795 176.015 83.965 177.155 ;
        RECT 84.155 176.985 86.590 177.155 ;
        RECT 84.235 176.015 84.485 176.815 ;
        RECT 85.130 176.185 85.460 176.985 ;
        RECT 85.760 176.015 86.090 176.815 ;
        RECT 86.260 176.185 86.590 176.985 ;
        RECT 86.965 177.105 87.715 177.625 ;
        RECT 87.885 177.275 88.635 177.795 ;
        RECT 89.355 177.745 89.990 177.915 ;
        RECT 90.195 177.745 91.205 177.915 ;
        RECT 91.375 177.765 91.705 178.565 ;
        RECT 92.025 177.795 95.535 178.565 ;
        RECT 89.820 177.575 89.990 177.745 ;
        RECT 90.705 177.715 91.205 177.745 ;
        RECT 89.270 177.335 89.650 177.575 ;
        RECT 89.820 177.405 90.320 177.575 ;
        RECT 86.965 176.015 88.635 177.105 ;
        RECT 88.805 176.015 89.095 177.180 ;
        RECT 89.820 177.165 89.990 177.405 ;
        RECT 90.710 177.205 91.205 177.715 ;
        RECT 89.275 176.995 89.990 177.165 ;
        RECT 90.195 177.035 91.205 177.205 ;
        RECT 89.275 176.185 89.605 176.995 ;
        RECT 89.775 176.015 90.015 176.815 ;
        RECT 90.195 176.185 90.365 177.035 ;
        RECT 90.535 176.015 90.865 176.815 ;
        RECT 91.035 176.185 91.205 177.035 ;
        RECT 91.375 176.015 91.705 177.165 ;
        RECT 92.025 177.105 93.715 177.625 ;
        RECT 93.885 177.275 95.535 177.795 ;
        RECT 95.910 177.785 96.410 178.395 ;
        RECT 95.705 177.325 96.055 177.575 ;
        RECT 96.240 177.155 96.410 177.785 ;
        RECT 97.040 177.915 97.370 178.395 ;
        RECT 97.540 178.105 97.765 178.565 ;
        RECT 97.935 177.915 98.265 178.395 ;
        RECT 97.040 177.745 98.265 177.915 ;
        RECT 98.455 177.765 98.705 178.565 ;
        RECT 98.875 177.765 99.215 178.395 ;
        RECT 96.580 177.375 96.910 177.575 ;
        RECT 97.080 177.375 97.410 177.575 ;
        RECT 97.580 177.375 98.000 177.575 ;
        RECT 98.175 177.405 98.870 177.575 ;
        RECT 98.175 177.155 98.345 177.405 ;
        RECT 99.040 177.155 99.215 177.765 ;
        RECT 92.025 176.015 95.535 177.105 ;
        RECT 95.910 176.985 98.345 177.155 ;
        RECT 95.910 176.185 96.240 176.985 ;
        RECT 96.410 176.015 96.740 176.815 ;
        RECT 97.040 176.185 97.370 176.985 ;
        RECT 98.015 176.015 98.265 176.815 ;
        RECT 98.535 176.015 98.705 177.155 ;
        RECT 98.875 176.185 99.215 177.155 ;
        RECT 99.390 177.855 99.645 178.385 ;
        RECT 99.815 178.105 100.120 178.565 ;
        RECT 100.365 178.185 101.435 178.355 ;
        RECT 99.390 177.205 99.600 177.855 ;
        RECT 100.365 177.830 100.685 178.185 ;
        RECT 100.360 177.655 100.685 177.830 ;
        RECT 99.770 177.355 100.685 177.655 ;
        RECT 100.855 177.615 101.095 178.015 ;
        RECT 101.265 177.955 101.435 178.185 ;
        RECT 101.605 178.125 101.795 178.565 ;
        RECT 101.965 178.115 102.915 178.395 ;
        RECT 103.135 178.205 103.485 178.375 ;
        RECT 101.265 177.785 101.795 177.955 ;
        RECT 99.770 177.325 100.510 177.355 ;
        RECT 99.390 176.325 99.645 177.205 ;
        RECT 99.815 176.015 100.120 177.155 ;
        RECT 100.340 176.735 100.510 177.325 ;
        RECT 100.855 177.245 101.395 177.615 ;
        RECT 101.575 177.505 101.795 177.785 ;
        RECT 101.965 177.335 102.135 178.115 ;
        RECT 101.730 177.165 102.135 177.335 ;
        RECT 102.305 177.325 102.655 177.945 ;
        RECT 101.730 177.075 101.900 177.165 ;
        RECT 102.825 177.155 103.035 177.945 ;
        RECT 100.680 176.905 101.900 177.075 ;
        RECT 102.360 176.995 103.035 177.155 ;
        RECT 100.340 176.565 101.140 176.735 ;
        RECT 100.460 176.015 100.790 176.395 ;
        RECT 100.970 176.275 101.140 176.565 ;
        RECT 101.730 176.525 101.900 176.905 ;
        RECT 102.070 176.985 103.035 176.995 ;
        RECT 103.225 177.815 103.485 178.205 ;
        RECT 103.695 178.105 104.025 178.565 ;
        RECT 104.900 178.175 105.755 178.345 ;
        RECT 105.960 178.175 106.455 178.345 ;
        RECT 106.625 178.205 106.955 178.565 ;
        RECT 103.225 177.125 103.395 177.815 ;
        RECT 103.565 177.465 103.735 177.645 ;
        RECT 103.905 177.635 104.695 177.885 ;
        RECT 104.900 177.465 105.070 178.175 ;
        RECT 105.240 177.665 105.595 177.885 ;
        RECT 103.565 177.295 105.255 177.465 ;
        RECT 102.070 176.695 102.530 176.985 ;
        RECT 103.225 176.955 104.725 177.125 ;
        RECT 103.225 176.815 103.395 176.955 ;
        RECT 102.835 176.645 103.395 176.815 ;
        RECT 101.310 176.015 101.560 176.475 ;
        RECT 101.730 176.185 102.600 176.525 ;
        RECT 102.835 176.185 103.005 176.645 ;
        RECT 103.840 176.615 104.915 176.785 ;
        RECT 103.175 176.015 103.545 176.475 ;
        RECT 103.840 176.275 104.010 176.615 ;
        RECT 104.180 176.015 104.510 176.445 ;
        RECT 104.745 176.275 104.915 176.615 ;
        RECT 105.085 176.515 105.255 177.295 ;
        RECT 105.425 177.075 105.595 177.665 ;
        RECT 105.765 177.265 106.115 177.885 ;
        RECT 105.425 176.685 105.890 177.075 ;
        RECT 106.285 176.815 106.455 178.175 ;
        RECT 106.625 176.985 107.085 178.035 ;
        RECT 106.060 176.645 106.455 176.815 ;
        RECT 106.060 176.515 106.230 176.645 ;
        RECT 105.085 176.185 105.765 176.515 ;
        RECT 105.980 176.185 106.230 176.515 ;
        RECT 106.400 176.015 106.650 176.475 ;
        RECT 106.820 176.200 107.145 176.985 ;
        RECT 107.315 176.185 107.485 178.305 ;
        RECT 107.655 178.185 107.985 178.565 ;
        RECT 108.155 178.015 108.410 178.305 ;
        RECT 107.660 177.845 108.410 178.015 ;
        RECT 107.660 176.855 107.890 177.845 ;
        RECT 108.585 177.765 108.925 178.395 ;
        RECT 109.095 177.765 109.345 178.565 ;
        RECT 109.535 177.915 109.865 178.395 ;
        RECT 110.035 178.105 110.260 178.565 ;
        RECT 110.430 177.915 110.760 178.395 ;
        RECT 108.060 177.025 108.410 177.675 ;
        RECT 108.585 177.155 108.760 177.765 ;
        RECT 109.535 177.745 110.760 177.915 ;
        RECT 111.390 177.785 111.890 178.395 ;
        RECT 112.725 177.795 114.395 178.565 ;
        RECT 114.565 177.840 114.855 178.565 ;
        RECT 115.025 177.795 118.535 178.565 ;
        RECT 108.930 177.405 109.625 177.575 ;
        RECT 109.455 177.155 109.625 177.405 ;
        RECT 109.800 177.375 110.220 177.575 ;
        RECT 110.390 177.375 110.720 177.575 ;
        RECT 110.890 177.375 111.220 177.575 ;
        RECT 111.390 177.155 111.560 177.785 ;
        RECT 111.745 177.325 112.095 177.575 ;
        RECT 107.660 176.685 108.410 176.855 ;
        RECT 107.655 176.015 107.985 176.515 ;
        RECT 108.155 176.185 108.410 176.685 ;
        RECT 108.585 176.185 108.925 177.155 ;
        RECT 109.095 176.015 109.265 177.155 ;
        RECT 109.455 176.985 111.890 177.155 ;
        RECT 109.535 176.015 109.785 176.815 ;
        RECT 110.430 176.185 110.760 176.985 ;
        RECT 111.060 176.015 111.390 176.815 ;
        RECT 111.560 176.185 111.890 176.985 ;
        RECT 112.725 177.105 113.475 177.625 ;
        RECT 113.645 177.275 114.395 177.795 ;
        RECT 112.725 176.015 114.395 177.105 ;
        RECT 114.565 176.015 114.855 177.180 ;
        RECT 115.025 177.105 116.715 177.625 ;
        RECT 116.885 177.275 118.535 177.795 ;
        RECT 118.745 177.745 118.975 178.565 ;
        RECT 119.145 177.765 119.475 178.395 ;
        RECT 118.725 177.325 119.055 177.575 ;
        RECT 119.225 177.165 119.475 177.765 ;
        RECT 119.645 177.745 119.855 178.565 ;
        RECT 120.545 177.795 122.215 178.565 ;
        RECT 122.475 178.015 122.645 178.395 ;
        RECT 122.825 178.185 123.155 178.565 ;
        RECT 122.475 177.845 123.140 178.015 ;
        RECT 123.335 177.890 123.595 178.395 ;
        RECT 115.025 176.015 118.535 177.105 ;
        RECT 118.745 176.015 118.975 177.155 ;
        RECT 119.145 176.185 119.475 177.165 ;
        RECT 119.645 176.015 119.855 177.155 ;
        RECT 120.545 177.105 121.295 177.625 ;
        RECT 121.465 177.275 122.215 177.795 ;
        RECT 122.405 177.295 122.735 177.665 ;
        RECT 122.970 177.590 123.140 177.845 ;
        RECT 122.970 177.260 123.255 177.590 ;
        RECT 122.970 177.115 123.140 177.260 ;
        RECT 120.545 176.015 122.215 177.105 ;
        RECT 122.475 176.945 123.140 177.115 ;
        RECT 123.425 177.090 123.595 177.890 ;
        RECT 123.765 177.795 126.355 178.565 ;
        RECT 126.525 177.815 127.735 178.565 ;
        RECT 122.475 176.185 122.645 176.945 ;
        RECT 122.825 176.015 123.155 176.775 ;
        RECT 123.325 176.185 123.595 177.090 ;
        RECT 123.765 177.105 124.975 177.625 ;
        RECT 125.145 177.275 126.355 177.795 ;
        RECT 126.525 177.105 127.045 177.645 ;
        RECT 127.215 177.275 127.735 177.815 ;
        RECT 123.765 176.015 126.355 177.105 ;
        RECT 126.525 176.015 127.735 177.105 ;
        RECT 20.640 175.845 127.820 176.015 ;
        RECT 20.725 174.755 21.935 175.845 ;
        RECT 20.725 174.045 21.245 174.585 ;
        RECT 21.415 174.215 21.935 174.755 ;
        RECT 22.565 174.755 24.235 175.845 ;
        RECT 22.565 174.235 23.315 174.755 ;
        RECT 24.405 174.680 24.695 175.845 ;
        RECT 24.870 175.175 25.125 175.675 ;
        RECT 25.295 175.345 25.625 175.845 ;
        RECT 24.870 175.005 25.620 175.175 ;
        RECT 23.485 174.065 24.235 174.585 ;
        RECT 24.870 174.185 25.220 174.835 ;
        RECT 20.725 173.295 21.935 174.045 ;
        RECT 22.565 173.295 24.235 174.065 ;
        RECT 24.405 173.295 24.695 174.020 ;
        RECT 25.390 174.015 25.620 175.005 ;
        RECT 24.870 173.845 25.620 174.015 ;
        RECT 24.870 173.555 25.125 173.845 ;
        RECT 25.295 173.295 25.625 173.675 ;
        RECT 25.795 173.555 25.965 175.675 ;
        RECT 26.135 174.875 26.460 175.660 ;
        RECT 26.630 175.385 26.880 175.845 ;
        RECT 27.050 175.345 27.300 175.675 ;
        RECT 27.515 175.345 28.195 175.675 ;
        RECT 27.050 175.215 27.220 175.345 ;
        RECT 26.825 175.045 27.220 175.215 ;
        RECT 26.195 173.825 26.655 174.875 ;
        RECT 26.825 173.685 26.995 175.045 ;
        RECT 27.390 174.785 27.855 175.175 ;
        RECT 27.165 173.975 27.515 174.595 ;
        RECT 27.685 174.195 27.855 174.785 ;
        RECT 28.025 174.565 28.195 175.345 ;
        RECT 28.365 175.245 28.535 175.585 ;
        RECT 28.770 175.415 29.100 175.845 ;
        RECT 29.270 175.245 29.440 175.585 ;
        RECT 29.735 175.385 30.105 175.845 ;
        RECT 28.365 175.075 29.440 175.245 ;
        RECT 30.275 175.215 30.445 175.675 ;
        RECT 30.680 175.335 31.550 175.675 ;
        RECT 31.720 175.385 31.970 175.845 ;
        RECT 29.885 175.045 30.445 175.215 ;
        RECT 29.885 174.905 30.055 175.045 ;
        RECT 28.555 174.735 30.055 174.905 ;
        RECT 30.750 174.875 31.210 175.165 ;
        RECT 28.025 174.395 29.715 174.565 ;
        RECT 27.685 173.975 28.040 174.195 ;
        RECT 28.210 173.685 28.380 174.395 ;
        RECT 28.585 173.975 29.375 174.225 ;
        RECT 29.545 174.215 29.715 174.395 ;
        RECT 29.885 174.045 30.055 174.735 ;
        RECT 26.325 173.295 26.655 173.655 ;
        RECT 26.825 173.515 27.320 173.685 ;
        RECT 27.525 173.515 28.380 173.685 ;
        RECT 29.255 173.295 29.585 173.755 ;
        RECT 29.795 173.655 30.055 174.045 ;
        RECT 30.245 174.865 31.210 174.875 ;
        RECT 31.380 174.955 31.550 175.335 ;
        RECT 32.140 175.295 32.310 175.585 ;
        RECT 32.490 175.465 32.820 175.845 ;
        RECT 32.140 175.125 32.940 175.295 ;
        RECT 30.245 174.705 30.920 174.865 ;
        RECT 31.380 174.785 32.600 174.955 ;
        RECT 30.245 173.915 30.455 174.705 ;
        RECT 31.380 174.695 31.550 174.785 ;
        RECT 30.625 173.915 30.975 174.535 ;
        RECT 31.145 174.525 31.550 174.695 ;
        RECT 31.145 173.745 31.315 174.525 ;
        RECT 31.485 174.075 31.705 174.355 ;
        RECT 31.885 174.245 32.425 174.615 ;
        RECT 32.770 174.535 32.940 175.125 ;
        RECT 33.160 174.705 33.465 175.845 ;
        RECT 33.635 174.655 33.890 175.535 ;
        RECT 32.770 174.505 33.510 174.535 ;
        RECT 31.485 173.905 32.015 174.075 ;
        RECT 29.795 173.485 30.145 173.655 ;
        RECT 30.365 173.465 31.315 173.745 ;
        RECT 31.485 173.295 31.675 173.735 ;
        RECT 31.845 173.675 32.015 173.905 ;
        RECT 32.185 173.845 32.425 174.245 ;
        RECT 32.595 174.205 33.510 174.505 ;
        RECT 32.595 174.030 32.920 174.205 ;
        RECT 32.595 173.675 32.915 174.030 ;
        RECT 33.680 174.005 33.890 174.655 ;
        RECT 34.525 174.755 36.195 175.845 ;
        RECT 34.525 174.235 35.275 174.755 ;
        RECT 36.365 174.705 36.705 175.675 ;
        RECT 36.875 174.705 37.045 175.845 ;
        RECT 37.315 175.045 37.565 175.845 ;
        RECT 38.210 174.875 38.540 175.675 ;
        RECT 38.840 175.045 39.170 175.845 ;
        RECT 39.340 174.875 39.670 175.675 ;
        RECT 37.235 174.705 39.670 174.875 ;
        RECT 40.250 174.875 40.580 175.675 ;
        RECT 40.750 175.045 41.080 175.845 ;
        RECT 41.380 174.875 41.710 175.675 ;
        RECT 42.355 175.045 42.605 175.845 ;
        RECT 40.250 174.705 42.685 174.875 ;
        RECT 42.875 174.705 43.045 175.845 ;
        RECT 43.215 174.705 43.555 175.675 ;
        RECT 44.650 175.410 49.995 175.845 ;
        RECT 35.445 174.065 36.195 174.585 ;
        RECT 31.845 173.505 32.915 173.675 ;
        RECT 33.160 173.295 33.465 173.755 ;
        RECT 33.635 173.475 33.890 174.005 ;
        RECT 34.525 173.295 36.195 174.065 ;
        RECT 36.365 174.145 36.540 174.705 ;
        RECT 37.235 174.455 37.405 174.705 ;
        RECT 36.710 174.285 37.405 174.455 ;
        RECT 37.580 174.285 38.000 174.485 ;
        RECT 38.170 174.285 38.500 174.485 ;
        RECT 38.670 174.285 39.000 174.485 ;
        RECT 36.365 174.095 36.595 174.145 ;
        RECT 36.365 173.465 36.705 174.095 ;
        RECT 36.875 173.295 37.125 174.095 ;
        RECT 37.315 173.945 38.540 174.115 ;
        RECT 37.315 173.465 37.645 173.945 ;
        RECT 37.815 173.295 38.040 173.755 ;
        RECT 38.210 173.465 38.540 173.945 ;
        RECT 39.170 174.075 39.340 174.705 ;
        RECT 39.525 174.285 39.875 174.535 ;
        RECT 40.045 174.285 40.395 174.535 ;
        RECT 40.580 174.075 40.750 174.705 ;
        RECT 40.920 174.285 41.250 174.485 ;
        RECT 41.420 174.285 41.750 174.485 ;
        RECT 41.920 174.285 42.340 174.485 ;
        RECT 42.515 174.455 42.685 174.705 ;
        RECT 42.515 174.285 43.210 174.455 ;
        RECT 39.170 173.465 39.670 174.075 ;
        RECT 40.250 173.465 40.750 174.075 ;
        RECT 41.380 173.945 42.605 174.115 ;
        RECT 43.380 174.095 43.555 174.705 ;
        RECT 46.240 174.160 46.590 175.410 ;
        RECT 50.165 174.680 50.455 175.845 ;
        RECT 50.625 174.755 53.215 175.845 ;
        RECT 41.380 173.465 41.710 173.945 ;
        RECT 41.880 173.295 42.105 173.755 ;
        RECT 42.275 173.465 42.605 173.945 ;
        RECT 42.795 173.295 43.045 174.095 ;
        RECT 43.215 173.465 43.555 174.095 ;
        RECT 48.070 173.840 48.410 174.670 ;
        RECT 50.625 174.235 51.835 174.755 ;
        RECT 53.385 174.705 53.725 175.675 ;
        RECT 53.895 174.705 54.065 175.845 ;
        RECT 54.335 175.045 54.585 175.845 ;
        RECT 55.230 174.875 55.560 175.675 ;
        RECT 55.860 175.045 56.190 175.845 ;
        RECT 56.360 174.875 56.690 175.675 ;
        RECT 54.255 174.705 56.690 174.875 ;
        RECT 57.065 174.705 57.405 175.675 ;
        RECT 57.575 174.705 57.745 175.845 ;
        RECT 58.015 175.045 58.265 175.845 ;
        RECT 58.910 174.875 59.240 175.675 ;
        RECT 59.540 175.045 59.870 175.845 ;
        RECT 60.040 174.875 60.370 175.675 ;
        RECT 57.935 174.705 60.370 174.875 ;
        RECT 60.805 174.705 61.015 175.845 ;
        RECT 52.005 174.065 53.215 174.585 ;
        RECT 44.650 173.295 49.995 173.840 ;
        RECT 50.165 173.295 50.455 174.020 ;
        RECT 50.625 173.295 53.215 174.065 ;
        RECT 53.385 174.145 53.560 174.705 ;
        RECT 54.255 174.455 54.425 174.705 ;
        RECT 53.730 174.285 54.425 174.455 ;
        RECT 54.600 174.285 55.020 174.485 ;
        RECT 55.190 174.285 55.520 174.485 ;
        RECT 55.690 174.285 56.020 174.485 ;
        RECT 53.385 174.095 53.615 174.145 ;
        RECT 53.385 173.465 53.725 174.095 ;
        RECT 53.895 173.295 54.145 174.095 ;
        RECT 54.335 173.945 55.560 174.115 ;
        RECT 54.335 173.465 54.665 173.945 ;
        RECT 54.835 173.295 55.060 173.755 ;
        RECT 55.230 173.465 55.560 173.945 ;
        RECT 56.190 174.075 56.360 174.705 ;
        RECT 56.545 174.285 56.895 174.535 ;
        RECT 57.065 174.095 57.240 174.705 ;
        RECT 57.935 174.455 58.105 174.705 ;
        RECT 57.410 174.285 58.105 174.455 ;
        RECT 58.280 174.285 58.700 174.485 ;
        RECT 58.870 174.285 59.200 174.485 ;
        RECT 59.370 174.285 59.700 174.485 ;
        RECT 56.190 173.465 56.690 174.075 ;
        RECT 57.065 173.465 57.405 174.095 ;
        RECT 57.575 173.295 57.825 174.095 ;
        RECT 58.015 173.945 59.240 174.115 ;
        RECT 58.015 173.465 58.345 173.945 ;
        RECT 58.515 173.295 58.740 173.755 ;
        RECT 58.910 173.465 59.240 173.945 ;
        RECT 59.870 174.075 60.040 174.705 ;
        RECT 61.185 174.695 61.515 175.675 ;
        RECT 61.685 174.705 61.915 175.845 ;
        RECT 62.590 175.410 67.935 175.845 ;
        RECT 60.225 174.285 60.575 174.535 ;
        RECT 59.870 173.465 60.370 174.075 ;
        RECT 60.805 173.295 61.015 174.115 ;
        RECT 61.185 174.095 61.435 174.695 ;
        RECT 61.605 174.285 61.935 174.535 ;
        RECT 64.180 174.160 64.530 175.410 ;
        RECT 68.110 174.695 68.370 175.845 ;
        RECT 68.545 174.770 68.800 175.675 ;
        RECT 68.970 175.085 69.300 175.845 ;
        RECT 69.515 174.915 69.685 175.675 ;
        RECT 61.185 173.465 61.515 174.095 ;
        RECT 61.685 173.295 61.915 174.115 ;
        RECT 66.010 173.840 66.350 174.670 ;
        RECT 62.590 173.295 67.935 173.840 ;
        RECT 68.110 173.295 68.370 174.135 ;
        RECT 68.545 174.040 68.715 174.770 ;
        RECT 68.970 174.745 69.685 174.915 ;
        RECT 70.015 174.905 70.275 175.675 ;
        RECT 70.445 175.075 70.775 175.845 ;
        RECT 70.945 175.505 72.065 175.675 ;
        RECT 70.945 174.905 71.135 175.505 ;
        RECT 68.970 174.535 69.140 174.745 ;
        RECT 70.015 174.735 71.135 174.905 ;
        RECT 71.305 174.920 71.635 175.335 ;
        RECT 71.805 175.310 72.065 175.505 ;
        RECT 72.295 175.125 72.625 175.845 ;
        RECT 72.795 174.920 72.985 175.675 ;
        RECT 73.155 175.125 73.485 175.845 ;
        RECT 73.655 174.920 73.915 175.675 ;
        RECT 74.085 175.385 74.345 175.845 ;
        RECT 71.305 174.750 73.915 174.920 ;
        RECT 68.885 174.205 69.140 174.535 ;
        RECT 68.545 173.465 68.800 174.040 ;
        RECT 68.970 174.015 69.140 174.205 ;
        RECT 69.420 174.195 69.775 174.565 ;
        RECT 70.005 174.455 70.900 174.505 ;
        RECT 70.005 174.285 70.955 174.455 ;
        RECT 71.125 174.285 72.095 174.565 ;
        RECT 72.555 174.285 73.415 174.575 ;
        RECT 68.970 173.845 69.685 174.015 ;
        RECT 70.005 173.975 70.345 174.285 ;
        RECT 68.970 173.295 69.300 173.675 ;
        RECT 69.515 173.465 69.685 173.845 ;
        RECT 70.515 173.845 73.055 174.055 ;
        RECT 70.515 173.725 70.705 173.845 ;
        RECT 73.225 173.675 73.415 174.100 ;
        RECT 73.585 173.880 73.915 174.750 ;
        RECT 74.085 174.205 74.375 175.180 ;
        RECT 74.605 174.705 74.815 175.845 ;
        RECT 74.985 174.695 75.315 175.675 ;
        RECT 75.485 174.705 75.715 175.845 ;
        RECT 72.295 173.655 73.415 173.675 ;
        RECT 70.015 173.295 70.345 173.655 ;
        RECT 70.875 173.295 71.205 173.655 ;
        RECT 71.735 173.295 72.065 173.655 ;
        RECT 72.295 173.465 74.365 173.655 ;
        RECT 74.605 173.295 74.815 174.115 ;
        RECT 74.985 174.095 75.235 174.695 ;
        RECT 75.925 174.680 76.215 175.845 ;
        RECT 75.405 174.285 75.735 174.535 ;
        RECT 74.985 173.465 75.315 174.095 ;
        RECT 75.485 173.295 75.715 174.115 ;
        RECT 76.385 174.035 76.645 175.660 ;
        RECT 78.395 175.395 78.725 175.845 ;
        RECT 76.825 175.005 79.435 175.215 ;
        RECT 76.825 174.205 77.045 175.005 ;
        RECT 77.285 174.205 77.585 174.825 ;
        RECT 77.755 174.205 78.085 174.825 ;
        RECT 78.255 174.205 78.575 174.825 ;
        RECT 78.745 174.205 79.095 174.825 ;
        RECT 79.265 174.035 79.435 175.005 ;
        RECT 80.065 174.755 81.735 175.845 ;
        RECT 80.065 174.235 80.815 174.755 ;
        RECT 81.905 174.705 82.245 175.675 ;
        RECT 82.415 174.705 82.585 175.845 ;
        RECT 82.855 175.045 83.105 175.845 ;
        RECT 83.750 174.875 84.080 175.675 ;
        RECT 84.380 175.045 84.710 175.845 ;
        RECT 84.880 174.875 85.210 175.675 ;
        RECT 85.675 175.175 85.845 175.675 ;
        RECT 86.015 175.345 86.345 175.845 ;
        RECT 85.675 175.005 86.340 175.175 ;
        RECT 82.775 174.705 85.210 174.875 ;
        RECT 80.985 174.065 81.735 174.585 ;
        RECT 75.925 173.295 76.215 174.020 ;
        RECT 76.385 173.865 78.225 174.035 ;
        RECT 76.655 173.295 76.985 173.690 ;
        RECT 77.155 173.510 77.355 173.865 ;
        RECT 77.525 173.295 77.855 173.695 ;
        RECT 78.025 173.520 78.225 173.865 ;
        RECT 78.395 173.295 78.725 174.035 ;
        RECT 78.960 173.865 79.435 174.035 ;
        RECT 78.960 173.615 79.130 173.865 ;
        RECT 80.065 173.295 81.735 174.065 ;
        RECT 81.905 174.145 82.080 174.705 ;
        RECT 82.775 174.455 82.945 174.705 ;
        RECT 82.250 174.285 82.945 174.455 ;
        RECT 83.120 174.285 83.540 174.485 ;
        RECT 83.710 174.285 84.040 174.485 ;
        RECT 84.210 174.285 84.540 174.485 ;
        RECT 81.905 174.095 82.135 174.145 ;
        RECT 81.905 173.465 82.245 174.095 ;
        RECT 82.415 173.295 82.665 174.095 ;
        RECT 82.855 173.945 84.080 174.115 ;
        RECT 82.855 173.465 83.185 173.945 ;
        RECT 83.355 173.295 83.580 173.755 ;
        RECT 83.750 173.465 84.080 173.945 ;
        RECT 84.710 174.075 84.880 174.705 ;
        RECT 85.065 174.285 85.415 174.535 ;
        RECT 85.590 174.185 85.940 174.835 ;
        RECT 84.710 173.465 85.210 174.075 ;
        RECT 86.110 174.015 86.340 175.005 ;
        RECT 85.675 173.845 86.340 174.015 ;
        RECT 85.675 173.555 85.845 173.845 ;
        RECT 86.015 173.295 86.345 173.675 ;
        RECT 86.515 173.555 86.740 175.675 ;
        RECT 86.955 175.345 87.285 175.845 ;
        RECT 87.455 175.175 87.625 175.675 ;
        RECT 87.860 175.460 88.690 175.630 ;
        RECT 88.930 175.465 89.310 175.845 ;
        RECT 86.930 175.005 87.625 175.175 ;
        RECT 86.930 174.035 87.100 175.005 ;
        RECT 87.270 174.215 87.680 174.835 ;
        RECT 87.850 174.785 88.350 175.165 ;
        RECT 86.930 173.845 87.625 174.035 ;
        RECT 87.850 173.915 88.070 174.785 ;
        RECT 88.520 174.615 88.690 175.460 ;
        RECT 89.490 175.295 89.660 175.585 ;
        RECT 89.830 175.465 90.160 175.845 ;
        RECT 90.630 175.375 91.260 175.625 ;
        RECT 91.440 175.465 91.860 175.845 ;
        RECT 91.090 175.295 91.260 175.375 ;
        RECT 92.060 175.295 92.300 175.585 ;
        RECT 88.860 175.045 90.230 175.295 ;
        RECT 88.860 174.785 89.110 175.045 ;
        RECT 89.620 174.615 89.870 174.775 ;
        RECT 88.520 174.445 89.870 174.615 ;
        RECT 88.520 174.405 88.940 174.445 ;
        RECT 88.250 173.855 88.600 174.225 ;
        RECT 86.955 173.295 87.285 173.675 ;
        RECT 87.455 173.515 87.625 173.845 ;
        RECT 88.770 173.675 88.940 174.405 ;
        RECT 90.040 174.275 90.230 175.045 ;
        RECT 89.110 173.945 89.520 174.275 ;
        RECT 89.810 173.935 90.230 174.275 ;
        RECT 90.400 174.865 90.920 175.175 ;
        RECT 91.090 175.125 92.300 175.295 ;
        RECT 92.530 175.155 92.860 175.845 ;
        RECT 90.400 174.105 90.570 174.865 ;
        RECT 90.740 174.275 90.920 174.685 ;
        RECT 91.090 174.615 91.260 175.125 ;
        RECT 93.030 174.975 93.200 175.585 ;
        RECT 93.470 175.125 93.800 175.635 ;
        RECT 93.030 174.955 93.350 174.975 ;
        RECT 91.430 174.785 93.350 174.955 ;
        RECT 91.090 174.445 92.990 174.615 ;
        RECT 91.320 174.105 91.650 174.225 ;
        RECT 90.400 173.935 91.650 174.105 ;
        RECT 87.925 173.475 88.940 173.675 ;
        RECT 89.110 173.295 89.520 173.735 ;
        RECT 89.810 173.505 90.060 173.935 ;
        RECT 90.260 173.295 90.580 173.755 ;
        RECT 91.820 173.685 91.990 174.445 ;
        RECT 92.660 174.385 92.990 174.445 ;
        RECT 92.180 174.215 92.510 174.275 ;
        RECT 92.180 173.945 92.840 174.215 ;
        RECT 93.160 173.890 93.350 174.785 ;
        RECT 91.140 173.515 91.990 173.685 ;
        RECT 92.190 173.295 92.850 173.775 ;
        RECT 93.030 173.560 93.350 173.890 ;
        RECT 93.550 174.535 93.800 175.125 ;
        RECT 93.980 175.045 94.265 175.845 ;
        RECT 94.445 174.865 94.700 175.535 ;
        RECT 93.550 174.205 94.350 174.535 ;
        RECT 93.550 173.555 93.800 174.205 ;
        RECT 94.520 174.145 94.700 174.865 ;
        RECT 95.705 174.755 97.375 175.845 ;
        RECT 97.545 175.085 98.060 175.495 ;
        RECT 98.295 175.085 98.465 175.845 ;
        RECT 98.635 175.505 100.665 175.675 ;
        RECT 95.705 174.235 96.455 174.755 ;
        RECT 94.520 174.005 94.785 174.145 ;
        RECT 96.625 174.065 97.375 174.585 ;
        RECT 97.545 174.275 97.885 175.085 ;
        RECT 98.635 174.840 98.805 175.505 ;
        RECT 99.200 175.165 100.325 175.335 ;
        RECT 98.055 174.650 98.805 174.840 ;
        RECT 98.975 174.825 99.985 174.995 ;
        RECT 97.545 174.105 98.775 174.275 ;
        RECT 94.445 173.975 94.785 174.005 ;
        RECT 93.980 173.295 94.265 173.755 ;
        RECT 94.445 173.475 94.700 173.975 ;
        RECT 95.705 173.295 97.375 174.065 ;
        RECT 97.820 173.500 98.065 174.105 ;
        RECT 98.285 173.295 98.795 173.830 ;
        RECT 98.975 173.465 99.165 174.825 ;
        RECT 99.335 174.485 99.610 174.625 ;
        RECT 99.335 174.315 99.615 174.485 ;
        RECT 99.335 173.465 99.610 174.315 ;
        RECT 99.815 174.025 99.985 174.825 ;
        RECT 100.155 174.035 100.325 175.165 ;
        RECT 100.495 174.535 100.665 175.505 ;
        RECT 100.835 174.705 101.005 175.845 ;
        RECT 101.175 174.705 101.510 175.675 ;
        RECT 100.495 174.205 100.690 174.535 ;
        RECT 100.915 174.205 101.170 174.535 ;
        RECT 100.915 174.035 101.085 174.205 ;
        RECT 101.340 174.035 101.510 174.705 ;
        RECT 101.685 174.680 101.975 175.845 ;
        RECT 102.605 174.755 104.275 175.845 ;
        RECT 104.535 174.915 104.705 175.675 ;
        RECT 104.885 175.085 105.215 175.845 ;
        RECT 102.605 174.235 103.355 174.755 ;
        RECT 104.535 174.745 105.200 174.915 ;
        RECT 105.385 174.770 105.655 175.675 ;
        RECT 105.030 174.600 105.200 174.745 ;
        RECT 103.525 174.065 104.275 174.585 ;
        RECT 104.465 174.195 104.795 174.565 ;
        RECT 105.030 174.270 105.315 174.600 ;
        RECT 100.155 173.865 101.085 174.035 ;
        RECT 100.155 173.830 100.330 173.865 ;
        RECT 99.800 173.465 100.330 173.830 ;
        RECT 100.755 173.295 101.085 173.695 ;
        RECT 101.255 173.465 101.510 174.035 ;
        RECT 101.685 173.295 101.975 174.020 ;
        RECT 102.605 173.295 104.275 174.065 ;
        RECT 105.030 174.015 105.200 174.270 ;
        RECT 104.535 173.845 105.200 174.015 ;
        RECT 105.485 173.970 105.655 174.770 ;
        RECT 106.285 174.755 107.955 175.845 ;
        RECT 108.330 174.875 108.660 175.675 ;
        RECT 108.830 175.045 109.160 175.845 ;
        RECT 109.460 174.875 109.790 175.675 ;
        RECT 110.435 175.045 110.685 175.845 ;
        RECT 106.285 174.235 107.035 174.755 ;
        RECT 108.330 174.705 110.765 174.875 ;
        RECT 110.955 174.705 111.125 175.845 ;
        RECT 111.295 174.705 111.635 175.675 ;
        RECT 107.205 174.065 107.955 174.585 ;
        RECT 108.125 174.285 108.475 174.535 ;
        RECT 108.660 174.075 108.830 174.705 ;
        RECT 109.000 174.285 109.330 174.485 ;
        RECT 109.500 174.285 109.830 174.485 ;
        RECT 110.000 174.285 110.420 174.485 ;
        RECT 110.595 174.455 110.765 174.705 ;
        RECT 110.595 174.285 111.290 174.455 ;
        RECT 111.460 174.145 111.635 174.705 ;
        RECT 104.535 173.465 104.705 173.845 ;
        RECT 104.885 173.295 105.215 173.675 ;
        RECT 105.395 173.465 105.655 173.970 ;
        RECT 106.285 173.295 107.955 174.065 ;
        RECT 108.330 173.465 108.830 174.075 ;
        RECT 109.460 173.945 110.685 174.115 ;
        RECT 111.405 174.095 111.635 174.145 ;
        RECT 111.805 175.085 112.320 175.495 ;
        RECT 112.555 175.085 112.725 175.845 ;
        RECT 112.895 175.505 114.925 175.675 ;
        RECT 111.805 174.275 112.145 175.085 ;
        RECT 112.895 174.840 113.065 175.505 ;
        RECT 113.460 175.165 114.585 175.335 ;
        RECT 112.315 174.650 113.065 174.840 ;
        RECT 113.235 174.825 114.245 174.995 ;
        RECT 111.805 174.105 113.035 174.275 ;
        RECT 109.460 173.465 109.790 173.945 ;
        RECT 109.960 173.295 110.185 173.755 ;
        RECT 110.355 173.465 110.685 173.945 ;
        RECT 110.875 173.295 111.125 174.095 ;
        RECT 111.295 173.465 111.635 174.095 ;
        RECT 112.080 173.500 112.325 174.105 ;
        RECT 112.545 173.295 113.055 173.830 ;
        RECT 113.235 173.465 113.425 174.825 ;
        RECT 113.595 174.485 113.870 174.625 ;
        RECT 113.595 174.315 113.875 174.485 ;
        RECT 113.595 173.465 113.870 174.315 ;
        RECT 114.075 174.025 114.245 174.825 ;
        RECT 114.415 174.035 114.585 175.165 ;
        RECT 114.755 174.535 114.925 175.505 ;
        RECT 115.095 174.705 115.265 175.845 ;
        RECT 115.435 174.705 115.770 175.675 ;
        RECT 114.755 174.205 114.950 174.535 ;
        RECT 115.175 174.205 115.430 174.535 ;
        RECT 115.175 174.035 115.345 174.205 ;
        RECT 115.600 174.035 115.770 174.705 ;
        RECT 114.415 173.865 115.345 174.035 ;
        RECT 114.415 173.830 114.590 173.865 ;
        RECT 114.060 173.465 114.590 173.830 ;
        RECT 115.015 173.295 115.345 173.695 ;
        RECT 115.515 173.465 115.770 174.035 ;
        RECT 115.950 174.655 116.205 175.535 ;
        RECT 116.375 174.705 116.680 175.845 ;
        RECT 117.020 175.465 117.350 175.845 ;
        RECT 117.530 175.295 117.700 175.585 ;
        RECT 117.870 175.385 118.120 175.845 ;
        RECT 116.900 175.125 117.700 175.295 ;
        RECT 118.290 175.335 119.160 175.675 ;
        RECT 115.950 174.005 116.160 174.655 ;
        RECT 116.900 174.535 117.070 175.125 ;
        RECT 118.290 174.955 118.460 175.335 ;
        RECT 119.395 175.215 119.565 175.675 ;
        RECT 119.735 175.385 120.105 175.845 ;
        RECT 120.400 175.245 120.570 175.585 ;
        RECT 120.740 175.415 121.070 175.845 ;
        RECT 121.305 175.245 121.475 175.585 ;
        RECT 117.240 174.785 118.460 174.955 ;
        RECT 118.630 174.875 119.090 175.165 ;
        RECT 119.395 175.045 119.955 175.215 ;
        RECT 120.400 175.075 121.475 175.245 ;
        RECT 121.645 175.345 122.325 175.675 ;
        RECT 122.540 175.345 122.790 175.675 ;
        RECT 122.960 175.385 123.210 175.845 ;
        RECT 119.785 174.905 119.955 175.045 ;
        RECT 118.630 174.865 119.595 174.875 ;
        RECT 118.290 174.695 118.460 174.785 ;
        RECT 118.920 174.705 119.595 174.865 ;
        RECT 116.330 174.505 117.070 174.535 ;
        RECT 116.330 174.205 117.245 174.505 ;
        RECT 116.920 174.030 117.245 174.205 ;
        RECT 115.950 173.475 116.205 174.005 ;
        RECT 116.375 173.295 116.680 173.755 ;
        RECT 116.925 173.675 117.245 174.030 ;
        RECT 117.415 174.245 117.955 174.615 ;
        RECT 118.290 174.525 118.695 174.695 ;
        RECT 117.415 173.845 117.655 174.245 ;
        RECT 118.135 174.075 118.355 174.355 ;
        RECT 117.825 173.905 118.355 174.075 ;
        RECT 117.825 173.675 117.995 173.905 ;
        RECT 118.525 173.745 118.695 174.525 ;
        RECT 118.865 173.915 119.215 174.535 ;
        RECT 119.385 173.915 119.595 174.705 ;
        RECT 119.785 174.735 121.285 174.905 ;
        RECT 119.785 174.045 119.955 174.735 ;
        RECT 121.645 174.565 121.815 175.345 ;
        RECT 122.620 175.215 122.790 175.345 ;
        RECT 120.125 174.395 121.815 174.565 ;
        RECT 121.985 174.785 122.450 175.175 ;
        RECT 122.620 175.045 123.015 175.215 ;
        RECT 120.125 174.215 120.295 174.395 ;
        RECT 116.925 173.505 117.995 173.675 ;
        RECT 118.165 173.295 118.355 173.735 ;
        RECT 118.525 173.465 119.475 173.745 ;
        RECT 119.785 173.655 120.045 174.045 ;
        RECT 120.465 173.975 121.255 174.225 ;
        RECT 119.695 173.485 120.045 173.655 ;
        RECT 120.255 173.295 120.585 173.755 ;
        RECT 121.460 173.685 121.630 174.395 ;
        RECT 121.985 174.195 122.155 174.785 ;
        RECT 121.800 173.975 122.155 174.195 ;
        RECT 122.325 173.975 122.675 174.595 ;
        RECT 122.845 173.685 123.015 175.045 ;
        RECT 123.380 174.875 123.705 175.660 ;
        RECT 123.185 173.825 123.645 174.875 ;
        RECT 121.460 173.515 122.315 173.685 ;
        RECT 122.520 173.515 123.015 173.685 ;
        RECT 123.185 173.295 123.515 173.655 ;
        RECT 123.875 173.555 124.045 175.675 ;
        RECT 124.215 175.345 124.545 175.845 ;
        RECT 124.715 175.175 124.970 175.675 ;
        RECT 124.220 175.005 124.970 175.175 ;
        RECT 124.220 174.015 124.450 175.005 ;
        RECT 124.620 174.185 124.970 174.835 ;
        RECT 125.145 174.755 126.355 175.845 ;
        RECT 126.525 174.755 127.735 175.845 ;
        RECT 125.145 174.215 125.665 174.755 ;
        RECT 125.835 174.045 126.355 174.585 ;
        RECT 126.525 174.215 127.045 174.755 ;
        RECT 127.215 174.045 127.735 174.585 ;
        RECT 124.220 173.845 124.970 174.015 ;
        RECT 124.215 173.295 124.545 173.675 ;
        RECT 124.715 173.555 124.970 173.845 ;
        RECT 125.145 173.295 126.355 174.045 ;
        RECT 126.525 173.295 127.735 174.045 ;
        RECT 20.640 173.125 127.820 173.295 ;
        RECT 20.725 172.375 21.935 173.125 ;
        RECT 20.725 171.835 21.245 172.375 ;
        RECT 22.105 172.355 23.775 173.125 ;
        RECT 21.415 171.665 21.935 172.205 ;
        RECT 20.725 170.575 21.935 171.665 ;
        RECT 22.105 171.665 22.855 172.185 ;
        RECT 23.025 171.835 23.775 172.355 ;
        RECT 24.005 172.305 24.215 173.125 ;
        RECT 24.385 172.325 24.715 172.955 ;
        RECT 24.385 171.725 24.635 172.325 ;
        RECT 24.885 172.305 25.115 173.125 ;
        RECT 25.365 172.305 25.595 173.125 ;
        RECT 25.765 172.325 26.095 172.955 ;
        RECT 24.805 171.885 25.135 172.135 ;
        RECT 25.345 171.885 25.675 172.135 ;
        RECT 25.845 171.725 26.095 172.325 ;
        RECT 26.265 172.305 26.475 173.125 ;
        RECT 26.710 172.415 26.965 172.945 ;
        RECT 27.135 172.665 27.440 173.125 ;
        RECT 27.685 172.745 28.755 172.915 ;
        RECT 22.105 170.575 23.775 171.665 ;
        RECT 24.005 170.575 24.215 171.715 ;
        RECT 24.385 170.745 24.715 171.725 ;
        RECT 24.885 170.575 25.115 171.715 ;
        RECT 25.365 170.575 25.595 171.715 ;
        RECT 25.765 170.745 26.095 171.725 ;
        RECT 26.710 171.765 26.920 172.415 ;
        RECT 27.685 172.390 28.005 172.745 ;
        RECT 27.680 172.215 28.005 172.390 ;
        RECT 27.090 171.915 28.005 172.215 ;
        RECT 28.175 172.175 28.415 172.575 ;
        RECT 28.585 172.515 28.755 172.745 ;
        RECT 28.925 172.685 29.115 173.125 ;
        RECT 29.285 172.675 30.235 172.955 ;
        RECT 30.455 172.765 30.805 172.935 ;
        RECT 28.585 172.345 29.115 172.515 ;
        RECT 27.090 171.885 27.830 171.915 ;
        RECT 26.265 170.575 26.475 171.715 ;
        RECT 26.710 170.885 26.965 171.765 ;
        RECT 27.135 170.575 27.440 171.715 ;
        RECT 27.660 171.295 27.830 171.885 ;
        RECT 28.175 171.805 28.715 172.175 ;
        RECT 28.895 172.065 29.115 172.345 ;
        RECT 29.285 171.895 29.455 172.675 ;
        RECT 29.050 171.725 29.455 171.895 ;
        RECT 29.625 171.885 29.975 172.505 ;
        RECT 29.050 171.635 29.220 171.725 ;
        RECT 30.145 171.715 30.355 172.505 ;
        RECT 28.000 171.465 29.220 171.635 ;
        RECT 29.680 171.555 30.355 171.715 ;
        RECT 27.660 171.125 28.460 171.295 ;
        RECT 27.780 170.575 28.110 170.955 ;
        RECT 28.290 170.835 28.460 171.125 ;
        RECT 29.050 171.085 29.220 171.465 ;
        RECT 29.390 171.545 30.355 171.555 ;
        RECT 30.545 172.375 30.805 172.765 ;
        RECT 31.015 172.665 31.345 173.125 ;
        RECT 32.220 172.735 33.075 172.905 ;
        RECT 33.280 172.735 33.775 172.905 ;
        RECT 33.945 172.765 34.275 173.125 ;
        RECT 30.545 171.685 30.715 172.375 ;
        RECT 30.885 172.025 31.055 172.205 ;
        RECT 31.225 172.195 32.015 172.445 ;
        RECT 32.220 172.025 32.390 172.735 ;
        RECT 32.560 172.225 32.915 172.445 ;
        RECT 30.885 171.855 32.575 172.025 ;
        RECT 29.390 171.255 29.850 171.545 ;
        RECT 30.545 171.515 32.045 171.685 ;
        RECT 30.545 171.375 30.715 171.515 ;
        RECT 30.155 171.205 30.715 171.375 ;
        RECT 28.630 170.575 28.880 171.035 ;
        RECT 29.050 170.745 29.920 171.085 ;
        RECT 30.155 170.745 30.325 171.205 ;
        RECT 31.160 171.175 32.235 171.345 ;
        RECT 30.495 170.575 30.865 171.035 ;
        RECT 31.160 170.835 31.330 171.175 ;
        RECT 31.500 170.575 31.830 171.005 ;
        RECT 32.065 170.835 32.235 171.175 ;
        RECT 32.405 171.075 32.575 171.855 ;
        RECT 32.745 171.635 32.915 172.225 ;
        RECT 33.085 171.825 33.435 172.445 ;
        RECT 32.745 171.245 33.210 171.635 ;
        RECT 33.605 171.375 33.775 172.735 ;
        RECT 33.945 171.545 34.405 172.595 ;
        RECT 33.380 171.205 33.775 171.375 ;
        RECT 33.380 171.075 33.550 171.205 ;
        RECT 32.405 170.745 33.085 171.075 ;
        RECT 33.300 170.745 33.550 171.075 ;
        RECT 33.720 170.575 33.970 171.035 ;
        RECT 34.140 170.760 34.465 171.545 ;
        RECT 34.635 170.745 34.805 172.865 ;
        RECT 34.975 172.745 35.305 173.125 ;
        RECT 35.475 172.575 35.730 172.865 ;
        RECT 34.980 172.405 35.730 172.575 ;
        RECT 34.980 171.415 35.210 172.405 ;
        RECT 35.905 172.375 37.115 173.125 ;
        RECT 37.285 172.400 37.575 173.125 ;
        RECT 35.380 171.585 35.730 172.235 ;
        RECT 35.905 171.665 36.425 172.205 ;
        RECT 36.595 171.835 37.115 172.375 ;
        RECT 38.665 172.355 42.175 173.125 ;
        RECT 34.980 171.245 35.730 171.415 ;
        RECT 34.975 170.575 35.305 171.075 ;
        RECT 35.475 170.745 35.730 171.245 ;
        RECT 35.905 170.575 37.115 171.665 ;
        RECT 37.285 170.575 37.575 171.740 ;
        RECT 38.665 171.665 40.355 172.185 ;
        RECT 40.525 171.835 42.175 172.355 ;
        RECT 42.385 172.305 42.615 173.125 ;
        RECT 42.785 172.325 43.115 172.955 ;
        RECT 42.365 171.885 42.695 172.135 ;
        RECT 42.865 171.725 43.115 172.325 ;
        RECT 43.285 172.305 43.495 173.125 ;
        RECT 43.725 172.325 44.065 172.955 ;
        RECT 44.235 172.325 44.485 173.125 ;
        RECT 44.675 172.475 45.005 172.955 ;
        RECT 45.175 172.665 45.400 173.125 ;
        RECT 45.570 172.475 45.900 172.955 ;
        RECT 38.665 170.575 42.175 171.665 ;
        RECT 42.385 170.575 42.615 171.715 ;
        RECT 42.785 170.745 43.115 171.725 ;
        RECT 43.725 171.715 43.900 172.325 ;
        RECT 44.675 172.305 45.900 172.475 ;
        RECT 46.530 172.345 47.030 172.955 ;
        RECT 47.405 172.615 47.710 173.125 ;
        RECT 44.070 171.965 44.765 172.135 ;
        RECT 44.595 171.715 44.765 171.965 ;
        RECT 44.940 171.935 45.360 172.135 ;
        RECT 45.530 171.935 45.860 172.135 ;
        RECT 46.030 171.935 46.360 172.135 ;
        RECT 46.530 171.715 46.700 172.345 ;
        RECT 46.885 171.885 47.235 172.135 ;
        RECT 47.405 171.885 47.720 172.445 ;
        RECT 47.890 172.135 48.140 172.945 ;
        RECT 48.310 172.600 48.570 173.125 ;
        RECT 48.750 172.135 49.000 172.945 ;
        RECT 49.170 172.565 49.430 173.125 ;
        RECT 49.600 172.475 49.860 172.930 ;
        RECT 50.030 172.645 50.290 173.125 ;
        RECT 50.460 172.475 50.720 172.930 ;
        RECT 50.890 172.645 51.150 173.125 ;
        RECT 51.320 172.475 51.580 172.930 ;
        RECT 51.750 172.645 51.995 173.125 ;
        RECT 52.165 172.475 52.440 172.930 ;
        RECT 52.610 172.645 52.855 173.125 ;
        RECT 53.025 172.475 53.285 172.930 ;
        RECT 53.465 172.645 53.715 173.125 ;
        RECT 53.885 172.475 54.145 172.930 ;
        RECT 54.325 172.645 54.575 173.125 ;
        RECT 54.745 172.475 55.005 172.930 ;
        RECT 55.185 172.645 55.445 173.125 ;
        RECT 55.615 172.475 55.875 172.930 ;
        RECT 56.045 172.645 56.345 173.125 ;
        RECT 57.530 172.580 62.875 173.125 ;
        RECT 49.600 172.305 56.345 172.475 ;
        RECT 47.890 171.885 55.010 172.135 ;
        RECT 43.285 170.575 43.495 171.715 ;
        RECT 43.725 170.745 44.065 171.715 ;
        RECT 44.235 170.575 44.405 171.715 ;
        RECT 44.595 171.545 47.030 171.715 ;
        RECT 44.675 170.575 44.925 171.375 ;
        RECT 45.570 170.745 45.900 171.545 ;
        RECT 46.200 170.575 46.530 171.375 ;
        RECT 46.700 170.745 47.030 171.545 ;
        RECT 47.415 170.575 47.710 171.385 ;
        RECT 47.890 170.745 48.135 171.885 ;
        RECT 48.310 170.575 48.570 171.385 ;
        RECT 48.750 170.750 49.000 171.885 ;
        RECT 55.180 171.765 56.345 172.305 ;
        RECT 55.180 171.715 56.375 171.765 ;
        RECT 49.600 171.595 56.375 171.715 ;
        RECT 49.600 171.490 56.345 171.595 ;
        RECT 49.600 171.475 55.005 171.490 ;
        RECT 49.170 170.580 49.430 171.375 ;
        RECT 49.600 170.750 49.860 171.475 ;
        RECT 50.030 170.580 50.290 171.305 ;
        RECT 50.460 170.750 50.720 171.475 ;
        RECT 50.890 170.580 51.150 171.305 ;
        RECT 51.320 170.750 51.580 171.475 ;
        RECT 51.750 170.580 52.010 171.305 ;
        RECT 52.180 170.750 52.440 171.475 ;
        RECT 52.610 170.580 52.855 171.305 ;
        RECT 53.025 170.750 53.285 171.475 ;
        RECT 53.470 170.580 53.715 171.305 ;
        RECT 53.885 170.750 54.145 171.475 ;
        RECT 54.330 170.580 54.575 171.305 ;
        RECT 54.745 170.750 55.005 171.475 ;
        RECT 55.190 170.580 55.445 171.305 ;
        RECT 55.615 170.750 55.905 171.490 ;
        RECT 49.170 170.575 55.445 170.580 ;
        RECT 56.075 170.575 56.345 171.320 ;
        RECT 59.120 171.010 59.470 172.260 ;
        RECT 60.950 171.750 61.290 172.580 ;
        RECT 63.045 172.400 63.335 173.125 ;
        RECT 63.970 172.580 69.315 173.125 ;
        RECT 57.530 170.575 62.875 171.010 ;
        RECT 63.045 170.575 63.335 171.740 ;
        RECT 65.560 171.010 65.910 172.260 ;
        RECT 67.390 171.750 67.730 172.580 ;
        RECT 69.790 172.555 69.960 172.805 ;
        RECT 69.485 172.385 69.960 172.555 ;
        RECT 70.195 172.385 70.525 173.125 ;
        RECT 70.695 172.555 70.895 172.900 ;
        RECT 71.065 172.725 71.395 173.125 ;
        RECT 71.565 172.555 71.765 172.910 ;
        RECT 71.935 172.730 72.265 173.125 ;
        RECT 72.705 172.625 72.965 172.955 ;
        RECT 73.275 172.745 73.605 173.125 ;
        RECT 73.785 172.785 75.265 172.955 ;
        RECT 70.695 172.385 72.535 172.555 ;
        RECT 69.485 171.415 69.655 172.385 ;
        RECT 69.825 171.595 70.175 172.215 ;
        RECT 70.345 171.595 70.665 172.215 ;
        RECT 70.835 171.595 71.165 172.215 ;
        RECT 71.335 171.595 71.635 172.215 ;
        RECT 71.875 171.415 72.095 172.215 ;
        RECT 69.485 171.205 72.095 171.415 ;
        RECT 63.970 170.575 69.315 171.010 ;
        RECT 70.195 170.575 70.525 171.025 ;
        RECT 72.275 170.760 72.535 172.385 ;
        RECT 72.705 171.925 72.875 172.625 ;
        RECT 73.785 172.455 74.185 172.785 ;
        RECT 73.225 172.265 73.435 172.445 ;
        RECT 73.225 172.095 73.845 172.265 ;
        RECT 74.015 171.975 74.185 172.455 ;
        RECT 74.375 172.285 74.925 172.615 ;
        RECT 72.705 171.755 73.835 171.925 ;
        RECT 74.015 171.805 74.585 171.975 ;
        RECT 72.705 171.075 72.875 171.755 ;
        RECT 73.665 171.635 73.835 171.755 ;
        RECT 73.045 171.255 73.395 171.585 ;
        RECT 73.665 171.465 74.245 171.635 ;
        RECT 74.415 171.295 74.585 171.805 ;
        RECT 73.845 171.125 74.585 171.295 ;
        RECT 74.755 171.295 74.925 172.285 ;
        RECT 75.095 171.885 75.265 172.785 ;
        RECT 75.515 172.215 75.700 172.795 ;
        RECT 75.970 172.215 76.165 172.790 ;
        RECT 76.375 172.745 76.705 173.125 ;
        RECT 75.515 171.885 75.745 172.215 ;
        RECT 75.970 171.885 76.225 172.215 ;
        RECT 75.515 171.575 75.700 171.885 ;
        RECT 75.970 171.575 76.165 171.885 ;
        RECT 76.535 171.295 76.705 172.215 ;
        RECT 74.755 171.125 76.705 171.295 ;
        RECT 72.705 170.745 72.965 171.075 ;
        RECT 73.275 170.575 73.605 170.955 ;
        RECT 73.845 170.745 74.035 171.125 ;
        RECT 74.285 170.575 74.615 170.955 ;
        RECT 74.825 170.745 74.995 171.125 ;
        RECT 75.190 170.575 75.520 170.955 ;
        RECT 75.780 170.745 75.950 171.125 ;
        RECT 76.375 170.575 76.705 170.955 ;
        RECT 76.875 170.745 77.135 172.955 ;
        RECT 77.770 172.580 83.115 173.125 ;
        RECT 79.360 171.010 79.710 172.260 ;
        RECT 81.190 171.750 81.530 172.580 ;
        RECT 83.375 172.575 83.545 172.955 ;
        RECT 83.725 172.745 84.055 173.125 ;
        RECT 83.375 172.405 84.040 172.575 ;
        RECT 84.235 172.450 84.495 172.955 ;
        RECT 83.305 171.855 83.635 172.225 ;
        RECT 83.870 172.150 84.040 172.405 ;
        RECT 83.870 171.820 84.155 172.150 ;
        RECT 83.870 171.675 84.040 171.820 ;
        RECT 83.375 171.505 84.040 171.675 ;
        RECT 84.325 171.650 84.495 172.450 ;
        RECT 77.770 170.575 83.115 171.010 ;
        RECT 83.375 170.745 83.545 171.505 ;
        RECT 83.725 170.575 84.055 171.335 ;
        RECT 84.225 170.745 84.495 171.650 ;
        RECT 84.670 172.385 84.925 172.955 ;
        RECT 85.095 172.725 85.425 173.125 ;
        RECT 85.850 172.590 86.380 172.955 ;
        RECT 85.850 172.555 86.025 172.590 ;
        RECT 85.095 172.385 86.025 172.555 ;
        RECT 86.570 172.445 86.845 172.955 ;
        RECT 84.670 171.715 84.840 172.385 ;
        RECT 85.095 172.215 85.265 172.385 ;
        RECT 85.010 171.885 85.265 172.215 ;
        RECT 85.490 171.885 85.685 172.215 ;
        RECT 84.670 170.745 85.005 171.715 ;
        RECT 85.175 170.575 85.345 171.715 ;
        RECT 85.515 170.915 85.685 171.885 ;
        RECT 85.855 171.255 86.025 172.385 ;
        RECT 86.195 171.595 86.365 172.395 ;
        RECT 86.565 172.275 86.845 172.445 ;
        RECT 86.570 171.795 86.845 172.275 ;
        RECT 87.015 171.595 87.205 172.955 ;
        RECT 87.385 172.590 87.895 173.125 ;
        RECT 88.115 172.315 88.360 172.920 ;
        RECT 88.805 172.400 89.095 173.125 ;
        RECT 87.405 172.145 88.635 172.315 ;
        RECT 90.245 172.305 90.455 173.125 ;
        RECT 90.625 172.325 90.955 172.955 ;
        RECT 86.195 171.425 87.205 171.595 ;
        RECT 87.375 171.580 88.125 171.770 ;
        RECT 85.855 171.085 86.980 171.255 ;
        RECT 87.375 170.915 87.545 171.580 ;
        RECT 88.295 171.335 88.635 172.145 ;
        RECT 85.515 170.745 87.545 170.915 ;
        RECT 87.715 170.575 87.885 171.335 ;
        RECT 88.120 170.925 88.635 171.335 ;
        RECT 88.805 170.575 89.095 171.740 ;
        RECT 90.625 171.725 90.875 172.325 ;
        RECT 91.125 172.305 91.355 173.125 ;
        RECT 91.565 172.355 93.235 173.125 ;
        RECT 91.045 171.885 91.375 172.135 ;
        RECT 90.245 170.575 90.455 171.715 ;
        RECT 90.625 170.745 90.955 171.725 ;
        RECT 91.125 170.575 91.355 171.715 ;
        RECT 91.565 171.665 92.315 172.185 ;
        RECT 92.485 171.835 93.235 172.355 ;
        RECT 93.465 172.305 93.675 173.125 ;
        RECT 93.845 172.325 94.175 172.955 ;
        RECT 93.845 171.725 94.095 172.325 ;
        RECT 94.345 172.305 94.575 173.125 ;
        RECT 95.245 172.355 98.755 173.125 ;
        RECT 98.925 172.615 99.230 173.125 ;
        RECT 94.265 171.885 94.595 172.135 ;
        RECT 91.565 170.575 93.235 171.665 ;
        RECT 93.465 170.575 93.675 171.715 ;
        RECT 93.845 170.745 94.175 171.725 ;
        RECT 94.345 170.575 94.575 171.715 ;
        RECT 95.245 171.665 96.935 172.185 ;
        RECT 97.105 171.835 98.755 172.355 ;
        RECT 98.925 171.885 99.240 172.445 ;
        RECT 99.410 172.135 99.660 172.945 ;
        RECT 99.830 172.600 100.090 173.125 ;
        RECT 100.270 172.135 100.520 172.945 ;
        RECT 100.690 172.565 100.950 173.125 ;
        RECT 101.120 172.475 101.380 172.930 ;
        RECT 101.550 172.645 101.810 173.125 ;
        RECT 101.980 172.475 102.240 172.930 ;
        RECT 102.410 172.645 102.670 173.125 ;
        RECT 102.840 172.475 103.100 172.930 ;
        RECT 103.270 172.645 103.515 173.125 ;
        RECT 103.685 172.475 103.960 172.930 ;
        RECT 104.130 172.645 104.375 173.125 ;
        RECT 104.545 172.475 104.805 172.930 ;
        RECT 104.985 172.645 105.235 173.125 ;
        RECT 105.405 172.475 105.665 172.930 ;
        RECT 105.845 172.645 106.095 173.125 ;
        RECT 106.265 172.475 106.525 172.930 ;
        RECT 106.705 172.645 106.965 173.125 ;
        RECT 107.135 172.475 107.395 172.930 ;
        RECT 107.565 172.645 107.865 173.125 ;
        RECT 109.050 172.580 114.395 173.125 ;
        RECT 101.120 172.445 107.865 172.475 ;
        RECT 101.120 172.305 107.895 172.445 ;
        RECT 106.700 172.275 107.895 172.305 ;
        RECT 99.410 171.885 106.530 172.135 ;
        RECT 95.245 170.575 98.755 171.665 ;
        RECT 98.935 170.575 99.230 171.385 ;
        RECT 99.410 170.745 99.655 171.885 ;
        RECT 99.830 170.575 100.090 171.385 ;
        RECT 100.270 170.750 100.520 171.885 ;
        RECT 106.700 171.715 107.865 172.275 ;
        RECT 101.120 171.490 107.865 171.715 ;
        RECT 101.120 171.475 106.525 171.490 ;
        RECT 100.690 170.580 100.950 171.375 ;
        RECT 101.120 170.750 101.380 171.475 ;
        RECT 101.550 170.580 101.810 171.305 ;
        RECT 101.980 170.750 102.240 171.475 ;
        RECT 102.410 170.580 102.670 171.305 ;
        RECT 102.840 170.750 103.100 171.475 ;
        RECT 103.270 170.580 103.530 171.305 ;
        RECT 103.700 170.750 103.960 171.475 ;
        RECT 104.130 170.580 104.375 171.305 ;
        RECT 104.545 170.750 104.805 171.475 ;
        RECT 104.990 170.580 105.235 171.305 ;
        RECT 105.405 170.750 105.665 171.475 ;
        RECT 105.850 170.580 106.095 171.305 ;
        RECT 106.265 170.750 106.525 171.475 ;
        RECT 106.710 170.580 106.965 171.305 ;
        RECT 107.135 170.750 107.425 171.490 ;
        RECT 100.690 170.575 106.965 170.580 ;
        RECT 107.595 170.575 107.865 171.320 ;
        RECT 110.640 171.010 110.990 172.260 ;
        RECT 112.470 171.750 112.810 172.580 ;
        RECT 114.565 172.400 114.855 173.125 ;
        RECT 116.220 172.315 116.465 172.920 ;
        RECT 116.685 172.590 117.195 173.125 ;
        RECT 115.945 172.145 117.175 172.315 ;
        RECT 109.050 170.575 114.395 171.010 ;
        RECT 114.565 170.575 114.855 171.740 ;
        RECT 115.945 171.335 116.285 172.145 ;
        RECT 116.455 171.580 117.205 171.770 ;
        RECT 115.945 170.925 116.460 171.335 ;
        RECT 116.695 170.575 116.865 171.335 ;
        RECT 117.035 170.915 117.205 171.580 ;
        RECT 117.375 171.595 117.565 172.955 ;
        RECT 117.735 172.445 118.010 172.955 ;
        RECT 118.200 172.590 118.730 172.955 ;
        RECT 119.155 172.725 119.485 173.125 ;
        RECT 118.555 172.555 118.730 172.590 ;
        RECT 117.735 172.275 118.015 172.445 ;
        RECT 117.735 171.795 118.010 172.275 ;
        RECT 118.215 171.595 118.385 172.395 ;
        RECT 117.375 171.425 118.385 171.595 ;
        RECT 118.555 172.385 119.485 172.555 ;
        RECT 119.655 172.385 119.910 172.955 ;
        RECT 120.635 172.575 120.805 172.955 ;
        RECT 120.985 172.745 121.315 173.125 ;
        RECT 120.635 172.405 121.300 172.575 ;
        RECT 121.495 172.450 121.755 172.955 ;
        RECT 121.930 172.725 122.265 173.125 ;
        RECT 122.435 172.555 122.640 172.955 ;
        RECT 122.850 172.645 123.125 173.125 ;
        RECT 123.335 172.625 123.595 172.955 ;
        RECT 118.555 171.255 118.725 172.385 ;
        RECT 119.315 172.215 119.485 172.385 ;
        RECT 117.600 171.085 118.725 171.255 ;
        RECT 118.895 171.885 119.090 172.215 ;
        RECT 119.315 171.885 119.570 172.215 ;
        RECT 118.895 170.915 119.065 171.885 ;
        RECT 119.740 171.715 119.910 172.385 ;
        RECT 120.565 171.855 120.895 172.225 ;
        RECT 121.130 172.150 121.300 172.405 ;
        RECT 117.035 170.745 119.065 170.915 ;
        RECT 119.235 170.575 119.405 171.715 ;
        RECT 119.575 170.745 119.910 171.715 ;
        RECT 121.130 171.820 121.415 172.150 ;
        RECT 121.130 171.675 121.300 171.820 ;
        RECT 120.635 171.505 121.300 171.675 ;
        RECT 121.585 171.650 121.755 172.450 ;
        RECT 120.635 170.745 120.805 171.505 ;
        RECT 120.985 170.575 121.315 171.335 ;
        RECT 121.485 170.745 121.755 171.650 ;
        RECT 121.955 172.385 122.640 172.555 ;
        RECT 121.955 171.355 122.295 172.385 ;
        RECT 122.465 171.715 122.715 172.215 ;
        RECT 122.895 171.885 123.255 172.465 ;
        RECT 123.425 171.715 123.595 172.625 ;
        RECT 123.765 172.355 126.355 173.125 ;
        RECT 126.525 172.375 127.735 173.125 ;
        RECT 122.465 171.545 123.595 171.715 ;
        RECT 121.955 171.180 122.620 171.355 ;
        RECT 121.930 170.575 122.265 171.000 ;
        RECT 122.435 170.775 122.620 171.180 ;
        RECT 122.825 170.575 123.155 171.355 ;
        RECT 123.325 170.775 123.595 171.545 ;
        RECT 123.765 171.665 124.975 172.185 ;
        RECT 125.145 171.835 126.355 172.355 ;
        RECT 126.525 171.665 127.045 172.205 ;
        RECT 127.215 171.835 127.735 172.375 ;
        RECT 123.765 170.575 126.355 171.665 ;
        RECT 126.525 170.575 127.735 171.665 ;
        RECT 20.640 170.405 127.820 170.575 ;
        RECT 20.725 169.315 21.935 170.405 ;
        RECT 20.725 168.605 21.245 169.145 ;
        RECT 21.415 168.775 21.935 169.315 ;
        RECT 23.115 169.475 23.285 170.235 ;
        RECT 23.465 169.645 23.795 170.405 ;
        RECT 23.115 169.305 23.780 169.475 ;
        RECT 23.965 169.330 24.235 170.235 ;
        RECT 23.610 169.160 23.780 169.305 ;
        RECT 23.045 168.755 23.375 169.125 ;
        RECT 23.610 168.830 23.895 169.160 ;
        RECT 20.725 167.855 21.935 168.605 ;
        RECT 23.610 168.575 23.780 168.830 ;
        RECT 23.115 168.405 23.780 168.575 ;
        RECT 24.065 168.530 24.235 169.330 ;
        RECT 24.405 169.240 24.695 170.405 ;
        RECT 24.955 169.660 25.225 170.405 ;
        RECT 25.855 170.400 32.130 170.405 ;
        RECT 25.395 169.490 25.685 170.230 ;
        RECT 25.855 169.675 26.110 170.400 ;
        RECT 26.295 169.505 26.555 170.230 ;
        RECT 26.725 169.675 26.970 170.400 ;
        RECT 27.155 169.505 27.415 170.230 ;
        RECT 27.585 169.675 27.830 170.400 ;
        RECT 28.015 169.505 28.275 170.230 ;
        RECT 28.445 169.675 28.690 170.400 ;
        RECT 28.860 169.505 29.120 170.230 ;
        RECT 29.290 169.675 29.550 170.400 ;
        RECT 29.720 169.505 29.980 170.230 ;
        RECT 30.150 169.675 30.410 170.400 ;
        RECT 30.580 169.505 30.840 170.230 ;
        RECT 31.010 169.675 31.270 170.400 ;
        RECT 31.440 169.505 31.700 170.230 ;
        RECT 31.870 169.605 32.130 170.400 ;
        RECT 26.295 169.490 31.700 169.505 ;
        RECT 24.955 169.265 31.700 169.490 ;
        RECT 24.955 168.675 26.120 169.265 ;
        RECT 32.300 169.095 32.550 170.230 ;
        RECT 32.730 169.595 32.990 170.405 ;
        RECT 33.165 169.095 33.410 170.235 ;
        RECT 33.590 169.595 33.885 170.405 ;
        RECT 34.070 169.215 34.325 170.095 ;
        RECT 34.495 169.265 34.800 170.405 ;
        RECT 35.140 170.025 35.470 170.405 ;
        RECT 35.650 169.855 35.820 170.145 ;
        RECT 35.990 169.945 36.240 170.405 ;
        RECT 35.020 169.685 35.820 169.855 ;
        RECT 36.410 169.895 37.280 170.235 ;
        RECT 26.290 168.845 33.410 169.095 ;
        RECT 23.115 168.025 23.285 168.405 ;
        RECT 23.465 167.855 23.795 168.235 ;
        RECT 23.975 168.025 24.235 168.530 ;
        RECT 24.405 167.855 24.695 168.580 ;
        RECT 24.955 168.505 31.700 168.675 ;
        RECT 24.955 167.855 25.255 168.335 ;
        RECT 25.425 168.050 25.685 168.505 ;
        RECT 25.855 167.855 26.115 168.335 ;
        RECT 26.295 168.050 26.555 168.505 ;
        RECT 26.725 167.855 26.975 168.335 ;
        RECT 27.155 168.050 27.415 168.505 ;
        RECT 27.585 167.855 27.835 168.335 ;
        RECT 28.015 168.050 28.275 168.505 ;
        RECT 28.445 167.855 28.690 168.335 ;
        RECT 28.860 168.050 29.135 168.505 ;
        RECT 29.305 167.855 29.550 168.335 ;
        RECT 29.720 168.050 29.980 168.505 ;
        RECT 30.150 167.855 30.410 168.335 ;
        RECT 30.580 168.050 30.840 168.505 ;
        RECT 31.010 167.855 31.270 168.335 ;
        RECT 31.440 168.050 31.700 168.505 ;
        RECT 31.870 167.855 32.130 168.415 ;
        RECT 32.300 168.035 32.550 168.845 ;
        RECT 32.730 167.855 32.990 168.380 ;
        RECT 33.160 168.035 33.410 168.845 ;
        RECT 33.580 168.535 33.895 169.095 ;
        RECT 34.070 168.565 34.280 169.215 ;
        RECT 35.020 169.095 35.190 169.685 ;
        RECT 36.410 169.515 36.580 169.895 ;
        RECT 37.515 169.775 37.685 170.235 ;
        RECT 37.855 169.945 38.225 170.405 ;
        RECT 38.520 169.805 38.690 170.145 ;
        RECT 38.860 169.975 39.190 170.405 ;
        RECT 39.425 169.805 39.595 170.145 ;
        RECT 35.360 169.345 36.580 169.515 ;
        RECT 36.750 169.435 37.210 169.725 ;
        RECT 37.515 169.605 38.075 169.775 ;
        RECT 38.520 169.635 39.595 169.805 ;
        RECT 39.765 169.905 40.445 170.235 ;
        RECT 40.660 169.905 40.910 170.235 ;
        RECT 41.080 169.945 41.330 170.405 ;
        RECT 37.905 169.465 38.075 169.605 ;
        RECT 36.750 169.425 37.715 169.435 ;
        RECT 36.410 169.255 36.580 169.345 ;
        RECT 37.040 169.265 37.715 169.425 ;
        RECT 34.450 169.065 35.190 169.095 ;
        RECT 34.450 168.765 35.365 169.065 ;
        RECT 35.040 168.590 35.365 168.765 ;
        RECT 33.590 167.855 33.895 168.365 ;
        RECT 34.070 168.035 34.325 168.565 ;
        RECT 34.495 167.855 34.800 168.315 ;
        RECT 35.045 168.235 35.365 168.590 ;
        RECT 35.535 168.805 36.075 169.175 ;
        RECT 36.410 169.085 36.815 169.255 ;
        RECT 35.535 168.405 35.775 168.805 ;
        RECT 36.255 168.635 36.475 168.915 ;
        RECT 35.945 168.465 36.475 168.635 ;
        RECT 35.945 168.235 36.115 168.465 ;
        RECT 36.645 168.305 36.815 169.085 ;
        RECT 36.985 168.475 37.335 169.095 ;
        RECT 37.505 168.475 37.715 169.265 ;
        RECT 37.905 169.295 39.405 169.465 ;
        RECT 37.905 168.605 38.075 169.295 ;
        RECT 39.765 169.125 39.935 169.905 ;
        RECT 40.740 169.775 40.910 169.905 ;
        RECT 38.245 168.955 39.935 169.125 ;
        RECT 40.105 169.345 40.570 169.735 ;
        RECT 40.740 169.605 41.135 169.775 ;
        RECT 38.245 168.775 38.415 168.955 ;
        RECT 35.045 168.065 36.115 168.235 ;
        RECT 36.285 167.855 36.475 168.295 ;
        RECT 36.645 168.025 37.595 168.305 ;
        RECT 37.905 168.215 38.165 168.605 ;
        RECT 38.585 168.535 39.375 168.785 ;
        RECT 37.815 168.045 38.165 168.215 ;
        RECT 38.375 167.855 38.705 168.315 ;
        RECT 39.580 168.245 39.750 168.955 ;
        RECT 40.105 168.755 40.275 169.345 ;
        RECT 39.920 168.535 40.275 168.755 ;
        RECT 40.445 168.535 40.795 169.155 ;
        RECT 40.965 168.245 41.135 169.605 ;
        RECT 41.500 169.435 41.825 170.220 ;
        RECT 41.305 168.385 41.765 169.435 ;
        RECT 39.580 168.075 40.435 168.245 ;
        RECT 40.640 168.075 41.135 168.245 ;
        RECT 41.305 167.855 41.635 168.215 ;
        RECT 41.995 168.115 42.165 170.235 ;
        RECT 42.335 169.905 42.665 170.405 ;
        RECT 42.835 169.735 43.090 170.235 ;
        RECT 42.340 169.565 43.090 169.735 ;
        RECT 43.325 169.570 43.580 170.405 ;
        RECT 42.340 168.575 42.570 169.565 ;
        RECT 43.750 169.400 44.010 170.205 ;
        RECT 44.180 169.570 44.440 170.405 ;
        RECT 44.610 169.400 44.865 170.205 ;
        RECT 42.740 168.745 43.090 169.395 ;
        RECT 43.265 169.230 44.865 169.400 ;
        RECT 46.025 169.645 46.540 170.055 ;
        RECT 46.775 169.645 46.945 170.405 ;
        RECT 47.115 170.065 49.145 170.235 ;
        RECT 43.265 168.665 43.545 169.230 ;
        RECT 43.715 168.835 44.935 169.060 ;
        RECT 46.025 168.835 46.365 169.645 ;
        RECT 47.115 169.400 47.285 170.065 ;
        RECT 47.680 169.725 48.805 169.895 ;
        RECT 46.535 169.210 47.285 169.400 ;
        RECT 47.455 169.385 48.465 169.555 ;
        RECT 46.025 168.665 47.255 168.835 ;
        RECT 42.340 168.405 43.090 168.575 ;
        RECT 43.265 168.495 43.995 168.665 ;
        RECT 42.335 167.855 42.665 168.235 ;
        RECT 42.835 168.115 43.090 168.405 ;
        RECT 43.270 167.855 43.600 168.325 ;
        RECT 43.770 168.050 43.995 168.495 ;
        RECT 44.165 167.855 44.460 168.380 ;
        RECT 46.300 168.060 46.545 168.665 ;
        RECT 46.765 167.855 47.275 168.390 ;
        RECT 47.455 168.025 47.645 169.385 ;
        RECT 47.815 169.045 48.090 169.185 ;
        RECT 47.815 168.875 48.095 169.045 ;
        RECT 47.815 168.025 48.090 168.875 ;
        RECT 48.295 168.585 48.465 169.385 ;
        RECT 48.635 168.595 48.805 169.725 ;
        RECT 48.975 169.095 49.145 170.065 ;
        RECT 49.315 169.265 49.485 170.405 ;
        RECT 49.655 169.265 49.990 170.235 ;
        RECT 48.975 168.765 49.170 169.095 ;
        RECT 49.395 168.765 49.650 169.095 ;
        RECT 49.395 168.595 49.565 168.765 ;
        RECT 49.820 168.595 49.990 169.265 ;
        RECT 50.165 169.240 50.455 170.405 ;
        RECT 50.680 169.535 50.965 170.405 ;
        RECT 51.135 169.775 51.395 170.235 ;
        RECT 51.570 169.945 51.825 170.405 ;
        RECT 51.995 169.775 52.255 170.235 ;
        RECT 51.135 169.605 52.255 169.775 ;
        RECT 52.425 169.605 52.735 170.405 ;
        RECT 51.135 169.355 51.395 169.605 ;
        RECT 52.905 169.435 53.215 170.235 ;
        RECT 53.385 169.570 53.770 170.405 ;
        RECT 48.635 168.425 49.565 168.595 ;
        RECT 48.635 168.390 48.810 168.425 ;
        RECT 48.280 168.025 48.810 168.390 ;
        RECT 49.235 167.855 49.565 168.255 ;
        RECT 49.735 168.025 49.990 168.595 ;
        RECT 50.640 169.185 51.395 169.355 ;
        RECT 52.185 169.265 53.215 169.435 ;
        RECT 53.940 169.400 54.200 170.205 ;
        RECT 54.370 169.570 54.630 170.405 ;
        RECT 54.800 169.400 55.055 170.205 ;
        RECT 55.230 169.570 55.490 170.405 ;
        RECT 55.660 169.400 55.915 170.205 ;
        RECT 56.090 169.570 56.435 170.405 ;
        RECT 50.640 168.675 51.045 169.185 ;
        RECT 52.185 169.015 52.355 169.265 ;
        RECT 51.215 168.845 52.355 169.015 ;
        RECT 50.165 167.855 50.455 168.580 ;
        RECT 50.640 168.505 52.290 168.675 ;
        RECT 52.525 168.525 52.875 169.095 ;
        RECT 50.685 167.855 50.965 168.335 ;
        RECT 51.135 168.115 51.395 168.505 ;
        RECT 51.570 167.855 51.825 168.335 ;
        RECT 51.995 168.115 52.290 168.505 ;
        RECT 53.045 168.355 53.215 169.265 ;
        RECT 53.385 169.230 56.415 169.400 ;
        RECT 57.675 169.255 58.005 170.405 ;
        RECT 58.175 169.385 58.345 170.235 ;
        RECT 58.515 169.605 58.845 170.405 ;
        RECT 59.015 169.385 59.185 170.235 ;
        RECT 59.365 169.605 59.605 170.405 ;
        RECT 59.775 169.425 60.105 170.235 ;
        RECT 53.385 168.665 53.685 169.230 ;
        RECT 53.860 168.835 56.075 169.060 ;
        RECT 56.245 168.665 56.415 169.230 ;
        RECT 53.385 168.495 56.415 168.665 ;
        RECT 58.175 169.215 59.185 169.385 ;
        RECT 59.390 169.255 60.105 169.425 ;
        RECT 60.435 169.255 60.765 170.405 ;
        RECT 60.935 169.385 61.105 170.235 ;
        RECT 61.275 169.605 61.605 170.405 ;
        RECT 61.775 169.385 61.945 170.235 ;
        RECT 62.125 169.605 62.365 170.405 ;
        RECT 62.535 169.425 62.865 170.235 ;
        RECT 63.100 169.535 63.385 170.405 ;
        RECT 63.555 169.775 63.815 170.235 ;
        RECT 63.990 169.945 64.245 170.405 ;
        RECT 64.415 169.775 64.675 170.235 ;
        RECT 63.555 169.605 64.675 169.775 ;
        RECT 64.845 169.605 65.155 170.405 ;
        RECT 58.175 168.675 58.670 169.215 ;
        RECT 59.390 169.015 59.560 169.255 ;
        RECT 60.935 169.215 61.945 169.385 ;
        RECT 62.150 169.255 62.865 169.425 ;
        RECT 63.555 169.355 63.815 169.605 ;
        RECT 65.325 169.435 65.635 170.235 ;
        RECT 59.060 168.845 59.560 169.015 ;
        RECT 59.730 168.845 60.110 169.085 ;
        RECT 59.390 168.675 59.560 168.845 ;
        RECT 60.935 168.675 61.430 169.215 ;
        RECT 62.150 169.015 62.320 169.255 ;
        RECT 63.060 169.185 63.815 169.355 ;
        RECT 64.605 169.265 65.635 169.435 ;
        RECT 61.820 168.845 62.320 169.015 ;
        RECT 62.490 168.845 62.870 169.085 ;
        RECT 62.150 168.675 62.320 168.845 ;
        RECT 63.060 168.675 63.465 169.185 ;
        RECT 64.605 169.015 64.775 169.265 ;
        RECT 63.635 168.845 64.775 169.015 ;
        RECT 52.470 167.855 52.745 168.335 ;
        RECT 52.915 168.025 53.215 168.355 ;
        RECT 53.905 167.855 54.205 168.325 ;
        RECT 54.375 168.050 54.630 168.495 ;
        RECT 54.800 167.855 55.060 168.325 ;
        RECT 55.230 168.050 55.490 168.495 ;
        RECT 55.660 167.855 55.955 168.325 ;
        RECT 57.675 167.855 58.005 168.655 ;
        RECT 58.175 168.505 59.185 168.675 ;
        RECT 59.390 168.505 60.025 168.675 ;
        RECT 58.175 168.025 58.345 168.505 ;
        RECT 58.515 167.855 58.845 168.335 ;
        RECT 59.015 168.025 59.185 168.505 ;
        RECT 59.435 167.855 59.675 168.335 ;
        RECT 59.855 168.025 60.025 168.505 ;
        RECT 60.435 167.855 60.765 168.655 ;
        RECT 60.935 168.505 61.945 168.675 ;
        RECT 62.150 168.505 62.785 168.675 ;
        RECT 63.060 168.505 64.710 168.675 ;
        RECT 64.945 168.525 65.295 169.095 ;
        RECT 60.935 168.025 61.105 168.505 ;
        RECT 61.275 167.855 61.605 168.335 ;
        RECT 61.775 168.025 61.945 168.505 ;
        RECT 62.195 167.855 62.435 168.335 ;
        RECT 62.615 168.025 62.785 168.505 ;
        RECT 63.105 167.855 63.385 168.335 ;
        RECT 63.555 168.115 63.815 168.505 ;
        RECT 63.990 167.855 64.245 168.335 ;
        RECT 64.415 168.115 64.710 168.505 ;
        RECT 65.465 168.355 65.635 169.265 ;
        RECT 66.265 169.315 67.935 170.405 ;
        RECT 68.110 169.970 73.455 170.405 ;
        RECT 66.265 168.795 67.015 169.315 ;
        RECT 67.185 168.625 67.935 169.145 ;
        RECT 69.700 168.720 70.050 169.970 ;
        RECT 73.630 169.255 73.890 170.405 ;
        RECT 74.065 169.330 74.320 170.235 ;
        RECT 74.490 169.645 74.820 170.405 ;
        RECT 75.035 169.475 75.205 170.235 ;
        RECT 64.890 167.855 65.165 168.335 ;
        RECT 65.335 168.025 65.635 168.355 ;
        RECT 66.265 167.855 67.935 168.625 ;
        RECT 71.530 168.400 71.870 169.230 ;
        RECT 68.110 167.855 73.455 168.400 ;
        RECT 73.630 167.855 73.890 168.695 ;
        RECT 74.065 168.600 74.235 169.330 ;
        RECT 74.490 169.305 75.205 169.475 ;
        RECT 74.490 169.095 74.660 169.305 ;
        RECT 75.925 169.240 76.215 170.405 ;
        RECT 76.385 169.315 78.055 170.405 ;
        RECT 78.225 169.435 78.535 170.235 ;
        RECT 78.705 169.605 79.015 170.405 ;
        RECT 79.185 169.775 79.445 170.235 ;
        RECT 79.615 169.945 79.870 170.405 ;
        RECT 80.045 169.775 80.305 170.235 ;
        RECT 79.185 169.605 80.305 169.775 ;
        RECT 74.405 168.765 74.660 169.095 ;
        RECT 74.065 168.025 74.320 168.600 ;
        RECT 74.490 168.575 74.660 168.765 ;
        RECT 74.940 168.755 75.295 169.125 ;
        RECT 76.385 168.795 77.135 169.315 ;
        RECT 78.225 169.265 79.255 169.435 ;
        RECT 77.305 168.625 78.055 169.145 ;
        RECT 74.490 168.405 75.205 168.575 ;
        RECT 74.490 167.855 74.820 168.235 ;
        RECT 75.035 168.025 75.205 168.405 ;
        RECT 75.925 167.855 76.215 168.580 ;
        RECT 76.385 167.855 78.055 168.625 ;
        RECT 78.225 168.355 78.395 169.265 ;
        RECT 78.565 168.525 78.915 169.095 ;
        RECT 79.085 169.015 79.255 169.265 ;
        RECT 80.045 169.355 80.305 169.605 ;
        RECT 80.475 169.535 80.760 170.405 ;
        RECT 80.045 169.185 80.800 169.355 ;
        RECT 79.085 168.845 80.225 169.015 ;
        RECT 80.395 168.675 80.800 169.185 ;
        RECT 80.985 169.315 83.575 170.405 ;
        RECT 83.745 169.645 84.260 170.055 ;
        RECT 84.495 169.645 84.665 170.405 ;
        RECT 84.835 170.065 86.865 170.235 ;
        RECT 80.985 168.795 82.195 169.315 ;
        RECT 79.150 168.505 80.800 168.675 ;
        RECT 82.365 168.625 83.575 169.145 ;
        RECT 83.745 168.835 84.085 169.645 ;
        RECT 84.835 169.400 85.005 170.065 ;
        RECT 85.400 169.725 86.525 169.895 ;
        RECT 84.255 169.210 85.005 169.400 ;
        RECT 85.175 169.385 86.185 169.555 ;
        RECT 83.745 168.665 84.975 168.835 ;
        RECT 78.225 168.025 78.525 168.355 ;
        RECT 78.695 167.855 78.970 168.335 ;
        RECT 79.150 168.115 79.445 168.505 ;
        RECT 79.615 167.855 79.870 168.335 ;
        RECT 80.045 168.115 80.305 168.505 ;
        RECT 80.475 167.855 80.755 168.335 ;
        RECT 80.985 167.855 83.575 168.625 ;
        RECT 84.020 168.060 84.265 168.665 ;
        RECT 84.485 167.855 84.995 168.390 ;
        RECT 85.175 168.025 85.365 169.385 ;
        RECT 85.535 168.365 85.810 169.185 ;
        RECT 86.015 168.585 86.185 169.385 ;
        RECT 86.355 168.595 86.525 169.725 ;
        RECT 86.695 169.095 86.865 170.065 ;
        RECT 87.035 169.265 87.205 170.405 ;
        RECT 87.375 169.265 87.710 170.235 ;
        RECT 87.975 169.660 88.245 170.405 ;
        RECT 88.875 170.400 95.150 170.405 ;
        RECT 88.415 169.490 88.705 170.230 ;
        RECT 88.875 169.675 89.130 170.400 ;
        RECT 89.315 169.505 89.575 170.230 ;
        RECT 89.745 169.675 89.990 170.400 ;
        RECT 90.175 169.505 90.435 170.230 ;
        RECT 90.605 169.675 90.850 170.400 ;
        RECT 91.035 169.505 91.295 170.230 ;
        RECT 91.465 169.675 91.710 170.400 ;
        RECT 91.880 169.505 92.140 170.230 ;
        RECT 92.310 169.675 92.570 170.400 ;
        RECT 92.740 169.505 93.000 170.230 ;
        RECT 93.170 169.675 93.430 170.400 ;
        RECT 93.600 169.505 93.860 170.230 ;
        RECT 94.030 169.675 94.290 170.400 ;
        RECT 94.460 169.505 94.720 170.230 ;
        RECT 94.890 169.605 95.150 170.400 ;
        RECT 89.315 169.490 94.720 169.505 ;
        RECT 86.695 168.765 86.890 169.095 ;
        RECT 87.115 168.765 87.370 169.095 ;
        RECT 87.115 168.595 87.285 168.765 ;
        RECT 87.540 168.595 87.710 169.265 ;
        RECT 86.355 168.425 87.285 168.595 ;
        RECT 86.355 168.390 86.530 168.425 ;
        RECT 85.535 168.195 85.815 168.365 ;
        RECT 85.535 168.025 85.810 168.195 ;
        RECT 86.000 168.025 86.530 168.390 ;
        RECT 86.955 167.855 87.285 168.255 ;
        RECT 87.455 168.025 87.710 168.595 ;
        RECT 87.975 169.265 94.720 169.490 ;
        RECT 87.975 168.675 89.140 169.265 ;
        RECT 95.320 169.095 95.570 170.230 ;
        RECT 95.750 169.595 96.010 170.405 ;
        RECT 96.185 169.095 96.430 170.235 ;
        RECT 96.610 169.595 96.905 170.405 ;
        RECT 97.085 169.315 98.755 170.405 ;
        RECT 89.310 168.845 96.430 169.095 ;
        RECT 87.975 168.505 94.720 168.675 ;
        RECT 87.975 167.855 88.275 168.335 ;
        RECT 88.445 168.050 88.705 168.505 ;
        RECT 88.875 167.855 89.135 168.335 ;
        RECT 89.315 168.050 89.575 168.505 ;
        RECT 89.745 167.855 89.995 168.335 ;
        RECT 90.175 168.050 90.435 168.505 ;
        RECT 90.605 167.855 90.855 168.335 ;
        RECT 91.035 168.050 91.295 168.505 ;
        RECT 91.465 167.855 91.710 168.335 ;
        RECT 91.880 168.050 92.155 168.505 ;
        RECT 92.325 167.855 92.570 168.335 ;
        RECT 92.740 168.050 93.000 168.505 ;
        RECT 93.170 167.855 93.430 168.335 ;
        RECT 93.600 168.050 93.860 168.505 ;
        RECT 94.030 167.855 94.290 168.335 ;
        RECT 94.460 168.050 94.720 168.505 ;
        RECT 94.890 167.855 95.150 168.415 ;
        RECT 95.320 168.035 95.570 168.845 ;
        RECT 95.750 167.855 96.010 168.380 ;
        RECT 96.180 168.035 96.430 168.845 ;
        RECT 96.600 168.535 96.915 169.095 ;
        RECT 97.085 168.795 97.835 169.315 ;
        RECT 98.965 169.265 99.195 170.405 ;
        RECT 99.365 169.255 99.695 170.235 ;
        RECT 99.865 169.265 100.075 170.405 ;
        RECT 100.305 169.315 101.515 170.405 ;
        RECT 98.005 168.625 98.755 169.145 ;
        RECT 98.945 168.845 99.275 169.095 ;
        RECT 96.610 167.855 96.915 168.365 ;
        RECT 97.085 167.855 98.755 168.625 ;
        RECT 98.965 167.855 99.195 168.675 ;
        RECT 99.445 168.655 99.695 169.255 ;
        RECT 100.305 168.775 100.825 169.315 ;
        RECT 101.685 169.240 101.975 170.405 ;
        RECT 102.235 169.475 102.405 170.235 ;
        RECT 102.585 169.645 102.915 170.405 ;
        RECT 102.235 169.305 102.900 169.475 ;
        RECT 103.085 169.330 103.355 170.235 ;
        RECT 102.730 169.160 102.900 169.305 ;
        RECT 99.365 168.025 99.695 168.655 ;
        RECT 99.865 167.855 100.075 168.675 ;
        RECT 100.995 168.605 101.515 169.145 ;
        RECT 102.165 168.755 102.495 169.125 ;
        RECT 102.730 168.830 103.015 169.160 ;
        RECT 100.305 167.855 101.515 168.605 ;
        RECT 101.685 167.855 101.975 168.580 ;
        RECT 102.730 168.575 102.900 168.830 ;
        RECT 102.235 168.405 102.900 168.575 ;
        RECT 103.185 168.530 103.355 169.330 ;
        RECT 103.565 169.265 103.795 170.405 ;
        RECT 103.965 169.255 104.295 170.235 ;
        RECT 104.465 169.265 104.675 170.405 ;
        RECT 105.420 169.535 105.705 170.405 ;
        RECT 105.875 169.775 106.135 170.235 ;
        RECT 106.310 169.945 106.565 170.405 ;
        RECT 106.735 169.775 106.995 170.235 ;
        RECT 105.875 169.605 106.995 169.775 ;
        RECT 107.165 169.605 107.475 170.405 ;
        RECT 105.875 169.355 106.135 169.605 ;
        RECT 107.645 169.435 107.955 170.235 ;
        RECT 103.545 168.845 103.875 169.095 ;
        RECT 102.235 168.025 102.405 168.405 ;
        RECT 102.585 167.855 102.915 168.235 ;
        RECT 103.095 168.025 103.355 168.530 ;
        RECT 103.565 167.855 103.795 168.675 ;
        RECT 104.045 168.655 104.295 169.255 ;
        RECT 105.380 169.185 106.135 169.355 ;
        RECT 106.925 169.265 107.955 169.435 ;
        RECT 105.380 168.675 105.785 169.185 ;
        RECT 106.925 169.015 107.095 169.265 ;
        RECT 105.955 168.845 107.095 169.015 ;
        RECT 103.965 168.025 104.295 168.655 ;
        RECT 104.465 167.855 104.675 168.675 ;
        RECT 105.380 168.505 107.030 168.675 ;
        RECT 107.265 168.525 107.615 169.095 ;
        RECT 105.425 167.855 105.705 168.335 ;
        RECT 105.875 168.115 106.135 168.505 ;
        RECT 106.310 167.855 106.565 168.335 ;
        RECT 106.735 168.115 107.030 168.505 ;
        RECT 107.785 168.355 107.955 169.265 ;
        RECT 108.125 169.315 109.795 170.405 ;
        RECT 108.125 168.795 108.875 169.315 ;
        RECT 110.025 169.265 110.235 170.405 ;
        RECT 110.405 169.255 110.735 170.235 ;
        RECT 110.905 169.265 111.135 170.405 ;
        RECT 111.345 169.645 111.860 170.055 ;
        RECT 112.095 169.645 112.265 170.405 ;
        RECT 112.435 170.065 114.465 170.235 ;
        RECT 109.045 168.625 109.795 169.145 ;
        RECT 107.210 167.855 107.485 168.335 ;
        RECT 107.655 168.025 107.955 168.355 ;
        RECT 108.125 167.855 109.795 168.625 ;
        RECT 110.025 167.855 110.235 168.675 ;
        RECT 110.405 168.655 110.655 169.255 ;
        RECT 110.825 168.845 111.155 169.095 ;
        RECT 111.345 168.835 111.685 169.645 ;
        RECT 112.435 169.400 112.605 170.065 ;
        RECT 113.000 169.725 114.125 169.895 ;
        RECT 111.855 169.210 112.605 169.400 ;
        RECT 112.775 169.385 113.785 169.555 ;
        RECT 110.405 168.025 110.735 168.655 ;
        RECT 110.905 167.855 111.135 168.675 ;
        RECT 111.345 168.665 112.575 168.835 ;
        RECT 111.620 168.060 111.865 168.665 ;
        RECT 112.085 167.855 112.595 168.390 ;
        RECT 112.775 168.025 112.965 169.385 ;
        RECT 113.135 168.705 113.410 169.185 ;
        RECT 113.135 168.535 113.415 168.705 ;
        RECT 113.615 168.585 113.785 169.385 ;
        RECT 113.955 168.595 114.125 169.725 ;
        RECT 114.295 169.095 114.465 170.065 ;
        RECT 114.635 169.265 114.805 170.405 ;
        RECT 114.975 169.265 115.310 170.235 ;
        RECT 114.295 168.765 114.490 169.095 ;
        RECT 114.715 168.765 114.970 169.095 ;
        RECT 114.715 168.595 114.885 168.765 ;
        RECT 115.140 168.595 115.310 169.265 ;
        RECT 115.485 169.315 116.695 170.405 ;
        RECT 115.485 168.775 116.005 169.315 ;
        RECT 116.905 169.265 117.135 170.405 ;
        RECT 117.305 169.255 117.635 170.235 ;
        RECT 117.805 169.265 118.015 170.405 ;
        RECT 118.395 169.255 118.725 170.405 ;
        RECT 118.895 169.385 119.065 170.235 ;
        RECT 119.235 169.605 119.565 170.405 ;
        RECT 119.735 169.385 119.905 170.235 ;
        RECT 120.085 169.605 120.325 170.405 ;
        RECT 120.495 169.425 120.825 170.235 ;
        RECT 121.010 169.970 126.355 170.405 ;
        RECT 116.175 168.605 116.695 169.145 ;
        RECT 116.885 168.845 117.215 169.095 ;
        RECT 113.135 168.025 113.410 168.535 ;
        RECT 113.955 168.425 114.885 168.595 ;
        RECT 113.955 168.390 114.130 168.425 ;
        RECT 113.600 168.025 114.130 168.390 ;
        RECT 114.555 167.855 114.885 168.255 ;
        RECT 115.055 168.025 115.310 168.595 ;
        RECT 115.485 167.855 116.695 168.605 ;
        RECT 116.905 167.855 117.135 168.675 ;
        RECT 117.385 168.655 117.635 169.255 ;
        RECT 118.895 169.215 119.905 169.385 ;
        RECT 120.110 169.255 120.825 169.425 ;
        RECT 118.895 168.705 119.390 169.215 ;
        RECT 120.110 169.015 120.280 169.255 ;
        RECT 119.780 168.845 120.280 169.015 ;
        RECT 120.450 168.845 120.830 169.085 ;
        RECT 118.895 168.675 119.395 168.705 ;
        RECT 120.110 168.675 120.280 168.845 ;
        RECT 122.600 168.720 122.950 169.970 ;
        RECT 126.525 169.315 127.735 170.405 ;
        RECT 117.305 168.025 117.635 168.655 ;
        RECT 117.805 167.855 118.015 168.675 ;
        RECT 118.395 167.855 118.725 168.655 ;
        RECT 118.895 168.505 119.905 168.675 ;
        RECT 120.110 168.505 120.745 168.675 ;
        RECT 118.895 168.025 119.065 168.505 ;
        RECT 119.235 167.855 119.565 168.335 ;
        RECT 119.735 168.025 119.905 168.505 ;
        RECT 120.155 167.855 120.395 168.335 ;
        RECT 120.575 168.025 120.745 168.505 ;
        RECT 124.430 168.400 124.770 169.230 ;
        RECT 126.525 168.775 127.045 169.315 ;
        RECT 127.215 168.605 127.735 169.145 ;
        RECT 121.010 167.855 126.355 168.400 ;
        RECT 126.525 167.855 127.735 168.605 ;
        RECT 20.640 167.685 127.820 167.855 ;
        RECT 20.725 166.935 21.935 167.685 ;
        RECT 22.110 167.140 27.455 167.685 ;
        RECT 20.725 166.395 21.245 166.935 ;
        RECT 21.415 166.225 21.935 166.765 ;
        RECT 20.725 165.135 21.935 166.225 ;
        RECT 23.700 165.570 24.050 166.820 ;
        RECT 25.530 166.310 25.870 167.140 ;
        RECT 27.630 166.945 27.885 167.515 ;
        RECT 28.055 167.285 28.385 167.685 ;
        RECT 28.810 167.150 29.340 167.515 ;
        RECT 28.810 167.115 28.985 167.150 ;
        RECT 28.055 166.945 28.985 167.115 ;
        RECT 29.530 167.005 29.805 167.515 ;
        RECT 27.630 166.275 27.800 166.945 ;
        RECT 28.055 166.775 28.225 166.945 ;
        RECT 27.970 166.445 28.225 166.775 ;
        RECT 28.450 166.445 28.645 166.775 ;
        RECT 22.110 165.135 27.455 165.570 ;
        RECT 27.630 165.305 27.965 166.275 ;
        RECT 28.135 165.135 28.305 166.275 ;
        RECT 28.475 165.475 28.645 166.445 ;
        RECT 28.815 165.815 28.985 166.945 ;
        RECT 29.155 166.155 29.325 166.955 ;
        RECT 29.525 166.835 29.805 167.005 ;
        RECT 29.530 166.355 29.805 166.835 ;
        RECT 29.975 166.155 30.165 167.515 ;
        RECT 30.345 167.150 30.855 167.685 ;
        RECT 31.075 166.875 31.320 167.480 ;
        RECT 32.690 166.945 32.945 167.515 ;
        RECT 33.115 167.285 33.445 167.685 ;
        RECT 33.870 167.150 34.400 167.515 ;
        RECT 33.870 167.115 34.045 167.150 ;
        RECT 33.115 166.945 34.045 167.115 ;
        RECT 30.365 166.705 31.595 166.875 ;
        RECT 29.155 165.985 30.165 166.155 ;
        RECT 30.335 166.140 31.085 166.330 ;
        RECT 28.815 165.645 29.940 165.815 ;
        RECT 30.335 165.475 30.505 166.140 ;
        RECT 31.255 165.895 31.595 166.705 ;
        RECT 28.475 165.305 30.505 165.475 ;
        RECT 30.675 165.135 30.845 165.895 ;
        RECT 31.080 165.485 31.595 165.895 ;
        RECT 32.690 166.275 32.860 166.945 ;
        RECT 33.115 166.775 33.285 166.945 ;
        RECT 33.030 166.445 33.285 166.775 ;
        RECT 33.510 166.445 33.705 166.775 ;
        RECT 32.690 165.305 33.025 166.275 ;
        RECT 33.195 165.135 33.365 166.275 ;
        RECT 33.535 165.475 33.705 166.445 ;
        RECT 33.875 165.815 34.045 166.945 ;
        RECT 34.215 166.155 34.385 166.955 ;
        RECT 34.590 166.665 34.865 167.515 ;
        RECT 34.585 166.495 34.865 166.665 ;
        RECT 34.590 166.355 34.865 166.495 ;
        RECT 35.035 166.155 35.225 167.515 ;
        RECT 35.405 167.150 35.915 167.685 ;
        RECT 36.135 166.875 36.380 167.480 ;
        RECT 37.285 166.960 37.575 167.685 ;
        RECT 37.745 166.935 38.955 167.685 ;
        RECT 39.215 167.135 39.385 167.515 ;
        RECT 39.565 167.305 39.895 167.685 ;
        RECT 39.215 166.965 39.880 167.135 ;
        RECT 40.075 167.010 40.335 167.515 ;
        RECT 35.425 166.705 36.655 166.875 ;
        RECT 34.215 165.985 35.225 166.155 ;
        RECT 35.395 166.140 36.145 166.330 ;
        RECT 33.875 165.645 35.000 165.815 ;
        RECT 35.395 165.475 35.565 166.140 ;
        RECT 36.315 165.895 36.655 166.705 ;
        RECT 33.535 165.305 35.565 165.475 ;
        RECT 35.735 165.135 35.905 165.895 ;
        RECT 36.140 165.485 36.655 165.895 ;
        RECT 37.285 165.135 37.575 166.300 ;
        RECT 37.745 166.225 38.265 166.765 ;
        RECT 38.435 166.395 38.955 166.935 ;
        RECT 39.145 166.415 39.475 166.785 ;
        RECT 39.710 166.710 39.880 166.965 ;
        RECT 39.710 166.380 39.995 166.710 ;
        RECT 39.710 166.235 39.880 166.380 ;
        RECT 37.745 165.135 38.955 166.225 ;
        RECT 39.215 166.065 39.880 166.235 ;
        RECT 40.165 166.210 40.335 167.010 ;
        RECT 39.215 165.305 39.385 166.065 ;
        RECT 39.565 165.135 39.895 165.895 ;
        RECT 40.065 165.305 40.335 166.210 ;
        RECT 40.510 166.975 40.765 167.505 ;
        RECT 40.935 167.225 41.240 167.685 ;
        RECT 41.485 167.305 42.555 167.475 ;
        RECT 40.510 166.325 40.720 166.975 ;
        RECT 41.485 166.950 41.805 167.305 ;
        RECT 41.480 166.775 41.805 166.950 ;
        RECT 40.890 166.475 41.805 166.775 ;
        RECT 41.975 166.735 42.215 167.135 ;
        RECT 42.385 167.075 42.555 167.305 ;
        RECT 42.725 167.245 42.915 167.685 ;
        RECT 43.085 167.235 44.035 167.515 ;
        RECT 44.255 167.325 44.605 167.495 ;
        RECT 42.385 166.905 42.915 167.075 ;
        RECT 40.890 166.445 41.630 166.475 ;
        RECT 40.510 165.445 40.765 166.325 ;
        RECT 40.935 165.135 41.240 166.275 ;
        RECT 41.460 165.855 41.630 166.445 ;
        RECT 41.975 166.365 42.515 166.735 ;
        RECT 42.695 166.625 42.915 166.905 ;
        RECT 43.085 166.455 43.255 167.235 ;
        RECT 42.850 166.285 43.255 166.455 ;
        RECT 43.425 166.445 43.775 167.065 ;
        RECT 42.850 166.195 43.020 166.285 ;
        RECT 43.945 166.275 44.155 167.065 ;
        RECT 41.800 166.025 43.020 166.195 ;
        RECT 43.480 166.115 44.155 166.275 ;
        RECT 41.460 165.685 42.260 165.855 ;
        RECT 41.580 165.135 41.910 165.515 ;
        RECT 42.090 165.395 42.260 165.685 ;
        RECT 42.850 165.645 43.020 166.025 ;
        RECT 43.190 166.105 44.155 166.115 ;
        RECT 44.345 166.935 44.605 167.325 ;
        RECT 44.815 167.225 45.145 167.685 ;
        RECT 46.020 167.295 46.875 167.465 ;
        RECT 47.080 167.295 47.575 167.465 ;
        RECT 47.745 167.325 48.075 167.685 ;
        RECT 44.345 166.245 44.515 166.935 ;
        RECT 44.685 166.585 44.855 166.765 ;
        RECT 45.025 166.755 45.815 167.005 ;
        RECT 46.020 166.585 46.190 167.295 ;
        RECT 46.360 166.785 46.715 167.005 ;
        RECT 44.685 166.415 46.375 166.585 ;
        RECT 43.190 165.815 43.650 166.105 ;
        RECT 44.345 166.075 45.845 166.245 ;
        RECT 44.345 165.935 44.515 166.075 ;
        RECT 43.955 165.765 44.515 165.935 ;
        RECT 42.430 165.135 42.680 165.595 ;
        RECT 42.850 165.305 43.720 165.645 ;
        RECT 43.955 165.305 44.125 165.765 ;
        RECT 44.960 165.735 46.035 165.905 ;
        RECT 44.295 165.135 44.665 165.595 ;
        RECT 44.960 165.395 45.130 165.735 ;
        RECT 45.300 165.135 45.630 165.565 ;
        RECT 45.865 165.395 46.035 165.735 ;
        RECT 46.205 165.635 46.375 166.415 ;
        RECT 46.545 166.195 46.715 166.785 ;
        RECT 46.885 166.385 47.235 167.005 ;
        RECT 46.545 165.805 47.010 166.195 ;
        RECT 47.405 165.935 47.575 167.295 ;
        RECT 47.745 166.105 48.205 167.155 ;
        RECT 47.180 165.765 47.575 165.935 ;
        RECT 47.180 165.635 47.350 165.765 ;
        RECT 46.205 165.305 46.885 165.635 ;
        RECT 47.100 165.305 47.350 165.635 ;
        RECT 47.520 165.135 47.770 165.595 ;
        RECT 47.940 165.320 48.265 166.105 ;
        RECT 48.435 165.305 48.605 167.425 ;
        RECT 48.775 167.305 49.105 167.685 ;
        RECT 49.275 167.135 49.530 167.425 ;
        RECT 48.780 166.965 49.530 167.135 ;
        RECT 49.710 166.975 49.965 167.505 ;
        RECT 50.135 167.225 50.440 167.685 ;
        RECT 50.685 167.305 51.755 167.475 ;
        RECT 48.780 165.975 49.010 166.965 ;
        RECT 49.180 166.145 49.530 166.795 ;
        RECT 49.710 166.325 49.920 166.975 ;
        RECT 50.685 166.950 51.005 167.305 ;
        RECT 50.680 166.775 51.005 166.950 ;
        RECT 50.090 166.475 51.005 166.775 ;
        RECT 51.175 166.735 51.415 167.135 ;
        RECT 51.585 167.075 51.755 167.305 ;
        RECT 51.925 167.245 52.115 167.685 ;
        RECT 52.285 167.235 53.235 167.515 ;
        RECT 53.455 167.325 53.805 167.495 ;
        RECT 51.585 166.905 52.115 167.075 ;
        RECT 50.090 166.445 50.830 166.475 ;
        RECT 48.780 165.805 49.530 165.975 ;
        RECT 48.775 165.135 49.105 165.635 ;
        RECT 49.275 165.305 49.530 165.805 ;
        RECT 49.710 165.445 49.965 166.325 ;
        RECT 50.135 165.135 50.440 166.275 ;
        RECT 50.660 165.855 50.830 166.445 ;
        RECT 51.175 166.365 51.715 166.735 ;
        RECT 51.895 166.625 52.115 166.905 ;
        RECT 52.285 166.455 52.455 167.235 ;
        RECT 52.050 166.285 52.455 166.455 ;
        RECT 52.625 166.445 52.975 167.065 ;
        RECT 52.050 166.195 52.220 166.285 ;
        RECT 53.145 166.275 53.355 167.065 ;
        RECT 51.000 166.025 52.220 166.195 ;
        RECT 52.680 166.115 53.355 166.275 ;
        RECT 50.660 165.685 51.460 165.855 ;
        RECT 50.780 165.135 51.110 165.515 ;
        RECT 51.290 165.395 51.460 165.685 ;
        RECT 52.050 165.645 52.220 166.025 ;
        RECT 52.390 166.105 53.355 166.115 ;
        RECT 53.545 166.935 53.805 167.325 ;
        RECT 54.015 167.225 54.345 167.685 ;
        RECT 55.220 167.295 56.075 167.465 ;
        RECT 56.280 167.295 56.775 167.465 ;
        RECT 56.945 167.325 57.275 167.685 ;
        RECT 53.545 166.245 53.715 166.935 ;
        RECT 53.885 166.585 54.055 166.765 ;
        RECT 54.225 166.755 55.015 167.005 ;
        RECT 55.220 166.585 55.390 167.295 ;
        RECT 55.560 166.785 55.915 167.005 ;
        RECT 53.885 166.415 55.575 166.585 ;
        RECT 52.390 165.815 52.850 166.105 ;
        RECT 53.545 166.075 55.045 166.245 ;
        RECT 53.545 165.935 53.715 166.075 ;
        RECT 53.155 165.765 53.715 165.935 ;
        RECT 51.630 165.135 51.880 165.595 ;
        RECT 52.050 165.305 52.920 165.645 ;
        RECT 53.155 165.305 53.325 165.765 ;
        RECT 54.160 165.735 55.235 165.905 ;
        RECT 53.495 165.135 53.865 165.595 ;
        RECT 54.160 165.395 54.330 165.735 ;
        RECT 54.500 165.135 54.830 165.565 ;
        RECT 55.065 165.395 55.235 165.735 ;
        RECT 55.405 165.635 55.575 166.415 ;
        RECT 55.745 166.195 55.915 166.785 ;
        RECT 56.085 166.385 56.435 167.005 ;
        RECT 55.745 165.805 56.210 166.195 ;
        RECT 56.605 165.935 56.775 167.295 ;
        RECT 56.945 166.105 57.405 167.155 ;
        RECT 56.380 165.765 56.775 165.935 ;
        RECT 56.380 165.635 56.550 165.765 ;
        RECT 55.405 165.305 56.085 165.635 ;
        RECT 56.300 165.305 56.550 165.635 ;
        RECT 56.720 165.135 56.970 165.595 ;
        RECT 57.140 165.320 57.465 166.105 ;
        RECT 57.635 165.305 57.805 167.425 ;
        RECT 57.975 167.305 58.305 167.685 ;
        RECT 58.475 167.135 58.730 167.425 ;
        RECT 57.980 166.965 58.730 167.135 ;
        RECT 57.980 165.975 58.210 166.965 ;
        RECT 58.905 166.935 60.115 167.685 ;
        RECT 58.380 166.145 58.730 166.795 ;
        RECT 58.905 166.225 59.425 166.765 ;
        RECT 59.595 166.395 60.115 166.935 ;
        RECT 60.375 167.035 60.545 167.515 ;
        RECT 60.725 167.205 60.965 167.685 ;
        RECT 61.215 167.035 61.385 167.515 ;
        RECT 61.555 167.205 61.885 167.685 ;
        RECT 62.055 167.035 62.225 167.515 ;
        RECT 60.375 166.865 61.010 167.035 ;
        RECT 61.215 166.865 62.225 167.035 ;
        RECT 62.395 166.885 62.725 167.685 ;
        RECT 63.045 166.960 63.335 167.685 ;
        RECT 64.515 167.135 64.685 167.515 ;
        RECT 64.865 167.305 65.195 167.685 ;
        RECT 64.515 166.965 65.180 167.135 ;
        RECT 65.375 167.010 65.635 167.515 ;
        RECT 60.840 166.695 61.010 166.865 ;
        RECT 60.290 166.455 60.670 166.695 ;
        RECT 60.840 166.525 61.340 166.695 ;
        RECT 60.840 166.285 61.010 166.525 ;
        RECT 61.730 166.325 62.225 166.865 ;
        RECT 64.445 166.415 64.775 166.785 ;
        RECT 65.010 166.710 65.180 166.965 ;
        RECT 57.980 165.805 58.730 165.975 ;
        RECT 57.975 165.135 58.305 165.635 ;
        RECT 58.475 165.305 58.730 165.805 ;
        RECT 58.905 165.135 60.115 166.225 ;
        RECT 60.295 166.115 61.010 166.285 ;
        RECT 61.215 166.155 62.225 166.325 ;
        RECT 65.010 166.380 65.295 166.710 ;
        RECT 60.295 165.305 60.625 166.115 ;
        RECT 60.795 165.135 61.035 165.935 ;
        RECT 61.215 165.305 61.385 166.155 ;
        RECT 61.555 165.135 61.885 165.935 ;
        RECT 62.055 165.305 62.225 166.155 ;
        RECT 62.395 165.135 62.725 166.285 ;
        RECT 63.045 165.135 63.335 166.300 ;
        RECT 65.010 166.235 65.180 166.380 ;
        RECT 64.515 166.065 65.180 166.235 ;
        RECT 65.465 166.210 65.635 167.010 ;
        RECT 66.265 166.915 68.855 167.685 ;
        RECT 69.030 167.140 74.375 167.685 ;
        RECT 74.555 167.155 74.885 167.515 ;
        RECT 75.055 167.325 75.385 167.685 ;
        RECT 75.585 167.155 75.915 167.515 ;
        RECT 64.515 165.305 64.685 166.065 ;
        RECT 64.865 165.135 65.195 165.895 ;
        RECT 65.365 165.305 65.635 166.210 ;
        RECT 66.265 166.225 67.475 166.745 ;
        RECT 67.645 166.395 68.855 166.915 ;
        RECT 66.265 165.135 68.855 166.225 ;
        RECT 70.620 165.570 70.970 166.820 ;
        RECT 72.450 166.310 72.790 167.140 ;
        RECT 74.555 166.945 75.915 167.155 ;
        RECT 76.425 166.925 77.135 167.515 ;
        RECT 74.545 166.445 74.855 166.775 ;
        RECT 75.065 166.445 75.440 166.775 ;
        RECT 75.760 166.445 76.255 166.775 ;
        RECT 69.030 165.135 74.375 165.570 ;
        RECT 74.555 165.135 74.885 166.195 ;
        RECT 75.065 165.520 75.235 166.445 ;
        RECT 75.405 165.955 75.735 166.175 ;
        RECT 75.930 166.155 76.255 166.445 ;
        RECT 76.430 166.155 76.760 166.695 ;
        RECT 76.930 165.955 77.135 166.925 ;
        RECT 77.305 166.915 78.975 167.685 ;
        RECT 75.405 165.725 77.135 165.955 ;
        RECT 75.405 165.325 75.735 165.725 ;
        RECT 75.905 165.135 76.235 165.495 ;
        RECT 76.435 165.305 77.135 165.725 ;
        RECT 77.305 166.225 78.055 166.745 ;
        RECT 78.225 166.395 78.975 166.915 ;
        RECT 79.520 166.975 79.775 167.505 ;
        RECT 79.955 167.225 80.240 167.685 ;
        RECT 77.305 165.135 78.975 166.225 ;
        RECT 79.520 166.115 79.700 166.975 ;
        RECT 80.420 166.775 80.670 167.425 ;
        RECT 79.870 166.445 80.670 166.775 ;
        RECT 79.520 165.645 79.775 166.115 ;
        RECT 79.435 165.475 79.775 165.645 ;
        RECT 79.520 165.445 79.775 165.475 ;
        RECT 79.955 165.135 80.240 165.935 ;
        RECT 80.420 165.855 80.670 166.445 ;
        RECT 80.870 167.090 81.190 167.420 ;
        RECT 81.370 167.205 82.030 167.685 ;
        RECT 82.230 167.295 83.080 167.465 ;
        RECT 80.870 166.195 81.060 167.090 ;
        RECT 81.380 166.765 82.040 167.035 ;
        RECT 81.710 166.705 82.040 166.765 ;
        RECT 81.230 166.535 81.560 166.595 ;
        RECT 82.230 166.535 82.400 167.295 ;
        RECT 83.640 167.225 83.960 167.685 ;
        RECT 84.160 167.045 84.410 167.475 ;
        RECT 84.700 167.245 85.110 167.685 ;
        RECT 85.280 167.305 86.295 167.505 ;
        RECT 82.570 166.875 83.820 167.045 ;
        RECT 82.570 166.755 82.900 166.875 ;
        RECT 81.230 166.365 83.130 166.535 ;
        RECT 80.870 166.025 82.790 166.195 ;
        RECT 80.870 166.005 81.190 166.025 ;
        RECT 80.420 165.345 80.750 165.855 ;
        RECT 81.020 165.395 81.190 166.005 ;
        RECT 82.960 165.855 83.130 166.365 ;
        RECT 83.300 166.295 83.480 166.705 ;
        RECT 83.650 166.115 83.820 166.875 ;
        RECT 81.360 165.135 81.690 165.825 ;
        RECT 81.920 165.685 83.130 165.855 ;
        RECT 83.300 165.805 83.820 166.115 ;
        RECT 83.990 166.705 84.410 167.045 ;
        RECT 84.700 166.705 85.110 167.035 ;
        RECT 83.990 165.935 84.180 166.705 ;
        RECT 85.280 166.575 85.450 167.305 ;
        RECT 86.595 167.135 86.765 167.465 ;
        RECT 86.935 167.305 87.265 167.685 ;
        RECT 85.620 166.755 85.970 167.125 ;
        RECT 85.280 166.535 85.700 166.575 ;
        RECT 84.350 166.365 85.700 166.535 ;
        RECT 84.350 166.205 84.600 166.365 ;
        RECT 85.110 165.935 85.360 166.195 ;
        RECT 83.990 165.685 85.360 165.935 ;
        RECT 81.920 165.395 82.160 165.685 ;
        RECT 82.960 165.605 83.130 165.685 ;
        RECT 82.360 165.135 82.780 165.515 ;
        RECT 82.960 165.355 83.590 165.605 ;
        RECT 84.060 165.135 84.390 165.515 ;
        RECT 84.560 165.395 84.730 165.685 ;
        RECT 85.530 165.520 85.700 166.365 ;
        RECT 86.150 166.195 86.370 167.065 ;
        RECT 86.595 166.945 87.290 167.135 ;
        RECT 85.870 165.815 86.370 166.195 ;
        RECT 86.540 166.145 86.950 166.765 ;
        RECT 87.120 165.975 87.290 166.945 ;
        RECT 86.595 165.805 87.290 165.975 ;
        RECT 84.910 165.135 85.290 165.515 ;
        RECT 85.530 165.350 86.360 165.520 ;
        RECT 86.595 165.305 86.765 165.805 ;
        RECT 86.935 165.135 87.265 165.635 ;
        RECT 87.480 165.305 87.705 167.425 ;
        RECT 87.875 167.305 88.205 167.685 ;
        RECT 88.375 167.135 88.545 167.425 ;
        RECT 87.880 166.965 88.545 167.135 ;
        RECT 87.880 165.975 88.110 166.965 ;
        RECT 88.805 166.960 89.095 167.685 ;
        RECT 89.265 167.010 89.525 167.515 ;
        RECT 89.705 167.305 90.035 167.685 ;
        RECT 90.215 167.135 90.385 167.515 ;
        RECT 88.280 166.145 88.630 166.795 ;
        RECT 87.880 165.805 88.545 165.975 ;
        RECT 87.875 165.135 88.205 165.635 ;
        RECT 88.375 165.305 88.545 165.805 ;
        RECT 88.805 165.135 89.095 166.300 ;
        RECT 89.265 166.210 89.435 167.010 ;
        RECT 89.720 166.965 90.385 167.135 ;
        RECT 89.720 166.710 89.890 166.965 ;
        RECT 90.705 166.865 90.915 167.685 ;
        RECT 91.085 166.885 91.415 167.515 ;
        RECT 89.605 166.380 89.890 166.710 ;
        RECT 90.125 166.415 90.455 166.785 ;
        RECT 89.720 166.235 89.890 166.380 ;
        RECT 91.085 166.285 91.335 166.885 ;
        RECT 91.585 166.865 91.815 167.685 ;
        RECT 92.115 167.135 92.285 167.515 ;
        RECT 92.465 167.305 92.795 167.685 ;
        RECT 92.115 166.965 92.780 167.135 ;
        RECT 92.975 167.010 93.235 167.515 ;
        RECT 93.870 167.215 94.200 167.685 ;
        RECT 94.370 167.045 94.595 167.490 ;
        RECT 94.765 167.160 95.060 167.685 ;
        RECT 91.505 166.445 91.835 166.695 ;
        RECT 92.045 166.415 92.375 166.785 ;
        RECT 92.610 166.710 92.780 166.965 ;
        RECT 92.610 166.380 92.895 166.710 ;
        RECT 89.265 165.305 89.535 166.210 ;
        RECT 89.720 166.065 90.385 166.235 ;
        RECT 89.705 165.135 90.035 165.895 ;
        RECT 90.215 165.305 90.385 166.065 ;
        RECT 90.705 165.135 90.915 166.275 ;
        RECT 91.085 165.305 91.415 166.285 ;
        RECT 91.585 165.135 91.815 166.275 ;
        RECT 92.610 166.235 92.780 166.380 ;
        RECT 92.115 166.065 92.780 166.235 ;
        RECT 93.065 166.210 93.235 167.010 ;
        RECT 92.115 165.305 92.285 166.065 ;
        RECT 92.465 165.135 92.795 165.895 ;
        RECT 92.965 165.305 93.235 166.210 ;
        RECT 93.865 166.875 94.595 167.045 ;
        RECT 96.080 166.975 96.335 167.505 ;
        RECT 96.515 167.225 96.800 167.685 ;
        RECT 93.865 166.310 94.145 166.875 ;
        RECT 94.315 166.480 95.535 166.705 ;
        RECT 93.865 166.140 95.465 166.310 ;
        RECT 93.925 165.135 94.180 165.970 ;
        RECT 94.350 165.335 94.610 166.140 ;
        RECT 94.780 165.135 95.040 165.970 ;
        RECT 95.210 165.335 95.465 166.140 ;
        RECT 96.080 166.115 96.260 166.975 ;
        RECT 96.980 166.775 97.230 167.425 ;
        RECT 96.430 166.445 97.230 166.775 ;
        RECT 96.080 165.645 96.335 166.115 ;
        RECT 95.995 165.475 96.335 165.645 ;
        RECT 96.080 165.445 96.335 165.475 ;
        RECT 96.515 165.135 96.800 165.935 ;
        RECT 96.980 165.855 97.230 166.445 ;
        RECT 97.430 167.090 97.750 167.420 ;
        RECT 97.930 167.205 98.590 167.685 ;
        RECT 98.790 167.295 99.640 167.465 ;
        RECT 97.430 166.195 97.620 167.090 ;
        RECT 97.940 166.765 98.600 167.035 ;
        RECT 98.270 166.705 98.600 166.765 ;
        RECT 97.790 166.535 98.120 166.595 ;
        RECT 98.790 166.535 98.960 167.295 ;
        RECT 100.200 167.225 100.520 167.685 ;
        RECT 100.720 167.045 100.970 167.475 ;
        RECT 101.260 167.245 101.670 167.685 ;
        RECT 101.840 167.305 102.855 167.505 ;
        RECT 99.130 166.875 100.380 167.045 ;
        RECT 99.130 166.755 99.460 166.875 ;
        RECT 97.790 166.365 99.690 166.535 ;
        RECT 97.430 166.025 99.350 166.195 ;
        RECT 97.430 166.005 97.750 166.025 ;
        RECT 96.980 165.345 97.310 165.855 ;
        RECT 97.580 165.395 97.750 166.005 ;
        RECT 99.520 165.855 99.690 166.365 ;
        RECT 99.860 166.295 100.040 166.705 ;
        RECT 100.210 166.115 100.380 166.875 ;
        RECT 97.920 165.135 98.250 165.825 ;
        RECT 98.480 165.685 99.690 165.855 ;
        RECT 99.860 165.805 100.380 166.115 ;
        RECT 100.550 166.705 100.970 167.045 ;
        RECT 101.260 166.705 101.670 167.035 ;
        RECT 100.550 165.935 100.740 166.705 ;
        RECT 101.840 166.575 102.010 167.305 ;
        RECT 103.155 167.135 103.325 167.465 ;
        RECT 103.495 167.305 103.825 167.685 ;
        RECT 102.180 166.755 102.530 167.125 ;
        RECT 101.840 166.535 102.260 166.575 ;
        RECT 100.910 166.365 102.260 166.535 ;
        RECT 100.910 166.205 101.160 166.365 ;
        RECT 101.670 165.935 101.920 166.195 ;
        RECT 100.550 165.685 101.920 165.935 ;
        RECT 98.480 165.395 98.720 165.685 ;
        RECT 99.520 165.605 99.690 165.685 ;
        RECT 98.920 165.135 99.340 165.515 ;
        RECT 99.520 165.355 100.150 165.605 ;
        RECT 100.620 165.135 100.950 165.515 ;
        RECT 101.120 165.395 101.290 165.685 ;
        RECT 102.090 165.520 102.260 166.365 ;
        RECT 102.710 166.195 102.930 167.065 ;
        RECT 103.155 166.945 103.850 167.135 ;
        RECT 102.430 165.815 102.930 166.195 ;
        RECT 103.100 166.145 103.510 166.765 ;
        RECT 103.680 165.975 103.850 166.945 ;
        RECT 103.155 165.805 103.850 165.975 ;
        RECT 101.470 165.135 101.850 165.515 ;
        RECT 102.090 165.350 102.920 165.520 ;
        RECT 103.155 165.305 103.325 165.805 ;
        RECT 103.495 165.135 103.825 165.635 ;
        RECT 104.040 165.305 104.265 167.425 ;
        RECT 104.435 167.305 104.765 167.685 ;
        RECT 104.935 167.135 105.105 167.425 ;
        RECT 104.440 166.965 105.105 167.135 ;
        RECT 105.370 166.975 105.625 167.505 ;
        RECT 105.795 167.225 106.100 167.685 ;
        RECT 106.345 167.305 107.415 167.475 ;
        RECT 104.440 165.975 104.670 166.965 ;
        RECT 104.840 166.145 105.190 166.795 ;
        RECT 105.370 166.325 105.580 166.975 ;
        RECT 106.345 166.950 106.665 167.305 ;
        RECT 106.340 166.775 106.665 166.950 ;
        RECT 105.750 166.475 106.665 166.775 ;
        RECT 106.835 166.735 107.075 167.135 ;
        RECT 107.245 167.075 107.415 167.305 ;
        RECT 107.585 167.245 107.775 167.685 ;
        RECT 107.945 167.235 108.895 167.515 ;
        RECT 109.115 167.325 109.465 167.495 ;
        RECT 107.245 166.905 107.775 167.075 ;
        RECT 105.750 166.445 106.490 166.475 ;
        RECT 104.440 165.805 105.105 165.975 ;
        RECT 104.435 165.135 104.765 165.635 ;
        RECT 104.935 165.305 105.105 165.805 ;
        RECT 105.370 165.445 105.625 166.325 ;
        RECT 105.795 165.135 106.100 166.275 ;
        RECT 106.320 165.855 106.490 166.445 ;
        RECT 106.835 166.365 107.375 166.735 ;
        RECT 107.555 166.625 107.775 166.905 ;
        RECT 107.945 166.455 108.115 167.235 ;
        RECT 107.710 166.285 108.115 166.455 ;
        RECT 108.285 166.445 108.635 167.065 ;
        RECT 107.710 166.195 107.880 166.285 ;
        RECT 108.805 166.275 109.015 167.065 ;
        RECT 106.660 166.025 107.880 166.195 ;
        RECT 108.340 166.115 109.015 166.275 ;
        RECT 106.320 165.685 107.120 165.855 ;
        RECT 106.440 165.135 106.770 165.515 ;
        RECT 106.950 165.395 107.120 165.685 ;
        RECT 107.710 165.645 107.880 166.025 ;
        RECT 108.050 166.105 109.015 166.115 ;
        RECT 109.205 166.935 109.465 167.325 ;
        RECT 109.675 167.225 110.005 167.685 ;
        RECT 110.880 167.295 111.735 167.465 ;
        RECT 111.940 167.295 112.435 167.465 ;
        RECT 112.605 167.325 112.935 167.685 ;
        RECT 109.205 166.245 109.375 166.935 ;
        RECT 109.545 166.585 109.715 166.765 ;
        RECT 109.885 166.755 110.675 167.005 ;
        RECT 110.880 166.585 111.050 167.295 ;
        RECT 111.220 166.785 111.575 167.005 ;
        RECT 109.545 166.415 111.235 166.585 ;
        RECT 108.050 165.815 108.510 166.105 ;
        RECT 109.205 166.075 110.705 166.245 ;
        RECT 109.205 165.935 109.375 166.075 ;
        RECT 108.815 165.765 109.375 165.935 ;
        RECT 107.290 165.135 107.540 165.595 ;
        RECT 107.710 165.305 108.580 165.645 ;
        RECT 108.815 165.305 108.985 165.765 ;
        RECT 109.820 165.735 110.895 165.905 ;
        RECT 109.155 165.135 109.525 165.595 ;
        RECT 109.820 165.395 109.990 165.735 ;
        RECT 110.160 165.135 110.490 165.565 ;
        RECT 110.725 165.395 110.895 165.735 ;
        RECT 111.065 165.635 111.235 166.415 ;
        RECT 111.405 166.195 111.575 166.785 ;
        RECT 111.745 166.385 112.095 167.005 ;
        RECT 111.405 165.805 111.870 166.195 ;
        RECT 112.265 165.935 112.435 167.295 ;
        RECT 112.605 166.105 113.065 167.155 ;
        RECT 112.040 165.765 112.435 165.935 ;
        RECT 112.040 165.635 112.210 165.765 ;
        RECT 111.065 165.305 111.745 165.635 ;
        RECT 111.960 165.305 112.210 165.635 ;
        RECT 112.380 165.135 112.630 165.595 ;
        RECT 112.800 165.320 113.125 166.105 ;
        RECT 113.295 165.305 113.465 167.425 ;
        RECT 113.635 167.305 113.965 167.685 ;
        RECT 114.135 167.135 114.390 167.425 ;
        RECT 113.640 166.965 114.390 167.135 ;
        RECT 113.640 165.975 113.870 166.965 ;
        RECT 114.565 166.960 114.855 167.685 ;
        RECT 115.490 166.975 115.745 167.505 ;
        RECT 115.915 167.225 116.220 167.685 ;
        RECT 116.465 167.305 117.535 167.475 ;
        RECT 114.040 166.145 114.390 166.795 ;
        RECT 115.490 166.325 115.700 166.975 ;
        RECT 116.465 166.950 116.785 167.305 ;
        RECT 116.460 166.775 116.785 166.950 ;
        RECT 115.870 166.475 116.785 166.775 ;
        RECT 116.955 166.735 117.195 167.135 ;
        RECT 117.365 167.075 117.535 167.305 ;
        RECT 117.705 167.245 117.895 167.685 ;
        RECT 118.065 167.235 119.015 167.515 ;
        RECT 119.235 167.325 119.585 167.495 ;
        RECT 117.365 166.905 117.895 167.075 ;
        RECT 115.870 166.445 116.610 166.475 ;
        RECT 113.640 165.805 114.390 165.975 ;
        RECT 113.635 165.135 113.965 165.635 ;
        RECT 114.135 165.305 114.390 165.805 ;
        RECT 114.565 165.135 114.855 166.300 ;
        RECT 115.490 165.445 115.745 166.325 ;
        RECT 115.915 165.135 116.220 166.275 ;
        RECT 116.440 165.855 116.610 166.445 ;
        RECT 116.955 166.365 117.495 166.735 ;
        RECT 117.675 166.625 117.895 166.905 ;
        RECT 118.065 166.455 118.235 167.235 ;
        RECT 117.830 166.285 118.235 166.455 ;
        RECT 118.405 166.445 118.755 167.065 ;
        RECT 117.830 166.195 118.000 166.285 ;
        RECT 118.925 166.275 119.135 167.065 ;
        RECT 116.780 166.025 118.000 166.195 ;
        RECT 118.460 166.115 119.135 166.275 ;
        RECT 116.440 165.685 117.240 165.855 ;
        RECT 116.560 165.135 116.890 165.515 ;
        RECT 117.070 165.395 117.240 165.685 ;
        RECT 117.830 165.645 118.000 166.025 ;
        RECT 118.170 166.105 119.135 166.115 ;
        RECT 119.325 166.935 119.585 167.325 ;
        RECT 119.795 167.225 120.125 167.685 ;
        RECT 121.000 167.295 121.855 167.465 ;
        RECT 122.060 167.295 122.555 167.465 ;
        RECT 122.725 167.325 123.055 167.685 ;
        RECT 119.325 166.245 119.495 166.935 ;
        RECT 119.665 166.585 119.835 166.765 ;
        RECT 120.005 166.755 120.795 167.005 ;
        RECT 121.000 166.585 121.170 167.295 ;
        RECT 121.340 166.785 121.695 167.005 ;
        RECT 119.665 166.415 121.355 166.585 ;
        RECT 118.170 165.815 118.630 166.105 ;
        RECT 119.325 166.075 120.825 166.245 ;
        RECT 119.325 165.935 119.495 166.075 ;
        RECT 118.935 165.765 119.495 165.935 ;
        RECT 117.410 165.135 117.660 165.595 ;
        RECT 117.830 165.305 118.700 165.645 ;
        RECT 118.935 165.305 119.105 165.765 ;
        RECT 119.940 165.735 121.015 165.905 ;
        RECT 119.275 165.135 119.645 165.595 ;
        RECT 119.940 165.395 120.110 165.735 ;
        RECT 120.280 165.135 120.610 165.565 ;
        RECT 120.845 165.395 121.015 165.735 ;
        RECT 121.185 165.635 121.355 166.415 ;
        RECT 121.525 166.195 121.695 166.785 ;
        RECT 121.865 166.385 122.215 167.005 ;
        RECT 121.525 165.805 121.990 166.195 ;
        RECT 122.385 165.935 122.555 167.295 ;
        RECT 122.725 166.105 123.185 167.155 ;
        RECT 122.160 165.765 122.555 165.935 ;
        RECT 122.160 165.635 122.330 165.765 ;
        RECT 121.185 165.305 121.865 165.635 ;
        RECT 122.080 165.305 122.330 165.635 ;
        RECT 122.500 165.135 122.750 165.595 ;
        RECT 122.920 165.320 123.245 166.105 ;
        RECT 123.415 165.305 123.585 167.425 ;
        RECT 123.755 167.305 124.085 167.685 ;
        RECT 124.255 167.135 124.510 167.425 ;
        RECT 123.760 166.965 124.510 167.135 ;
        RECT 123.760 165.975 123.990 166.965 ;
        RECT 124.685 166.915 126.355 167.685 ;
        RECT 126.525 166.935 127.735 167.685 ;
        RECT 124.160 166.145 124.510 166.795 ;
        RECT 124.685 166.225 125.435 166.745 ;
        RECT 125.605 166.395 126.355 166.915 ;
        RECT 126.525 166.225 127.045 166.765 ;
        RECT 127.215 166.395 127.735 166.935 ;
        RECT 123.760 165.805 124.510 165.975 ;
        RECT 123.755 165.135 124.085 165.635 ;
        RECT 124.255 165.305 124.510 165.805 ;
        RECT 124.685 165.135 126.355 166.225 ;
        RECT 126.525 165.135 127.735 166.225 ;
        RECT 20.640 164.965 127.820 165.135 ;
        RECT 20.725 163.875 21.935 164.965 ;
        RECT 20.725 163.165 21.245 163.705 ;
        RECT 21.415 163.335 21.935 163.875 ;
        RECT 22.565 163.875 24.235 164.965 ;
        RECT 22.565 163.355 23.315 163.875 ;
        RECT 24.405 163.800 24.695 164.965 ;
        RECT 25.385 163.825 25.595 164.965 ;
        RECT 25.765 163.815 26.095 164.795 ;
        RECT 26.265 163.825 26.495 164.965 ;
        RECT 26.705 164.205 27.220 164.615 ;
        RECT 27.455 164.205 27.625 164.965 ;
        RECT 27.795 164.625 29.825 164.795 ;
        RECT 23.485 163.185 24.235 163.705 ;
        RECT 20.725 162.415 21.935 163.165 ;
        RECT 22.565 162.415 24.235 163.185 ;
        RECT 24.405 162.415 24.695 163.140 ;
        RECT 25.385 162.415 25.595 163.235 ;
        RECT 25.765 163.215 26.015 163.815 ;
        RECT 26.185 163.405 26.515 163.655 ;
        RECT 26.705 163.395 27.045 164.205 ;
        RECT 27.795 163.960 27.965 164.625 ;
        RECT 28.360 164.285 29.485 164.455 ;
        RECT 27.215 163.770 27.965 163.960 ;
        RECT 28.135 163.945 29.145 164.115 ;
        RECT 25.765 162.585 26.095 163.215 ;
        RECT 26.265 162.415 26.495 163.235 ;
        RECT 26.705 163.225 27.935 163.395 ;
        RECT 26.980 162.620 27.225 163.225 ;
        RECT 27.445 162.415 27.955 162.950 ;
        RECT 28.135 162.585 28.325 163.945 ;
        RECT 28.495 163.265 28.770 163.745 ;
        RECT 28.495 163.095 28.775 163.265 ;
        RECT 28.975 163.145 29.145 163.945 ;
        RECT 29.315 163.155 29.485 164.285 ;
        RECT 29.655 163.655 29.825 164.625 ;
        RECT 29.995 163.825 30.165 164.965 ;
        RECT 30.335 163.825 30.670 164.795 ;
        RECT 31.395 164.035 31.565 164.795 ;
        RECT 31.745 164.205 32.075 164.965 ;
        RECT 31.395 163.865 32.060 164.035 ;
        RECT 32.245 163.890 32.515 164.795 ;
        RECT 29.655 163.325 29.850 163.655 ;
        RECT 30.075 163.325 30.330 163.655 ;
        RECT 30.075 163.155 30.245 163.325 ;
        RECT 30.500 163.155 30.670 163.825 ;
        RECT 31.890 163.720 32.060 163.865 ;
        RECT 31.325 163.315 31.655 163.685 ;
        RECT 31.890 163.390 32.175 163.720 ;
        RECT 28.495 162.585 28.770 163.095 ;
        RECT 29.315 162.985 30.245 163.155 ;
        RECT 29.315 162.950 29.490 162.985 ;
        RECT 28.960 162.585 29.490 162.950 ;
        RECT 29.915 162.415 30.245 162.815 ;
        RECT 30.415 162.585 30.670 163.155 ;
        RECT 31.890 163.135 32.060 163.390 ;
        RECT 31.395 162.965 32.060 163.135 ;
        RECT 32.345 163.090 32.515 163.890 ;
        RECT 32.725 163.825 32.955 164.965 ;
        RECT 33.125 163.815 33.455 164.795 ;
        RECT 33.625 163.825 33.835 164.965 ;
        RECT 34.070 164.530 39.415 164.965 ;
        RECT 32.705 163.405 33.035 163.655 ;
        RECT 31.395 162.585 31.565 162.965 ;
        RECT 31.745 162.415 32.075 162.795 ;
        RECT 32.255 162.585 32.515 163.090 ;
        RECT 32.725 162.415 32.955 163.235 ;
        RECT 33.205 163.215 33.455 163.815 ;
        RECT 35.660 163.280 36.010 164.530 ;
        RECT 39.590 163.825 39.925 164.795 ;
        RECT 40.095 163.825 40.265 164.965 ;
        RECT 40.435 164.625 42.465 164.795 ;
        RECT 33.125 162.585 33.455 163.215 ;
        RECT 33.625 162.415 33.835 163.235 ;
        RECT 37.490 162.960 37.830 163.790 ;
        RECT 39.590 163.155 39.760 163.825 ;
        RECT 40.435 163.655 40.605 164.625 ;
        RECT 39.930 163.325 40.185 163.655 ;
        RECT 40.410 163.325 40.605 163.655 ;
        RECT 40.775 164.285 41.900 164.455 ;
        RECT 40.015 163.155 40.185 163.325 ;
        RECT 40.775 163.155 40.945 164.285 ;
        RECT 34.070 162.415 39.415 162.960 ;
        RECT 39.590 162.585 39.845 163.155 ;
        RECT 40.015 162.985 40.945 163.155 ;
        RECT 41.115 163.945 42.125 164.115 ;
        RECT 41.115 163.145 41.285 163.945 ;
        RECT 41.490 163.265 41.765 163.745 ;
        RECT 41.485 163.095 41.765 163.265 ;
        RECT 40.770 162.950 40.945 162.985 ;
        RECT 40.015 162.415 40.345 162.815 ;
        RECT 40.770 162.585 41.300 162.950 ;
        RECT 41.490 162.585 41.765 163.095 ;
        RECT 41.935 162.585 42.125 163.945 ;
        RECT 42.295 163.960 42.465 164.625 ;
        RECT 42.635 164.205 42.805 164.965 ;
        RECT 43.040 164.205 43.555 164.615 ;
        RECT 42.295 163.770 43.045 163.960 ;
        RECT 43.215 163.395 43.555 164.205 ;
        RECT 42.325 163.225 43.555 163.395 ;
        RECT 43.725 163.875 44.935 164.965 ;
        RECT 45.105 163.875 48.615 164.965 ;
        RECT 48.785 163.890 49.055 164.795 ;
        RECT 49.225 164.205 49.555 164.965 ;
        RECT 49.735 164.035 49.905 164.795 ;
        RECT 43.725 163.335 44.245 163.875 ;
        RECT 42.305 162.415 42.815 162.950 ;
        RECT 43.035 162.620 43.280 163.225 ;
        RECT 44.415 163.165 44.935 163.705 ;
        RECT 45.105 163.355 46.795 163.875 ;
        RECT 46.965 163.185 48.615 163.705 ;
        RECT 43.725 162.415 44.935 163.165 ;
        RECT 45.105 162.415 48.615 163.185 ;
        RECT 48.785 163.090 48.955 163.890 ;
        RECT 49.240 163.865 49.905 164.035 ;
        RECT 49.240 163.720 49.410 163.865 ;
        RECT 50.165 163.800 50.455 164.965 ;
        RECT 51.085 163.875 52.755 164.965 ;
        RECT 49.125 163.390 49.410 163.720 ;
        RECT 49.240 163.135 49.410 163.390 ;
        RECT 49.645 163.315 49.975 163.685 ;
        RECT 51.085 163.355 51.835 163.875 ;
        RECT 52.985 163.825 53.195 164.965 ;
        RECT 53.365 163.815 53.695 164.795 ;
        RECT 53.865 163.825 54.095 164.965 ;
        RECT 54.395 164.035 54.565 164.795 ;
        RECT 54.745 164.205 55.075 164.965 ;
        RECT 54.395 163.865 55.060 164.035 ;
        RECT 55.245 163.890 55.515 164.795 ;
        RECT 52.005 163.185 52.755 163.705 ;
        RECT 48.785 162.585 49.045 163.090 ;
        RECT 49.240 162.965 49.905 163.135 ;
        RECT 49.225 162.415 49.555 162.795 ;
        RECT 49.735 162.585 49.905 162.965 ;
        RECT 50.165 162.415 50.455 163.140 ;
        RECT 51.085 162.415 52.755 163.185 ;
        RECT 52.985 162.415 53.195 163.235 ;
        RECT 53.365 163.215 53.615 163.815 ;
        RECT 54.890 163.720 55.060 163.865 ;
        RECT 53.785 163.405 54.115 163.655 ;
        RECT 54.325 163.315 54.655 163.685 ;
        RECT 54.890 163.390 55.175 163.720 ;
        RECT 53.365 162.585 53.695 163.215 ;
        RECT 53.865 162.415 54.095 163.235 ;
        RECT 54.890 163.135 55.060 163.390 ;
        RECT 54.395 162.965 55.060 163.135 ;
        RECT 55.345 163.090 55.515 163.890 ;
        RECT 55.685 163.875 56.895 164.965 ;
        RECT 55.685 163.335 56.205 163.875 ;
        RECT 57.105 163.825 57.335 164.965 ;
        RECT 57.505 163.815 57.835 164.795 ;
        RECT 58.005 163.825 58.215 164.965 ;
        RECT 58.820 163.985 59.075 164.655 ;
        RECT 59.255 164.165 59.540 164.965 ;
        RECT 59.720 164.245 60.050 164.755 ;
        RECT 56.375 163.165 56.895 163.705 ;
        RECT 57.085 163.405 57.415 163.655 ;
        RECT 54.395 162.585 54.565 162.965 ;
        RECT 54.745 162.415 55.075 162.795 ;
        RECT 55.255 162.585 55.515 163.090 ;
        RECT 55.685 162.415 56.895 163.165 ;
        RECT 57.105 162.415 57.335 163.235 ;
        RECT 57.585 163.215 57.835 163.815 ;
        RECT 57.505 162.585 57.835 163.215 ;
        RECT 58.005 162.415 58.215 163.235 ;
        RECT 58.820 163.125 59.000 163.985 ;
        RECT 59.720 163.655 59.970 164.245 ;
        RECT 60.320 164.095 60.490 164.705 ;
        RECT 60.660 164.275 60.990 164.965 ;
        RECT 61.220 164.415 61.460 164.705 ;
        RECT 61.660 164.585 62.080 164.965 ;
        RECT 62.260 164.495 62.890 164.745 ;
        RECT 63.360 164.585 63.690 164.965 ;
        RECT 62.260 164.415 62.430 164.495 ;
        RECT 63.860 164.415 64.030 164.705 ;
        RECT 64.210 164.585 64.590 164.965 ;
        RECT 64.830 164.580 65.660 164.750 ;
        RECT 61.220 164.245 62.430 164.415 ;
        RECT 59.170 163.325 59.970 163.655 ;
        RECT 58.820 162.925 59.075 163.125 ;
        RECT 58.735 162.755 59.075 162.925 ;
        RECT 58.820 162.595 59.075 162.755 ;
        RECT 59.255 162.415 59.540 162.875 ;
        RECT 59.720 162.675 59.970 163.325 ;
        RECT 60.170 164.075 60.490 164.095 ;
        RECT 60.170 163.905 62.090 164.075 ;
        RECT 60.170 163.010 60.360 163.905 ;
        RECT 62.260 163.735 62.430 164.245 ;
        RECT 62.600 163.985 63.120 164.295 ;
        RECT 60.530 163.565 62.430 163.735 ;
        RECT 60.530 163.505 60.860 163.565 ;
        RECT 61.010 163.335 61.340 163.395 ;
        RECT 60.680 163.065 61.340 163.335 ;
        RECT 60.170 162.680 60.490 163.010 ;
        RECT 60.670 162.415 61.330 162.895 ;
        RECT 61.530 162.805 61.700 163.565 ;
        RECT 62.600 163.395 62.780 163.805 ;
        RECT 61.870 163.225 62.200 163.345 ;
        RECT 62.950 163.225 63.120 163.985 ;
        RECT 61.870 163.055 63.120 163.225 ;
        RECT 63.290 164.165 64.660 164.415 ;
        RECT 63.290 163.395 63.480 164.165 ;
        RECT 64.410 163.905 64.660 164.165 ;
        RECT 63.650 163.735 63.900 163.895 ;
        RECT 64.830 163.735 65.000 164.580 ;
        RECT 65.895 164.295 66.065 164.795 ;
        RECT 66.235 164.465 66.565 164.965 ;
        RECT 65.170 163.905 65.670 164.285 ;
        RECT 65.895 164.125 66.590 164.295 ;
        RECT 63.650 163.565 65.000 163.735 ;
        RECT 64.580 163.525 65.000 163.565 ;
        RECT 63.290 163.055 63.710 163.395 ;
        RECT 64.000 163.065 64.410 163.395 ;
        RECT 61.530 162.635 62.380 162.805 ;
        RECT 62.940 162.415 63.260 162.875 ;
        RECT 63.460 162.625 63.710 163.055 ;
        RECT 64.000 162.415 64.410 162.855 ;
        RECT 64.580 162.795 64.750 163.525 ;
        RECT 64.920 162.975 65.270 163.345 ;
        RECT 65.450 163.035 65.670 163.905 ;
        RECT 65.840 163.335 66.250 163.955 ;
        RECT 66.420 163.155 66.590 164.125 ;
        RECT 65.895 162.965 66.590 163.155 ;
        RECT 64.580 162.595 65.595 162.795 ;
        RECT 65.895 162.635 66.065 162.965 ;
        RECT 66.235 162.415 66.565 162.795 ;
        RECT 66.780 162.675 67.005 164.795 ;
        RECT 67.175 164.465 67.505 164.965 ;
        RECT 67.675 164.295 67.845 164.795 ;
        RECT 67.180 164.125 67.845 164.295 ;
        RECT 67.180 163.135 67.410 164.125 ;
        RECT 67.580 163.305 67.930 163.955 ;
        RECT 68.105 163.875 70.695 164.965 ;
        RECT 68.105 163.355 69.315 163.875 ;
        RECT 70.870 163.815 71.130 164.965 ;
        RECT 71.305 163.890 71.560 164.795 ;
        RECT 71.730 164.205 72.060 164.965 ;
        RECT 72.275 164.035 72.445 164.795 ;
        RECT 69.485 163.185 70.695 163.705 ;
        RECT 67.180 162.965 67.845 163.135 ;
        RECT 67.175 162.415 67.505 162.795 ;
        RECT 67.675 162.675 67.845 162.965 ;
        RECT 68.105 162.415 70.695 163.185 ;
        RECT 70.870 162.415 71.130 163.255 ;
        RECT 71.305 163.160 71.475 163.890 ;
        RECT 71.730 163.865 72.445 164.035 ;
        RECT 72.795 164.035 72.965 164.795 ;
        RECT 73.180 164.205 73.510 164.965 ;
        RECT 72.795 163.865 73.510 164.035 ;
        RECT 73.680 163.890 73.935 164.795 ;
        RECT 71.730 163.655 71.900 163.865 ;
        RECT 71.645 163.325 71.900 163.655 ;
        RECT 71.305 162.585 71.560 163.160 ;
        RECT 71.730 163.135 71.900 163.325 ;
        RECT 72.180 163.315 72.535 163.685 ;
        RECT 72.705 163.315 73.060 163.685 ;
        RECT 73.340 163.655 73.510 163.865 ;
        RECT 73.340 163.325 73.595 163.655 ;
        RECT 73.340 163.135 73.510 163.325 ;
        RECT 73.765 163.160 73.935 163.890 ;
        RECT 74.110 163.815 74.370 164.965 ;
        RECT 74.545 163.875 75.755 164.965 ;
        RECT 74.545 163.335 75.065 163.875 ;
        RECT 75.925 163.800 76.215 164.965 ;
        RECT 76.850 164.530 82.195 164.965 ;
        RECT 71.730 162.965 72.445 163.135 ;
        RECT 71.730 162.415 72.060 162.795 ;
        RECT 72.275 162.585 72.445 162.965 ;
        RECT 72.795 162.965 73.510 163.135 ;
        RECT 72.795 162.585 72.965 162.965 ;
        RECT 73.180 162.415 73.510 162.795 ;
        RECT 73.680 162.585 73.935 163.160 ;
        RECT 74.110 162.415 74.370 163.255 ;
        RECT 75.235 163.165 75.755 163.705 ;
        RECT 78.440 163.280 78.790 164.530 ;
        RECT 82.365 164.205 82.880 164.615 ;
        RECT 83.115 164.205 83.285 164.965 ;
        RECT 83.455 164.625 85.485 164.795 ;
        RECT 74.545 162.415 75.755 163.165 ;
        RECT 75.925 162.415 76.215 163.140 ;
        RECT 80.270 162.960 80.610 163.790 ;
        RECT 82.365 163.395 82.705 164.205 ;
        RECT 83.455 163.960 83.625 164.625 ;
        RECT 84.020 164.285 85.145 164.455 ;
        RECT 82.875 163.770 83.625 163.960 ;
        RECT 83.795 163.945 84.805 164.115 ;
        RECT 82.365 163.225 83.595 163.395 ;
        RECT 76.850 162.415 82.195 162.960 ;
        RECT 82.640 162.620 82.885 163.225 ;
        RECT 83.105 162.415 83.615 162.950 ;
        RECT 83.795 162.585 83.985 163.945 ;
        RECT 84.155 163.265 84.430 163.745 ;
        RECT 84.155 163.095 84.435 163.265 ;
        RECT 84.635 163.145 84.805 163.945 ;
        RECT 84.975 163.155 85.145 164.285 ;
        RECT 85.315 163.655 85.485 164.625 ;
        RECT 85.655 163.825 85.825 164.965 ;
        RECT 85.995 163.825 86.330 164.795 ;
        RECT 85.315 163.325 85.510 163.655 ;
        RECT 85.735 163.325 85.990 163.655 ;
        RECT 85.735 163.155 85.905 163.325 ;
        RECT 86.160 163.155 86.330 163.825 ;
        RECT 84.155 162.585 84.430 163.095 ;
        RECT 84.975 162.985 85.905 163.155 ;
        RECT 84.975 162.950 85.150 162.985 ;
        RECT 84.620 162.585 85.150 162.950 ;
        RECT 85.575 162.415 85.905 162.815 ;
        RECT 86.075 162.585 86.330 163.155 ;
        RECT 86.880 163.985 87.135 164.655 ;
        RECT 87.315 164.165 87.600 164.965 ;
        RECT 87.780 164.245 88.110 164.755 ;
        RECT 86.880 163.125 87.060 163.985 ;
        RECT 87.780 163.655 88.030 164.245 ;
        RECT 88.380 164.095 88.550 164.705 ;
        RECT 88.720 164.275 89.050 164.965 ;
        RECT 89.280 164.415 89.520 164.705 ;
        RECT 89.720 164.585 90.140 164.965 ;
        RECT 90.320 164.495 90.950 164.745 ;
        RECT 91.420 164.585 91.750 164.965 ;
        RECT 90.320 164.415 90.490 164.495 ;
        RECT 91.920 164.415 92.090 164.705 ;
        RECT 92.270 164.585 92.650 164.965 ;
        RECT 92.890 164.580 93.720 164.750 ;
        RECT 89.280 164.245 90.490 164.415 ;
        RECT 87.230 163.325 88.030 163.655 ;
        RECT 86.880 162.925 87.135 163.125 ;
        RECT 86.795 162.755 87.135 162.925 ;
        RECT 86.880 162.595 87.135 162.755 ;
        RECT 87.315 162.415 87.600 162.875 ;
        RECT 87.780 162.675 88.030 163.325 ;
        RECT 88.230 164.075 88.550 164.095 ;
        RECT 88.230 163.905 90.150 164.075 ;
        RECT 88.230 163.010 88.420 163.905 ;
        RECT 90.320 163.735 90.490 164.245 ;
        RECT 90.660 163.985 91.180 164.295 ;
        RECT 88.590 163.565 90.490 163.735 ;
        RECT 88.590 163.505 88.920 163.565 ;
        RECT 89.070 163.335 89.400 163.395 ;
        RECT 88.740 163.065 89.400 163.335 ;
        RECT 88.230 162.680 88.550 163.010 ;
        RECT 88.730 162.415 89.390 162.895 ;
        RECT 89.590 162.805 89.760 163.565 ;
        RECT 90.660 163.395 90.840 163.805 ;
        RECT 89.930 163.225 90.260 163.345 ;
        RECT 91.010 163.225 91.180 163.985 ;
        RECT 89.930 163.055 91.180 163.225 ;
        RECT 91.350 164.165 92.720 164.415 ;
        RECT 91.350 163.395 91.540 164.165 ;
        RECT 92.470 163.905 92.720 164.165 ;
        RECT 91.710 163.735 91.960 163.895 ;
        RECT 92.890 163.735 93.060 164.580 ;
        RECT 93.955 164.295 94.125 164.795 ;
        RECT 94.295 164.465 94.625 164.965 ;
        RECT 93.230 163.905 93.730 164.285 ;
        RECT 93.955 164.125 94.650 164.295 ;
        RECT 91.710 163.565 93.060 163.735 ;
        RECT 92.640 163.525 93.060 163.565 ;
        RECT 91.350 163.055 91.770 163.395 ;
        RECT 92.060 163.065 92.470 163.395 ;
        RECT 89.590 162.635 90.440 162.805 ;
        RECT 91.000 162.415 91.320 162.875 ;
        RECT 91.520 162.625 91.770 163.055 ;
        RECT 92.060 162.415 92.470 162.855 ;
        RECT 92.640 162.795 92.810 163.525 ;
        RECT 92.980 162.975 93.330 163.345 ;
        RECT 93.510 163.035 93.730 163.905 ;
        RECT 93.900 163.335 94.310 163.955 ;
        RECT 94.480 163.155 94.650 164.125 ;
        RECT 93.955 162.965 94.650 163.155 ;
        RECT 92.640 162.595 93.655 162.795 ;
        RECT 93.955 162.635 94.125 162.965 ;
        RECT 94.295 162.415 94.625 162.795 ;
        RECT 94.840 162.675 95.065 164.795 ;
        RECT 95.235 164.465 95.565 164.965 ;
        RECT 95.735 164.295 95.905 164.795 ;
        RECT 95.240 164.125 95.905 164.295 ;
        RECT 95.240 163.135 95.470 164.125 ;
        RECT 95.640 163.305 95.990 163.955 ;
        RECT 96.165 163.875 97.375 164.965 ;
        RECT 97.545 164.205 98.060 164.615 ;
        RECT 98.295 164.205 98.465 164.965 ;
        RECT 98.635 164.625 100.665 164.795 ;
        RECT 96.165 163.335 96.685 163.875 ;
        RECT 96.855 163.165 97.375 163.705 ;
        RECT 97.545 163.395 97.885 164.205 ;
        RECT 98.635 163.960 98.805 164.625 ;
        RECT 99.200 164.285 100.325 164.455 ;
        RECT 98.055 163.770 98.805 163.960 ;
        RECT 98.975 163.945 99.985 164.115 ;
        RECT 97.545 163.225 98.775 163.395 ;
        RECT 95.240 162.965 95.905 163.135 ;
        RECT 95.235 162.415 95.565 162.795 ;
        RECT 95.735 162.675 95.905 162.965 ;
        RECT 96.165 162.415 97.375 163.165 ;
        RECT 97.820 162.620 98.065 163.225 ;
        RECT 98.285 162.415 98.795 162.950 ;
        RECT 98.975 162.585 99.165 163.945 ;
        RECT 99.335 162.925 99.610 163.745 ;
        RECT 99.815 163.145 99.985 163.945 ;
        RECT 100.155 163.155 100.325 164.285 ;
        RECT 100.495 163.655 100.665 164.625 ;
        RECT 100.835 163.825 101.005 164.965 ;
        RECT 101.175 163.825 101.510 164.795 ;
        RECT 100.495 163.325 100.690 163.655 ;
        RECT 100.915 163.325 101.170 163.655 ;
        RECT 100.915 163.155 101.085 163.325 ;
        RECT 101.340 163.155 101.510 163.825 ;
        RECT 101.685 163.800 101.975 164.965 ;
        RECT 102.520 163.985 102.775 164.655 ;
        RECT 102.955 164.165 103.240 164.965 ;
        RECT 103.420 164.245 103.750 164.755 ;
        RECT 100.155 162.985 101.085 163.155 ;
        RECT 100.155 162.950 100.330 162.985 ;
        RECT 99.335 162.755 99.615 162.925 ;
        RECT 99.335 162.585 99.610 162.755 ;
        RECT 99.800 162.585 100.330 162.950 ;
        RECT 100.755 162.415 101.085 162.815 ;
        RECT 101.255 162.585 101.510 163.155 ;
        RECT 101.685 162.415 101.975 163.140 ;
        RECT 102.520 163.125 102.700 163.985 ;
        RECT 103.420 163.655 103.670 164.245 ;
        RECT 104.020 164.095 104.190 164.705 ;
        RECT 104.360 164.275 104.690 164.965 ;
        RECT 104.920 164.415 105.160 164.705 ;
        RECT 105.360 164.585 105.780 164.965 ;
        RECT 105.960 164.495 106.590 164.745 ;
        RECT 107.060 164.585 107.390 164.965 ;
        RECT 105.960 164.415 106.130 164.495 ;
        RECT 107.560 164.415 107.730 164.705 ;
        RECT 107.910 164.585 108.290 164.965 ;
        RECT 108.530 164.580 109.360 164.750 ;
        RECT 104.920 164.245 106.130 164.415 ;
        RECT 102.870 163.325 103.670 163.655 ;
        RECT 102.520 162.925 102.775 163.125 ;
        RECT 102.435 162.755 102.775 162.925 ;
        RECT 102.520 162.595 102.775 162.755 ;
        RECT 102.955 162.415 103.240 162.875 ;
        RECT 103.420 162.675 103.670 163.325 ;
        RECT 103.870 164.075 104.190 164.095 ;
        RECT 103.870 163.905 105.790 164.075 ;
        RECT 103.870 163.010 104.060 163.905 ;
        RECT 105.960 163.735 106.130 164.245 ;
        RECT 106.300 163.985 106.820 164.295 ;
        RECT 104.230 163.565 106.130 163.735 ;
        RECT 104.230 163.505 104.560 163.565 ;
        RECT 104.710 163.335 105.040 163.395 ;
        RECT 104.380 163.065 105.040 163.335 ;
        RECT 103.870 162.680 104.190 163.010 ;
        RECT 104.370 162.415 105.030 162.895 ;
        RECT 105.230 162.805 105.400 163.565 ;
        RECT 106.300 163.395 106.480 163.805 ;
        RECT 105.570 163.225 105.900 163.345 ;
        RECT 106.650 163.225 106.820 163.985 ;
        RECT 105.570 163.055 106.820 163.225 ;
        RECT 106.990 164.165 108.360 164.415 ;
        RECT 106.990 163.395 107.180 164.165 ;
        RECT 108.110 163.905 108.360 164.165 ;
        RECT 107.350 163.735 107.600 163.895 ;
        RECT 108.530 163.735 108.700 164.580 ;
        RECT 109.595 164.295 109.765 164.795 ;
        RECT 109.935 164.465 110.265 164.965 ;
        RECT 108.870 163.905 109.370 164.285 ;
        RECT 109.595 164.125 110.290 164.295 ;
        RECT 107.350 163.565 108.700 163.735 ;
        RECT 108.280 163.525 108.700 163.565 ;
        RECT 106.990 163.055 107.410 163.395 ;
        RECT 107.700 163.065 108.110 163.395 ;
        RECT 105.230 162.635 106.080 162.805 ;
        RECT 106.640 162.415 106.960 162.875 ;
        RECT 107.160 162.625 107.410 163.055 ;
        RECT 107.700 162.415 108.110 162.855 ;
        RECT 108.280 162.795 108.450 163.525 ;
        RECT 108.620 162.975 108.970 163.345 ;
        RECT 109.150 163.035 109.370 163.905 ;
        RECT 109.540 163.335 109.950 163.955 ;
        RECT 110.120 163.155 110.290 164.125 ;
        RECT 109.595 162.965 110.290 163.155 ;
        RECT 108.280 162.595 109.295 162.795 ;
        RECT 109.595 162.635 109.765 162.965 ;
        RECT 109.935 162.415 110.265 162.795 ;
        RECT 110.480 162.675 110.705 164.795 ;
        RECT 110.875 164.465 111.205 164.965 ;
        RECT 111.375 164.295 111.545 164.795 ;
        RECT 110.880 164.125 111.545 164.295 ;
        RECT 110.880 163.135 111.110 164.125 ;
        RECT 111.280 163.305 111.630 163.955 ;
        RECT 112.265 163.875 113.935 164.965 ;
        RECT 114.105 163.890 114.375 164.795 ;
        RECT 114.545 164.205 114.875 164.965 ;
        RECT 115.055 164.035 115.225 164.795 ;
        RECT 112.265 163.355 113.015 163.875 ;
        RECT 113.185 163.185 113.935 163.705 ;
        RECT 110.880 162.965 111.545 163.135 ;
        RECT 110.875 162.415 111.205 162.795 ;
        RECT 111.375 162.675 111.545 162.965 ;
        RECT 112.265 162.415 113.935 163.185 ;
        RECT 114.105 163.090 114.275 163.890 ;
        RECT 114.560 163.865 115.225 164.035 ;
        RECT 115.485 164.205 116.000 164.615 ;
        RECT 116.235 164.205 116.405 164.965 ;
        RECT 116.575 164.625 118.605 164.795 ;
        RECT 114.560 163.720 114.730 163.865 ;
        RECT 114.445 163.390 114.730 163.720 ;
        RECT 114.560 163.135 114.730 163.390 ;
        RECT 114.965 163.315 115.295 163.685 ;
        RECT 115.485 163.395 115.825 164.205 ;
        RECT 116.575 163.960 116.745 164.625 ;
        RECT 117.140 164.285 118.265 164.455 ;
        RECT 115.995 163.770 116.745 163.960 ;
        RECT 116.915 163.945 117.925 164.115 ;
        RECT 115.485 163.225 116.715 163.395 ;
        RECT 114.105 162.585 114.365 163.090 ;
        RECT 114.560 162.965 115.225 163.135 ;
        RECT 114.545 162.415 114.875 162.795 ;
        RECT 115.055 162.585 115.225 162.965 ;
        RECT 115.760 162.620 116.005 163.225 ;
        RECT 116.225 162.415 116.735 162.950 ;
        RECT 116.915 162.585 117.105 163.945 ;
        RECT 117.275 163.265 117.550 163.745 ;
        RECT 117.275 163.095 117.555 163.265 ;
        RECT 117.755 163.145 117.925 163.945 ;
        RECT 118.095 163.155 118.265 164.285 ;
        RECT 118.435 163.655 118.605 164.625 ;
        RECT 118.775 163.825 118.945 164.965 ;
        RECT 119.115 163.825 119.450 164.795 ;
        RECT 120.635 164.035 120.805 164.795 ;
        RECT 120.985 164.205 121.315 164.965 ;
        RECT 120.635 163.865 121.300 164.035 ;
        RECT 121.485 163.890 121.755 164.795 ;
        RECT 118.435 163.325 118.630 163.655 ;
        RECT 118.855 163.325 119.110 163.655 ;
        RECT 118.855 163.155 119.025 163.325 ;
        RECT 119.280 163.155 119.450 163.825 ;
        RECT 121.130 163.720 121.300 163.865 ;
        RECT 120.565 163.315 120.895 163.685 ;
        RECT 121.130 163.390 121.415 163.720 ;
        RECT 117.275 162.585 117.550 163.095 ;
        RECT 118.095 162.985 119.025 163.155 ;
        RECT 118.095 162.950 118.270 162.985 ;
        RECT 117.740 162.585 118.270 162.950 ;
        RECT 118.695 162.415 119.025 162.815 ;
        RECT 119.195 162.585 119.450 163.155 ;
        RECT 121.130 163.135 121.300 163.390 ;
        RECT 120.635 162.965 121.300 163.135 ;
        RECT 121.585 163.090 121.755 163.890 ;
        RECT 122.845 163.875 126.355 164.965 ;
        RECT 126.525 163.875 127.735 164.965 ;
        RECT 122.845 163.355 124.535 163.875 ;
        RECT 124.705 163.185 126.355 163.705 ;
        RECT 126.525 163.335 127.045 163.875 ;
        RECT 120.635 162.585 120.805 162.965 ;
        RECT 120.985 162.415 121.315 162.795 ;
        RECT 121.495 162.585 121.755 163.090 ;
        RECT 122.845 162.415 126.355 163.185 ;
        RECT 127.215 163.165 127.735 163.705 ;
        RECT 126.525 162.415 127.735 163.165 ;
        RECT 20.640 162.245 127.820 162.415 ;
        RECT 20.725 161.495 21.935 162.245 ;
        RECT 23.400 161.905 23.655 162.065 ;
        RECT 23.315 161.735 23.655 161.905 ;
        RECT 23.835 161.785 24.120 162.245 ;
        RECT 23.400 161.535 23.655 161.735 ;
        RECT 20.725 160.955 21.245 161.495 ;
        RECT 21.415 160.785 21.935 161.325 ;
        RECT 20.725 159.695 21.935 160.785 ;
        RECT 23.400 160.675 23.580 161.535 ;
        RECT 24.300 161.335 24.550 161.985 ;
        RECT 23.750 161.005 24.550 161.335 ;
        RECT 23.400 160.005 23.655 160.675 ;
        RECT 23.835 159.695 24.120 160.495 ;
        RECT 24.300 160.415 24.550 161.005 ;
        RECT 24.750 161.650 25.070 161.980 ;
        RECT 25.250 161.765 25.910 162.245 ;
        RECT 26.110 161.855 26.960 162.025 ;
        RECT 24.750 160.755 24.940 161.650 ;
        RECT 25.260 161.325 25.920 161.595 ;
        RECT 25.590 161.265 25.920 161.325 ;
        RECT 25.110 161.095 25.440 161.155 ;
        RECT 26.110 161.095 26.280 161.855 ;
        RECT 27.520 161.785 27.840 162.245 ;
        RECT 28.040 161.605 28.290 162.035 ;
        RECT 28.580 161.805 28.990 162.245 ;
        RECT 29.160 161.865 30.175 162.065 ;
        RECT 26.450 161.435 27.700 161.605 ;
        RECT 26.450 161.315 26.780 161.435 ;
        RECT 25.110 160.925 27.010 161.095 ;
        RECT 24.750 160.585 26.670 160.755 ;
        RECT 24.750 160.565 25.070 160.585 ;
        RECT 24.300 159.905 24.630 160.415 ;
        RECT 24.900 159.955 25.070 160.565 ;
        RECT 26.840 160.415 27.010 160.925 ;
        RECT 27.180 160.855 27.360 161.265 ;
        RECT 27.530 160.675 27.700 161.435 ;
        RECT 25.240 159.695 25.570 160.385 ;
        RECT 25.800 160.245 27.010 160.415 ;
        RECT 27.180 160.365 27.700 160.675 ;
        RECT 27.870 161.265 28.290 161.605 ;
        RECT 28.580 161.265 28.990 161.595 ;
        RECT 27.870 160.495 28.060 161.265 ;
        RECT 29.160 161.135 29.330 161.865 ;
        RECT 30.475 161.695 30.645 162.025 ;
        RECT 30.815 161.865 31.145 162.245 ;
        RECT 29.500 161.315 29.850 161.685 ;
        RECT 29.160 161.095 29.580 161.135 ;
        RECT 28.230 160.925 29.580 161.095 ;
        RECT 28.230 160.765 28.480 160.925 ;
        RECT 28.990 160.495 29.240 160.755 ;
        RECT 27.870 160.245 29.240 160.495 ;
        RECT 25.800 159.955 26.040 160.245 ;
        RECT 26.840 160.165 27.010 160.245 ;
        RECT 26.240 159.695 26.660 160.075 ;
        RECT 26.840 159.915 27.470 160.165 ;
        RECT 27.940 159.695 28.270 160.075 ;
        RECT 28.440 159.955 28.610 160.245 ;
        RECT 29.410 160.080 29.580 160.925 ;
        RECT 30.030 160.755 30.250 161.625 ;
        RECT 30.475 161.505 31.170 161.695 ;
        RECT 29.750 160.375 30.250 160.755 ;
        RECT 30.420 160.705 30.830 161.325 ;
        RECT 31.000 160.535 31.170 161.505 ;
        RECT 30.475 160.365 31.170 160.535 ;
        RECT 28.790 159.695 29.170 160.075 ;
        RECT 29.410 159.910 30.240 160.080 ;
        RECT 30.475 159.865 30.645 160.365 ;
        RECT 30.815 159.695 31.145 160.195 ;
        RECT 31.360 159.865 31.585 161.985 ;
        RECT 31.755 161.865 32.085 162.245 ;
        RECT 32.255 161.695 32.425 161.985 ;
        RECT 31.760 161.525 32.425 161.695 ;
        RECT 32.685 161.570 32.945 162.075 ;
        RECT 33.125 161.865 33.455 162.245 ;
        RECT 33.635 161.695 33.805 162.075 ;
        RECT 31.760 160.535 31.990 161.525 ;
        RECT 32.160 160.705 32.510 161.355 ;
        RECT 32.685 160.770 32.855 161.570 ;
        RECT 33.140 161.525 33.805 161.695 ;
        RECT 33.140 161.270 33.310 161.525 ;
        RECT 34.065 161.475 35.735 162.245 ;
        RECT 33.025 160.940 33.310 161.270 ;
        RECT 33.545 160.975 33.875 161.345 ;
        RECT 33.140 160.795 33.310 160.940 ;
        RECT 31.760 160.365 32.425 160.535 ;
        RECT 31.755 159.695 32.085 160.195 ;
        RECT 32.255 159.865 32.425 160.365 ;
        RECT 32.685 159.865 32.955 160.770 ;
        RECT 33.140 160.625 33.805 160.795 ;
        RECT 33.125 159.695 33.455 160.455 ;
        RECT 33.635 159.865 33.805 160.625 ;
        RECT 34.065 160.785 34.815 161.305 ;
        RECT 34.985 160.955 35.735 161.475 ;
        RECT 35.945 161.425 36.175 162.245 ;
        RECT 36.345 161.445 36.675 162.075 ;
        RECT 35.925 161.005 36.255 161.255 ;
        RECT 36.425 160.845 36.675 161.445 ;
        RECT 36.845 161.425 37.055 162.245 ;
        RECT 37.285 161.520 37.575 162.245 ;
        RECT 37.950 161.465 38.450 162.075 ;
        RECT 37.745 161.005 38.095 161.255 ;
        RECT 34.065 159.695 35.735 160.785 ;
        RECT 35.945 159.695 36.175 160.835 ;
        RECT 36.345 159.865 36.675 160.845 ;
        RECT 36.845 159.695 37.055 160.835 ;
        RECT 37.285 159.695 37.575 160.860 ;
        RECT 38.280 160.835 38.450 161.465 ;
        RECT 39.080 161.595 39.410 162.075 ;
        RECT 39.580 161.785 39.805 162.245 ;
        RECT 39.975 161.595 40.305 162.075 ;
        RECT 39.080 161.425 40.305 161.595 ;
        RECT 40.495 161.445 40.745 162.245 ;
        RECT 40.915 161.445 41.255 162.075 ;
        RECT 41.630 161.465 42.130 162.075 ;
        RECT 38.620 161.055 38.950 161.255 ;
        RECT 39.120 161.055 39.450 161.255 ;
        RECT 39.620 161.055 40.040 161.255 ;
        RECT 40.215 161.085 40.910 161.255 ;
        RECT 40.215 160.835 40.385 161.085 ;
        RECT 41.080 160.885 41.255 161.445 ;
        RECT 41.425 161.005 41.775 161.255 ;
        RECT 41.025 160.835 41.255 160.885 ;
        RECT 41.960 160.835 42.130 161.465 ;
        RECT 42.760 161.595 43.090 162.075 ;
        RECT 43.260 161.785 43.485 162.245 ;
        RECT 43.655 161.595 43.985 162.075 ;
        RECT 42.760 161.425 43.985 161.595 ;
        RECT 44.175 161.445 44.425 162.245 ;
        RECT 44.595 161.445 44.935 162.075 ;
        RECT 45.310 161.465 45.810 162.075 ;
        RECT 42.300 161.055 42.630 161.255 ;
        RECT 42.800 161.055 43.130 161.255 ;
        RECT 43.300 161.055 43.720 161.255 ;
        RECT 43.895 161.085 44.590 161.255 ;
        RECT 43.895 160.835 44.065 161.085 ;
        RECT 44.760 160.835 44.935 161.445 ;
        RECT 45.105 161.005 45.455 161.255 ;
        RECT 45.640 160.835 45.810 161.465 ;
        RECT 46.440 161.595 46.770 162.075 ;
        RECT 46.940 161.785 47.165 162.245 ;
        RECT 47.335 161.595 47.665 162.075 ;
        RECT 46.440 161.425 47.665 161.595 ;
        RECT 47.855 161.445 48.105 162.245 ;
        RECT 48.275 161.445 48.615 162.075 ;
        RECT 45.980 161.055 46.310 161.255 ;
        RECT 46.480 161.055 46.810 161.255 ;
        RECT 46.980 161.055 47.400 161.255 ;
        RECT 47.575 161.085 48.270 161.255 ;
        RECT 47.575 160.835 47.745 161.085 ;
        RECT 48.440 160.835 48.615 161.445 ;
        RECT 49.060 161.435 49.305 162.040 ;
        RECT 49.525 161.710 50.035 162.245 ;
        RECT 37.950 160.665 40.385 160.835 ;
        RECT 37.950 159.865 38.280 160.665 ;
        RECT 38.450 159.695 38.780 160.495 ;
        RECT 39.080 159.865 39.410 160.665 ;
        RECT 40.055 159.695 40.305 160.495 ;
        RECT 40.575 159.695 40.745 160.835 ;
        RECT 40.915 159.865 41.255 160.835 ;
        RECT 41.630 160.665 44.065 160.835 ;
        RECT 41.630 159.865 41.960 160.665 ;
        RECT 42.130 159.695 42.460 160.495 ;
        RECT 42.760 159.865 43.090 160.665 ;
        RECT 43.735 159.695 43.985 160.495 ;
        RECT 44.255 159.695 44.425 160.835 ;
        RECT 44.595 159.865 44.935 160.835 ;
        RECT 45.310 160.665 47.745 160.835 ;
        RECT 45.310 159.865 45.640 160.665 ;
        RECT 45.810 159.695 46.140 160.495 ;
        RECT 46.440 159.865 46.770 160.665 ;
        RECT 47.415 159.695 47.665 160.495 ;
        RECT 47.935 159.695 48.105 160.835 ;
        RECT 48.275 159.865 48.615 160.835 ;
        RECT 48.785 161.265 50.015 161.435 ;
        RECT 48.785 160.455 49.125 161.265 ;
        RECT 49.295 160.700 50.045 160.890 ;
        RECT 48.785 160.045 49.300 160.455 ;
        RECT 49.535 159.695 49.705 160.455 ;
        RECT 49.875 160.035 50.045 160.700 ;
        RECT 50.215 160.715 50.405 162.075 ;
        RECT 50.575 161.225 50.850 162.075 ;
        RECT 51.040 161.710 51.570 162.075 ;
        RECT 51.995 161.845 52.325 162.245 ;
        RECT 51.395 161.675 51.570 161.710 ;
        RECT 50.575 161.055 50.855 161.225 ;
        RECT 50.575 160.915 50.850 161.055 ;
        RECT 51.055 160.715 51.225 161.515 ;
        RECT 50.215 160.545 51.225 160.715 ;
        RECT 51.395 161.505 52.325 161.675 ;
        RECT 52.495 161.505 52.750 162.075 ;
        RECT 53.390 161.700 58.735 162.245 ;
        RECT 51.395 160.375 51.565 161.505 ;
        RECT 52.155 161.335 52.325 161.505 ;
        RECT 50.440 160.205 51.565 160.375 ;
        RECT 51.735 161.005 51.930 161.335 ;
        RECT 52.155 161.005 52.410 161.335 ;
        RECT 51.735 160.035 51.905 161.005 ;
        RECT 52.580 160.835 52.750 161.505 ;
        RECT 49.875 159.865 51.905 160.035 ;
        RECT 52.075 159.695 52.245 160.835 ;
        RECT 52.415 159.865 52.750 160.835 ;
        RECT 54.980 160.130 55.330 161.380 ;
        RECT 56.810 160.870 57.150 161.700 ;
        RECT 59.180 161.435 59.425 162.040 ;
        RECT 59.645 161.710 60.155 162.245 ;
        RECT 58.905 161.265 60.135 161.435 ;
        RECT 58.905 160.455 59.245 161.265 ;
        RECT 59.415 160.700 60.165 160.890 ;
        RECT 53.390 159.695 58.735 160.130 ;
        RECT 58.905 160.045 59.420 160.455 ;
        RECT 59.655 159.695 59.825 160.455 ;
        RECT 59.995 160.035 60.165 160.700 ;
        RECT 60.335 160.715 60.525 162.075 ;
        RECT 60.695 161.225 60.970 162.075 ;
        RECT 61.160 161.710 61.690 162.075 ;
        RECT 62.115 161.845 62.445 162.245 ;
        RECT 61.515 161.675 61.690 161.710 ;
        RECT 60.695 161.055 60.975 161.225 ;
        RECT 60.695 160.915 60.970 161.055 ;
        RECT 61.175 160.715 61.345 161.515 ;
        RECT 60.335 160.545 61.345 160.715 ;
        RECT 61.515 161.505 62.445 161.675 ;
        RECT 62.615 161.505 62.870 162.075 ;
        RECT 63.045 161.520 63.335 162.245 ;
        RECT 61.515 160.375 61.685 161.505 ;
        RECT 62.275 161.335 62.445 161.505 ;
        RECT 60.560 160.205 61.685 160.375 ;
        RECT 61.855 161.005 62.050 161.335 ;
        RECT 62.275 161.005 62.530 161.335 ;
        RECT 61.855 160.035 62.025 161.005 ;
        RECT 62.700 160.835 62.870 161.505 ;
        RECT 63.965 161.475 65.635 162.245 ;
        RECT 59.995 159.865 62.025 160.035 ;
        RECT 62.195 159.695 62.365 160.835 ;
        RECT 62.535 159.865 62.870 160.835 ;
        RECT 63.045 159.695 63.335 160.860 ;
        RECT 63.965 160.785 64.715 161.305 ;
        RECT 64.885 160.955 65.635 161.475 ;
        RECT 65.845 161.425 66.075 162.245 ;
        RECT 66.245 161.445 66.575 162.075 ;
        RECT 65.825 161.005 66.155 161.255 ;
        RECT 66.325 160.845 66.575 161.445 ;
        RECT 66.745 161.425 66.955 162.245 ;
        RECT 67.185 161.475 68.855 162.245 ;
        RECT 63.965 159.695 65.635 160.785 ;
        RECT 65.845 159.695 66.075 160.835 ;
        RECT 66.245 159.865 66.575 160.845 ;
        RECT 66.745 159.695 66.955 160.835 ;
        RECT 67.185 160.785 67.935 161.305 ;
        RECT 68.105 160.955 68.855 161.475 ;
        RECT 69.030 161.405 69.290 162.245 ;
        RECT 69.465 161.500 69.720 162.075 ;
        RECT 69.890 161.865 70.220 162.245 ;
        RECT 70.435 161.695 70.605 162.075 ;
        RECT 69.890 161.525 70.605 161.695 ;
        RECT 67.185 159.695 68.855 160.785 ;
        RECT 69.030 159.695 69.290 160.845 ;
        RECT 69.465 160.770 69.635 161.500 ;
        RECT 69.890 161.335 70.060 161.525 ;
        RECT 70.870 161.405 71.130 162.245 ;
        RECT 71.305 161.500 71.560 162.075 ;
        RECT 71.730 161.865 72.060 162.245 ;
        RECT 72.275 161.695 72.445 162.075 ;
        RECT 71.730 161.525 72.445 161.695 ;
        RECT 72.795 161.695 72.965 162.075 ;
        RECT 73.180 161.865 73.510 162.245 ;
        RECT 72.795 161.525 73.510 161.695 ;
        RECT 69.805 161.005 70.060 161.335 ;
        RECT 69.890 160.795 70.060 161.005 ;
        RECT 70.340 160.975 70.695 161.345 ;
        RECT 69.465 159.865 69.720 160.770 ;
        RECT 69.890 160.625 70.605 160.795 ;
        RECT 69.890 159.695 70.220 160.455 ;
        RECT 70.435 159.865 70.605 160.625 ;
        RECT 70.870 159.695 71.130 160.845 ;
        RECT 71.305 160.770 71.475 161.500 ;
        RECT 71.730 161.335 71.900 161.525 ;
        RECT 71.645 161.005 71.900 161.335 ;
        RECT 71.730 160.795 71.900 161.005 ;
        RECT 72.180 160.975 72.535 161.345 ;
        RECT 72.705 160.975 73.060 161.345 ;
        RECT 73.340 161.335 73.510 161.525 ;
        RECT 73.680 161.500 73.935 162.075 ;
        RECT 73.340 161.005 73.595 161.335 ;
        RECT 73.340 160.795 73.510 161.005 ;
        RECT 71.305 159.865 71.560 160.770 ;
        RECT 71.730 160.625 72.445 160.795 ;
        RECT 71.730 159.695 72.060 160.455 ;
        RECT 72.275 159.865 72.445 160.625 ;
        RECT 72.795 160.625 73.510 160.795 ;
        RECT 73.765 160.770 73.935 161.500 ;
        RECT 74.110 161.405 74.370 162.245 ;
        RECT 74.550 161.405 74.810 162.245 ;
        RECT 74.985 161.500 75.240 162.075 ;
        RECT 75.410 161.865 75.740 162.245 ;
        RECT 75.955 161.695 76.125 162.075 ;
        RECT 75.410 161.525 76.125 161.695 ;
        RECT 72.795 159.865 72.965 160.625 ;
        RECT 73.180 159.695 73.510 160.455 ;
        RECT 73.680 159.865 73.935 160.770 ;
        RECT 74.110 159.695 74.370 160.845 ;
        RECT 74.550 159.695 74.810 160.845 ;
        RECT 74.985 160.770 75.155 161.500 ;
        RECT 75.410 161.335 75.580 161.525 ;
        RECT 77.305 161.475 80.815 162.245 ;
        RECT 75.325 161.005 75.580 161.335 ;
        RECT 75.410 160.795 75.580 161.005 ;
        RECT 75.860 160.975 76.215 161.345 ;
        RECT 74.985 159.865 75.240 160.770 ;
        RECT 75.410 160.625 76.125 160.795 ;
        RECT 75.410 159.695 75.740 160.455 ;
        RECT 75.955 159.865 76.125 160.625 ;
        RECT 77.305 160.785 78.995 161.305 ;
        RECT 79.165 160.955 80.815 161.475 ;
        RECT 80.985 161.445 81.325 162.075 ;
        RECT 81.495 161.445 81.745 162.245 ;
        RECT 81.935 161.595 82.265 162.075 ;
        RECT 82.435 161.785 82.660 162.245 ;
        RECT 82.830 161.595 83.160 162.075 ;
        RECT 80.985 160.835 81.160 161.445 ;
        RECT 81.935 161.425 83.160 161.595 ;
        RECT 83.790 161.465 84.290 162.075 ;
        RECT 85.125 161.475 88.635 162.245 ;
        RECT 88.805 161.520 89.095 162.245 ;
        RECT 89.725 161.475 91.395 162.245 ;
        RECT 91.570 161.700 96.915 162.245 ;
        RECT 97.090 161.700 102.435 162.245 ;
        RECT 81.330 161.085 82.025 161.255 ;
        RECT 81.855 160.835 82.025 161.085 ;
        RECT 82.200 161.055 82.620 161.255 ;
        RECT 82.790 161.055 83.120 161.255 ;
        RECT 83.290 161.055 83.620 161.255 ;
        RECT 83.790 160.835 83.960 161.465 ;
        RECT 84.145 161.005 84.495 161.255 ;
        RECT 77.305 159.695 80.815 160.785 ;
        RECT 80.985 159.865 81.325 160.835 ;
        RECT 81.495 159.695 81.665 160.835 ;
        RECT 81.855 160.665 84.290 160.835 ;
        RECT 81.935 159.695 82.185 160.495 ;
        RECT 82.830 159.865 83.160 160.665 ;
        RECT 83.460 159.695 83.790 160.495 ;
        RECT 83.960 159.865 84.290 160.665 ;
        RECT 85.125 160.785 86.815 161.305 ;
        RECT 86.985 160.955 88.635 161.475 ;
        RECT 85.125 159.695 88.635 160.785 ;
        RECT 88.805 159.695 89.095 160.860 ;
        RECT 89.725 160.785 90.475 161.305 ;
        RECT 90.645 160.955 91.395 161.475 ;
        RECT 89.725 159.695 91.395 160.785 ;
        RECT 93.160 160.130 93.510 161.380 ;
        RECT 94.990 160.870 95.330 161.700 ;
        RECT 98.680 160.130 99.030 161.380 ;
        RECT 100.510 160.870 100.850 161.700 ;
        RECT 102.695 161.695 102.865 162.075 ;
        RECT 103.045 161.865 103.375 162.245 ;
        RECT 102.695 161.525 103.360 161.695 ;
        RECT 103.555 161.570 103.815 162.075 ;
        RECT 102.625 160.975 102.955 161.345 ;
        RECT 103.190 161.270 103.360 161.525 ;
        RECT 103.190 160.940 103.475 161.270 ;
        RECT 103.190 160.795 103.360 160.940 ;
        RECT 102.695 160.625 103.360 160.795 ;
        RECT 103.645 160.770 103.815 161.570 ;
        RECT 91.570 159.695 96.915 160.130 ;
        RECT 97.090 159.695 102.435 160.130 ;
        RECT 102.695 159.865 102.865 160.625 ;
        RECT 103.045 159.695 103.375 160.455 ;
        RECT 103.545 159.865 103.815 160.770 ;
        RECT 103.990 161.505 104.245 162.075 ;
        RECT 104.415 161.845 104.745 162.245 ;
        RECT 105.170 161.710 105.700 162.075 ;
        RECT 105.890 161.905 106.165 162.075 ;
        RECT 105.885 161.735 106.165 161.905 ;
        RECT 105.170 161.675 105.345 161.710 ;
        RECT 104.415 161.505 105.345 161.675 ;
        RECT 103.990 160.835 104.160 161.505 ;
        RECT 104.415 161.335 104.585 161.505 ;
        RECT 104.330 161.005 104.585 161.335 ;
        RECT 104.810 161.005 105.005 161.335 ;
        RECT 103.990 159.865 104.325 160.835 ;
        RECT 104.495 159.695 104.665 160.835 ;
        RECT 104.835 160.035 105.005 161.005 ;
        RECT 105.175 160.375 105.345 161.505 ;
        RECT 105.515 160.715 105.685 161.515 ;
        RECT 105.890 160.915 106.165 161.735 ;
        RECT 106.335 160.715 106.525 162.075 ;
        RECT 106.705 161.710 107.215 162.245 ;
        RECT 107.435 161.435 107.680 162.040 ;
        RECT 109.050 161.700 114.395 162.245 ;
        RECT 106.725 161.265 107.955 161.435 ;
        RECT 105.515 160.545 106.525 160.715 ;
        RECT 106.695 160.700 107.445 160.890 ;
        RECT 105.175 160.205 106.300 160.375 ;
        RECT 106.695 160.035 106.865 160.700 ;
        RECT 107.615 160.455 107.955 161.265 ;
        RECT 104.835 159.865 106.865 160.035 ;
        RECT 107.035 159.695 107.205 160.455 ;
        RECT 107.440 160.045 107.955 160.455 ;
        RECT 110.640 160.130 110.990 161.380 ;
        RECT 112.470 160.870 112.810 161.700 ;
        RECT 114.565 161.520 114.855 162.245 ;
        RECT 115.025 161.495 116.235 162.245 ;
        RECT 109.050 159.695 114.395 160.130 ;
        RECT 114.565 159.695 114.855 160.860 ;
        RECT 115.025 160.785 115.545 161.325 ;
        RECT 115.715 160.955 116.235 161.495 ;
        RECT 116.495 161.595 116.665 162.075 ;
        RECT 116.845 161.765 117.085 162.245 ;
        RECT 117.335 161.595 117.505 162.075 ;
        RECT 117.675 161.765 118.005 162.245 ;
        RECT 118.175 161.595 118.345 162.075 ;
        RECT 116.495 161.425 117.130 161.595 ;
        RECT 117.335 161.425 118.345 161.595 ;
        RECT 118.515 161.445 118.845 162.245 ;
        RECT 119.165 161.475 120.835 162.245 ;
        RECT 121.010 161.700 126.355 162.245 ;
        RECT 116.960 161.255 117.130 161.425 ;
        RECT 116.410 161.015 116.790 161.255 ;
        RECT 116.960 161.085 117.460 161.255 ;
        RECT 116.960 160.845 117.130 161.085 ;
        RECT 117.850 160.885 118.345 161.425 ;
        RECT 115.025 159.695 116.235 160.785 ;
        RECT 116.415 160.675 117.130 160.845 ;
        RECT 117.335 160.715 118.345 160.885 ;
        RECT 116.415 159.865 116.745 160.675 ;
        RECT 116.915 159.695 117.155 160.495 ;
        RECT 117.335 159.865 117.505 160.715 ;
        RECT 117.675 159.695 118.005 160.495 ;
        RECT 118.175 159.865 118.345 160.715 ;
        RECT 118.515 159.695 118.845 160.845 ;
        RECT 119.165 160.785 119.915 161.305 ;
        RECT 120.085 160.955 120.835 161.475 ;
        RECT 119.165 159.695 120.835 160.785 ;
        RECT 122.600 160.130 122.950 161.380 ;
        RECT 124.430 160.870 124.770 161.700 ;
        RECT 126.525 161.495 127.735 162.245 ;
        RECT 126.525 160.785 127.045 161.325 ;
        RECT 127.215 160.955 127.735 161.495 ;
        RECT 121.010 159.695 126.355 160.130 ;
        RECT 126.525 159.695 127.735 160.785 ;
        RECT 20.640 159.525 127.820 159.695 ;
        RECT 20.725 158.435 21.935 159.525 ;
        RECT 20.725 157.725 21.245 158.265 ;
        RECT 21.415 157.895 21.935 158.435 ;
        RECT 22.565 158.435 24.235 159.525 ;
        RECT 22.565 157.915 23.315 158.435 ;
        RECT 24.405 158.360 24.695 159.525 ;
        RECT 25.845 158.385 26.055 159.525 ;
        RECT 26.225 158.375 26.555 159.355 ;
        RECT 26.725 158.385 26.955 159.525 ;
        RECT 27.165 158.765 27.680 159.175 ;
        RECT 27.915 158.765 28.085 159.525 ;
        RECT 28.255 159.185 30.285 159.355 ;
        RECT 23.485 157.745 24.235 158.265 ;
        RECT 20.725 156.975 21.935 157.725 ;
        RECT 22.565 156.975 24.235 157.745 ;
        RECT 24.405 156.975 24.695 157.700 ;
        RECT 25.845 156.975 26.055 157.795 ;
        RECT 26.225 157.775 26.475 158.375 ;
        RECT 26.645 157.965 26.975 158.215 ;
        RECT 27.165 157.955 27.505 158.765 ;
        RECT 28.255 158.520 28.425 159.185 ;
        RECT 28.820 158.845 29.945 159.015 ;
        RECT 27.675 158.330 28.425 158.520 ;
        RECT 28.595 158.505 29.605 158.675 ;
        RECT 26.225 157.145 26.555 157.775 ;
        RECT 26.725 156.975 26.955 157.795 ;
        RECT 27.165 157.785 28.395 157.955 ;
        RECT 27.440 157.180 27.685 157.785 ;
        RECT 27.905 156.975 28.415 157.510 ;
        RECT 28.595 157.145 28.785 158.505 ;
        RECT 28.955 157.485 29.230 158.305 ;
        RECT 29.435 157.705 29.605 158.505 ;
        RECT 29.775 157.715 29.945 158.845 ;
        RECT 30.115 158.215 30.285 159.185 ;
        RECT 30.455 158.385 30.625 159.525 ;
        RECT 30.795 158.385 31.130 159.355 ;
        RECT 30.115 157.885 30.310 158.215 ;
        RECT 30.535 157.885 30.790 158.215 ;
        RECT 30.535 157.715 30.705 157.885 ;
        RECT 30.960 157.715 31.130 158.385 ;
        RECT 31.305 158.435 33.895 159.525 ;
        RECT 34.440 159.185 34.695 159.215 ;
        RECT 34.355 159.015 34.695 159.185 ;
        RECT 34.440 158.545 34.695 159.015 ;
        RECT 34.875 158.725 35.160 159.525 ;
        RECT 35.340 158.805 35.670 159.315 ;
        RECT 31.305 157.915 32.515 158.435 ;
        RECT 32.685 157.745 33.895 158.265 ;
        RECT 29.775 157.545 30.705 157.715 ;
        RECT 29.775 157.510 29.950 157.545 ;
        RECT 28.955 157.315 29.235 157.485 ;
        RECT 28.955 157.145 29.230 157.315 ;
        RECT 29.420 157.145 29.950 157.510 ;
        RECT 30.375 156.975 30.705 157.375 ;
        RECT 30.875 157.145 31.130 157.715 ;
        RECT 31.305 156.975 33.895 157.745 ;
        RECT 34.440 157.685 34.620 158.545 ;
        RECT 35.340 158.215 35.590 158.805 ;
        RECT 35.940 158.655 36.110 159.265 ;
        RECT 36.280 158.835 36.610 159.525 ;
        RECT 36.840 158.975 37.080 159.265 ;
        RECT 37.280 159.145 37.700 159.525 ;
        RECT 37.880 159.055 38.510 159.305 ;
        RECT 38.980 159.145 39.310 159.525 ;
        RECT 37.880 158.975 38.050 159.055 ;
        RECT 39.480 158.975 39.650 159.265 ;
        RECT 39.830 159.145 40.210 159.525 ;
        RECT 40.450 159.140 41.280 159.310 ;
        RECT 36.840 158.805 38.050 158.975 ;
        RECT 34.790 157.885 35.590 158.215 ;
        RECT 34.440 157.155 34.695 157.685 ;
        RECT 34.875 156.975 35.160 157.435 ;
        RECT 35.340 157.235 35.590 157.885 ;
        RECT 35.790 158.635 36.110 158.655 ;
        RECT 35.790 158.465 37.710 158.635 ;
        RECT 35.790 157.570 35.980 158.465 ;
        RECT 37.880 158.295 38.050 158.805 ;
        RECT 38.220 158.545 38.740 158.855 ;
        RECT 36.150 158.125 38.050 158.295 ;
        RECT 36.150 158.065 36.480 158.125 ;
        RECT 36.630 157.895 36.960 157.955 ;
        RECT 36.300 157.625 36.960 157.895 ;
        RECT 35.790 157.240 36.110 157.570 ;
        RECT 36.290 156.975 36.950 157.455 ;
        RECT 37.150 157.365 37.320 158.125 ;
        RECT 38.220 157.955 38.400 158.365 ;
        RECT 37.490 157.785 37.820 157.905 ;
        RECT 38.570 157.785 38.740 158.545 ;
        RECT 37.490 157.615 38.740 157.785 ;
        RECT 38.910 158.725 40.280 158.975 ;
        RECT 38.910 157.955 39.100 158.725 ;
        RECT 40.030 158.465 40.280 158.725 ;
        RECT 39.270 158.295 39.520 158.455 ;
        RECT 40.450 158.295 40.620 159.140 ;
        RECT 41.515 158.855 41.685 159.355 ;
        RECT 41.855 159.025 42.185 159.525 ;
        RECT 40.790 158.465 41.290 158.845 ;
        RECT 41.515 158.685 42.210 158.855 ;
        RECT 39.270 158.125 40.620 158.295 ;
        RECT 40.200 158.085 40.620 158.125 ;
        RECT 38.910 157.615 39.330 157.955 ;
        RECT 39.620 157.625 40.030 157.955 ;
        RECT 37.150 157.195 38.000 157.365 ;
        RECT 38.560 156.975 38.880 157.435 ;
        RECT 39.080 157.185 39.330 157.615 ;
        RECT 39.620 156.975 40.030 157.415 ;
        RECT 40.200 157.355 40.370 158.085 ;
        RECT 40.540 157.535 40.890 157.905 ;
        RECT 41.070 157.595 41.290 158.465 ;
        RECT 41.460 157.895 41.870 158.515 ;
        RECT 42.040 157.715 42.210 158.685 ;
        RECT 41.515 157.525 42.210 157.715 ;
        RECT 40.200 157.155 41.215 157.355 ;
        RECT 41.515 157.195 41.685 157.525 ;
        RECT 41.855 156.975 42.185 157.355 ;
        RECT 42.400 157.235 42.625 159.355 ;
        RECT 42.795 159.025 43.125 159.525 ;
        RECT 43.295 158.855 43.465 159.355 ;
        RECT 42.800 158.685 43.465 158.855 ;
        RECT 42.800 157.695 43.030 158.685 ;
        RECT 43.200 157.865 43.550 158.515 ;
        RECT 43.725 158.435 46.315 159.525 ;
        RECT 46.690 158.555 47.020 159.355 ;
        RECT 47.190 158.725 47.520 159.525 ;
        RECT 47.820 158.555 48.150 159.355 ;
        RECT 48.795 158.725 49.045 159.525 ;
        RECT 43.725 157.915 44.935 158.435 ;
        RECT 46.690 158.385 49.125 158.555 ;
        RECT 49.315 158.385 49.485 159.525 ;
        RECT 49.655 158.385 49.995 159.355 ;
        RECT 45.105 157.745 46.315 158.265 ;
        RECT 46.485 157.965 46.835 158.215 ;
        RECT 47.020 157.755 47.190 158.385 ;
        RECT 47.360 157.965 47.690 158.165 ;
        RECT 47.860 157.965 48.190 158.165 ;
        RECT 48.360 157.965 48.780 158.165 ;
        RECT 48.955 158.135 49.125 158.385 ;
        RECT 48.955 157.965 49.650 158.135 ;
        RECT 42.800 157.525 43.465 157.695 ;
        RECT 42.795 156.975 43.125 157.355 ;
        RECT 43.295 157.235 43.465 157.525 ;
        RECT 43.725 156.975 46.315 157.745 ;
        RECT 46.690 157.145 47.190 157.755 ;
        RECT 47.820 157.625 49.045 157.795 ;
        RECT 49.820 157.775 49.995 158.385 ;
        RECT 50.165 158.360 50.455 159.525 ;
        RECT 50.625 158.385 50.965 159.355 ;
        RECT 51.135 158.385 51.305 159.525 ;
        RECT 51.575 158.725 51.825 159.525 ;
        RECT 52.470 158.555 52.800 159.355 ;
        RECT 53.100 158.725 53.430 159.525 ;
        RECT 53.600 158.555 53.930 159.355 ;
        RECT 51.495 158.385 53.930 158.555 ;
        RECT 54.765 158.435 57.355 159.525 ;
        RECT 47.820 157.145 48.150 157.625 ;
        RECT 48.320 156.975 48.545 157.435 ;
        RECT 48.715 157.145 49.045 157.625 ;
        RECT 49.235 156.975 49.485 157.775 ;
        RECT 49.655 157.145 49.995 157.775 ;
        RECT 50.625 157.775 50.800 158.385 ;
        RECT 51.495 158.135 51.665 158.385 ;
        RECT 50.970 157.965 51.665 158.135 ;
        RECT 51.840 157.965 52.260 158.165 ;
        RECT 52.430 157.965 52.760 158.165 ;
        RECT 52.930 157.965 53.260 158.165 ;
        RECT 50.165 156.975 50.455 157.700 ;
        RECT 50.625 157.145 50.965 157.775 ;
        RECT 51.135 156.975 51.385 157.775 ;
        RECT 51.575 157.625 52.800 157.795 ;
        RECT 51.575 157.145 51.905 157.625 ;
        RECT 52.075 156.975 52.300 157.435 ;
        RECT 52.470 157.145 52.800 157.625 ;
        RECT 53.430 157.755 53.600 158.385 ;
        RECT 53.785 157.965 54.135 158.215 ;
        RECT 54.765 157.915 55.975 158.435 ;
        RECT 57.585 158.385 57.795 159.525 ;
        RECT 57.965 158.375 58.295 159.355 ;
        RECT 58.465 158.385 58.695 159.525 ;
        RECT 58.905 158.765 59.420 159.175 ;
        RECT 59.655 158.765 59.825 159.525 ;
        RECT 59.995 159.185 62.025 159.355 ;
        RECT 53.430 157.145 53.930 157.755 ;
        RECT 56.145 157.745 57.355 158.265 ;
        RECT 54.765 156.975 57.355 157.745 ;
        RECT 57.585 156.975 57.795 157.795 ;
        RECT 57.965 157.775 58.215 158.375 ;
        RECT 58.385 157.965 58.715 158.215 ;
        RECT 58.905 157.955 59.245 158.765 ;
        RECT 59.995 158.520 60.165 159.185 ;
        RECT 60.560 158.845 61.685 159.015 ;
        RECT 59.415 158.330 60.165 158.520 ;
        RECT 60.335 158.505 61.345 158.675 ;
        RECT 57.965 157.145 58.295 157.775 ;
        RECT 58.465 156.975 58.695 157.795 ;
        RECT 58.905 157.785 60.135 157.955 ;
        RECT 59.180 157.180 59.425 157.785 ;
        RECT 59.645 156.975 60.155 157.510 ;
        RECT 60.335 157.145 60.525 158.505 ;
        RECT 60.695 157.825 60.970 158.305 ;
        RECT 60.695 157.655 60.975 157.825 ;
        RECT 61.175 157.705 61.345 158.505 ;
        RECT 61.515 157.715 61.685 158.845 ;
        RECT 61.855 158.215 62.025 159.185 ;
        RECT 62.195 158.385 62.365 159.525 ;
        RECT 62.535 158.385 62.870 159.355 ;
        RECT 61.855 157.885 62.050 158.215 ;
        RECT 62.275 157.885 62.530 158.215 ;
        RECT 62.275 157.715 62.445 157.885 ;
        RECT 62.700 157.715 62.870 158.385 ;
        RECT 63.420 158.545 63.675 159.215 ;
        RECT 63.855 158.725 64.140 159.525 ;
        RECT 64.320 158.805 64.650 159.315 ;
        RECT 63.420 157.825 63.600 158.545 ;
        RECT 64.320 158.215 64.570 158.805 ;
        RECT 64.920 158.655 65.090 159.265 ;
        RECT 65.260 158.835 65.590 159.525 ;
        RECT 65.820 158.975 66.060 159.265 ;
        RECT 66.260 159.145 66.680 159.525 ;
        RECT 66.860 159.055 67.490 159.305 ;
        RECT 67.960 159.145 68.290 159.525 ;
        RECT 66.860 158.975 67.030 159.055 ;
        RECT 68.460 158.975 68.630 159.265 ;
        RECT 68.810 159.145 69.190 159.525 ;
        RECT 69.430 159.140 70.260 159.310 ;
        RECT 65.820 158.805 67.030 158.975 ;
        RECT 63.770 157.885 64.570 158.215 ;
        RECT 60.695 157.145 60.970 157.655 ;
        RECT 61.515 157.545 62.445 157.715 ;
        RECT 61.515 157.510 61.690 157.545 ;
        RECT 61.160 157.145 61.690 157.510 ;
        RECT 62.115 156.975 62.445 157.375 ;
        RECT 62.615 157.145 62.870 157.715 ;
        RECT 63.335 157.685 63.600 157.825 ;
        RECT 63.335 157.655 63.675 157.685 ;
        RECT 63.420 157.155 63.675 157.655 ;
        RECT 63.855 156.975 64.140 157.435 ;
        RECT 64.320 157.235 64.570 157.885 ;
        RECT 64.770 158.635 65.090 158.655 ;
        RECT 64.770 158.465 66.690 158.635 ;
        RECT 64.770 157.570 64.960 158.465 ;
        RECT 66.860 158.295 67.030 158.805 ;
        RECT 67.200 158.545 67.720 158.855 ;
        RECT 65.130 158.125 67.030 158.295 ;
        RECT 65.130 158.065 65.460 158.125 ;
        RECT 65.610 157.895 65.940 157.955 ;
        RECT 65.280 157.625 65.940 157.895 ;
        RECT 64.770 157.240 65.090 157.570 ;
        RECT 65.270 156.975 65.930 157.455 ;
        RECT 66.130 157.365 66.300 158.125 ;
        RECT 67.200 157.955 67.380 158.365 ;
        RECT 66.470 157.785 66.800 157.905 ;
        RECT 67.550 157.785 67.720 158.545 ;
        RECT 66.470 157.615 67.720 157.785 ;
        RECT 67.890 158.725 69.260 158.975 ;
        RECT 67.890 157.955 68.080 158.725 ;
        RECT 69.010 158.465 69.260 158.725 ;
        RECT 68.250 158.295 68.500 158.455 ;
        RECT 69.430 158.295 69.600 159.140 ;
        RECT 70.495 158.855 70.665 159.355 ;
        RECT 70.835 159.025 71.165 159.525 ;
        RECT 69.770 158.465 70.270 158.845 ;
        RECT 70.495 158.685 71.190 158.855 ;
        RECT 68.250 158.125 69.600 158.295 ;
        RECT 69.180 158.085 69.600 158.125 ;
        RECT 67.890 157.615 68.310 157.955 ;
        RECT 68.600 157.625 69.010 157.955 ;
        RECT 66.130 157.195 66.980 157.365 ;
        RECT 67.540 156.975 67.860 157.435 ;
        RECT 68.060 157.185 68.310 157.615 ;
        RECT 68.600 156.975 69.010 157.415 ;
        RECT 69.180 157.355 69.350 158.085 ;
        RECT 69.520 157.535 69.870 157.905 ;
        RECT 70.050 157.595 70.270 158.465 ;
        RECT 70.440 157.895 70.850 158.515 ;
        RECT 71.020 157.715 71.190 158.685 ;
        RECT 70.495 157.525 71.190 157.715 ;
        RECT 69.180 157.155 70.195 157.355 ;
        RECT 70.495 157.195 70.665 157.525 ;
        RECT 70.835 156.975 71.165 157.355 ;
        RECT 71.380 157.235 71.605 159.355 ;
        RECT 71.775 159.025 72.105 159.525 ;
        RECT 72.275 158.855 72.445 159.355 ;
        RECT 71.780 158.685 72.445 158.855 ;
        RECT 71.780 157.695 72.010 158.685 ;
        RECT 72.180 157.865 72.530 158.515 ;
        RECT 73.175 158.465 73.505 159.525 ;
        RECT 73.685 158.215 73.855 159.185 ;
        RECT 74.025 158.935 74.355 159.335 ;
        RECT 74.525 159.165 74.855 159.525 ;
        RECT 75.055 158.935 75.755 159.355 ;
        RECT 74.025 158.705 75.755 158.935 ;
        RECT 74.025 158.485 74.355 158.705 ;
        RECT 74.550 158.215 74.875 158.505 ;
        RECT 73.165 157.885 73.475 158.215 ;
        RECT 73.685 157.885 74.060 158.215 ;
        RECT 74.380 157.885 74.875 158.215 ;
        RECT 75.050 157.965 75.380 158.505 ;
        RECT 75.550 157.735 75.755 158.705 ;
        RECT 75.925 158.360 76.215 159.525 ;
        RECT 77.305 158.385 77.645 159.355 ;
        RECT 77.815 158.385 77.985 159.525 ;
        RECT 78.255 158.725 78.505 159.525 ;
        RECT 79.150 158.555 79.480 159.355 ;
        RECT 79.780 158.725 80.110 159.525 ;
        RECT 80.280 158.555 80.610 159.355 ;
        RECT 78.175 158.385 80.610 158.555 ;
        RECT 80.985 158.385 81.325 159.355 ;
        RECT 81.495 158.385 81.665 159.525 ;
        RECT 81.935 158.725 82.185 159.525 ;
        RECT 82.830 158.555 83.160 159.355 ;
        RECT 83.460 158.725 83.790 159.525 ;
        RECT 83.960 158.555 84.290 159.355 ;
        RECT 81.855 158.385 84.290 158.555 ;
        RECT 84.665 158.435 87.255 159.525 ;
        RECT 87.430 159.090 92.775 159.525 ;
        RECT 71.780 157.525 72.445 157.695 ;
        RECT 71.775 156.975 72.105 157.355 ;
        RECT 72.275 157.235 72.445 157.525 ;
        RECT 73.175 157.505 74.535 157.715 ;
        RECT 73.175 157.145 73.505 157.505 ;
        RECT 73.675 156.975 74.005 157.335 ;
        RECT 74.205 157.145 74.535 157.505 ;
        RECT 75.045 157.145 75.755 157.735 ;
        RECT 77.305 157.775 77.480 158.385 ;
        RECT 78.175 158.135 78.345 158.385 ;
        RECT 77.650 157.965 78.345 158.135 ;
        RECT 78.520 157.965 78.940 158.165 ;
        RECT 79.110 157.965 79.440 158.165 ;
        RECT 79.610 157.965 79.940 158.165 ;
        RECT 75.925 156.975 76.215 157.700 ;
        RECT 77.305 157.145 77.645 157.775 ;
        RECT 77.815 156.975 78.065 157.775 ;
        RECT 78.255 157.625 79.480 157.795 ;
        RECT 78.255 157.145 78.585 157.625 ;
        RECT 78.755 156.975 78.980 157.435 ;
        RECT 79.150 157.145 79.480 157.625 ;
        RECT 80.110 157.755 80.280 158.385 ;
        RECT 80.465 157.965 80.815 158.215 ;
        RECT 80.985 157.775 81.160 158.385 ;
        RECT 81.855 158.135 82.025 158.385 ;
        RECT 81.330 157.965 82.025 158.135 ;
        RECT 82.200 157.965 82.620 158.165 ;
        RECT 82.790 157.965 83.120 158.165 ;
        RECT 83.290 157.965 83.620 158.165 ;
        RECT 80.110 157.145 80.610 157.755 ;
        RECT 80.985 157.145 81.325 157.775 ;
        RECT 81.495 156.975 81.745 157.775 ;
        RECT 81.935 157.625 83.160 157.795 ;
        RECT 81.935 157.145 82.265 157.625 ;
        RECT 82.435 156.975 82.660 157.435 ;
        RECT 82.830 157.145 83.160 157.625 ;
        RECT 83.790 157.755 83.960 158.385 ;
        RECT 84.145 157.965 84.495 158.215 ;
        RECT 84.665 157.915 85.875 158.435 ;
        RECT 83.790 157.145 84.290 157.755 ;
        RECT 86.045 157.745 87.255 158.265 ;
        RECT 89.020 157.840 89.370 159.090 ;
        RECT 93.005 158.385 93.215 159.525 ;
        RECT 93.385 158.375 93.715 159.355 ;
        RECT 93.885 158.385 94.115 159.525 ;
        RECT 94.325 158.435 95.995 159.525 ;
        RECT 96.170 159.090 101.515 159.525 ;
        RECT 84.665 156.975 87.255 157.745 ;
        RECT 90.850 157.520 91.190 158.350 ;
        RECT 87.430 156.975 92.775 157.520 ;
        RECT 93.005 156.975 93.215 157.795 ;
        RECT 93.385 157.775 93.635 158.375 ;
        RECT 93.805 157.965 94.135 158.215 ;
        RECT 94.325 157.915 95.075 158.435 ;
        RECT 93.385 157.145 93.715 157.775 ;
        RECT 93.885 156.975 94.115 157.795 ;
        RECT 95.245 157.745 95.995 158.265 ;
        RECT 97.760 157.840 98.110 159.090 ;
        RECT 101.685 158.360 101.975 159.525 ;
        RECT 102.145 158.435 103.355 159.525 ;
        RECT 103.525 158.435 107.035 159.525 ;
        RECT 107.410 158.555 107.740 159.355 ;
        RECT 107.910 158.725 108.240 159.525 ;
        RECT 108.540 158.555 108.870 159.355 ;
        RECT 109.515 158.725 109.765 159.525 ;
        RECT 94.325 156.975 95.995 157.745 ;
        RECT 99.590 157.520 99.930 158.350 ;
        RECT 102.145 157.895 102.665 158.435 ;
        RECT 102.835 157.725 103.355 158.265 ;
        RECT 103.525 157.915 105.215 158.435 ;
        RECT 107.410 158.385 109.845 158.555 ;
        RECT 110.035 158.385 110.205 159.525 ;
        RECT 110.375 158.385 110.715 159.355 ;
        RECT 105.385 157.745 107.035 158.265 ;
        RECT 107.205 157.965 107.555 158.215 ;
        RECT 107.740 157.755 107.910 158.385 ;
        RECT 108.080 157.965 108.410 158.165 ;
        RECT 108.580 157.965 108.910 158.165 ;
        RECT 109.080 157.965 109.500 158.165 ;
        RECT 109.675 158.135 109.845 158.385 ;
        RECT 109.675 157.965 110.370 158.135 ;
        RECT 96.170 156.975 101.515 157.520 ;
        RECT 101.685 156.975 101.975 157.700 ;
        RECT 102.145 156.975 103.355 157.725 ;
        RECT 103.525 156.975 107.035 157.745 ;
        RECT 107.410 157.145 107.910 157.755 ;
        RECT 108.540 157.625 109.765 157.795 ;
        RECT 110.540 157.775 110.715 158.385 ;
        RECT 108.540 157.145 108.870 157.625 ;
        RECT 109.040 156.975 109.265 157.435 ;
        RECT 109.435 157.145 109.765 157.625 ;
        RECT 109.955 156.975 110.205 157.775 ;
        RECT 110.375 157.145 110.715 157.775 ;
        RECT 110.885 158.385 111.225 159.355 ;
        RECT 111.395 158.385 111.565 159.525 ;
        RECT 111.835 158.725 112.085 159.525 ;
        RECT 112.730 158.555 113.060 159.355 ;
        RECT 113.360 158.725 113.690 159.525 ;
        RECT 113.860 158.555 114.190 159.355 ;
        RECT 115.490 159.090 120.835 159.525 ;
        RECT 121.010 159.090 126.355 159.525 ;
        RECT 111.755 158.385 114.190 158.555 ;
        RECT 110.885 157.775 111.060 158.385 ;
        RECT 111.755 158.135 111.925 158.385 ;
        RECT 111.230 157.965 111.925 158.135 ;
        RECT 112.100 157.965 112.520 158.165 ;
        RECT 112.690 157.965 113.020 158.165 ;
        RECT 113.190 157.965 113.520 158.165 ;
        RECT 110.885 157.145 111.225 157.775 ;
        RECT 111.395 156.975 111.645 157.775 ;
        RECT 111.835 157.625 113.060 157.795 ;
        RECT 111.835 157.145 112.165 157.625 ;
        RECT 112.335 156.975 112.560 157.435 ;
        RECT 112.730 157.145 113.060 157.625 ;
        RECT 113.690 157.755 113.860 158.385 ;
        RECT 114.045 157.965 114.395 158.215 ;
        RECT 117.080 157.840 117.430 159.090 ;
        RECT 113.690 157.145 114.190 157.755 ;
        RECT 118.910 157.520 119.250 158.350 ;
        RECT 122.600 157.840 122.950 159.090 ;
        RECT 126.525 158.435 127.735 159.525 ;
        RECT 124.430 157.520 124.770 158.350 ;
        RECT 126.525 157.895 127.045 158.435 ;
        RECT 127.215 157.725 127.735 158.265 ;
        RECT 115.490 156.975 120.835 157.520 ;
        RECT 121.010 156.975 126.355 157.520 ;
        RECT 126.525 156.975 127.735 157.725 ;
        RECT 20.640 156.805 127.820 156.975 ;
        RECT 20.725 156.055 21.935 156.805 ;
        RECT 23.400 156.465 23.655 156.625 ;
        RECT 23.315 156.295 23.655 156.465 ;
        RECT 23.835 156.345 24.120 156.805 ;
        RECT 23.400 156.095 23.655 156.295 ;
        RECT 20.725 155.515 21.245 156.055 ;
        RECT 21.415 155.345 21.935 155.885 ;
        RECT 20.725 154.255 21.935 155.345 ;
        RECT 23.400 155.235 23.580 156.095 ;
        RECT 24.300 155.895 24.550 156.545 ;
        RECT 23.750 155.565 24.550 155.895 ;
        RECT 23.400 154.565 23.655 155.235 ;
        RECT 23.835 154.255 24.120 155.055 ;
        RECT 24.300 154.975 24.550 155.565 ;
        RECT 24.750 156.210 25.070 156.540 ;
        RECT 25.250 156.325 25.910 156.805 ;
        RECT 26.110 156.415 26.960 156.585 ;
        RECT 24.750 155.315 24.940 156.210 ;
        RECT 25.260 155.885 25.920 156.155 ;
        RECT 25.590 155.825 25.920 155.885 ;
        RECT 25.110 155.655 25.440 155.715 ;
        RECT 26.110 155.655 26.280 156.415 ;
        RECT 27.520 156.345 27.840 156.805 ;
        RECT 28.040 156.165 28.290 156.595 ;
        RECT 28.580 156.365 28.990 156.805 ;
        RECT 29.160 156.425 30.175 156.625 ;
        RECT 26.450 155.995 27.700 156.165 ;
        RECT 26.450 155.875 26.780 155.995 ;
        RECT 25.110 155.485 27.010 155.655 ;
        RECT 24.750 155.145 26.670 155.315 ;
        RECT 24.750 155.125 25.070 155.145 ;
        RECT 24.300 154.465 24.630 154.975 ;
        RECT 24.900 154.515 25.070 155.125 ;
        RECT 26.840 154.975 27.010 155.485 ;
        RECT 27.180 155.415 27.360 155.825 ;
        RECT 27.530 155.235 27.700 155.995 ;
        RECT 25.240 154.255 25.570 154.945 ;
        RECT 25.800 154.805 27.010 154.975 ;
        RECT 27.180 154.925 27.700 155.235 ;
        RECT 27.870 155.825 28.290 156.165 ;
        RECT 28.580 155.825 28.990 156.155 ;
        RECT 27.870 155.055 28.060 155.825 ;
        RECT 29.160 155.695 29.330 156.425 ;
        RECT 30.475 156.255 30.645 156.585 ;
        RECT 30.815 156.425 31.145 156.805 ;
        RECT 29.500 155.875 29.850 156.245 ;
        RECT 29.160 155.655 29.580 155.695 ;
        RECT 28.230 155.485 29.580 155.655 ;
        RECT 28.230 155.325 28.480 155.485 ;
        RECT 28.990 155.055 29.240 155.315 ;
        RECT 27.870 154.805 29.240 155.055 ;
        RECT 25.800 154.515 26.040 154.805 ;
        RECT 26.840 154.725 27.010 154.805 ;
        RECT 26.240 154.255 26.660 154.635 ;
        RECT 26.840 154.475 27.470 154.725 ;
        RECT 27.940 154.255 28.270 154.635 ;
        RECT 28.440 154.515 28.610 154.805 ;
        RECT 29.410 154.640 29.580 155.485 ;
        RECT 30.030 155.315 30.250 156.185 ;
        RECT 30.475 156.065 31.170 156.255 ;
        RECT 29.750 154.935 30.250 155.315 ;
        RECT 30.420 155.265 30.830 155.885 ;
        RECT 31.000 155.095 31.170 156.065 ;
        RECT 30.475 154.925 31.170 155.095 ;
        RECT 28.790 154.255 29.170 154.635 ;
        RECT 29.410 154.470 30.240 154.640 ;
        RECT 30.475 154.425 30.645 154.925 ;
        RECT 30.815 154.255 31.145 154.755 ;
        RECT 31.360 154.425 31.585 156.545 ;
        RECT 31.755 156.425 32.085 156.805 ;
        RECT 32.255 156.255 32.425 156.545 ;
        RECT 31.760 156.085 32.425 156.255 ;
        RECT 32.685 156.130 32.945 156.635 ;
        RECT 33.125 156.425 33.455 156.805 ;
        RECT 33.635 156.255 33.805 156.635 ;
        RECT 31.760 155.095 31.990 156.085 ;
        RECT 32.160 155.265 32.510 155.915 ;
        RECT 32.685 155.330 32.855 156.130 ;
        RECT 33.140 156.085 33.805 156.255 ;
        RECT 33.140 155.830 33.310 156.085 ;
        RECT 34.525 156.035 37.115 156.805 ;
        RECT 37.285 156.080 37.575 156.805 ;
        RECT 33.025 155.500 33.310 155.830 ;
        RECT 33.545 155.535 33.875 155.905 ;
        RECT 33.140 155.355 33.310 155.500 ;
        RECT 31.760 154.925 32.425 155.095 ;
        RECT 31.755 154.255 32.085 154.755 ;
        RECT 32.255 154.425 32.425 154.925 ;
        RECT 32.685 154.425 32.955 155.330 ;
        RECT 33.140 155.185 33.805 155.355 ;
        RECT 33.125 154.255 33.455 155.015 ;
        RECT 33.635 154.425 33.805 155.185 ;
        RECT 34.525 155.345 35.735 155.865 ;
        RECT 35.905 155.515 37.115 156.035 ;
        RECT 38.020 155.995 38.265 156.600 ;
        RECT 38.485 156.270 38.995 156.805 ;
        RECT 37.745 155.825 38.975 155.995 ;
        RECT 34.525 154.255 37.115 155.345 ;
        RECT 37.285 154.255 37.575 155.420 ;
        RECT 37.745 155.015 38.085 155.825 ;
        RECT 38.255 155.260 39.005 155.450 ;
        RECT 37.745 154.605 38.260 155.015 ;
        RECT 38.495 154.255 38.665 155.015 ;
        RECT 38.835 154.595 39.005 155.260 ;
        RECT 39.175 155.275 39.365 156.635 ;
        RECT 39.535 156.125 39.810 156.635 ;
        RECT 40.000 156.270 40.530 156.635 ;
        RECT 40.955 156.405 41.285 156.805 ;
        RECT 40.355 156.235 40.530 156.270 ;
        RECT 39.535 155.955 39.815 156.125 ;
        RECT 39.535 155.475 39.810 155.955 ;
        RECT 40.015 155.275 40.185 156.075 ;
        RECT 39.175 155.105 40.185 155.275 ;
        RECT 40.355 156.065 41.285 156.235 ;
        RECT 41.455 156.065 41.710 156.635 ;
        RECT 40.355 154.935 40.525 156.065 ;
        RECT 41.115 155.895 41.285 156.065 ;
        RECT 39.400 154.765 40.525 154.935 ;
        RECT 40.695 155.565 40.890 155.895 ;
        RECT 41.115 155.565 41.370 155.895 ;
        RECT 40.695 154.595 40.865 155.565 ;
        RECT 41.540 155.395 41.710 156.065 ;
        RECT 38.835 154.425 40.865 154.595 ;
        RECT 41.035 154.255 41.205 155.395 ;
        RECT 41.375 154.425 41.710 155.395 ;
        RECT 41.885 156.130 42.145 156.635 ;
        RECT 42.325 156.425 42.655 156.805 ;
        RECT 42.835 156.255 43.005 156.635 ;
        RECT 41.885 155.330 42.055 156.130 ;
        RECT 42.340 156.085 43.005 156.255 ;
        RECT 42.340 155.830 42.510 156.085 ;
        RECT 43.265 156.035 44.935 156.805 ;
        RECT 42.225 155.500 42.510 155.830 ;
        RECT 42.745 155.535 43.075 155.905 ;
        RECT 42.340 155.355 42.510 155.500 ;
        RECT 41.885 154.425 42.155 155.330 ;
        RECT 42.340 155.185 43.005 155.355 ;
        RECT 42.325 154.255 42.655 155.015 ;
        RECT 42.835 154.425 43.005 155.185 ;
        RECT 43.265 155.345 44.015 155.865 ;
        RECT 44.185 155.515 44.935 156.035 ;
        RECT 45.310 156.025 45.810 156.635 ;
        RECT 45.105 155.565 45.455 155.815 ;
        RECT 45.640 155.395 45.810 156.025 ;
        RECT 46.440 156.155 46.770 156.635 ;
        RECT 46.940 156.345 47.165 156.805 ;
        RECT 47.335 156.155 47.665 156.635 ;
        RECT 46.440 155.985 47.665 156.155 ;
        RECT 47.855 156.005 48.105 156.805 ;
        RECT 48.275 156.005 48.615 156.635 ;
        RECT 49.705 156.035 53.215 156.805 ;
        RECT 45.980 155.615 46.310 155.815 ;
        RECT 46.480 155.615 46.810 155.815 ;
        RECT 46.980 155.615 47.400 155.815 ;
        RECT 47.575 155.645 48.270 155.815 ;
        RECT 47.575 155.395 47.745 155.645 ;
        RECT 48.440 155.395 48.615 156.005 ;
        RECT 43.265 154.255 44.935 155.345 ;
        RECT 45.310 155.225 47.745 155.395 ;
        RECT 45.310 154.425 45.640 155.225 ;
        RECT 45.810 154.255 46.140 155.055 ;
        RECT 46.440 154.425 46.770 155.225 ;
        RECT 47.415 154.255 47.665 155.055 ;
        RECT 47.935 154.255 48.105 155.395 ;
        RECT 48.275 154.425 48.615 155.395 ;
        RECT 49.705 155.345 51.395 155.865 ;
        RECT 51.565 155.515 53.215 156.035 ;
        RECT 53.760 156.095 54.015 156.625 ;
        RECT 54.195 156.345 54.480 156.805 ;
        RECT 49.705 154.255 53.215 155.345 ;
        RECT 53.760 155.235 53.940 156.095 ;
        RECT 54.660 155.895 54.910 156.545 ;
        RECT 54.110 155.565 54.910 155.895 ;
        RECT 53.760 154.765 54.015 155.235 ;
        RECT 53.675 154.595 54.015 154.765 ;
        RECT 53.760 154.565 54.015 154.595 ;
        RECT 54.195 154.255 54.480 155.055 ;
        RECT 54.660 154.975 54.910 155.565 ;
        RECT 55.110 156.210 55.430 156.540 ;
        RECT 55.610 156.325 56.270 156.805 ;
        RECT 56.470 156.415 57.320 156.585 ;
        RECT 55.110 155.315 55.300 156.210 ;
        RECT 55.620 155.885 56.280 156.155 ;
        RECT 55.950 155.825 56.280 155.885 ;
        RECT 55.470 155.655 55.800 155.715 ;
        RECT 56.470 155.655 56.640 156.415 ;
        RECT 57.880 156.345 58.200 156.805 ;
        RECT 58.400 156.165 58.650 156.595 ;
        RECT 58.940 156.365 59.350 156.805 ;
        RECT 59.520 156.425 60.535 156.625 ;
        RECT 56.810 155.995 58.060 156.165 ;
        RECT 56.810 155.875 57.140 155.995 ;
        RECT 55.470 155.485 57.370 155.655 ;
        RECT 55.110 155.145 57.030 155.315 ;
        RECT 55.110 155.125 55.430 155.145 ;
        RECT 54.660 154.465 54.990 154.975 ;
        RECT 55.260 154.515 55.430 155.125 ;
        RECT 57.200 154.975 57.370 155.485 ;
        RECT 57.540 155.415 57.720 155.825 ;
        RECT 57.890 155.235 58.060 155.995 ;
        RECT 55.600 154.255 55.930 154.945 ;
        RECT 56.160 154.805 57.370 154.975 ;
        RECT 57.540 154.925 58.060 155.235 ;
        RECT 58.230 155.825 58.650 156.165 ;
        RECT 58.940 155.825 59.350 156.155 ;
        RECT 58.230 155.055 58.420 155.825 ;
        RECT 59.520 155.695 59.690 156.425 ;
        RECT 60.835 156.255 61.005 156.585 ;
        RECT 61.175 156.425 61.505 156.805 ;
        RECT 59.860 155.875 60.210 156.245 ;
        RECT 59.520 155.655 59.940 155.695 ;
        RECT 58.590 155.485 59.940 155.655 ;
        RECT 58.590 155.325 58.840 155.485 ;
        RECT 59.350 155.055 59.600 155.315 ;
        RECT 58.230 154.805 59.600 155.055 ;
        RECT 56.160 154.515 56.400 154.805 ;
        RECT 57.200 154.725 57.370 154.805 ;
        RECT 56.600 154.255 57.020 154.635 ;
        RECT 57.200 154.475 57.830 154.725 ;
        RECT 58.300 154.255 58.630 154.635 ;
        RECT 58.800 154.515 58.970 154.805 ;
        RECT 59.770 154.640 59.940 155.485 ;
        RECT 60.390 155.315 60.610 156.185 ;
        RECT 60.835 156.065 61.530 156.255 ;
        RECT 60.110 154.935 60.610 155.315 ;
        RECT 60.780 155.265 61.190 155.885 ;
        RECT 61.360 155.095 61.530 156.065 ;
        RECT 60.835 154.925 61.530 155.095 ;
        RECT 59.150 154.255 59.530 154.635 ;
        RECT 59.770 154.470 60.600 154.640 ;
        RECT 60.835 154.425 61.005 154.925 ;
        RECT 61.175 154.255 61.505 154.755 ;
        RECT 61.720 154.425 61.945 156.545 ;
        RECT 62.115 156.425 62.445 156.805 ;
        RECT 62.615 156.255 62.785 156.545 ;
        RECT 62.120 156.085 62.785 156.255 ;
        RECT 62.120 155.095 62.350 156.085 ;
        RECT 63.045 156.080 63.335 156.805 ;
        RECT 63.505 156.130 63.765 156.635 ;
        RECT 63.945 156.425 64.275 156.805 ;
        RECT 64.455 156.255 64.625 156.635 ;
        RECT 62.520 155.265 62.870 155.915 ;
        RECT 62.120 154.925 62.785 155.095 ;
        RECT 62.115 154.255 62.445 154.755 ;
        RECT 62.615 154.425 62.785 154.925 ;
        RECT 63.045 154.255 63.335 155.420 ;
        RECT 63.505 155.330 63.675 156.130 ;
        RECT 63.960 156.085 64.625 156.255 ;
        RECT 63.960 155.830 64.130 156.085 ;
        RECT 64.885 156.035 66.555 156.805 ;
        RECT 66.815 156.255 66.985 156.635 ;
        RECT 67.165 156.425 67.495 156.805 ;
        RECT 66.815 156.085 67.480 156.255 ;
        RECT 67.675 156.130 67.935 156.635 ;
        RECT 63.845 155.500 64.130 155.830 ;
        RECT 64.365 155.535 64.695 155.905 ;
        RECT 63.960 155.355 64.130 155.500 ;
        RECT 63.505 154.425 63.775 155.330 ;
        RECT 63.960 155.185 64.625 155.355 ;
        RECT 63.945 154.255 64.275 155.015 ;
        RECT 64.455 154.425 64.625 155.185 ;
        RECT 64.885 155.345 65.635 155.865 ;
        RECT 65.805 155.515 66.555 156.035 ;
        RECT 66.745 155.535 67.075 155.905 ;
        RECT 67.310 155.830 67.480 156.085 ;
        RECT 67.310 155.500 67.595 155.830 ;
        RECT 67.310 155.355 67.480 155.500 ;
        RECT 64.885 154.255 66.555 155.345 ;
        RECT 66.815 155.185 67.480 155.355 ;
        RECT 67.765 155.330 67.935 156.130 ;
        RECT 68.110 155.965 68.370 156.805 ;
        RECT 68.545 156.060 68.800 156.635 ;
        RECT 68.970 156.425 69.300 156.805 ;
        RECT 69.515 156.255 69.685 156.635 ;
        RECT 68.970 156.085 69.685 156.255 ;
        RECT 66.815 154.425 66.985 155.185 ;
        RECT 67.165 154.255 67.495 155.015 ;
        RECT 67.665 154.425 67.935 155.330 ;
        RECT 68.110 154.255 68.370 155.405 ;
        RECT 68.545 155.330 68.715 156.060 ;
        RECT 68.970 155.895 69.140 156.085 ;
        RECT 69.950 155.965 70.210 156.805 ;
        RECT 70.385 156.060 70.640 156.635 ;
        RECT 70.810 156.425 71.140 156.805 ;
        RECT 71.355 156.255 71.525 156.635 ;
        RECT 72.765 156.325 73.045 156.805 ;
        RECT 70.810 156.085 71.525 156.255 ;
        RECT 73.215 156.155 73.475 156.545 ;
        RECT 73.650 156.325 73.905 156.805 ;
        RECT 74.075 156.155 74.370 156.545 ;
        RECT 74.550 156.325 74.825 156.805 ;
        RECT 74.995 156.305 75.295 156.635 ;
        RECT 68.885 155.565 69.140 155.895 ;
        RECT 68.970 155.355 69.140 155.565 ;
        RECT 69.420 155.535 69.775 155.905 ;
        RECT 68.545 154.425 68.800 155.330 ;
        RECT 68.970 155.185 69.685 155.355 ;
        RECT 68.970 154.255 69.300 155.015 ;
        RECT 69.515 154.425 69.685 155.185 ;
        RECT 69.950 154.255 70.210 155.405 ;
        RECT 70.385 155.330 70.555 156.060 ;
        RECT 70.810 155.895 70.980 156.085 ;
        RECT 72.720 155.985 74.370 156.155 ;
        RECT 70.725 155.565 70.980 155.895 ;
        RECT 70.810 155.355 70.980 155.565 ;
        RECT 71.260 155.535 71.615 155.905 ;
        RECT 72.720 155.475 73.125 155.985 ;
        RECT 73.295 155.645 74.435 155.815 ;
        RECT 70.385 154.425 70.640 155.330 ;
        RECT 70.810 155.185 71.525 155.355 ;
        RECT 72.720 155.305 73.475 155.475 ;
        RECT 70.810 154.255 71.140 155.015 ;
        RECT 71.355 154.425 71.525 155.185 ;
        RECT 72.760 154.255 73.045 155.125 ;
        RECT 73.215 155.055 73.475 155.305 ;
        RECT 74.265 155.395 74.435 155.645 ;
        RECT 74.605 155.565 74.955 156.135 ;
        RECT 75.125 155.395 75.295 156.305 ;
        RECT 75.555 156.255 75.725 156.635 ;
        RECT 75.940 156.425 76.270 156.805 ;
        RECT 75.555 156.085 76.270 156.255 ;
        RECT 75.465 155.535 75.820 155.905 ;
        RECT 76.100 155.895 76.270 156.085 ;
        RECT 76.440 156.060 76.695 156.635 ;
        RECT 76.100 155.565 76.355 155.895 ;
        RECT 74.265 155.225 75.295 155.395 ;
        RECT 76.100 155.355 76.270 155.565 ;
        RECT 73.215 154.885 74.335 155.055 ;
        RECT 73.215 154.425 73.475 154.885 ;
        RECT 73.650 154.255 73.905 154.715 ;
        RECT 74.075 154.425 74.335 154.885 ;
        RECT 74.505 154.255 74.815 155.055 ;
        RECT 74.985 154.425 75.295 155.225 ;
        RECT 75.555 155.185 76.270 155.355 ;
        RECT 76.525 155.330 76.695 156.060 ;
        RECT 76.870 155.965 77.130 156.805 ;
        RECT 77.305 156.055 78.515 156.805 ;
        RECT 75.555 154.425 75.725 155.185 ;
        RECT 75.940 154.255 76.270 155.015 ;
        RECT 76.440 154.425 76.695 155.330 ;
        RECT 76.870 154.255 77.130 155.405 ;
        RECT 77.305 155.345 77.825 155.885 ;
        RECT 77.995 155.515 78.515 156.055 ;
        RECT 78.685 156.305 78.985 156.635 ;
        RECT 79.155 156.325 79.430 156.805 ;
        RECT 78.685 155.395 78.855 156.305 ;
        RECT 79.610 156.155 79.905 156.545 ;
        RECT 80.075 156.325 80.330 156.805 ;
        RECT 80.505 156.155 80.765 156.545 ;
        RECT 80.935 156.325 81.215 156.805 ;
        RECT 79.025 155.565 79.375 156.135 ;
        RECT 79.610 155.985 81.260 156.155 ;
        RECT 79.545 155.645 80.685 155.815 ;
        RECT 79.545 155.395 79.715 155.645 ;
        RECT 80.855 155.475 81.260 155.985 ;
        RECT 77.305 154.255 78.515 155.345 ;
        RECT 78.685 155.225 79.715 155.395 ;
        RECT 80.505 155.305 81.260 155.475 ;
        RECT 81.445 156.005 81.785 156.635 ;
        RECT 81.955 156.005 82.205 156.805 ;
        RECT 82.395 156.155 82.725 156.635 ;
        RECT 82.895 156.345 83.120 156.805 ;
        RECT 83.290 156.155 83.620 156.635 ;
        RECT 81.445 155.955 81.675 156.005 ;
        RECT 82.395 155.985 83.620 156.155 ;
        RECT 84.250 156.025 84.750 156.635 ;
        RECT 85.125 156.035 88.635 156.805 ;
        RECT 88.805 156.080 89.095 156.805 ;
        RECT 89.640 156.095 89.895 156.625 ;
        RECT 90.075 156.345 90.360 156.805 ;
        RECT 81.445 155.395 81.620 155.955 ;
        RECT 81.790 155.645 82.485 155.815 ;
        RECT 82.315 155.395 82.485 155.645 ;
        RECT 82.660 155.615 83.080 155.815 ;
        RECT 83.250 155.615 83.580 155.815 ;
        RECT 83.750 155.615 84.080 155.815 ;
        RECT 84.250 155.395 84.420 156.025 ;
        RECT 84.605 155.565 84.955 155.815 ;
        RECT 78.685 154.425 78.995 155.225 ;
        RECT 80.505 155.055 80.765 155.305 ;
        RECT 79.165 154.255 79.475 155.055 ;
        RECT 79.645 154.885 80.765 155.055 ;
        RECT 79.645 154.425 79.905 154.885 ;
        RECT 80.075 154.255 80.330 154.715 ;
        RECT 80.505 154.425 80.765 154.885 ;
        RECT 80.935 154.255 81.220 155.125 ;
        RECT 81.445 154.425 81.785 155.395 ;
        RECT 81.955 154.255 82.125 155.395 ;
        RECT 82.315 155.225 84.750 155.395 ;
        RECT 82.395 154.255 82.645 155.055 ;
        RECT 83.290 154.425 83.620 155.225 ;
        RECT 83.920 154.255 84.250 155.055 ;
        RECT 84.420 154.425 84.750 155.225 ;
        RECT 85.125 155.345 86.815 155.865 ;
        RECT 86.985 155.515 88.635 156.035 ;
        RECT 85.125 154.255 88.635 155.345 ;
        RECT 88.805 154.255 89.095 155.420 ;
        RECT 89.640 155.235 89.820 156.095 ;
        RECT 90.540 155.895 90.790 156.545 ;
        RECT 89.990 155.565 90.790 155.895 ;
        RECT 89.640 154.765 89.895 155.235 ;
        RECT 89.555 154.595 89.895 154.765 ;
        RECT 89.640 154.565 89.895 154.595 ;
        RECT 90.075 154.255 90.360 155.055 ;
        RECT 90.540 154.975 90.790 155.565 ;
        RECT 90.990 156.210 91.310 156.540 ;
        RECT 91.490 156.325 92.150 156.805 ;
        RECT 92.350 156.415 93.200 156.585 ;
        RECT 90.990 155.315 91.180 156.210 ;
        RECT 91.500 155.885 92.160 156.155 ;
        RECT 91.830 155.825 92.160 155.885 ;
        RECT 91.350 155.655 91.680 155.715 ;
        RECT 92.350 155.655 92.520 156.415 ;
        RECT 93.760 156.345 94.080 156.805 ;
        RECT 94.280 156.165 94.530 156.595 ;
        RECT 94.820 156.365 95.230 156.805 ;
        RECT 95.400 156.425 96.415 156.625 ;
        RECT 92.690 155.995 93.940 156.165 ;
        RECT 92.690 155.875 93.020 155.995 ;
        RECT 91.350 155.485 93.250 155.655 ;
        RECT 90.990 155.145 92.910 155.315 ;
        RECT 90.990 155.125 91.310 155.145 ;
        RECT 90.540 154.465 90.870 154.975 ;
        RECT 91.140 154.515 91.310 155.125 ;
        RECT 93.080 154.975 93.250 155.485 ;
        RECT 93.420 155.415 93.600 155.825 ;
        RECT 93.770 155.235 93.940 155.995 ;
        RECT 91.480 154.255 91.810 154.945 ;
        RECT 92.040 154.805 93.250 154.975 ;
        RECT 93.420 154.925 93.940 155.235 ;
        RECT 94.110 155.825 94.530 156.165 ;
        RECT 94.820 155.825 95.230 156.155 ;
        RECT 94.110 155.055 94.300 155.825 ;
        RECT 95.400 155.695 95.570 156.425 ;
        RECT 96.715 156.255 96.885 156.585 ;
        RECT 97.055 156.425 97.385 156.805 ;
        RECT 95.740 155.875 96.090 156.245 ;
        RECT 95.400 155.655 95.820 155.695 ;
        RECT 94.470 155.485 95.820 155.655 ;
        RECT 94.470 155.325 94.720 155.485 ;
        RECT 95.230 155.055 95.480 155.315 ;
        RECT 94.110 154.805 95.480 155.055 ;
        RECT 92.040 154.515 92.280 154.805 ;
        RECT 93.080 154.725 93.250 154.805 ;
        RECT 92.480 154.255 92.900 154.635 ;
        RECT 93.080 154.475 93.710 154.725 ;
        RECT 94.180 154.255 94.510 154.635 ;
        RECT 94.680 154.515 94.850 154.805 ;
        RECT 95.650 154.640 95.820 155.485 ;
        RECT 96.270 155.315 96.490 156.185 ;
        RECT 96.715 156.065 97.410 156.255 ;
        RECT 95.990 154.935 96.490 155.315 ;
        RECT 96.660 155.265 97.070 155.885 ;
        RECT 97.240 155.095 97.410 156.065 ;
        RECT 96.715 154.925 97.410 155.095 ;
        RECT 95.030 154.255 95.410 154.635 ;
        RECT 95.650 154.470 96.480 154.640 ;
        RECT 96.715 154.425 96.885 154.925 ;
        RECT 97.055 154.255 97.385 154.755 ;
        RECT 97.600 154.425 97.825 156.545 ;
        RECT 97.995 156.425 98.325 156.805 ;
        RECT 98.495 156.255 98.665 156.545 ;
        RECT 98.000 156.085 98.665 156.255 ;
        RECT 98.000 155.095 98.230 156.085 ;
        RECT 99.385 156.005 99.725 156.635 ;
        RECT 99.895 156.005 100.145 156.805 ;
        RECT 100.335 156.155 100.665 156.635 ;
        RECT 100.835 156.345 101.060 156.805 ;
        RECT 101.230 156.155 101.560 156.635 ;
        RECT 98.400 155.265 98.750 155.915 ;
        RECT 99.385 155.395 99.560 156.005 ;
        RECT 100.335 155.985 101.560 156.155 ;
        RECT 102.190 156.025 102.690 156.635 ;
        RECT 103.525 156.035 106.115 156.805 ;
        RECT 99.730 155.645 100.425 155.815 ;
        RECT 100.255 155.395 100.425 155.645 ;
        RECT 100.600 155.615 101.020 155.815 ;
        RECT 101.190 155.615 101.520 155.815 ;
        RECT 101.690 155.615 102.020 155.815 ;
        RECT 102.190 155.395 102.360 156.025 ;
        RECT 102.545 155.565 102.895 155.815 ;
        RECT 98.000 154.925 98.665 155.095 ;
        RECT 97.995 154.255 98.325 154.755 ;
        RECT 98.495 154.425 98.665 154.925 ;
        RECT 99.385 154.425 99.725 155.395 ;
        RECT 99.895 154.255 100.065 155.395 ;
        RECT 100.255 155.225 102.690 155.395 ;
        RECT 100.335 154.255 100.585 155.055 ;
        RECT 101.230 154.425 101.560 155.225 ;
        RECT 101.860 154.255 102.190 155.055 ;
        RECT 102.360 154.425 102.690 155.225 ;
        RECT 103.525 155.345 104.735 155.865 ;
        RECT 104.905 155.515 106.115 156.035 ;
        RECT 106.285 156.005 106.625 156.635 ;
        RECT 106.795 156.005 107.045 156.805 ;
        RECT 107.235 156.155 107.565 156.635 ;
        RECT 107.735 156.345 107.960 156.805 ;
        RECT 108.130 156.155 108.460 156.635 ;
        RECT 106.285 155.395 106.460 156.005 ;
        RECT 107.235 155.985 108.460 156.155 ;
        RECT 109.090 156.025 109.590 156.635 ;
        RECT 106.630 155.645 107.325 155.815 ;
        RECT 107.155 155.395 107.325 155.645 ;
        RECT 107.500 155.615 107.920 155.815 ;
        RECT 108.090 155.615 108.420 155.815 ;
        RECT 108.590 155.615 108.920 155.815 ;
        RECT 109.090 155.395 109.260 156.025 ;
        RECT 109.965 156.005 110.305 156.635 ;
        RECT 110.475 156.005 110.725 156.805 ;
        RECT 110.915 156.155 111.245 156.635 ;
        RECT 111.415 156.345 111.640 156.805 ;
        RECT 111.810 156.155 112.140 156.635 ;
        RECT 109.445 155.565 109.795 155.815 ;
        RECT 109.965 155.395 110.140 156.005 ;
        RECT 110.915 155.985 112.140 156.155 ;
        RECT 112.770 156.025 113.270 156.635 ;
        RECT 114.565 156.080 114.855 156.805 ;
        RECT 110.310 155.645 111.005 155.815 ;
        RECT 110.835 155.395 111.005 155.645 ;
        RECT 111.180 155.615 111.600 155.815 ;
        RECT 111.770 155.615 112.100 155.815 ;
        RECT 112.270 155.615 112.600 155.815 ;
        RECT 112.770 155.395 112.940 156.025 ;
        RECT 115.985 155.985 116.215 156.805 ;
        RECT 116.385 156.005 116.715 156.635 ;
        RECT 113.125 155.565 113.475 155.815 ;
        RECT 115.965 155.565 116.295 155.815 ;
        RECT 103.525 154.255 106.115 155.345 ;
        RECT 106.285 154.425 106.625 155.395 ;
        RECT 106.795 154.255 106.965 155.395 ;
        RECT 107.155 155.225 109.590 155.395 ;
        RECT 107.235 154.255 107.485 155.055 ;
        RECT 108.130 154.425 108.460 155.225 ;
        RECT 108.760 154.255 109.090 155.055 ;
        RECT 109.260 154.425 109.590 155.225 ;
        RECT 109.965 154.425 110.305 155.395 ;
        RECT 110.475 154.255 110.645 155.395 ;
        RECT 110.835 155.225 113.270 155.395 ;
        RECT 110.915 154.255 111.165 155.055 ;
        RECT 111.810 154.425 112.140 155.225 ;
        RECT 112.440 154.255 112.770 155.055 ;
        RECT 112.940 154.425 113.270 155.225 ;
        RECT 114.565 154.255 114.855 155.420 ;
        RECT 116.465 155.405 116.715 156.005 ;
        RECT 116.885 155.985 117.095 156.805 ;
        RECT 117.330 156.095 117.585 156.625 ;
        RECT 117.755 156.345 118.060 156.805 ;
        RECT 118.305 156.425 119.375 156.595 ;
        RECT 115.985 154.255 116.215 155.395 ;
        RECT 116.385 154.425 116.715 155.405 ;
        RECT 117.330 155.445 117.540 156.095 ;
        RECT 118.305 156.070 118.625 156.425 ;
        RECT 118.300 155.895 118.625 156.070 ;
        RECT 117.710 155.595 118.625 155.895 ;
        RECT 118.795 155.855 119.035 156.255 ;
        RECT 119.205 156.195 119.375 156.425 ;
        RECT 119.545 156.365 119.735 156.805 ;
        RECT 119.905 156.355 120.855 156.635 ;
        RECT 121.075 156.445 121.425 156.615 ;
        RECT 119.205 156.025 119.735 156.195 ;
        RECT 117.710 155.565 118.450 155.595 ;
        RECT 116.885 154.255 117.095 155.395 ;
        RECT 117.330 154.565 117.585 155.445 ;
        RECT 117.755 154.255 118.060 155.395 ;
        RECT 118.280 154.975 118.450 155.565 ;
        RECT 118.795 155.485 119.335 155.855 ;
        RECT 119.515 155.745 119.735 156.025 ;
        RECT 119.905 155.575 120.075 156.355 ;
        RECT 119.670 155.405 120.075 155.575 ;
        RECT 120.245 155.565 120.595 156.185 ;
        RECT 119.670 155.315 119.840 155.405 ;
        RECT 120.765 155.395 120.975 156.185 ;
        RECT 118.620 155.145 119.840 155.315 ;
        RECT 120.300 155.235 120.975 155.395 ;
        RECT 118.280 154.805 119.080 154.975 ;
        RECT 118.400 154.255 118.730 154.635 ;
        RECT 118.910 154.515 119.080 154.805 ;
        RECT 119.670 154.765 119.840 155.145 ;
        RECT 120.010 155.225 120.975 155.235 ;
        RECT 121.165 156.055 121.425 156.445 ;
        RECT 121.635 156.345 121.965 156.805 ;
        RECT 122.840 156.415 123.695 156.585 ;
        RECT 123.900 156.415 124.395 156.585 ;
        RECT 124.565 156.445 124.895 156.805 ;
        RECT 121.165 155.365 121.335 156.055 ;
        RECT 121.505 155.705 121.675 155.885 ;
        RECT 121.845 155.875 122.635 156.125 ;
        RECT 122.840 155.705 123.010 156.415 ;
        RECT 123.180 155.905 123.535 156.125 ;
        RECT 121.505 155.535 123.195 155.705 ;
        RECT 120.010 154.935 120.470 155.225 ;
        RECT 121.165 155.195 122.665 155.365 ;
        RECT 121.165 155.055 121.335 155.195 ;
        RECT 120.775 154.885 121.335 155.055 ;
        RECT 119.250 154.255 119.500 154.715 ;
        RECT 119.670 154.425 120.540 154.765 ;
        RECT 120.775 154.425 120.945 154.885 ;
        RECT 121.780 154.855 122.855 155.025 ;
        RECT 121.115 154.255 121.485 154.715 ;
        RECT 121.780 154.515 121.950 154.855 ;
        RECT 122.120 154.255 122.450 154.685 ;
        RECT 122.685 154.515 122.855 154.855 ;
        RECT 123.025 154.755 123.195 155.535 ;
        RECT 123.365 155.315 123.535 155.905 ;
        RECT 123.705 155.505 124.055 156.125 ;
        RECT 123.365 154.925 123.830 155.315 ;
        RECT 124.225 155.055 124.395 156.415 ;
        RECT 124.565 155.225 125.025 156.275 ;
        RECT 124.000 154.885 124.395 155.055 ;
        RECT 124.000 154.755 124.170 154.885 ;
        RECT 123.025 154.425 123.705 154.755 ;
        RECT 123.920 154.425 124.170 154.755 ;
        RECT 124.340 154.255 124.590 154.715 ;
        RECT 124.760 154.440 125.085 155.225 ;
        RECT 125.255 154.425 125.425 156.545 ;
        RECT 125.595 156.425 125.925 156.805 ;
        RECT 126.095 156.255 126.350 156.545 ;
        RECT 125.600 156.085 126.350 156.255 ;
        RECT 125.600 155.095 125.830 156.085 ;
        RECT 126.525 156.055 127.735 156.805 ;
        RECT 126.000 155.265 126.350 155.915 ;
        RECT 126.525 155.345 127.045 155.885 ;
        RECT 127.215 155.515 127.735 156.055 ;
        RECT 125.600 154.925 126.350 155.095 ;
        RECT 125.595 154.255 125.925 154.755 ;
        RECT 126.095 154.425 126.350 154.925 ;
        RECT 126.525 154.255 127.735 155.345 ;
        RECT 20.640 154.085 127.820 154.255 ;
        RECT 20.725 152.995 21.935 154.085 ;
        RECT 20.725 152.285 21.245 152.825 ;
        RECT 21.415 152.455 21.935 152.995 ;
        RECT 22.565 152.995 24.235 154.085 ;
        RECT 22.565 152.475 23.315 152.995 ;
        RECT 24.405 152.920 24.695 154.085 ;
        RECT 25.875 153.155 26.045 153.915 ;
        RECT 26.225 153.325 26.555 154.085 ;
        RECT 25.875 152.985 26.540 153.155 ;
        RECT 26.725 153.010 26.995 153.915 ;
        RECT 26.370 152.840 26.540 152.985 ;
        RECT 23.485 152.305 24.235 152.825 ;
        RECT 25.805 152.435 26.135 152.805 ;
        RECT 26.370 152.510 26.655 152.840 ;
        RECT 20.725 151.535 21.935 152.285 ;
        RECT 22.565 151.535 24.235 152.305 ;
        RECT 24.405 151.535 24.695 152.260 ;
        RECT 26.370 152.255 26.540 152.510 ;
        RECT 25.875 152.085 26.540 152.255 ;
        RECT 26.825 152.210 26.995 153.010 ;
        RECT 25.875 151.705 26.045 152.085 ;
        RECT 26.225 151.535 26.555 151.915 ;
        RECT 26.735 151.705 26.995 152.210 ;
        RECT 27.170 152.945 27.505 153.915 ;
        RECT 27.675 152.945 27.845 154.085 ;
        RECT 28.015 153.745 30.045 153.915 ;
        RECT 27.170 152.275 27.340 152.945 ;
        RECT 28.015 152.775 28.185 153.745 ;
        RECT 27.510 152.445 27.765 152.775 ;
        RECT 27.990 152.445 28.185 152.775 ;
        RECT 28.355 153.405 29.480 153.575 ;
        RECT 27.595 152.275 27.765 152.445 ;
        RECT 28.355 152.275 28.525 153.405 ;
        RECT 27.170 151.705 27.425 152.275 ;
        RECT 27.595 152.105 28.525 152.275 ;
        RECT 28.695 153.065 29.705 153.235 ;
        RECT 28.695 152.265 28.865 153.065 ;
        RECT 28.350 152.070 28.525 152.105 ;
        RECT 27.595 151.535 27.925 151.935 ;
        RECT 28.350 151.705 28.880 152.070 ;
        RECT 29.070 152.045 29.345 152.865 ;
        RECT 29.065 151.875 29.345 152.045 ;
        RECT 29.070 151.705 29.345 151.875 ;
        RECT 29.515 151.705 29.705 153.065 ;
        RECT 29.875 153.080 30.045 153.745 ;
        RECT 30.215 153.325 30.385 154.085 ;
        RECT 30.620 153.325 31.135 153.735 ;
        RECT 31.770 153.650 37.115 154.085 ;
        RECT 37.290 153.650 42.635 154.085 ;
        RECT 29.875 152.890 30.625 153.080 ;
        RECT 30.795 152.515 31.135 153.325 ;
        RECT 29.905 152.345 31.135 152.515 ;
        RECT 33.360 152.400 33.710 153.650 ;
        RECT 29.885 151.535 30.395 152.070 ;
        RECT 30.615 151.740 30.860 152.345 ;
        RECT 35.190 152.080 35.530 152.910 ;
        RECT 38.880 152.400 39.230 153.650 ;
        RECT 42.805 152.945 43.145 153.915 ;
        RECT 43.315 152.945 43.485 154.085 ;
        RECT 43.755 153.285 44.005 154.085 ;
        RECT 44.650 153.115 44.980 153.915 ;
        RECT 45.280 153.285 45.610 154.085 ;
        RECT 45.780 153.115 46.110 153.915 ;
        RECT 43.675 152.945 46.110 153.115 ;
        RECT 47.405 152.945 47.675 153.915 ;
        RECT 47.885 153.285 48.165 154.085 ;
        RECT 48.335 153.575 49.990 153.865 ;
        RECT 48.400 153.235 49.990 153.405 ;
        RECT 48.400 153.115 48.570 153.235 ;
        RECT 47.845 152.945 48.570 153.115 ;
        RECT 40.710 152.080 41.050 152.910 ;
        RECT 42.805 152.335 42.980 152.945 ;
        RECT 43.675 152.695 43.845 152.945 ;
        RECT 43.150 152.525 43.845 152.695 ;
        RECT 44.020 152.525 44.440 152.725 ;
        RECT 44.610 152.525 44.940 152.725 ;
        RECT 45.110 152.525 45.440 152.725 ;
        RECT 31.770 151.535 37.115 152.080 ;
        RECT 37.290 151.535 42.635 152.080 ;
        RECT 42.805 151.705 43.145 152.335 ;
        RECT 43.315 151.535 43.565 152.335 ;
        RECT 43.755 152.185 44.980 152.355 ;
        RECT 43.755 151.705 44.085 152.185 ;
        RECT 44.255 151.535 44.480 151.995 ;
        RECT 44.650 151.705 44.980 152.185 ;
        RECT 45.610 152.315 45.780 152.945 ;
        RECT 45.965 152.525 46.315 152.775 ;
        RECT 45.610 151.705 46.110 152.315 ;
        RECT 47.405 152.210 47.575 152.945 ;
        RECT 47.845 152.775 48.015 152.945 ;
        RECT 48.760 152.895 49.475 153.065 ;
        RECT 49.670 152.945 49.990 153.235 ;
        RECT 50.165 152.920 50.455 154.085 ;
        RECT 50.625 152.945 50.895 153.915 ;
        RECT 51.105 153.285 51.385 154.085 ;
        RECT 51.555 153.575 53.210 153.865 ;
        RECT 51.620 153.235 53.210 153.405 ;
        RECT 51.620 153.115 51.790 153.235 ;
        RECT 51.065 152.945 51.790 153.115 ;
        RECT 47.745 152.445 48.015 152.775 ;
        RECT 48.185 152.445 48.590 152.775 ;
        RECT 48.760 152.445 49.470 152.895 ;
        RECT 47.845 152.275 48.015 152.445 ;
        RECT 47.405 151.865 47.675 152.210 ;
        RECT 47.845 152.105 49.455 152.275 ;
        RECT 49.640 152.205 49.990 152.775 ;
        RECT 47.865 151.535 48.245 151.935 ;
        RECT 48.415 151.755 48.585 152.105 ;
        RECT 48.755 151.535 49.085 151.935 ;
        RECT 49.285 151.755 49.455 152.105 ;
        RECT 49.655 151.535 49.985 152.035 ;
        RECT 50.165 151.535 50.455 152.260 ;
        RECT 50.625 152.210 50.795 152.945 ;
        RECT 51.065 152.775 51.235 152.945 ;
        RECT 50.965 152.445 51.235 152.775 ;
        RECT 51.405 152.445 51.810 152.775 ;
        RECT 51.980 152.445 52.690 153.065 ;
        RECT 52.890 152.945 53.210 153.235 ;
        RECT 53.385 152.945 53.725 153.915 ;
        RECT 53.895 152.945 54.065 154.085 ;
        RECT 54.335 153.285 54.585 154.085 ;
        RECT 55.230 153.115 55.560 153.915 ;
        RECT 55.860 153.285 56.190 154.085 ;
        RECT 56.360 153.115 56.690 153.915 ;
        RECT 54.255 152.945 56.690 153.115 ;
        RECT 57.065 152.945 57.405 153.915 ;
        RECT 57.575 152.945 57.745 154.085 ;
        RECT 58.015 153.285 58.265 154.085 ;
        RECT 58.910 153.115 59.240 153.915 ;
        RECT 59.540 153.285 59.870 154.085 ;
        RECT 60.040 153.115 60.370 153.915 ;
        RECT 57.935 152.945 60.370 153.115 ;
        RECT 61.205 153.325 61.720 153.735 ;
        RECT 61.955 153.325 62.125 154.085 ;
        RECT 62.295 153.745 64.325 153.915 ;
        RECT 51.065 152.275 51.235 152.445 ;
        RECT 50.625 151.865 50.895 152.210 ;
        RECT 51.065 152.105 52.675 152.275 ;
        RECT 52.860 152.205 53.210 152.775 ;
        RECT 53.385 152.385 53.560 152.945 ;
        RECT 54.255 152.695 54.425 152.945 ;
        RECT 53.730 152.525 54.425 152.695 ;
        RECT 54.600 152.525 55.020 152.725 ;
        RECT 55.190 152.525 55.520 152.725 ;
        RECT 55.690 152.525 56.020 152.725 ;
        RECT 53.385 152.335 53.615 152.385 ;
        RECT 51.085 151.535 51.465 151.935 ;
        RECT 51.635 151.755 51.805 152.105 ;
        RECT 51.975 151.535 52.305 151.935 ;
        RECT 52.505 151.755 52.675 152.105 ;
        RECT 52.875 151.535 53.205 152.035 ;
        RECT 53.385 151.705 53.725 152.335 ;
        RECT 53.895 151.535 54.145 152.335 ;
        RECT 54.335 152.185 55.560 152.355 ;
        RECT 54.335 151.705 54.665 152.185 ;
        RECT 54.835 151.535 55.060 151.995 ;
        RECT 55.230 151.705 55.560 152.185 ;
        RECT 56.190 152.315 56.360 152.945 ;
        RECT 57.065 152.895 57.295 152.945 ;
        RECT 56.545 152.525 56.895 152.775 ;
        RECT 57.065 152.335 57.240 152.895 ;
        RECT 57.935 152.695 58.105 152.945 ;
        RECT 57.410 152.525 58.105 152.695 ;
        RECT 58.280 152.525 58.700 152.725 ;
        RECT 58.870 152.525 59.200 152.725 ;
        RECT 59.370 152.525 59.700 152.725 ;
        RECT 56.190 151.705 56.690 152.315 ;
        RECT 57.065 151.705 57.405 152.335 ;
        RECT 57.575 151.535 57.825 152.335 ;
        RECT 58.015 152.185 59.240 152.355 ;
        RECT 58.015 151.705 58.345 152.185 ;
        RECT 58.515 151.535 58.740 151.995 ;
        RECT 58.910 151.705 59.240 152.185 ;
        RECT 59.870 152.315 60.040 152.945 ;
        RECT 60.225 152.525 60.575 152.775 ;
        RECT 61.205 152.515 61.545 153.325 ;
        RECT 62.295 153.080 62.465 153.745 ;
        RECT 62.860 153.405 63.985 153.575 ;
        RECT 61.715 152.890 62.465 153.080 ;
        RECT 62.635 153.065 63.645 153.235 ;
        RECT 61.205 152.345 62.435 152.515 ;
        RECT 59.870 151.705 60.370 152.315 ;
        RECT 61.480 151.740 61.725 152.345 ;
        RECT 61.945 151.535 62.455 152.070 ;
        RECT 62.635 151.705 62.825 153.065 ;
        RECT 62.995 152.045 63.270 152.865 ;
        RECT 63.475 152.265 63.645 153.065 ;
        RECT 63.815 152.275 63.985 153.405 ;
        RECT 64.155 152.775 64.325 153.745 ;
        RECT 64.495 152.945 64.665 154.085 ;
        RECT 64.835 152.945 65.170 153.915 ;
        RECT 65.435 153.340 65.705 154.085 ;
        RECT 66.335 154.080 72.610 154.085 ;
        RECT 65.875 153.170 66.165 153.910 ;
        RECT 66.335 153.355 66.590 154.080 ;
        RECT 66.775 153.185 67.035 153.910 ;
        RECT 67.205 153.355 67.450 154.080 ;
        RECT 67.635 153.185 67.895 153.910 ;
        RECT 68.065 153.355 68.310 154.080 ;
        RECT 68.495 153.185 68.755 153.910 ;
        RECT 68.925 153.355 69.170 154.080 ;
        RECT 69.340 153.185 69.600 153.910 ;
        RECT 69.770 153.355 70.030 154.080 ;
        RECT 70.200 153.185 70.460 153.910 ;
        RECT 70.630 153.355 70.890 154.080 ;
        RECT 71.060 153.185 71.320 153.910 ;
        RECT 71.490 153.355 71.750 154.080 ;
        RECT 71.920 153.185 72.180 153.910 ;
        RECT 72.350 153.285 72.610 154.080 ;
        RECT 66.775 153.170 72.180 153.185 ;
        RECT 65.435 153.065 72.180 153.170 ;
        RECT 64.155 152.445 64.350 152.775 ;
        RECT 64.575 152.445 64.830 152.775 ;
        RECT 64.575 152.275 64.745 152.445 ;
        RECT 65.000 152.275 65.170 152.945 ;
        RECT 65.405 152.945 72.180 153.065 ;
        RECT 65.405 152.895 66.600 152.945 ;
        RECT 63.815 152.105 64.745 152.275 ;
        RECT 63.815 152.070 63.990 152.105 ;
        RECT 62.995 151.875 63.275 152.045 ;
        RECT 62.995 151.705 63.270 151.875 ;
        RECT 63.460 151.705 63.990 152.070 ;
        RECT 64.415 151.535 64.745 151.935 ;
        RECT 64.915 151.705 65.170 152.275 ;
        RECT 65.435 152.355 66.600 152.895 ;
        RECT 72.780 152.775 73.030 153.910 ;
        RECT 73.210 153.275 73.470 154.085 ;
        RECT 73.645 152.775 73.890 153.915 ;
        RECT 74.070 153.275 74.365 154.085 ;
        RECT 74.545 152.995 75.755 154.085 ;
        RECT 66.770 152.525 73.890 152.775 ;
        RECT 65.435 152.185 72.180 152.355 ;
        RECT 65.435 151.535 65.735 152.015 ;
        RECT 65.905 151.730 66.165 152.185 ;
        RECT 66.335 151.535 66.595 152.015 ;
        RECT 66.775 151.730 67.035 152.185 ;
        RECT 67.205 151.535 67.455 152.015 ;
        RECT 67.635 151.730 67.895 152.185 ;
        RECT 68.065 151.535 68.315 152.015 ;
        RECT 68.495 151.730 68.755 152.185 ;
        RECT 68.925 151.535 69.170 152.015 ;
        RECT 69.340 151.730 69.615 152.185 ;
        RECT 69.785 151.535 70.030 152.015 ;
        RECT 70.200 151.730 70.460 152.185 ;
        RECT 70.630 151.535 70.890 152.015 ;
        RECT 71.060 151.730 71.320 152.185 ;
        RECT 71.490 151.535 71.750 152.015 ;
        RECT 71.920 151.730 72.180 152.185 ;
        RECT 72.350 151.535 72.610 152.095 ;
        RECT 72.780 151.715 73.030 152.525 ;
        RECT 73.210 151.535 73.470 152.060 ;
        RECT 73.640 151.715 73.890 152.525 ;
        RECT 74.060 152.215 74.375 152.775 ;
        RECT 74.545 152.455 75.065 152.995 ;
        RECT 75.925 152.920 76.215 154.085 ;
        RECT 76.475 153.155 76.645 153.915 ;
        RECT 76.860 153.325 77.190 154.085 ;
        RECT 76.475 152.985 77.190 153.155 ;
        RECT 77.360 153.010 77.615 153.915 ;
        RECT 75.235 152.285 75.755 152.825 ;
        RECT 76.385 152.435 76.740 152.805 ;
        RECT 77.020 152.775 77.190 152.985 ;
        RECT 77.020 152.445 77.275 152.775 ;
        RECT 74.070 151.535 74.375 152.045 ;
        RECT 74.545 151.535 75.755 152.285 ;
        RECT 75.925 151.535 76.215 152.260 ;
        RECT 77.020 152.255 77.190 152.445 ;
        RECT 77.445 152.280 77.615 153.010 ;
        RECT 77.790 152.935 78.050 154.085 ;
        RECT 78.225 152.995 79.895 154.085 ;
        RECT 78.225 152.475 78.975 152.995 ;
        RECT 80.065 152.945 80.335 153.915 ;
        RECT 80.545 153.285 80.825 154.085 ;
        RECT 80.995 153.575 82.650 153.865 ;
        RECT 81.060 153.235 82.650 153.405 ;
        RECT 81.060 153.115 81.230 153.235 ;
        RECT 80.505 152.945 81.230 153.115 ;
        RECT 76.475 152.085 77.190 152.255 ;
        RECT 76.475 151.705 76.645 152.085 ;
        RECT 76.860 151.535 77.190 151.915 ;
        RECT 77.360 151.705 77.615 152.280 ;
        RECT 77.790 151.535 78.050 152.375 ;
        RECT 79.145 152.305 79.895 152.825 ;
        RECT 78.225 151.535 79.895 152.305 ;
        RECT 80.065 152.210 80.235 152.945 ;
        RECT 80.505 152.775 80.675 152.945 ;
        RECT 81.420 152.895 82.135 153.065 ;
        RECT 82.330 152.945 82.650 153.235 ;
        RECT 82.825 152.945 83.165 153.915 ;
        RECT 83.335 152.945 83.505 154.085 ;
        RECT 83.775 153.285 84.025 154.085 ;
        RECT 84.670 153.115 85.000 153.915 ;
        RECT 85.300 153.285 85.630 154.085 ;
        RECT 85.800 153.115 86.130 153.915 ;
        RECT 83.695 152.945 86.130 153.115 ;
        RECT 86.565 152.945 86.775 154.085 ;
        RECT 80.405 152.445 80.675 152.775 ;
        RECT 80.845 152.445 81.250 152.775 ;
        RECT 81.420 152.445 82.130 152.895 ;
        RECT 80.505 152.275 80.675 152.445 ;
        RECT 80.065 151.865 80.335 152.210 ;
        RECT 80.505 152.105 82.115 152.275 ;
        RECT 82.300 152.205 82.650 152.775 ;
        RECT 82.825 152.385 83.000 152.945 ;
        RECT 83.695 152.695 83.865 152.945 ;
        RECT 83.170 152.525 83.865 152.695 ;
        RECT 84.040 152.525 84.460 152.725 ;
        RECT 84.630 152.525 84.960 152.725 ;
        RECT 85.130 152.525 85.460 152.725 ;
        RECT 82.825 152.335 83.055 152.385 ;
        RECT 80.525 151.535 80.905 151.935 ;
        RECT 81.075 151.755 81.245 152.105 ;
        RECT 81.415 151.535 81.745 151.935 ;
        RECT 81.945 151.755 82.115 152.105 ;
        RECT 82.315 151.535 82.645 152.035 ;
        RECT 82.825 151.705 83.165 152.335 ;
        RECT 83.335 151.535 83.585 152.335 ;
        RECT 83.775 152.185 85.000 152.355 ;
        RECT 83.775 151.705 84.105 152.185 ;
        RECT 84.275 151.535 84.500 151.995 ;
        RECT 84.670 151.705 85.000 152.185 ;
        RECT 85.630 152.315 85.800 152.945 ;
        RECT 86.945 152.935 87.275 153.915 ;
        RECT 87.445 152.945 87.675 154.085 ;
        RECT 88.260 153.105 88.515 153.775 ;
        RECT 88.695 153.285 88.980 154.085 ;
        RECT 89.160 153.365 89.490 153.875 ;
        RECT 85.985 152.525 86.335 152.775 ;
        RECT 85.630 151.705 86.130 152.315 ;
        RECT 86.565 151.535 86.775 152.355 ;
        RECT 86.945 152.335 87.195 152.935 ;
        RECT 87.365 152.525 87.695 152.775 ;
        RECT 86.945 151.705 87.275 152.335 ;
        RECT 87.445 151.535 87.675 152.355 ;
        RECT 88.260 152.245 88.440 153.105 ;
        RECT 89.160 152.775 89.410 153.365 ;
        RECT 89.760 153.215 89.930 153.825 ;
        RECT 90.100 153.395 90.430 154.085 ;
        RECT 90.660 153.535 90.900 153.825 ;
        RECT 91.100 153.705 91.520 154.085 ;
        RECT 91.700 153.615 92.330 153.865 ;
        RECT 92.800 153.705 93.130 154.085 ;
        RECT 91.700 153.535 91.870 153.615 ;
        RECT 93.300 153.535 93.470 153.825 ;
        RECT 93.650 153.705 94.030 154.085 ;
        RECT 94.270 153.700 95.100 153.870 ;
        RECT 90.660 153.365 91.870 153.535 ;
        RECT 88.610 152.445 89.410 152.775 ;
        RECT 88.260 152.045 88.515 152.245 ;
        RECT 88.175 151.875 88.515 152.045 ;
        RECT 88.260 151.715 88.515 151.875 ;
        RECT 88.695 151.535 88.980 151.995 ;
        RECT 89.160 151.795 89.410 152.445 ;
        RECT 89.610 153.195 89.930 153.215 ;
        RECT 89.610 153.025 91.530 153.195 ;
        RECT 89.610 152.130 89.800 153.025 ;
        RECT 91.700 152.855 91.870 153.365 ;
        RECT 92.040 153.105 92.560 153.415 ;
        RECT 89.970 152.685 91.870 152.855 ;
        RECT 89.970 152.625 90.300 152.685 ;
        RECT 90.450 152.455 90.780 152.515 ;
        RECT 90.120 152.185 90.780 152.455 ;
        RECT 89.610 151.800 89.930 152.130 ;
        RECT 90.110 151.535 90.770 152.015 ;
        RECT 90.970 151.925 91.140 152.685 ;
        RECT 92.040 152.515 92.220 152.925 ;
        RECT 91.310 152.345 91.640 152.465 ;
        RECT 92.390 152.345 92.560 153.105 ;
        RECT 91.310 152.175 92.560 152.345 ;
        RECT 92.730 153.285 94.100 153.535 ;
        RECT 92.730 152.515 92.920 153.285 ;
        RECT 93.850 153.025 94.100 153.285 ;
        RECT 93.090 152.855 93.340 153.015 ;
        RECT 94.270 152.855 94.440 153.700 ;
        RECT 95.335 153.415 95.505 153.915 ;
        RECT 95.675 153.585 96.005 154.085 ;
        RECT 94.610 153.025 95.110 153.405 ;
        RECT 95.335 153.245 96.030 153.415 ;
        RECT 93.090 152.685 94.440 152.855 ;
        RECT 94.020 152.645 94.440 152.685 ;
        RECT 92.730 152.175 93.150 152.515 ;
        RECT 93.440 152.185 93.850 152.515 ;
        RECT 90.970 151.755 91.820 151.925 ;
        RECT 92.380 151.535 92.700 151.995 ;
        RECT 92.900 151.745 93.150 152.175 ;
        RECT 93.440 151.535 93.850 151.975 ;
        RECT 94.020 151.915 94.190 152.645 ;
        RECT 94.360 152.095 94.710 152.465 ;
        RECT 94.890 152.155 95.110 153.025 ;
        RECT 95.280 152.455 95.690 153.075 ;
        RECT 95.860 152.275 96.030 153.245 ;
        RECT 95.335 152.085 96.030 152.275 ;
        RECT 94.020 151.715 95.035 151.915 ;
        RECT 95.335 151.755 95.505 152.085 ;
        RECT 95.675 151.535 96.005 151.915 ;
        RECT 96.220 151.795 96.445 153.915 ;
        RECT 96.615 153.585 96.945 154.085 ;
        RECT 97.115 153.415 97.285 153.915 ;
        RECT 96.620 153.245 97.285 153.415 ;
        RECT 97.545 153.325 98.060 153.735 ;
        RECT 98.295 153.325 98.465 154.085 ;
        RECT 98.635 153.745 100.665 153.915 ;
        RECT 96.620 152.255 96.850 153.245 ;
        RECT 97.020 152.425 97.370 153.075 ;
        RECT 97.545 152.515 97.885 153.325 ;
        RECT 98.635 153.080 98.805 153.745 ;
        RECT 99.200 153.405 100.325 153.575 ;
        RECT 98.055 152.890 98.805 153.080 ;
        RECT 98.975 153.065 99.985 153.235 ;
        RECT 97.545 152.345 98.775 152.515 ;
        RECT 96.620 152.085 97.285 152.255 ;
        RECT 96.615 151.535 96.945 151.915 ;
        RECT 97.115 151.795 97.285 152.085 ;
        RECT 97.820 151.740 98.065 152.345 ;
        RECT 98.285 151.535 98.795 152.070 ;
        RECT 98.975 151.705 99.165 153.065 ;
        RECT 99.335 152.385 99.610 152.865 ;
        RECT 99.335 152.215 99.615 152.385 ;
        RECT 99.815 152.265 99.985 153.065 ;
        RECT 100.155 152.275 100.325 153.405 ;
        RECT 100.495 152.775 100.665 153.745 ;
        RECT 100.835 152.945 101.005 154.085 ;
        RECT 101.175 152.945 101.510 153.915 ;
        RECT 100.495 152.445 100.690 152.775 ;
        RECT 100.915 152.445 101.170 152.775 ;
        RECT 100.915 152.275 101.085 152.445 ;
        RECT 101.340 152.275 101.510 152.945 ;
        RECT 101.685 152.920 101.975 154.085 ;
        RECT 102.205 152.945 102.415 154.085 ;
        RECT 102.585 152.935 102.915 153.915 ;
        RECT 103.085 152.945 103.315 154.085 ;
        RECT 103.615 153.155 103.785 153.915 ;
        RECT 103.965 153.325 104.295 154.085 ;
        RECT 103.615 152.985 104.280 153.155 ;
        RECT 104.465 153.010 104.735 153.915 ;
        RECT 99.335 151.705 99.610 152.215 ;
        RECT 100.155 152.105 101.085 152.275 ;
        RECT 100.155 152.070 100.330 152.105 ;
        RECT 99.800 151.705 100.330 152.070 ;
        RECT 100.755 151.535 101.085 151.935 ;
        RECT 101.255 151.705 101.510 152.275 ;
        RECT 101.685 151.535 101.975 152.260 ;
        RECT 102.205 151.535 102.415 152.355 ;
        RECT 102.585 152.335 102.835 152.935 ;
        RECT 104.110 152.840 104.280 152.985 ;
        RECT 103.005 152.525 103.335 152.775 ;
        RECT 103.545 152.435 103.875 152.805 ;
        RECT 104.110 152.510 104.395 152.840 ;
        RECT 102.585 151.705 102.915 152.335 ;
        RECT 103.085 151.535 103.315 152.355 ;
        RECT 104.110 152.255 104.280 152.510 ;
        RECT 103.615 152.085 104.280 152.255 ;
        RECT 104.565 152.210 104.735 153.010 ;
        RECT 105.570 153.115 105.900 153.915 ;
        RECT 106.070 153.285 106.400 154.085 ;
        RECT 106.700 153.115 107.030 153.915 ;
        RECT 107.675 153.285 107.925 154.085 ;
        RECT 105.570 152.945 108.005 153.115 ;
        RECT 108.195 152.945 108.365 154.085 ;
        RECT 108.535 152.945 108.875 153.915 ;
        RECT 109.250 153.115 109.580 153.915 ;
        RECT 109.750 153.285 110.080 154.085 ;
        RECT 110.380 153.115 110.710 153.915 ;
        RECT 111.355 153.285 111.605 154.085 ;
        RECT 109.250 152.945 111.685 153.115 ;
        RECT 111.875 152.945 112.045 154.085 ;
        RECT 112.215 152.945 112.555 153.915 ;
        RECT 105.365 152.525 105.715 152.775 ;
        RECT 105.900 152.315 106.070 152.945 ;
        RECT 106.240 152.525 106.570 152.725 ;
        RECT 106.740 152.525 107.070 152.725 ;
        RECT 107.240 152.525 107.660 152.725 ;
        RECT 107.835 152.695 108.005 152.945 ;
        RECT 107.835 152.525 108.530 152.695 ;
        RECT 103.615 151.705 103.785 152.085 ;
        RECT 103.965 151.535 104.295 151.915 ;
        RECT 104.475 151.705 104.735 152.210 ;
        RECT 105.570 151.705 106.070 152.315 ;
        RECT 106.700 152.185 107.925 152.355 ;
        RECT 108.700 152.335 108.875 152.945 ;
        RECT 109.045 152.525 109.395 152.775 ;
        RECT 106.700 151.705 107.030 152.185 ;
        RECT 107.200 151.535 107.425 151.995 ;
        RECT 107.595 151.705 107.925 152.185 ;
        RECT 108.115 151.535 108.365 152.335 ;
        RECT 108.535 151.705 108.875 152.335 ;
        RECT 109.580 152.315 109.750 152.945 ;
        RECT 109.920 152.525 110.250 152.725 ;
        RECT 110.420 152.525 110.750 152.725 ;
        RECT 110.920 152.525 111.340 152.725 ;
        RECT 111.515 152.695 111.685 152.945 ;
        RECT 111.515 152.525 112.210 152.695 ;
        RECT 109.250 151.705 109.750 152.315 ;
        RECT 110.380 152.185 111.605 152.355 ;
        RECT 112.380 152.335 112.555 152.945 ;
        RECT 112.725 153.325 113.240 153.735 ;
        RECT 113.475 153.325 113.645 154.085 ;
        RECT 113.815 153.745 115.845 153.915 ;
        RECT 112.725 152.515 113.065 153.325 ;
        RECT 113.815 153.080 113.985 153.745 ;
        RECT 114.380 153.405 115.505 153.575 ;
        RECT 113.235 152.890 113.985 153.080 ;
        RECT 114.155 153.065 115.165 153.235 ;
        RECT 112.725 152.345 113.955 152.515 ;
        RECT 110.380 151.705 110.710 152.185 ;
        RECT 110.880 151.535 111.105 151.995 ;
        RECT 111.275 151.705 111.605 152.185 ;
        RECT 111.795 151.535 112.045 152.335 ;
        RECT 112.215 151.705 112.555 152.335 ;
        RECT 113.000 151.740 113.245 152.345 ;
        RECT 113.465 151.535 113.975 152.070 ;
        RECT 114.155 151.705 114.345 153.065 ;
        RECT 114.515 152.045 114.790 152.865 ;
        RECT 114.995 152.265 115.165 153.065 ;
        RECT 115.335 152.275 115.505 153.405 ;
        RECT 115.675 152.775 115.845 153.745 ;
        RECT 116.015 152.945 116.185 154.085 ;
        RECT 116.355 152.945 116.690 153.915 ;
        RECT 115.675 152.445 115.870 152.775 ;
        RECT 116.095 152.445 116.350 152.775 ;
        RECT 116.095 152.275 116.265 152.445 ;
        RECT 116.520 152.275 116.690 152.945 ;
        RECT 116.865 153.325 117.380 153.735 ;
        RECT 117.615 153.325 117.785 154.085 ;
        RECT 117.955 153.745 119.985 153.915 ;
        RECT 116.865 152.515 117.205 153.325 ;
        RECT 117.955 153.080 118.125 153.745 ;
        RECT 118.520 153.405 119.645 153.575 ;
        RECT 117.375 152.890 118.125 153.080 ;
        RECT 118.295 153.065 119.305 153.235 ;
        RECT 116.865 152.345 118.095 152.515 ;
        RECT 115.335 152.105 116.265 152.275 ;
        RECT 115.335 152.070 115.510 152.105 ;
        RECT 114.515 151.875 114.795 152.045 ;
        RECT 114.515 151.705 114.790 151.875 ;
        RECT 114.980 151.705 115.510 152.070 ;
        RECT 115.935 151.535 116.265 151.935 ;
        RECT 116.435 151.705 116.690 152.275 ;
        RECT 117.140 151.740 117.385 152.345 ;
        RECT 117.605 151.535 118.115 152.070 ;
        RECT 118.295 151.705 118.485 153.065 ;
        RECT 118.655 152.725 118.930 152.865 ;
        RECT 118.655 152.555 118.935 152.725 ;
        RECT 118.655 151.705 118.930 152.555 ;
        RECT 119.135 152.265 119.305 153.065 ;
        RECT 119.475 152.275 119.645 153.405 ;
        RECT 119.815 152.775 119.985 153.745 ;
        RECT 120.155 152.945 120.325 154.085 ;
        RECT 120.495 152.945 120.830 153.915 ;
        RECT 121.095 153.155 121.265 153.915 ;
        RECT 121.445 153.325 121.775 154.085 ;
        RECT 121.095 152.985 121.760 153.155 ;
        RECT 121.945 153.010 122.215 153.915 ;
        RECT 119.815 152.445 120.010 152.775 ;
        RECT 120.235 152.445 120.490 152.775 ;
        RECT 120.235 152.275 120.405 152.445 ;
        RECT 120.660 152.275 120.830 152.945 ;
        RECT 121.590 152.840 121.760 152.985 ;
        RECT 121.025 152.435 121.355 152.805 ;
        RECT 121.590 152.510 121.875 152.840 ;
        RECT 119.475 152.105 120.405 152.275 ;
        RECT 119.475 152.070 119.650 152.105 ;
        RECT 119.120 151.705 119.650 152.070 ;
        RECT 120.075 151.535 120.405 151.935 ;
        RECT 120.575 151.705 120.830 152.275 ;
        RECT 121.590 152.255 121.760 152.510 ;
        RECT 121.095 152.085 121.760 152.255 ;
        RECT 122.045 152.210 122.215 153.010 ;
        RECT 122.475 153.155 122.645 153.915 ;
        RECT 122.825 153.325 123.155 154.085 ;
        RECT 122.475 152.985 123.140 153.155 ;
        RECT 123.325 153.010 123.595 153.915 ;
        RECT 122.970 152.840 123.140 152.985 ;
        RECT 122.405 152.435 122.735 152.805 ;
        RECT 122.970 152.510 123.255 152.840 ;
        RECT 122.970 152.255 123.140 152.510 ;
        RECT 121.095 151.705 121.265 152.085 ;
        RECT 121.445 151.535 121.775 151.915 ;
        RECT 121.955 151.705 122.215 152.210 ;
        RECT 122.475 152.085 123.140 152.255 ;
        RECT 123.425 152.210 123.595 153.010 ;
        RECT 123.765 152.995 126.355 154.085 ;
        RECT 126.525 152.995 127.735 154.085 ;
        RECT 123.765 152.475 124.975 152.995 ;
        RECT 125.145 152.305 126.355 152.825 ;
        RECT 126.525 152.455 127.045 152.995 ;
        RECT 122.475 151.705 122.645 152.085 ;
        RECT 122.825 151.535 123.155 151.915 ;
        RECT 123.335 151.705 123.595 152.210 ;
        RECT 123.765 151.535 126.355 152.305 ;
        RECT 127.215 152.285 127.735 152.825 ;
        RECT 126.525 151.535 127.735 152.285 ;
        RECT 20.640 151.365 127.820 151.535 ;
        RECT 20.725 150.615 21.935 151.365 ;
        RECT 22.480 151.025 22.735 151.185 ;
        RECT 22.395 150.855 22.735 151.025 ;
        RECT 22.915 150.905 23.200 151.365 ;
        RECT 22.480 150.655 22.735 150.855 ;
        RECT 20.725 150.075 21.245 150.615 ;
        RECT 21.415 149.905 21.935 150.445 ;
        RECT 20.725 148.815 21.935 149.905 ;
        RECT 22.480 149.795 22.660 150.655 ;
        RECT 23.380 150.455 23.630 151.105 ;
        RECT 22.830 150.125 23.630 150.455 ;
        RECT 22.480 149.125 22.735 149.795 ;
        RECT 22.915 148.815 23.200 149.615 ;
        RECT 23.380 149.535 23.630 150.125 ;
        RECT 23.830 150.770 24.150 151.100 ;
        RECT 24.330 150.885 24.990 151.365 ;
        RECT 25.190 150.975 26.040 151.145 ;
        RECT 23.830 149.875 24.020 150.770 ;
        RECT 24.340 150.445 25.000 150.715 ;
        RECT 24.670 150.385 25.000 150.445 ;
        RECT 24.190 150.215 24.520 150.275 ;
        RECT 25.190 150.215 25.360 150.975 ;
        RECT 26.600 150.905 26.920 151.365 ;
        RECT 27.120 150.725 27.370 151.155 ;
        RECT 27.660 150.925 28.070 151.365 ;
        RECT 28.240 150.985 29.255 151.185 ;
        RECT 25.530 150.555 26.780 150.725 ;
        RECT 25.530 150.435 25.860 150.555 ;
        RECT 24.190 150.045 26.090 150.215 ;
        RECT 23.830 149.705 25.750 149.875 ;
        RECT 23.830 149.685 24.150 149.705 ;
        RECT 23.380 149.025 23.710 149.535 ;
        RECT 23.980 149.075 24.150 149.685 ;
        RECT 25.920 149.535 26.090 150.045 ;
        RECT 26.260 149.975 26.440 150.385 ;
        RECT 26.610 149.795 26.780 150.555 ;
        RECT 24.320 148.815 24.650 149.505 ;
        RECT 24.880 149.365 26.090 149.535 ;
        RECT 26.260 149.485 26.780 149.795 ;
        RECT 26.950 150.385 27.370 150.725 ;
        RECT 27.660 150.385 28.070 150.715 ;
        RECT 26.950 149.615 27.140 150.385 ;
        RECT 28.240 150.255 28.410 150.985 ;
        RECT 29.555 150.815 29.725 151.145 ;
        RECT 29.895 150.985 30.225 151.365 ;
        RECT 28.580 150.435 28.930 150.805 ;
        RECT 28.240 150.215 28.660 150.255 ;
        RECT 27.310 150.045 28.660 150.215 ;
        RECT 27.310 149.885 27.560 150.045 ;
        RECT 28.070 149.615 28.320 149.875 ;
        RECT 26.950 149.365 28.320 149.615 ;
        RECT 24.880 149.075 25.120 149.365 ;
        RECT 25.920 149.285 26.090 149.365 ;
        RECT 25.320 148.815 25.740 149.195 ;
        RECT 25.920 149.035 26.550 149.285 ;
        RECT 27.020 148.815 27.350 149.195 ;
        RECT 27.520 149.075 27.690 149.365 ;
        RECT 28.490 149.200 28.660 150.045 ;
        RECT 29.110 149.875 29.330 150.745 ;
        RECT 29.555 150.625 30.250 150.815 ;
        RECT 28.830 149.495 29.330 149.875 ;
        RECT 29.500 149.825 29.910 150.445 ;
        RECT 30.080 149.655 30.250 150.625 ;
        RECT 29.555 149.485 30.250 149.655 ;
        RECT 27.870 148.815 28.250 149.195 ;
        RECT 28.490 149.030 29.320 149.200 ;
        RECT 29.555 148.985 29.725 149.485 ;
        RECT 29.895 148.815 30.225 149.315 ;
        RECT 30.440 148.985 30.665 151.105 ;
        RECT 30.835 150.985 31.165 151.365 ;
        RECT 31.335 150.815 31.505 151.105 ;
        RECT 30.840 150.645 31.505 150.815 ;
        RECT 30.840 149.655 31.070 150.645 ;
        RECT 32.040 150.555 32.285 151.160 ;
        RECT 32.505 150.830 33.015 151.365 ;
        RECT 31.240 149.825 31.590 150.475 ;
        RECT 31.765 150.385 32.995 150.555 ;
        RECT 30.840 149.485 31.505 149.655 ;
        RECT 30.835 148.815 31.165 149.315 ;
        RECT 31.335 148.985 31.505 149.485 ;
        RECT 31.765 149.575 32.105 150.385 ;
        RECT 32.275 149.820 33.025 150.010 ;
        RECT 31.765 149.165 32.280 149.575 ;
        RECT 32.515 148.815 32.685 149.575 ;
        RECT 32.855 149.155 33.025 149.820 ;
        RECT 33.195 149.835 33.385 151.195 ;
        RECT 33.555 150.685 33.830 151.195 ;
        RECT 34.020 150.830 34.550 151.195 ;
        RECT 34.975 150.965 35.305 151.365 ;
        RECT 34.375 150.795 34.550 150.830 ;
        RECT 33.555 150.515 33.835 150.685 ;
        RECT 33.555 150.035 33.830 150.515 ;
        RECT 34.035 149.835 34.205 150.635 ;
        RECT 33.195 149.665 34.205 149.835 ;
        RECT 34.375 150.625 35.305 150.795 ;
        RECT 35.475 150.625 35.730 151.195 ;
        RECT 34.375 149.495 34.545 150.625 ;
        RECT 35.135 150.455 35.305 150.625 ;
        RECT 33.420 149.325 34.545 149.495 ;
        RECT 34.715 150.125 34.910 150.455 ;
        RECT 35.135 150.125 35.390 150.455 ;
        RECT 34.715 149.155 34.885 150.125 ;
        RECT 35.560 149.955 35.730 150.625 ;
        RECT 32.855 148.985 34.885 149.155 ;
        RECT 35.055 148.815 35.225 149.955 ;
        RECT 35.395 148.985 35.730 149.955 ;
        RECT 35.905 150.690 36.165 151.195 ;
        RECT 36.345 150.985 36.675 151.365 ;
        RECT 36.855 150.815 37.025 151.195 ;
        RECT 35.905 149.890 36.075 150.690 ;
        RECT 36.360 150.645 37.025 150.815 ;
        RECT 36.360 150.390 36.530 150.645 ;
        RECT 37.285 150.640 37.575 151.365 ;
        RECT 37.745 150.595 39.415 151.365 ;
        RECT 36.245 150.060 36.530 150.390 ;
        RECT 36.765 150.095 37.095 150.465 ;
        RECT 36.360 149.915 36.530 150.060 ;
        RECT 35.905 148.985 36.175 149.890 ;
        RECT 36.360 149.745 37.025 149.915 ;
        RECT 36.345 148.815 36.675 149.575 ;
        RECT 36.855 148.985 37.025 149.745 ;
        RECT 37.285 148.815 37.575 149.980 ;
        RECT 37.745 149.905 38.495 150.425 ;
        RECT 38.665 150.075 39.415 150.595 ;
        RECT 39.585 150.565 39.925 151.195 ;
        RECT 40.095 150.565 40.345 151.365 ;
        RECT 40.535 150.715 40.865 151.195 ;
        RECT 41.035 150.905 41.260 151.365 ;
        RECT 41.430 150.715 41.760 151.195 ;
        RECT 39.585 149.955 39.760 150.565 ;
        RECT 40.535 150.545 41.760 150.715 ;
        RECT 42.390 150.585 42.890 151.195 ;
        RECT 39.930 150.205 40.625 150.375 ;
        RECT 40.455 149.955 40.625 150.205 ;
        RECT 40.800 150.175 41.220 150.375 ;
        RECT 41.390 150.175 41.720 150.375 ;
        RECT 41.890 150.175 42.220 150.375 ;
        RECT 42.390 149.955 42.560 150.585 ;
        RECT 43.265 150.565 43.605 151.195 ;
        RECT 43.775 150.565 44.025 151.365 ;
        RECT 44.215 150.715 44.545 151.195 ;
        RECT 44.715 150.905 44.940 151.365 ;
        RECT 45.110 150.715 45.440 151.195 ;
        RECT 42.745 150.125 43.095 150.375 ;
        RECT 43.265 149.955 43.440 150.565 ;
        RECT 44.215 150.545 45.440 150.715 ;
        RECT 46.070 150.585 46.570 151.195 ;
        RECT 46.945 150.615 48.155 151.365 ;
        RECT 43.610 150.205 44.305 150.375 ;
        RECT 44.135 149.955 44.305 150.205 ;
        RECT 44.480 150.175 44.900 150.375 ;
        RECT 45.070 150.175 45.400 150.375 ;
        RECT 45.570 150.175 45.900 150.375 ;
        RECT 46.070 149.955 46.240 150.585 ;
        RECT 46.425 150.125 46.775 150.375 ;
        RECT 37.745 148.815 39.415 149.905 ;
        RECT 39.585 148.985 39.925 149.955 ;
        RECT 40.095 148.815 40.265 149.955 ;
        RECT 40.455 149.785 42.890 149.955 ;
        RECT 40.535 148.815 40.785 149.615 ;
        RECT 41.430 148.985 41.760 149.785 ;
        RECT 42.060 148.815 42.390 149.615 ;
        RECT 42.560 148.985 42.890 149.785 ;
        RECT 43.265 148.985 43.605 149.955 ;
        RECT 43.775 148.815 43.945 149.955 ;
        RECT 44.135 149.785 46.570 149.955 ;
        RECT 44.215 148.815 44.465 149.615 ;
        RECT 45.110 148.985 45.440 149.785 ;
        RECT 45.740 148.815 46.070 149.615 ;
        RECT 46.240 148.985 46.570 149.785 ;
        RECT 46.945 149.905 47.465 150.445 ;
        RECT 47.635 150.075 48.155 150.615 ;
        RECT 48.325 150.595 51.835 151.365 ;
        RECT 52.010 150.820 57.355 151.365 ;
        RECT 57.530 150.820 62.875 151.365 ;
        RECT 48.325 149.905 50.015 150.425 ;
        RECT 50.185 150.075 51.835 150.595 ;
        RECT 46.945 148.815 48.155 149.905 ;
        RECT 48.325 148.815 51.835 149.905 ;
        RECT 53.600 149.250 53.950 150.500 ;
        RECT 55.430 149.990 55.770 150.820 ;
        RECT 59.120 149.250 59.470 150.500 ;
        RECT 60.950 149.990 61.290 150.820 ;
        RECT 63.045 150.640 63.335 151.365 ;
        RECT 63.965 150.595 66.555 151.365 ;
        RECT 52.010 148.815 57.355 149.250 ;
        RECT 57.530 148.815 62.875 149.250 ;
        RECT 63.045 148.815 63.335 149.980 ;
        RECT 63.965 149.905 65.175 150.425 ;
        RECT 65.345 150.075 66.555 150.595 ;
        RECT 66.765 150.545 66.995 151.365 ;
        RECT 67.165 150.565 67.495 151.195 ;
        RECT 66.745 150.125 67.075 150.375 ;
        RECT 67.245 149.965 67.495 150.565 ;
        RECT 67.665 150.545 67.875 151.365 ;
        RECT 68.565 150.595 70.235 151.365 ;
        RECT 70.495 150.815 70.665 151.195 ;
        RECT 70.845 150.985 71.175 151.365 ;
        RECT 70.495 150.645 71.160 150.815 ;
        RECT 71.355 150.690 71.615 151.195 ;
        RECT 63.965 148.815 66.555 149.905 ;
        RECT 66.765 148.815 66.995 149.955 ;
        RECT 67.165 148.985 67.495 149.965 ;
        RECT 67.665 148.815 67.875 149.955 ;
        RECT 68.565 149.905 69.315 150.425 ;
        RECT 69.485 150.075 70.235 150.595 ;
        RECT 70.425 150.095 70.755 150.465 ;
        RECT 70.990 150.390 71.160 150.645 ;
        RECT 70.990 150.060 71.275 150.390 ;
        RECT 70.990 149.915 71.160 150.060 ;
        RECT 68.565 148.815 70.235 149.905 ;
        RECT 70.495 149.745 71.160 149.915 ;
        RECT 71.445 149.890 71.615 150.690 ;
        RECT 71.790 150.525 72.050 151.365 ;
        RECT 72.225 150.620 72.480 151.195 ;
        RECT 72.650 150.985 72.980 151.365 ;
        RECT 73.195 150.815 73.365 151.195 ;
        RECT 72.650 150.645 73.365 150.815 ;
        RECT 73.715 150.815 73.885 151.195 ;
        RECT 74.100 150.985 74.430 151.365 ;
        RECT 73.715 150.645 74.430 150.815 ;
        RECT 70.495 148.985 70.665 149.745 ;
        RECT 70.845 148.815 71.175 149.575 ;
        RECT 71.345 148.985 71.615 149.890 ;
        RECT 71.790 148.815 72.050 149.965 ;
        RECT 72.225 149.890 72.395 150.620 ;
        RECT 72.650 150.455 72.820 150.645 ;
        RECT 72.565 150.125 72.820 150.455 ;
        RECT 72.650 149.915 72.820 150.125 ;
        RECT 73.100 150.095 73.455 150.465 ;
        RECT 73.625 150.095 73.980 150.465 ;
        RECT 74.260 150.455 74.430 150.645 ;
        RECT 74.600 150.620 74.855 151.195 ;
        RECT 74.260 150.125 74.515 150.455 ;
        RECT 74.260 149.915 74.430 150.125 ;
        RECT 72.225 148.985 72.480 149.890 ;
        RECT 72.650 149.745 73.365 149.915 ;
        RECT 72.650 148.815 72.980 149.575 ;
        RECT 73.195 148.985 73.365 149.745 ;
        RECT 73.715 149.745 74.430 149.915 ;
        RECT 74.685 149.890 74.855 150.620 ;
        RECT 75.030 150.525 75.290 151.365 ;
        RECT 75.465 150.595 78.055 151.365 ;
        RECT 73.715 148.985 73.885 149.745 ;
        RECT 74.100 148.815 74.430 149.575 ;
        RECT 74.600 148.985 74.855 149.890 ;
        RECT 75.030 148.815 75.290 149.965 ;
        RECT 75.465 149.905 76.675 150.425 ;
        RECT 76.845 150.075 78.055 150.595 ;
        RECT 78.225 150.690 78.495 151.035 ;
        RECT 78.685 150.965 79.065 151.365 ;
        RECT 79.235 150.795 79.405 151.145 ;
        RECT 79.575 150.965 79.905 151.365 ;
        RECT 80.105 150.795 80.275 151.145 ;
        RECT 80.475 150.865 80.805 151.365 ;
        RECT 78.225 149.955 78.395 150.690 ;
        RECT 78.665 150.625 80.275 150.795 ;
        RECT 78.665 150.455 78.835 150.625 ;
        RECT 78.565 150.125 78.835 150.455 ;
        RECT 79.005 150.125 79.410 150.455 ;
        RECT 78.665 149.955 78.835 150.125 ;
        RECT 75.465 148.815 78.055 149.905 ;
        RECT 78.225 148.985 78.495 149.955 ;
        RECT 78.665 149.785 79.390 149.955 ;
        RECT 79.580 149.835 80.290 150.455 ;
        RECT 80.460 150.125 80.810 150.695 ;
        RECT 80.985 150.565 81.325 151.195 ;
        RECT 81.495 150.565 81.745 151.365 ;
        RECT 81.935 150.715 82.265 151.195 ;
        RECT 82.435 150.905 82.660 151.365 ;
        RECT 82.830 150.715 83.160 151.195 ;
        RECT 80.985 150.515 81.215 150.565 ;
        RECT 81.935 150.545 83.160 150.715 ;
        RECT 83.790 150.585 84.290 151.195 ;
        RECT 80.985 149.955 81.160 150.515 ;
        RECT 81.330 150.205 82.025 150.375 ;
        RECT 81.855 149.955 82.025 150.205 ;
        RECT 82.200 150.175 82.620 150.375 ;
        RECT 82.790 150.175 83.120 150.375 ;
        RECT 83.290 150.175 83.620 150.375 ;
        RECT 83.790 149.955 83.960 150.585 ;
        RECT 84.940 150.555 85.185 151.160 ;
        RECT 85.405 150.830 85.915 151.365 ;
        RECT 84.665 150.385 85.895 150.555 ;
        RECT 84.145 150.125 84.495 150.375 ;
        RECT 79.220 149.665 79.390 149.785 ;
        RECT 80.490 149.665 80.810 149.955 ;
        RECT 78.705 148.815 78.985 149.615 ;
        RECT 79.220 149.495 80.810 149.665 ;
        RECT 79.155 149.035 80.810 149.325 ;
        RECT 80.985 148.985 81.325 149.955 ;
        RECT 81.495 148.815 81.665 149.955 ;
        RECT 81.855 149.785 84.290 149.955 ;
        RECT 81.935 148.815 82.185 149.615 ;
        RECT 82.830 148.985 83.160 149.785 ;
        RECT 83.460 148.815 83.790 149.615 ;
        RECT 83.960 148.985 84.290 149.785 ;
        RECT 84.665 149.575 85.005 150.385 ;
        RECT 85.175 149.820 85.925 150.010 ;
        RECT 84.665 149.165 85.180 149.575 ;
        RECT 85.415 148.815 85.585 149.575 ;
        RECT 85.755 149.155 85.925 149.820 ;
        RECT 86.095 149.835 86.285 151.195 ;
        RECT 86.455 150.345 86.730 151.195 ;
        RECT 86.920 150.830 87.450 151.195 ;
        RECT 87.875 150.965 88.205 151.365 ;
        RECT 87.275 150.795 87.450 150.830 ;
        RECT 86.455 150.175 86.735 150.345 ;
        RECT 86.455 150.035 86.730 150.175 ;
        RECT 86.935 149.835 87.105 150.635 ;
        RECT 86.095 149.665 87.105 149.835 ;
        RECT 87.275 150.625 88.205 150.795 ;
        RECT 88.375 150.625 88.630 151.195 ;
        RECT 88.805 150.640 89.095 151.365 ;
        RECT 87.275 149.495 87.445 150.625 ;
        RECT 88.035 150.455 88.205 150.625 ;
        RECT 86.320 149.325 87.445 149.495 ;
        RECT 87.615 150.125 87.810 150.455 ;
        RECT 88.035 150.125 88.290 150.455 ;
        RECT 87.615 149.155 87.785 150.125 ;
        RECT 88.460 149.955 88.630 150.625 ;
        RECT 89.540 150.555 89.785 151.160 ;
        RECT 90.005 150.830 90.515 151.365 ;
        RECT 89.265 150.385 90.495 150.555 ;
        RECT 85.755 148.985 87.785 149.155 ;
        RECT 87.955 148.815 88.125 149.955 ;
        RECT 88.295 148.985 88.630 149.955 ;
        RECT 88.805 148.815 89.095 149.980 ;
        RECT 89.265 149.575 89.605 150.385 ;
        RECT 89.775 149.820 90.525 150.010 ;
        RECT 89.265 149.165 89.780 149.575 ;
        RECT 90.015 148.815 90.185 149.575 ;
        RECT 90.355 149.155 90.525 149.820 ;
        RECT 90.695 149.835 90.885 151.195 ;
        RECT 91.055 150.685 91.330 151.195 ;
        RECT 91.520 150.830 92.050 151.195 ;
        RECT 92.475 150.965 92.805 151.365 ;
        RECT 91.875 150.795 92.050 150.830 ;
        RECT 91.055 150.515 91.335 150.685 ;
        RECT 91.055 150.035 91.330 150.515 ;
        RECT 91.535 149.835 91.705 150.635 ;
        RECT 90.695 149.665 91.705 149.835 ;
        RECT 91.875 150.625 92.805 150.795 ;
        RECT 92.975 150.625 93.230 151.195 ;
        RECT 93.495 150.815 93.665 151.195 ;
        RECT 93.845 150.985 94.175 151.365 ;
        RECT 93.495 150.645 94.160 150.815 ;
        RECT 94.355 150.690 94.615 151.195 ;
        RECT 91.875 149.495 92.045 150.625 ;
        RECT 92.635 150.455 92.805 150.625 ;
        RECT 90.920 149.325 92.045 149.495 ;
        RECT 92.215 150.125 92.410 150.455 ;
        RECT 92.635 150.125 92.890 150.455 ;
        RECT 92.215 149.155 92.385 150.125 ;
        RECT 93.060 149.955 93.230 150.625 ;
        RECT 93.425 150.095 93.755 150.465 ;
        RECT 93.990 150.390 94.160 150.645 ;
        RECT 90.355 148.985 92.385 149.155 ;
        RECT 92.555 148.815 92.725 149.955 ;
        RECT 92.895 148.985 93.230 149.955 ;
        RECT 93.990 150.060 94.275 150.390 ;
        RECT 93.990 149.915 94.160 150.060 ;
        RECT 93.495 149.745 94.160 149.915 ;
        RECT 94.445 149.890 94.615 150.690 ;
        RECT 94.875 150.815 95.045 151.195 ;
        RECT 95.225 150.985 95.555 151.365 ;
        RECT 94.875 150.645 95.540 150.815 ;
        RECT 95.735 150.690 95.995 151.195 ;
        RECT 94.805 150.095 95.135 150.465 ;
        RECT 95.370 150.390 95.540 150.645 ;
        RECT 95.370 150.060 95.655 150.390 ;
        RECT 95.370 149.915 95.540 150.060 ;
        RECT 93.495 148.985 93.665 149.745 ;
        RECT 93.845 148.815 94.175 149.575 ;
        RECT 94.345 148.985 94.615 149.890 ;
        RECT 94.875 149.745 95.540 149.915 ;
        RECT 95.825 149.890 95.995 150.690 ;
        RECT 96.625 150.595 98.295 151.365 ;
        RECT 94.875 148.985 95.045 149.745 ;
        RECT 95.225 148.815 95.555 149.575 ;
        RECT 95.725 148.985 95.995 149.890 ;
        RECT 96.625 149.905 97.375 150.425 ;
        RECT 97.545 150.075 98.295 150.595 ;
        RECT 98.470 150.655 98.725 151.185 ;
        RECT 98.895 150.905 99.200 151.365 ;
        RECT 99.445 150.985 100.515 151.155 ;
        RECT 98.470 150.005 98.680 150.655 ;
        RECT 99.445 150.630 99.765 150.985 ;
        RECT 99.440 150.455 99.765 150.630 ;
        RECT 98.850 150.155 99.765 150.455 ;
        RECT 99.935 150.415 100.175 150.815 ;
        RECT 100.345 150.755 100.515 150.985 ;
        RECT 100.685 150.925 100.875 151.365 ;
        RECT 101.045 150.915 101.995 151.195 ;
        RECT 102.215 151.005 102.565 151.175 ;
        RECT 100.345 150.585 100.875 150.755 ;
        RECT 98.850 150.125 99.590 150.155 ;
        RECT 96.625 148.815 98.295 149.905 ;
        RECT 98.470 149.125 98.725 150.005 ;
        RECT 98.895 148.815 99.200 149.955 ;
        RECT 99.420 149.535 99.590 150.125 ;
        RECT 99.935 150.045 100.475 150.415 ;
        RECT 100.655 150.305 100.875 150.585 ;
        RECT 101.045 150.135 101.215 150.915 ;
        RECT 100.810 149.965 101.215 150.135 ;
        RECT 101.385 150.125 101.735 150.745 ;
        RECT 100.810 149.875 100.980 149.965 ;
        RECT 101.905 149.955 102.115 150.745 ;
        RECT 99.760 149.705 100.980 149.875 ;
        RECT 101.440 149.795 102.115 149.955 ;
        RECT 99.420 149.365 100.220 149.535 ;
        RECT 99.540 148.815 99.870 149.195 ;
        RECT 100.050 149.075 100.220 149.365 ;
        RECT 100.810 149.325 100.980 149.705 ;
        RECT 101.150 149.785 102.115 149.795 ;
        RECT 102.305 150.615 102.565 151.005 ;
        RECT 102.775 150.905 103.105 151.365 ;
        RECT 103.980 150.975 104.835 151.145 ;
        RECT 105.040 150.975 105.535 151.145 ;
        RECT 105.705 151.005 106.035 151.365 ;
        RECT 102.305 149.925 102.475 150.615 ;
        RECT 102.645 150.265 102.815 150.445 ;
        RECT 102.985 150.435 103.775 150.685 ;
        RECT 103.980 150.265 104.150 150.975 ;
        RECT 104.320 150.465 104.675 150.685 ;
        RECT 102.645 150.095 104.335 150.265 ;
        RECT 101.150 149.495 101.610 149.785 ;
        RECT 102.305 149.755 103.805 149.925 ;
        RECT 102.305 149.615 102.475 149.755 ;
        RECT 101.915 149.445 102.475 149.615 ;
        RECT 100.390 148.815 100.640 149.275 ;
        RECT 100.810 148.985 101.680 149.325 ;
        RECT 101.915 148.985 102.085 149.445 ;
        RECT 102.920 149.415 103.995 149.585 ;
        RECT 102.255 148.815 102.625 149.275 ;
        RECT 102.920 149.075 103.090 149.415 ;
        RECT 103.260 148.815 103.590 149.245 ;
        RECT 103.825 149.075 103.995 149.415 ;
        RECT 104.165 149.315 104.335 150.095 ;
        RECT 104.505 149.875 104.675 150.465 ;
        RECT 104.845 150.065 105.195 150.685 ;
        RECT 104.505 149.485 104.970 149.875 ;
        RECT 105.365 149.615 105.535 150.975 ;
        RECT 105.705 149.785 106.165 150.835 ;
        RECT 105.140 149.445 105.535 149.615 ;
        RECT 105.140 149.315 105.310 149.445 ;
        RECT 104.165 148.985 104.845 149.315 ;
        RECT 105.060 148.985 105.310 149.315 ;
        RECT 105.480 148.815 105.730 149.275 ;
        RECT 105.900 149.000 106.225 149.785 ;
        RECT 106.395 148.985 106.565 151.105 ;
        RECT 106.735 150.985 107.065 151.365 ;
        RECT 107.235 150.815 107.490 151.105 ;
        RECT 106.740 150.645 107.490 150.815 ;
        RECT 106.740 149.655 106.970 150.645 ;
        RECT 107.665 150.615 108.875 151.365 ;
        RECT 107.140 149.825 107.490 150.475 ;
        RECT 107.665 149.905 108.185 150.445 ;
        RECT 108.355 150.075 108.875 150.615 ;
        RECT 109.045 150.565 109.385 151.195 ;
        RECT 109.555 150.565 109.805 151.365 ;
        RECT 109.995 150.715 110.325 151.195 ;
        RECT 110.495 150.905 110.720 151.365 ;
        RECT 110.890 150.715 111.220 151.195 ;
        RECT 109.045 149.955 109.220 150.565 ;
        RECT 109.995 150.545 111.220 150.715 ;
        RECT 111.850 150.585 112.350 151.195 ;
        RECT 112.725 150.595 114.395 151.365 ;
        RECT 114.565 150.640 114.855 151.365 ;
        RECT 115.025 150.595 116.695 151.365 ;
        RECT 109.390 150.205 110.085 150.375 ;
        RECT 109.915 149.955 110.085 150.205 ;
        RECT 110.260 150.175 110.680 150.375 ;
        RECT 110.850 150.175 111.180 150.375 ;
        RECT 111.350 150.175 111.680 150.375 ;
        RECT 111.850 149.955 112.020 150.585 ;
        RECT 112.205 150.125 112.555 150.375 ;
        RECT 106.740 149.485 107.490 149.655 ;
        RECT 106.735 148.815 107.065 149.315 ;
        RECT 107.235 148.985 107.490 149.485 ;
        RECT 107.665 148.815 108.875 149.905 ;
        RECT 109.045 148.985 109.385 149.955 ;
        RECT 109.555 148.815 109.725 149.955 ;
        RECT 109.915 149.785 112.350 149.955 ;
        RECT 109.995 148.815 110.245 149.615 ;
        RECT 110.890 148.985 111.220 149.785 ;
        RECT 111.520 148.815 111.850 149.615 ;
        RECT 112.020 148.985 112.350 149.785 ;
        RECT 112.725 149.905 113.475 150.425 ;
        RECT 113.645 150.075 114.395 150.595 ;
        RECT 112.725 148.815 114.395 149.905 ;
        RECT 114.565 148.815 114.855 149.980 ;
        RECT 115.025 149.905 115.775 150.425 ;
        RECT 115.945 150.075 116.695 150.595 ;
        RECT 117.240 150.655 117.495 151.185 ;
        RECT 117.675 150.905 117.960 151.365 ;
        RECT 115.025 148.815 116.695 149.905 ;
        RECT 117.240 149.795 117.420 150.655 ;
        RECT 118.140 150.455 118.390 151.105 ;
        RECT 117.590 150.125 118.390 150.455 ;
        RECT 117.240 149.325 117.495 149.795 ;
        RECT 117.155 149.155 117.495 149.325 ;
        RECT 117.240 149.125 117.495 149.155 ;
        RECT 117.675 148.815 117.960 149.615 ;
        RECT 118.140 149.535 118.390 150.125 ;
        RECT 118.590 150.770 118.910 151.100 ;
        RECT 119.090 150.885 119.750 151.365 ;
        RECT 119.950 150.975 120.800 151.145 ;
        RECT 118.590 149.875 118.780 150.770 ;
        RECT 119.100 150.445 119.760 150.715 ;
        RECT 119.430 150.385 119.760 150.445 ;
        RECT 118.950 150.215 119.280 150.275 ;
        RECT 119.950 150.215 120.120 150.975 ;
        RECT 121.360 150.905 121.680 151.365 ;
        RECT 121.880 150.725 122.130 151.155 ;
        RECT 122.420 150.925 122.830 151.365 ;
        RECT 123.000 150.985 124.015 151.185 ;
        RECT 120.290 150.555 121.540 150.725 ;
        RECT 120.290 150.435 120.620 150.555 ;
        RECT 118.950 150.045 120.850 150.215 ;
        RECT 118.590 149.705 120.510 149.875 ;
        RECT 118.590 149.685 118.910 149.705 ;
        RECT 118.140 149.025 118.470 149.535 ;
        RECT 118.740 149.075 118.910 149.685 ;
        RECT 120.680 149.535 120.850 150.045 ;
        RECT 121.020 149.975 121.200 150.385 ;
        RECT 121.370 149.795 121.540 150.555 ;
        RECT 119.080 148.815 119.410 149.505 ;
        RECT 119.640 149.365 120.850 149.535 ;
        RECT 121.020 149.485 121.540 149.795 ;
        RECT 121.710 150.385 122.130 150.725 ;
        RECT 122.420 150.385 122.830 150.715 ;
        RECT 121.710 149.615 121.900 150.385 ;
        RECT 123.000 150.255 123.170 150.985 ;
        RECT 124.315 150.815 124.485 151.145 ;
        RECT 124.655 150.985 124.985 151.365 ;
        RECT 123.340 150.435 123.690 150.805 ;
        RECT 123.000 150.215 123.420 150.255 ;
        RECT 122.070 150.045 123.420 150.215 ;
        RECT 122.070 149.885 122.320 150.045 ;
        RECT 122.830 149.615 123.080 149.875 ;
        RECT 121.710 149.365 123.080 149.615 ;
        RECT 119.640 149.075 119.880 149.365 ;
        RECT 120.680 149.285 120.850 149.365 ;
        RECT 120.080 148.815 120.500 149.195 ;
        RECT 120.680 149.035 121.310 149.285 ;
        RECT 121.780 148.815 122.110 149.195 ;
        RECT 122.280 149.075 122.450 149.365 ;
        RECT 123.250 149.200 123.420 150.045 ;
        RECT 123.870 149.875 124.090 150.745 ;
        RECT 124.315 150.625 125.010 150.815 ;
        RECT 123.590 149.495 124.090 149.875 ;
        RECT 124.260 149.825 124.670 150.445 ;
        RECT 124.840 149.655 125.010 150.625 ;
        RECT 124.315 149.485 125.010 149.655 ;
        RECT 122.630 148.815 123.010 149.195 ;
        RECT 123.250 149.030 124.080 149.200 ;
        RECT 124.315 148.985 124.485 149.485 ;
        RECT 124.655 148.815 124.985 149.315 ;
        RECT 125.200 148.985 125.425 151.105 ;
        RECT 125.595 150.985 125.925 151.365 ;
        RECT 126.095 150.815 126.265 151.105 ;
        RECT 125.600 150.645 126.265 150.815 ;
        RECT 125.600 149.655 125.830 150.645 ;
        RECT 126.525 150.615 127.735 151.365 ;
        RECT 126.000 149.825 126.350 150.475 ;
        RECT 126.525 149.905 127.045 150.445 ;
        RECT 127.215 150.075 127.735 150.615 ;
        RECT 125.600 149.485 126.265 149.655 ;
        RECT 125.595 148.815 125.925 149.315 ;
        RECT 126.095 148.985 126.265 149.485 ;
        RECT 126.525 148.815 127.735 149.905 ;
        RECT 20.640 148.645 127.820 148.815 ;
        RECT 20.725 147.555 21.935 148.645 ;
        RECT 20.725 146.845 21.245 147.385 ;
        RECT 21.415 147.015 21.935 147.555 ;
        RECT 22.565 147.555 24.235 148.645 ;
        RECT 22.565 147.035 23.315 147.555 ;
        RECT 24.405 147.480 24.695 148.645 ;
        RECT 25.385 147.505 25.595 148.645 ;
        RECT 25.765 147.495 26.095 148.475 ;
        RECT 26.265 147.505 26.495 148.645 ;
        RECT 27.080 148.305 27.335 148.335 ;
        RECT 26.995 148.135 27.335 148.305 ;
        RECT 27.080 147.665 27.335 148.135 ;
        RECT 27.515 147.845 27.800 148.645 ;
        RECT 27.980 147.925 28.310 148.435 ;
        RECT 23.485 146.865 24.235 147.385 ;
        RECT 20.725 146.095 21.935 146.845 ;
        RECT 22.565 146.095 24.235 146.865 ;
        RECT 24.405 146.095 24.695 146.820 ;
        RECT 25.385 146.095 25.595 146.915 ;
        RECT 25.765 146.895 26.015 147.495 ;
        RECT 26.185 147.085 26.515 147.335 ;
        RECT 25.765 146.265 26.095 146.895 ;
        RECT 26.265 146.095 26.495 146.915 ;
        RECT 27.080 146.805 27.260 147.665 ;
        RECT 27.980 147.335 28.230 147.925 ;
        RECT 28.580 147.775 28.750 148.385 ;
        RECT 28.920 147.955 29.250 148.645 ;
        RECT 29.480 148.095 29.720 148.385 ;
        RECT 29.920 148.265 30.340 148.645 ;
        RECT 30.520 148.175 31.150 148.425 ;
        RECT 31.620 148.265 31.950 148.645 ;
        RECT 30.520 148.095 30.690 148.175 ;
        RECT 32.120 148.095 32.290 148.385 ;
        RECT 32.470 148.265 32.850 148.645 ;
        RECT 33.090 148.260 33.920 148.430 ;
        RECT 29.480 147.925 30.690 148.095 ;
        RECT 27.430 147.005 28.230 147.335 ;
        RECT 27.080 146.275 27.335 146.805 ;
        RECT 27.515 146.095 27.800 146.555 ;
        RECT 27.980 146.355 28.230 147.005 ;
        RECT 28.430 147.755 28.750 147.775 ;
        RECT 28.430 147.585 30.350 147.755 ;
        RECT 28.430 146.690 28.620 147.585 ;
        RECT 30.520 147.415 30.690 147.925 ;
        RECT 30.860 147.665 31.380 147.975 ;
        RECT 28.790 147.245 30.690 147.415 ;
        RECT 28.790 147.185 29.120 147.245 ;
        RECT 29.270 147.015 29.600 147.075 ;
        RECT 28.940 146.745 29.600 147.015 ;
        RECT 28.430 146.360 28.750 146.690 ;
        RECT 28.930 146.095 29.590 146.575 ;
        RECT 29.790 146.485 29.960 147.245 ;
        RECT 30.860 147.075 31.040 147.485 ;
        RECT 30.130 146.905 30.460 147.025 ;
        RECT 31.210 146.905 31.380 147.665 ;
        RECT 30.130 146.735 31.380 146.905 ;
        RECT 31.550 147.845 32.920 148.095 ;
        RECT 31.550 147.075 31.740 147.845 ;
        RECT 32.670 147.585 32.920 147.845 ;
        RECT 31.910 147.415 32.160 147.575 ;
        RECT 33.090 147.415 33.260 148.260 ;
        RECT 34.155 147.975 34.325 148.475 ;
        RECT 34.495 148.145 34.825 148.645 ;
        RECT 33.430 147.585 33.930 147.965 ;
        RECT 34.155 147.805 34.850 147.975 ;
        RECT 31.910 147.245 33.260 147.415 ;
        RECT 32.840 147.205 33.260 147.245 ;
        RECT 31.550 146.735 31.970 147.075 ;
        RECT 32.260 146.745 32.670 147.075 ;
        RECT 29.790 146.315 30.640 146.485 ;
        RECT 31.200 146.095 31.520 146.555 ;
        RECT 31.720 146.305 31.970 146.735 ;
        RECT 32.260 146.095 32.670 146.535 ;
        RECT 32.840 146.475 33.010 147.205 ;
        RECT 33.180 146.655 33.530 147.025 ;
        RECT 33.710 146.715 33.930 147.585 ;
        RECT 34.100 147.015 34.510 147.635 ;
        RECT 34.680 146.835 34.850 147.805 ;
        RECT 34.155 146.645 34.850 146.835 ;
        RECT 32.840 146.275 33.855 146.475 ;
        RECT 34.155 146.315 34.325 146.645 ;
        RECT 34.495 146.095 34.825 146.475 ;
        RECT 35.040 146.355 35.265 148.475 ;
        RECT 35.435 148.145 35.765 148.645 ;
        RECT 35.935 147.975 36.105 148.475 ;
        RECT 35.440 147.805 36.105 147.975 ;
        RECT 35.440 146.815 35.670 147.805 ;
        RECT 35.840 146.985 36.190 147.635 ;
        RECT 36.825 147.555 39.415 148.645 ;
        RECT 36.825 147.035 38.035 147.555 ;
        RECT 39.585 147.505 39.925 148.475 ;
        RECT 40.095 147.505 40.265 148.645 ;
        RECT 40.535 147.845 40.785 148.645 ;
        RECT 41.430 147.675 41.760 148.475 ;
        RECT 42.060 147.845 42.390 148.645 ;
        RECT 42.560 147.675 42.890 148.475 ;
        RECT 40.455 147.505 42.890 147.675 ;
        RECT 43.265 147.555 44.475 148.645 ;
        RECT 44.650 148.210 49.995 148.645 ;
        RECT 38.205 146.865 39.415 147.385 ;
        RECT 35.440 146.645 36.105 146.815 ;
        RECT 35.435 146.095 35.765 146.475 ;
        RECT 35.935 146.355 36.105 146.645 ;
        RECT 36.825 146.095 39.415 146.865 ;
        RECT 39.585 146.895 39.760 147.505 ;
        RECT 40.455 147.255 40.625 147.505 ;
        RECT 39.930 147.085 40.625 147.255 ;
        RECT 40.800 147.085 41.220 147.285 ;
        RECT 41.390 147.085 41.720 147.285 ;
        RECT 41.890 147.085 42.220 147.285 ;
        RECT 39.585 146.265 39.925 146.895 ;
        RECT 40.095 146.095 40.345 146.895 ;
        RECT 40.535 146.745 41.760 146.915 ;
        RECT 40.535 146.265 40.865 146.745 ;
        RECT 41.035 146.095 41.260 146.555 ;
        RECT 41.430 146.265 41.760 146.745 ;
        RECT 42.390 146.875 42.560 147.505 ;
        RECT 42.745 147.085 43.095 147.335 ;
        RECT 43.265 147.015 43.785 147.555 ;
        RECT 42.390 146.265 42.890 146.875 ;
        RECT 43.955 146.845 44.475 147.385 ;
        RECT 46.240 146.960 46.590 148.210 ;
        RECT 50.165 147.480 50.455 148.645 ;
        RECT 51.085 147.505 51.355 148.475 ;
        RECT 51.565 147.845 51.845 148.645 ;
        RECT 52.015 148.135 53.670 148.425 ;
        RECT 52.080 147.795 53.670 147.965 ;
        RECT 52.080 147.675 52.250 147.795 ;
        RECT 51.525 147.505 52.250 147.675 ;
        RECT 43.265 146.095 44.475 146.845 ;
        RECT 48.070 146.640 48.410 147.470 ;
        RECT 44.650 146.095 49.995 146.640 ;
        RECT 50.165 146.095 50.455 146.820 ;
        RECT 51.085 146.770 51.255 147.505 ;
        RECT 51.525 147.335 51.695 147.505 ;
        RECT 52.440 147.455 53.155 147.625 ;
        RECT 53.350 147.505 53.670 147.795 ;
        RECT 53.845 147.505 54.185 148.475 ;
        RECT 54.355 147.505 54.525 148.645 ;
        RECT 54.795 147.845 55.045 148.645 ;
        RECT 55.690 147.675 56.020 148.475 ;
        RECT 56.320 147.845 56.650 148.645 ;
        RECT 56.820 147.675 57.150 148.475 ;
        RECT 54.715 147.505 57.150 147.675 ;
        RECT 57.525 147.505 57.865 148.475 ;
        RECT 58.035 147.505 58.205 148.645 ;
        RECT 58.475 147.845 58.725 148.645 ;
        RECT 59.370 147.675 59.700 148.475 ;
        RECT 60.000 147.845 60.330 148.645 ;
        RECT 60.500 147.675 60.830 148.475 ;
        RECT 58.395 147.505 60.830 147.675 ;
        RECT 61.265 147.505 61.475 148.645 ;
        RECT 51.425 147.005 51.695 147.335 ;
        RECT 51.865 147.005 52.270 147.335 ;
        RECT 52.440 147.005 53.150 147.455 ;
        RECT 51.525 146.835 51.695 147.005 ;
        RECT 51.085 146.425 51.355 146.770 ;
        RECT 51.525 146.665 53.135 146.835 ;
        RECT 53.320 146.765 53.670 147.335 ;
        RECT 53.845 146.895 54.020 147.505 ;
        RECT 54.715 147.255 54.885 147.505 ;
        RECT 54.190 147.085 54.885 147.255 ;
        RECT 55.060 147.085 55.480 147.285 ;
        RECT 55.650 147.085 55.980 147.285 ;
        RECT 56.150 147.085 56.480 147.285 ;
        RECT 51.545 146.095 51.925 146.495 ;
        RECT 52.095 146.315 52.265 146.665 ;
        RECT 52.435 146.095 52.765 146.495 ;
        RECT 52.965 146.315 53.135 146.665 ;
        RECT 53.335 146.095 53.665 146.595 ;
        RECT 53.845 146.265 54.185 146.895 ;
        RECT 54.355 146.095 54.605 146.895 ;
        RECT 54.795 146.745 56.020 146.915 ;
        RECT 54.795 146.265 55.125 146.745 ;
        RECT 55.295 146.095 55.520 146.555 ;
        RECT 55.690 146.265 56.020 146.745 ;
        RECT 56.650 146.875 56.820 147.505 ;
        RECT 57.005 147.085 57.355 147.335 ;
        RECT 57.525 146.945 57.700 147.505 ;
        RECT 58.395 147.255 58.565 147.505 ;
        RECT 57.870 147.085 58.565 147.255 ;
        RECT 58.740 147.085 59.160 147.285 ;
        RECT 59.330 147.085 59.660 147.285 ;
        RECT 59.830 147.085 60.160 147.285 ;
        RECT 57.525 146.895 57.755 146.945 ;
        RECT 56.650 146.265 57.150 146.875 ;
        RECT 57.525 146.265 57.865 146.895 ;
        RECT 58.035 146.095 58.285 146.895 ;
        RECT 58.475 146.745 59.700 146.915 ;
        RECT 58.475 146.265 58.805 146.745 ;
        RECT 58.975 146.095 59.200 146.555 ;
        RECT 59.370 146.265 59.700 146.745 ;
        RECT 60.330 146.875 60.500 147.505 ;
        RECT 61.645 147.495 61.975 148.475 ;
        RECT 62.145 147.505 62.375 148.645 ;
        RECT 62.585 147.555 65.175 148.645 ;
        RECT 60.685 147.085 61.035 147.335 ;
        RECT 60.330 146.265 60.830 146.875 ;
        RECT 61.265 146.095 61.475 146.915 ;
        RECT 61.645 146.895 61.895 147.495 ;
        RECT 62.065 147.085 62.395 147.335 ;
        RECT 62.585 147.035 63.795 147.555 ;
        RECT 65.350 147.455 65.605 148.335 ;
        RECT 65.775 147.505 66.080 148.645 ;
        RECT 66.420 148.265 66.750 148.645 ;
        RECT 66.930 148.095 67.100 148.385 ;
        RECT 67.270 148.185 67.520 148.645 ;
        RECT 66.300 147.925 67.100 148.095 ;
        RECT 67.690 148.135 68.560 148.475 ;
        RECT 61.645 146.265 61.975 146.895 ;
        RECT 62.145 146.095 62.375 146.915 ;
        RECT 63.965 146.865 65.175 147.385 ;
        RECT 62.585 146.095 65.175 146.865 ;
        RECT 65.350 146.805 65.560 147.455 ;
        RECT 66.300 147.335 66.470 147.925 ;
        RECT 67.690 147.755 67.860 148.135 ;
        RECT 68.795 148.015 68.965 148.475 ;
        RECT 69.135 148.185 69.505 148.645 ;
        RECT 69.800 148.045 69.970 148.385 ;
        RECT 70.140 148.215 70.470 148.645 ;
        RECT 70.705 148.045 70.875 148.385 ;
        RECT 66.640 147.585 67.860 147.755 ;
        RECT 68.030 147.675 68.490 147.965 ;
        RECT 68.795 147.845 69.355 148.015 ;
        RECT 69.800 147.875 70.875 148.045 ;
        RECT 71.045 148.145 71.725 148.475 ;
        RECT 71.940 148.145 72.190 148.475 ;
        RECT 72.360 148.185 72.610 148.645 ;
        RECT 69.185 147.705 69.355 147.845 ;
        RECT 68.030 147.665 68.995 147.675 ;
        RECT 67.690 147.495 67.860 147.585 ;
        RECT 68.320 147.505 68.995 147.665 ;
        RECT 65.730 147.305 66.470 147.335 ;
        RECT 65.730 147.005 66.645 147.305 ;
        RECT 66.320 146.830 66.645 147.005 ;
        RECT 65.350 146.275 65.605 146.805 ;
        RECT 65.775 146.095 66.080 146.555 ;
        RECT 66.325 146.475 66.645 146.830 ;
        RECT 66.815 147.045 67.355 147.415 ;
        RECT 67.690 147.325 68.095 147.495 ;
        RECT 66.815 146.645 67.055 147.045 ;
        RECT 67.535 146.875 67.755 147.155 ;
        RECT 67.225 146.705 67.755 146.875 ;
        RECT 67.225 146.475 67.395 146.705 ;
        RECT 67.925 146.545 68.095 147.325 ;
        RECT 68.265 146.715 68.615 147.335 ;
        RECT 68.785 146.715 68.995 147.505 ;
        RECT 69.185 147.535 70.685 147.705 ;
        RECT 69.185 146.845 69.355 147.535 ;
        RECT 71.045 147.365 71.215 148.145 ;
        RECT 72.020 148.015 72.190 148.145 ;
        RECT 69.525 147.195 71.215 147.365 ;
        RECT 71.385 147.585 71.850 147.975 ;
        RECT 72.020 147.845 72.415 148.015 ;
        RECT 69.525 147.015 69.695 147.195 ;
        RECT 66.325 146.305 67.395 146.475 ;
        RECT 67.565 146.095 67.755 146.535 ;
        RECT 67.925 146.265 68.875 146.545 ;
        RECT 69.185 146.455 69.445 146.845 ;
        RECT 69.865 146.775 70.655 147.025 ;
        RECT 69.095 146.285 69.445 146.455 ;
        RECT 69.655 146.095 69.985 146.555 ;
        RECT 70.860 146.485 71.030 147.195 ;
        RECT 71.385 146.995 71.555 147.585 ;
        RECT 71.200 146.775 71.555 146.995 ;
        RECT 71.725 146.775 72.075 147.395 ;
        RECT 72.245 146.485 72.415 147.845 ;
        RECT 72.780 147.675 73.105 148.460 ;
        RECT 72.585 146.625 73.045 147.675 ;
        RECT 70.860 146.315 71.715 146.485 ;
        RECT 71.920 146.315 72.415 146.485 ;
        RECT 72.585 146.095 72.915 146.455 ;
        RECT 73.275 146.355 73.445 148.475 ;
        RECT 73.615 148.145 73.945 148.645 ;
        RECT 74.115 147.975 74.370 148.475 ;
        RECT 73.620 147.805 74.370 147.975 ;
        RECT 73.620 146.815 73.850 147.805 ;
        RECT 74.020 146.985 74.370 147.635 ;
        RECT 74.545 147.555 75.755 148.645 ;
        RECT 74.545 147.015 75.065 147.555 ;
        RECT 75.925 147.480 76.215 148.645 ;
        RECT 76.385 147.555 77.595 148.645 ;
        RECT 77.765 147.555 81.275 148.645 ;
        RECT 81.450 148.135 83.105 148.425 ;
        RECT 81.450 147.795 83.040 147.965 ;
        RECT 83.275 147.845 83.555 148.645 ;
        RECT 75.235 146.845 75.755 147.385 ;
        RECT 76.385 147.015 76.905 147.555 ;
        RECT 77.075 146.845 77.595 147.385 ;
        RECT 77.765 147.035 79.455 147.555 ;
        RECT 81.450 147.505 81.770 147.795 ;
        RECT 82.870 147.675 83.040 147.795 ;
        RECT 79.625 146.865 81.275 147.385 ;
        RECT 73.620 146.645 74.370 146.815 ;
        RECT 73.615 146.095 73.945 146.475 ;
        RECT 74.115 146.355 74.370 146.645 ;
        RECT 74.545 146.095 75.755 146.845 ;
        RECT 75.925 146.095 76.215 146.820 ;
        RECT 76.385 146.095 77.595 146.845 ;
        RECT 77.765 146.095 81.275 146.865 ;
        RECT 81.450 146.765 81.800 147.335 ;
        RECT 81.970 147.005 82.680 147.625 ;
        RECT 82.870 147.505 83.595 147.675 ;
        RECT 83.765 147.505 84.035 148.475 ;
        RECT 85.130 148.210 90.475 148.645 ;
        RECT 90.650 148.210 95.995 148.645 ;
        RECT 96.170 148.210 101.515 148.645 ;
        RECT 83.425 147.335 83.595 147.505 ;
        RECT 82.850 147.005 83.255 147.335 ;
        RECT 83.425 147.005 83.695 147.335 ;
        RECT 83.425 146.835 83.595 147.005 ;
        RECT 81.985 146.665 83.595 146.835 ;
        RECT 83.865 146.770 84.035 147.505 ;
        RECT 86.720 146.960 87.070 148.210 ;
        RECT 81.455 146.095 81.785 146.595 ;
        RECT 81.985 146.315 82.155 146.665 ;
        RECT 82.355 146.095 82.685 146.495 ;
        RECT 82.855 146.315 83.025 146.665 ;
        RECT 83.195 146.095 83.575 146.495 ;
        RECT 83.765 146.425 84.035 146.770 ;
        RECT 88.550 146.640 88.890 147.470 ;
        RECT 92.240 146.960 92.590 148.210 ;
        RECT 94.070 146.640 94.410 147.470 ;
        RECT 97.760 146.960 98.110 148.210 ;
        RECT 101.685 147.480 101.975 148.645 ;
        RECT 102.145 147.555 105.655 148.645 ;
        RECT 99.590 146.640 99.930 147.470 ;
        RECT 102.145 147.035 103.835 147.555 ;
        RECT 105.825 147.505 106.095 148.475 ;
        RECT 106.305 147.845 106.585 148.645 ;
        RECT 106.755 148.135 108.410 148.425 ;
        RECT 106.820 147.795 108.410 147.965 ;
        RECT 106.820 147.675 106.990 147.795 ;
        RECT 106.265 147.505 106.990 147.675 ;
        RECT 104.005 146.865 105.655 147.385 ;
        RECT 85.130 146.095 90.475 146.640 ;
        RECT 90.650 146.095 95.995 146.640 ;
        RECT 96.170 146.095 101.515 146.640 ;
        RECT 101.685 146.095 101.975 146.820 ;
        RECT 102.145 146.095 105.655 146.865 ;
        RECT 105.825 146.770 105.995 147.505 ;
        RECT 106.265 147.335 106.435 147.505 ;
        RECT 106.165 147.005 106.435 147.335 ;
        RECT 106.605 147.005 107.010 147.335 ;
        RECT 107.180 147.005 107.890 147.625 ;
        RECT 108.090 147.505 108.410 147.795 ;
        RECT 108.585 147.505 108.855 148.475 ;
        RECT 109.065 147.845 109.345 148.645 ;
        RECT 109.515 148.135 111.170 148.425 ;
        RECT 109.580 147.795 111.170 147.965 ;
        RECT 109.580 147.675 109.750 147.795 ;
        RECT 109.025 147.505 109.750 147.675 ;
        RECT 106.265 146.835 106.435 147.005 ;
        RECT 105.825 146.425 106.095 146.770 ;
        RECT 106.265 146.665 107.875 146.835 ;
        RECT 108.060 146.765 108.410 147.335 ;
        RECT 108.585 146.770 108.755 147.505 ;
        RECT 109.025 147.335 109.195 147.505 ;
        RECT 109.940 147.455 110.655 147.625 ;
        RECT 110.850 147.505 111.170 147.795 ;
        RECT 111.345 147.505 111.685 148.475 ;
        RECT 111.855 147.505 112.025 148.645 ;
        RECT 112.295 147.845 112.545 148.645 ;
        RECT 113.190 147.675 113.520 148.475 ;
        RECT 113.820 147.845 114.150 148.645 ;
        RECT 114.320 147.675 114.650 148.475 ;
        RECT 112.215 147.505 114.650 147.675 ;
        RECT 115.025 147.555 116.235 148.645 ;
        RECT 116.405 147.555 119.915 148.645 ;
        RECT 108.925 147.005 109.195 147.335 ;
        RECT 109.365 147.005 109.770 147.335 ;
        RECT 109.940 147.005 110.650 147.455 ;
        RECT 109.025 146.835 109.195 147.005 ;
        RECT 106.285 146.095 106.665 146.495 ;
        RECT 106.835 146.315 107.005 146.665 ;
        RECT 107.175 146.095 107.505 146.495 ;
        RECT 107.705 146.315 107.875 146.665 ;
        RECT 108.075 146.095 108.405 146.595 ;
        RECT 108.585 146.425 108.855 146.770 ;
        RECT 109.025 146.665 110.635 146.835 ;
        RECT 110.820 146.765 111.170 147.335 ;
        RECT 111.345 146.945 111.520 147.505 ;
        RECT 112.215 147.255 112.385 147.505 ;
        RECT 111.690 147.085 112.385 147.255 ;
        RECT 112.560 147.085 112.980 147.285 ;
        RECT 113.150 147.085 113.480 147.285 ;
        RECT 113.650 147.085 113.980 147.285 ;
        RECT 111.345 146.895 111.575 146.945 ;
        RECT 109.045 146.095 109.425 146.495 ;
        RECT 109.595 146.315 109.765 146.665 ;
        RECT 109.935 146.095 110.265 146.495 ;
        RECT 110.465 146.315 110.635 146.665 ;
        RECT 110.835 146.095 111.165 146.595 ;
        RECT 111.345 146.265 111.685 146.895 ;
        RECT 111.855 146.095 112.105 146.895 ;
        RECT 112.295 146.745 113.520 146.915 ;
        RECT 112.295 146.265 112.625 146.745 ;
        RECT 112.795 146.095 113.020 146.555 ;
        RECT 113.190 146.265 113.520 146.745 ;
        RECT 114.150 146.875 114.320 147.505 ;
        RECT 114.505 147.085 114.855 147.335 ;
        RECT 115.025 147.015 115.545 147.555 ;
        RECT 114.150 146.265 114.650 146.875 ;
        RECT 115.715 146.845 116.235 147.385 ;
        RECT 116.405 147.035 118.095 147.555 ;
        RECT 120.125 147.505 120.355 148.645 ;
        RECT 120.525 147.495 120.855 148.475 ;
        RECT 121.025 147.505 121.235 148.645 ;
        RECT 121.465 147.555 122.675 148.645 ;
        RECT 122.845 147.555 126.355 148.645 ;
        RECT 126.525 147.555 127.735 148.645 ;
        RECT 118.265 146.865 119.915 147.385 ;
        RECT 120.105 147.085 120.435 147.335 ;
        RECT 115.025 146.095 116.235 146.845 ;
        RECT 116.405 146.095 119.915 146.865 ;
        RECT 120.125 146.095 120.355 146.915 ;
        RECT 120.605 146.895 120.855 147.495 ;
        RECT 121.465 147.015 121.985 147.555 ;
        RECT 120.525 146.265 120.855 146.895 ;
        RECT 121.025 146.095 121.235 146.915 ;
        RECT 122.155 146.845 122.675 147.385 ;
        RECT 122.845 147.035 124.535 147.555 ;
        RECT 124.705 146.865 126.355 147.385 ;
        RECT 126.525 147.015 127.045 147.555 ;
        RECT 121.465 146.095 122.675 146.845 ;
        RECT 122.845 146.095 126.355 146.865 ;
        RECT 127.215 146.845 127.735 147.385 ;
        RECT 126.525 146.095 127.735 146.845 ;
        RECT 20.640 145.925 127.820 146.095 ;
        RECT 20.725 145.175 21.935 145.925 ;
        RECT 20.725 144.635 21.245 145.175 ;
        RECT 22.565 145.155 24.235 145.925 ;
        RECT 24.410 145.380 29.755 145.925 ;
        RECT 21.415 144.465 21.935 145.005 ;
        RECT 20.725 143.375 21.935 144.465 ;
        RECT 22.565 144.465 23.315 144.985 ;
        RECT 23.485 144.635 24.235 145.155 ;
        RECT 22.565 143.375 24.235 144.465 ;
        RECT 26.000 143.810 26.350 145.060 ;
        RECT 27.830 144.550 28.170 145.380 ;
        RECT 29.965 145.105 30.195 145.925 ;
        RECT 30.365 145.125 30.695 145.755 ;
        RECT 29.945 144.685 30.275 144.935 ;
        RECT 30.445 144.525 30.695 145.125 ;
        RECT 30.865 145.105 31.075 145.925 ;
        RECT 31.770 145.380 37.115 145.925 ;
        RECT 24.410 143.375 29.755 143.810 ;
        RECT 29.965 143.375 30.195 144.515 ;
        RECT 30.365 143.545 30.695 144.525 ;
        RECT 30.865 143.375 31.075 144.515 ;
        RECT 33.360 143.810 33.710 145.060 ;
        RECT 35.190 144.550 35.530 145.380 ;
        RECT 37.285 145.200 37.575 145.925 ;
        RECT 37.745 145.155 39.415 145.925 ;
        RECT 31.770 143.375 37.115 143.810 ;
        RECT 37.285 143.375 37.575 144.540 ;
        RECT 37.745 144.465 38.495 144.985 ;
        RECT 38.665 144.635 39.415 145.155 ;
        RECT 39.585 145.250 39.855 145.595 ;
        RECT 40.045 145.525 40.425 145.925 ;
        RECT 40.595 145.355 40.765 145.705 ;
        RECT 40.935 145.525 41.265 145.925 ;
        RECT 41.465 145.355 41.635 145.705 ;
        RECT 41.835 145.425 42.165 145.925 ;
        RECT 39.585 144.515 39.755 145.250 ;
        RECT 40.025 145.185 41.635 145.355 ;
        RECT 40.025 145.015 40.195 145.185 ;
        RECT 39.925 144.685 40.195 145.015 ;
        RECT 40.365 144.685 40.770 145.015 ;
        RECT 40.025 144.515 40.195 144.685 ;
        RECT 40.940 144.565 41.650 145.015 ;
        RECT 41.820 144.685 42.170 145.255 ;
        RECT 42.345 145.250 42.615 145.595 ;
        RECT 42.805 145.525 43.185 145.925 ;
        RECT 43.355 145.355 43.525 145.705 ;
        RECT 43.695 145.525 44.025 145.925 ;
        RECT 44.225 145.355 44.395 145.705 ;
        RECT 44.595 145.425 44.925 145.925 ;
        RECT 37.745 143.375 39.415 144.465 ;
        RECT 39.585 143.545 39.855 144.515 ;
        RECT 40.025 144.345 40.750 144.515 ;
        RECT 40.940 144.395 41.655 144.565 ;
        RECT 42.345 144.515 42.515 145.250 ;
        RECT 42.785 145.185 44.395 145.355 ;
        RECT 42.785 145.015 42.955 145.185 ;
        RECT 42.685 144.685 42.955 145.015 ;
        RECT 43.125 144.685 43.530 145.015 ;
        RECT 42.785 144.515 42.955 144.685 ;
        RECT 40.580 144.225 40.750 144.345 ;
        RECT 41.850 144.225 42.170 144.515 ;
        RECT 40.065 143.375 40.345 144.175 ;
        RECT 40.580 144.055 42.170 144.225 ;
        RECT 40.515 143.595 42.170 143.885 ;
        RECT 42.345 143.545 42.615 144.515 ;
        RECT 42.785 144.345 43.510 144.515 ;
        RECT 43.700 144.395 44.410 145.015 ;
        RECT 44.580 144.685 44.930 145.255 ;
        RECT 45.105 145.250 45.375 145.595 ;
        RECT 45.565 145.525 45.945 145.925 ;
        RECT 46.115 145.355 46.285 145.705 ;
        RECT 46.455 145.525 46.785 145.925 ;
        RECT 46.985 145.355 47.155 145.705 ;
        RECT 47.355 145.425 47.685 145.925 ;
        RECT 45.105 144.515 45.275 145.250 ;
        RECT 45.545 145.185 47.155 145.355 ;
        RECT 45.545 145.015 45.715 145.185 ;
        RECT 45.445 144.685 45.715 145.015 ;
        RECT 45.885 144.685 46.290 145.015 ;
        RECT 45.545 144.515 45.715 144.685 ;
        RECT 43.340 144.225 43.510 144.345 ;
        RECT 44.610 144.225 44.930 144.515 ;
        RECT 42.825 143.375 43.105 144.175 ;
        RECT 43.340 144.055 44.930 144.225 ;
        RECT 43.275 143.595 44.930 143.885 ;
        RECT 45.105 143.545 45.375 144.515 ;
        RECT 45.545 144.345 46.270 144.515 ;
        RECT 46.460 144.395 47.170 145.015 ;
        RECT 47.340 144.685 47.690 145.255 ;
        RECT 47.865 145.250 48.135 145.595 ;
        RECT 48.325 145.525 48.705 145.925 ;
        RECT 48.875 145.355 49.045 145.705 ;
        RECT 49.215 145.525 49.545 145.925 ;
        RECT 49.745 145.355 49.915 145.705 ;
        RECT 50.115 145.425 50.445 145.925 ;
        RECT 47.865 144.515 48.035 145.250 ;
        RECT 48.305 145.185 49.915 145.355 ;
        RECT 48.305 145.015 48.475 145.185 ;
        RECT 48.205 144.685 48.475 145.015 ;
        RECT 48.645 144.685 49.050 145.015 ;
        RECT 48.305 144.515 48.475 144.685 ;
        RECT 49.220 144.565 49.930 145.015 ;
        RECT 50.100 144.685 50.450 145.255 ;
        RECT 50.625 145.125 50.965 145.755 ;
        RECT 51.135 145.125 51.385 145.925 ;
        RECT 51.575 145.275 51.905 145.755 ;
        RECT 52.075 145.465 52.300 145.925 ;
        RECT 52.470 145.275 52.800 145.755 ;
        RECT 46.100 144.225 46.270 144.345 ;
        RECT 47.370 144.225 47.690 144.515 ;
        RECT 45.585 143.375 45.865 144.175 ;
        RECT 46.100 144.055 47.690 144.225 ;
        RECT 46.035 143.595 47.690 143.885 ;
        RECT 47.865 143.545 48.135 144.515 ;
        RECT 48.305 144.345 49.030 144.515 ;
        RECT 49.220 144.395 49.935 144.565 ;
        RECT 50.625 144.515 50.800 145.125 ;
        RECT 51.575 145.105 52.800 145.275 ;
        RECT 53.430 145.145 53.930 145.755 ;
        RECT 50.970 144.765 51.665 144.935 ;
        RECT 51.495 144.515 51.665 144.765 ;
        RECT 51.840 144.735 52.260 144.935 ;
        RECT 52.430 144.735 52.760 144.935 ;
        RECT 52.930 144.735 53.260 144.935 ;
        RECT 53.430 144.515 53.600 145.145 ;
        RECT 54.305 145.125 54.645 145.755 ;
        RECT 54.815 145.125 55.065 145.925 ;
        RECT 55.255 145.275 55.585 145.755 ;
        RECT 55.755 145.465 55.980 145.925 ;
        RECT 56.150 145.275 56.480 145.755 ;
        RECT 53.785 144.685 54.135 144.935 ;
        RECT 54.305 144.515 54.480 145.125 ;
        RECT 55.255 145.105 56.480 145.275 ;
        RECT 57.110 145.145 57.610 145.755 ;
        RECT 54.650 144.765 55.345 144.935 ;
        RECT 55.175 144.515 55.345 144.765 ;
        RECT 55.520 144.735 55.940 144.935 ;
        RECT 56.110 144.735 56.440 144.935 ;
        RECT 56.610 144.735 56.940 144.935 ;
        RECT 57.110 144.515 57.280 145.145 ;
        RECT 59.180 145.115 59.425 145.720 ;
        RECT 59.645 145.390 60.155 145.925 ;
        RECT 58.905 144.945 60.135 145.115 ;
        RECT 57.465 144.685 57.815 144.935 ;
        RECT 48.860 144.225 49.030 144.345 ;
        RECT 50.130 144.225 50.450 144.515 ;
        RECT 48.345 143.375 48.625 144.175 ;
        RECT 48.860 144.055 50.450 144.225 ;
        RECT 48.795 143.595 50.450 143.885 ;
        RECT 50.625 143.545 50.965 144.515 ;
        RECT 51.135 143.375 51.305 144.515 ;
        RECT 51.495 144.345 53.930 144.515 ;
        RECT 51.575 143.375 51.825 144.175 ;
        RECT 52.470 143.545 52.800 144.345 ;
        RECT 53.100 143.375 53.430 144.175 ;
        RECT 53.600 143.545 53.930 144.345 ;
        RECT 54.305 143.545 54.645 144.515 ;
        RECT 54.815 143.375 54.985 144.515 ;
        RECT 55.175 144.345 57.610 144.515 ;
        RECT 55.255 143.375 55.505 144.175 ;
        RECT 56.150 143.545 56.480 144.345 ;
        RECT 56.780 143.375 57.110 144.175 ;
        RECT 57.280 143.545 57.610 144.345 ;
        RECT 58.905 144.135 59.245 144.945 ;
        RECT 59.415 144.380 60.165 144.570 ;
        RECT 58.905 143.725 59.420 144.135 ;
        RECT 59.655 143.375 59.825 144.135 ;
        RECT 59.995 143.715 60.165 144.380 ;
        RECT 60.335 144.395 60.525 145.755 ;
        RECT 60.695 145.585 60.970 145.755 ;
        RECT 60.695 145.415 60.975 145.585 ;
        RECT 60.695 144.595 60.970 145.415 ;
        RECT 61.160 145.390 61.690 145.755 ;
        RECT 62.115 145.525 62.445 145.925 ;
        RECT 61.515 145.355 61.690 145.390 ;
        RECT 61.175 144.395 61.345 145.195 ;
        RECT 60.335 144.225 61.345 144.395 ;
        RECT 61.515 145.185 62.445 145.355 ;
        RECT 62.615 145.185 62.870 145.755 ;
        RECT 63.045 145.200 63.335 145.925 ;
        RECT 61.515 144.055 61.685 145.185 ;
        RECT 62.275 145.015 62.445 145.185 ;
        RECT 60.560 143.885 61.685 144.055 ;
        RECT 61.855 144.685 62.050 145.015 ;
        RECT 62.275 144.685 62.530 145.015 ;
        RECT 61.855 143.715 62.025 144.685 ;
        RECT 62.700 144.515 62.870 145.185 ;
        RECT 64.425 145.125 64.765 145.755 ;
        RECT 64.935 145.125 65.185 145.925 ;
        RECT 65.375 145.275 65.705 145.755 ;
        RECT 65.875 145.465 66.100 145.925 ;
        RECT 66.270 145.275 66.600 145.755 ;
        RECT 59.995 143.545 62.025 143.715 ;
        RECT 62.195 143.375 62.365 144.515 ;
        RECT 62.535 143.545 62.870 144.515 ;
        RECT 63.045 143.375 63.335 144.540 ;
        RECT 64.425 144.515 64.600 145.125 ;
        RECT 65.375 145.105 66.600 145.275 ;
        RECT 67.230 145.145 67.730 145.755 ;
        RECT 64.770 144.765 65.465 144.935 ;
        RECT 65.295 144.515 65.465 144.765 ;
        RECT 65.640 144.735 66.060 144.935 ;
        RECT 66.230 144.735 66.560 144.935 ;
        RECT 66.730 144.735 67.060 144.935 ;
        RECT 67.230 144.515 67.400 145.145 ;
        RECT 68.380 145.115 68.625 145.720 ;
        RECT 68.845 145.390 69.355 145.925 ;
        RECT 68.105 144.945 69.335 145.115 ;
        RECT 67.585 144.685 67.935 144.935 ;
        RECT 64.425 143.545 64.765 144.515 ;
        RECT 64.935 143.375 65.105 144.515 ;
        RECT 65.295 144.345 67.730 144.515 ;
        RECT 65.375 143.375 65.625 144.175 ;
        RECT 66.270 143.545 66.600 144.345 ;
        RECT 66.900 143.375 67.230 144.175 ;
        RECT 67.400 143.545 67.730 144.345 ;
        RECT 68.105 144.135 68.445 144.945 ;
        RECT 68.615 144.380 69.365 144.570 ;
        RECT 68.105 143.725 68.620 144.135 ;
        RECT 68.855 143.375 69.025 144.135 ;
        RECT 69.195 143.715 69.365 144.380 ;
        RECT 69.535 144.395 69.725 145.755 ;
        RECT 69.895 144.905 70.170 145.755 ;
        RECT 70.360 145.390 70.890 145.755 ;
        RECT 71.315 145.525 71.645 145.925 ;
        RECT 70.715 145.355 70.890 145.390 ;
        RECT 69.895 144.735 70.175 144.905 ;
        RECT 69.895 144.595 70.170 144.735 ;
        RECT 70.375 144.395 70.545 145.195 ;
        RECT 69.535 144.225 70.545 144.395 ;
        RECT 70.715 145.185 71.645 145.355 ;
        RECT 71.815 145.185 72.070 145.755 ;
        RECT 70.715 144.055 70.885 145.185 ;
        RECT 71.475 145.015 71.645 145.185 ;
        RECT 69.760 143.885 70.885 144.055 ;
        RECT 71.055 144.685 71.250 145.015 ;
        RECT 71.475 144.685 71.730 145.015 ;
        RECT 71.055 143.715 71.225 144.685 ;
        RECT 71.900 144.515 72.070 145.185 ;
        RECT 72.305 145.105 72.515 145.925 ;
        RECT 72.685 145.125 73.015 145.755 ;
        RECT 72.685 144.525 72.935 145.125 ;
        RECT 73.185 145.105 73.415 145.925 ;
        RECT 73.625 145.175 74.835 145.925 ;
        RECT 73.105 144.685 73.435 144.935 ;
        RECT 69.195 143.545 71.225 143.715 ;
        RECT 71.395 143.375 71.565 144.515 ;
        RECT 71.735 143.545 72.070 144.515 ;
        RECT 72.305 143.375 72.515 144.515 ;
        RECT 72.685 143.545 73.015 144.525 ;
        RECT 73.185 143.375 73.415 144.515 ;
        RECT 73.625 144.465 74.145 145.005 ;
        RECT 74.315 144.635 74.835 145.175 ;
        RECT 75.005 145.155 78.515 145.925 ;
        RECT 75.005 144.465 76.695 144.985 ;
        RECT 76.865 144.635 78.515 145.155 ;
        RECT 78.890 145.145 79.390 145.755 ;
        RECT 78.685 144.685 79.035 144.935 ;
        RECT 79.220 144.515 79.390 145.145 ;
        RECT 80.020 145.275 80.350 145.755 ;
        RECT 80.520 145.465 80.745 145.925 ;
        RECT 80.915 145.275 81.245 145.755 ;
        RECT 80.020 145.105 81.245 145.275 ;
        RECT 81.435 145.125 81.685 145.925 ;
        RECT 81.855 145.125 82.195 145.755 ;
        RECT 79.560 144.735 79.890 144.935 ;
        RECT 80.060 144.735 80.390 144.935 ;
        RECT 80.560 144.735 80.980 144.935 ;
        RECT 81.155 144.765 81.850 144.935 ;
        RECT 81.155 144.515 81.325 144.765 ;
        RECT 82.020 144.515 82.195 145.125 ;
        RECT 73.625 143.375 74.835 144.465 ;
        RECT 75.005 143.375 78.515 144.465 ;
        RECT 78.890 144.345 81.325 144.515 ;
        RECT 78.890 143.545 79.220 144.345 ;
        RECT 79.390 143.375 79.720 144.175 ;
        RECT 80.020 143.545 80.350 144.345 ;
        RECT 80.995 143.375 81.245 144.175 ;
        RECT 81.515 143.375 81.685 144.515 ;
        RECT 81.855 143.545 82.195 144.515 ;
        RECT 82.365 145.125 82.705 145.755 ;
        RECT 82.875 145.125 83.125 145.925 ;
        RECT 83.315 145.275 83.645 145.755 ;
        RECT 83.815 145.465 84.040 145.925 ;
        RECT 84.210 145.275 84.540 145.755 ;
        RECT 82.365 144.515 82.540 145.125 ;
        RECT 83.315 145.105 84.540 145.275 ;
        RECT 85.170 145.145 85.670 145.755 ;
        RECT 86.045 145.155 88.635 145.925 ;
        RECT 88.805 145.200 89.095 145.925 ;
        RECT 90.185 145.155 93.695 145.925 ;
        RECT 93.870 145.380 99.215 145.925 ;
        RECT 99.390 145.380 104.735 145.925 ;
        RECT 104.910 145.380 110.255 145.925 ;
        RECT 110.435 145.425 110.765 145.925 ;
        RECT 82.710 144.765 83.405 144.935 ;
        RECT 83.235 144.515 83.405 144.765 ;
        RECT 83.580 144.735 84.000 144.935 ;
        RECT 84.170 144.735 84.500 144.935 ;
        RECT 84.670 144.735 85.000 144.935 ;
        RECT 85.170 144.515 85.340 145.145 ;
        RECT 85.525 144.685 85.875 144.935 ;
        RECT 82.365 143.545 82.705 144.515 ;
        RECT 82.875 143.375 83.045 144.515 ;
        RECT 83.235 144.345 85.670 144.515 ;
        RECT 83.315 143.375 83.565 144.175 ;
        RECT 84.210 143.545 84.540 144.345 ;
        RECT 84.840 143.375 85.170 144.175 ;
        RECT 85.340 143.545 85.670 144.345 ;
        RECT 86.045 144.465 87.255 144.985 ;
        RECT 87.425 144.635 88.635 145.155 ;
        RECT 86.045 143.375 88.635 144.465 ;
        RECT 88.805 143.375 89.095 144.540 ;
        RECT 90.185 144.465 91.875 144.985 ;
        RECT 92.045 144.635 93.695 145.155 ;
        RECT 90.185 143.375 93.695 144.465 ;
        RECT 95.460 143.810 95.810 145.060 ;
        RECT 97.290 144.550 97.630 145.380 ;
        RECT 100.980 143.810 101.330 145.060 ;
        RECT 102.810 144.550 103.150 145.380 ;
        RECT 106.500 143.810 106.850 145.060 ;
        RECT 108.330 144.550 108.670 145.380 ;
        RECT 110.965 145.355 111.135 145.705 ;
        RECT 111.335 145.525 111.665 145.925 ;
        RECT 111.835 145.355 112.005 145.705 ;
        RECT 112.175 145.525 112.555 145.925 ;
        RECT 110.430 144.685 110.780 145.255 ;
        RECT 110.965 145.185 112.575 145.355 ;
        RECT 112.745 145.250 113.015 145.595 ;
        RECT 112.405 145.015 112.575 145.185 ;
        RECT 110.430 144.225 110.750 144.515 ;
        RECT 110.950 144.395 111.660 145.015 ;
        RECT 111.830 144.685 112.235 145.015 ;
        RECT 112.405 144.685 112.675 145.015 ;
        RECT 112.405 144.515 112.575 144.685 ;
        RECT 112.845 144.515 113.015 145.250 ;
        RECT 113.185 145.175 114.395 145.925 ;
        RECT 114.565 145.200 114.855 145.925 ;
        RECT 111.850 144.345 112.575 144.515 ;
        RECT 111.850 144.225 112.020 144.345 ;
        RECT 110.430 144.055 112.020 144.225 ;
        RECT 93.870 143.375 99.215 143.810 ;
        RECT 99.390 143.375 104.735 143.810 ;
        RECT 104.910 143.375 110.255 143.810 ;
        RECT 110.430 143.595 112.085 143.885 ;
        RECT 112.255 143.375 112.535 144.175 ;
        RECT 112.745 143.545 113.015 144.515 ;
        RECT 113.185 144.465 113.705 145.005 ;
        RECT 113.875 144.635 114.395 145.175 ;
        RECT 115.025 145.155 117.615 145.925 ;
        RECT 113.185 143.375 114.395 144.465 ;
        RECT 114.565 143.375 114.855 144.540 ;
        RECT 115.025 144.465 116.235 144.985 ;
        RECT 116.405 144.635 117.615 145.155 ;
        RECT 117.825 145.105 118.055 145.925 ;
        RECT 118.225 145.125 118.555 145.755 ;
        RECT 117.805 144.685 118.135 144.935 ;
        RECT 118.305 144.525 118.555 145.125 ;
        RECT 118.725 145.105 118.935 145.925 ;
        RECT 119.665 145.105 119.895 145.925 ;
        RECT 120.065 145.125 120.395 145.755 ;
        RECT 119.645 144.685 119.975 144.935 ;
        RECT 120.145 144.525 120.395 145.125 ;
        RECT 120.565 145.105 120.775 145.925 ;
        RECT 121.010 145.380 126.355 145.925 ;
        RECT 115.025 143.375 117.615 144.465 ;
        RECT 117.825 143.375 118.055 144.515 ;
        RECT 118.225 143.545 118.555 144.525 ;
        RECT 118.725 143.375 118.935 144.515 ;
        RECT 119.665 143.375 119.895 144.515 ;
        RECT 120.065 143.545 120.395 144.525 ;
        RECT 120.565 143.375 120.775 144.515 ;
        RECT 122.600 143.810 122.950 145.060 ;
        RECT 124.430 144.550 124.770 145.380 ;
        RECT 126.525 145.175 127.735 145.925 ;
        RECT 126.525 144.465 127.045 145.005 ;
        RECT 127.215 144.635 127.735 145.175 ;
        RECT 121.010 143.375 126.355 143.810 ;
        RECT 126.525 143.375 127.735 144.465 ;
        RECT 20.640 143.205 127.820 143.375 ;
        RECT 20.725 142.115 21.935 143.205 ;
        RECT 20.725 141.405 21.245 141.945 ;
        RECT 21.415 141.575 21.935 142.115 ;
        RECT 22.565 142.115 24.235 143.205 ;
        RECT 22.565 141.595 23.315 142.115 ;
        RECT 24.405 142.040 24.695 143.205 ;
        RECT 25.330 142.770 30.675 143.205 ;
        RECT 30.850 142.770 36.195 143.205 ;
        RECT 36.370 142.770 41.715 143.205 ;
        RECT 23.485 141.425 24.235 141.945 ;
        RECT 26.920 141.520 27.270 142.770 ;
        RECT 20.725 140.655 21.935 141.405 ;
        RECT 22.565 140.655 24.235 141.425 ;
        RECT 24.405 140.655 24.695 141.380 ;
        RECT 28.750 141.200 29.090 142.030 ;
        RECT 32.440 141.520 32.790 142.770 ;
        RECT 34.270 141.200 34.610 142.030 ;
        RECT 37.960 141.520 38.310 142.770 ;
        RECT 41.885 142.065 42.155 143.035 ;
        RECT 42.365 142.405 42.645 143.205 ;
        RECT 42.815 142.695 44.470 142.985 ;
        RECT 44.845 142.535 45.125 143.205 ;
        RECT 42.880 142.355 44.470 142.525 ;
        RECT 42.880 142.235 43.050 142.355 ;
        RECT 42.325 142.065 43.050 142.235 ;
        RECT 39.790 141.200 40.130 142.030 ;
        RECT 41.885 141.330 42.055 142.065 ;
        RECT 42.325 141.895 42.495 142.065 ;
        RECT 42.225 141.565 42.495 141.895 ;
        RECT 42.665 141.565 43.070 141.895 ;
        RECT 43.240 141.565 43.950 142.185 ;
        RECT 44.150 142.065 44.470 142.355 ;
        RECT 45.295 142.315 45.595 142.865 ;
        RECT 45.795 142.485 46.125 143.205 ;
        RECT 46.315 142.485 46.775 143.035 ;
        RECT 44.660 141.895 44.925 142.255 ;
        RECT 45.295 142.145 46.235 142.315 ;
        RECT 46.065 141.895 46.235 142.145 ;
        RECT 42.325 141.395 42.495 141.565 ;
        RECT 25.330 140.655 30.675 141.200 ;
        RECT 30.850 140.655 36.195 141.200 ;
        RECT 36.370 140.655 41.715 141.200 ;
        RECT 41.885 140.985 42.155 141.330 ;
        RECT 42.325 141.225 43.935 141.395 ;
        RECT 44.120 141.325 44.470 141.895 ;
        RECT 44.660 141.645 45.335 141.895 ;
        RECT 45.555 141.645 45.895 141.895 ;
        RECT 46.065 141.565 46.355 141.895 ;
        RECT 46.065 141.475 46.235 141.565 ;
        RECT 42.345 140.655 42.725 141.055 ;
        RECT 42.895 140.875 43.065 141.225 ;
        RECT 43.235 140.655 43.565 141.055 ;
        RECT 43.765 140.875 43.935 141.225 ;
        RECT 44.845 141.285 46.235 141.475 ;
        RECT 44.135 140.655 44.465 141.155 ;
        RECT 44.845 140.925 45.175 141.285 ;
        RECT 46.525 141.115 46.775 142.485 ;
        RECT 47.405 142.115 49.995 143.205 ;
        RECT 47.405 141.595 48.615 142.115 ;
        RECT 50.165 142.040 50.455 143.205 ;
        RECT 50.630 142.770 55.975 143.205 ;
        RECT 48.785 141.425 49.995 141.945 ;
        RECT 52.220 141.520 52.570 142.770 ;
        RECT 56.520 142.225 56.775 142.895 ;
        RECT 56.955 142.405 57.240 143.205 ;
        RECT 57.420 142.485 57.750 142.995 ;
        RECT 45.795 140.655 46.045 141.115 ;
        RECT 46.215 140.825 46.775 141.115 ;
        RECT 47.405 140.655 49.995 141.425 ;
        RECT 50.165 140.655 50.455 141.380 ;
        RECT 54.050 141.200 54.390 142.030 ;
        RECT 56.520 141.365 56.700 142.225 ;
        RECT 57.420 141.895 57.670 142.485 ;
        RECT 58.020 142.335 58.190 142.945 ;
        RECT 58.360 142.515 58.690 143.205 ;
        RECT 58.920 142.655 59.160 142.945 ;
        RECT 59.360 142.825 59.780 143.205 ;
        RECT 59.960 142.735 60.590 142.985 ;
        RECT 61.060 142.825 61.390 143.205 ;
        RECT 59.960 142.655 60.130 142.735 ;
        RECT 61.560 142.655 61.730 142.945 ;
        RECT 61.910 142.825 62.290 143.205 ;
        RECT 62.530 142.820 63.360 142.990 ;
        RECT 58.920 142.485 60.130 142.655 ;
        RECT 56.870 141.565 57.670 141.895 ;
        RECT 50.630 140.655 55.975 141.200 ;
        RECT 56.520 141.165 56.775 141.365 ;
        RECT 56.435 140.995 56.775 141.165 ;
        RECT 56.520 140.835 56.775 140.995 ;
        RECT 56.955 140.655 57.240 141.115 ;
        RECT 57.420 140.915 57.670 141.565 ;
        RECT 57.870 142.315 58.190 142.335 ;
        RECT 57.870 142.145 59.790 142.315 ;
        RECT 57.870 141.250 58.060 142.145 ;
        RECT 59.960 141.975 60.130 142.485 ;
        RECT 60.300 142.225 60.820 142.535 ;
        RECT 58.230 141.805 60.130 141.975 ;
        RECT 58.230 141.745 58.560 141.805 ;
        RECT 58.710 141.575 59.040 141.635 ;
        RECT 58.380 141.305 59.040 141.575 ;
        RECT 57.870 140.920 58.190 141.250 ;
        RECT 58.370 140.655 59.030 141.135 ;
        RECT 59.230 141.045 59.400 141.805 ;
        RECT 60.300 141.635 60.480 142.045 ;
        RECT 59.570 141.465 59.900 141.585 ;
        RECT 60.650 141.465 60.820 142.225 ;
        RECT 59.570 141.295 60.820 141.465 ;
        RECT 60.990 142.405 62.360 142.655 ;
        RECT 60.990 141.635 61.180 142.405 ;
        RECT 62.110 142.145 62.360 142.405 ;
        RECT 61.350 141.975 61.600 142.135 ;
        RECT 62.530 141.975 62.700 142.820 ;
        RECT 63.595 142.535 63.765 143.035 ;
        RECT 63.935 142.705 64.265 143.205 ;
        RECT 62.870 142.145 63.370 142.525 ;
        RECT 63.595 142.365 64.290 142.535 ;
        RECT 61.350 141.805 62.700 141.975 ;
        RECT 62.280 141.765 62.700 141.805 ;
        RECT 60.990 141.295 61.410 141.635 ;
        RECT 61.700 141.305 62.110 141.635 ;
        RECT 59.230 140.875 60.080 141.045 ;
        RECT 60.640 140.655 60.960 141.115 ;
        RECT 61.160 140.865 61.410 141.295 ;
        RECT 61.700 140.655 62.110 141.095 ;
        RECT 62.280 141.035 62.450 141.765 ;
        RECT 62.620 141.215 62.970 141.585 ;
        RECT 63.150 141.275 63.370 142.145 ;
        RECT 63.540 141.575 63.950 142.195 ;
        RECT 64.120 141.395 64.290 142.365 ;
        RECT 63.595 141.205 64.290 141.395 ;
        RECT 62.280 140.835 63.295 141.035 ;
        RECT 63.595 140.875 63.765 141.205 ;
        RECT 63.935 140.655 64.265 141.035 ;
        RECT 64.480 140.915 64.705 143.035 ;
        RECT 64.875 142.705 65.205 143.205 ;
        RECT 65.375 142.535 65.545 143.035 ;
        RECT 64.880 142.365 65.545 142.535 ;
        RECT 64.880 141.375 65.110 142.365 ;
        RECT 66.640 142.225 66.895 142.895 ;
        RECT 67.075 142.405 67.360 143.205 ;
        RECT 67.540 142.485 67.870 142.995 ;
        RECT 65.280 141.545 65.630 142.195 ;
        RECT 66.640 142.185 66.820 142.225 ;
        RECT 66.555 142.015 66.820 142.185 ;
        RECT 64.880 141.205 65.545 141.375 ;
        RECT 64.875 140.655 65.205 141.035 ;
        RECT 65.375 140.915 65.545 141.205 ;
        RECT 66.640 141.365 66.820 142.015 ;
        RECT 67.540 141.895 67.790 142.485 ;
        RECT 68.140 142.335 68.310 142.945 ;
        RECT 68.480 142.515 68.810 143.205 ;
        RECT 69.040 142.655 69.280 142.945 ;
        RECT 69.480 142.825 69.900 143.205 ;
        RECT 70.080 142.735 70.710 142.985 ;
        RECT 71.180 142.825 71.510 143.205 ;
        RECT 70.080 142.655 70.250 142.735 ;
        RECT 71.680 142.655 71.850 142.945 ;
        RECT 72.030 142.825 72.410 143.205 ;
        RECT 72.650 142.820 73.480 142.990 ;
        RECT 69.040 142.485 70.250 142.655 ;
        RECT 66.990 141.565 67.790 141.895 ;
        RECT 66.640 140.835 66.895 141.365 ;
        RECT 67.075 140.655 67.360 141.115 ;
        RECT 67.540 140.915 67.790 141.565 ;
        RECT 67.990 142.315 68.310 142.335 ;
        RECT 67.990 142.145 69.910 142.315 ;
        RECT 67.990 141.250 68.180 142.145 ;
        RECT 70.080 141.975 70.250 142.485 ;
        RECT 70.420 142.225 70.940 142.535 ;
        RECT 68.350 141.805 70.250 141.975 ;
        RECT 68.350 141.745 68.680 141.805 ;
        RECT 68.830 141.575 69.160 141.635 ;
        RECT 68.500 141.305 69.160 141.575 ;
        RECT 67.990 140.920 68.310 141.250 ;
        RECT 68.490 140.655 69.150 141.135 ;
        RECT 69.350 141.045 69.520 141.805 ;
        RECT 70.420 141.635 70.600 142.045 ;
        RECT 69.690 141.465 70.020 141.585 ;
        RECT 70.770 141.465 70.940 142.225 ;
        RECT 69.690 141.295 70.940 141.465 ;
        RECT 71.110 142.405 72.480 142.655 ;
        RECT 71.110 141.635 71.300 142.405 ;
        RECT 72.230 142.145 72.480 142.405 ;
        RECT 71.470 141.975 71.720 142.135 ;
        RECT 72.650 141.975 72.820 142.820 ;
        RECT 73.715 142.535 73.885 143.035 ;
        RECT 74.055 142.705 74.385 143.205 ;
        RECT 72.990 142.145 73.490 142.525 ;
        RECT 73.715 142.365 74.410 142.535 ;
        RECT 71.470 141.805 72.820 141.975 ;
        RECT 72.400 141.765 72.820 141.805 ;
        RECT 71.110 141.295 71.530 141.635 ;
        RECT 71.820 141.305 72.230 141.635 ;
        RECT 69.350 140.875 70.200 141.045 ;
        RECT 70.760 140.655 71.080 141.115 ;
        RECT 71.280 140.865 71.530 141.295 ;
        RECT 71.820 140.655 72.230 141.095 ;
        RECT 72.400 141.035 72.570 141.765 ;
        RECT 72.740 141.215 73.090 141.585 ;
        RECT 73.270 141.275 73.490 142.145 ;
        RECT 73.660 141.575 74.070 142.195 ;
        RECT 74.240 141.395 74.410 142.365 ;
        RECT 73.715 141.205 74.410 141.395 ;
        RECT 72.400 140.835 73.415 141.035 ;
        RECT 73.715 140.875 73.885 141.205 ;
        RECT 74.055 140.655 74.385 141.035 ;
        RECT 74.600 140.915 74.825 143.035 ;
        RECT 74.995 142.705 75.325 143.205 ;
        RECT 75.495 142.535 75.665 143.035 ;
        RECT 75.000 142.365 75.665 142.535 ;
        RECT 75.000 141.375 75.230 142.365 ;
        RECT 75.400 141.545 75.750 142.195 ;
        RECT 75.925 142.040 76.215 143.205 ;
        RECT 76.845 142.115 79.435 143.205 ;
        RECT 76.845 141.595 78.055 142.115 ;
        RECT 79.605 142.065 79.875 143.035 ;
        RECT 80.085 142.405 80.365 143.205 ;
        RECT 80.535 142.695 82.190 142.985 ;
        RECT 80.600 142.355 82.190 142.525 ;
        RECT 80.600 142.235 80.770 142.355 ;
        RECT 80.045 142.065 80.770 142.235 ;
        RECT 78.225 141.425 79.435 141.945 ;
        RECT 75.000 141.205 75.665 141.375 ;
        RECT 74.995 140.655 75.325 141.035 ;
        RECT 75.495 140.915 75.665 141.205 ;
        RECT 75.925 140.655 76.215 141.380 ;
        RECT 76.845 140.655 79.435 141.425 ;
        RECT 79.605 141.330 79.775 142.065 ;
        RECT 80.045 141.895 80.215 142.065 ;
        RECT 80.960 142.015 81.675 142.185 ;
        RECT 81.870 142.065 82.190 142.355 ;
        RECT 82.365 142.445 82.880 142.855 ;
        RECT 83.115 142.445 83.285 143.205 ;
        RECT 83.455 142.865 85.485 143.035 ;
        RECT 79.945 141.565 80.215 141.895 ;
        RECT 80.385 141.565 80.790 141.895 ;
        RECT 80.960 141.565 81.670 142.015 ;
        RECT 80.045 141.395 80.215 141.565 ;
        RECT 79.605 140.985 79.875 141.330 ;
        RECT 80.045 141.225 81.655 141.395 ;
        RECT 81.840 141.325 82.190 141.895 ;
        RECT 82.365 141.635 82.705 142.445 ;
        RECT 83.455 142.200 83.625 142.865 ;
        RECT 84.020 142.525 85.145 142.695 ;
        RECT 82.875 142.010 83.625 142.200 ;
        RECT 83.795 142.185 84.805 142.355 ;
        RECT 82.365 141.465 83.595 141.635 ;
        RECT 80.065 140.655 80.445 141.055 ;
        RECT 80.615 140.875 80.785 141.225 ;
        RECT 80.955 140.655 81.285 141.055 ;
        RECT 81.485 140.875 81.655 141.225 ;
        RECT 81.855 140.655 82.185 141.155 ;
        RECT 82.640 140.860 82.885 141.465 ;
        RECT 83.105 140.655 83.615 141.190 ;
        RECT 83.795 140.825 83.985 142.185 ;
        RECT 84.155 141.165 84.430 141.985 ;
        RECT 84.635 141.385 84.805 142.185 ;
        RECT 84.975 141.395 85.145 142.525 ;
        RECT 85.315 141.895 85.485 142.865 ;
        RECT 85.655 142.065 85.825 143.205 ;
        RECT 85.995 142.065 86.330 143.035 ;
        RECT 86.880 142.865 87.135 142.895 ;
        RECT 86.795 142.695 87.135 142.865 ;
        RECT 85.315 141.565 85.510 141.895 ;
        RECT 85.735 141.565 85.990 141.895 ;
        RECT 85.735 141.395 85.905 141.565 ;
        RECT 86.160 141.395 86.330 142.065 ;
        RECT 84.975 141.225 85.905 141.395 ;
        RECT 84.975 141.190 85.150 141.225 ;
        RECT 84.155 140.995 84.435 141.165 ;
        RECT 84.155 140.825 84.430 140.995 ;
        RECT 84.620 140.825 85.150 141.190 ;
        RECT 85.575 140.655 85.905 141.055 ;
        RECT 86.075 140.825 86.330 141.395 ;
        RECT 86.880 142.225 87.135 142.695 ;
        RECT 87.315 142.405 87.600 143.205 ;
        RECT 87.780 142.485 88.110 142.995 ;
        RECT 86.880 141.365 87.060 142.225 ;
        RECT 87.780 141.895 88.030 142.485 ;
        RECT 88.380 142.335 88.550 142.945 ;
        RECT 88.720 142.515 89.050 143.205 ;
        RECT 89.280 142.655 89.520 142.945 ;
        RECT 89.720 142.825 90.140 143.205 ;
        RECT 90.320 142.735 90.950 142.985 ;
        RECT 91.420 142.825 91.750 143.205 ;
        RECT 90.320 142.655 90.490 142.735 ;
        RECT 91.920 142.655 92.090 142.945 ;
        RECT 92.270 142.825 92.650 143.205 ;
        RECT 92.890 142.820 93.720 142.990 ;
        RECT 89.280 142.485 90.490 142.655 ;
        RECT 87.230 141.565 88.030 141.895 ;
        RECT 86.880 140.835 87.135 141.365 ;
        RECT 87.315 140.655 87.600 141.115 ;
        RECT 87.780 140.915 88.030 141.565 ;
        RECT 88.230 142.315 88.550 142.335 ;
        RECT 88.230 142.145 90.150 142.315 ;
        RECT 88.230 141.250 88.420 142.145 ;
        RECT 90.320 141.975 90.490 142.485 ;
        RECT 90.660 142.225 91.180 142.535 ;
        RECT 88.590 141.805 90.490 141.975 ;
        RECT 88.590 141.745 88.920 141.805 ;
        RECT 89.070 141.575 89.400 141.635 ;
        RECT 88.740 141.305 89.400 141.575 ;
        RECT 88.230 140.920 88.550 141.250 ;
        RECT 88.730 140.655 89.390 141.135 ;
        RECT 89.590 141.045 89.760 141.805 ;
        RECT 90.660 141.635 90.840 142.045 ;
        RECT 89.930 141.465 90.260 141.585 ;
        RECT 91.010 141.465 91.180 142.225 ;
        RECT 89.930 141.295 91.180 141.465 ;
        RECT 91.350 142.405 92.720 142.655 ;
        RECT 91.350 141.635 91.540 142.405 ;
        RECT 92.470 142.145 92.720 142.405 ;
        RECT 91.710 141.975 91.960 142.135 ;
        RECT 92.890 141.975 93.060 142.820 ;
        RECT 93.955 142.535 94.125 143.035 ;
        RECT 94.295 142.705 94.625 143.205 ;
        RECT 93.230 142.145 93.730 142.525 ;
        RECT 93.955 142.365 94.650 142.535 ;
        RECT 91.710 141.805 93.060 141.975 ;
        RECT 92.640 141.765 93.060 141.805 ;
        RECT 91.350 141.295 91.770 141.635 ;
        RECT 92.060 141.305 92.470 141.635 ;
        RECT 89.590 140.875 90.440 141.045 ;
        RECT 91.000 140.655 91.320 141.115 ;
        RECT 91.520 140.865 91.770 141.295 ;
        RECT 92.060 140.655 92.470 141.095 ;
        RECT 92.640 141.035 92.810 141.765 ;
        RECT 92.980 141.215 93.330 141.585 ;
        RECT 93.510 141.275 93.730 142.145 ;
        RECT 93.900 141.575 94.310 142.195 ;
        RECT 94.480 141.395 94.650 142.365 ;
        RECT 93.955 141.205 94.650 141.395 ;
        RECT 92.640 140.835 93.655 141.035 ;
        RECT 93.955 140.875 94.125 141.205 ;
        RECT 94.295 140.655 94.625 141.035 ;
        RECT 94.840 140.915 95.065 143.035 ;
        RECT 95.235 142.705 95.565 143.205 ;
        RECT 95.735 142.535 95.905 143.035 ;
        RECT 95.240 142.365 95.905 142.535 ;
        RECT 95.240 141.375 95.470 142.365 ;
        RECT 95.640 141.545 95.990 142.195 ;
        RECT 96.625 142.130 96.895 143.035 ;
        RECT 97.065 142.445 97.395 143.205 ;
        RECT 97.575 142.275 97.745 143.035 ;
        RECT 95.240 141.205 95.905 141.375 ;
        RECT 95.235 140.655 95.565 141.035 ;
        RECT 95.735 140.915 95.905 141.205 ;
        RECT 96.625 141.330 96.795 142.130 ;
        RECT 97.080 142.105 97.745 142.275 ;
        RECT 98.210 142.235 98.540 143.035 ;
        RECT 98.710 142.405 99.040 143.205 ;
        RECT 99.340 142.235 99.670 143.035 ;
        RECT 100.315 142.405 100.565 143.205 ;
        RECT 97.080 141.960 97.250 142.105 ;
        RECT 98.210 142.065 100.645 142.235 ;
        RECT 100.835 142.065 101.005 143.205 ;
        RECT 101.175 142.065 101.515 143.035 ;
        RECT 96.965 141.630 97.250 141.960 ;
        RECT 97.080 141.375 97.250 141.630 ;
        RECT 97.485 141.555 97.815 141.925 ;
        RECT 98.005 141.645 98.355 141.895 ;
        RECT 98.540 141.435 98.710 142.065 ;
        RECT 98.880 141.645 99.210 141.845 ;
        RECT 99.380 141.645 99.710 141.845 ;
        RECT 99.880 141.645 100.300 141.845 ;
        RECT 100.475 141.815 100.645 142.065 ;
        RECT 100.475 141.645 101.170 141.815 ;
        RECT 96.625 140.825 96.885 141.330 ;
        RECT 97.080 141.205 97.745 141.375 ;
        RECT 97.065 140.655 97.395 141.035 ;
        RECT 97.575 140.825 97.745 141.205 ;
        RECT 98.210 140.825 98.710 141.435 ;
        RECT 99.340 141.305 100.565 141.475 ;
        RECT 101.340 141.455 101.515 142.065 ;
        RECT 101.685 142.040 101.975 143.205 ;
        RECT 102.185 142.065 102.415 143.205 ;
        RECT 102.585 142.055 102.915 143.035 ;
        RECT 103.085 142.065 103.295 143.205 ;
        RECT 103.985 142.445 104.500 142.855 ;
        RECT 104.735 142.445 104.905 143.205 ;
        RECT 105.075 142.865 107.105 143.035 ;
        RECT 102.165 141.645 102.495 141.895 ;
        RECT 99.340 140.825 99.670 141.305 ;
        RECT 99.840 140.655 100.065 141.115 ;
        RECT 100.235 140.825 100.565 141.305 ;
        RECT 100.755 140.655 101.005 141.455 ;
        RECT 101.175 140.825 101.515 141.455 ;
        RECT 101.685 140.655 101.975 141.380 ;
        RECT 102.185 140.655 102.415 141.475 ;
        RECT 102.665 141.455 102.915 142.055 ;
        RECT 103.985 141.635 104.325 142.445 ;
        RECT 105.075 142.200 105.245 142.865 ;
        RECT 105.640 142.525 106.765 142.695 ;
        RECT 104.495 142.010 105.245 142.200 ;
        RECT 105.415 142.185 106.425 142.355 ;
        RECT 102.585 140.825 102.915 141.455 ;
        RECT 103.085 140.655 103.295 141.475 ;
        RECT 103.985 141.465 105.215 141.635 ;
        RECT 104.260 140.860 104.505 141.465 ;
        RECT 104.725 140.655 105.235 141.190 ;
        RECT 105.415 140.825 105.605 142.185 ;
        RECT 105.775 141.505 106.050 141.985 ;
        RECT 105.775 141.335 106.055 141.505 ;
        RECT 106.255 141.385 106.425 142.185 ;
        RECT 106.595 141.395 106.765 142.525 ;
        RECT 106.935 141.895 107.105 142.865 ;
        RECT 107.275 142.065 107.445 143.205 ;
        RECT 107.615 142.065 107.950 143.035 ;
        RECT 109.250 142.235 109.580 143.035 ;
        RECT 109.750 142.405 110.080 143.205 ;
        RECT 110.380 142.235 110.710 143.035 ;
        RECT 111.355 142.405 111.605 143.205 ;
        RECT 109.250 142.065 111.685 142.235 ;
        RECT 111.875 142.065 112.045 143.205 ;
        RECT 112.215 142.065 112.555 143.035 ;
        RECT 106.935 141.565 107.130 141.895 ;
        RECT 107.355 141.565 107.610 141.895 ;
        RECT 107.355 141.395 107.525 141.565 ;
        RECT 107.780 141.395 107.950 142.065 ;
        RECT 109.045 141.645 109.395 141.895 ;
        RECT 109.580 141.435 109.750 142.065 ;
        RECT 109.920 141.645 110.250 141.845 ;
        RECT 110.420 141.645 110.750 141.845 ;
        RECT 110.920 141.645 111.340 141.845 ;
        RECT 111.515 141.815 111.685 142.065 ;
        RECT 111.515 141.645 112.210 141.815 ;
        RECT 105.775 140.825 106.050 141.335 ;
        RECT 106.595 141.225 107.525 141.395 ;
        RECT 106.595 141.190 106.770 141.225 ;
        RECT 106.240 140.825 106.770 141.190 ;
        RECT 107.195 140.655 107.525 141.055 ;
        RECT 107.695 140.825 107.950 141.395 ;
        RECT 109.250 140.825 109.750 141.435 ;
        RECT 110.380 141.305 111.605 141.475 ;
        RECT 112.380 141.455 112.555 142.065 ;
        RECT 112.725 142.445 113.240 142.855 ;
        RECT 113.475 142.445 113.645 143.205 ;
        RECT 113.815 142.865 115.845 143.035 ;
        RECT 112.725 141.635 113.065 142.445 ;
        RECT 113.815 142.200 113.985 142.865 ;
        RECT 114.380 142.525 115.505 142.695 ;
        RECT 113.235 142.010 113.985 142.200 ;
        RECT 114.155 142.185 115.165 142.355 ;
        RECT 112.725 141.465 113.955 141.635 ;
        RECT 110.380 140.825 110.710 141.305 ;
        RECT 110.880 140.655 111.105 141.115 ;
        RECT 111.275 140.825 111.605 141.305 ;
        RECT 111.795 140.655 112.045 141.455 ;
        RECT 112.215 140.825 112.555 141.455 ;
        RECT 113.000 140.860 113.245 141.465 ;
        RECT 113.465 140.655 113.975 141.190 ;
        RECT 114.155 140.825 114.345 142.185 ;
        RECT 114.515 141.845 114.790 141.985 ;
        RECT 114.515 141.675 114.795 141.845 ;
        RECT 114.515 140.825 114.790 141.675 ;
        RECT 114.995 141.385 115.165 142.185 ;
        RECT 115.335 141.395 115.505 142.525 ;
        RECT 115.675 141.895 115.845 142.865 ;
        RECT 116.015 142.065 116.185 143.205 ;
        RECT 116.355 142.065 116.690 143.035 ;
        RECT 115.675 141.565 115.870 141.895 ;
        RECT 116.095 141.565 116.350 141.895 ;
        RECT 116.095 141.395 116.265 141.565 ;
        RECT 116.520 141.395 116.690 142.065 ;
        RECT 117.240 142.225 117.495 142.895 ;
        RECT 117.675 142.405 117.960 143.205 ;
        RECT 118.140 142.485 118.470 142.995 ;
        RECT 117.240 141.505 117.420 142.225 ;
        RECT 118.140 141.895 118.390 142.485 ;
        RECT 118.740 142.335 118.910 142.945 ;
        RECT 119.080 142.515 119.410 143.205 ;
        RECT 119.640 142.655 119.880 142.945 ;
        RECT 120.080 142.825 120.500 143.205 ;
        RECT 120.680 142.735 121.310 142.985 ;
        RECT 121.780 142.825 122.110 143.205 ;
        RECT 120.680 142.655 120.850 142.735 ;
        RECT 122.280 142.655 122.450 142.945 ;
        RECT 122.630 142.825 123.010 143.205 ;
        RECT 123.250 142.820 124.080 142.990 ;
        RECT 119.640 142.485 120.850 142.655 ;
        RECT 117.590 141.565 118.390 141.895 ;
        RECT 115.335 141.225 116.265 141.395 ;
        RECT 115.335 141.190 115.510 141.225 ;
        RECT 114.980 140.825 115.510 141.190 ;
        RECT 115.935 140.655 116.265 141.055 ;
        RECT 116.435 140.825 116.690 141.395 ;
        RECT 117.155 141.365 117.420 141.505 ;
        RECT 117.155 141.335 117.495 141.365 ;
        RECT 117.240 140.835 117.495 141.335 ;
        RECT 117.675 140.655 117.960 141.115 ;
        RECT 118.140 140.915 118.390 141.565 ;
        RECT 118.590 142.315 118.910 142.335 ;
        RECT 118.590 142.145 120.510 142.315 ;
        RECT 118.590 141.250 118.780 142.145 ;
        RECT 120.680 141.975 120.850 142.485 ;
        RECT 121.020 142.225 121.540 142.535 ;
        RECT 118.950 141.805 120.850 141.975 ;
        RECT 118.950 141.745 119.280 141.805 ;
        RECT 119.430 141.575 119.760 141.635 ;
        RECT 119.100 141.305 119.760 141.575 ;
        RECT 118.590 140.920 118.910 141.250 ;
        RECT 119.090 140.655 119.750 141.135 ;
        RECT 119.950 141.045 120.120 141.805 ;
        RECT 121.020 141.635 121.200 142.045 ;
        RECT 120.290 141.465 120.620 141.585 ;
        RECT 121.370 141.465 121.540 142.225 ;
        RECT 120.290 141.295 121.540 141.465 ;
        RECT 121.710 142.405 123.080 142.655 ;
        RECT 121.710 141.635 121.900 142.405 ;
        RECT 122.830 142.145 123.080 142.405 ;
        RECT 122.070 141.975 122.320 142.135 ;
        RECT 123.250 141.975 123.420 142.820 ;
        RECT 124.315 142.535 124.485 143.035 ;
        RECT 124.655 142.705 124.985 143.205 ;
        RECT 123.590 142.145 124.090 142.525 ;
        RECT 124.315 142.365 125.010 142.535 ;
        RECT 122.070 141.805 123.420 141.975 ;
        RECT 123.000 141.765 123.420 141.805 ;
        RECT 121.710 141.295 122.130 141.635 ;
        RECT 122.420 141.305 122.830 141.635 ;
        RECT 119.950 140.875 120.800 141.045 ;
        RECT 121.360 140.655 121.680 141.115 ;
        RECT 121.880 140.865 122.130 141.295 ;
        RECT 122.420 140.655 122.830 141.095 ;
        RECT 123.000 141.035 123.170 141.765 ;
        RECT 123.340 141.215 123.690 141.585 ;
        RECT 123.870 141.275 124.090 142.145 ;
        RECT 124.260 141.575 124.670 142.195 ;
        RECT 124.840 141.395 125.010 142.365 ;
        RECT 124.315 141.205 125.010 141.395 ;
        RECT 123.000 140.835 124.015 141.035 ;
        RECT 124.315 140.875 124.485 141.205 ;
        RECT 124.655 140.655 124.985 141.035 ;
        RECT 125.200 140.915 125.425 143.035 ;
        RECT 125.595 142.705 125.925 143.205 ;
        RECT 126.095 142.535 126.265 143.035 ;
        RECT 125.600 142.365 126.265 142.535 ;
        RECT 125.600 141.375 125.830 142.365 ;
        RECT 126.000 141.545 126.350 142.195 ;
        RECT 126.525 142.115 127.735 143.205 ;
        RECT 126.525 141.575 127.045 142.115 ;
        RECT 127.215 141.405 127.735 141.945 ;
        RECT 125.600 141.205 126.265 141.375 ;
        RECT 125.595 140.655 125.925 141.035 ;
        RECT 126.095 140.915 126.265 141.205 ;
        RECT 126.525 140.655 127.735 141.405 ;
        RECT 20.640 140.485 127.820 140.655 ;
        RECT 20.725 139.735 21.935 140.485 ;
        RECT 23.400 139.775 23.655 140.305 ;
        RECT 23.835 140.025 24.120 140.485 ;
        RECT 20.725 139.195 21.245 139.735 ;
        RECT 21.415 139.025 21.935 139.565 ;
        RECT 20.725 137.935 21.935 139.025 ;
        RECT 23.400 138.915 23.580 139.775 ;
        RECT 24.300 139.575 24.550 140.225 ;
        RECT 23.750 139.245 24.550 139.575 ;
        RECT 23.400 138.445 23.655 138.915 ;
        RECT 23.315 138.275 23.655 138.445 ;
        RECT 23.400 138.245 23.655 138.275 ;
        RECT 23.835 137.935 24.120 138.735 ;
        RECT 24.300 138.655 24.550 139.245 ;
        RECT 24.750 139.890 25.070 140.220 ;
        RECT 25.250 140.005 25.910 140.485 ;
        RECT 26.110 140.095 26.960 140.265 ;
        RECT 24.750 138.995 24.940 139.890 ;
        RECT 25.260 139.565 25.920 139.835 ;
        RECT 25.590 139.505 25.920 139.565 ;
        RECT 25.110 139.335 25.440 139.395 ;
        RECT 26.110 139.335 26.280 140.095 ;
        RECT 27.520 140.025 27.840 140.485 ;
        RECT 28.040 139.845 28.290 140.275 ;
        RECT 28.580 140.045 28.990 140.485 ;
        RECT 29.160 140.105 30.175 140.305 ;
        RECT 26.450 139.675 27.700 139.845 ;
        RECT 26.450 139.555 26.780 139.675 ;
        RECT 25.110 139.165 27.010 139.335 ;
        RECT 24.750 138.825 26.670 138.995 ;
        RECT 24.750 138.805 25.070 138.825 ;
        RECT 24.300 138.145 24.630 138.655 ;
        RECT 24.900 138.195 25.070 138.805 ;
        RECT 26.840 138.655 27.010 139.165 ;
        RECT 27.180 139.095 27.360 139.505 ;
        RECT 27.530 138.915 27.700 139.675 ;
        RECT 25.240 137.935 25.570 138.625 ;
        RECT 25.800 138.485 27.010 138.655 ;
        RECT 27.180 138.605 27.700 138.915 ;
        RECT 27.870 139.505 28.290 139.845 ;
        RECT 28.580 139.505 28.990 139.835 ;
        RECT 27.870 138.735 28.060 139.505 ;
        RECT 29.160 139.375 29.330 140.105 ;
        RECT 30.475 139.935 30.645 140.265 ;
        RECT 30.815 140.105 31.145 140.485 ;
        RECT 29.500 139.555 29.850 139.925 ;
        RECT 29.160 139.335 29.580 139.375 ;
        RECT 28.230 139.165 29.580 139.335 ;
        RECT 28.230 139.005 28.480 139.165 ;
        RECT 28.990 138.735 29.240 138.995 ;
        RECT 27.870 138.485 29.240 138.735 ;
        RECT 25.800 138.195 26.040 138.485 ;
        RECT 26.840 138.405 27.010 138.485 ;
        RECT 26.240 137.935 26.660 138.315 ;
        RECT 26.840 138.155 27.470 138.405 ;
        RECT 27.940 137.935 28.270 138.315 ;
        RECT 28.440 138.195 28.610 138.485 ;
        RECT 29.410 138.320 29.580 139.165 ;
        RECT 30.030 138.995 30.250 139.865 ;
        RECT 30.475 139.745 31.170 139.935 ;
        RECT 29.750 138.615 30.250 138.995 ;
        RECT 30.420 138.945 30.830 139.565 ;
        RECT 31.000 138.775 31.170 139.745 ;
        RECT 30.475 138.605 31.170 138.775 ;
        RECT 28.790 137.935 29.170 138.315 ;
        RECT 29.410 138.150 30.240 138.320 ;
        RECT 30.475 138.105 30.645 138.605 ;
        RECT 30.815 137.935 31.145 138.435 ;
        RECT 31.360 138.105 31.585 140.225 ;
        RECT 31.755 140.105 32.085 140.485 ;
        RECT 32.255 139.935 32.425 140.225 ;
        RECT 31.760 139.765 32.425 139.935 ;
        RECT 32.685 139.810 32.945 140.315 ;
        RECT 33.125 140.105 33.455 140.485 ;
        RECT 33.635 139.935 33.805 140.315 ;
        RECT 31.760 138.775 31.990 139.765 ;
        RECT 32.160 138.945 32.510 139.595 ;
        RECT 32.685 139.010 32.855 139.810 ;
        RECT 33.140 139.765 33.805 139.935 ;
        RECT 33.140 139.510 33.310 139.765 ;
        RECT 34.065 139.735 35.275 140.485 ;
        RECT 33.025 139.180 33.310 139.510 ;
        RECT 33.545 139.215 33.875 139.585 ;
        RECT 33.140 139.035 33.310 139.180 ;
        RECT 31.760 138.605 32.425 138.775 ;
        RECT 31.755 137.935 32.085 138.435 ;
        RECT 32.255 138.105 32.425 138.605 ;
        RECT 32.685 138.105 32.955 139.010 ;
        RECT 33.140 138.865 33.805 139.035 ;
        RECT 33.125 137.935 33.455 138.695 ;
        RECT 33.635 138.105 33.805 138.865 ;
        RECT 34.065 139.025 34.585 139.565 ;
        RECT 34.755 139.195 35.275 139.735 ;
        RECT 35.485 139.665 35.715 140.485 ;
        RECT 35.885 139.685 36.215 140.315 ;
        RECT 35.465 139.245 35.795 139.495 ;
        RECT 35.965 139.085 36.215 139.685 ;
        RECT 36.385 139.665 36.595 140.485 ;
        RECT 37.285 139.760 37.575 140.485 ;
        RECT 38.205 139.715 40.795 140.485 ;
        RECT 34.065 137.935 35.275 139.025 ;
        RECT 35.485 137.935 35.715 139.075 ;
        RECT 35.885 138.105 36.215 139.085 ;
        RECT 36.385 137.935 36.595 139.075 ;
        RECT 37.285 137.935 37.575 139.100 ;
        RECT 38.205 139.025 39.415 139.545 ;
        RECT 39.585 139.195 40.795 139.715 ;
        RECT 40.965 139.810 41.225 140.315 ;
        RECT 41.405 140.105 41.735 140.485 ;
        RECT 41.915 139.935 42.085 140.315 ;
        RECT 38.205 137.935 40.795 139.025 ;
        RECT 40.965 139.010 41.135 139.810 ;
        RECT 41.420 139.765 42.085 139.935 ;
        RECT 42.545 139.855 42.875 140.215 ;
        RECT 43.495 140.025 43.745 140.485 ;
        RECT 43.915 140.025 44.475 140.315 ;
        RECT 41.420 139.510 41.590 139.765 ;
        RECT 42.545 139.665 43.935 139.855 ;
        RECT 41.305 139.180 41.590 139.510 ;
        RECT 41.825 139.215 42.155 139.585 ;
        RECT 43.765 139.575 43.935 139.665 ;
        RECT 42.360 139.245 43.035 139.495 ;
        RECT 43.255 139.245 43.595 139.495 ;
        RECT 43.765 139.245 44.055 139.575 ;
        RECT 41.420 139.035 41.590 139.180 ;
        RECT 40.965 138.105 41.235 139.010 ;
        RECT 41.420 138.865 42.085 139.035 ;
        RECT 42.360 138.885 42.625 139.245 ;
        RECT 43.765 138.995 43.935 139.245 ;
        RECT 41.405 137.935 41.735 138.695 ;
        RECT 41.915 138.105 42.085 138.865 ;
        RECT 42.995 138.825 43.935 138.995 ;
        RECT 42.545 137.935 42.825 138.605 ;
        RECT 42.995 138.275 43.295 138.825 ;
        RECT 44.225 138.655 44.475 140.025 ;
        RECT 44.845 139.855 45.175 140.215 ;
        RECT 45.795 140.025 46.045 140.485 ;
        RECT 46.215 140.025 46.775 140.315 ;
        RECT 44.845 139.665 46.235 139.855 ;
        RECT 46.065 139.575 46.235 139.665 ;
        RECT 44.660 139.245 45.335 139.495 ;
        RECT 45.555 139.245 45.895 139.495 ;
        RECT 46.065 139.245 46.355 139.575 ;
        RECT 44.660 138.885 44.925 139.245 ;
        RECT 46.065 138.995 46.235 139.245 ;
        RECT 43.495 137.935 43.825 138.655 ;
        RECT 44.015 138.105 44.475 138.655 ;
        RECT 45.295 138.825 46.235 138.995 ;
        RECT 44.845 137.935 45.125 138.605 ;
        RECT 45.295 138.275 45.595 138.825 ;
        RECT 46.525 138.655 46.775 140.025 ;
        RECT 46.945 139.715 49.535 140.485 ;
        RECT 45.795 137.935 46.125 138.655 ;
        RECT 46.315 138.105 46.775 138.655 ;
        RECT 46.945 139.025 48.155 139.545 ;
        RECT 48.325 139.195 49.535 139.715 ;
        RECT 49.705 140.025 50.265 140.315 ;
        RECT 50.435 140.025 50.685 140.485 ;
        RECT 46.945 137.935 49.535 139.025 ;
        RECT 49.705 138.655 49.955 140.025 ;
        RECT 51.305 139.855 51.635 140.215 ;
        RECT 50.245 139.665 51.635 139.855 ;
        RECT 52.005 140.025 52.565 140.315 ;
        RECT 52.735 140.025 52.985 140.485 ;
        RECT 50.245 139.575 50.415 139.665 ;
        RECT 50.125 139.245 50.415 139.575 ;
        RECT 50.585 139.245 50.925 139.495 ;
        RECT 51.145 139.245 51.820 139.495 ;
        RECT 50.245 138.995 50.415 139.245 ;
        RECT 50.245 138.825 51.185 138.995 ;
        RECT 51.555 138.885 51.820 139.245 ;
        RECT 49.705 138.105 50.165 138.655 ;
        RECT 50.355 137.935 50.685 138.655 ;
        RECT 50.885 138.275 51.185 138.825 ;
        RECT 52.005 138.655 52.255 140.025 ;
        RECT 53.605 139.855 53.935 140.215 ;
        RECT 52.545 139.665 53.935 139.855 ;
        RECT 54.305 139.715 55.975 140.485 ;
        RECT 56.150 139.940 61.495 140.485 ;
        RECT 52.545 139.575 52.715 139.665 ;
        RECT 52.425 139.245 52.715 139.575 ;
        RECT 52.885 139.245 53.225 139.495 ;
        RECT 53.445 139.245 54.120 139.495 ;
        RECT 52.545 138.995 52.715 139.245 ;
        RECT 52.545 138.825 53.485 138.995 ;
        RECT 53.855 138.885 54.120 139.245 ;
        RECT 54.305 139.025 55.055 139.545 ;
        RECT 55.225 139.195 55.975 139.715 ;
        RECT 51.355 137.935 51.635 138.605 ;
        RECT 52.005 138.105 52.465 138.655 ;
        RECT 52.655 137.935 52.985 138.655 ;
        RECT 53.185 138.275 53.485 138.825 ;
        RECT 53.655 137.935 53.935 138.605 ;
        RECT 54.305 137.935 55.975 139.025 ;
        RECT 57.740 138.370 58.090 139.620 ;
        RECT 59.570 139.110 59.910 139.940 ;
        RECT 61.755 139.935 61.925 140.315 ;
        RECT 62.105 140.105 62.435 140.485 ;
        RECT 61.755 139.765 62.420 139.935 ;
        RECT 62.615 139.810 62.875 140.315 ;
        RECT 61.685 139.215 62.015 139.585 ;
        RECT 62.250 139.510 62.420 139.765 ;
        RECT 62.250 139.180 62.535 139.510 ;
        RECT 62.250 139.035 62.420 139.180 ;
        RECT 61.755 138.865 62.420 139.035 ;
        RECT 62.705 139.010 62.875 139.810 ;
        RECT 63.045 139.760 63.335 140.485 ;
        RECT 63.505 139.715 66.095 140.485 ;
        RECT 56.150 137.935 61.495 138.370 ;
        RECT 61.755 138.105 61.925 138.865 ;
        RECT 62.105 137.935 62.435 138.695 ;
        RECT 62.605 138.105 62.875 139.010 ;
        RECT 63.045 137.935 63.335 139.100 ;
        RECT 63.505 139.025 64.715 139.545 ;
        RECT 64.885 139.195 66.095 139.715 ;
        RECT 66.265 139.685 66.605 140.315 ;
        RECT 66.775 139.685 67.025 140.485 ;
        RECT 67.215 139.835 67.545 140.315 ;
        RECT 67.715 140.025 67.940 140.485 ;
        RECT 68.110 139.835 68.440 140.315 ;
        RECT 66.265 139.635 66.495 139.685 ;
        RECT 67.215 139.665 68.440 139.835 ;
        RECT 69.070 139.705 69.570 140.315 ;
        RECT 69.950 139.720 70.405 140.485 ;
        RECT 70.680 140.105 71.980 140.315 ;
        RECT 72.235 140.125 72.565 140.485 ;
        RECT 71.810 139.955 71.980 140.105 ;
        RECT 72.735 139.985 72.995 140.315 ;
        RECT 72.765 139.975 72.995 139.985 ;
        RECT 66.265 139.075 66.440 139.635 ;
        RECT 66.610 139.325 67.305 139.495 ;
        RECT 67.135 139.075 67.305 139.325 ;
        RECT 67.480 139.295 67.900 139.495 ;
        RECT 68.070 139.295 68.400 139.495 ;
        RECT 68.570 139.295 68.900 139.495 ;
        RECT 69.070 139.075 69.240 139.705 ;
        RECT 70.880 139.495 71.100 139.895 ;
        RECT 69.425 139.245 69.775 139.495 ;
        RECT 69.945 139.295 70.435 139.495 ;
        RECT 70.625 139.285 71.100 139.495 ;
        RECT 71.345 139.495 71.555 139.895 ;
        RECT 71.810 139.830 72.565 139.955 ;
        RECT 71.810 139.785 72.655 139.830 ;
        RECT 72.385 139.665 72.655 139.785 ;
        RECT 71.345 139.285 71.675 139.495 ;
        RECT 71.845 139.225 72.255 139.530 ;
        RECT 63.505 137.935 66.095 139.025 ;
        RECT 66.265 138.105 66.605 139.075 ;
        RECT 66.775 137.935 66.945 139.075 ;
        RECT 67.135 138.905 69.570 139.075 ;
        RECT 67.215 137.935 67.465 138.735 ;
        RECT 68.110 138.105 68.440 138.905 ;
        RECT 68.740 137.935 69.070 138.735 ;
        RECT 69.240 138.105 69.570 138.905 ;
        RECT 69.950 139.055 71.125 139.115 ;
        RECT 72.485 139.090 72.655 139.665 ;
        RECT 72.455 139.055 72.655 139.090 ;
        RECT 69.950 138.945 72.655 139.055 ;
        RECT 69.950 138.325 70.205 138.945 ;
        RECT 70.795 138.885 72.595 138.945 ;
        RECT 70.795 138.855 71.125 138.885 ;
        RECT 72.825 138.785 72.995 139.975 ;
        RECT 73.625 139.715 75.295 140.485 ;
        RECT 75.470 139.940 80.815 140.485 ;
        RECT 70.455 138.685 70.640 138.775 ;
        RECT 71.230 138.685 72.065 138.695 ;
        RECT 70.455 138.485 72.065 138.685 ;
        RECT 70.455 138.445 70.685 138.485 ;
        RECT 69.950 138.105 70.285 138.325 ;
        RECT 71.290 137.935 71.645 138.315 ;
        RECT 71.815 138.105 72.065 138.485 ;
        RECT 72.315 137.935 72.565 138.715 ;
        RECT 72.735 138.105 72.995 138.785 ;
        RECT 73.625 139.025 74.375 139.545 ;
        RECT 74.545 139.195 75.295 139.715 ;
        RECT 73.625 137.935 75.295 139.025 ;
        RECT 77.060 138.370 77.410 139.620 ;
        RECT 78.890 139.110 79.230 139.940 ;
        RECT 81.185 139.855 81.515 140.215 ;
        RECT 82.135 140.025 82.385 140.485 ;
        RECT 82.555 140.025 83.115 140.315 ;
        RECT 81.185 139.665 82.575 139.855 ;
        RECT 82.405 139.575 82.575 139.665 ;
        RECT 81.000 139.245 81.675 139.495 ;
        RECT 81.895 139.245 82.235 139.495 ;
        RECT 82.405 139.245 82.695 139.575 ;
        RECT 81.000 138.885 81.265 139.245 ;
        RECT 82.405 138.995 82.575 139.245 ;
        RECT 81.635 138.825 82.575 138.995 ;
        RECT 75.470 137.935 80.815 138.370 ;
        RECT 81.185 137.935 81.465 138.605 ;
        RECT 81.635 138.275 81.935 138.825 ;
        RECT 82.865 138.655 83.115 140.025 ;
        RECT 83.745 139.715 87.255 140.485 ;
        RECT 82.135 137.935 82.465 138.655 ;
        RECT 82.655 138.105 83.115 138.655 ;
        RECT 83.745 139.025 85.435 139.545 ;
        RECT 85.605 139.195 87.255 139.715 ;
        RECT 87.465 139.665 87.695 140.485 ;
        RECT 87.865 139.685 88.195 140.315 ;
        RECT 87.445 139.245 87.775 139.495 ;
        RECT 87.945 139.085 88.195 139.685 ;
        RECT 88.365 139.665 88.575 140.485 ;
        RECT 88.805 139.760 89.095 140.485 ;
        RECT 90.100 139.775 90.355 140.305 ;
        RECT 90.535 140.025 90.820 140.485 ;
        RECT 83.745 137.935 87.255 139.025 ;
        RECT 87.465 137.935 87.695 139.075 ;
        RECT 87.865 138.105 88.195 139.085 ;
        RECT 88.365 137.935 88.575 139.075 ;
        RECT 88.805 137.935 89.095 139.100 ;
        RECT 90.100 138.915 90.280 139.775 ;
        RECT 91.000 139.575 91.250 140.225 ;
        RECT 90.450 139.245 91.250 139.575 ;
        RECT 90.100 138.445 90.355 138.915 ;
        RECT 90.015 138.275 90.355 138.445 ;
        RECT 90.100 138.245 90.355 138.275 ;
        RECT 90.535 137.935 90.820 138.735 ;
        RECT 91.000 138.655 91.250 139.245 ;
        RECT 91.450 139.890 91.770 140.220 ;
        RECT 91.950 140.005 92.610 140.485 ;
        RECT 92.810 140.095 93.660 140.265 ;
        RECT 91.450 138.995 91.640 139.890 ;
        RECT 91.960 139.565 92.620 139.835 ;
        RECT 92.290 139.505 92.620 139.565 ;
        RECT 91.810 139.335 92.140 139.395 ;
        RECT 92.810 139.335 92.980 140.095 ;
        RECT 94.220 140.025 94.540 140.485 ;
        RECT 94.740 139.845 94.990 140.275 ;
        RECT 95.280 140.045 95.690 140.485 ;
        RECT 95.860 140.105 96.875 140.305 ;
        RECT 93.150 139.675 94.400 139.845 ;
        RECT 93.150 139.555 93.480 139.675 ;
        RECT 91.810 139.165 93.710 139.335 ;
        RECT 91.450 138.825 93.370 138.995 ;
        RECT 91.450 138.805 91.770 138.825 ;
        RECT 91.000 138.145 91.330 138.655 ;
        RECT 91.600 138.195 91.770 138.805 ;
        RECT 93.540 138.655 93.710 139.165 ;
        RECT 93.880 139.095 94.060 139.505 ;
        RECT 94.230 138.915 94.400 139.675 ;
        RECT 91.940 137.935 92.270 138.625 ;
        RECT 92.500 138.485 93.710 138.655 ;
        RECT 93.880 138.605 94.400 138.915 ;
        RECT 94.570 139.505 94.990 139.845 ;
        RECT 95.280 139.505 95.690 139.835 ;
        RECT 94.570 138.735 94.760 139.505 ;
        RECT 95.860 139.375 96.030 140.105 ;
        RECT 97.175 139.935 97.345 140.265 ;
        RECT 97.515 140.105 97.845 140.485 ;
        RECT 96.200 139.555 96.550 139.925 ;
        RECT 95.860 139.335 96.280 139.375 ;
        RECT 94.930 139.165 96.280 139.335 ;
        RECT 94.930 139.005 95.180 139.165 ;
        RECT 95.690 138.735 95.940 138.995 ;
        RECT 94.570 138.485 95.940 138.735 ;
        RECT 92.500 138.195 92.740 138.485 ;
        RECT 93.540 138.405 93.710 138.485 ;
        RECT 92.940 137.935 93.360 138.315 ;
        RECT 93.540 138.155 94.170 138.405 ;
        RECT 94.640 137.935 94.970 138.315 ;
        RECT 95.140 138.195 95.310 138.485 ;
        RECT 96.110 138.320 96.280 139.165 ;
        RECT 96.730 138.995 96.950 139.865 ;
        RECT 97.175 139.745 97.870 139.935 ;
        RECT 96.450 138.615 96.950 138.995 ;
        RECT 97.120 138.945 97.530 139.565 ;
        RECT 97.700 138.775 97.870 139.745 ;
        RECT 97.175 138.605 97.870 138.775 ;
        RECT 95.490 137.935 95.870 138.315 ;
        RECT 96.110 138.150 96.940 138.320 ;
        RECT 97.175 138.105 97.345 138.605 ;
        RECT 97.515 137.935 97.845 138.435 ;
        RECT 98.060 138.105 98.285 140.225 ;
        RECT 98.455 140.105 98.785 140.485 ;
        RECT 98.955 139.935 99.125 140.225 ;
        RECT 98.460 139.765 99.125 139.935 ;
        RECT 99.760 139.775 100.015 140.305 ;
        RECT 100.195 140.025 100.480 140.485 ;
        RECT 98.460 138.775 98.690 139.765 ;
        RECT 98.860 138.945 99.210 139.595 ;
        RECT 99.760 138.915 99.940 139.775 ;
        RECT 100.660 139.575 100.910 140.225 ;
        RECT 100.110 139.245 100.910 139.575 ;
        RECT 98.460 138.605 99.125 138.775 ;
        RECT 98.455 137.935 98.785 138.435 ;
        RECT 98.955 138.105 99.125 138.605 ;
        RECT 99.760 138.445 100.015 138.915 ;
        RECT 99.675 138.275 100.015 138.445 ;
        RECT 99.760 138.245 100.015 138.275 ;
        RECT 100.195 137.935 100.480 138.735 ;
        RECT 100.660 138.655 100.910 139.245 ;
        RECT 101.110 139.890 101.430 140.220 ;
        RECT 101.610 140.005 102.270 140.485 ;
        RECT 102.470 140.095 103.320 140.265 ;
        RECT 101.110 138.995 101.300 139.890 ;
        RECT 101.620 139.565 102.280 139.835 ;
        RECT 101.950 139.505 102.280 139.565 ;
        RECT 101.470 139.335 101.800 139.395 ;
        RECT 102.470 139.335 102.640 140.095 ;
        RECT 103.880 140.025 104.200 140.485 ;
        RECT 104.400 139.845 104.650 140.275 ;
        RECT 104.940 140.045 105.350 140.485 ;
        RECT 105.520 140.105 106.535 140.305 ;
        RECT 102.810 139.675 104.060 139.845 ;
        RECT 102.810 139.555 103.140 139.675 ;
        RECT 101.470 139.165 103.370 139.335 ;
        RECT 101.110 138.825 103.030 138.995 ;
        RECT 101.110 138.805 101.430 138.825 ;
        RECT 100.660 138.145 100.990 138.655 ;
        RECT 101.260 138.195 101.430 138.805 ;
        RECT 103.200 138.655 103.370 139.165 ;
        RECT 103.540 139.095 103.720 139.505 ;
        RECT 103.890 138.915 104.060 139.675 ;
        RECT 101.600 137.935 101.930 138.625 ;
        RECT 102.160 138.485 103.370 138.655 ;
        RECT 103.540 138.605 104.060 138.915 ;
        RECT 104.230 139.505 104.650 139.845 ;
        RECT 104.940 139.505 105.350 139.835 ;
        RECT 104.230 138.735 104.420 139.505 ;
        RECT 105.520 139.375 105.690 140.105 ;
        RECT 106.835 139.935 107.005 140.265 ;
        RECT 107.175 140.105 107.505 140.485 ;
        RECT 105.860 139.555 106.210 139.925 ;
        RECT 105.520 139.335 105.940 139.375 ;
        RECT 104.590 139.165 105.940 139.335 ;
        RECT 104.590 139.005 104.840 139.165 ;
        RECT 105.350 138.735 105.600 138.995 ;
        RECT 104.230 138.485 105.600 138.735 ;
        RECT 102.160 138.195 102.400 138.485 ;
        RECT 103.200 138.405 103.370 138.485 ;
        RECT 102.600 137.935 103.020 138.315 ;
        RECT 103.200 138.155 103.830 138.405 ;
        RECT 104.300 137.935 104.630 138.315 ;
        RECT 104.800 138.195 104.970 138.485 ;
        RECT 105.770 138.320 105.940 139.165 ;
        RECT 106.390 138.995 106.610 139.865 ;
        RECT 106.835 139.745 107.530 139.935 ;
        RECT 106.110 138.615 106.610 138.995 ;
        RECT 106.780 138.945 107.190 139.565 ;
        RECT 107.360 138.775 107.530 139.745 ;
        RECT 106.835 138.605 107.530 138.775 ;
        RECT 105.150 137.935 105.530 138.315 ;
        RECT 105.770 138.150 106.600 138.320 ;
        RECT 106.835 138.105 107.005 138.605 ;
        RECT 107.175 137.935 107.505 138.435 ;
        RECT 107.720 138.105 107.945 140.225 ;
        RECT 108.115 140.105 108.445 140.485 ;
        RECT 108.615 139.935 108.785 140.225 ;
        RECT 108.120 139.765 108.785 139.935 ;
        RECT 109.045 139.810 109.305 140.315 ;
        RECT 109.485 140.105 109.815 140.485 ;
        RECT 109.995 139.935 110.165 140.315 ;
        RECT 108.120 138.775 108.350 139.765 ;
        RECT 108.520 138.945 108.870 139.595 ;
        RECT 109.045 139.010 109.215 139.810 ;
        RECT 109.500 139.765 110.165 139.935 ;
        RECT 109.500 139.510 109.670 139.765 ;
        RECT 110.700 139.675 110.945 140.280 ;
        RECT 111.165 139.950 111.675 140.485 ;
        RECT 109.385 139.180 109.670 139.510 ;
        RECT 109.905 139.215 110.235 139.585 ;
        RECT 110.425 139.505 111.655 139.675 ;
        RECT 109.500 139.035 109.670 139.180 ;
        RECT 108.120 138.605 108.785 138.775 ;
        RECT 108.115 137.935 108.445 138.435 ;
        RECT 108.615 138.105 108.785 138.605 ;
        RECT 109.045 138.105 109.315 139.010 ;
        RECT 109.500 138.865 110.165 139.035 ;
        RECT 109.485 137.935 109.815 138.695 ;
        RECT 109.995 138.105 110.165 138.865 ;
        RECT 110.425 138.695 110.765 139.505 ;
        RECT 110.935 138.940 111.685 139.130 ;
        RECT 110.425 138.285 110.940 138.695 ;
        RECT 111.175 137.935 111.345 138.695 ;
        RECT 111.515 138.275 111.685 138.940 ;
        RECT 111.855 138.955 112.045 140.315 ;
        RECT 112.215 140.145 112.490 140.315 ;
        RECT 112.215 139.975 112.495 140.145 ;
        RECT 112.215 139.155 112.490 139.975 ;
        RECT 112.680 139.950 113.210 140.315 ;
        RECT 113.635 140.085 113.965 140.485 ;
        RECT 113.035 139.915 113.210 139.950 ;
        RECT 112.695 138.955 112.865 139.755 ;
        RECT 111.855 138.785 112.865 138.955 ;
        RECT 113.035 139.745 113.965 139.915 ;
        RECT 114.135 139.745 114.390 140.315 ;
        RECT 114.565 139.760 114.855 140.485 ;
        RECT 115.400 139.775 115.655 140.305 ;
        RECT 115.835 140.025 116.120 140.485 ;
        RECT 113.035 138.615 113.205 139.745 ;
        RECT 113.795 139.575 113.965 139.745 ;
        RECT 112.080 138.445 113.205 138.615 ;
        RECT 113.375 139.245 113.570 139.575 ;
        RECT 113.795 139.245 114.050 139.575 ;
        RECT 113.375 138.275 113.545 139.245 ;
        RECT 114.220 139.075 114.390 139.745 ;
        RECT 115.400 139.125 115.580 139.775 ;
        RECT 116.300 139.575 116.550 140.225 ;
        RECT 115.750 139.245 116.550 139.575 ;
        RECT 111.515 138.105 113.545 138.275 ;
        RECT 113.715 137.935 113.885 139.075 ;
        RECT 114.055 138.105 114.390 139.075 ;
        RECT 114.565 137.935 114.855 139.100 ;
        RECT 115.315 138.955 115.580 139.125 ;
        RECT 115.400 138.915 115.580 138.955 ;
        RECT 115.400 138.245 115.655 138.915 ;
        RECT 115.835 137.935 116.120 138.735 ;
        RECT 116.300 138.655 116.550 139.245 ;
        RECT 116.750 139.890 117.070 140.220 ;
        RECT 117.250 140.005 117.910 140.485 ;
        RECT 118.110 140.095 118.960 140.265 ;
        RECT 116.750 138.995 116.940 139.890 ;
        RECT 117.260 139.565 117.920 139.835 ;
        RECT 117.590 139.505 117.920 139.565 ;
        RECT 117.110 139.335 117.440 139.395 ;
        RECT 118.110 139.335 118.280 140.095 ;
        RECT 119.520 140.025 119.840 140.485 ;
        RECT 120.040 139.845 120.290 140.275 ;
        RECT 120.580 140.045 120.990 140.485 ;
        RECT 121.160 140.105 122.175 140.305 ;
        RECT 118.450 139.675 119.700 139.845 ;
        RECT 118.450 139.555 118.780 139.675 ;
        RECT 117.110 139.165 119.010 139.335 ;
        RECT 116.750 138.825 118.670 138.995 ;
        RECT 116.750 138.805 117.070 138.825 ;
        RECT 116.300 138.145 116.630 138.655 ;
        RECT 116.900 138.195 117.070 138.805 ;
        RECT 118.840 138.655 119.010 139.165 ;
        RECT 119.180 139.095 119.360 139.505 ;
        RECT 119.530 138.915 119.700 139.675 ;
        RECT 117.240 137.935 117.570 138.625 ;
        RECT 117.800 138.485 119.010 138.655 ;
        RECT 119.180 138.605 119.700 138.915 ;
        RECT 119.870 139.505 120.290 139.845 ;
        RECT 120.580 139.505 120.990 139.835 ;
        RECT 119.870 138.735 120.060 139.505 ;
        RECT 121.160 139.375 121.330 140.105 ;
        RECT 122.475 139.935 122.645 140.265 ;
        RECT 122.815 140.105 123.145 140.485 ;
        RECT 121.500 139.555 121.850 139.925 ;
        RECT 121.160 139.335 121.580 139.375 ;
        RECT 120.230 139.165 121.580 139.335 ;
        RECT 120.230 139.005 120.480 139.165 ;
        RECT 120.990 138.735 121.240 138.995 ;
        RECT 119.870 138.485 121.240 138.735 ;
        RECT 117.800 138.195 118.040 138.485 ;
        RECT 118.840 138.405 119.010 138.485 ;
        RECT 118.240 137.935 118.660 138.315 ;
        RECT 118.840 138.155 119.470 138.405 ;
        RECT 119.940 137.935 120.270 138.315 ;
        RECT 120.440 138.195 120.610 138.485 ;
        RECT 121.410 138.320 121.580 139.165 ;
        RECT 122.030 138.995 122.250 139.865 ;
        RECT 122.475 139.745 123.170 139.935 ;
        RECT 121.750 138.615 122.250 138.995 ;
        RECT 122.420 138.945 122.830 139.565 ;
        RECT 123.000 138.775 123.170 139.745 ;
        RECT 122.475 138.605 123.170 138.775 ;
        RECT 120.790 137.935 121.170 138.315 ;
        RECT 121.410 138.150 122.240 138.320 ;
        RECT 122.475 138.105 122.645 138.605 ;
        RECT 122.815 137.935 123.145 138.435 ;
        RECT 123.360 138.105 123.585 140.225 ;
        RECT 123.755 140.105 124.085 140.485 ;
        RECT 124.255 139.935 124.425 140.225 ;
        RECT 123.760 139.765 124.425 139.935 ;
        RECT 123.760 138.775 123.990 139.765 ;
        RECT 124.685 139.715 126.355 140.485 ;
        RECT 126.525 139.735 127.735 140.485 ;
        RECT 124.160 138.945 124.510 139.595 ;
        RECT 124.685 139.025 125.435 139.545 ;
        RECT 125.605 139.195 126.355 139.715 ;
        RECT 126.525 139.025 127.045 139.565 ;
        RECT 127.215 139.195 127.735 139.735 ;
        RECT 123.760 138.605 124.425 138.775 ;
        RECT 123.755 137.935 124.085 138.435 ;
        RECT 124.255 138.105 124.425 138.605 ;
        RECT 124.685 137.935 126.355 139.025 ;
        RECT 126.525 137.935 127.735 139.025 ;
        RECT 20.640 137.765 127.820 137.935 ;
        RECT 20.725 136.675 21.935 137.765 ;
        RECT 20.725 135.965 21.245 136.505 ;
        RECT 21.415 136.135 21.935 136.675 ;
        RECT 22.565 136.675 24.235 137.765 ;
        RECT 22.565 136.155 23.315 136.675 ;
        RECT 24.405 136.600 24.695 137.765 ;
        RECT 24.865 136.675 26.535 137.765 ;
        RECT 23.485 135.985 24.235 136.505 ;
        RECT 24.865 136.155 25.615 136.675 ;
        RECT 26.765 136.625 26.975 137.765 ;
        RECT 27.145 136.615 27.475 137.595 ;
        RECT 27.645 136.625 27.875 137.765 ;
        RECT 28.085 137.005 28.600 137.415 ;
        RECT 28.835 137.005 29.005 137.765 ;
        RECT 29.175 137.425 31.205 137.595 ;
        RECT 25.785 135.985 26.535 136.505 ;
        RECT 20.725 135.215 21.935 135.965 ;
        RECT 22.565 135.215 24.235 135.985 ;
        RECT 24.405 135.215 24.695 135.940 ;
        RECT 24.865 135.215 26.535 135.985 ;
        RECT 26.765 135.215 26.975 136.035 ;
        RECT 27.145 136.015 27.395 136.615 ;
        RECT 27.565 136.205 27.895 136.455 ;
        RECT 28.085 136.195 28.425 137.005 ;
        RECT 29.175 136.760 29.345 137.425 ;
        RECT 29.740 137.085 30.865 137.255 ;
        RECT 28.595 136.570 29.345 136.760 ;
        RECT 29.515 136.745 30.525 136.915 ;
        RECT 27.145 135.385 27.475 136.015 ;
        RECT 27.645 135.215 27.875 136.035 ;
        RECT 28.085 136.025 29.315 136.195 ;
        RECT 28.360 135.420 28.605 136.025 ;
        RECT 28.825 135.215 29.335 135.750 ;
        RECT 29.515 135.385 29.705 136.745 ;
        RECT 29.875 136.405 30.150 136.545 ;
        RECT 29.875 136.235 30.155 136.405 ;
        RECT 29.875 135.385 30.150 136.235 ;
        RECT 30.355 135.945 30.525 136.745 ;
        RECT 30.695 135.955 30.865 137.085 ;
        RECT 31.035 136.455 31.205 137.425 ;
        RECT 31.375 136.625 31.545 137.765 ;
        RECT 31.715 136.625 32.050 137.595 ;
        RECT 31.035 136.125 31.230 136.455 ;
        RECT 31.455 136.125 31.710 136.455 ;
        RECT 31.455 135.955 31.625 136.125 ;
        RECT 31.880 135.955 32.050 136.625 ;
        RECT 30.695 135.785 31.625 135.955 ;
        RECT 30.695 135.750 30.870 135.785 ;
        RECT 30.340 135.385 30.870 135.750 ;
        RECT 31.295 135.215 31.625 135.615 ;
        RECT 31.795 135.385 32.050 135.955 ;
        RECT 32.600 136.785 32.855 137.455 ;
        RECT 33.035 136.965 33.320 137.765 ;
        RECT 33.500 137.045 33.830 137.555 ;
        RECT 32.600 135.925 32.780 136.785 ;
        RECT 33.500 136.455 33.750 137.045 ;
        RECT 34.100 136.895 34.270 137.505 ;
        RECT 34.440 137.075 34.770 137.765 ;
        RECT 35.000 137.215 35.240 137.505 ;
        RECT 35.440 137.385 35.860 137.765 ;
        RECT 36.040 137.295 36.670 137.545 ;
        RECT 37.140 137.385 37.470 137.765 ;
        RECT 36.040 137.215 36.210 137.295 ;
        RECT 37.640 137.215 37.810 137.505 ;
        RECT 37.990 137.385 38.370 137.765 ;
        RECT 38.610 137.380 39.440 137.550 ;
        RECT 35.000 137.045 36.210 137.215 ;
        RECT 32.950 136.125 33.750 136.455 ;
        RECT 32.600 135.725 32.855 135.925 ;
        RECT 32.515 135.555 32.855 135.725 ;
        RECT 32.600 135.395 32.855 135.555 ;
        RECT 33.035 135.215 33.320 135.675 ;
        RECT 33.500 135.475 33.750 136.125 ;
        RECT 33.950 136.875 34.270 136.895 ;
        RECT 33.950 136.705 35.870 136.875 ;
        RECT 33.950 135.810 34.140 136.705 ;
        RECT 36.040 136.535 36.210 137.045 ;
        RECT 36.380 136.785 36.900 137.095 ;
        RECT 34.310 136.365 36.210 136.535 ;
        RECT 34.310 136.305 34.640 136.365 ;
        RECT 34.790 136.135 35.120 136.195 ;
        RECT 34.460 135.865 35.120 136.135 ;
        RECT 33.950 135.480 34.270 135.810 ;
        RECT 34.450 135.215 35.110 135.695 ;
        RECT 35.310 135.605 35.480 136.365 ;
        RECT 36.380 136.195 36.560 136.605 ;
        RECT 35.650 136.025 35.980 136.145 ;
        RECT 36.730 136.025 36.900 136.785 ;
        RECT 35.650 135.855 36.900 136.025 ;
        RECT 37.070 136.965 38.440 137.215 ;
        RECT 37.070 136.195 37.260 136.965 ;
        RECT 38.190 136.705 38.440 136.965 ;
        RECT 37.430 136.535 37.680 136.695 ;
        RECT 38.610 136.535 38.780 137.380 ;
        RECT 39.675 137.095 39.845 137.595 ;
        RECT 40.015 137.265 40.345 137.765 ;
        RECT 38.950 136.705 39.450 137.085 ;
        RECT 39.675 136.925 40.370 137.095 ;
        RECT 37.430 136.365 38.780 136.535 ;
        RECT 38.360 136.325 38.780 136.365 ;
        RECT 37.070 135.855 37.490 136.195 ;
        RECT 37.780 135.865 38.190 136.195 ;
        RECT 35.310 135.435 36.160 135.605 ;
        RECT 36.720 135.215 37.040 135.675 ;
        RECT 37.240 135.425 37.490 135.855 ;
        RECT 37.780 135.215 38.190 135.655 ;
        RECT 38.360 135.595 38.530 136.325 ;
        RECT 38.700 135.775 39.050 136.145 ;
        RECT 39.230 135.835 39.450 136.705 ;
        RECT 39.620 136.135 40.030 136.755 ;
        RECT 40.200 135.955 40.370 136.925 ;
        RECT 39.675 135.765 40.370 135.955 ;
        RECT 38.360 135.395 39.375 135.595 ;
        RECT 39.675 135.435 39.845 135.765 ;
        RECT 40.015 135.215 40.345 135.595 ;
        RECT 40.560 135.475 40.785 137.595 ;
        RECT 40.955 137.265 41.285 137.765 ;
        RECT 41.455 137.095 41.625 137.595 ;
        RECT 40.960 136.925 41.625 137.095 ;
        RECT 40.960 135.935 41.190 136.925 ;
        RECT 41.360 136.105 41.710 136.755 ;
        RECT 41.890 136.625 42.225 137.595 ;
        RECT 42.395 136.625 42.565 137.765 ;
        RECT 42.735 137.425 44.765 137.595 ;
        RECT 41.890 135.955 42.060 136.625 ;
        RECT 42.735 136.455 42.905 137.425 ;
        RECT 42.230 136.125 42.485 136.455 ;
        RECT 42.710 136.125 42.905 136.455 ;
        RECT 43.075 137.085 44.200 137.255 ;
        RECT 42.315 135.955 42.485 136.125 ;
        RECT 43.075 135.955 43.245 137.085 ;
        RECT 40.960 135.765 41.625 135.935 ;
        RECT 40.955 135.215 41.285 135.595 ;
        RECT 41.455 135.475 41.625 135.765 ;
        RECT 41.890 135.385 42.145 135.955 ;
        RECT 42.315 135.785 43.245 135.955 ;
        RECT 43.415 136.745 44.425 136.915 ;
        RECT 43.415 135.945 43.585 136.745 ;
        RECT 43.790 136.065 44.065 136.545 ;
        RECT 43.785 135.895 44.065 136.065 ;
        RECT 43.070 135.750 43.245 135.785 ;
        RECT 42.315 135.215 42.645 135.615 ;
        RECT 43.070 135.385 43.600 135.750 ;
        RECT 43.790 135.385 44.065 135.895 ;
        RECT 44.235 135.385 44.425 136.745 ;
        RECT 44.595 136.760 44.765 137.425 ;
        RECT 44.935 137.005 45.105 137.765 ;
        RECT 45.340 137.005 45.855 137.415 ;
        RECT 44.595 136.570 45.345 136.760 ;
        RECT 45.515 136.195 45.855 137.005 ;
        RECT 44.625 136.025 45.855 136.195 ;
        RECT 46.485 136.675 48.155 137.765 ;
        RECT 46.485 136.155 47.235 136.675 ;
        RECT 48.385 136.625 48.595 137.765 ;
        RECT 48.765 136.615 49.095 137.595 ;
        RECT 49.265 136.625 49.495 137.765 ;
        RECT 44.605 135.215 45.115 135.750 ;
        RECT 45.335 135.420 45.580 136.025 ;
        RECT 47.405 135.985 48.155 136.505 ;
        RECT 46.485 135.215 48.155 135.985 ;
        RECT 48.385 135.215 48.595 136.035 ;
        RECT 48.765 136.015 49.015 136.615 ;
        RECT 50.165 136.600 50.455 137.765 ;
        RECT 51.085 136.690 51.355 137.595 ;
        RECT 51.525 137.005 51.855 137.765 ;
        RECT 52.035 136.835 52.205 137.595 ;
        RECT 49.185 136.205 49.515 136.455 ;
        RECT 48.765 135.385 49.095 136.015 ;
        RECT 49.265 135.215 49.495 136.035 ;
        RECT 50.165 135.215 50.455 135.940 ;
        RECT 51.085 135.890 51.255 136.690 ;
        RECT 51.540 136.665 52.205 136.835 ;
        RECT 52.465 137.045 52.925 137.595 ;
        RECT 53.115 137.045 53.445 137.765 ;
        RECT 51.540 136.520 51.710 136.665 ;
        RECT 51.425 136.190 51.710 136.520 ;
        RECT 51.540 135.935 51.710 136.190 ;
        RECT 51.945 136.115 52.275 136.485 ;
        RECT 51.085 135.385 51.345 135.890 ;
        RECT 51.540 135.765 52.205 135.935 ;
        RECT 51.525 135.215 51.855 135.595 ;
        RECT 52.035 135.385 52.205 135.765 ;
        RECT 52.465 135.675 52.715 137.045 ;
        RECT 53.645 136.875 53.945 137.425 ;
        RECT 54.115 137.095 54.395 137.765 ;
        RECT 55.280 136.895 55.565 137.765 ;
        RECT 55.735 137.135 55.995 137.595 ;
        RECT 56.170 137.305 56.425 137.765 ;
        RECT 56.595 137.135 56.855 137.595 ;
        RECT 55.735 136.965 56.855 137.135 ;
        RECT 57.025 136.965 57.335 137.765 ;
        RECT 53.005 136.705 53.945 136.875 ;
        RECT 53.005 136.455 53.175 136.705 ;
        RECT 54.315 136.455 54.580 136.815 ;
        RECT 55.735 136.715 55.995 136.965 ;
        RECT 57.505 136.795 57.815 137.595 ;
        RECT 58.910 137.330 64.255 137.765 ;
        RECT 52.885 136.125 53.175 136.455 ;
        RECT 53.345 136.205 53.685 136.455 ;
        RECT 53.905 136.205 54.580 136.455 ;
        RECT 55.240 136.545 55.995 136.715 ;
        RECT 56.785 136.625 57.815 136.795 ;
        RECT 53.005 136.035 53.175 136.125 ;
        RECT 55.240 136.035 55.645 136.545 ;
        RECT 56.785 136.375 56.955 136.625 ;
        RECT 55.815 136.205 56.955 136.375 ;
        RECT 53.005 135.845 54.395 136.035 ;
        RECT 55.240 135.865 56.890 136.035 ;
        RECT 57.125 135.885 57.475 136.455 ;
        RECT 52.465 135.385 53.025 135.675 ;
        RECT 53.195 135.215 53.445 135.675 ;
        RECT 54.065 135.485 54.395 135.845 ;
        RECT 55.285 135.215 55.565 135.695 ;
        RECT 55.735 135.475 55.995 135.865 ;
        RECT 56.170 135.215 56.425 135.695 ;
        RECT 56.595 135.475 56.890 135.865 ;
        RECT 57.645 135.715 57.815 136.625 ;
        RECT 60.500 136.080 60.850 137.330 ;
        RECT 64.425 136.625 64.765 137.595 ;
        RECT 64.935 136.625 65.105 137.765 ;
        RECT 65.375 136.965 65.625 137.765 ;
        RECT 66.270 136.795 66.600 137.595 ;
        RECT 66.900 136.965 67.230 137.765 ;
        RECT 67.400 136.795 67.730 137.595 ;
        RECT 65.295 136.625 67.730 136.795 ;
        RECT 69.025 136.675 72.535 137.765 ;
        RECT 72.710 137.340 73.045 137.765 ;
        RECT 73.215 137.160 73.400 137.565 ;
        RECT 72.735 136.985 73.400 137.160 ;
        RECT 73.605 136.985 73.935 137.765 ;
        RECT 62.330 135.760 62.670 136.590 ;
        RECT 64.425 136.575 64.655 136.625 ;
        RECT 64.425 136.015 64.600 136.575 ;
        RECT 65.295 136.375 65.465 136.625 ;
        RECT 64.770 136.205 65.465 136.375 ;
        RECT 65.640 136.205 66.060 136.405 ;
        RECT 66.230 136.205 66.560 136.405 ;
        RECT 66.730 136.205 67.060 136.405 ;
        RECT 57.070 135.215 57.345 135.695 ;
        RECT 57.515 135.385 57.815 135.715 ;
        RECT 58.910 135.215 64.255 135.760 ;
        RECT 64.425 135.385 64.765 136.015 ;
        RECT 64.935 135.215 65.185 136.015 ;
        RECT 65.375 135.865 66.600 136.035 ;
        RECT 65.375 135.385 65.705 135.865 ;
        RECT 65.875 135.215 66.100 135.675 ;
        RECT 66.270 135.385 66.600 135.865 ;
        RECT 67.230 135.995 67.400 136.625 ;
        RECT 67.585 136.205 67.935 136.455 ;
        RECT 69.025 136.155 70.715 136.675 ;
        RECT 67.230 135.385 67.730 135.995 ;
        RECT 70.885 135.985 72.535 136.505 ;
        RECT 69.025 135.215 72.535 135.985 ;
        RECT 72.735 135.955 73.075 136.985 ;
        RECT 74.105 136.795 74.375 137.565 ;
        RECT 73.245 136.625 74.375 136.795 ;
        RECT 73.245 136.125 73.495 136.625 ;
        RECT 72.735 135.785 73.420 135.955 ;
        RECT 73.675 135.875 74.035 136.455 ;
        RECT 72.710 135.215 73.045 135.615 ;
        RECT 73.215 135.385 73.420 135.785 ;
        RECT 74.205 135.715 74.375 136.625 ;
        RECT 74.545 136.675 75.755 137.765 ;
        RECT 74.545 136.135 75.065 136.675 ;
        RECT 75.925 136.600 76.215 137.765 ;
        RECT 76.385 136.675 78.055 137.765 ;
        RECT 78.425 137.095 78.705 137.765 ;
        RECT 78.875 136.875 79.175 137.425 ;
        RECT 79.375 137.045 79.705 137.765 ;
        RECT 79.895 137.045 80.355 137.595 ;
        RECT 75.235 135.965 75.755 136.505 ;
        RECT 76.385 136.155 77.135 136.675 ;
        RECT 77.305 135.985 78.055 136.505 ;
        RECT 78.240 136.455 78.505 136.815 ;
        RECT 78.875 136.705 79.815 136.875 ;
        RECT 79.645 136.455 79.815 136.705 ;
        RECT 78.240 136.205 78.915 136.455 ;
        RECT 79.135 136.205 79.475 136.455 ;
        RECT 79.645 136.125 79.935 136.455 ;
        RECT 79.645 136.035 79.815 136.125 ;
        RECT 73.630 135.215 73.905 135.695 ;
        RECT 74.115 135.385 74.375 135.715 ;
        RECT 74.545 135.215 75.755 135.965 ;
        RECT 75.925 135.215 76.215 135.940 ;
        RECT 76.385 135.215 78.055 135.985 ;
        RECT 78.425 135.845 79.815 136.035 ;
        RECT 78.425 135.485 78.755 135.845 ;
        RECT 80.105 135.675 80.355 137.045 ;
        RECT 79.375 135.215 79.625 135.675 ;
        RECT 79.795 135.385 80.355 135.675 ;
        RECT 80.525 137.045 80.985 137.595 ;
        RECT 81.175 137.045 81.505 137.765 ;
        RECT 80.525 135.675 80.775 137.045 ;
        RECT 81.705 136.875 82.005 137.425 ;
        RECT 82.175 137.095 82.455 137.765 ;
        RECT 81.065 136.705 82.005 136.875 ;
        RECT 82.825 137.045 83.285 137.595 ;
        RECT 83.475 137.045 83.805 137.765 ;
        RECT 81.065 136.455 81.235 136.705 ;
        RECT 82.375 136.455 82.640 136.815 ;
        RECT 80.945 136.125 81.235 136.455 ;
        RECT 81.405 136.205 81.745 136.455 ;
        RECT 81.965 136.205 82.640 136.455 ;
        RECT 81.065 136.035 81.235 136.125 ;
        RECT 81.065 135.845 82.455 136.035 ;
        RECT 80.525 135.385 81.085 135.675 ;
        RECT 81.255 135.215 81.505 135.675 ;
        RECT 82.125 135.485 82.455 135.845 ;
        RECT 82.825 135.675 83.075 137.045 ;
        RECT 84.005 136.875 84.305 137.425 ;
        RECT 84.475 137.095 84.755 137.765 ;
        RECT 83.365 136.705 84.305 136.875 ;
        RECT 85.215 136.835 85.385 137.595 ;
        RECT 85.565 137.005 85.895 137.765 ;
        RECT 83.365 136.455 83.535 136.705 ;
        RECT 84.675 136.455 84.940 136.815 ;
        RECT 85.215 136.665 85.880 136.835 ;
        RECT 86.065 136.690 86.335 137.595 ;
        RECT 85.710 136.520 85.880 136.665 ;
        RECT 83.245 136.125 83.535 136.455 ;
        RECT 83.705 136.205 84.045 136.455 ;
        RECT 84.265 136.205 84.940 136.455 ;
        RECT 83.365 136.035 83.535 136.125 ;
        RECT 85.145 136.115 85.475 136.485 ;
        RECT 85.710 136.190 85.995 136.520 ;
        RECT 83.365 135.845 84.755 136.035 ;
        RECT 85.710 135.935 85.880 136.190 ;
        RECT 82.825 135.385 83.385 135.675 ;
        RECT 83.555 135.215 83.805 135.675 ;
        RECT 84.425 135.485 84.755 135.845 ;
        RECT 85.215 135.765 85.880 135.935 ;
        RECT 86.165 135.890 86.335 136.690 ;
        RECT 86.965 136.675 90.475 137.765 ;
        RECT 86.965 136.155 88.655 136.675 ;
        RECT 90.685 136.625 90.915 137.765 ;
        RECT 91.085 136.615 91.415 137.595 ;
        RECT 91.585 136.625 91.795 137.765 ;
        RECT 92.115 136.835 92.285 137.595 ;
        RECT 92.465 137.005 92.795 137.765 ;
        RECT 92.115 136.665 92.780 136.835 ;
        RECT 92.965 136.690 93.235 137.595 ;
        RECT 88.825 135.985 90.475 136.505 ;
        RECT 90.665 136.205 90.995 136.455 ;
        RECT 85.215 135.385 85.385 135.765 ;
        RECT 85.565 135.215 85.895 135.595 ;
        RECT 86.075 135.385 86.335 135.890 ;
        RECT 86.965 135.215 90.475 135.985 ;
        RECT 90.685 135.215 90.915 136.035 ;
        RECT 91.165 136.015 91.415 136.615 ;
        RECT 92.610 136.520 92.780 136.665 ;
        RECT 92.045 136.115 92.375 136.485 ;
        RECT 92.610 136.190 92.895 136.520 ;
        RECT 91.085 135.385 91.415 136.015 ;
        RECT 91.585 135.215 91.795 136.035 ;
        RECT 92.610 135.935 92.780 136.190 ;
        RECT 92.115 135.765 92.780 135.935 ;
        RECT 93.065 135.890 93.235 136.690 ;
        RECT 94.325 137.005 94.840 137.415 ;
        RECT 95.075 137.005 95.245 137.765 ;
        RECT 95.415 137.425 97.445 137.595 ;
        RECT 94.325 136.195 94.665 137.005 ;
        RECT 95.415 136.760 95.585 137.425 ;
        RECT 95.980 137.085 97.105 137.255 ;
        RECT 94.835 136.570 95.585 136.760 ;
        RECT 95.755 136.745 96.765 136.915 ;
        RECT 94.325 136.025 95.555 136.195 ;
        RECT 92.115 135.385 92.285 135.765 ;
        RECT 92.465 135.215 92.795 135.595 ;
        RECT 92.975 135.385 93.235 135.890 ;
        RECT 94.600 135.420 94.845 136.025 ;
        RECT 95.065 135.215 95.575 135.750 ;
        RECT 95.755 135.385 95.945 136.745 ;
        RECT 96.115 136.065 96.390 136.545 ;
        RECT 96.115 135.895 96.395 136.065 ;
        RECT 96.595 135.945 96.765 136.745 ;
        RECT 96.935 135.955 97.105 137.085 ;
        RECT 97.275 136.455 97.445 137.425 ;
        RECT 97.615 136.625 97.785 137.765 ;
        RECT 97.955 136.625 98.290 137.595 ;
        RECT 97.275 136.125 97.470 136.455 ;
        RECT 97.695 136.125 97.950 136.455 ;
        RECT 97.695 135.955 97.865 136.125 ;
        RECT 98.120 135.955 98.290 136.625 ;
        RECT 96.115 135.385 96.390 135.895 ;
        RECT 96.935 135.785 97.865 135.955 ;
        RECT 96.935 135.750 97.110 135.785 ;
        RECT 96.580 135.385 97.110 135.750 ;
        RECT 97.535 135.215 97.865 135.615 ;
        RECT 98.035 135.385 98.290 135.955 ;
        RECT 98.465 136.625 98.735 137.595 ;
        RECT 98.945 136.965 99.225 137.765 ;
        RECT 99.395 137.255 101.050 137.545 ;
        RECT 99.460 136.915 101.050 137.085 ;
        RECT 99.460 136.795 99.630 136.915 ;
        RECT 98.905 136.625 99.630 136.795 ;
        RECT 98.465 135.890 98.635 136.625 ;
        RECT 98.905 136.455 99.075 136.625 ;
        RECT 98.805 136.125 99.075 136.455 ;
        RECT 99.245 136.125 99.650 136.455 ;
        RECT 99.820 136.125 100.530 136.745 ;
        RECT 100.730 136.625 101.050 136.915 ;
        RECT 101.685 136.600 101.975 137.765 ;
        RECT 102.145 136.675 104.735 137.765 ;
        RECT 98.905 135.955 99.075 136.125 ;
        RECT 98.465 135.545 98.735 135.890 ;
        RECT 98.905 135.785 100.515 135.955 ;
        RECT 100.700 135.885 101.050 136.455 ;
        RECT 102.145 136.155 103.355 136.675 ;
        RECT 104.905 136.625 105.175 137.595 ;
        RECT 105.385 136.965 105.665 137.765 ;
        RECT 105.835 137.255 107.490 137.545 ;
        RECT 105.900 136.915 107.490 137.085 ;
        RECT 105.900 136.795 106.070 136.915 ;
        RECT 105.345 136.625 106.070 136.795 ;
        RECT 103.525 135.985 104.735 136.505 ;
        RECT 98.925 135.215 99.305 135.615 ;
        RECT 99.475 135.435 99.645 135.785 ;
        RECT 99.815 135.215 100.145 135.615 ;
        RECT 100.345 135.435 100.515 135.785 ;
        RECT 100.715 135.215 101.045 135.715 ;
        RECT 101.685 135.215 101.975 135.940 ;
        RECT 102.145 135.215 104.735 135.985 ;
        RECT 104.905 135.890 105.075 136.625 ;
        RECT 105.345 136.455 105.515 136.625 ;
        RECT 106.260 136.575 106.975 136.745 ;
        RECT 107.170 136.625 107.490 136.915 ;
        RECT 107.665 136.625 108.005 137.595 ;
        RECT 108.175 136.625 108.345 137.765 ;
        RECT 108.615 136.965 108.865 137.765 ;
        RECT 109.510 136.795 109.840 137.595 ;
        RECT 110.140 136.965 110.470 137.765 ;
        RECT 110.640 136.795 110.970 137.595 ;
        RECT 108.535 136.625 110.970 136.795 ;
        RECT 111.345 136.625 111.615 137.595 ;
        RECT 111.825 136.965 112.105 137.765 ;
        RECT 112.275 137.255 113.930 137.545 ;
        RECT 114.110 137.330 119.455 137.765 ;
        RECT 112.340 136.915 113.930 137.085 ;
        RECT 112.340 136.795 112.510 136.915 ;
        RECT 111.785 136.625 112.510 136.795 ;
        RECT 105.245 136.125 105.515 136.455 ;
        RECT 105.685 136.125 106.090 136.455 ;
        RECT 106.260 136.125 106.970 136.575 ;
        RECT 105.345 135.955 105.515 136.125 ;
        RECT 104.905 135.545 105.175 135.890 ;
        RECT 105.345 135.785 106.955 135.955 ;
        RECT 107.140 135.885 107.490 136.455 ;
        RECT 107.665 136.065 107.840 136.625 ;
        RECT 108.535 136.375 108.705 136.625 ;
        RECT 108.010 136.205 108.705 136.375 ;
        RECT 108.880 136.205 109.300 136.405 ;
        RECT 109.470 136.205 109.800 136.405 ;
        RECT 109.970 136.205 110.300 136.405 ;
        RECT 107.665 136.015 107.895 136.065 ;
        RECT 105.365 135.215 105.745 135.615 ;
        RECT 105.915 135.435 106.085 135.785 ;
        RECT 106.255 135.215 106.585 135.615 ;
        RECT 106.785 135.435 106.955 135.785 ;
        RECT 107.155 135.215 107.485 135.715 ;
        RECT 107.665 135.385 108.005 136.015 ;
        RECT 108.175 135.215 108.425 136.015 ;
        RECT 108.615 135.865 109.840 136.035 ;
        RECT 108.615 135.385 108.945 135.865 ;
        RECT 109.115 135.215 109.340 135.675 ;
        RECT 109.510 135.385 109.840 135.865 ;
        RECT 110.470 135.995 110.640 136.625 ;
        RECT 110.825 136.205 111.175 136.455 ;
        RECT 110.470 135.385 110.970 135.995 ;
        RECT 111.345 135.890 111.515 136.625 ;
        RECT 111.785 136.455 111.955 136.625 ;
        RECT 112.700 136.575 113.415 136.745 ;
        RECT 113.610 136.625 113.930 136.915 ;
        RECT 111.685 136.125 111.955 136.455 ;
        RECT 112.125 136.125 112.530 136.455 ;
        RECT 112.700 136.125 113.410 136.575 ;
        RECT 111.785 135.955 111.955 136.125 ;
        RECT 111.345 135.545 111.615 135.890 ;
        RECT 111.785 135.785 113.395 135.955 ;
        RECT 113.580 135.885 113.930 136.455 ;
        RECT 115.700 136.080 116.050 137.330 ;
        RECT 119.715 136.835 119.885 137.595 ;
        RECT 120.065 137.005 120.395 137.765 ;
        RECT 119.715 136.665 120.380 136.835 ;
        RECT 120.565 136.690 120.835 137.595 ;
        RECT 111.805 135.215 112.185 135.615 ;
        RECT 112.355 135.435 112.525 135.785 ;
        RECT 112.695 135.215 113.025 135.615 ;
        RECT 113.225 135.435 113.395 135.785 ;
        RECT 117.530 135.760 117.870 136.590 ;
        RECT 120.210 136.520 120.380 136.665 ;
        RECT 119.645 136.115 119.975 136.485 ;
        RECT 120.210 136.190 120.495 136.520 ;
        RECT 120.210 135.935 120.380 136.190 ;
        RECT 119.715 135.765 120.380 135.935 ;
        RECT 120.665 135.890 120.835 136.690 ;
        RECT 122.015 136.835 122.185 137.595 ;
        RECT 122.365 137.005 122.695 137.765 ;
        RECT 122.015 136.665 122.680 136.835 ;
        RECT 122.865 136.690 123.135 137.595 ;
        RECT 122.510 136.520 122.680 136.665 ;
        RECT 121.945 136.115 122.275 136.485 ;
        RECT 122.510 136.190 122.795 136.520 ;
        RECT 122.510 135.935 122.680 136.190 ;
        RECT 113.595 135.215 113.925 135.715 ;
        RECT 114.110 135.215 119.455 135.760 ;
        RECT 119.715 135.385 119.885 135.765 ;
        RECT 120.065 135.215 120.395 135.595 ;
        RECT 120.575 135.385 120.835 135.890 ;
        RECT 122.015 135.765 122.680 135.935 ;
        RECT 122.965 135.890 123.135 136.690 ;
        RECT 123.765 136.675 126.355 137.765 ;
        RECT 126.525 136.675 127.735 137.765 ;
        RECT 123.765 136.155 124.975 136.675 ;
        RECT 125.145 135.985 126.355 136.505 ;
        RECT 126.525 136.135 127.045 136.675 ;
        RECT 122.015 135.385 122.185 135.765 ;
        RECT 122.365 135.215 122.695 135.595 ;
        RECT 122.875 135.385 123.135 135.890 ;
        RECT 123.765 135.215 126.355 135.985 ;
        RECT 127.215 135.965 127.735 136.505 ;
        RECT 126.525 135.215 127.735 135.965 ;
        RECT 20.640 135.045 127.820 135.215 ;
        RECT 20.725 134.295 21.935 135.045 ;
        RECT 22.480 134.705 22.735 134.865 ;
        RECT 22.395 134.535 22.735 134.705 ;
        RECT 22.915 134.585 23.200 135.045 ;
        RECT 22.480 134.335 22.735 134.535 ;
        RECT 20.725 133.755 21.245 134.295 ;
        RECT 21.415 133.585 21.935 134.125 ;
        RECT 20.725 132.495 21.935 133.585 ;
        RECT 22.480 133.475 22.660 134.335 ;
        RECT 23.380 134.135 23.630 134.785 ;
        RECT 22.830 133.805 23.630 134.135 ;
        RECT 22.480 132.805 22.735 133.475 ;
        RECT 22.915 132.495 23.200 133.295 ;
        RECT 23.380 133.215 23.630 133.805 ;
        RECT 23.830 134.450 24.150 134.780 ;
        RECT 24.330 134.565 24.990 135.045 ;
        RECT 25.190 134.655 26.040 134.825 ;
        RECT 23.830 133.555 24.020 134.450 ;
        RECT 24.340 134.125 25.000 134.395 ;
        RECT 24.670 134.065 25.000 134.125 ;
        RECT 24.190 133.895 24.520 133.955 ;
        RECT 25.190 133.895 25.360 134.655 ;
        RECT 26.600 134.585 26.920 135.045 ;
        RECT 27.120 134.405 27.370 134.835 ;
        RECT 27.660 134.605 28.070 135.045 ;
        RECT 28.240 134.665 29.255 134.865 ;
        RECT 25.530 134.235 26.780 134.405 ;
        RECT 25.530 134.115 25.860 134.235 ;
        RECT 24.190 133.725 26.090 133.895 ;
        RECT 23.830 133.385 25.750 133.555 ;
        RECT 23.830 133.365 24.150 133.385 ;
        RECT 23.380 132.705 23.710 133.215 ;
        RECT 23.980 132.755 24.150 133.365 ;
        RECT 25.920 133.215 26.090 133.725 ;
        RECT 26.260 133.655 26.440 134.065 ;
        RECT 26.610 133.475 26.780 134.235 ;
        RECT 24.320 132.495 24.650 133.185 ;
        RECT 24.880 133.045 26.090 133.215 ;
        RECT 26.260 133.165 26.780 133.475 ;
        RECT 26.950 134.065 27.370 134.405 ;
        RECT 27.660 134.065 28.070 134.395 ;
        RECT 26.950 133.295 27.140 134.065 ;
        RECT 28.240 133.935 28.410 134.665 ;
        RECT 29.555 134.495 29.725 134.825 ;
        RECT 29.895 134.665 30.225 135.045 ;
        RECT 28.580 134.115 28.930 134.485 ;
        RECT 28.240 133.895 28.660 133.935 ;
        RECT 27.310 133.725 28.660 133.895 ;
        RECT 27.310 133.565 27.560 133.725 ;
        RECT 28.070 133.295 28.320 133.555 ;
        RECT 26.950 133.045 28.320 133.295 ;
        RECT 24.880 132.755 25.120 133.045 ;
        RECT 25.920 132.965 26.090 133.045 ;
        RECT 25.320 132.495 25.740 132.875 ;
        RECT 25.920 132.715 26.550 132.965 ;
        RECT 27.020 132.495 27.350 132.875 ;
        RECT 27.520 132.755 27.690 133.045 ;
        RECT 28.490 132.880 28.660 133.725 ;
        RECT 29.110 133.555 29.330 134.425 ;
        RECT 29.555 134.305 30.250 134.495 ;
        RECT 28.830 133.175 29.330 133.555 ;
        RECT 29.500 133.505 29.910 134.125 ;
        RECT 30.080 133.335 30.250 134.305 ;
        RECT 29.555 133.165 30.250 133.335 ;
        RECT 27.870 132.495 28.250 132.875 ;
        RECT 28.490 132.710 29.320 132.880 ;
        RECT 29.555 132.665 29.725 133.165 ;
        RECT 29.895 132.495 30.225 132.995 ;
        RECT 30.440 132.665 30.665 134.785 ;
        RECT 30.835 134.665 31.165 135.045 ;
        RECT 31.335 134.495 31.505 134.785 ;
        RECT 30.840 134.325 31.505 134.495 ;
        RECT 31.765 134.370 32.025 134.875 ;
        RECT 32.205 134.665 32.535 135.045 ;
        RECT 32.715 134.495 32.885 134.875 ;
        RECT 30.840 133.335 31.070 134.325 ;
        RECT 31.240 133.505 31.590 134.155 ;
        RECT 31.765 133.570 31.935 134.370 ;
        RECT 32.220 134.325 32.885 134.495 ;
        RECT 32.220 134.070 32.390 134.325 ;
        RECT 33.145 134.295 34.355 135.045 ;
        RECT 32.105 133.740 32.390 134.070 ;
        RECT 32.625 133.775 32.955 134.145 ;
        RECT 32.220 133.595 32.390 133.740 ;
        RECT 30.840 133.165 31.505 133.335 ;
        RECT 30.835 132.495 31.165 132.995 ;
        RECT 31.335 132.665 31.505 133.165 ;
        RECT 31.765 132.665 32.035 133.570 ;
        RECT 32.220 133.425 32.885 133.595 ;
        RECT 32.205 132.495 32.535 133.255 ;
        RECT 32.715 132.665 32.885 133.425 ;
        RECT 33.145 133.585 33.665 134.125 ;
        RECT 33.835 133.755 34.355 134.295 ;
        RECT 34.525 134.370 34.795 134.715 ;
        RECT 34.985 134.645 35.365 135.045 ;
        RECT 35.535 134.475 35.705 134.825 ;
        RECT 35.875 134.645 36.205 135.045 ;
        RECT 36.405 134.475 36.575 134.825 ;
        RECT 36.775 134.545 37.105 135.045 ;
        RECT 34.525 133.635 34.695 134.370 ;
        RECT 34.965 134.305 36.575 134.475 ;
        RECT 34.965 134.135 35.135 134.305 ;
        RECT 34.865 133.805 35.135 134.135 ;
        RECT 35.305 133.805 35.710 134.135 ;
        RECT 34.965 133.635 35.135 133.805 ;
        RECT 35.880 133.685 36.590 134.135 ;
        RECT 36.760 133.805 37.110 134.375 ;
        RECT 37.285 134.320 37.575 135.045 ;
        RECT 37.750 134.575 38.080 135.045 ;
        RECT 38.250 134.405 38.475 134.850 ;
        RECT 38.645 134.520 38.940 135.045 ;
        RECT 37.745 134.235 38.475 134.405 ;
        RECT 39.585 134.370 39.855 134.715 ;
        RECT 40.045 134.645 40.425 135.045 ;
        RECT 40.595 134.475 40.765 134.825 ;
        RECT 40.935 134.645 41.265 135.045 ;
        RECT 41.465 134.475 41.635 134.825 ;
        RECT 41.835 134.545 42.165 135.045 ;
        RECT 43.265 134.535 43.570 135.045 ;
        RECT 33.145 132.495 34.355 133.585 ;
        RECT 34.525 132.665 34.795 133.635 ;
        RECT 34.965 133.465 35.690 133.635 ;
        RECT 35.880 133.515 36.595 133.685 ;
        RECT 37.745 133.670 38.025 134.235 ;
        RECT 38.195 133.840 39.415 134.065 ;
        RECT 35.520 133.345 35.690 133.465 ;
        RECT 36.790 133.345 37.110 133.635 ;
        RECT 35.005 132.495 35.285 133.295 ;
        RECT 35.520 133.175 37.110 133.345 ;
        RECT 35.455 132.715 37.110 133.005 ;
        RECT 37.285 132.495 37.575 133.660 ;
        RECT 37.745 133.500 39.345 133.670 ;
        RECT 37.805 132.495 38.060 133.330 ;
        RECT 38.230 132.695 38.490 133.500 ;
        RECT 38.660 132.495 38.920 133.330 ;
        RECT 39.090 132.695 39.345 133.500 ;
        RECT 39.585 133.635 39.755 134.370 ;
        RECT 40.025 134.305 41.635 134.475 ;
        RECT 40.025 134.135 40.195 134.305 ;
        RECT 39.925 133.805 40.195 134.135 ;
        RECT 40.365 133.805 40.770 134.135 ;
        RECT 40.025 133.635 40.195 133.805 ;
        RECT 39.585 132.665 39.855 133.635 ;
        RECT 40.025 133.465 40.750 133.635 ;
        RECT 40.940 133.515 41.650 134.135 ;
        RECT 41.820 133.805 42.170 134.375 ;
        RECT 43.265 133.805 43.580 134.365 ;
        RECT 43.750 134.055 44.000 134.865 ;
        RECT 44.170 134.520 44.430 135.045 ;
        RECT 44.610 134.055 44.860 134.865 ;
        RECT 45.030 134.485 45.290 135.045 ;
        RECT 45.460 134.395 45.720 134.850 ;
        RECT 45.890 134.565 46.150 135.045 ;
        RECT 46.320 134.395 46.580 134.850 ;
        RECT 46.750 134.565 47.010 135.045 ;
        RECT 47.180 134.395 47.440 134.850 ;
        RECT 47.610 134.565 47.855 135.045 ;
        RECT 48.025 134.395 48.300 134.850 ;
        RECT 48.470 134.565 48.715 135.045 ;
        RECT 48.885 134.395 49.145 134.850 ;
        RECT 49.325 134.565 49.575 135.045 ;
        RECT 49.745 134.395 50.005 134.850 ;
        RECT 50.185 134.565 50.435 135.045 ;
        RECT 50.605 134.395 50.865 134.850 ;
        RECT 51.045 134.565 51.305 135.045 ;
        RECT 51.475 134.395 51.735 134.850 ;
        RECT 51.905 134.565 52.205 135.045 ;
        RECT 45.460 134.225 52.205 134.395 ;
        RECT 43.750 133.805 50.870 134.055 ;
        RECT 40.580 133.345 40.750 133.465 ;
        RECT 41.850 133.345 42.170 133.635 ;
        RECT 40.065 132.495 40.345 133.295 ;
        RECT 40.580 133.175 42.170 133.345 ;
        RECT 40.515 132.715 42.170 133.005 ;
        RECT 43.275 132.495 43.570 133.305 ;
        RECT 43.750 132.665 43.995 133.805 ;
        RECT 44.170 132.495 44.430 133.305 ;
        RECT 44.610 132.670 44.860 133.805 ;
        RECT 51.040 133.635 52.205 134.225 ;
        RECT 45.460 133.410 52.205 133.635 ;
        RECT 52.470 134.305 52.725 134.875 ;
        RECT 52.895 134.645 53.225 135.045 ;
        RECT 53.650 134.510 54.180 134.875 ;
        RECT 53.650 134.475 53.825 134.510 ;
        RECT 52.895 134.305 53.825 134.475 ;
        RECT 52.470 133.635 52.640 134.305 ;
        RECT 52.895 134.135 53.065 134.305 ;
        RECT 52.810 133.805 53.065 134.135 ;
        RECT 53.290 133.805 53.485 134.135 ;
        RECT 45.460 133.395 50.865 133.410 ;
        RECT 45.030 132.500 45.290 133.295 ;
        RECT 45.460 132.670 45.720 133.395 ;
        RECT 45.890 132.500 46.150 133.225 ;
        RECT 46.320 132.670 46.580 133.395 ;
        RECT 46.750 132.500 47.010 133.225 ;
        RECT 47.180 132.670 47.440 133.395 ;
        RECT 47.610 132.500 47.870 133.225 ;
        RECT 48.040 132.670 48.300 133.395 ;
        RECT 48.470 132.500 48.715 133.225 ;
        RECT 48.885 132.670 49.145 133.395 ;
        RECT 49.330 132.500 49.575 133.225 ;
        RECT 49.745 132.670 50.005 133.395 ;
        RECT 50.190 132.500 50.435 133.225 ;
        RECT 50.605 132.670 50.865 133.395 ;
        RECT 51.050 132.500 51.305 133.225 ;
        RECT 51.475 132.670 51.765 133.410 ;
        RECT 45.030 132.495 51.305 132.500 ;
        RECT 51.935 132.495 52.205 133.240 ;
        RECT 52.470 132.665 52.805 133.635 ;
        RECT 52.975 132.495 53.145 133.635 ;
        RECT 53.315 132.835 53.485 133.805 ;
        RECT 53.655 133.175 53.825 134.305 ;
        RECT 53.995 133.515 54.165 134.315 ;
        RECT 54.370 134.025 54.645 134.875 ;
        RECT 54.365 133.855 54.645 134.025 ;
        RECT 54.370 133.715 54.645 133.855 ;
        RECT 54.815 133.515 55.005 134.875 ;
        RECT 55.185 134.510 55.695 135.045 ;
        RECT 55.915 134.235 56.160 134.840 ;
        RECT 56.605 134.370 56.865 134.875 ;
        RECT 57.045 134.665 57.375 135.045 ;
        RECT 57.555 134.495 57.725 134.875 ;
        RECT 55.205 134.065 56.435 134.235 ;
        RECT 53.995 133.345 55.005 133.515 ;
        RECT 55.175 133.500 55.925 133.690 ;
        RECT 53.655 133.005 54.780 133.175 ;
        RECT 55.175 132.835 55.345 133.500 ;
        RECT 56.095 133.255 56.435 134.065 ;
        RECT 53.315 132.665 55.345 132.835 ;
        RECT 55.515 132.495 55.685 133.255 ;
        RECT 55.920 132.845 56.435 133.255 ;
        RECT 56.605 133.570 56.775 134.370 ;
        RECT 57.060 134.325 57.725 134.495 ;
        RECT 57.060 134.070 57.230 134.325 ;
        RECT 59.180 134.235 59.425 134.840 ;
        RECT 59.645 134.510 60.155 135.045 ;
        RECT 56.945 133.740 57.230 134.070 ;
        RECT 57.465 133.775 57.795 134.145 ;
        RECT 58.905 134.065 60.135 134.235 ;
        RECT 57.060 133.595 57.230 133.740 ;
        RECT 56.605 132.665 56.875 133.570 ;
        RECT 57.060 133.425 57.725 133.595 ;
        RECT 57.045 132.495 57.375 133.255 ;
        RECT 57.555 132.665 57.725 133.425 ;
        RECT 58.905 133.255 59.245 134.065 ;
        RECT 59.415 133.500 60.165 133.690 ;
        RECT 58.905 132.845 59.420 133.255 ;
        RECT 59.655 132.495 59.825 133.255 ;
        RECT 59.995 132.835 60.165 133.500 ;
        RECT 60.335 133.515 60.525 134.875 ;
        RECT 60.695 134.025 60.970 134.875 ;
        RECT 61.160 134.510 61.690 134.875 ;
        RECT 62.115 134.645 62.445 135.045 ;
        RECT 61.515 134.475 61.690 134.510 ;
        RECT 60.695 133.855 60.975 134.025 ;
        RECT 60.695 133.715 60.970 133.855 ;
        RECT 61.175 133.515 61.345 134.315 ;
        RECT 60.335 133.345 61.345 133.515 ;
        RECT 61.515 134.305 62.445 134.475 ;
        RECT 62.615 134.305 62.870 134.875 ;
        RECT 63.045 134.320 63.335 135.045 ;
        RECT 61.515 133.175 61.685 134.305 ;
        RECT 62.275 134.135 62.445 134.305 ;
        RECT 60.560 133.005 61.685 133.175 ;
        RECT 61.855 133.805 62.050 134.135 ;
        RECT 62.275 133.805 62.530 134.135 ;
        RECT 61.855 132.835 62.025 133.805 ;
        RECT 62.700 133.635 62.870 134.305 ;
        RECT 63.505 134.295 64.715 135.045 ;
        RECT 59.995 132.665 62.025 132.835 ;
        RECT 62.195 132.495 62.365 133.635 ;
        RECT 62.535 132.665 62.870 133.635 ;
        RECT 63.045 132.495 63.335 133.660 ;
        RECT 63.505 133.585 64.025 134.125 ;
        RECT 64.195 133.755 64.715 134.295 ;
        RECT 64.885 134.245 65.225 134.875 ;
        RECT 65.395 134.245 65.645 135.045 ;
        RECT 65.835 134.395 66.165 134.875 ;
        RECT 66.335 134.585 66.560 135.045 ;
        RECT 66.730 134.395 67.060 134.875 ;
        RECT 64.885 134.195 65.115 134.245 ;
        RECT 65.835 134.225 67.060 134.395 ;
        RECT 67.690 134.265 68.190 134.875 ;
        RECT 68.565 134.275 71.155 135.045 ;
        RECT 71.330 134.645 71.665 135.045 ;
        RECT 71.835 134.475 72.040 134.875 ;
        RECT 72.250 134.565 72.525 135.045 ;
        RECT 72.735 134.545 72.995 134.875 ;
        RECT 64.885 133.635 65.060 134.195 ;
        RECT 65.230 133.885 65.925 134.055 ;
        RECT 65.755 133.635 65.925 133.885 ;
        RECT 66.100 133.855 66.520 134.055 ;
        RECT 66.690 133.855 67.020 134.055 ;
        RECT 67.190 133.855 67.520 134.055 ;
        RECT 67.690 133.635 67.860 134.265 ;
        RECT 68.045 133.805 68.395 134.055 ;
        RECT 63.505 132.495 64.715 133.585 ;
        RECT 64.885 132.665 65.225 133.635 ;
        RECT 65.395 132.495 65.565 133.635 ;
        RECT 65.755 133.465 68.190 133.635 ;
        RECT 65.835 132.495 66.085 133.295 ;
        RECT 66.730 132.665 67.060 133.465 ;
        RECT 67.360 132.495 67.690 133.295 ;
        RECT 67.860 132.665 68.190 133.465 ;
        RECT 68.565 133.585 69.775 134.105 ;
        RECT 69.945 133.755 71.155 134.275 ;
        RECT 71.355 134.305 72.040 134.475 ;
        RECT 68.565 132.495 71.155 133.585 ;
        RECT 71.355 133.275 71.695 134.305 ;
        RECT 71.865 133.635 72.115 134.135 ;
        RECT 72.295 133.805 72.655 134.385 ;
        RECT 72.825 133.635 72.995 134.545 ;
        RECT 71.865 133.465 72.995 133.635 ;
        RECT 71.355 133.100 72.020 133.275 ;
        RECT 71.330 132.495 71.665 132.920 ;
        RECT 71.835 132.695 72.020 133.100 ;
        RECT 72.225 132.495 72.555 133.275 ;
        RECT 72.725 132.695 72.995 133.465 ;
        RECT 73.165 134.585 73.725 134.875 ;
        RECT 73.895 134.585 74.145 135.045 ;
        RECT 73.165 133.215 73.415 134.585 ;
        RECT 74.765 134.415 75.095 134.775 ;
        RECT 73.705 134.225 75.095 134.415 ;
        RECT 75.925 134.275 78.515 135.045 ;
        RECT 73.705 134.135 73.875 134.225 ;
        RECT 73.585 133.805 73.875 134.135 ;
        RECT 74.045 133.805 74.385 134.055 ;
        RECT 74.605 133.805 75.280 134.055 ;
        RECT 73.705 133.555 73.875 133.805 ;
        RECT 73.705 133.385 74.645 133.555 ;
        RECT 75.015 133.445 75.280 133.805 ;
        RECT 75.925 133.585 77.135 134.105 ;
        RECT 77.305 133.755 78.515 134.275 ;
        RECT 79.060 134.335 79.315 134.865 ;
        RECT 79.495 134.585 79.780 135.045 ;
        RECT 73.165 132.665 73.625 133.215 ;
        RECT 73.815 132.495 74.145 133.215 ;
        RECT 74.345 132.835 74.645 133.385 ;
        RECT 74.815 132.495 75.095 133.165 ;
        RECT 75.925 132.495 78.515 133.585 ;
        RECT 79.060 133.475 79.240 134.335 ;
        RECT 79.960 134.135 80.210 134.785 ;
        RECT 79.410 133.805 80.210 134.135 ;
        RECT 79.060 133.005 79.315 133.475 ;
        RECT 78.975 132.835 79.315 133.005 ;
        RECT 79.060 132.805 79.315 132.835 ;
        RECT 79.495 132.495 79.780 133.295 ;
        RECT 79.960 133.215 80.210 133.805 ;
        RECT 80.410 134.450 80.730 134.780 ;
        RECT 80.910 134.565 81.570 135.045 ;
        RECT 81.770 134.655 82.620 134.825 ;
        RECT 80.410 133.555 80.600 134.450 ;
        RECT 80.920 134.125 81.580 134.395 ;
        RECT 81.250 134.065 81.580 134.125 ;
        RECT 80.770 133.895 81.100 133.955 ;
        RECT 81.770 133.895 81.940 134.655 ;
        RECT 83.180 134.585 83.500 135.045 ;
        RECT 83.700 134.405 83.950 134.835 ;
        RECT 84.240 134.605 84.650 135.045 ;
        RECT 84.820 134.665 85.835 134.865 ;
        RECT 82.110 134.235 83.360 134.405 ;
        RECT 82.110 134.115 82.440 134.235 ;
        RECT 80.770 133.725 82.670 133.895 ;
        RECT 80.410 133.385 82.330 133.555 ;
        RECT 80.410 133.365 80.730 133.385 ;
        RECT 79.960 132.705 80.290 133.215 ;
        RECT 80.560 132.755 80.730 133.365 ;
        RECT 82.500 133.215 82.670 133.725 ;
        RECT 82.840 133.655 83.020 134.065 ;
        RECT 83.190 133.475 83.360 134.235 ;
        RECT 80.900 132.495 81.230 133.185 ;
        RECT 81.460 133.045 82.670 133.215 ;
        RECT 82.840 133.165 83.360 133.475 ;
        RECT 83.530 134.065 83.950 134.405 ;
        RECT 84.240 134.065 84.650 134.395 ;
        RECT 83.530 133.295 83.720 134.065 ;
        RECT 84.820 133.935 84.990 134.665 ;
        RECT 86.135 134.495 86.305 134.825 ;
        RECT 86.475 134.665 86.805 135.045 ;
        RECT 85.160 134.115 85.510 134.485 ;
        RECT 84.820 133.895 85.240 133.935 ;
        RECT 83.890 133.725 85.240 133.895 ;
        RECT 83.890 133.565 84.140 133.725 ;
        RECT 84.650 133.295 84.900 133.555 ;
        RECT 83.530 133.045 84.900 133.295 ;
        RECT 81.460 132.755 81.700 133.045 ;
        RECT 82.500 132.965 82.670 133.045 ;
        RECT 81.900 132.495 82.320 132.875 ;
        RECT 82.500 132.715 83.130 132.965 ;
        RECT 83.600 132.495 83.930 132.875 ;
        RECT 84.100 132.755 84.270 133.045 ;
        RECT 85.070 132.880 85.240 133.725 ;
        RECT 85.690 133.555 85.910 134.425 ;
        RECT 86.135 134.305 86.830 134.495 ;
        RECT 85.410 133.175 85.910 133.555 ;
        RECT 86.080 133.505 86.490 134.125 ;
        RECT 86.660 133.335 86.830 134.305 ;
        RECT 86.135 133.165 86.830 133.335 ;
        RECT 84.450 132.495 84.830 132.875 ;
        RECT 85.070 132.710 85.900 132.880 ;
        RECT 86.135 132.665 86.305 133.165 ;
        RECT 86.475 132.495 86.805 132.995 ;
        RECT 87.020 132.665 87.245 134.785 ;
        RECT 87.415 134.665 87.745 135.045 ;
        RECT 87.915 134.495 88.085 134.785 ;
        RECT 87.420 134.325 88.085 134.495 ;
        RECT 87.420 133.335 87.650 134.325 ;
        RECT 88.805 134.320 89.095 135.045 ;
        RECT 90.190 134.500 95.535 135.045 ;
        RECT 95.710 134.500 101.055 135.045 ;
        RECT 101.230 134.500 106.575 135.045 ;
        RECT 87.820 133.505 88.170 134.155 ;
        RECT 87.420 133.165 88.085 133.335 ;
        RECT 87.415 132.495 87.745 132.995 ;
        RECT 87.915 132.665 88.085 133.165 ;
        RECT 88.805 132.495 89.095 133.660 ;
        RECT 91.780 132.930 92.130 134.180 ;
        RECT 93.610 133.670 93.950 134.500 ;
        RECT 97.300 132.930 97.650 134.180 ;
        RECT 99.130 133.670 99.470 134.500 ;
        RECT 102.820 132.930 103.170 134.180 ;
        RECT 104.650 133.670 104.990 134.500 ;
        RECT 106.945 134.415 107.275 134.775 ;
        RECT 107.895 134.585 108.145 135.045 ;
        RECT 108.315 134.585 108.875 134.875 ;
        RECT 106.945 134.225 108.335 134.415 ;
        RECT 108.165 134.135 108.335 134.225 ;
        RECT 106.760 133.805 107.435 134.055 ;
        RECT 107.655 133.805 107.995 134.055 ;
        RECT 108.165 133.805 108.455 134.135 ;
        RECT 106.760 133.445 107.025 133.805 ;
        RECT 108.165 133.555 108.335 133.805 ;
        RECT 107.395 133.385 108.335 133.555 ;
        RECT 90.190 132.495 95.535 132.930 ;
        RECT 95.710 132.495 101.055 132.930 ;
        RECT 101.230 132.495 106.575 132.930 ;
        RECT 106.945 132.495 107.225 133.165 ;
        RECT 107.395 132.835 107.695 133.385 ;
        RECT 108.625 133.215 108.875 134.585 ;
        RECT 107.895 132.495 108.225 133.215 ;
        RECT 108.415 132.665 108.875 133.215 ;
        RECT 109.045 134.585 109.605 134.875 ;
        RECT 109.775 134.585 110.025 135.045 ;
        RECT 109.045 133.215 109.295 134.585 ;
        RECT 110.645 134.415 110.975 134.775 ;
        RECT 109.585 134.225 110.975 134.415 ;
        RECT 111.805 134.585 112.365 134.875 ;
        RECT 112.535 134.585 112.785 135.045 ;
        RECT 109.585 134.135 109.755 134.225 ;
        RECT 109.465 133.805 109.755 134.135 ;
        RECT 109.925 133.805 110.265 134.055 ;
        RECT 110.485 133.805 111.160 134.055 ;
        RECT 109.585 133.555 109.755 133.805 ;
        RECT 109.585 133.385 110.525 133.555 ;
        RECT 110.895 133.445 111.160 133.805 ;
        RECT 109.045 132.665 109.505 133.215 ;
        RECT 109.695 132.495 110.025 133.215 ;
        RECT 110.225 132.835 110.525 133.385 ;
        RECT 111.805 133.215 112.055 134.585 ;
        RECT 113.405 134.415 113.735 134.775 ;
        RECT 112.345 134.225 113.735 134.415 ;
        RECT 114.565 134.320 114.855 135.045 ;
        RECT 115.490 134.500 120.835 135.045 ;
        RECT 121.010 134.500 126.355 135.045 ;
        RECT 112.345 134.135 112.515 134.225 ;
        RECT 112.225 133.805 112.515 134.135 ;
        RECT 112.685 133.805 113.025 134.055 ;
        RECT 113.245 133.805 113.920 134.055 ;
        RECT 112.345 133.555 112.515 133.805 ;
        RECT 112.345 133.385 113.285 133.555 ;
        RECT 113.655 133.445 113.920 133.805 ;
        RECT 110.695 132.495 110.975 133.165 ;
        RECT 111.805 132.665 112.265 133.215 ;
        RECT 112.455 132.495 112.785 133.215 ;
        RECT 112.985 132.835 113.285 133.385 ;
        RECT 113.455 132.495 113.735 133.165 ;
        RECT 114.565 132.495 114.855 133.660 ;
        RECT 117.080 132.930 117.430 134.180 ;
        RECT 118.910 133.670 119.250 134.500 ;
        RECT 122.600 132.930 122.950 134.180 ;
        RECT 124.430 133.670 124.770 134.500 ;
        RECT 126.525 134.295 127.735 135.045 ;
        RECT 126.525 133.585 127.045 134.125 ;
        RECT 127.215 133.755 127.735 134.295 ;
        RECT 115.490 132.495 120.835 132.930 ;
        RECT 121.010 132.495 126.355 132.930 ;
        RECT 126.525 132.495 127.735 133.585 ;
        RECT 20.640 132.325 127.820 132.495 ;
        RECT 20.725 131.235 21.935 132.325 ;
        RECT 20.725 130.525 21.245 131.065 ;
        RECT 21.415 130.695 21.935 131.235 ;
        RECT 22.565 131.235 24.235 132.325 ;
        RECT 22.565 130.715 23.315 131.235 ;
        RECT 24.405 131.160 24.695 132.325 ;
        RECT 25.845 131.185 26.055 132.325 ;
        RECT 26.225 131.175 26.555 132.155 ;
        RECT 26.725 131.185 26.955 132.325 ;
        RECT 27.165 131.565 27.680 131.975 ;
        RECT 27.915 131.565 28.085 132.325 ;
        RECT 28.255 131.985 30.285 132.155 ;
        RECT 23.485 130.545 24.235 131.065 ;
        RECT 20.725 129.775 21.935 130.525 ;
        RECT 22.565 129.775 24.235 130.545 ;
        RECT 24.405 129.775 24.695 130.500 ;
        RECT 25.845 129.775 26.055 130.595 ;
        RECT 26.225 130.575 26.475 131.175 ;
        RECT 26.645 130.765 26.975 131.015 ;
        RECT 27.165 130.755 27.505 131.565 ;
        RECT 28.255 131.320 28.425 131.985 ;
        RECT 28.820 131.645 29.945 131.815 ;
        RECT 27.675 131.130 28.425 131.320 ;
        RECT 28.595 131.305 29.605 131.475 ;
        RECT 26.225 129.945 26.555 130.575 ;
        RECT 26.725 129.775 26.955 130.595 ;
        RECT 27.165 130.585 28.395 130.755 ;
        RECT 27.440 129.980 27.685 130.585 ;
        RECT 27.905 129.775 28.415 130.310 ;
        RECT 28.595 129.945 28.785 131.305 ;
        RECT 28.955 130.965 29.230 131.105 ;
        RECT 28.955 130.795 29.235 130.965 ;
        RECT 28.955 129.945 29.230 130.795 ;
        RECT 29.435 130.505 29.605 131.305 ;
        RECT 29.775 130.515 29.945 131.645 ;
        RECT 30.115 131.015 30.285 131.985 ;
        RECT 30.455 131.185 30.625 132.325 ;
        RECT 30.795 131.185 31.130 132.155 ;
        RECT 31.395 131.580 31.665 132.325 ;
        RECT 32.295 132.320 38.570 132.325 ;
        RECT 31.835 131.410 32.125 132.150 ;
        RECT 32.295 131.595 32.550 132.320 ;
        RECT 32.735 131.425 32.995 132.150 ;
        RECT 33.165 131.595 33.410 132.320 ;
        RECT 33.595 131.425 33.855 132.150 ;
        RECT 34.025 131.595 34.270 132.320 ;
        RECT 34.455 131.425 34.715 132.150 ;
        RECT 34.885 131.595 35.130 132.320 ;
        RECT 35.300 131.425 35.560 132.150 ;
        RECT 35.730 131.595 35.990 132.320 ;
        RECT 36.160 131.425 36.420 132.150 ;
        RECT 36.590 131.595 36.850 132.320 ;
        RECT 37.020 131.425 37.280 132.150 ;
        RECT 37.450 131.595 37.710 132.320 ;
        RECT 37.880 131.425 38.140 132.150 ;
        RECT 38.310 131.525 38.570 132.320 ;
        RECT 32.735 131.410 38.140 131.425 ;
        RECT 31.395 131.305 38.140 131.410 ;
        RECT 30.115 130.685 30.310 131.015 ;
        RECT 30.535 130.685 30.790 131.015 ;
        RECT 30.535 130.515 30.705 130.685 ;
        RECT 30.960 130.515 31.130 131.185 ;
        RECT 31.365 131.185 38.140 131.305 ;
        RECT 31.365 131.135 32.560 131.185 ;
        RECT 29.775 130.345 30.705 130.515 ;
        RECT 29.775 130.310 29.950 130.345 ;
        RECT 29.420 129.945 29.950 130.310 ;
        RECT 30.375 129.775 30.705 130.175 ;
        RECT 30.875 129.945 31.130 130.515 ;
        RECT 31.395 130.595 32.560 131.135 ;
        RECT 38.740 131.015 38.990 132.150 ;
        RECT 39.170 131.515 39.430 132.325 ;
        RECT 39.605 131.015 39.850 132.155 ;
        RECT 40.030 131.515 40.325 132.325 ;
        RECT 40.880 131.985 41.135 132.015 ;
        RECT 40.795 131.815 41.135 131.985 ;
        RECT 40.880 131.345 41.135 131.815 ;
        RECT 41.315 131.525 41.600 132.325 ;
        RECT 41.780 131.605 42.110 132.115 ;
        RECT 32.730 130.765 39.850 131.015 ;
        RECT 31.395 130.425 38.140 130.595 ;
        RECT 31.395 129.775 31.695 130.255 ;
        RECT 31.865 129.970 32.125 130.425 ;
        RECT 32.295 129.775 32.555 130.255 ;
        RECT 32.735 129.970 32.995 130.425 ;
        RECT 33.165 129.775 33.415 130.255 ;
        RECT 33.595 129.970 33.855 130.425 ;
        RECT 34.025 129.775 34.275 130.255 ;
        RECT 34.455 129.970 34.715 130.425 ;
        RECT 34.885 129.775 35.130 130.255 ;
        RECT 35.300 129.970 35.575 130.425 ;
        RECT 35.745 129.775 35.990 130.255 ;
        RECT 36.160 129.970 36.420 130.425 ;
        RECT 36.590 129.775 36.850 130.255 ;
        RECT 37.020 129.970 37.280 130.425 ;
        RECT 37.450 129.775 37.710 130.255 ;
        RECT 37.880 129.970 38.140 130.425 ;
        RECT 38.310 129.775 38.570 130.335 ;
        RECT 38.740 129.955 38.990 130.765 ;
        RECT 39.170 129.775 39.430 130.300 ;
        RECT 39.600 129.955 39.850 130.765 ;
        RECT 40.020 130.455 40.335 131.015 ;
        RECT 40.880 130.485 41.060 131.345 ;
        RECT 41.780 131.015 42.030 131.605 ;
        RECT 42.380 131.455 42.550 132.065 ;
        RECT 42.720 131.635 43.050 132.325 ;
        RECT 43.280 131.775 43.520 132.065 ;
        RECT 43.720 131.945 44.140 132.325 ;
        RECT 44.320 131.855 44.950 132.105 ;
        RECT 45.420 131.945 45.750 132.325 ;
        RECT 44.320 131.775 44.490 131.855 ;
        RECT 45.920 131.775 46.090 132.065 ;
        RECT 46.270 131.945 46.650 132.325 ;
        RECT 46.890 131.940 47.720 132.110 ;
        RECT 43.280 131.605 44.490 131.775 ;
        RECT 41.230 130.685 42.030 131.015 ;
        RECT 40.030 129.775 40.335 130.285 ;
        RECT 40.880 129.955 41.135 130.485 ;
        RECT 41.315 129.775 41.600 130.235 ;
        RECT 41.780 130.035 42.030 130.685 ;
        RECT 42.230 131.435 42.550 131.455 ;
        RECT 42.230 131.265 44.150 131.435 ;
        RECT 42.230 130.370 42.420 131.265 ;
        RECT 44.320 131.095 44.490 131.605 ;
        RECT 44.660 131.345 45.180 131.655 ;
        RECT 42.590 130.925 44.490 131.095 ;
        RECT 42.590 130.865 42.920 130.925 ;
        RECT 43.070 130.695 43.400 130.755 ;
        RECT 42.740 130.425 43.400 130.695 ;
        RECT 42.230 130.040 42.550 130.370 ;
        RECT 42.730 129.775 43.390 130.255 ;
        RECT 43.590 130.165 43.760 130.925 ;
        RECT 44.660 130.755 44.840 131.165 ;
        RECT 43.930 130.585 44.260 130.705 ;
        RECT 45.010 130.585 45.180 131.345 ;
        RECT 43.930 130.415 45.180 130.585 ;
        RECT 45.350 131.525 46.720 131.775 ;
        RECT 45.350 130.755 45.540 131.525 ;
        RECT 46.470 131.265 46.720 131.525 ;
        RECT 45.710 131.095 45.960 131.255 ;
        RECT 46.890 131.095 47.060 131.940 ;
        RECT 47.955 131.655 48.125 132.155 ;
        RECT 48.295 131.825 48.625 132.325 ;
        RECT 47.230 131.265 47.730 131.645 ;
        RECT 47.955 131.485 48.650 131.655 ;
        RECT 45.710 130.925 47.060 131.095 ;
        RECT 46.640 130.885 47.060 130.925 ;
        RECT 45.350 130.415 45.770 130.755 ;
        RECT 46.060 130.425 46.470 130.755 ;
        RECT 43.590 129.995 44.440 130.165 ;
        RECT 45.000 129.775 45.320 130.235 ;
        RECT 45.520 129.985 45.770 130.415 ;
        RECT 46.060 129.775 46.470 130.215 ;
        RECT 46.640 130.155 46.810 130.885 ;
        RECT 46.980 130.335 47.330 130.705 ;
        RECT 47.510 130.395 47.730 131.265 ;
        RECT 47.900 130.695 48.310 131.315 ;
        RECT 48.480 130.515 48.650 131.485 ;
        RECT 47.955 130.325 48.650 130.515 ;
        RECT 46.640 129.955 47.655 130.155 ;
        RECT 47.955 129.995 48.125 130.325 ;
        RECT 48.295 129.775 48.625 130.155 ;
        RECT 48.840 130.035 49.065 132.155 ;
        RECT 49.235 131.825 49.565 132.325 ;
        RECT 49.735 131.655 49.905 132.155 ;
        RECT 49.240 131.485 49.905 131.655 ;
        RECT 49.240 130.495 49.470 131.485 ;
        RECT 49.640 130.665 49.990 131.315 ;
        RECT 50.165 131.160 50.455 132.325 ;
        RECT 51.145 131.185 51.355 132.325 ;
        RECT 51.525 131.175 51.855 132.155 ;
        RECT 52.025 131.185 52.255 132.325 ;
        RECT 52.465 131.565 52.980 131.975 ;
        RECT 53.215 131.565 53.385 132.325 ;
        RECT 53.555 131.985 55.585 132.155 ;
        RECT 49.240 130.325 49.905 130.495 ;
        RECT 49.235 129.775 49.565 130.155 ;
        RECT 49.735 130.035 49.905 130.325 ;
        RECT 50.165 129.775 50.455 130.500 ;
        RECT 51.145 129.775 51.355 130.595 ;
        RECT 51.525 130.575 51.775 131.175 ;
        RECT 51.945 130.765 52.275 131.015 ;
        RECT 52.465 130.755 52.805 131.565 ;
        RECT 53.555 131.320 53.725 131.985 ;
        RECT 54.120 131.645 55.245 131.815 ;
        RECT 52.975 131.130 53.725 131.320 ;
        RECT 53.895 131.305 54.905 131.475 ;
        RECT 51.525 129.945 51.855 130.575 ;
        RECT 52.025 129.775 52.255 130.595 ;
        RECT 52.465 130.585 53.695 130.755 ;
        RECT 52.740 129.980 52.985 130.585 ;
        RECT 53.205 129.775 53.715 130.310 ;
        RECT 53.895 129.945 54.085 131.305 ;
        RECT 54.255 130.285 54.530 131.105 ;
        RECT 54.735 130.505 54.905 131.305 ;
        RECT 55.075 130.515 55.245 131.645 ;
        RECT 55.415 131.015 55.585 131.985 ;
        RECT 55.755 131.185 55.925 132.325 ;
        RECT 56.095 131.185 56.430 132.155 ;
        RECT 56.605 131.490 56.990 132.325 ;
        RECT 57.160 131.320 57.420 132.125 ;
        RECT 57.590 131.490 57.850 132.325 ;
        RECT 58.020 131.320 58.275 132.125 ;
        RECT 58.450 131.490 58.710 132.325 ;
        RECT 58.880 131.320 59.135 132.125 ;
        RECT 59.310 131.490 59.655 132.325 ;
        RECT 55.415 130.685 55.610 131.015 ;
        RECT 55.835 130.685 56.090 131.015 ;
        RECT 55.835 130.515 56.005 130.685 ;
        RECT 56.260 130.515 56.430 131.185 ;
        RECT 55.075 130.345 56.005 130.515 ;
        RECT 55.075 130.310 55.250 130.345 ;
        RECT 54.255 130.115 54.535 130.285 ;
        RECT 54.255 129.945 54.530 130.115 ;
        RECT 54.720 129.945 55.250 130.310 ;
        RECT 55.675 129.775 56.005 130.175 ;
        RECT 56.175 129.945 56.430 130.515 ;
        RECT 56.605 131.150 59.635 131.320 ;
        RECT 56.605 130.585 56.905 131.150 ;
        RECT 57.080 130.755 59.295 130.980 ;
        RECT 59.465 130.585 59.635 131.150 ;
        RECT 59.825 131.235 63.335 132.325 ;
        RECT 63.505 131.250 63.775 132.155 ;
        RECT 63.945 131.565 64.275 132.325 ;
        RECT 64.455 131.395 64.625 132.155 ;
        RECT 59.825 130.715 61.515 131.235 ;
        RECT 56.605 130.415 59.635 130.585 ;
        RECT 61.685 130.545 63.335 131.065 ;
        RECT 57.125 129.775 57.425 130.245 ;
        RECT 57.595 129.970 57.850 130.415 ;
        RECT 58.020 129.775 58.280 130.245 ;
        RECT 58.450 129.970 58.710 130.415 ;
        RECT 58.880 129.775 59.175 130.245 ;
        RECT 59.825 129.775 63.335 130.545 ;
        RECT 63.505 130.450 63.675 131.250 ;
        RECT 63.960 131.225 64.625 131.395 ;
        RECT 65.345 131.235 67.935 132.325 ;
        RECT 68.105 131.565 68.620 131.975 ;
        RECT 68.855 131.565 69.025 132.325 ;
        RECT 69.195 131.985 71.225 132.155 ;
        RECT 63.960 131.080 64.130 131.225 ;
        RECT 63.845 130.750 64.130 131.080 ;
        RECT 63.960 130.495 64.130 130.750 ;
        RECT 64.365 130.675 64.695 131.045 ;
        RECT 65.345 130.715 66.555 131.235 ;
        RECT 66.725 130.545 67.935 131.065 ;
        RECT 68.105 130.755 68.445 131.565 ;
        RECT 69.195 131.320 69.365 131.985 ;
        RECT 69.760 131.645 70.885 131.815 ;
        RECT 68.615 131.130 69.365 131.320 ;
        RECT 69.535 131.305 70.545 131.475 ;
        RECT 68.105 130.585 69.335 130.755 ;
        RECT 63.505 129.945 63.765 130.450 ;
        RECT 63.960 130.325 64.625 130.495 ;
        RECT 63.945 129.775 64.275 130.155 ;
        RECT 64.455 129.945 64.625 130.325 ;
        RECT 65.345 129.775 67.935 130.545 ;
        RECT 68.380 129.980 68.625 130.585 ;
        RECT 68.845 129.775 69.355 130.310 ;
        RECT 69.535 129.945 69.725 131.305 ;
        RECT 69.895 130.285 70.170 131.105 ;
        RECT 70.375 130.505 70.545 131.305 ;
        RECT 70.715 130.515 70.885 131.645 ;
        RECT 71.055 131.015 71.225 131.985 ;
        RECT 71.395 131.185 71.565 132.325 ;
        RECT 71.735 131.185 72.070 132.155 ;
        RECT 71.055 130.685 71.250 131.015 ;
        RECT 71.475 130.685 71.730 131.015 ;
        RECT 71.475 130.515 71.645 130.685 ;
        RECT 71.900 130.515 72.070 131.185 ;
        RECT 70.715 130.345 71.645 130.515 ;
        RECT 70.715 130.310 70.890 130.345 ;
        RECT 69.895 130.115 70.175 130.285 ;
        RECT 69.895 129.945 70.170 130.115 ;
        RECT 70.360 129.945 70.890 130.310 ;
        RECT 71.315 129.775 71.645 130.175 ;
        RECT 71.815 129.945 72.070 130.515 ;
        RECT 73.165 131.355 73.475 132.155 ;
        RECT 73.645 131.525 73.955 132.325 ;
        RECT 74.125 131.695 74.385 132.155 ;
        RECT 74.555 131.865 74.810 132.325 ;
        RECT 74.985 131.695 75.245 132.155 ;
        RECT 74.125 131.525 75.245 131.695 ;
        RECT 73.165 131.185 74.195 131.355 ;
        RECT 73.165 130.275 73.335 131.185 ;
        RECT 73.505 130.445 73.855 131.015 ;
        RECT 74.025 130.935 74.195 131.185 ;
        RECT 74.985 131.275 75.245 131.525 ;
        RECT 75.415 131.455 75.700 132.325 ;
        RECT 74.985 131.105 75.740 131.275 ;
        RECT 75.925 131.160 76.215 132.325 ;
        RECT 76.425 131.185 76.655 132.325 ;
        RECT 76.825 131.175 77.155 132.155 ;
        RECT 77.325 131.185 77.535 132.325 ;
        RECT 77.770 131.185 78.105 132.155 ;
        RECT 78.275 131.185 78.445 132.325 ;
        RECT 78.615 131.985 80.645 132.155 ;
        RECT 74.025 130.765 75.165 130.935 ;
        RECT 75.335 130.595 75.740 131.105 ;
        RECT 76.405 130.765 76.735 131.015 ;
        RECT 74.090 130.425 75.740 130.595 ;
        RECT 73.165 129.945 73.465 130.275 ;
        RECT 73.635 129.775 73.910 130.255 ;
        RECT 74.090 130.035 74.385 130.425 ;
        RECT 74.555 129.775 74.810 130.255 ;
        RECT 74.985 130.035 75.245 130.425 ;
        RECT 75.415 129.775 75.695 130.255 ;
        RECT 75.925 129.775 76.215 130.500 ;
        RECT 76.425 129.775 76.655 130.595 ;
        RECT 76.905 130.575 77.155 131.175 ;
        RECT 76.825 129.945 77.155 130.575 ;
        RECT 77.325 129.775 77.535 130.595 ;
        RECT 77.770 130.515 77.940 131.185 ;
        RECT 78.615 131.015 78.785 131.985 ;
        RECT 78.110 130.685 78.365 131.015 ;
        RECT 78.590 130.685 78.785 131.015 ;
        RECT 78.955 131.645 80.080 131.815 ;
        RECT 78.195 130.515 78.365 130.685 ;
        RECT 78.955 130.515 79.125 131.645 ;
        RECT 77.770 129.945 78.025 130.515 ;
        RECT 78.195 130.345 79.125 130.515 ;
        RECT 79.295 131.305 80.305 131.475 ;
        RECT 79.295 130.505 79.465 131.305 ;
        RECT 78.950 130.310 79.125 130.345 ;
        RECT 78.195 129.775 78.525 130.175 ;
        RECT 78.950 129.945 79.480 130.310 ;
        RECT 79.670 130.285 79.945 131.105 ;
        RECT 79.665 130.115 79.945 130.285 ;
        RECT 79.670 129.945 79.945 130.115 ;
        RECT 80.115 129.945 80.305 131.305 ;
        RECT 80.475 131.320 80.645 131.985 ;
        RECT 80.815 131.565 80.985 132.325 ;
        RECT 81.220 131.565 81.735 131.975 ;
        RECT 80.475 131.130 81.225 131.320 ;
        RECT 81.395 130.755 81.735 131.565 ;
        RECT 80.505 130.585 81.735 130.755 ;
        RECT 81.905 131.565 82.420 131.975 ;
        RECT 82.655 131.565 82.825 132.325 ;
        RECT 82.995 131.985 85.025 132.155 ;
        RECT 81.905 130.755 82.245 131.565 ;
        RECT 82.995 131.320 83.165 131.985 ;
        RECT 83.560 131.645 84.685 131.815 ;
        RECT 82.415 131.130 83.165 131.320 ;
        RECT 83.335 131.305 84.345 131.475 ;
        RECT 81.905 130.585 83.135 130.755 ;
        RECT 80.485 129.775 80.995 130.310 ;
        RECT 81.215 129.980 81.460 130.585 ;
        RECT 82.180 129.980 82.425 130.585 ;
        RECT 82.645 129.775 83.155 130.310 ;
        RECT 83.335 129.945 83.525 131.305 ;
        RECT 83.695 130.965 83.970 131.105 ;
        RECT 83.695 130.795 83.975 130.965 ;
        RECT 83.695 129.945 83.970 130.795 ;
        RECT 84.175 130.505 84.345 131.305 ;
        RECT 84.515 130.515 84.685 131.645 ;
        RECT 84.855 131.015 85.025 131.985 ;
        RECT 85.195 131.185 85.365 132.325 ;
        RECT 85.535 131.185 85.870 132.155 ;
        RECT 84.855 130.685 85.050 131.015 ;
        RECT 85.275 130.685 85.530 131.015 ;
        RECT 85.275 130.515 85.445 130.685 ;
        RECT 85.700 130.515 85.870 131.185 ;
        RECT 86.045 131.235 87.715 132.325 ;
        RECT 87.890 131.890 93.235 132.325 ;
        RECT 86.045 130.715 86.795 131.235 ;
        RECT 86.965 130.545 87.715 131.065 ;
        RECT 89.480 130.640 89.830 131.890 ;
        RECT 93.445 131.185 93.675 132.325 ;
        RECT 93.845 131.175 94.175 132.155 ;
        RECT 94.345 131.185 94.555 132.325 ;
        RECT 94.785 131.565 95.300 131.975 ;
        RECT 95.535 131.565 95.705 132.325 ;
        RECT 95.875 131.985 97.905 132.155 ;
        RECT 84.515 130.345 85.445 130.515 ;
        RECT 84.515 130.310 84.690 130.345 ;
        RECT 84.160 129.945 84.690 130.310 ;
        RECT 85.115 129.775 85.445 130.175 ;
        RECT 85.615 129.945 85.870 130.515 ;
        RECT 86.045 129.775 87.715 130.545 ;
        RECT 91.310 130.320 91.650 131.150 ;
        RECT 93.425 130.765 93.755 131.015 ;
        RECT 87.890 129.775 93.235 130.320 ;
        RECT 93.445 129.775 93.675 130.595 ;
        RECT 93.925 130.575 94.175 131.175 ;
        RECT 94.785 130.755 95.125 131.565 ;
        RECT 95.875 131.320 96.045 131.985 ;
        RECT 96.440 131.645 97.565 131.815 ;
        RECT 95.295 131.130 96.045 131.320 ;
        RECT 96.215 131.305 97.225 131.475 ;
        RECT 93.845 129.945 94.175 130.575 ;
        RECT 94.345 129.775 94.555 130.595 ;
        RECT 94.785 130.585 96.015 130.755 ;
        RECT 95.060 129.980 95.305 130.585 ;
        RECT 95.525 129.775 96.035 130.310 ;
        RECT 96.215 129.945 96.405 131.305 ;
        RECT 96.575 130.625 96.850 131.105 ;
        RECT 96.575 130.455 96.855 130.625 ;
        RECT 97.055 130.505 97.225 131.305 ;
        RECT 97.395 130.515 97.565 131.645 ;
        RECT 97.735 131.015 97.905 131.985 ;
        RECT 98.075 131.185 98.245 132.325 ;
        RECT 98.415 131.185 98.750 132.155 ;
        RECT 97.735 130.685 97.930 131.015 ;
        RECT 98.155 130.685 98.410 131.015 ;
        RECT 98.155 130.515 98.325 130.685 ;
        RECT 98.580 130.515 98.750 131.185 ;
        RECT 96.575 129.945 96.850 130.455 ;
        RECT 97.395 130.345 98.325 130.515 ;
        RECT 97.395 130.310 97.570 130.345 ;
        RECT 97.040 129.945 97.570 130.310 ;
        RECT 97.995 129.775 98.325 130.175 ;
        RECT 98.495 129.945 98.750 130.515 ;
        RECT 98.925 131.250 99.195 132.155 ;
        RECT 99.365 131.565 99.695 132.325 ;
        RECT 99.875 131.395 100.045 132.155 ;
        RECT 98.925 130.450 99.095 131.250 ;
        RECT 99.380 131.225 100.045 131.395 ;
        RECT 100.305 131.235 101.515 132.325 ;
        RECT 99.380 131.080 99.550 131.225 ;
        RECT 99.265 130.750 99.550 131.080 ;
        RECT 99.380 130.495 99.550 130.750 ;
        RECT 99.785 130.675 100.115 131.045 ;
        RECT 100.305 130.695 100.825 131.235 ;
        RECT 101.685 131.160 101.975 132.325 ;
        RECT 102.145 131.235 103.355 132.325 ;
        RECT 103.580 131.455 103.865 132.325 ;
        RECT 104.035 131.695 104.295 132.155 ;
        RECT 104.470 131.865 104.725 132.325 ;
        RECT 104.895 131.695 105.155 132.155 ;
        RECT 104.035 131.525 105.155 131.695 ;
        RECT 105.325 131.525 105.635 132.325 ;
        RECT 104.035 131.275 104.295 131.525 ;
        RECT 105.805 131.355 106.115 132.155 ;
        RECT 100.995 130.525 101.515 131.065 ;
        RECT 102.145 130.695 102.665 131.235 ;
        RECT 103.540 131.105 104.295 131.275 ;
        RECT 105.085 131.185 106.115 131.355 ;
        RECT 102.835 130.525 103.355 131.065 ;
        RECT 98.925 129.945 99.185 130.450 ;
        RECT 99.380 130.325 100.045 130.495 ;
        RECT 99.365 129.775 99.695 130.155 ;
        RECT 99.875 129.945 100.045 130.325 ;
        RECT 100.305 129.775 101.515 130.525 ;
        RECT 101.685 129.775 101.975 130.500 ;
        RECT 102.145 129.775 103.355 130.525 ;
        RECT 103.540 130.595 103.945 131.105 ;
        RECT 105.085 130.935 105.255 131.185 ;
        RECT 104.115 130.765 105.255 130.935 ;
        RECT 103.540 130.425 105.190 130.595 ;
        RECT 105.425 130.445 105.775 131.015 ;
        RECT 103.585 129.775 103.865 130.255 ;
        RECT 104.035 130.035 104.295 130.425 ;
        RECT 104.470 129.775 104.725 130.255 ;
        RECT 104.895 130.035 105.190 130.425 ;
        RECT 105.945 130.275 106.115 131.185 ;
        RECT 105.370 129.775 105.645 130.255 ;
        RECT 105.815 129.945 106.115 130.275 ;
        RECT 106.285 131.605 106.745 132.155 ;
        RECT 106.935 131.605 107.265 132.325 ;
        RECT 106.285 130.235 106.535 131.605 ;
        RECT 107.465 131.435 107.765 131.985 ;
        RECT 107.935 131.655 108.215 132.325 ;
        RECT 106.825 131.265 107.765 131.435 ;
        RECT 106.825 131.015 106.995 131.265 ;
        RECT 108.135 131.015 108.400 131.375 ;
        RECT 106.705 130.685 106.995 131.015 ;
        RECT 107.165 130.765 107.505 131.015 ;
        RECT 107.725 130.765 108.400 131.015 ;
        RECT 108.585 131.235 110.255 132.325 ;
        RECT 110.425 131.565 110.940 131.975 ;
        RECT 111.175 131.565 111.345 132.325 ;
        RECT 111.515 131.985 113.545 132.155 ;
        RECT 108.585 130.715 109.335 131.235 ;
        RECT 106.825 130.595 106.995 130.685 ;
        RECT 106.825 130.405 108.215 130.595 ;
        RECT 109.505 130.545 110.255 131.065 ;
        RECT 110.425 130.755 110.765 131.565 ;
        RECT 111.515 131.320 111.685 131.985 ;
        RECT 112.080 131.645 113.205 131.815 ;
        RECT 110.935 131.130 111.685 131.320 ;
        RECT 111.855 131.305 112.865 131.475 ;
        RECT 110.425 130.585 111.655 130.755 ;
        RECT 106.285 129.945 106.845 130.235 ;
        RECT 107.015 129.775 107.265 130.235 ;
        RECT 107.885 130.045 108.215 130.405 ;
        RECT 108.585 129.775 110.255 130.545 ;
        RECT 110.700 129.980 110.945 130.585 ;
        RECT 111.165 129.775 111.675 130.310 ;
        RECT 111.855 129.945 112.045 131.305 ;
        RECT 112.215 130.285 112.490 131.105 ;
        RECT 112.695 130.505 112.865 131.305 ;
        RECT 113.035 130.515 113.205 131.645 ;
        RECT 113.375 131.015 113.545 131.985 ;
        RECT 113.715 131.185 113.885 132.325 ;
        RECT 114.055 131.185 114.390 132.155 ;
        RECT 113.375 130.685 113.570 131.015 ;
        RECT 113.795 130.685 114.050 131.015 ;
        RECT 113.795 130.515 113.965 130.685 ;
        RECT 114.220 130.515 114.390 131.185 ;
        RECT 114.565 131.235 118.075 132.325 ;
        RECT 114.565 130.715 116.255 131.235 ;
        RECT 118.285 131.185 118.515 132.325 ;
        RECT 118.685 131.175 119.015 132.155 ;
        RECT 119.185 131.185 119.395 132.325 ;
        RECT 120.635 131.395 120.805 132.155 ;
        RECT 120.985 131.565 121.315 132.325 ;
        RECT 120.635 131.225 121.300 131.395 ;
        RECT 121.485 131.250 121.755 132.155 ;
        RECT 116.425 130.545 118.075 131.065 ;
        RECT 118.265 130.765 118.595 131.015 ;
        RECT 113.035 130.345 113.965 130.515 ;
        RECT 113.035 130.310 113.210 130.345 ;
        RECT 112.215 130.115 112.495 130.285 ;
        RECT 112.215 129.945 112.490 130.115 ;
        RECT 112.680 129.945 113.210 130.310 ;
        RECT 113.635 129.775 113.965 130.175 ;
        RECT 114.135 129.945 114.390 130.515 ;
        RECT 114.565 129.775 118.075 130.545 ;
        RECT 118.285 129.775 118.515 130.595 ;
        RECT 118.765 130.575 119.015 131.175 ;
        RECT 121.130 131.080 121.300 131.225 ;
        RECT 120.565 130.675 120.895 131.045 ;
        RECT 121.130 130.750 121.415 131.080 ;
        RECT 118.685 129.945 119.015 130.575 ;
        RECT 119.185 129.775 119.395 130.595 ;
        RECT 121.130 130.495 121.300 130.750 ;
        RECT 120.635 130.325 121.300 130.495 ;
        RECT 121.585 130.450 121.755 131.250 ;
        RECT 122.845 131.235 126.355 132.325 ;
        RECT 126.525 131.235 127.735 132.325 ;
        RECT 122.845 130.715 124.535 131.235 ;
        RECT 124.705 130.545 126.355 131.065 ;
        RECT 126.525 130.695 127.045 131.235 ;
        RECT 120.635 129.945 120.805 130.325 ;
        RECT 120.985 129.775 121.315 130.155 ;
        RECT 121.495 129.945 121.755 130.450 ;
        RECT 122.845 129.775 126.355 130.545 ;
        RECT 127.215 130.525 127.735 131.065 ;
        RECT 126.525 129.775 127.735 130.525 ;
        RECT 20.640 129.605 127.820 129.775 ;
        RECT 20.725 128.855 21.935 129.605 ;
        RECT 22.570 129.060 27.915 129.605 ;
        RECT 20.725 128.315 21.245 128.855 ;
        RECT 21.415 128.145 21.935 128.685 ;
        RECT 20.725 127.055 21.935 128.145 ;
        RECT 24.160 127.490 24.510 128.740 ;
        RECT 25.990 128.230 26.330 129.060 ;
        RECT 28.360 128.795 28.605 129.400 ;
        RECT 28.825 129.070 29.335 129.605 ;
        RECT 28.085 128.625 29.315 128.795 ;
        RECT 28.085 127.815 28.425 128.625 ;
        RECT 28.595 128.060 29.345 128.250 ;
        RECT 22.570 127.055 27.915 127.490 ;
        RECT 28.085 127.405 28.600 127.815 ;
        RECT 28.835 127.055 29.005 127.815 ;
        RECT 29.175 127.395 29.345 128.060 ;
        RECT 29.515 128.075 29.705 129.435 ;
        RECT 29.875 128.585 30.150 129.435 ;
        RECT 30.340 129.070 30.870 129.435 ;
        RECT 31.295 129.205 31.625 129.605 ;
        RECT 30.695 129.035 30.870 129.070 ;
        RECT 29.875 128.415 30.155 128.585 ;
        RECT 29.875 128.275 30.150 128.415 ;
        RECT 30.355 128.075 30.525 128.875 ;
        RECT 29.515 127.905 30.525 128.075 ;
        RECT 30.695 128.865 31.625 129.035 ;
        RECT 31.795 128.865 32.050 129.435 ;
        RECT 30.695 127.735 30.865 128.865 ;
        RECT 31.455 128.695 31.625 128.865 ;
        RECT 29.740 127.565 30.865 127.735 ;
        RECT 31.035 128.365 31.230 128.695 ;
        RECT 31.455 128.365 31.710 128.695 ;
        RECT 31.035 127.395 31.205 128.365 ;
        RECT 31.880 128.195 32.050 128.865 ;
        RECT 32.885 128.975 33.215 129.335 ;
        RECT 33.835 129.145 34.085 129.605 ;
        RECT 34.255 129.145 34.815 129.435 ;
        RECT 32.885 128.785 34.275 128.975 ;
        RECT 34.105 128.695 34.275 128.785 ;
        RECT 29.175 127.225 31.205 127.395 ;
        RECT 31.375 127.055 31.545 128.195 ;
        RECT 31.715 127.225 32.050 128.195 ;
        RECT 32.700 128.365 33.375 128.615 ;
        RECT 33.595 128.365 33.935 128.615 ;
        RECT 34.105 128.365 34.395 128.695 ;
        RECT 32.700 128.005 32.965 128.365 ;
        RECT 34.105 128.115 34.275 128.365 ;
        RECT 33.335 127.945 34.275 128.115 ;
        RECT 32.885 127.055 33.165 127.725 ;
        RECT 33.335 127.395 33.635 127.945 ;
        RECT 34.565 127.775 34.815 129.145 ;
        RECT 35.185 128.975 35.515 129.335 ;
        RECT 36.135 129.145 36.385 129.605 ;
        RECT 36.555 129.145 37.115 129.435 ;
        RECT 35.185 128.785 36.575 128.975 ;
        RECT 36.405 128.695 36.575 128.785 ;
        RECT 35.000 128.365 35.675 128.615 ;
        RECT 35.895 128.365 36.235 128.615 ;
        RECT 36.405 128.365 36.695 128.695 ;
        RECT 35.000 128.005 35.265 128.365 ;
        RECT 36.405 128.115 36.575 128.365 ;
        RECT 33.835 127.055 34.165 127.775 ;
        RECT 34.355 127.225 34.815 127.775 ;
        RECT 35.635 127.945 36.575 128.115 ;
        RECT 35.185 127.055 35.465 127.725 ;
        RECT 35.635 127.395 35.935 127.945 ;
        RECT 36.865 127.775 37.115 129.145 ;
        RECT 37.285 128.880 37.575 129.605 ;
        RECT 38.205 129.145 38.765 129.435 ;
        RECT 38.935 129.145 39.185 129.605 ;
        RECT 36.135 127.055 36.465 127.775 ;
        RECT 36.655 127.225 37.115 127.775 ;
        RECT 37.285 127.055 37.575 128.220 ;
        RECT 38.205 127.775 38.455 129.145 ;
        RECT 39.805 128.975 40.135 129.335 ;
        RECT 38.745 128.785 40.135 128.975 ;
        RECT 41.625 128.975 41.955 129.335 ;
        RECT 42.575 129.145 42.825 129.605 ;
        RECT 42.995 129.145 43.555 129.435 ;
        RECT 44.100 129.265 44.355 129.425 ;
        RECT 41.625 128.785 43.015 128.975 ;
        RECT 38.745 128.695 38.915 128.785 ;
        RECT 38.625 128.365 38.915 128.695 ;
        RECT 42.845 128.695 43.015 128.785 ;
        RECT 39.085 128.365 39.425 128.615 ;
        RECT 39.645 128.365 40.320 128.615 ;
        RECT 38.745 128.115 38.915 128.365 ;
        RECT 38.745 127.945 39.685 128.115 ;
        RECT 40.055 128.005 40.320 128.365 ;
        RECT 41.440 128.365 42.115 128.615 ;
        RECT 42.335 128.365 42.675 128.615 ;
        RECT 42.845 128.365 43.135 128.695 ;
        RECT 41.440 128.005 41.705 128.365 ;
        RECT 42.845 128.115 43.015 128.365 ;
        RECT 38.205 127.225 38.665 127.775 ;
        RECT 38.855 127.055 39.185 127.775 ;
        RECT 39.385 127.395 39.685 127.945 ;
        RECT 42.075 127.945 43.015 128.115 ;
        RECT 39.855 127.055 40.135 127.725 ;
        RECT 41.625 127.055 41.905 127.725 ;
        RECT 42.075 127.395 42.375 127.945 ;
        RECT 43.305 127.775 43.555 129.145 ;
        RECT 44.015 129.095 44.355 129.265 ;
        RECT 44.535 129.145 44.820 129.605 ;
        RECT 42.575 127.055 42.905 127.775 ;
        RECT 43.095 127.225 43.555 127.775 ;
        RECT 44.100 128.895 44.355 129.095 ;
        RECT 44.100 128.035 44.280 128.895 ;
        RECT 45.000 128.695 45.250 129.345 ;
        RECT 44.450 128.365 45.250 128.695 ;
        RECT 44.100 127.365 44.355 128.035 ;
        RECT 44.535 127.055 44.820 127.855 ;
        RECT 45.000 127.775 45.250 128.365 ;
        RECT 45.450 129.010 45.770 129.340 ;
        RECT 45.950 129.125 46.610 129.605 ;
        RECT 46.810 129.215 47.660 129.385 ;
        RECT 45.450 128.115 45.640 129.010 ;
        RECT 45.960 128.685 46.620 128.955 ;
        RECT 46.290 128.625 46.620 128.685 ;
        RECT 45.810 128.455 46.140 128.515 ;
        RECT 46.810 128.455 46.980 129.215 ;
        RECT 48.220 129.145 48.540 129.605 ;
        RECT 48.740 128.965 48.990 129.395 ;
        RECT 49.280 129.165 49.690 129.605 ;
        RECT 49.860 129.225 50.875 129.425 ;
        RECT 47.150 128.795 48.400 128.965 ;
        RECT 47.150 128.675 47.480 128.795 ;
        RECT 45.810 128.285 47.710 128.455 ;
        RECT 45.450 127.945 47.370 128.115 ;
        RECT 45.450 127.925 45.770 127.945 ;
        RECT 45.000 127.265 45.330 127.775 ;
        RECT 45.600 127.315 45.770 127.925 ;
        RECT 47.540 127.775 47.710 128.285 ;
        RECT 47.880 128.215 48.060 128.625 ;
        RECT 48.230 128.035 48.400 128.795 ;
        RECT 45.940 127.055 46.270 127.745 ;
        RECT 46.500 127.605 47.710 127.775 ;
        RECT 47.880 127.725 48.400 128.035 ;
        RECT 48.570 128.625 48.990 128.965 ;
        RECT 49.280 128.625 49.690 128.955 ;
        RECT 48.570 127.855 48.760 128.625 ;
        RECT 49.860 128.495 50.030 129.225 ;
        RECT 51.175 129.055 51.345 129.385 ;
        RECT 51.515 129.225 51.845 129.605 ;
        RECT 50.200 128.675 50.550 129.045 ;
        RECT 49.860 128.455 50.280 128.495 ;
        RECT 48.930 128.285 50.280 128.455 ;
        RECT 48.930 128.125 49.180 128.285 ;
        RECT 49.690 127.855 49.940 128.115 ;
        RECT 48.570 127.605 49.940 127.855 ;
        RECT 46.500 127.315 46.740 127.605 ;
        RECT 47.540 127.525 47.710 127.605 ;
        RECT 46.940 127.055 47.360 127.435 ;
        RECT 47.540 127.275 48.170 127.525 ;
        RECT 48.640 127.055 48.970 127.435 ;
        RECT 49.140 127.315 49.310 127.605 ;
        RECT 50.110 127.440 50.280 128.285 ;
        RECT 50.730 128.115 50.950 128.985 ;
        RECT 51.175 128.865 51.870 129.055 ;
        RECT 50.450 127.735 50.950 128.115 ;
        RECT 51.120 128.065 51.530 128.685 ;
        RECT 51.700 127.895 51.870 128.865 ;
        RECT 51.175 127.725 51.870 127.895 ;
        RECT 49.490 127.055 49.870 127.435 ;
        RECT 50.110 127.270 50.940 127.440 ;
        RECT 51.175 127.225 51.345 127.725 ;
        RECT 51.515 127.055 51.845 127.555 ;
        RECT 52.060 127.225 52.285 129.345 ;
        RECT 52.455 129.225 52.785 129.605 ;
        RECT 52.955 129.055 53.125 129.345 ;
        RECT 53.760 129.265 54.015 129.425 ;
        RECT 53.675 129.095 54.015 129.265 ;
        RECT 54.195 129.145 54.480 129.605 ;
        RECT 52.460 128.885 53.125 129.055 ;
        RECT 53.760 128.895 54.015 129.095 ;
        RECT 52.460 127.895 52.690 128.885 ;
        RECT 52.860 128.065 53.210 128.715 ;
        RECT 53.760 128.035 53.940 128.895 ;
        RECT 54.660 128.695 54.910 129.345 ;
        RECT 54.110 128.365 54.910 128.695 ;
        RECT 52.460 127.725 53.125 127.895 ;
        RECT 52.455 127.055 52.785 127.555 ;
        RECT 52.955 127.225 53.125 127.725 ;
        RECT 53.760 127.365 54.015 128.035 ;
        RECT 54.195 127.055 54.480 127.855 ;
        RECT 54.660 127.775 54.910 128.365 ;
        RECT 55.110 129.010 55.430 129.340 ;
        RECT 55.610 129.125 56.270 129.605 ;
        RECT 56.470 129.215 57.320 129.385 ;
        RECT 55.110 128.115 55.300 129.010 ;
        RECT 55.620 128.685 56.280 128.955 ;
        RECT 55.950 128.625 56.280 128.685 ;
        RECT 55.470 128.455 55.800 128.515 ;
        RECT 56.470 128.455 56.640 129.215 ;
        RECT 57.880 129.145 58.200 129.605 ;
        RECT 58.400 128.965 58.650 129.395 ;
        RECT 58.940 129.165 59.350 129.605 ;
        RECT 59.520 129.225 60.535 129.425 ;
        RECT 56.810 128.795 58.060 128.965 ;
        RECT 56.810 128.675 57.140 128.795 ;
        RECT 55.470 128.285 57.370 128.455 ;
        RECT 55.110 127.945 57.030 128.115 ;
        RECT 55.110 127.925 55.430 127.945 ;
        RECT 54.660 127.265 54.990 127.775 ;
        RECT 55.260 127.315 55.430 127.925 ;
        RECT 57.200 127.775 57.370 128.285 ;
        RECT 57.540 128.215 57.720 128.625 ;
        RECT 57.890 128.035 58.060 128.795 ;
        RECT 55.600 127.055 55.930 127.745 ;
        RECT 56.160 127.605 57.370 127.775 ;
        RECT 57.540 127.725 58.060 128.035 ;
        RECT 58.230 128.625 58.650 128.965 ;
        RECT 58.940 128.625 59.350 128.955 ;
        RECT 58.230 127.855 58.420 128.625 ;
        RECT 59.520 128.495 59.690 129.225 ;
        RECT 60.835 129.055 61.005 129.385 ;
        RECT 61.175 129.225 61.505 129.605 ;
        RECT 59.860 128.675 60.210 129.045 ;
        RECT 59.520 128.455 59.940 128.495 ;
        RECT 58.590 128.285 59.940 128.455 ;
        RECT 58.590 128.125 58.840 128.285 ;
        RECT 59.350 127.855 59.600 128.115 ;
        RECT 58.230 127.605 59.600 127.855 ;
        RECT 56.160 127.315 56.400 127.605 ;
        RECT 57.200 127.525 57.370 127.605 ;
        RECT 56.600 127.055 57.020 127.435 ;
        RECT 57.200 127.275 57.830 127.525 ;
        RECT 58.300 127.055 58.630 127.435 ;
        RECT 58.800 127.315 58.970 127.605 ;
        RECT 59.770 127.440 59.940 128.285 ;
        RECT 60.390 128.115 60.610 128.985 ;
        RECT 60.835 128.865 61.530 129.055 ;
        RECT 60.110 127.735 60.610 128.115 ;
        RECT 60.780 128.065 61.190 128.685 ;
        RECT 61.360 127.895 61.530 128.865 ;
        RECT 60.835 127.725 61.530 127.895 ;
        RECT 59.150 127.055 59.530 127.435 ;
        RECT 59.770 127.270 60.600 127.440 ;
        RECT 60.835 127.225 61.005 127.725 ;
        RECT 61.175 127.055 61.505 127.555 ;
        RECT 61.720 127.225 61.945 129.345 ;
        RECT 62.115 129.225 62.445 129.605 ;
        RECT 62.615 129.055 62.785 129.345 ;
        RECT 62.120 128.885 62.785 129.055 ;
        RECT 62.120 127.895 62.350 128.885 ;
        RECT 63.045 128.880 63.335 129.605 ;
        RECT 63.565 128.785 63.775 129.605 ;
        RECT 63.945 128.805 64.275 129.435 ;
        RECT 62.520 128.065 62.870 128.715 ;
        RECT 62.120 127.725 62.785 127.895 ;
        RECT 62.115 127.055 62.445 127.555 ;
        RECT 62.615 127.225 62.785 127.725 ;
        RECT 63.045 127.055 63.335 128.220 ;
        RECT 63.945 128.205 64.195 128.805 ;
        RECT 64.445 128.785 64.675 129.605 ;
        RECT 65.345 128.835 67.015 129.605 ;
        RECT 67.560 129.265 67.815 129.425 ;
        RECT 67.475 129.095 67.815 129.265 ;
        RECT 67.995 129.145 68.280 129.605 ;
        RECT 64.365 128.365 64.695 128.615 ;
        RECT 63.565 127.055 63.775 128.195 ;
        RECT 63.945 127.225 64.275 128.205 ;
        RECT 64.445 127.055 64.675 128.195 ;
        RECT 65.345 128.145 66.095 128.665 ;
        RECT 66.265 128.315 67.015 128.835 ;
        RECT 67.560 128.895 67.815 129.095 ;
        RECT 65.345 127.055 67.015 128.145 ;
        RECT 67.560 128.035 67.740 128.895 ;
        RECT 68.460 128.695 68.710 129.345 ;
        RECT 67.910 128.365 68.710 128.695 ;
        RECT 67.560 127.365 67.815 128.035 ;
        RECT 67.995 127.055 68.280 127.855 ;
        RECT 68.460 127.775 68.710 128.365 ;
        RECT 68.910 129.010 69.230 129.340 ;
        RECT 69.410 129.125 70.070 129.605 ;
        RECT 70.270 129.215 71.120 129.385 ;
        RECT 68.910 128.115 69.100 129.010 ;
        RECT 69.420 128.685 70.080 128.955 ;
        RECT 69.750 128.625 70.080 128.685 ;
        RECT 69.270 128.455 69.600 128.515 ;
        RECT 70.270 128.455 70.440 129.215 ;
        RECT 71.680 129.145 72.000 129.605 ;
        RECT 72.200 128.965 72.450 129.395 ;
        RECT 72.740 129.165 73.150 129.605 ;
        RECT 73.320 129.225 74.335 129.425 ;
        RECT 70.610 128.795 71.860 128.965 ;
        RECT 70.610 128.675 70.940 128.795 ;
        RECT 69.270 128.285 71.170 128.455 ;
        RECT 68.910 127.945 70.830 128.115 ;
        RECT 68.910 127.925 69.230 127.945 ;
        RECT 68.460 127.265 68.790 127.775 ;
        RECT 69.060 127.315 69.230 127.925 ;
        RECT 71.000 127.775 71.170 128.285 ;
        RECT 71.340 128.215 71.520 128.625 ;
        RECT 71.690 128.035 71.860 128.795 ;
        RECT 69.400 127.055 69.730 127.745 ;
        RECT 69.960 127.605 71.170 127.775 ;
        RECT 71.340 127.725 71.860 128.035 ;
        RECT 72.030 128.625 72.450 128.965 ;
        RECT 72.740 128.625 73.150 128.955 ;
        RECT 72.030 127.855 72.220 128.625 ;
        RECT 73.320 128.495 73.490 129.225 ;
        RECT 74.635 129.055 74.805 129.385 ;
        RECT 74.975 129.225 75.305 129.605 ;
        RECT 73.660 128.675 74.010 129.045 ;
        RECT 73.320 128.455 73.740 128.495 ;
        RECT 72.390 128.285 73.740 128.455 ;
        RECT 72.390 128.125 72.640 128.285 ;
        RECT 73.150 127.855 73.400 128.115 ;
        RECT 72.030 127.605 73.400 127.855 ;
        RECT 69.960 127.315 70.200 127.605 ;
        RECT 71.000 127.525 71.170 127.605 ;
        RECT 70.400 127.055 70.820 127.435 ;
        RECT 71.000 127.275 71.630 127.525 ;
        RECT 72.100 127.055 72.430 127.435 ;
        RECT 72.600 127.315 72.770 127.605 ;
        RECT 73.570 127.440 73.740 128.285 ;
        RECT 74.190 128.115 74.410 128.985 ;
        RECT 74.635 128.865 75.330 129.055 ;
        RECT 73.910 127.735 74.410 128.115 ;
        RECT 74.580 128.065 74.990 128.685 ;
        RECT 75.160 127.895 75.330 128.865 ;
        RECT 74.635 127.725 75.330 127.895 ;
        RECT 72.950 127.055 73.330 127.435 ;
        RECT 73.570 127.270 74.400 127.440 ;
        RECT 74.635 127.225 74.805 127.725 ;
        RECT 74.975 127.055 75.305 127.555 ;
        RECT 75.520 127.225 75.745 129.345 ;
        RECT 75.915 129.225 76.245 129.605 ;
        RECT 76.415 129.055 76.585 129.345 ;
        RECT 75.920 128.885 76.585 129.055 ;
        RECT 75.920 127.895 76.150 128.885 ;
        RECT 76.845 128.835 79.435 129.605 ;
        RECT 79.605 129.095 79.910 129.605 ;
        RECT 76.320 128.065 76.670 128.715 ;
        RECT 76.845 128.145 78.055 128.665 ;
        RECT 78.225 128.315 79.435 128.835 ;
        RECT 79.605 128.365 79.920 128.925 ;
        RECT 80.090 128.615 80.340 129.425 ;
        RECT 80.510 129.080 80.770 129.605 ;
        RECT 80.950 128.615 81.200 129.425 ;
        RECT 81.370 129.045 81.630 129.605 ;
        RECT 81.800 128.955 82.060 129.410 ;
        RECT 82.230 129.125 82.490 129.605 ;
        RECT 82.660 128.955 82.920 129.410 ;
        RECT 83.090 129.125 83.350 129.605 ;
        RECT 83.520 128.955 83.780 129.410 ;
        RECT 83.950 129.125 84.195 129.605 ;
        RECT 84.365 128.955 84.640 129.410 ;
        RECT 84.810 129.125 85.055 129.605 ;
        RECT 85.225 128.955 85.485 129.410 ;
        RECT 85.665 129.125 85.915 129.605 ;
        RECT 86.085 128.955 86.345 129.410 ;
        RECT 86.525 129.125 86.775 129.605 ;
        RECT 86.945 128.955 87.205 129.410 ;
        RECT 87.385 129.125 87.645 129.605 ;
        RECT 87.815 128.955 88.075 129.410 ;
        RECT 88.245 129.125 88.545 129.605 ;
        RECT 81.800 128.785 88.545 128.955 ;
        RECT 88.805 128.880 89.095 129.605 ;
        RECT 89.725 128.835 92.315 129.605 ;
        RECT 92.575 129.055 92.745 129.345 ;
        RECT 92.915 129.225 93.245 129.605 ;
        RECT 92.575 128.885 93.240 129.055 ;
        RECT 80.090 128.365 87.210 128.615 ;
        RECT 75.920 127.725 76.585 127.895 ;
        RECT 75.915 127.055 76.245 127.555 ;
        RECT 76.415 127.225 76.585 127.725 ;
        RECT 76.845 127.055 79.435 128.145 ;
        RECT 79.615 127.055 79.910 127.865 ;
        RECT 80.090 127.225 80.335 128.365 ;
        RECT 80.510 127.055 80.770 127.865 ;
        RECT 80.950 127.230 81.200 128.365 ;
        RECT 87.380 128.195 88.545 128.785 ;
        RECT 81.800 127.970 88.545 128.195 ;
        RECT 81.800 127.955 87.205 127.970 ;
        RECT 81.370 127.060 81.630 127.855 ;
        RECT 81.800 127.230 82.060 127.955 ;
        RECT 82.230 127.060 82.490 127.785 ;
        RECT 82.660 127.230 82.920 127.955 ;
        RECT 83.090 127.060 83.350 127.785 ;
        RECT 83.520 127.230 83.780 127.955 ;
        RECT 83.950 127.060 84.210 127.785 ;
        RECT 84.380 127.230 84.640 127.955 ;
        RECT 84.810 127.060 85.055 127.785 ;
        RECT 85.225 127.230 85.485 127.955 ;
        RECT 85.670 127.060 85.915 127.785 ;
        RECT 86.085 127.230 86.345 127.955 ;
        RECT 86.530 127.060 86.775 127.785 ;
        RECT 86.945 127.230 87.205 127.955 ;
        RECT 87.390 127.060 87.645 127.785 ;
        RECT 87.815 127.230 88.105 127.970 ;
        RECT 81.370 127.055 87.645 127.060 ;
        RECT 88.275 127.055 88.545 127.800 ;
        RECT 88.805 127.055 89.095 128.220 ;
        RECT 89.725 128.145 90.935 128.665 ;
        RECT 91.105 128.315 92.315 128.835 ;
        RECT 89.725 127.055 92.315 128.145 ;
        RECT 92.490 128.065 92.840 128.715 ;
        RECT 93.010 127.895 93.240 128.885 ;
        RECT 92.575 127.725 93.240 127.895 ;
        RECT 92.575 127.225 92.745 127.725 ;
        RECT 92.915 127.055 93.245 127.555 ;
        RECT 93.415 127.225 93.640 129.345 ;
        RECT 93.855 129.225 94.185 129.605 ;
        RECT 94.355 129.055 94.525 129.385 ;
        RECT 94.825 129.225 95.840 129.425 ;
        RECT 93.830 128.865 94.525 129.055 ;
        RECT 93.830 127.895 94.000 128.865 ;
        RECT 94.170 128.065 94.580 128.685 ;
        RECT 94.750 128.115 94.970 128.985 ;
        RECT 95.150 128.675 95.500 129.045 ;
        RECT 95.670 128.495 95.840 129.225 ;
        RECT 96.010 129.165 96.420 129.605 ;
        RECT 96.710 128.965 96.960 129.395 ;
        RECT 97.160 129.145 97.480 129.605 ;
        RECT 98.040 129.215 98.890 129.385 ;
        RECT 96.010 128.625 96.420 128.955 ;
        RECT 96.710 128.625 97.130 128.965 ;
        RECT 95.420 128.455 95.840 128.495 ;
        RECT 95.420 128.285 96.770 128.455 ;
        RECT 93.830 127.725 94.525 127.895 ;
        RECT 94.750 127.735 95.250 128.115 ;
        RECT 93.855 127.055 94.185 127.555 ;
        RECT 94.355 127.225 94.525 127.725 ;
        RECT 95.420 127.440 95.590 128.285 ;
        RECT 96.520 128.125 96.770 128.285 ;
        RECT 95.760 127.855 96.010 128.115 ;
        RECT 96.940 127.855 97.130 128.625 ;
        RECT 95.760 127.605 97.130 127.855 ;
        RECT 97.300 128.795 98.550 128.965 ;
        RECT 97.300 128.035 97.470 128.795 ;
        RECT 98.220 128.675 98.550 128.795 ;
        RECT 97.640 128.215 97.820 128.625 ;
        RECT 98.720 128.455 98.890 129.215 ;
        RECT 99.090 129.125 99.750 129.605 ;
        RECT 99.930 129.010 100.250 129.340 ;
        RECT 99.080 128.685 99.740 128.955 ;
        RECT 99.080 128.625 99.410 128.685 ;
        RECT 99.560 128.455 99.890 128.515 ;
        RECT 97.990 128.285 99.890 128.455 ;
        RECT 97.300 127.725 97.820 128.035 ;
        RECT 97.990 127.775 98.160 128.285 ;
        RECT 100.060 128.115 100.250 129.010 ;
        RECT 98.330 127.945 100.250 128.115 ;
        RECT 99.930 127.925 100.250 127.945 ;
        RECT 100.450 128.695 100.700 129.345 ;
        RECT 100.880 129.145 101.165 129.605 ;
        RECT 101.345 129.265 101.600 129.425 ;
        RECT 101.345 129.095 101.685 129.265 ;
        RECT 102.145 129.095 102.450 129.605 ;
        RECT 101.345 128.895 101.600 129.095 ;
        RECT 100.450 128.365 101.250 128.695 ;
        RECT 97.990 127.605 99.200 127.775 ;
        RECT 94.760 127.270 95.590 127.440 ;
        RECT 95.830 127.055 96.210 127.435 ;
        RECT 96.390 127.315 96.560 127.605 ;
        RECT 97.990 127.525 98.160 127.605 ;
        RECT 96.730 127.055 97.060 127.435 ;
        RECT 97.530 127.275 98.160 127.525 ;
        RECT 98.340 127.055 98.760 127.435 ;
        RECT 98.960 127.315 99.200 127.605 ;
        RECT 99.430 127.055 99.760 127.745 ;
        RECT 99.930 127.315 100.100 127.925 ;
        RECT 100.450 127.775 100.700 128.365 ;
        RECT 101.420 128.035 101.600 128.895 ;
        RECT 102.145 128.365 102.460 128.925 ;
        RECT 102.630 128.615 102.880 129.425 ;
        RECT 103.050 129.080 103.310 129.605 ;
        RECT 103.490 128.615 103.740 129.425 ;
        RECT 103.910 129.045 104.170 129.605 ;
        RECT 104.340 128.955 104.600 129.410 ;
        RECT 104.770 129.125 105.030 129.605 ;
        RECT 105.200 128.955 105.460 129.410 ;
        RECT 105.630 129.125 105.890 129.605 ;
        RECT 106.060 128.955 106.320 129.410 ;
        RECT 106.490 129.125 106.735 129.605 ;
        RECT 106.905 128.955 107.180 129.410 ;
        RECT 107.350 129.125 107.595 129.605 ;
        RECT 107.765 128.955 108.025 129.410 ;
        RECT 108.205 129.125 108.455 129.605 ;
        RECT 108.625 128.955 108.885 129.410 ;
        RECT 109.065 129.125 109.315 129.605 ;
        RECT 109.485 128.955 109.745 129.410 ;
        RECT 109.925 129.125 110.185 129.605 ;
        RECT 110.355 128.955 110.615 129.410 ;
        RECT 110.785 129.125 111.085 129.605 ;
        RECT 111.545 128.975 111.875 129.335 ;
        RECT 112.495 129.145 112.745 129.605 ;
        RECT 112.915 129.145 113.475 129.435 ;
        RECT 104.340 128.785 111.085 128.955 ;
        RECT 111.545 128.785 112.935 128.975 ;
        RECT 102.630 128.365 109.750 128.615 ;
        RECT 100.370 127.265 100.700 127.775 ;
        RECT 100.880 127.055 101.165 127.855 ;
        RECT 101.345 127.365 101.600 128.035 ;
        RECT 102.155 127.055 102.450 127.865 ;
        RECT 102.630 127.225 102.875 128.365 ;
        RECT 103.050 127.055 103.310 127.865 ;
        RECT 103.490 127.230 103.740 128.365 ;
        RECT 109.920 128.195 111.085 128.785 ;
        RECT 112.765 128.695 112.935 128.785 ;
        RECT 104.340 127.970 111.085 128.195 ;
        RECT 111.360 128.365 112.035 128.615 ;
        RECT 112.255 128.365 112.595 128.615 ;
        RECT 112.765 128.365 113.055 128.695 ;
        RECT 111.360 128.005 111.625 128.365 ;
        RECT 112.765 128.115 112.935 128.365 ;
        RECT 104.340 127.955 109.745 127.970 ;
        RECT 103.910 127.060 104.170 127.855 ;
        RECT 104.340 127.230 104.600 127.955 ;
        RECT 104.770 127.060 105.030 127.785 ;
        RECT 105.200 127.230 105.460 127.955 ;
        RECT 105.630 127.060 105.890 127.785 ;
        RECT 106.060 127.230 106.320 127.955 ;
        RECT 106.490 127.060 106.750 127.785 ;
        RECT 106.920 127.230 107.180 127.955 ;
        RECT 107.350 127.060 107.595 127.785 ;
        RECT 107.765 127.230 108.025 127.955 ;
        RECT 108.210 127.060 108.455 127.785 ;
        RECT 108.625 127.230 108.885 127.955 ;
        RECT 109.070 127.060 109.315 127.785 ;
        RECT 109.485 127.230 109.745 127.955 ;
        RECT 109.930 127.060 110.185 127.785 ;
        RECT 110.355 127.230 110.645 127.970 ;
        RECT 111.995 127.945 112.935 128.115 ;
        RECT 103.910 127.055 110.185 127.060 ;
        RECT 110.815 127.055 111.085 127.800 ;
        RECT 111.545 127.055 111.825 127.725 ;
        RECT 111.995 127.395 112.295 127.945 ;
        RECT 113.225 127.775 113.475 129.145 ;
        RECT 114.565 128.880 114.855 129.605 ;
        RECT 115.860 128.925 116.115 129.425 ;
        RECT 116.295 129.145 116.580 129.605 ;
        RECT 115.775 128.895 116.115 128.925 ;
        RECT 115.775 128.755 116.040 128.895 ;
        RECT 112.495 127.055 112.825 127.775 ;
        RECT 113.015 127.225 113.475 127.775 ;
        RECT 114.565 127.055 114.855 128.220 ;
        RECT 115.860 128.035 116.040 128.755 ;
        RECT 116.760 128.695 117.010 129.345 ;
        RECT 116.210 128.365 117.010 128.695 ;
        RECT 115.860 127.365 116.115 128.035 ;
        RECT 116.295 127.055 116.580 127.855 ;
        RECT 116.760 127.775 117.010 128.365 ;
        RECT 117.210 129.010 117.530 129.340 ;
        RECT 117.710 129.125 118.370 129.605 ;
        RECT 118.570 129.215 119.420 129.385 ;
        RECT 117.210 128.115 117.400 129.010 ;
        RECT 117.720 128.685 118.380 128.955 ;
        RECT 118.050 128.625 118.380 128.685 ;
        RECT 117.570 128.455 117.900 128.515 ;
        RECT 118.570 128.455 118.740 129.215 ;
        RECT 119.980 129.145 120.300 129.605 ;
        RECT 120.500 128.965 120.750 129.395 ;
        RECT 121.040 129.165 121.450 129.605 ;
        RECT 121.620 129.225 122.635 129.425 ;
        RECT 118.910 128.795 120.160 128.965 ;
        RECT 118.910 128.675 119.240 128.795 ;
        RECT 117.570 128.285 119.470 128.455 ;
        RECT 117.210 127.945 119.130 128.115 ;
        RECT 117.210 127.925 117.530 127.945 ;
        RECT 116.760 127.265 117.090 127.775 ;
        RECT 117.360 127.315 117.530 127.925 ;
        RECT 119.300 127.775 119.470 128.285 ;
        RECT 119.640 128.215 119.820 128.625 ;
        RECT 119.990 128.035 120.160 128.795 ;
        RECT 117.700 127.055 118.030 127.745 ;
        RECT 118.260 127.605 119.470 127.775 ;
        RECT 119.640 127.725 120.160 128.035 ;
        RECT 120.330 128.625 120.750 128.965 ;
        RECT 121.040 128.625 121.450 128.955 ;
        RECT 120.330 127.855 120.520 128.625 ;
        RECT 121.620 128.495 121.790 129.225 ;
        RECT 122.935 129.055 123.105 129.385 ;
        RECT 123.275 129.225 123.605 129.605 ;
        RECT 121.960 128.675 122.310 129.045 ;
        RECT 121.620 128.455 122.040 128.495 ;
        RECT 120.690 128.285 122.040 128.455 ;
        RECT 120.690 128.125 120.940 128.285 ;
        RECT 121.450 127.855 121.700 128.115 ;
        RECT 120.330 127.605 121.700 127.855 ;
        RECT 118.260 127.315 118.500 127.605 ;
        RECT 119.300 127.525 119.470 127.605 ;
        RECT 118.700 127.055 119.120 127.435 ;
        RECT 119.300 127.275 119.930 127.525 ;
        RECT 120.400 127.055 120.730 127.435 ;
        RECT 120.900 127.315 121.070 127.605 ;
        RECT 121.870 127.440 122.040 128.285 ;
        RECT 122.490 128.115 122.710 128.985 ;
        RECT 122.935 128.865 123.630 129.055 ;
        RECT 122.210 127.735 122.710 128.115 ;
        RECT 122.880 128.065 123.290 128.685 ;
        RECT 123.460 127.895 123.630 128.865 ;
        RECT 122.935 127.725 123.630 127.895 ;
        RECT 121.250 127.055 121.630 127.435 ;
        RECT 121.870 127.270 122.700 127.440 ;
        RECT 122.935 127.225 123.105 127.725 ;
        RECT 123.275 127.055 123.605 127.555 ;
        RECT 123.820 127.225 124.045 129.345 ;
        RECT 124.215 129.225 124.545 129.605 ;
        RECT 124.715 129.055 124.885 129.345 ;
        RECT 124.220 128.885 124.885 129.055 ;
        RECT 124.220 127.895 124.450 128.885 ;
        RECT 125.145 128.855 126.355 129.605 ;
        RECT 126.525 128.855 127.735 129.605 ;
        RECT 124.620 128.065 124.970 128.715 ;
        RECT 125.145 128.145 125.665 128.685 ;
        RECT 125.835 128.315 126.355 128.855 ;
        RECT 126.525 128.145 127.045 128.685 ;
        RECT 127.215 128.315 127.735 128.855 ;
        RECT 124.220 127.725 124.885 127.895 ;
        RECT 124.215 127.055 124.545 127.555 ;
        RECT 124.715 127.225 124.885 127.725 ;
        RECT 125.145 127.055 126.355 128.145 ;
        RECT 126.525 127.055 127.735 128.145 ;
        RECT 20.640 126.885 127.820 127.055 ;
        RECT 20.725 125.795 21.935 126.885 ;
        RECT 20.725 125.085 21.245 125.625 ;
        RECT 21.415 125.255 21.935 125.795 ;
        RECT 23.085 125.745 23.295 126.885 ;
        RECT 23.465 125.735 23.795 126.715 ;
        RECT 23.965 125.745 24.195 126.885 ;
        RECT 20.725 124.335 21.935 125.085 ;
        RECT 23.085 124.335 23.295 125.155 ;
        RECT 23.465 125.135 23.715 125.735 ;
        RECT 24.405 125.720 24.695 126.885 ;
        RECT 24.905 125.745 25.135 126.885 ;
        RECT 25.305 125.735 25.635 126.715 ;
        RECT 25.805 125.745 26.015 126.885 ;
        RECT 26.335 125.955 26.505 126.715 ;
        RECT 26.685 126.125 27.015 126.885 ;
        RECT 26.335 125.785 27.000 125.955 ;
        RECT 27.185 125.810 27.455 126.715 ;
        RECT 23.885 125.325 24.215 125.575 ;
        RECT 24.885 125.325 25.215 125.575 ;
        RECT 23.465 124.505 23.795 125.135 ;
        RECT 23.965 124.335 24.195 125.155 ;
        RECT 24.405 124.335 24.695 125.060 ;
        RECT 24.905 124.335 25.135 125.155 ;
        RECT 25.385 125.135 25.635 125.735 ;
        RECT 26.830 125.640 27.000 125.785 ;
        RECT 26.265 125.235 26.595 125.605 ;
        RECT 26.830 125.310 27.115 125.640 ;
        RECT 25.305 124.505 25.635 125.135 ;
        RECT 25.805 124.335 26.015 125.155 ;
        RECT 26.830 125.055 27.000 125.310 ;
        RECT 26.335 124.885 27.000 125.055 ;
        RECT 27.285 125.010 27.455 125.810 ;
        RECT 26.335 124.505 26.505 124.885 ;
        RECT 26.685 124.335 27.015 124.715 ;
        RECT 27.195 124.505 27.455 125.010 ;
        RECT 27.630 125.745 27.965 126.715 ;
        RECT 28.135 125.745 28.305 126.885 ;
        RECT 28.475 126.545 30.505 126.715 ;
        RECT 27.630 125.075 27.800 125.745 ;
        RECT 28.475 125.575 28.645 126.545 ;
        RECT 27.970 125.245 28.225 125.575 ;
        RECT 28.450 125.245 28.645 125.575 ;
        RECT 28.815 126.205 29.940 126.375 ;
        RECT 28.055 125.075 28.225 125.245 ;
        RECT 28.815 125.075 28.985 126.205 ;
        RECT 27.630 124.505 27.885 125.075 ;
        RECT 28.055 124.905 28.985 125.075 ;
        RECT 29.155 125.865 30.165 126.035 ;
        RECT 29.155 125.065 29.325 125.865 ;
        RECT 28.810 124.870 28.985 124.905 ;
        RECT 28.055 124.335 28.385 124.735 ;
        RECT 28.810 124.505 29.340 124.870 ;
        RECT 29.530 124.845 29.805 125.665 ;
        RECT 29.525 124.675 29.805 124.845 ;
        RECT 29.530 124.505 29.805 124.675 ;
        RECT 29.975 124.505 30.165 125.865 ;
        RECT 30.335 125.880 30.505 126.545 ;
        RECT 30.675 126.125 30.845 126.885 ;
        RECT 33.060 126.545 33.315 126.575 ;
        RECT 31.080 126.125 31.595 126.535 ;
        RECT 32.975 126.375 33.315 126.545 ;
        RECT 30.335 125.690 31.085 125.880 ;
        RECT 31.255 125.315 31.595 126.125 ;
        RECT 30.365 125.145 31.595 125.315 ;
        RECT 33.060 125.905 33.315 126.375 ;
        RECT 33.495 126.085 33.780 126.885 ;
        RECT 33.960 126.165 34.290 126.675 ;
        RECT 30.345 124.335 30.855 124.870 ;
        RECT 31.075 124.540 31.320 125.145 ;
        RECT 33.060 125.045 33.240 125.905 ;
        RECT 33.960 125.575 34.210 126.165 ;
        RECT 34.560 126.015 34.730 126.625 ;
        RECT 34.900 126.195 35.230 126.885 ;
        RECT 35.460 126.335 35.700 126.625 ;
        RECT 35.900 126.505 36.320 126.885 ;
        RECT 36.500 126.415 37.130 126.665 ;
        RECT 37.600 126.505 37.930 126.885 ;
        RECT 36.500 126.335 36.670 126.415 ;
        RECT 38.100 126.335 38.270 126.625 ;
        RECT 38.450 126.505 38.830 126.885 ;
        RECT 39.070 126.500 39.900 126.670 ;
        RECT 35.460 126.165 36.670 126.335 ;
        RECT 33.410 125.245 34.210 125.575 ;
        RECT 33.060 124.515 33.315 125.045 ;
        RECT 33.495 124.335 33.780 124.795 ;
        RECT 33.960 124.595 34.210 125.245 ;
        RECT 34.410 125.995 34.730 126.015 ;
        RECT 34.410 125.825 36.330 125.995 ;
        RECT 34.410 124.930 34.600 125.825 ;
        RECT 36.500 125.655 36.670 126.165 ;
        RECT 36.840 125.905 37.360 126.215 ;
        RECT 34.770 125.485 36.670 125.655 ;
        RECT 34.770 125.425 35.100 125.485 ;
        RECT 35.250 125.255 35.580 125.315 ;
        RECT 34.920 124.985 35.580 125.255 ;
        RECT 34.410 124.600 34.730 124.930 ;
        RECT 34.910 124.335 35.570 124.815 ;
        RECT 35.770 124.725 35.940 125.485 ;
        RECT 36.840 125.315 37.020 125.725 ;
        RECT 36.110 125.145 36.440 125.265 ;
        RECT 37.190 125.145 37.360 125.905 ;
        RECT 36.110 124.975 37.360 125.145 ;
        RECT 37.530 126.085 38.900 126.335 ;
        RECT 37.530 125.315 37.720 126.085 ;
        RECT 38.650 125.825 38.900 126.085 ;
        RECT 37.890 125.655 38.140 125.815 ;
        RECT 39.070 125.655 39.240 126.500 ;
        RECT 40.135 126.215 40.305 126.715 ;
        RECT 40.475 126.385 40.805 126.885 ;
        RECT 39.410 125.825 39.910 126.205 ;
        RECT 40.135 126.045 40.830 126.215 ;
        RECT 37.890 125.485 39.240 125.655 ;
        RECT 38.820 125.445 39.240 125.485 ;
        RECT 37.530 124.975 37.950 125.315 ;
        RECT 38.240 124.985 38.650 125.315 ;
        RECT 35.770 124.555 36.620 124.725 ;
        RECT 37.180 124.335 37.500 124.795 ;
        RECT 37.700 124.545 37.950 124.975 ;
        RECT 38.240 124.335 38.650 124.775 ;
        RECT 38.820 124.715 38.990 125.445 ;
        RECT 39.160 124.895 39.510 125.265 ;
        RECT 39.690 124.955 39.910 125.825 ;
        RECT 40.080 125.255 40.490 125.875 ;
        RECT 40.660 125.075 40.830 126.045 ;
        RECT 40.135 124.885 40.830 125.075 ;
        RECT 38.820 124.515 39.835 124.715 ;
        RECT 40.135 124.555 40.305 124.885 ;
        RECT 40.475 124.335 40.805 124.715 ;
        RECT 41.020 124.595 41.245 126.715 ;
        RECT 41.415 126.385 41.745 126.885 ;
        RECT 41.915 126.215 42.085 126.715 ;
        RECT 41.420 126.045 42.085 126.215 ;
        RECT 42.805 126.125 43.320 126.535 ;
        RECT 43.555 126.125 43.725 126.885 ;
        RECT 43.895 126.545 45.925 126.715 ;
        RECT 41.420 125.055 41.650 126.045 ;
        RECT 41.820 125.225 42.170 125.875 ;
        RECT 42.805 125.315 43.145 126.125 ;
        RECT 43.895 125.880 44.065 126.545 ;
        RECT 44.460 126.205 45.585 126.375 ;
        RECT 43.315 125.690 44.065 125.880 ;
        RECT 44.235 125.865 45.245 126.035 ;
        RECT 42.805 125.145 44.035 125.315 ;
        RECT 41.420 124.885 42.085 125.055 ;
        RECT 41.415 124.335 41.745 124.715 ;
        RECT 41.915 124.595 42.085 124.885 ;
        RECT 43.080 124.540 43.325 125.145 ;
        RECT 43.545 124.335 44.055 124.870 ;
        RECT 44.235 124.505 44.425 125.865 ;
        RECT 44.595 124.845 44.870 125.665 ;
        RECT 45.075 125.065 45.245 125.865 ;
        RECT 45.415 125.075 45.585 126.205 ;
        RECT 45.755 125.575 45.925 126.545 ;
        RECT 46.095 125.745 46.265 126.885 ;
        RECT 46.435 125.745 46.770 126.715 ;
        RECT 45.755 125.245 45.950 125.575 ;
        RECT 46.175 125.245 46.430 125.575 ;
        RECT 46.175 125.075 46.345 125.245 ;
        RECT 46.600 125.075 46.770 125.745 ;
        RECT 47.405 125.795 49.995 126.885 ;
        RECT 47.405 125.275 48.615 125.795 ;
        RECT 50.165 125.720 50.455 126.885 ;
        RECT 50.625 126.125 51.140 126.535 ;
        RECT 51.375 126.125 51.545 126.885 ;
        RECT 51.715 126.545 53.745 126.715 ;
        RECT 48.785 125.105 49.995 125.625 ;
        RECT 50.625 125.315 50.965 126.125 ;
        RECT 51.715 125.880 51.885 126.545 ;
        RECT 52.280 126.205 53.405 126.375 ;
        RECT 51.135 125.690 51.885 125.880 ;
        RECT 52.055 125.865 53.065 126.035 ;
        RECT 50.625 125.145 51.855 125.315 ;
        RECT 45.415 124.905 46.345 125.075 ;
        RECT 45.415 124.870 45.590 124.905 ;
        RECT 44.595 124.675 44.875 124.845 ;
        RECT 44.595 124.505 44.870 124.675 ;
        RECT 45.060 124.505 45.590 124.870 ;
        RECT 46.015 124.335 46.345 124.735 ;
        RECT 46.515 124.505 46.770 125.075 ;
        RECT 47.405 124.335 49.995 125.105 ;
        RECT 50.165 124.335 50.455 125.060 ;
        RECT 50.900 124.540 51.145 125.145 ;
        RECT 51.365 124.335 51.875 124.870 ;
        RECT 52.055 124.505 52.245 125.865 ;
        RECT 52.415 124.845 52.690 125.665 ;
        RECT 52.895 125.065 53.065 125.865 ;
        RECT 53.235 125.075 53.405 126.205 ;
        RECT 53.575 125.575 53.745 126.545 ;
        RECT 53.915 125.745 54.085 126.885 ;
        RECT 54.255 125.745 54.590 126.715 ;
        RECT 55.690 126.450 61.035 126.885 ;
        RECT 53.575 125.245 53.770 125.575 ;
        RECT 53.995 125.245 54.250 125.575 ;
        RECT 53.995 125.075 54.165 125.245 ;
        RECT 54.420 125.075 54.590 125.745 ;
        RECT 57.280 125.200 57.630 126.450 ;
        RECT 61.205 126.125 61.720 126.535 ;
        RECT 61.955 126.125 62.125 126.885 ;
        RECT 62.295 126.545 64.325 126.715 ;
        RECT 53.235 124.905 54.165 125.075 ;
        RECT 53.235 124.870 53.410 124.905 ;
        RECT 52.415 124.675 52.695 124.845 ;
        RECT 52.415 124.505 52.690 124.675 ;
        RECT 52.880 124.505 53.410 124.870 ;
        RECT 53.835 124.335 54.165 124.735 ;
        RECT 54.335 124.505 54.590 125.075 ;
        RECT 59.110 124.880 59.450 125.710 ;
        RECT 61.205 125.315 61.545 126.125 ;
        RECT 62.295 125.880 62.465 126.545 ;
        RECT 62.860 126.205 63.985 126.375 ;
        RECT 61.715 125.690 62.465 125.880 ;
        RECT 62.635 125.865 63.645 126.035 ;
        RECT 61.205 125.145 62.435 125.315 ;
        RECT 55.690 124.335 61.035 124.880 ;
        RECT 61.480 124.540 61.725 125.145 ;
        RECT 61.945 124.335 62.455 124.870 ;
        RECT 62.635 124.505 62.825 125.865 ;
        RECT 62.995 125.525 63.270 125.665 ;
        RECT 62.995 125.355 63.275 125.525 ;
        RECT 62.995 124.505 63.270 125.355 ;
        RECT 63.475 125.065 63.645 125.865 ;
        RECT 63.815 125.075 63.985 126.205 ;
        RECT 64.155 125.575 64.325 126.545 ;
        RECT 64.495 125.745 64.665 126.885 ;
        RECT 64.835 125.745 65.170 126.715 ;
        RECT 64.155 125.245 64.350 125.575 ;
        RECT 64.575 125.245 64.830 125.575 ;
        RECT 64.575 125.075 64.745 125.245 ;
        RECT 65.000 125.075 65.170 125.745 ;
        RECT 65.345 125.795 66.555 126.885 ;
        RECT 66.725 126.125 67.240 126.535 ;
        RECT 67.475 126.125 67.645 126.885 ;
        RECT 67.815 126.545 69.845 126.715 ;
        RECT 65.345 125.255 65.865 125.795 ;
        RECT 66.035 125.085 66.555 125.625 ;
        RECT 66.725 125.315 67.065 126.125 ;
        RECT 67.815 125.880 67.985 126.545 ;
        RECT 68.380 126.205 69.505 126.375 ;
        RECT 67.235 125.690 67.985 125.880 ;
        RECT 68.155 125.865 69.165 126.035 ;
        RECT 66.725 125.145 67.955 125.315 ;
        RECT 63.815 124.905 64.745 125.075 ;
        RECT 63.815 124.870 63.990 124.905 ;
        RECT 63.460 124.505 63.990 124.870 ;
        RECT 64.415 124.335 64.745 124.735 ;
        RECT 64.915 124.505 65.170 125.075 ;
        RECT 65.345 124.335 66.555 125.085 ;
        RECT 67.000 124.540 67.245 125.145 ;
        RECT 67.465 124.335 67.975 124.870 ;
        RECT 68.155 124.505 68.345 125.865 ;
        RECT 68.515 124.845 68.790 125.665 ;
        RECT 68.995 125.065 69.165 125.865 ;
        RECT 69.335 125.075 69.505 126.205 ;
        RECT 69.675 125.575 69.845 126.545 ;
        RECT 70.015 125.745 70.185 126.885 ;
        RECT 70.355 125.745 70.690 126.715 ;
        RECT 70.925 125.745 71.135 126.885 ;
        RECT 69.675 125.245 69.870 125.575 ;
        RECT 70.095 125.245 70.350 125.575 ;
        RECT 70.095 125.075 70.265 125.245 ;
        RECT 70.520 125.075 70.690 125.745 ;
        RECT 71.305 125.735 71.635 126.715 ;
        RECT 71.805 125.745 72.035 126.885 ;
        RECT 72.795 125.955 72.965 126.715 ;
        RECT 73.145 126.125 73.475 126.885 ;
        RECT 72.795 125.785 73.460 125.955 ;
        RECT 73.645 125.810 73.915 126.715 ;
        RECT 69.335 124.905 70.265 125.075 ;
        RECT 69.335 124.870 69.510 124.905 ;
        RECT 68.515 124.675 68.795 124.845 ;
        RECT 68.515 124.505 68.790 124.675 ;
        RECT 68.980 124.505 69.510 124.870 ;
        RECT 69.935 124.335 70.265 124.735 ;
        RECT 70.435 124.505 70.690 125.075 ;
        RECT 70.925 124.335 71.135 125.155 ;
        RECT 71.305 125.135 71.555 125.735 ;
        RECT 73.290 125.640 73.460 125.785 ;
        RECT 71.725 125.325 72.055 125.575 ;
        RECT 72.725 125.235 73.055 125.605 ;
        RECT 73.290 125.310 73.575 125.640 ;
        RECT 71.305 124.505 71.635 125.135 ;
        RECT 71.805 124.335 72.035 125.155 ;
        RECT 73.290 125.055 73.460 125.310 ;
        RECT 72.795 124.885 73.460 125.055 ;
        RECT 73.745 125.010 73.915 125.810 ;
        RECT 74.635 125.955 74.805 126.715 ;
        RECT 74.985 126.125 75.315 126.885 ;
        RECT 74.635 125.785 75.300 125.955 ;
        RECT 75.485 125.810 75.755 126.715 ;
        RECT 75.130 125.640 75.300 125.785 ;
        RECT 74.565 125.235 74.895 125.605 ;
        RECT 75.130 125.310 75.415 125.640 ;
        RECT 75.130 125.055 75.300 125.310 ;
        RECT 72.795 124.505 72.965 124.885 ;
        RECT 73.145 124.335 73.475 124.715 ;
        RECT 73.655 124.505 73.915 125.010 ;
        RECT 74.635 124.885 75.300 125.055 ;
        RECT 75.585 125.010 75.755 125.810 ;
        RECT 75.925 125.720 76.215 126.885 ;
        RECT 77.345 125.745 77.575 126.885 ;
        RECT 77.745 125.735 78.075 126.715 ;
        RECT 78.245 125.745 78.455 126.885 ;
        RECT 79.060 126.545 79.315 126.575 ;
        RECT 78.975 126.375 79.315 126.545 ;
        RECT 79.060 125.905 79.315 126.375 ;
        RECT 79.495 126.085 79.780 126.885 ;
        RECT 79.960 126.165 80.290 126.675 ;
        RECT 77.325 125.325 77.655 125.575 ;
        RECT 74.635 124.505 74.805 124.885 ;
        RECT 74.985 124.335 75.315 124.715 ;
        RECT 75.495 124.505 75.755 125.010 ;
        RECT 75.925 124.335 76.215 125.060 ;
        RECT 77.345 124.335 77.575 125.155 ;
        RECT 77.825 125.135 78.075 125.735 ;
        RECT 77.745 124.505 78.075 125.135 ;
        RECT 78.245 124.335 78.455 125.155 ;
        RECT 79.060 125.045 79.240 125.905 ;
        RECT 79.960 125.575 80.210 126.165 ;
        RECT 80.560 126.015 80.730 126.625 ;
        RECT 80.900 126.195 81.230 126.885 ;
        RECT 81.460 126.335 81.700 126.625 ;
        RECT 81.900 126.505 82.320 126.885 ;
        RECT 82.500 126.415 83.130 126.665 ;
        RECT 83.600 126.505 83.930 126.885 ;
        RECT 82.500 126.335 82.670 126.415 ;
        RECT 84.100 126.335 84.270 126.625 ;
        RECT 84.450 126.505 84.830 126.885 ;
        RECT 85.070 126.500 85.900 126.670 ;
        RECT 81.460 126.165 82.670 126.335 ;
        RECT 79.410 125.245 80.210 125.575 ;
        RECT 79.060 124.515 79.315 125.045 ;
        RECT 79.495 124.335 79.780 124.795 ;
        RECT 79.960 124.595 80.210 125.245 ;
        RECT 80.410 125.995 80.730 126.015 ;
        RECT 80.410 125.825 82.330 125.995 ;
        RECT 80.410 124.930 80.600 125.825 ;
        RECT 82.500 125.655 82.670 126.165 ;
        RECT 82.840 125.905 83.360 126.215 ;
        RECT 80.770 125.485 82.670 125.655 ;
        RECT 80.770 125.425 81.100 125.485 ;
        RECT 81.250 125.255 81.580 125.315 ;
        RECT 80.920 124.985 81.580 125.255 ;
        RECT 80.410 124.600 80.730 124.930 ;
        RECT 80.910 124.335 81.570 124.815 ;
        RECT 81.770 124.725 81.940 125.485 ;
        RECT 82.840 125.315 83.020 125.725 ;
        RECT 82.110 125.145 82.440 125.265 ;
        RECT 83.190 125.145 83.360 125.905 ;
        RECT 82.110 124.975 83.360 125.145 ;
        RECT 83.530 126.085 84.900 126.335 ;
        RECT 83.530 125.315 83.720 126.085 ;
        RECT 84.650 125.825 84.900 126.085 ;
        RECT 83.890 125.655 84.140 125.815 ;
        RECT 85.070 125.655 85.240 126.500 ;
        RECT 86.135 126.215 86.305 126.715 ;
        RECT 86.475 126.385 86.805 126.885 ;
        RECT 85.410 125.825 85.910 126.205 ;
        RECT 86.135 126.045 86.830 126.215 ;
        RECT 83.890 125.485 85.240 125.655 ;
        RECT 84.820 125.445 85.240 125.485 ;
        RECT 83.530 124.975 83.950 125.315 ;
        RECT 84.240 124.985 84.650 125.315 ;
        RECT 81.770 124.555 82.620 124.725 ;
        RECT 83.180 124.335 83.500 124.795 ;
        RECT 83.700 124.545 83.950 124.975 ;
        RECT 84.240 124.335 84.650 124.775 ;
        RECT 84.820 124.715 84.990 125.445 ;
        RECT 85.160 124.895 85.510 125.265 ;
        RECT 85.690 124.955 85.910 125.825 ;
        RECT 86.080 125.255 86.490 125.875 ;
        RECT 86.660 125.075 86.830 126.045 ;
        RECT 86.135 124.885 86.830 125.075 ;
        RECT 84.820 124.515 85.835 124.715 ;
        RECT 86.135 124.555 86.305 124.885 ;
        RECT 86.475 124.335 86.805 124.715 ;
        RECT 87.020 124.595 87.245 126.715 ;
        RECT 87.415 126.385 87.745 126.885 ;
        RECT 87.915 126.215 88.085 126.715 ;
        RECT 87.420 126.045 88.085 126.215 ;
        RECT 87.420 125.055 87.650 126.045 ;
        RECT 87.820 125.225 88.170 125.875 ;
        RECT 89.305 125.745 89.535 126.885 ;
        RECT 89.705 125.735 90.035 126.715 ;
        RECT 90.205 125.745 90.415 126.885 ;
        RECT 90.650 125.745 90.985 126.715 ;
        RECT 91.155 125.745 91.325 126.885 ;
        RECT 91.495 126.545 93.525 126.715 ;
        RECT 89.285 125.325 89.615 125.575 ;
        RECT 87.420 124.885 88.085 125.055 ;
        RECT 87.415 124.335 87.745 124.715 ;
        RECT 87.915 124.595 88.085 124.885 ;
        RECT 89.305 124.335 89.535 125.155 ;
        RECT 89.785 125.135 90.035 125.735 ;
        RECT 89.705 124.505 90.035 125.135 ;
        RECT 90.205 124.335 90.415 125.155 ;
        RECT 90.650 125.075 90.820 125.745 ;
        RECT 91.495 125.575 91.665 126.545 ;
        RECT 90.990 125.245 91.245 125.575 ;
        RECT 91.470 125.245 91.665 125.575 ;
        RECT 91.835 126.205 92.960 126.375 ;
        RECT 91.075 125.075 91.245 125.245 ;
        RECT 91.835 125.075 92.005 126.205 ;
        RECT 90.650 124.505 90.905 125.075 ;
        RECT 91.075 124.905 92.005 125.075 ;
        RECT 92.175 125.865 93.185 126.035 ;
        RECT 92.175 125.065 92.345 125.865 ;
        RECT 92.550 125.185 92.825 125.665 ;
        RECT 92.545 125.015 92.825 125.185 ;
        RECT 91.830 124.870 92.005 124.905 ;
        RECT 91.075 124.335 91.405 124.735 ;
        RECT 91.830 124.505 92.360 124.870 ;
        RECT 92.550 124.505 92.825 125.015 ;
        RECT 92.995 124.505 93.185 125.865 ;
        RECT 93.355 125.880 93.525 126.545 ;
        RECT 93.695 126.125 93.865 126.885 ;
        RECT 94.100 126.125 94.615 126.535 ;
        RECT 93.355 125.690 94.105 125.880 ;
        RECT 94.275 125.315 94.615 126.125 ;
        RECT 93.385 125.145 94.615 125.315 ;
        RECT 94.785 125.795 97.375 126.885 ;
        RECT 97.545 126.125 98.060 126.535 ;
        RECT 98.295 126.125 98.465 126.885 ;
        RECT 98.635 126.545 100.665 126.715 ;
        RECT 94.785 125.275 95.995 125.795 ;
        RECT 93.365 124.335 93.875 124.870 ;
        RECT 94.095 124.540 94.340 125.145 ;
        RECT 96.165 125.105 97.375 125.625 ;
        RECT 97.545 125.315 97.885 126.125 ;
        RECT 98.635 125.880 98.805 126.545 ;
        RECT 99.200 126.205 100.325 126.375 ;
        RECT 98.055 125.690 98.805 125.880 ;
        RECT 98.975 125.865 99.985 126.035 ;
        RECT 97.545 125.145 98.775 125.315 ;
        RECT 94.785 124.335 97.375 125.105 ;
        RECT 97.820 124.540 98.065 125.145 ;
        RECT 98.285 124.335 98.795 124.870 ;
        RECT 98.975 124.505 99.165 125.865 ;
        RECT 99.335 124.845 99.610 125.665 ;
        RECT 99.815 125.065 99.985 125.865 ;
        RECT 100.155 125.075 100.325 126.205 ;
        RECT 100.495 125.575 100.665 126.545 ;
        RECT 100.835 125.745 101.005 126.885 ;
        RECT 101.175 125.745 101.510 126.715 ;
        RECT 100.495 125.245 100.690 125.575 ;
        RECT 100.915 125.245 101.170 125.575 ;
        RECT 100.915 125.075 101.085 125.245 ;
        RECT 101.340 125.075 101.510 125.745 ;
        RECT 101.685 125.720 101.975 126.885 ;
        RECT 102.145 126.165 102.605 126.715 ;
        RECT 102.795 126.165 103.125 126.885 ;
        RECT 100.155 124.905 101.085 125.075 ;
        RECT 100.155 124.870 100.330 124.905 ;
        RECT 99.335 124.675 99.615 124.845 ;
        RECT 99.335 124.505 99.610 124.675 ;
        RECT 99.800 124.505 100.330 124.870 ;
        RECT 100.755 124.335 101.085 124.735 ;
        RECT 101.255 124.505 101.510 125.075 ;
        RECT 101.685 124.335 101.975 125.060 ;
        RECT 102.145 124.795 102.395 126.165 ;
        RECT 103.325 125.995 103.625 126.545 ;
        RECT 103.795 126.215 104.075 126.885 ;
        RECT 102.685 125.825 103.625 125.995 ;
        RECT 102.685 125.575 102.855 125.825 ;
        RECT 103.995 125.575 104.260 125.935 ;
        RECT 104.485 125.745 104.715 126.885 ;
        RECT 104.885 125.735 105.215 126.715 ;
        RECT 105.385 125.745 105.595 126.885 ;
        RECT 106.285 126.125 106.800 126.535 ;
        RECT 107.035 126.125 107.205 126.885 ;
        RECT 107.375 126.545 109.405 126.715 ;
        RECT 102.565 125.245 102.855 125.575 ;
        RECT 103.025 125.325 103.365 125.575 ;
        RECT 103.585 125.325 104.260 125.575 ;
        RECT 104.465 125.325 104.795 125.575 ;
        RECT 102.685 125.155 102.855 125.245 ;
        RECT 102.685 124.965 104.075 125.155 ;
        RECT 102.145 124.505 102.705 124.795 ;
        RECT 102.875 124.335 103.125 124.795 ;
        RECT 103.745 124.605 104.075 124.965 ;
        RECT 104.485 124.335 104.715 125.155 ;
        RECT 104.965 125.135 105.215 125.735 ;
        RECT 106.285 125.315 106.625 126.125 ;
        RECT 107.375 125.880 107.545 126.545 ;
        RECT 107.940 126.205 109.065 126.375 ;
        RECT 106.795 125.690 107.545 125.880 ;
        RECT 107.715 125.865 108.725 126.035 ;
        RECT 104.885 124.505 105.215 125.135 ;
        RECT 105.385 124.335 105.595 125.155 ;
        RECT 106.285 125.145 107.515 125.315 ;
        RECT 106.560 124.540 106.805 125.145 ;
        RECT 107.025 124.335 107.535 124.870 ;
        RECT 107.715 124.505 107.905 125.865 ;
        RECT 108.075 125.525 108.350 125.665 ;
        RECT 108.075 125.355 108.355 125.525 ;
        RECT 108.075 124.505 108.350 125.355 ;
        RECT 108.555 125.065 108.725 125.865 ;
        RECT 108.895 125.075 109.065 126.205 ;
        RECT 109.235 125.575 109.405 126.545 ;
        RECT 109.575 125.745 109.745 126.885 ;
        RECT 109.915 125.745 110.250 126.715 ;
        RECT 109.235 125.245 109.430 125.575 ;
        RECT 109.655 125.245 109.910 125.575 ;
        RECT 109.655 125.075 109.825 125.245 ;
        RECT 110.080 125.075 110.250 125.745 ;
        RECT 110.885 126.125 111.400 126.535 ;
        RECT 111.635 126.125 111.805 126.885 ;
        RECT 111.975 126.545 114.005 126.715 ;
        RECT 110.885 125.315 111.225 126.125 ;
        RECT 111.975 125.880 112.145 126.545 ;
        RECT 112.540 126.205 113.665 126.375 ;
        RECT 111.395 125.690 112.145 125.880 ;
        RECT 112.315 125.865 113.325 126.035 ;
        RECT 110.885 125.145 112.115 125.315 ;
        RECT 108.895 124.905 109.825 125.075 ;
        RECT 108.895 124.870 109.070 124.905 ;
        RECT 108.540 124.505 109.070 124.870 ;
        RECT 109.495 124.335 109.825 124.735 ;
        RECT 109.995 124.505 110.250 125.075 ;
        RECT 111.160 124.540 111.405 125.145 ;
        RECT 111.625 124.335 112.135 124.870 ;
        RECT 112.315 124.505 112.505 125.865 ;
        RECT 112.675 125.525 112.950 125.665 ;
        RECT 112.675 125.355 112.955 125.525 ;
        RECT 112.675 124.505 112.950 125.355 ;
        RECT 113.155 125.065 113.325 125.865 ;
        RECT 113.495 125.075 113.665 126.205 ;
        RECT 113.835 125.575 114.005 126.545 ;
        RECT 114.175 125.745 114.345 126.885 ;
        RECT 114.515 125.745 114.850 126.715 ;
        RECT 113.835 125.245 114.030 125.575 ;
        RECT 114.255 125.245 114.510 125.575 ;
        RECT 114.255 125.075 114.425 125.245 ;
        RECT 114.680 125.075 114.850 125.745 ;
        RECT 115.400 125.905 115.655 126.575 ;
        RECT 115.835 126.085 116.120 126.885 ;
        RECT 116.300 126.165 116.630 126.675 ;
        RECT 115.400 125.525 115.580 125.905 ;
        RECT 116.300 125.575 116.550 126.165 ;
        RECT 116.900 126.015 117.070 126.625 ;
        RECT 117.240 126.195 117.570 126.885 ;
        RECT 117.800 126.335 118.040 126.625 ;
        RECT 118.240 126.505 118.660 126.885 ;
        RECT 118.840 126.415 119.470 126.665 ;
        RECT 119.940 126.505 120.270 126.885 ;
        RECT 118.840 126.335 119.010 126.415 ;
        RECT 120.440 126.335 120.610 126.625 ;
        RECT 120.790 126.505 121.170 126.885 ;
        RECT 121.410 126.500 122.240 126.670 ;
        RECT 117.800 126.165 119.010 126.335 ;
        RECT 115.315 125.355 115.580 125.525 ;
        RECT 113.495 124.905 114.425 125.075 ;
        RECT 113.495 124.870 113.670 124.905 ;
        RECT 113.140 124.505 113.670 124.870 ;
        RECT 114.095 124.335 114.425 124.735 ;
        RECT 114.595 124.505 114.850 125.075 ;
        RECT 115.400 125.045 115.580 125.355 ;
        RECT 115.750 125.245 116.550 125.575 ;
        RECT 115.400 124.515 115.655 125.045 ;
        RECT 115.835 124.335 116.120 124.795 ;
        RECT 116.300 124.595 116.550 125.245 ;
        RECT 116.750 125.995 117.070 126.015 ;
        RECT 116.750 125.825 118.670 125.995 ;
        RECT 116.750 124.930 116.940 125.825 ;
        RECT 118.840 125.655 119.010 126.165 ;
        RECT 119.180 125.905 119.700 126.215 ;
        RECT 117.110 125.485 119.010 125.655 ;
        RECT 117.110 125.425 117.440 125.485 ;
        RECT 117.590 125.255 117.920 125.315 ;
        RECT 117.260 124.985 117.920 125.255 ;
        RECT 116.750 124.600 117.070 124.930 ;
        RECT 117.250 124.335 117.910 124.815 ;
        RECT 118.110 124.725 118.280 125.485 ;
        RECT 119.180 125.315 119.360 125.725 ;
        RECT 118.450 125.145 118.780 125.265 ;
        RECT 119.530 125.145 119.700 125.905 ;
        RECT 118.450 124.975 119.700 125.145 ;
        RECT 119.870 126.085 121.240 126.335 ;
        RECT 119.870 125.315 120.060 126.085 ;
        RECT 120.990 125.825 121.240 126.085 ;
        RECT 120.230 125.655 120.480 125.815 ;
        RECT 121.410 125.655 121.580 126.500 ;
        RECT 122.475 126.215 122.645 126.715 ;
        RECT 122.815 126.385 123.145 126.885 ;
        RECT 121.750 125.825 122.250 126.205 ;
        RECT 122.475 126.045 123.170 126.215 ;
        RECT 120.230 125.485 121.580 125.655 ;
        RECT 121.160 125.445 121.580 125.485 ;
        RECT 119.870 124.975 120.290 125.315 ;
        RECT 120.580 124.985 120.990 125.315 ;
        RECT 118.110 124.555 118.960 124.725 ;
        RECT 119.520 124.335 119.840 124.795 ;
        RECT 120.040 124.545 120.290 124.975 ;
        RECT 120.580 124.335 120.990 124.775 ;
        RECT 121.160 124.715 121.330 125.445 ;
        RECT 121.500 124.895 121.850 125.265 ;
        RECT 122.030 124.955 122.250 125.825 ;
        RECT 122.420 125.255 122.830 125.875 ;
        RECT 123.000 125.075 123.170 126.045 ;
        RECT 122.475 124.885 123.170 125.075 ;
        RECT 121.160 124.515 122.175 124.715 ;
        RECT 122.475 124.555 122.645 124.885 ;
        RECT 122.815 124.335 123.145 124.715 ;
        RECT 123.360 124.595 123.585 126.715 ;
        RECT 123.755 126.385 124.085 126.885 ;
        RECT 124.255 126.215 124.425 126.715 ;
        RECT 123.760 126.045 124.425 126.215 ;
        RECT 123.760 125.055 123.990 126.045 ;
        RECT 124.160 125.225 124.510 125.875 ;
        RECT 124.685 125.810 124.955 126.715 ;
        RECT 125.125 126.125 125.455 126.885 ;
        RECT 125.635 125.955 125.805 126.715 ;
        RECT 123.760 124.885 124.425 125.055 ;
        RECT 123.755 124.335 124.085 124.715 ;
        RECT 124.255 124.595 124.425 124.885 ;
        RECT 124.685 125.010 124.855 125.810 ;
        RECT 125.140 125.785 125.805 125.955 ;
        RECT 126.525 125.795 127.735 126.885 ;
        RECT 125.140 125.640 125.310 125.785 ;
        RECT 125.025 125.310 125.310 125.640 ;
        RECT 125.140 125.055 125.310 125.310 ;
        RECT 125.545 125.235 125.875 125.605 ;
        RECT 126.525 125.255 127.045 125.795 ;
        RECT 127.215 125.085 127.735 125.625 ;
        RECT 124.685 124.505 124.945 125.010 ;
        RECT 125.140 124.885 125.805 125.055 ;
        RECT 125.125 124.335 125.455 124.715 ;
        RECT 125.635 124.505 125.805 124.885 ;
        RECT 126.525 124.335 127.735 125.085 ;
        RECT 20.640 124.165 127.820 124.335 ;
        RECT 20.725 123.415 21.935 124.165 ;
        RECT 22.940 123.825 23.195 123.985 ;
        RECT 22.855 123.655 23.195 123.825 ;
        RECT 23.375 123.705 23.660 124.165 ;
        RECT 22.940 123.455 23.195 123.655 ;
        RECT 20.725 122.875 21.245 123.415 ;
        RECT 21.415 122.705 21.935 123.245 ;
        RECT 20.725 121.615 21.935 122.705 ;
        RECT 22.940 122.595 23.120 123.455 ;
        RECT 23.840 123.255 24.090 123.905 ;
        RECT 23.290 122.925 24.090 123.255 ;
        RECT 22.940 121.925 23.195 122.595 ;
        RECT 23.375 121.615 23.660 122.415 ;
        RECT 23.840 122.335 24.090 122.925 ;
        RECT 24.290 123.570 24.610 123.900 ;
        RECT 24.790 123.685 25.450 124.165 ;
        RECT 25.650 123.775 26.500 123.945 ;
        RECT 24.290 122.675 24.480 123.570 ;
        RECT 24.800 123.245 25.460 123.515 ;
        RECT 25.130 123.185 25.460 123.245 ;
        RECT 24.650 123.015 24.980 123.075 ;
        RECT 25.650 123.015 25.820 123.775 ;
        RECT 27.060 123.705 27.380 124.165 ;
        RECT 27.580 123.525 27.830 123.955 ;
        RECT 28.120 123.725 28.530 124.165 ;
        RECT 28.700 123.785 29.715 123.985 ;
        RECT 25.990 123.355 27.240 123.525 ;
        RECT 25.990 123.235 26.320 123.355 ;
        RECT 24.650 122.845 26.550 123.015 ;
        RECT 24.290 122.505 26.210 122.675 ;
        RECT 24.290 122.485 24.610 122.505 ;
        RECT 23.840 121.825 24.170 122.335 ;
        RECT 24.440 121.875 24.610 122.485 ;
        RECT 26.380 122.335 26.550 122.845 ;
        RECT 26.720 122.775 26.900 123.185 ;
        RECT 27.070 122.595 27.240 123.355 ;
        RECT 24.780 121.615 25.110 122.305 ;
        RECT 25.340 122.165 26.550 122.335 ;
        RECT 26.720 122.285 27.240 122.595 ;
        RECT 27.410 123.185 27.830 123.525 ;
        RECT 28.120 123.185 28.530 123.515 ;
        RECT 27.410 122.415 27.600 123.185 ;
        RECT 28.700 123.055 28.870 123.785 ;
        RECT 30.015 123.615 30.185 123.945 ;
        RECT 30.355 123.785 30.685 124.165 ;
        RECT 29.040 123.235 29.390 123.605 ;
        RECT 28.700 123.015 29.120 123.055 ;
        RECT 27.770 122.845 29.120 123.015 ;
        RECT 27.770 122.685 28.020 122.845 ;
        RECT 28.530 122.415 28.780 122.675 ;
        RECT 27.410 122.165 28.780 122.415 ;
        RECT 25.340 121.875 25.580 122.165 ;
        RECT 26.380 122.085 26.550 122.165 ;
        RECT 25.780 121.615 26.200 121.995 ;
        RECT 26.380 121.835 27.010 122.085 ;
        RECT 27.480 121.615 27.810 121.995 ;
        RECT 27.980 121.875 28.150 122.165 ;
        RECT 28.950 122.000 29.120 122.845 ;
        RECT 29.570 122.675 29.790 123.545 ;
        RECT 30.015 123.425 30.710 123.615 ;
        RECT 29.290 122.295 29.790 122.675 ;
        RECT 29.960 122.625 30.370 123.245 ;
        RECT 30.540 122.455 30.710 123.425 ;
        RECT 30.015 122.285 30.710 122.455 ;
        RECT 28.330 121.615 28.710 121.995 ;
        RECT 28.950 121.830 29.780 122.000 ;
        RECT 30.015 121.785 30.185 122.285 ;
        RECT 30.355 121.615 30.685 122.115 ;
        RECT 30.900 121.785 31.125 123.905 ;
        RECT 31.295 123.785 31.625 124.165 ;
        RECT 31.795 123.615 31.965 123.905 ;
        RECT 31.300 123.445 31.965 123.615 ;
        RECT 31.300 122.455 31.530 123.445 ;
        RECT 33.420 123.355 33.665 123.960 ;
        RECT 33.885 123.630 34.395 124.165 ;
        RECT 31.700 122.625 32.050 123.275 ;
        RECT 33.145 123.185 34.375 123.355 ;
        RECT 31.300 122.285 31.965 122.455 ;
        RECT 31.295 121.615 31.625 122.115 ;
        RECT 31.795 121.785 31.965 122.285 ;
        RECT 33.145 122.375 33.485 123.185 ;
        RECT 33.655 122.620 34.405 122.810 ;
        RECT 33.145 121.965 33.660 122.375 ;
        RECT 33.895 121.615 34.065 122.375 ;
        RECT 34.235 121.955 34.405 122.620 ;
        RECT 34.575 122.635 34.765 123.995 ;
        RECT 34.935 123.485 35.210 123.995 ;
        RECT 35.400 123.630 35.930 123.995 ;
        RECT 36.355 123.765 36.685 124.165 ;
        RECT 35.755 123.595 35.930 123.630 ;
        RECT 34.935 123.315 35.215 123.485 ;
        RECT 34.935 122.835 35.210 123.315 ;
        RECT 35.415 122.635 35.585 123.435 ;
        RECT 34.575 122.465 35.585 122.635 ;
        RECT 35.755 123.425 36.685 123.595 ;
        RECT 36.855 123.425 37.110 123.995 ;
        RECT 37.285 123.440 37.575 124.165 ;
        RECT 37.835 123.615 38.005 123.995 ;
        RECT 38.185 123.785 38.515 124.165 ;
        RECT 37.835 123.445 38.500 123.615 ;
        RECT 38.695 123.490 38.955 123.995 ;
        RECT 35.755 122.295 35.925 123.425 ;
        RECT 36.515 123.255 36.685 123.425 ;
        RECT 34.800 122.125 35.925 122.295 ;
        RECT 36.095 122.925 36.290 123.255 ;
        RECT 36.515 122.925 36.770 123.255 ;
        RECT 36.095 121.955 36.265 122.925 ;
        RECT 36.940 122.755 37.110 123.425 ;
        RECT 37.765 122.895 38.095 123.265 ;
        RECT 38.330 123.190 38.500 123.445 ;
        RECT 38.330 122.860 38.615 123.190 ;
        RECT 34.235 121.785 36.265 121.955 ;
        RECT 36.435 121.615 36.605 122.755 ;
        RECT 36.775 121.785 37.110 122.755 ;
        RECT 37.285 121.615 37.575 122.780 ;
        RECT 38.330 122.715 38.500 122.860 ;
        RECT 37.835 122.545 38.500 122.715 ;
        RECT 38.785 122.690 38.955 123.490 ;
        RECT 37.835 121.785 38.005 122.545 ;
        RECT 38.185 121.615 38.515 122.375 ;
        RECT 38.685 121.785 38.955 122.690 ;
        RECT 39.500 123.455 39.755 123.985 ;
        RECT 39.935 123.705 40.220 124.165 ;
        RECT 39.500 122.595 39.680 123.455 ;
        RECT 40.400 123.255 40.650 123.905 ;
        RECT 39.850 122.925 40.650 123.255 ;
        RECT 39.500 122.125 39.755 122.595 ;
        RECT 39.415 121.955 39.755 122.125 ;
        RECT 39.500 121.925 39.755 121.955 ;
        RECT 39.935 121.615 40.220 122.415 ;
        RECT 40.400 122.335 40.650 122.925 ;
        RECT 40.850 123.570 41.170 123.900 ;
        RECT 41.350 123.685 42.010 124.165 ;
        RECT 42.210 123.775 43.060 123.945 ;
        RECT 40.850 122.675 41.040 123.570 ;
        RECT 41.360 123.245 42.020 123.515 ;
        RECT 41.690 123.185 42.020 123.245 ;
        RECT 41.210 123.015 41.540 123.075 ;
        RECT 42.210 123.015 42.380 123.775 ;
        RECT 43.620 123.705 43.940 124.165 ;
        RECT 44.140 123.525 44.390 123.955 ;
        RECT 44.680 123.725 45.090 124.165 ;
        RECT 45.260 123.785 46.275 123.985 ;
        RECT 42.550 123.355 43.800 123.525 ;
        RECT 42.550 123.235 42.880 123.355 ;
        RECT 41.210 122.845 43.110 123.015 ;
        RECT 40.850 122.505 42.770 122.675 ;
        RECT 40.850 122.485 41.170 122.505 ;
        RECT 40.400 121.825 40.730 122.335 ;
        RECT 41.000 121.875 41.170 122.485 ;
        RECT 42.940 122.335 43.110 122.845 ;
        RECT 43.280 122.775 43.460 123.185 ;
        RECT 43.630 122.595 43.800 123.355 ;
        RECT 41.340 121.615 41.670 122.305 ;
        RECT 41.900 122.165 43.110 122.335 ;
        RECT 43.280 122.285 43.800 122.595 ;
        RECT 43.970 123.185 44.390 123.525 ;
        RECT 44.680 123.185 45.090 123.515 ;
        RECT 43.970 122.415 44.160 123.185 ;
        RECT 45.260 123.055 45.430 123.785 ;
        RECT 46.575 123.615 46.745 123.945 ;
        RECT 46.915 123.785 47.245 124.165 ;
        RECT 45.600 123.235 45.950 123.605 ;
        RECT 45.260 123.015 45.680 123.055 ;
        RECT 44.330 122.845 45.680 123.015 ;
        RECT 44.330 122.685 44.580 122.845 ;
        RECT 45.090 122.415 45.340 122.675 ;
        RECT 43.970 122.165 45.340 122.415 ;
        RECT 41.900 121.875 42.140 122.165 ;
        RECT 42.940 122.085 43.110 122.165 ;
        RECT 42.340 121.615 42.760 121.995 ;
        RECT 42.940 121.835 43.570 122.085 ;
        RECT 44.040 121.615 44.370 121.995 ;
        RECT 44.540 121.875 44.710 122.165 ;
        RECT 45.510 122.000 45.680 122.845 ;
        RECT 46.130 122.675 46.350 123.545 ;
        RECT 46.575 123.425 47.270 123.615 ;
        RECT 45.850 122.295 46.350 122.675 ;
        RECT 46.520 122.625 46.930 123.245 ;
        RECT 47.100 122.455 47.270 123.425 ;
        RECT 46.575 122.285 47.270 122.455 ;
        RECT 44.890 121.615 45.270 121.995 ;
        RECT 45.510 121.830 46.340 122.000 ;
        RECT 46.575 121.785 46.745 122.285 ;
        RECT 46.915 121.615 47.245 122.115 ;
        RECT 47.460 121.785 47.685 123.905 ;
        RECT 47.855 123.785 48.185 124.165 ;
        RECT 48.355 123.615 48.525 123.905 ;
        RECT 49.160 123.825 49.415 123.985 ;
        RECT 49.075 123.655 49.415 123.825 ;
        RECT 49.595 123.705 49.880 124.165 ;
        RECT 47.860 123.445 48.525 123.615 ;
        RECT 49.160 123.455 49.415 123.655 ;
        RECT 47.860 122.455 48.090 123.445 ;
        RECT 48.260 122.625 48.610 123.275 ;
        RECT 49.160 122.595 49.340 123.455 ;
        RECT 50.060 123.255 50.310 123.905 ;
        RECT 49.510 122.925 50.310 123.255 ;
        RECT 47.860 122.285 48.525 122.455 ;
        RECT 47.855 121.615 48.185 122.115 ;
        RECT 48.355 121.785 48.525 122.285 ;
        RECT 49.160 121.925 49.415 122.595 ;
        RECT 49.595 121.615 49.880 122.415 ;
        RECT 50.060 122.335 50.310 122.925 ;
        RECT 50.510 123.570 50.830 123.900 ;
        RECT 51.010 123.685 51.670 124.165 ;
        RECT 51.870 123.775 52.720 123.945 ;
        RECT 50.510 122.675 50.700 123.570 ;
        RECT 51.020 123.245 51.680 123.515 ;
        RECT 51.350 123.185 51.680 123.245 ;
        RECT 50.870 123.015 51.200 123.075 ;
        RECT 51.870 123.015 52.040 123.775 ;
        RECT 53.280 123.705 53.600 124.165 ;
        RECT 53.800 123.525 54.050 123.955 ;
        RECT 54.340 123.725 54.750 124.165 ;
        RECT 54.920 123.785 55.935 123.985 ;
        RECT 52.210 123.355 53.460 123.525 ;
        RECT 52.210 123.235 52.540 123.355 ;
        RECT 50.870 122.845 52.770 123.015 ;
        RECT 50.510 122.505 52.430 122.675 ;
        RECT 50.510 122.485 50.830 122.505 ;
        RECT 50.060 121.825 50.390 122.335 ;
        RECT 50.660 121.875 50.830 122.485 ;
        RECT 52.600 122.335 52.770 122.845 ;
        RECT 52.940 122.775 53.120 123.185 ;
        RECT 53.290 122.595 53.460 123.355 ;
        RECT 51.000 121.615 51.330 122.305 ;
        RECT 51.560 122.165 52.770 122.335 ;
        RECT 52.940 122.285 53.460 122.595 ;
        RECT 53.630 123.185 54.050 123.525 ;
        RECT 54.340 123.185 54.750 123.515 ;
        RECT 53.630 122.415 53.820 123.185 ;
        RECT 54.920 123.055 55.090 123.785 ;
        RECT 56.235 123.615 56.405 123.945 ;
        RECT 56.575 123.785 56.905 124.165 ;
        RECT 55.260 123.235 55.610 123.605 ;
        RECT 54.920 123.015 55.340 123.055 ;
        RECT 53.990 122.845 55.340 123.015 ;
        RECT 53.990 122.685 54.240 122.845 ;
        RECT 54.750 122.415 55.000 122.675 ;
        RECT 53.630 122.165 55.000 122.415 ;
        RECT 51.560 121.875 51.800 122.165 ;
        RECT 52.600 122.085 52.770 122.165 ;
        RECT 52.000 121.615 52.420 121.995 ;
        RECT 52.600 121.835 53.230 122.085 ;
        RECT 53.700 121.615 54.030 121.995 ;
        RECT 54.200 121.875 54.370 122.165 ;
        RECT 55.170 122.000 55.340 122.845 ;
        RECT 55.790 122.675 56.010 123.545 ;
        RECT 56.235 123.425 56.930 123.615 ;
        RECT 55.510 122.295 56.010 122.675 ;
        RECT 56.180 122.625 56.590 123.245 ;
        RECT 56.760 122.455 56.930 123.425 ;
        RECT 56.235 122.285 56.930 122.455 ;
        RECT 54.550 121.615 54.930 121.995 ;
        RECT 55.170 121.830 56.000 122.000 ;
        RECT 56.235 121.785 56.405 122.285 ;
        RECT 56.575 121.615 56.905 122.115 ;
        RECT 57.120 121.785 57.345 123.905 ;
        RECT 57.515 123.785 57.845 124.165 ;
        RECT 58.015 123.615 58.185 123.905 ;
        RECT 57.520 123.445 58.185 123.615 ;
        RECT 57.520 122.455 57.750 123.445 ;
        RECT 58.905 123.395 61.495 124.165 ;
        RECT 57.920 122.625 58.270 123.275 ;
        RECT 58.905 122.705 60.115 123.225 ;
        RECT 60.285 122.875 61.495 123.395 ;
        RECT 61.705 123.345 61.935 124.165 ;
        RECT 62.105 123.365 62.435 123.995 ;
        RECT 61.685 122.925 62.015 123.175 ;
        RECT 62.185 122.765 62.435 123.365 ;
        RECT 62.605 123.345 62.815 124.165 ;
        RECT 63.045 123.440 63.335 124.165 ;
        RECT 64.425 123.490 64.685 123.995 ;
        RECT 64.865 123.785 65.195 124.165 ;
        RECT 65.375 123.615 65.545 123.995 ;
        RECT 66.180 123.825 66.435 123.985 ;
        RECT 66.095 123.655 66.435 123.825 ;
        RECT 66.615 123.705 66.900 124.165 ;
        RECT 57.520 122.285 58.185 122.455 ;
        RECT 57.515 121.615 57.845 122.115 ;
        RECT 58.015 121.785 58.185 122.285 ;
        RECT 58.905 121.615 61.495 122.705 ;
        RECT 61.705 121.615 61.935 122.755 ;
        RECT 62.105 121.785 62.435 122.765 ;
        RECT 62.605 121.615 62.815 122.755 ;
        RECT 63.045 121.615 63.335 122.780 ;
        RECT 64.425 122.690 64.595 123.490 ;
        RECT 64.880 123.445 65.545 123.615 ;
        RECT 66.180 123.455 66.435 123.655 ;
        RECT 64.880 123.190 65.050 123.445 ;
        RECT 64.765 122.860 65.050 123.190 ;
        RECT 65.285 122.895 65.615 123.265 ;
        RECT 64.880 122.715 65.050 122.860 ;
        RECT 64.425 121.785 64.695 122.690 ;
        RECT 64.880 122.545 65.545 122.715 ;
        RECT 64.865 121.615 65.195 122.375 ;
        RECT 65.375 121.785 65.545 122.545 ;
        RECT 66.180 122.595 66.360 123.455 ;
        RECT 67.080 123.255 67.330 123.905 ;
        RECT 66.530 122.925 67.330 123.255 ;
        RECT 66.180 121.925 66.435 122.595 ;
        RECT 66.615 121.615 66.900 122.415 ;
        RECT 67.080 122.335 67.330 122.925 ;
        RECT 67.530 123.570 67.850 123.900 ;
        RECT 68.030 123.685 68.690 124.165 ;
        RECT 68.890 123.775 69.740 123.945 ;
        RECT 67.530 122.675 67.720 123.570 ;
        RECT 68.040 123.245 68.700 123.515 ;
        RECT 68.370 123.185 68.700 123.245 ;
        RECT 67.890 123.015 68.220 123.075 ;
        RECT 68.890 123.015 69.060 123.775 ;
        RECT 70.300 123.705 70.620 124.165 ;
        RECT 70.820 123.525 71.070 123.955 ;
        RECT 71.360 123.725 71.770 124.165 ;
        RECT 71.940 123.785 72.955 123.985 ;
        RECT 69.230 123.355 70.480 123.525 ;
        RECT 69.230 123.235 69.560 123.355 ;
        RECT 67.890 122.845 69.790 123.015 ;
        RECT 67.530 122.505 69.450 122.675 ;
        RECT 67.530 122.485 67.850 122.505 ;
        RECT 67.080 121.825 67.410 122.335 ;
        RECT 67.680 121.875 67.850 122.485 ;
        RECT 69.620 122.335 69.790 122.845 ;
        RECT 69.960 122.775 70.140 123.185 ;
        RECT 70.310 122.595 70.480 123.355 ;
        RECT 68.020 121.615 68.350 122.305 ;
        RECT 68.580 122.165 69.790 122.335 ;
        RECT 69.960 122.285 70.480 122.595 ;
        RECT 70.650 123.185 71.070 123.525 ;
        RECT 71.360 123.185 71.770 123.515 ;
        RECT 70.650 122.415 70.840 123.185 ;
        RECT 71.940 123.055 72.110 123.785 ;
        RECT 73.255 123.615 73.425 123.945 ;
        RECT 73.595 123.785 73.925 124.165 ;
        RECT 72.280 123.235 72.630 123.605 ;
        RECT 71.940 123.015 72.360 123.055 ;
        RECT 71.010 122.845 72.360 123.015 ;
        RECT 71.010 122.685 71.260 122.845 ;
        RECT 71.770 122.415 72.020 122.675 ;
        RECT 70.650 122.165 72.020 122.415 ;
        RECT 68.580 121.875 68.820 122.165 ;
        RECT 69.620 122.085 69.790 122.165 ;
        RECT 69.020 121.615 69.440 121.995 ;
        RECT 69.620 121.835 70.250 122.085 ;
        RECT 70.720 121.615 71.050 121.995 ;
        RECT 71.220 121.875 71.390 122.165 ;
        RECT 72.190 122.000 72.360 122.845 ;
        RECT 72.810 122.675 73.030 123.545 ;
        RECT 73.255 123.425 73.950 123.615 ;
        RECT 72.530 122.295 73.030 122.675 ;
        RECT 73.200 122.625 73.610 123.245 ;
        RECT 73.780 122.455 73.950 123.425 ;
        RECT 73.255 122.285 73.950 122.455 ;
        RECT 71.570 121.615 71.950 121.995 ;
        RECT 72.190 121.830 73.020 122.000 ;
        RECT 73.255 121.785 73.425 122.285 ;
        RECT 73.595 121.615 73.925 122.115 ;
        RECT 74.140 121.785 74.365 123.905 ;
        RECT 74.535 123.785 74.865 124.165 ;
        RECT 75.035 123.615 75.205 123.905 ;
        RECT 74.540 123.445 75.205 123.615 ;
        RECT 76.015 123.615 76.185 123.905 ;
        RECT 76.355 123.785 76.685 124.165 ;
        RECT 76.015 123.445 76.680 123.615 ;
        RECT 74.540 122.455 74.770 123.445 ;
        RECT 74.940 122.625 75.290 123.275 ;
        RECT 75.930 122.625 76.280 123.275 ;
        RECT 76.450 122.455 76.680 123.445 ;
        RECT 74.540 122.285 75.205 122.455 ;
        RECT 74.535 121.615 74.865 122.115 ;
        RECT 75.035 121.785 75.205 122.285 ;
        RECT 76.015 122.285 76.680 122.455 ;
        RECT 76.015 121.785 76.185 122.285 ;
        RECT 76.355 121.615 76.685 122.115 ;
        RECT 76.855 121.785 77.080 123.905 ;
        RECT 77.295 123.785 77.625 124.165 ;
        RECT 77.795 123.615 77.965 123.945 ;
        RECT 78.265 123.785 79.280 123.985 ;
        RECT 77.270 123.425 77.965 123.615 ;
        RECT 77.270 122.455 77.440 123.425 ;
        RECT 77.610 122.625 78.020 123.245 ;
        RECT 78.190 122.675 78.410 123.545 ;
        RECT 78.590 123.235 78.940 123.605 ;
        RECT 79.110 123.055 79.280 123.785 ;
        RECT 79.450 123.725 79.860 124.165 ;
        RECT 80.150 123.525 80.400 123.955 ;
        RECT 80.600 123.705 80.920 124.165 ;
        RECT 81.480 123.775 82.330 123.945 ;
        RECT 79.450 123.185 79.860 123.515 ;
        RECT 80.150 123.185 80.570 123.525 ;
        RECT 78.860 123.015 79.280 123.055 ;
        RECT 78.860 122.845 80.210 123.015 ;
        RECT 77.270 122.285 77.965 122.455 ;
        RECT 78.190 122.295 78.690 122.675 ;
        RECT 77.295 121.615 77.625 122.115 ;
        RECT 77.795 121.785 77.965 122.285 ;
        RECT 78.860 122.000 79.030 122.845 ;
        RECT 79.960 122.685 80.210 122.845 ;
        RECT 79.200 122.415 79.450 122.675 ;
        RECT 80.380 122.415 80.570 123.185 ;
        RECT 79.200 122.165 80.570 122.415 ;
        RECT 80.740 123.355 81.990 123.525 ;
        RECT 80.740 122.595 80.910 123.355 ;
        RECT 81.660 123.235 81.990 123.355 ;
        RECT 81.080 122.775 81.260 123.185 ;
        RECT 82.160 123.015 82.330 123.775 ;
        RECT 82.530 123.685 83.190 124.165 ;
        RECT 83.370 123.570 83.690 123.900 ;
        RECT 82.520 123.245 83.180 123.515 ;
        RECT 82.520 123.185 82.850 123.245 ;
        RECT 83.000 123.015 83.330 123.075 ;
        RECT 81.430 122.845 83.330 123.015 ;
        RECT 80.740 122.285 81.260 122.595 ;
        RECT 81.430 122.335 81.600 122.845 ;
        RECT 83.500 122.675 83.690 123.570 ;
        RECT 81.770 122.505 83.690 122.675 ;
        RECT 83.370 122.485 83.690 122.505 ;
        RECT 83.890 123.255 84.140 123.905 ;
        RECT 84.320 123.705 84.605 124.165 ;
        RECT 84.785 123.825 85.040 123.985 ;
        RECT 84.785 123.655 85.125 123.825 ;
        RECT 84.785 123.455 85.040 123.655 ;
        RECT 83.890 122.925 84.690 123.255 ;
        RECT 81.430 122.165 82.640 122.335 ;
        RECT 78.200 121.830 79.030 122.000 ;
        RECT 79.270 121.615 79.650 121.995 ;
        RECT 79.830 121.875 80.000 122.165 ;
        RECT 81.430 122.085 81.600 122.165 ;
        RECT 80.170 121.615 80.500 121.995 ;
        RECT 80.970 121.835 81.600 122.085 ;
        RECT 81.780 121.615 82.200 121.995 ;
        RECT 82.400 121.875 82.640 122.165 ;
        RECT 82.870 121.615 83.200 122.305 ;
        RECT 83.370 121.875 83.540 122.485 ;
        RECT 83.890 122.335 84.140 122.925 ;
        RECT 84.860 122.595 85.040 123.455 ;
        RECT 85.645 123.345 85.855 124.165 ;
        RECT 86.025 123.365 86.355 123.995 ;
        RECT 86.025 122.765 86.275 123.365 ;
        RECT 86.525 123.345 86.755 124.165 ;
        RECT 86.965 123.490 87.225 123.995 ;
        RECT 87.405 123.785 87.735 124.165 ;
        RECT 87.915 123.615 88.085 123.995 ;
        RECT 86.445 122.925 86.775 123.175 ;
        RECT 83.810 121.825 84.140 122.335 ;
        RECT 84.320 121.615 84.605 122.415 ;
        RECT 84.785 121.925 85.040 122.595 ;
        RECT 85.645 121.615 85.855 122.755 ;
        RECT 86.025 121.785 86.355 122.765 ;
        RECT 86.525 121.615 86.755 122.755 ;
        RECT 86.965 122.690 87.135 123.490 ;
        RECT 87.420 123.445 88.085 123.615 ;
        RECT 87.420 123.190 87.590 123.445 ;
        RECT 88.805 123.440 89.095 124.165 ;
        RECT 89.305 123.345 89.535 124.165 ;
        RECT 89.705 123.365 90.035 123.995 ;
        RECT 87.305 122.860 87.590 123.190 ;
        RECT 87.825 122.895 88.155 123.265 ;
        RECT 89.285 122.925 89.615 123.175 ;
        RECT 87.420 122.715 87.590 122.860 ;
        RECT 86.965 121.785 87.235 122.690 ;
        RECT 87.420 122.545 88.085 122.715 ;
        RECT 87.405 121.615 87.735 122.375 ;
        RECT 87.915 121.785 88.085 122.545 ;
        RECT 88.805 121.615 89.095 122.780 ;
        RECT 89.785 122.765 90.035 123.365 ;
        RECT 90.205 123.345 90.415 124.165 ;
        RECT 90.735 123.615 90.905 123.995 ;
        RECT 91.085 123.785 91.415 124.165 ;
        RECT 90.735 123.445 91.400 123.615 ;
        RECT 91.595 123.490 91.855 123.995 ;
        RECT 92.400 123.825 92.655 123.985 ;
        RECT 92.315 123.655 92.655 123.825 ;
        RECT 92.835 123.705 93.120 124.165 ;
        RECT 90.665 122.895 90.995 123.265 ;
        RECT 91.230 123.190 91.400 123.445 ;
        RECT 89.305 121.615 89.535 122.755 ;
        RECT 89.705 121.785 90.035 122.765 ;
        RECT 91.230 122.860 91.515 123.190 ;
        RECT 90.205 121.615 90.415 122.755 ;
        RECT 91.230 122.715 91.400 122.860 ;
        RECT 90.735 122.545 91.400 122.715 ;
        RECT 91.685 122.690 91.855 123.490 ;
        RECT 90.735 121.785 90.905 122.545 ;
        RECT 91.085 121.615 91.415 122.375 ;
        RECT 91.585 121.785 91.855 122.690 ;
        RECT 92.400 123.455 92.655 123.655 ;
        RECT 92.400 122.595 92.580 123.455 ;
        RECT 93.300 123.255 93.550 123.905 ;
        RECT 92.750 122.925 93.550 123.255 ;
        RECT 92.400 121.925 92.655 122.595 ;
        RECT 92.835 121.615 93.120 122.415 ;
        RECT 93.300 122.335 93.550 122.925 ;
        RECT 93.750 123.570 94.070 123.900 ;
        RECT 94.250 123.685 94.910 124.165 ;
        RECT 95.110 123.775 95.960 123.945 ;
        RECT 93.750 122.675 93.940 123.570 ;
        RECT 94.260 123.245 94.920 123.515 ;
        RECT 94.590 123.185 94.920 123.245 ;
        RECT 94.110 123.015 94.440 123.075 ;
        RECT 95.110 123.015 95.280 123.775 ;
        RECT 96.520 123.705 96.840 124.165 ;
        RECT 97.040 123.525 97.290 123.955 ;
        RECT 97.580 123.725 97.990 124.165 ;
        RECT 98.160 123.785 99.175 123.985 ;
        RECT 95.450 123.355 96.700 123.525 ;
        RECT 95.450 123.235 95.780 123.355 ;
        RECT 94.110 122.845 96.010 123.015 ;
        RECT 93.750 122.505 95.670 122.675 ;
        RECT 93.750 122.485 94.070 122.505 ;
        RECT 93.300 121.825 93.630 122.335 ;
        RECT 93.900 121.875 94.070 122.485 ;
        RECT 95.840 122.335 96.010 122.845 ;
        RECT 96.180 122.775 96.360 123.185 ;
        RECT 96.530 122.595 96.700 123.355 ;
        RECT 94.240 121.615 94.570 122.305 ;
        RECT 94.800 122.165 96.010 122.335 ;
        RECT 96.180 122.285 96.700 122.595 ;
        RECT 96.870 123.185 97.290 123.525 ;
        RECT 97.580 123.185 97.990 123.515 ;
        RECT 96.870 122.415 97.060 123.185 ;
        RECT 98.160 123.055 98.330 123.785 ;
        RECT 99.475 123.615 99.645 123.945 ;
        RECT 99.815 123.785 100.145 124.165 ;
        RECT 98.500 123.235 98.850 123.605 ;
        RECT 98.160 123.015 98.580 123.055 ;
        RECT 97.230 122.845 98.580 123.015 ;
        RECT 97.230 122.685 97.480 122.845 ;
        RECT 97.990 122.415 98.240 122.675 ;
        RECT 96.870 122.165 98.240 122.415 ;
        RECT 94.800 121.875 95.040 122.165 ;
        RECT 95.840 122.085 96.010 122.165 ;
        RECT 95.240 121.615 95.660 121.995 ;
        RECT 95.840 121.835 96.470 122.085 ;
        RECT 96.940 121.615 97.270 121.995 ;
        RECT 97.440 121.875 97.610 122.165 ;
        RECT 98.410 122.000 98.580 122.845 ;
        RECT 99.030 122.675 99.250 123.545 ;
        RECT 99.475 123.425 100.170 123.615 ;
        RECT 98.750 122.295 99.250 122.675 ;
        RECT 99.420 122.625 99.830 123.245 ;
        RECT 100.000 122.455 100.170 123.425 ;
        RECT 99.475 122.285 100.170 122.455 ;
        RECT 97.790 121.615 98.170 121.995 ;
        RECT 98.410 121.830 99.240 122.000 ;
        RECT 99.475 121.785 99.645 122.285 ;
        RECT 99.815 121.615 100.145 122.115 ;
        RECT 100.360 121.785 100.585 123.905 ;
        RECT 100.755 123.785 101.085 124.165 ;
        RECT 101.255 123.615 101.425 123.905 ;
        RECT 100.760 123.445 101.425 123.615 ;
        RECT 102.060 123.455 102.315 123.985 ;
        RECT 102.495 123.705 102.780 124.165 ;
        RECT 100.760 122.455 100.990 123.445 ;
        RECT 101.160 122.625 101.510 123.275 ;
        RECT 102.060 122.805 102.240 123.455 ;
        RECT 102.960 123.255 103.210 123.905 ;
        RECT 102.410 122.925 103.210 123.255 ;
        RECT 101.975 122.635 102.240 122.805 ;
        RECT 102.060 122.595 102.240 122.635 ;
        RECT 100.760 122.285 101.425 122.455 ;
        RECT 100.755 121.615 101.085 122.115 ;
        RECT 101.255 121.785 101.425 122.285 ;
        RECT 102.060 121.925 102.315 122.595 ;
        RECT 102.495 121.615 102.780 122.415 ;
        RECT 102.960 122.335 103.210 122.925 ;
        RECT 103.410 123.570 103.730 123.900 ;
        RECT 103.910 123.685 104.570 124.165 ;
        RECT 104.770 123.775 105.620 123.945 ;
        RECT 103.410 122.675 103.600 123.570 ;
        RECT 103.920 123.245 104.580 123.515 ;
        RECT 104.250 123.185 104.580 123.245 ;
        RECT 103.770 123.015 104.100 123.075 ;
        RECT 104.770 123.015 104.940 123.775 ;
        RECT 106.180 123.705 106.500 124.165 ;
        RECT 106.700 123.525 106.950 123.955 ;
        RECT 107.240 123.725 107.650 124.165 ;
        RECT 107.820 123.785 108.835 123.985 ;
        RECT 105.110 123.355 106.360 123.525 ;
        RECT 105.110 123.235 105.440 123.355 ;
        RECT 103.770 122.845 105.670 123.015 ;
        RECT 103.410 122.505 105.330 122.675 ;
        RECT 103.410 122.485 103.730 122.505 ;
        RECT 102.960 121.825 103.290 122.335 ;
        RECT 103.560 121.875 103.730 122.485 ;
        RECT 105.500 122.335 105.670 122.845 ;
        RECT 105.840 122.775 106.020 123.185 ;
        RECT 106.190 122.595 106.360 123.355 ;
        RECT 103.900 121.615 104.230 122.305 ;
        RECT 104.460 122.165 105.670 122.335 ;
        RECT 105.840 122.285 106.360 122.595 ;
        RECT 106.530 123.185 106.950 123.525 ;
        RECT 107.240 123.185 107.650 123.515 ;
        RECT 106.530 122.415 106.720 123.185 ;
        RECT 107.820 123.055 107.990 123.785 ;
        RECT 109.135 123.615 109.305 123.945 ;
        RECT 109.475 123.785 109.805 124.165 ;
        RECT 108.160 123.235 108.510 123.605 ;
        RECT 107.820 123.015 108.240 123.055 ;
        RECT 106.890 122.845 108.240 123.015 ;
        RECT 106.890 122.685 107.140 122.845 ;
        RECT 107.650 122.415 107.900 122.675 ;
        RECT 106.530 122.165 107.900 122.415 ;
        RECT 104.460 121.875 104.700 122.165 ;
        RECT 105.500 122.085 105.670 122.165 ;
        RECT 104.900 121.615 105.320 121.995 ;
        RECT 105.500 121.835 106.130 122.085 ;
        RECT 106.600 121.615 106.930 121.995 ;
        RECT 107.100 121.875 107.270 122.165 ;
        RECT 108.070 122.000 108.240 122.845 ;
        RECT 108.690 122.675 108.910 123.545 ;
        RECT 109.135 123.425 109.830 123.615 ;
        RECT 108.410 122.295 108.910 122.675 ;
        RECT 109.080 122.625 109.490 123.245 ;
        RECT 109.660 122.455 109.830 123.425 ;
        RECT 109.135 122.285 109.830 122.455 ;
        RECT 107.450 121.615 107.830 121.995 ;
        RECT 108.070 121.830 108.900 122.000 ;
        RECT 109.135 121.785 109.305 122.285 ;
        RECT 109.475 121.615 109.805 122.115 ;
        RECT 110.020 121.785 110.245 123.905 ;
        RECT 110.415 123.785 110.745 124.165 ;
        RECT 110.915 123.615 111.085 123.905 ;
        RECT 110.420 123.445 111.085 123.615 ;
        RECT 111.345 123.490 111.605 123.995 ;
        RECT 111.785 123.785 112.115 124.165 ;
        RECT 112.295 123.615 112.465 123.995 ;
        RECT 110.420 122.455 110.650 123.445 ;
        RECT 110.820 122.625 111.170 123.275 ;
        RECT 111.345 122.690 111.515 123.490 ;
        RECT 111.800 123.445 112.465 123.615 ;
        RECT 111.800 123.190 111.970 123.445 ;
        RECT 112.785 123.345 112.995 124.165 ;
        RECT 113.165 123.365 113.495 123.995 ;
        RECT 111.685 122.860 111.970 123.190 ;
        RECT 112.205 122.895 112.535 123.265 ;
        RECT 111.800 122.715 111.970 122.860 ;
        RECT 113.165 122.765 113.415 123.365 ;
        RECT 113.665 123.345 113.895 124.165 ;
        RECT 114.565 123.440 114.855 124.165 ;
        RECT 115.030 123.425 115.285 123.995 ;
        RECT 115.455 123.765 115.785 124.165 ;
        RECT 116.210 123.630 116.740 123.995 ;
        RECT 116.210 123.595 116.385 123.630 ;
        RECT 115.455 123.425 116.385 123.595 ;
        RECT 113.585 122.925 113.915 123.175 ;
        RECT 110.420 122.285 111.085 122.455 ;
        RECT 110.415 121.615 110.745 122.115 ;
        RECT 110.915 121.785 111.085 122.285 ;
        RECT 111.345 121.785 111.615 122.690 ;
        RECT 111.800 122.545 112.465 122.715 ;
        RECT 111.785 121.615 112.115 122.375 ;
        RECT 112.295 121.785 112.465 122.545 ;
        RECT 112.785 121.615 112.995 122.755 ;
        RECT 113.165 121.785 113.495 122.765 ;
        RECT 113.665 121.615 113.895 122.755 ;
        RECT 114.565 121.615 114.855 122.780 ;
        RECT 115.030 122.755 115.200 123.425 ;
        RECT 115.455 123.255 115.625 123.425 ;
        RECT 115.370 122.925 115.625 123.255 ;
        RECT 115.850 122.925 116.045 123.255 ;
        RECT 115.030 121.785 115.365 122.755 ;
        RECT 115.535 121.615 115.705 122.755 ;
        RECT 115.875 121.955 116.045 122.925 ;
        RECT 116.215 122.295 116.385 123.425 ;
        RECT 116.555 122.635 116.725 123.435 ;
        RECT 116.930 123.145 117.205 123.995 ;
        RECT 116.925 122.975 117.205 123.145 ;
        RECT 116.930 122.835 117.205 122.975 ;
        RECT 117.375 122.635 117.565 123.995 ;
        RECT 117.745 123.630 118.255 124.165 ;
        RECT 118.475 123.355 118.720 123.960 ;
        RECT 117.765 123.185 118.995 123.355 ;
        RECT 119.205 123.345 119.435 124.165 ;
        RECT 119.605 123.365 119.935 123.995 ;
        RECT 116.555 122.465 117.565 122.635 ;
        RECT 117.735 122.620 118.485 122.810 ;
        RECT 116.215 122.125 117.340 122.295 ;
        RECT 117.735 121.955 117.905 122.620 ;
        RECT 118.655 122.375 118.995 123.185 ;
        RECT 119.185 122.925 119.515 123.175 ;
        RECT 119.685 122.765 119.935 123.365 ;
        RECT 120.105 123.345 120.315 124.165 ;
        RECT 121.010 123.620 126.355 124.165 ;
        RECT 115.875 121.785 117.905 121.955 ;
        RECT 118.075 121.615 118.245 122.375 ;
        RECT 118.480 121.965 118.995 122.375 ;
        RECT 119.205 121.615 119.435 122.755 ;
        RECT 119.605 121.785 119.935 122.765 ;
        RECT 120.105 121.615 120.315 122.755 ;
        RECT 122.600 122.050 122.950 123.300 ;
        RECT 124.430 122.790 124.770 123.620 ;
        RECT 126.525 123.415 127.735 124.165 ;
        RECT 126.525 122.705 127.045 123.245 ;
        RECT 127.215 122.875 127.735 123.415 ;
        RECT 121.010 121.615 126.355 122.050 ;
        RECT 126.525 121.615 127.735 122.705 ;
        RECT 20.640 121.445 127.820 121.615 ;
        RECT 20.725 120.355 21.935 121.445 ;
        RECT 20.725 119.645 21.245 120.185 ;
        RECT 21.415 119.815 21.935 120.355 ;
        RECT 22.565 120.355 24.235 121.445 ;
        RECT 22.565 119.835 23.315 120.355 ;
        RECT 24.405 120.280 24.695 121.445 ;
        RECT 25.240 121.105 25.495 121.135 ;
        RECT 25.155 120.935 25.495 121.105 ;
        RECT 25.240 120.465 25.495 120.935 ;
        RECT 25.675 120.645 25.960 121.445 ;
        RECT 26.140 120.725 26.470 121.235 ;
        RECT 23.485 119.665 24.235 120.185 ;
        RECT 20.725 118.895 21.935 119.645 ;
        RECT 22.565 118.895 24.235 119.665 ;
        RECT 24.405 118.895 24.695 119.620 ;
        RECT 25.240 119.605 25.420 120.465 ;
        RECT 26.140 120.135 26.390 120.725 ;
        RECT 26.740 120.575 26.910 121.185 ;
        RECT 27.080 120.755 27.410 121.445 ;
        RECT 27.640 120.895 27.880 121.185 ;
        RECT 28.080 121.065 28.500 121.445 ;
        RECT 28.680 120.975 29.310 121.225 ;
        RECT 29.780 121.065 30.110 121.445 ;
        RECT 28.680 120.895 28.850 120.975 ;
        RECT 30.280 120.895 30.450 121.185 ;
        RECT 30.630 121.065 31.010 121.445 ;
        RECT 31.250 121.060 32.080 121.230 ;
        RECT 27.640 120.725 28.850 120.895 ;
        RECT 25.590 119.805 26.390 120.135 ;
        RECT 25.240 119.075 25.495 119.605 ;
        RECT 25.675 118.895 25.960 119.355 ;
        RECT 26.140 119.155 26.390 119.805 ;
        RECT 26.590 120.555 26.910 120.575 ;
        RECT 26.590 120.385 28.510 120.555 ;
        RECT 26.590 119.490 26.780 120.385 ;
        RECT 28.680 120.215 28.850 120.725 ;
        RECT 29.020 120.465 29.540 120.775 ;
        RECT 26.950 120.045 28.850 120.215 ;
        RECT 26.950 119.985 27.280 120.045 ;
        RECT 27.430 119.815 27.760 119.875 ;
        RECT 27.100 119.545 27.760 119.815 ;
        RECT 26.590 119.160 26.910 119.490 ;
        RECT 27.090 118.895 27.750 119.375 ;
        RECT 27.950 119.285 28.120 120.045 ;
        RECT 29.020 119.875 29.200 120.285 ;
        RECT 28.290 119.705 28.620 119.825 ;
        RECT 29.370 119.705 29.540 120.465 ;
        RECT 28.290 119.535 29.540 119.705 ;
        RECT 29.710 120.645 31.080 120.895 ;
        RECT 29.710 119.875 29.900 120.645 ;
        RECT 30.830 120.385 31.080 120.645 ;
        RECT 30.070 120.215 30.320 120.375 ;
        RECT 31.250 120.215 31.420 121.060 ;
        RECT 32.315 120.775 32.485 121.275 ;
        RECT 32.655 120.945 32.985 121.445 ;
        RECT 31.590 120.385 32.090 120.765 ;
        RECT 32.315 120.605 33.010 120.775 ;
        RECT 30.070 120.045 31.420 120.215 ;
        RECT 31.000 120.005 31.420 120.045 ;
        RECT 29.710 119.535 30.130 119.875 ;
        RECT 30.420 119.545 30.830 119.875 ;
        RECT 27.950 119.115 28.800 119.285 ;
        RECT 29.360 118.895 29.680 119.355 ;
        RECT 29.880 119.105 30.130 119.535 ;
        RECT 30.420 118.895 30.830 119.335 ;
        RECT 31.000 119.275 31.170 120.005 ;
        RECT 31.340 119.455 31.690 119.825 ;
        RECT 31.870 119.515 32.090 120.385 ;
        RECT 32.260 119.815 32.670 120.435 ;
        RECT 32.840 119.635 33.010 120.605 ;
        RECT 32.315 119.445 33.010 119.635 ;
        RECT 31.000 119.075 32.015 119.275 ;
        RECT 32.315 119.115 32.485 119.445 ;
        RECT 32.655 118.895 32.985 119.275 ;
        RECT 33.200 119.155 33.425 121.275 ;
        RECT 33.595 120.945 33.925 121.445 ;
        RECT 34.095 120.775 34.265 121.275 ;
        RECT 33.600 120.605 34.265 120.775 ;
        RECT 33.600 119.615 33.830 120.605 ;
        RECT 34.000 119.785 34.350 120.435 ;
        RECT 34.525 120.355 35.735 121.445 ;
        RECT 34.525 119.815 35.045 120.355 ;
        RECT 35.945 120.305 36.175 121.445 ;
        RECT 36.345 120.295 36.675 121.275 ;
        RECT 36.845 120.305 37.055 121.445 ;
        RECT 37.290 121.010 42.635 121.445 ;
        RECT 35.215 119.645 35.735 120.185 ;
        RECT 35.925 119.885 36.255 120.135 ;
        RECT 33.600 119.445 34.265 119.615 ;
        RECT 33.595 118.895 33.925 119.275 ;
        RECT 34.095 119.155 34.265 119.445 ;
        RECT 34.525 118.895 35.735 119.645 ;
        RECT 35.945 118.895 36.175 119.715 ;
        RECT 36.425 119.695 36.675 120.295 ;
        RECT 38.880 119.760 39.230 121.010 ;
        RECT 42.865 120.305 43.075 121.445 ;
        RECT 43.245 120.295 43.575 121.275 ;
        RECT 43.745 120.305 43.975 121.445 ;
        RECT 44.185 120.355 45.855 121.445 ;
        RECT 46.115 120.515 46.285 121.275 ;
        RECT 46.465 120.685 46.795 121.445 ;
        RECT 36.345 119.065 36.675 119.695 ;
        RECT 36.845 118.895 37.055 119.715 ;
        RECT 40.710 119.440 41.050 120.270 ;
        RECT 37.290 118.895 42.635 119.440 ;
        RECT 42.865 118.895 43.075 119.715 ;
        RECT 43.245 119.695 43.495 120.295 ;
        RECT 43.665 119.885 43.995 120.135 ;
        RECT 44.185 119.835 44.935 120.355 ;
        RECT 46.115 120.345 46.780 120.515 ;
        RECT 46.965 120.370 47.235 121.275 ;
        RECT 46.610 120.200 46.780 120.345 ;
        RECT 43.245 119.065 43.575 119.695 ;
        RECT 43.745 118.895 43.975 119.715 ;
        RECT 45.105 119.665 45.855 120.185 ;
        RECT 46.045 119.795 46.375 120.165 ;
        RECT 46.610 119.870 46.895 120.200 ;
        RECT 44.185 118.895 45.855 119.665 ;
        RECT 46.610 119.615 46.780 119.870 ;
        RECT 46.115 119.445 46.780 119.615 ;
        RECT 47.065 119.570 47.235 120.370 ;
        RECT 47.405 120.355 49.995 121.445 ;
        RECT 47.405 119.835 48.615 120.355 ;
        RECT 50.165 120.280 50.455 121.445 ;
        RECT 50.625 120.355 52.295 121.445 ;
        RECT 48.785 119.665 49.995 120.185 ;
        RECT 50.625 119.835 51.375 120.355 ;
        RECT 52.525 120.305 52.735 121.445 ;
        RECT 52.905 120.295 53.235 121.275 ;
        RECT 53.405 120.305 53.635 121.445 ;
        RECT 54.855 120.515 55.025 121.275 ;
        RECT 55.205 120.685 55.535 121.445 ;
        RECT 54.855 120.345 55.520 120.515 ;
        RECT 55.705 120.370 55.975 121.275 ;
        RECT 51.545 119.665 52.295 120.185 ;
        RECT 46.115 119.065 46.285 119.445 ;
        RECT 46.465 118.895 46.795 119.275 ;
        RECT 46.975 119.065 47.235 119.570 ;
        RECT 47.405 118.895 49.995 119.665 ;
        RECT 50.165 118.895 50.455 119.620 ;
        RECT 50.625 118.895 52.295 119.665 ;
        RECT 52.525 118.895 52.735 119.715 ;
        RECT 52.905 119.695 53.155 120.295 ;
        RECT 55.350 120.200 55.520 120.345 ;
        RECT 53.325 119.885 53.655 120.135 ;
        RECT 54.785 119.795 55.115 120.165 ;
        RECT 55.350 119.870 55.635 120.200 ;
        RECT 52.905 119.065 53.235 119.695 ;
        RECT 53.405 118.895 53.635 119.715 ;
        RECT 55.350 119.615 55.520 119.870 ;
        RECT 54.855 119.445 55.520 119.615 ;
        RECT 55.805 119.570 55.975 120.370 ;
        RECT 56.755 120.295 57.085 121.445 ;
        RECT 57.255 120.425 57.425 121.275 ;
        RECT 57.595 120.645 57.925 121.445 ;
        RECT 58.095 120.425 58.265 121.275 ;
        RECT 58.445 120.645 58.685 121.445 ;
        RECT 58.855 120.465 59.185 121.275 ;
        RECT 59.915 120.775 60.085 121.275 ;
        RECT 60.255 120.945 60.585 121.445 ;
        RECT 59.915 120.605 60.580 120.775 ;
        RECT 57.255 120.255 58.265 120.425 ;
        RECT 58.470 120.295 59.185 120.465 ;
        RECT 57.255 119.715 57.750 120.255 ;
        RECT 58.470 120.055 58.640 120.295 ;
        RECT 58.140 119.885 58.640 120.055 ;
        RECT 58.810 119.885 59.190 120.125 ;
        RECT 58.470 119.715 58.640 119.885 ;
        RECT 59.830 119.785 60.180 120.435 ;
        RECT 54.855 119.065 55.025 119.445 ;
        RECT 55.205 118.895 55.535 119.275 ;
        RECT 55.715 119.065 55.975 119.570 ;
        RECT 56.755 118.895 57.085 119.695 ;
        RECT 57.255 119.545 58.265 119.715 ;
        RECT 58.470 119.545 59.105 119.715 ;
        RECT 60.350 119.615 60.580 120.605 ;
        RECT 57.255 119.065 57.425 119.545 ;
        RECT 57.595 118.895 57.925 119.375 ;
        RECT 58.095 119.065 58.265 119.545 ;
        RECT 58.515 118.895 58.755 119.375 ;
        RECT 58.935 119.065 59.105 119.545 ;
        RECT 59.915 119.445 60.580 119.615 ;
        RECT 59.915 119.155 60.085 119.445 ;
        RECT 60.255 118.895 60.585 119.275 ;
        RECT 60.755 119.155 60.980 121.275 ;
        RECT 61.195 120.945 61.525 121.445 ;
        RECT 61.695 120.775 61.865 121.275 ;
        RECT 62.100 121.060 62.930 121.230 ;
        RECT 63.170 121.065 63.550 121.445 ;
        RECT 61.170 120.605 61.865 120.775 ;
        RECT 61.170 119.635 61.340 120.605 ;
        RECT 61.510 119.815 61.920 120.435 ;
        RECT 62.090 120.385 62.590 120.765 ;
        RECT 61.170 119.445 61.865 119.635 ;
        RECT 62.090 119.515 62.310 120.385 ;
        RECT 62.760 120.215 62.930 121.060 ;
        RECT 63.730 120.895 63.900 121.185 ;
        RECT 64.070 121.065 64.400 121.445 ;
        RECT 64.870 120.975 65.500 121.225 ;
        RECT 65.680 121.065 66.100 121.445 ;
        RECT 65.330 120.895 65.500 120.975 ;
        RECT 66.300 120.895 66.540 121.185 ;
        RECT 63.100 120.645 64.470 120.895 ;
        RECT 63.100 120.385 63.350 120.645 ;
        RECT 63.860 120.215 64.110 120.375 ;
        RECT 62.760 120.045 64.110 120.215 ;
        RECT 62.760 120.005 63.180 120.045 ;
        RECT 62.490 119.455 62.840 119.825 ;
        RECT 61.195 118.895 61.525 119.275 ;
        RECT 61.695 119.115 61.865 119.445 ;
        RECT 63.010 119.275 63.180 120.005 ;
        RECT 64.280 119.875 64.470 120.645 ;
        RECT 63.350 119.545 63.760 119.875 ;
        RECT 64.050 119.535 64.470 119.875 ;
        RECT 64.640 120.465 65.160 120.775 ;
        RECT 65.330 120.725 66.540 120.895 ;
        RECT 66.770 120.755 67.100 121.445 ;
        RECT 64.640 119.705 64.810 120.465 ;
        RECT 64.980 119.875 65.160 120.285 ;
        RECT 65.330 120.215 65.500 120.725 ;
        RECT 67.270 120.575 67.440 121.185 ;
        RECT 67.710 120.725 68.040 121.235 ;
        RECT 67.270 120.555 67.590 120.575 ;
        RECT 65.670 120.385 67.590 120.555 ;
        RECT 65.330 120.045 67.230 120.215 ;
        RECT 65.560 119.705 65.890 119.825 ;
        RECT 64.640 119.535 65.890 119.705 ;
        RECT 62.165 119.075 63.180 119.275 ;
        RECT 63.350 118.895 63.760 119.335 ;
        RECT 64.050 119.105 64.300 119.535 ;
        RECT 64.500 118.895 64.820 119.355 ;
        RECT 66.060 119.285 66.230 120.045 ;
        RECT 66.900 119.985 67.230 120.045 ;
        RECT 66.420 119.815 66.750 119.875 ;
        RECT 66.420 119.545 67.080 119.815 ;
        RECT 67.400 119.490 67.590 120.385 ;
        RECT 65.380 119.115 66.230 119.285 ;
        RECT 66.430 118.895 67.090 119.375 ;
        RECT 67.270 119.160 67.590 119.490 ;
        RECT 67.790 120.135 68.040 120.725 ;
        RECT 68.220 120.645 68.505 121.445 ;
        RECT 68.685 121.105 68.940 121.135 ;
        RECT 68.685 120.935 69.025 121.105 ;
        RECT 68.685 120.465 68.940 120.935 ;
        RECT 67.790 119.805 68.590 120.135 ;
        RECT 67.790 119.155 68.040 119.805 ;
        RECT 68.760 119.605 68.940 120.465 ;
        RECT 69.545 120.305 69.755 121.445 ;
        RECT 69.925 120.295 70.255 121.275 ;
        RECT 70.425 120.305 70.655 121.445 ;
        RECT 71.415 120.515 71.585 121.275 ;
        RECT 71.765 120.685 72.095 121.445 ;
        RECT 71.415 120.345 72.080 120.515 ;
        RECT 72.265 120.370 72.535 121.275 ;
        RECT 68.220 118.895 68.505 119.355 ;
        RECT 68.685 119.075 68.940 119.605 ;
        RECT 69.545 118.895 69.755 119.715 ;
        RECT 69.925 119.695 70.175 120.295 ;
        RECT 71.910 120.200 72.080 120.345 ;
        RECT 70.345 119.885 70.675 120.135 ;
        RECT 71.345 119.795 71.675 120.165 ;
        RECT 71.910 119.870 72.195 120.200 ;
        RECT 69.925 119.065 70.255 119.695 ;
        RECT 70.425 118.895 70.655 119.715 ;
        RECT 71.910 119.615 72.080 119.870 ;
        RECT 71.415 119.445 72.080 119.615 ;
        RECT 72.365 119.570 72.535 120.370 ;
        RECT 73.165 120.355 75.755 121.445 ;
        RECT 73.165 119.835 74.375 120.355 ;
        RECT 75.925 120.280 76.215 121.445 ;
        RECT 76.390 121.010 81.735 121.445 ;
        RECT 74.545 119.665 75.755 120.185 ;
        RECT 77.980 119.760 78.330 121.010 ;
        RECT 81.905 120.685 82.420 121.095 ;
        RECT 82.655 120.685 82.825 121.445 ;
        RECT 82.995 121.105 85.025 121.275 ;
        RECT 71.415 119.065 71.585 119.445 ;
        RECT 71.765 118.895 72.095 119.275 ;
        RECT 72.275 119.065 72.535 119.570 ;
        RECT 73.165 118.895 75.755 119.665 ;
        RECT 75.925 118.895 76.215 119.620 ;
        RECT 79.810 119.440 80.150 120.270 ;
        RECT 81.905 119.875 82.245 120.685 ;
        RECT 82.995 120.440 83.165 121.105 ;
        RECT 83.560 120.765 84.685 120.935 ;
        RECT 82.415 120.250 83.165 120.440 ;
        RECT 83.335 120.425 84.345 120.595 ;
        RECT 81.905 119.705 83.135 119.875 ;
        RECT 76.390 118.895 81.735 119.440 ;
        RECT 82.180 119.100 82.425 119.705 ;
        RECT 82.645 118.895 83.155 119.430 ;
        RECT 83.335 119.065 83.525 120.425 ;
        RECT 83.695 120.085 83.970 120.225 ;
        RECT 83.695 119.915 83.975 120.085 ;
        RECT 83.695 119.065 83.970 119.915 ;
        RECT 84.175 119.625 84.345 120.425 ;
        RECT 84.515 119.635 84.685 120.765 ;
        RECT 84.855 120.135 85.025 121.105 ;
        RECT 85.195 120.305 85.365 121.445 ;
        RECT 85.535 120.305 85.870 121.275 ;
        RECT 86.420 120.465 86.675 121.135 ;
        RECT 86.855 120.645 87.140 121.445 ;
        RECT 87.320 120.725 87.650 121.235 ;
        RECT 86.420 120.425 86.600 120.465 ;
        RECT 84.855 119.805 85.050 120.135 ;
        RECT 85.275 119.805 85.530 120.135 ;
        RECT 85.275 119.635 85.445 119.805 ;
        RECT 85.700 119.635 85.870 120.305 ;
        RECT 86.335 120.255 86.600 120.425 ;
        RECT 84.515 119.465 85.445 119.635 ;
        RECT 84.515 119.430 84.690 119.465 ;
        RECT 84.160 119.065 84.690 119.430 ;
        RECT 85.115 118.895 85.445 119.295 ;
        RECT 85.615 119.065 85.870 119.635 ;
        RECT 86.420 119.605 86.600 120.255 ;
        RECT 87.320 120.135 87.570 120.725 ;
        RECT 87.920 120.575 88.090 121.185 ;
        RECT 88.260 120.755 88.590 121.445 ;
        RECT 88.820 120.895 89.060 121.185 ;
        RECT 89.260 121.065 89.680 121.445 ;
        RECT 89.860 120.975 90.490 121.225 ;
        RECT 90.960 121.065 91.290 121.445 ;
        RECT 89.860 120.895 90.030 120.975 ;
        RECT 91.460 120.895 91.630 121.185 ;
        RECT 91.810 121.065 92.190 121.445 ;
        RECT 92.430 121.060 93.260 121.230 ;
        RECT 88.820 120.725 90.030 120.895 ;
        RECT 86.770 119.805 87.570 120.135 ;
        RECT 86.420 119.075 86.675 119.605 ;
        RECT 86.855 118.895 87.140 119.355 ;
        RECT 87.320 119.155 87.570 119.805 ;
        RECT 87.770 120.555 88.090 120.575 ;
        RECT 87.770 120.385 89.690 120.555 ;
        RECT 87.770 119.490 87.960 120.385 ;
        RECT 89.860 120.215 90.030 120.725 ;
        RECT 90.200 120.465 90.720 120.775 ;
        RECT 88.130 120.045 90.030 120.215 ;
        RECT 88.130 119.985 88.460 120.045 ;
        RECT 88.610 119.815 88.940 119.875 ;
        RECT 88.280 119.545 88.940 119.815 ;
        RECT 87.770 119.160 88.090 119.490 ;
        RECT 88.270 118.895 88.930 119.375 ;
        RECT 89.130 119.285 89.300 120.045 ;
        RECT 90.200 119.875 90.380 120.285 ;
        RECT 89.470 119.705 89.800 119.825 ;
        RECT 90.550 119.705 90.720 120.465 ;
        RECT 89.470 119.535 90.720 119.705 ;
        RECT 90.890 120.645 92.260 120.895 ;
        RECT 90.890 119.875 91.080 120.645 ;
        RECT 92.010 120.385 92.260 120.645 ;
        RECT 91.250 120.215 91.500 120.375 ;
        RECT 92.430 120.215 92.600 121.060 ;
        RECT 93.495 120.775 93.665 121.275 ;
        RECT 93.835 120.945 94.165 121.445 ;
        RECT 92.770 120.385 93.270 120.765 ;
        RECT 93.495 120.605 94.190 120.775 ;
        RECT 91.250 120.045 92.600 120.215 ;
        RECT 92.180 120.005 92.600 120.045 ;
        RECT 90.890 119.535 91.310 119.875 ;
        RECT 91.600 119.545 92.010 119.875 ;
        RECT 89.130 119.115 89.980 119.285 ;
        RECT 90.540 118.895 90.860 119.355 ;
        RECT 91.060 119.105 91.310 119.535 ;
        RECT 91.600 118.895 92.010 119.335 ;
        RECT 92.180 119.275 92.350 120.005 ;
        RECT 92.520 119.455 92.870 119.825 ;
        RECT 93.050 119.515 93.270 120.385 ;
        RECT 93.440 119.815 93.850 120.435 ;
        RECT 94.020 119.635 94.190 120.605 ;
        RECT 93.495 119.445 94.190 119.635 ;
        RECT 92.180 119.075 93.195 119.275 ;
        RECT 93.495 119.115 93.665 119.445 ;
        RECT 93.835 118.895 94.165 119.275 ;
        RECT 94.380 119.155 94.605 121.275 ;
        RECT 94.775 120.945 95.105 121.445 ;
        RECT 95.275 120.775 95.445 121.275 ;
        RECT 94.780 120.605 95.445 120.775 ;
        RECT 94.780 119.615 95.010 120.605 ;
        RECT 95.180 119.785 95.530 120.435 ;
        RECT 96.625 120.355 100.135 121.445 ;
        RECT 100.305 120.370 100.575 121.275 ;
        RECT 100.745 120.685 101.075 121.445 ;
        RECT 101.255 120.515 101.425 121.275 ;
        RECT 96.625 119.835 98.315 120.355 ;
        RECT 98.485 119.665 100.135 120.185 ;
        RECT 94.780 119.445 95.445 119.615 ;
        RECT 94.775 118.895 95.105 119.275 ;
        RECT 95.275 119.155 95.445 119.445 ;
        RECT 96.625 118.895 100.135 119.665 ;
        RECT 100.305 119.570 100.475 120.370 ;
        RECT 100.760 120.345 101.425 120.515 ;
        RECT 100.760 120.200 100.930 120.345 ;
        RECT 101.685 120.280 101.975 121.445 ;
        RECT 102.610 121.010 107.955 121.445 ;
        RECT 108.500 121.105 108.755 121.135 ;
        RECT 100.645 119.870 100.930 120.200 ;
        RECT 100.760 119.615 100.930 119.870 ;
        RECT 101.165 119.795 101.495 120.165 ;
        RECT 104.200 119.760 104.550 121.010 ;
        RECT 108.415 120.935 108.755 121.105 ;
        RECT 108.500 120.465 108.755 120.935 ;
        RECT 108.935 120.645 109.220 121.445 ;
        RECT 109.400 120.725 109.730 121.235 ;
        RECT 100.305 119.065 100.565 119.570 ;
        RECT 100.760 119.445 101.425 119.615 ;
        RECT 100.745 118.895 101.075 119.275 ;
        RECT 101.255 119.065 101.425 119.445 ;
        RECT 101.685 118.895 101.975 119.620 ;
        RECT 106.030 119.440 106.370 120.270 ;
        RECT 108.500 119.605 108.680 120.465 ;
        RECT 109.400 120.135 109.650 120.725 ;
        RECT 110.000 120.575 110.170 121.185 ;
        RECT 110.340 120.755 110.670 121.445 ;
        RECT 110.900 120.895 111.140 121.185 ;
        RECT 111.340 121.065 111.760 121.445 ;
        RECT 111.940 120.975 112.570 121.225 ;
        RECT 113.040 121.065 113.370 121.445 ;
        RECT 111.940 120.895 112.110 120.975 ;
        RECT 113.540 120.895 113.710 121.185 ;
        RECT 113.890 121.065 114.270 121.445 ;
        RECT 114.510 121.060 115.340 121.230 ;
        RECT 110.900 120.725 112.110 120.895 ;
        RECT 108.850 119.805 109.650 120.135 ;
        RECT 102.610 118.895 107.955 119.440 ;
        RECT 108.500 119.075 108.755 119.605 ;
        RECT 108.935 118.895 109.220 119.355 ;
        RECT 109.400 119.155 109.650 119.805 ;
        RECT 109.850 120.555 110.170 120.575 ;
        RECT 109.850 120.385 111.770 120.555 ;
        RECT 109.850 119.490 110.040 120.385 ;
        RECT 111.940 120.215 112.110 120.725 ;
        RECT 112.280 120.465 112.800 120.775 ;
        RECT 110.210 120.045 112.110 120.215 ;
        RECT 110.210 119.985 110.540 120.045 ;
        RECT 110.690 119.815 111.020 119.875 ;
        RECT 110.360 119.545 111.020 119.815 ;
        RECT 109.850 119.160 110.170 119.490 ;
        RECT 110.350 118.895 111.010 119.375 ;
        RECT 111.210 119.285 111.380 120.045 ;
        RECT 112.280 119.875 112.460 120.285 ;
        RECT 111.550 119.705 111.880 119.825 ;
        RECT 112.630 119.705 112.800 120.465 ;
        RECT 111.550 119.535 112.800 119.705 ;
        RECT 112.970 120.645 114.340 120.895 ;
        RECT 112.970 119.875 113.160 120.645 ;
        RECT 114.090 120.385 114.340 120.645 ;
        RECT 113.330 120.215 113.580 120.375 ;
        RECT 114.510 120.215 114.680 121.060 ;
        RECT 115.575 120.775 115.745 121.275 ;
        RECT 115.915 120.945 116.245 121.445 ;
        RECT 114.850 120.385 115.350 120.765 ;
        RECT 115.575 120.605 116.270 120.775 ;
        RECT 113.330 120.045 114.680 120.215 ;
        RECT 114.260 120.005 114.680 120.045 ;
        RECT 112.970 119.535 113.390 119.875 ;
        RECT 113.680 119.545 114.090 119.875 ;
        RECT 111.210 119.115 112.060 119.285 ;
        RECT 112.620 118.895 112.940 119.355 ;
        RECT 113.140 119.105 113.390 119.535 ;
        RECT 113.680 118.895 114.090 119.335 ;
        RECT 114.260 119.275 114.430 120.005 ;
        RECT 114.600 119.455 114.950 119.825 ;
        RECT 115.130 119.515 115.350 120.385 ;
        RECT 115.520 119.815 115.930 120.435 ;
        RECT 116.100 119.635 116.270 120.605 ;
        RECT 115.575 119.445 116.270 119.635 ;
        RECT 114.260 119.075 115.275 119.275 ;
        RECT 115.575 119.115 115.745 119.445 ;
        RECT 115.915 118.895 116.245 119.275 ;
        RECT 116.460 119.155 116.685 121.275 ;
        RECT 116.855 120.945 117.185 121.445 ;
        RECT 117.355 120.775 117.525 121.275 ;
        RECT 116.860 120.605 117.525 120.775 ;
        RECT 116.860 119.615 117.090 120.605 ;
        RECT 117.260 119.785 117.610 120.435 ;
        RECT 118.245 120.355 120.835 121.445 ;
        RECT 121.010 121.010 126.355 121.445 ;
        RECT 118.245 119.835 119.455 120.355 ;
        RECT 119.625 119.665 120.835 120.185 ;
        RECT 122.600 119.760 122.950 121.010 ;
        RECT 126.525 120.355 127.735 121.445 ;
        RECT 116.860 119.445 117.525 119.615 ;
        RECT 116.855 118.895 117.185 119.275 ;
        RECT 117.355 119.155 117.525 119.445 ;
        RECT 118.245 118.895 120.835 119.665 ;
        RECT 124.430 119.440 124.770 120.270 ;
        RECT 126.525 119.815 127.045 120.355 ;
        RECT 127.215 119.645 127.735 120.185 ;
        RECT 121.010 118.895 126.355 119.440 ;
        RECT 126.525 118.895 127.735 119.645 ;
        RECT 20.640 118.725 127.820 118.895 ;
        RECT 20.725 117.975 21.935 118.725 ;
        RECT 20.725 117.435 21.245 117.975 ;
        RECT 22.105 117.955 25.615 118.725 ;
        RECT 25.790 118.180 31.135 118.725 ;
        RECT 21.415 117.265 21.935 117.805 ;
        RECT 20.725 116.175 21.935 117.265 ;
        RECT 22.105 117.265 23.795 117.785 ;
        RECT 23.965 117.435 25.615 117.955 ;
        RECT 22.105 116.175 25.615 117.265 ;
        RECT 27.380 116.610 27.730 117.860 ;
        RECT 29.210 117.350 29.550 118.180 ;
        RECT 31.395 118.175 31.565 118.555 ;
        RECT 31.745 118.345 32.075 118.725 ;
        RECT 31.395 118.005 32.060 118.175 ;
        RECT 32.255 118.050 32.515 118.555 ;
        RECT 31.325 117.455 31.655 117.825 ;
        RECT 31.890 117.750 32.060 118.005 ;
        RECT 31.890 117.420 32.175 117.750 ;
        RECT 31.890 117.275 32.060 117.420 ;
        RECT 31.395 117.105 32.060 117.275 ;
        RECT 32.345 117.250 32.515 118.050 ;
        RECT 33.605 117.955 37.115 118.725 ;
        RECT 37.285 118.000 37.575 118.725 ;
        RECT 38.205 117.955 40.795 118.725 ;
        RECT 40.970 118.180 46.315 118.725 ;
        RECT 46.490 118.180 51.835 118.725 ;
        RECT 52.010 118.180 57.355 118.725 ;
        RECT 57.530 118.180 62.875 118.725 ;
        RECT 25.790 116.175 31.135 116.610 ;
        RECT 31.395 116.345 31.565 117.105 ;
        RECT 31.745 116.175 32.075 116.935 ;
        RECT 32.245 116.345 32.515 117.250 ;
        RECT 33.605 117.265 35.295 117.785 ;
        RECT 35.465 117.435 37.115 117.955 ;
        RECT 33.605 116.175 37.115 117.265 ;
        RECT 37.285 116.175 37.575 117.340 ;
        RECT 38.205 117.265 39.415 117.785 ;
        RECT 39.585 117.435 40.795 117.955 ;
        RECT 38.205 116.175 40.795 117.265 ;
        RECT 42.560 116.610 42.910 117.860 ;
        RECT 44.390 117.350 44.730 118.180 ;
        RECT 48.080 116.610 48.430 117.860 ;
        RECT 49.910 117.350 50.250 118.180 ;
        RECT 53.600 116.610 53.950 117.860 ;
        RECT 55.430 117.350 55.770 118.180 ;
        RECT 59.120 116.610 59.470 117.860 ;
        RECT 60.950 117.350 61.290 118.180 ;
        RECT 63.045 118.000 63.335 118.725 ;
        RECT 63.965 117.955 66.555 118.725 ;
        RECT 66.730 118.180 72.075 118.725 ;
        RECT 72.250 118.180 77.595 118.725 ;
        RECT 77.770 118.180 83.115 118.725 ;
        RECT 83.290 118.180 88.635 118.725 ;
        RECT 40.970 116.175 46.315 116.610 ;
        RECT 46.490 116.175 51.835 116.610 ;
        RECT 52.010 116.175 57.355 116.610 ;
        RECT 57.530 116.175 62.875 116.610 ;
        RECT 63.045 116.175 63.335 117.340 ;
        RECT 63.965 117.265 65.175 117.785 ;
        RECT 65.345 117.435 66.555 117.955 ;
        RECT 63.965 116.175 66.555 117.265 ;
        RECT 68.320 116.610 68.670 117.860 ;
        RECT 70.150 117.350 70.490 118.180 ;
        RECT 73.840 116.610 74.190 117.860 ;
        RECT 75.670 117.350 76.010 118.180 ;
        RECT 79.360 116.610 79.710 117.860 ;
        RECT 81.190 117.350 81.530 118.180 ;
        RECT 84.880 116.610 85.230 117.860 ;
        RECT 86.710 117.350 87.050 118.180 ;
        RECT 88.805 118.000 89.095 118.725 ;
        RECT 89.725 117.955 92.315 118.725 ;
        RECT 92.490 118.180 97.835 118.725 ;
        RECT 98.010 118.180 103.355 118.725 ;
        RECT 103.530 118.180 108.875 118.725 ;
        RECT 109.050 118.180 114.395 118.725 ;
        RECT 66.730 116.175 72.075 116.610 ;
        RECT 72.250 116.175 77.595 116.610 ;
        RECT 77.770 116.175 83.115 116.610 ;
        RECT 83.290 116.175 88.635 116.610 ;
        RECT 88.805 116.175 89.095 117.340 ;
        RECT 89.725 117.265 90.935 117.785 ;
        RECT 91.105 117.435 92.315 117.955 ;
        RECT 89.725 116.175 92.315 117.265 ;
        RECT 94.080 116.610 94.430 117.860 ;
        RECT 95.910 117.350 96.250 118.180 ;
        RECT 99.600 116.610 99.950 117.860 ;
        RECT 101.430 117.350 101.770 118.180 ;
        RECT 105.120 116.610 105.470 117.860 ;
        RECT 106.950 117.350 107.290 118.180 ;
        RECT 110.640 116.610 110.990 117.860 ;
        RECT 112.470 117.350 112.810 118.180 ;
        RECT 114.565 118.000 114.855 118.725 ;
        RECT 115.115 118.175 115.285 118.555 ;
        RECT 115.465 118.345 115.795 118.725 ;
        RECT 115.115 118.005 115.780 118.175 ;
        RECT 115.975 118.050 116.235 118.555 ;
        RECT 115.045 117.455 115.375 117.825 ;
        RECT 115.610 117.750 115.780 118.005 ;
        RECT 115.610 117.420 115.895 117.750 ;
        RECT 92.490 116.175 97.835 116.610 ;
        RECT 98.010 116.175 103.355 116.610 ;
        RECT 103.530 116.175 108.875 116.610 ;
        RECT 109.050 116.175 114.395 116.610 ;
        RECT 114.565 116.175 114.855 117.340 ;
        RECT 115.610 117.275 115.780 117.420 ;
        RECT 115.115 117.105 115.780 117.275 ;
        RECT 116.065 117.250 116.235 118.050 ;
        RECT 116.865 117.955 119.455 118.725 ;
        RECT 115.115 116.345 115.285 117.105 ;
        RECT 115.465 116.175 115.795 116.935 ;
        RECT 115.965 116.345 116.235 117.250 ;
        RECT 116.865 117.265 118.075 117.785 ;
        RECT 118.245 117.435 119.455 117.955 ;
        RECT 119.665 117.905 119.895 118.725 ;
        RECT 120.065 117.925 120.395 118.555 ;
        RECT 119.645 117.485 119.975 117.735 ;
        RECT 120.145 117.325 120.395 117.925 ;
        RECT 120.565 117.905 120.775 118.725 ;
        RECT 121.095 118.175 121.265 118.555 ;
        RECT 121.445 118.345 121.775 118.725 ;
        RECT 121.095 118.005 121.760 118.175 ;
        RECT 121.955 118.050 122.215 118.555 ;
        RECT 121.025 117.455 121.355 117.825 ;
        RECT 121.590 117.750 121.760 118.005 ;
        RECT 116.865 116.175 119.455 117.265 ;
        RECT 119.665 116.175 119.895 117.315 ;
        RECT 120.065 116.345 120.395 117.325 ;
        RECT 121.590 117.420 121.875 117.750 ;
        RECT 120.565 116.175 120.775 117.315 ;
        RECT 121.590 117.275 121.760 117.420 ;
        RECT 121.095 117.105 121.760 117.275 ;
        RECT 122.045 117.250 122.215 118.050 ;
        RECT 121.095 116.345 121.265 117.105 ;
        RECT 121.445 116.175 121.775 116.935 ;
        RECT 121.945 116.345 122.215 117.250 ;
        RECT 122.385 118.050 122.645 118.555 ;
        RECT 122.825 118.345 123.155 118.725 ;
        RECT 123.335 118.175 123.505 118.555 ;
        RECT 122.385 117.250 122.555 118.050 ;
        RECT 122.840 118.005 123.505 118.175 ;
        RECT 122.840 117.750 123.010 118.005 ;
        RECT 123.765 117.955 126.355 118.725 ;
        RECT 126.525 117.975 127.735 118.725 ;
        RECT 122.725 117.420 123.010 117.750 ;
        RECT 123.245 117.455 123.575 117.825 ;
        RECT 122.840 117.275 123.010 117.420 ;
        RECT 122.385 116.345 122.655 117.250 ;
        RECT 122.840 117.105 123.505 117.275 ;
        RECT 122.825 116.175 123.155 116.935 ;
        RECT 123.335 116.345 123.505 117.105 ;
        RECT 123.765 117.265 124.975 117.785 ;
        RECT 125.145 117.435 126.355 117.955 ;
        RECT 126.525 117.265 127.045 117.805 ;
        RECT 127.215 117.435 127.735 117.975 ;
        RECT 123.765 116.175 126.355 117.265 ;
        RECT 126.525 116.175 127.735 117.265 ;
        RECT 20.640 116.005 127.820 116.175 ;
        RECT 20.725 114.915 21.935 116.005 ;
        RECT 20.725 114.205 21.245 114.745 ;
        RECT 21.415 114.375 21.935 114.915 ;
        RECT 22.565 114.915 24.235 116.005 ;
        RECT 22.565 114.395 23.315 114.915 ;
        RECT 24.405 114.840 24.695 116.005 ;
        RECT 24.865 114.915 26.535 116.005 ;
        RECT 23.485 114.225 24.235 114.745 ;
        RECT 24.865 114.395 25.615 114.915 ;
        RECT 26.710 114.815 26.965 115.695 ;
        RECT 27.135 114.865 27.440 116.005 ;
        RECT 27.780 115.625 28.110 116.005 ;
        RECT 28.290 115.455 28.460 115.745 ;
        RECT 28.630 115.545 28.880 116.005 ;
        RECT 27.660 115.285 28.460 115.455 ;
        RECT 29.050 115.495 29.920 115.835 ;
        RECT 25.785 114.225 26.535 114.745 ;
        RECT 20.725 113.455 21.935 114.205 ;
        RECT 22.565 113.455 24.235 114.225 ;
        RECT 24.405 113.455 24.695 114.180 ;
        RECT 24.865 113.455 26.535 114.225 ;
        RECT 26.710 114.165 26.920 114.815 ;
        RECT 27.660 114.695 27.830 115.285 ;
        RECT 29.050 115.115 29.220 115.495 ;
        RECT 30.155 115.375 30.325 115.835 ;
        RECT 30.495 115.545 30.865 116.005 ;
        RECT 31.160 115.405 31.330 115.745 ;
        RECT 31.500 115.575 31.830 116.005 ;
        RECT 32.065 115.405 32.235 115.745 ;
        RECT 28.000 114.945 29.220 115.115 ;
        RECT 29.390 115.035 29.850 115.325 ;
        RECT 30.155 115.205 30.715 115.375 ;
        RECT 31.160 115.235 32.235 115.405 ;
        RECT 32.405 115.505 33.085 115.835 ;
        RECT 33.300 115.505 33.550 115.835 ;
        RECT 33.720 115.545 33.970 116.005 ;
        RECT 30.545 115.065 30.715 115.205 ;
        RECT 29.390 115.025 30.355 115.035 ;
        RECT 29.050 114.855 29.220 114.945 ;
        RECT 29.680 114.865 30.355 115.025 ;
        RECT 27.090 114.665 27.830 114.695 ;
        RECT 27.090 114.365 28.005 114.665 ;
        RECT 27.680 114.190 28.005 114.365 ;
        RECT 26.710 113.635 26.965 114.165 ;
        RECT 27.135 113.455 27.440 113.915 ;
        RECT 27.685 113.835 28.005 114.190 ;
        RECT 28.175 114.405 28.715 114.775 ;
        RECT 29.050 114.685 29.455 114.855 ;
        RECT 28.175 114.005 28.415 114.405 ;
        RECT 28.895 114.235 29.115 114.515 ;
        RECT 28.585 114.065 29.115 114.235 ;
        RECT 28.585 113.835 28.755 114.065 ;
        RECT 29.285 113.905 29.455 114.685 ;
        RECT 29.625 114.075 29.975 114.695 ;
        RECT 30.145 114.075 30.355 114.865 ;
        RECT 30.545 114.895 32.045 115.065 ;
        RECT 30.545 114.205 30.715 114.895 ;
        RECT 32.405 114.725 32.575 115.505 ;
        RECT 33.380 115.375 33.550 115.505 ;
        RECT 30.885 114.555 32.575 114.725 ;
        RECT 32.745 114.945 33.210 115.335 ;
        RECT 33.380 115.205 33.775 115.375 ;
        RECT 30.885 114.375 31.055 114.555 ;
        RECT 27.685 113.665 28.755 113.835 ;
        RECT 28.925 113.455 29.115 113.895 ;
        RECT 29.285 113.625 30.235 113.905 ;
        RECT 30.545 113.815 30.805 114.205 ;
        RECT 31.225 114.135 32.015 114.385 ;
        RECT 30.455 113.645 30.805 113.815 ;
        RECT 31.015 113.455 31.345 113.915 ;
        RECT 32.220 113.845 32.390 114.555 ;
        RECT 32.745 114.355 32.915 114.945 ;
        RECT 32.560 114.135 32.915 114.355 ;
        RECT 33.085 114.135 33.435 114.755 ;
        RECT 33.605 113.845 33.775 115.205 ;
        RECT 34.140 115.035 34.465 115.820 ;
        RECT 33.945 113.985 34.405 115.035 ;
        RECT 32.220 113.675 33.075 113.845 ;
        RECT 33.280 113.675 33.775 113.845 ;
        RECT 33.945 113.455 34.275 113.815 ;
        RECT 34.635 113.715 34.805 115.835 ;
        RECT 34.975 115.505 35.305 116.005 ;
        RECT 35.475 115.335 35.730 115.835 ;
        RECT 34.980 115.165 35.730 115.335 ;
        RECT 34.980 114.175 35.210 115.165 ;
        RECT 35.380 114.345 35.730 114.995 ;
        RECT 35.905 114.930 36.175 115.835 ;
        RECT 36.345 115.245 36.675 116.005 ;
        RECT 36.855 115.075 37.025 115.835 ;
        RECT 34.980 114.005 35.730 114.175 ;
        RECT 34.975 113.455 35.305 113.835 ;
        RECT 35.475 113.715 35.730 114.005 ;
        RECT 35.905 114.130 36.075 114.930 ;
        RECT 36.360 114.905 37.025 115.075 ;
        RECT 37.285 114.930 37.555 115.835 ;
        RECT 37.725 115.245 38.055 116.005 ;
        RECT 38.235 115.075 38.405 115.835 ;
        RECT 36.360 114.760 36.530 114.905 ;
        RECT 36.245 114.430 36.530 114.760 ;
        RECT 36.360 114.175 36.530 114.430 ;
        RECT 36.765 114.355 37.095 114.725 ;
        RECT 35.905 113.625 36.165 114.130 ;
        RECT 36.360 114.005 37.025 114.175 ;
        RECT 36.345 113.455 36.675 113.835 ;
        RECT 36.855 113.625 37.025 114.005 ;
        RECT 37.285 114.130 37.455 114.930 ;
        RECT 37.740 114.905 38.405 115.075 ;
        RECT 37.740 114.760 37.910 114.905 ;
        RECT 38.725 114.865 38.935 116.005 ;
        RECT 37.625 114.430 37.910 114.760 ;
        RECT 39.105 114.855 39.435 115.835 ;
        RECT 39.605 114.865 39.835 116.005 ;
        RECT 40.050 115.570 45.395 116.005 ;
        RECT 37.740 114.175 37.910 114.430 ;
        RECT 38.145 114.355 38.475 114.725 ;
        RECT 37.285 113.625 37.545 114.130 ;
        RECT 37.740 114.005 38.405 114.175 ;
        RECT 37.725 113.455 38.055 113.835 ;
        RECT 38.235 113.625 38.405 114.005 ;
        RECT 38.725 113.455 38.935 114.275 ;
        RECT 39.105 114.255 39.355 114.855 ;
        RECT 39.525 114.445 39.855 114.695 ;
        RECT 41.640 114.320 41.990 115.570 ;
        RECT 45.655 115.075 45.825 115.835 ;
        RECT 46.005 115.245 46.335 116.005 ;
        RECT 45.655 114.905 46.320 115.075 ;
        RECT 46.505 114.930 46.775 115.835 ;
        RECT 39.105 113.625 39.435 114.255 ;
        RECT 39.605 113.455 39.835 114.275 ;
        RECT 43.470 114.000 43.810 114.830 ;
        RECT 46.150 114.760 46.320 114.905 ;
        RECT 45.585 114.355 45.915 114.725 ;
        RECT 46.150 114.430 46.435 114.760 ;
        RECT 46.150 114.175 46.320 114.430 ;
        RECT 45.655 114.005 46.320 114.175 ;
        RECT 46.605 114.130 46.775 114.930 ;
        RECT 46.945 114.915 48.155 116.005 ;
        RECT 46.945 114.375 47.465 114.915 ;
        RECT 48.385 114.865 48.595 116.005 ;
        RECT 48.765 114.855 49.095 115.835 ;
        RECT 49.265 114.865 49.495 116.005 ;
        RECT 47.635 114.205 48.155 114.745 ;
        RECT 40.050 113.455 45.395 114.000 ;
        RECT 45.655 113.625 45.825 114.005 ;
        RECT 46.005 113.455 46.335 113.835 ;
        RECT 46.515 113.625 46.775 114.130 ;
        RECT 46.945 113.455 48.155 114.205 ;
        RECT 48.385 113.455 48.595 114.275 ;
        RECT 48.765 114.255 49.015 114.855 ;
        RECT 50.165 114.840 50.455 116.005 ;
        RECT 51.085 114.915 53.675 116.005 ;
        RECT 53.935 115.075 54.105 115.835 ;
        RECT 54.285 115.245 54.615 116.005 ;
        RECT 49.185 114.445 49.515 114.695 ;
        RECT 51.085 114.395 52.295 114.915 ;
        RECT 53.935 114.905 54.600 115.075 ;
        RECT 54.785 114.930 55.055 115.835 ;
        RECT 54.430 114.760 54.600 114.905 ;
        RECT 48.765 113.625 49.095 114.255 ;
        RECT 49.265 113.455 49.495 114.275 ;
        RECT 52.465 114.225 53.675 114.745 ;
        RECT 53.865 114.355 54.195 114.725 ;
        RECT 54.430 114.430 54.715 114.760 ;
        RECT 50.165 113.455 50.455 114.180 ;
        RECT 51.085 113.455 53.675 114.225 ;
        RECT 54.430 114.175 54.600 114.430 ;
        RECT 53.935 114.005 54.600 114.175 ;
        RECT 54.885 114.130 55.055 114.930 ;
        RECT 55.225 114.915 56.895 116.005 ;
        RECT 57.070 115.570 62.415 116.005 ;
        RECT 55.225 114.395 55.975 114.915 ;
        RECT 56.145 114.225 56.895 114.745 ;
        RECT 58.660 114.320 59.010 115.570 ;
        RECT 62.595 115.025 62.925 115.835 ;
        RECT 63.095 115.205 63.335 116.005 ;
        RECT 62.595 114.855 63.310 115.025 ;
        RECT 53.935 113.625 54.105 114.005 ;
        RECT 54.285 113.455 54.615 113.835 ;
        RECT 54.795 113.625 55.055 114.130 ;
        RECT 55.225 113.455 56.895 114.225 ;
        RECT 60.490 114.000 60.830 114.830 ;
        RECT 62.590 114.445 62.970 114.685 ;
        RECT 63.140 114.615 63.310 114.855 ;
        RECT 63.515 114.985 63.685 115.835 ;
        RECT 63.855 115.205 64.185 116.005 ;
        RECT 64.355 114.985 64.525 115.835 ;
        RECT 63.515 114.815 64.525 114.985 ;
        RECT 64.695 114.855 65.025 116.005 ;
        RECT 65.350 115.570 70.695 116.005 ;
        RECT 63.140 114.445 63.640 114.615 ;
        RECT 63.140 114.275 63.310 114.445 ;
        RECT 64.030 114.305 64.525 114.815 ;
        RECT 66.940 114.320 67.290 115.570 ;
        RECT 70.955 115.075 71.125 115.835 ;
        RECT 71.305 115.245 71.635 116.005 ;
        RECT 70.955 114.905 71.620 115.075 ;
        RECT 71.805 114.930 72.075 115.835 ;
        RECT 64.025 114.275 64.525 114.305 ;
        RECT 62.675 114.105 63.310 114.275 ;
        RECT 63.515 114.105 64.525 114.275 ;
        RECT 57.070 113.455 62.415 114.000 ;
        RECT 62.675 113.625 62.845 114.105 ;
        RECT 63.025 113.455 63.265 113.935 ;
        RECT 63.515 113.625 63.685 114.105 ;
        RECT 63.855 113.455 64.185 113.935 ;
        RECT 64.355 113.625 64.525 114.105 ;
        RECT 64.695 113.455 65.025 114.255 ;
        RECT 68.770 114.000 69.110 114.830 ;
        RECT 71.450 114.760 71.620 114.905 ;
        RECT 70.885 114.355 71.215 114.725 ;
        RECT 71.450 114.430 71.735 114.760 ;
        RECT 71.450 114.175 71.620 114.430 ;
        RECT 70.955 114.005 71.620 114.175 ;
        RECT 71.905 114.130 72.075 114.930 ;
        RECT 72.245 114.915 75.755 116.005 ;
        RECT 72.245 114.395 73.935 114.915 ;
        RECT 75.925 114.840 76.215 116.005 ;
        RECT 76.845 114.915 78.515 116.005 ;
        RECT 74.105 114.225 75.755 114.745 ;
        RECT 76.845 114.395 77.595 114.915 ;
        RECT 78.745 114.865 78.955 116.005 ;
        RECT 79.125 114.855 79.455 115.835 ;
        RECT 79.625 114.865 79.855 116.005 ;
        RECT 80.105 114.865 80.335 116.005 ;
        RECT 80.505 114.855 80.835 115.835 ;
        RECT 81.005 114.865 81.215 116.005 ;
        RECT 81.535 115.075 81.705 115.835 ;
        RECT 81.885 115.245 82.215 116.005 ;
        RECT 81.535 114.905 82.200 115.075 ;
        RECT 82.385 114.930 82.655 115.835 ;
        RECT 77.765 114.225 78.515 114.745 ;
        RECT 65.350 113.455 70.695 114.000 ;
        RECT 70.955 113.625 71.125 114.005 ;
        RECT 71.305 113.455 71.635 113.835 ;
        RECT 71.815 113.625 72.075 114.130 ;
        RECT 72.245 113.455 75.755 114.225 ;
        RECT 75.925 113.455 76.215 114.180 ;
        RECT 76.845 113.455 78.515 114.225 ;
        RECT 78.745 113.455 78.955 114.275 ;
        RECT 79.125 114.255 79.375 114.855 ;
        RECT 79.545 114.445 79.875 114.695 ;
        RECT 80.085 114.445 80.415 114.695 ;
        RECT 79.125 113.625 79.455 114.255 ;
        RECT 79.625 113.455 79.855 114.275 ;
        RECT 80.105 113.455 80.335 114.275 ;
        RECT 80.585 114.255 80.835 114.855 ;
        RECT 82.030 114.760 82.200 114.905 ;
        RECT 81.465 114.355 81.795 114.725 ;
        RECT 82.030 114.430 82.315 114.760 ;
        RECT 80.505 113.625 80.835 114.255 ;
        RECT 81.005 113.455 81.215 114.275 ;
        RECT 82.030 114.175 82.200 114.430 ;
        RECT 81.535 114.005 82.200 114.175 ;
        RECT 82.485 114.130 82.655 114.930 ;
        RECT 83.295 115.025 83.625 115.835 ;
        RECT 83.795 115.205 84.035 116.005 ;
        RECT 83.295 114.855 84.010 115.025 ;
        RECT 83.290 114.445 83.670 114.685 ;
        RECT 83.840 114.615 84.010 114.855 ;
        RECT 84.215 114.985 84.385 115.835 ;
        RECT 84.555 115.205 84.885 116.005 ;
        RECT 85.055 114.985 85.225 115.835 ;
        RECT 84.215 114.815 85.225 114.985 ;
        RECT 85.395 114.855 85.725 116.005 ;
        RECT 86.135 115.075 86.305 115.835 ;
        RECT 86.485 115.245 86.815 116.005 ;
        RECT 86.135 114.905 86.800 115.075 ;
        RECT 86.985 114.930 87.255 115.835 ;
        RECT 87.890 115.570 93.235 116.005 ;
        RECT 83.840 114.445 84.340 114.615 ;
        RECT 83.840 114.275 84.010 114.445 ;
        RECT 84.730 114.305 85.225 114.815 ;
        RECT 86.630 114.760 86.800 114.905 ;
        RECT 86.065 114.355 86.395 114.725 ;
        RECT 86.630 114.430 86.915 114.760 ;
        RECT 84.725 114.275 85.225 114.305 ;
        RECT 81.535 113.625 81.705 114.005 ;
        RECT 81.885 113.455 82.215 113.835 ;
        RECT 82.395 113.625 82.655 114.130 ;
        RECT 83.375 114.105 84.010 114.275 ;
        RECT 84.215 114.105 85.225 114.275 ;
        RECT 83.375 113.625 83.545 114.105 ;
        RECT 83.725 113.455 83.965 113.935 ;
        RECT 84.215 113.625 84.385 114.105 ;
        RECT 84.555 113.455 84.885 113.935 ;
        RECT 85.055 113.625 85.225 114.105 ;
        RECT 85.395 113.455 85.725 114.255 ;
        RECT 86.630 114.175 86.800 114.430 ;
        RECT 86.135 114.005 86.800 114.175 ;
        RECT 87.085 114.130 87.255 114.930 ;
        RECT 89.480 114.320 89.830 115.570 ;
        RECT 93.465 114.865 93.675 116.005 ;
        RECT 93.845 114.855 94.175 115.835 ;
        RECT 94.345 114.865 94.575 116.005 ;
        RECT 94.875 115.075 95.045 115.835 ;
        RECT 95.225 115.245 95.555 116.005 ;
        RECT 94.875 114.905 95.540 115.075 ;
        RECT 95.725 114.930 95.995 115.835 ;
        RECT 86.135 113.625 86.305 114.005 ;
        RECT 86.485 113.455 86.815 113.835 ;
        RECT 86.995 113.625 87.255 114.130 ;
        RECT 91.310 114.000 91.650 114.830 ;
        RECT 87.890 113.455 93.235 114.000 ;
        RECT 93.465 113.455 93.675 114.275 ;
        RECT 93.845 114.255 94.095 114.855 ;
        RECT 95.370 114.760 95.540 114.905 ;
        RECT 94.265 114.445 94.595 114.695 ;
        RECT 94.805 114.355 95.135 114.725 ;
        RECT 95.370 114.430 95.655 114.760 ;
        RECT 93.845 113.625 94.175 114.255 ;
        RECT 94.345 113.455 94.575 114.275 ;
        RECT 95.370 114.175 95.540 114.430 ;
        RECT 94.875 114.005 95.540 114.175 ;
        RECT 95.825 114.130 95.995 114.930 ;
        RECT 96.165 114.915 97.375 116.005 ;
        RECT 96.165 114.375 96.685 114.915 ;
        RECT 97.585 114.865 97.815 116.005 ;
        RECT 97.985 114.855 98.315 115.835 ;
        RECT 98.485 114.865 98.695 116.005 ;
        RECT 98.925 114.915 101.515 116.005 ;
        RECT 96.855 114.205 97.375 114.745 ;
        RECT 97.565 114.445 97.895 114.695 ;
        RECT 94.875 113.625 95.045 114.005 ;
        RECT 95.225 113.455 95.555 113.835 ;
        RECT 95.735 113.625 95.995 114.130 ;
        RECT 96.165 113.455 97.375 114.205 ;
        RECT 97.585 113.455 97.815 114.275 ;
        RECT 98.065 114.255 98.315 114.855 ;
        RECT 98.925 114.395 100.135 114.915 ;
        RECT 101.685 114.840 101.975 116.005 ;
        RECT 102.605 114.915 104.275 116.005 ;
        RECT 97.985 113.625 98.315 114.255 ;
        RECT 98.485 113.455 98.695 114.275 ;
        RECT 100.305 114.225 101.515 114.745 ;
        RECT 102.605 114.395 103.355 114.915 ;
        RECT 104.505 114.865 104.715 116.005 ;
        RECT 104.885 114.855 105.215 115.835 ;
        RECT 105.385 114.865 105.615 116.005 ;
        RECT 106.835 115.075 107.005 115.835 ;
        RECT 107.185 115.245 107.515 116.005 ;
        RECT 106.835 114.905 107.500 115.075 ;
        RECT 107.685 114.930 107.955 115.835 ;
        RECT 103.525 114.225 104.275 114.745 ;
        RECT 98.925 113.455 101.515 114.225 ;
        RECT 101.685 113.455 101.975 114.180 ;
        RECT 102.605 113.455 104.275 114.225 ;
        RECT 104.505 113.455 104.715 114.275 ;
        RECT 104.885 114.255 105.135 114.855 ;
        RECT 107.330 114.760 107.500 114.905 ;
        RECT 105.305 114.445 105.635 114.695 ;
        RECT 106.765 114.355 107.095 114.725 ;
        RECT 107.330 114.430 107.615 114.760 ;
        RECT 104.885 113.625 105.215 114.255 ;
        RECT 105.385 113.455 105.615 114.275 ;
        RECT 107.330 114.175 107.500 114.430 ;
        RECT 106.835 114.005 107.500 114.175 ;
        RECT 107.785 114.130 107.955 114.930 ;
        RECT 108.185 114.865 108.395 116.005 ;
        RECT 108.565 114.855 108.895 115.835 ;
        RECT 109.065 114.865 109.295 116.005 ;
        RECT 110.430 115.570 115.775 116.005 ;
        RECT 106.835 113.625 107.005 114.005 ;
        RECT 107.185 113.455 107.515 113.835 ;
        RECT 107.695 113.625 107.955 114.130 ;
        RECT 108.185 113.455 108.395 114.275 ;
        RECT 108.565 114.255 108.815 114.855 ;
        RECT 108.985 114.445 109.315 114.695 ;
        RECT 112.020 114.320 112.370 115.570 ;
        RECT 115.985 114.865 116.215 116.005 ;
        RECT 116.385 114.855 116.715 115.835 ;
        RECT 116.885 114.865 117.095 116.005 ;
        RECT 117.330 115.335 117.585 115.835 ;
        RECT 117.755 115.505 118.085 116.005 ;
        RECT 117.330 115.165 118.080 115.335 ;
        RECT 108.565 113.625 108.895 114.255 ;
        RECT 109.065 113.455 109.295 114.275 ;
        RECT 113.850 114.000 114.190 114.830 ;
        RECT 115.965 114.445 116.295 114.695 ;
        RECT 110.430 113.455 115.775 114.000 ;
        RECT 115.985 113.455 116.215 114.275 ;
        RECT 116.465 114.255 116.715 114.855 ;
        RECT 117.330 114.345 117.680 114.995 ;
        RECT 116.385 113.625 116.715 114.255 ;
        RECT 116.885 113.455 117.095 114.275 ;
        RECT 117.850 114.175 118.080 115.165 ;
        RECT 117.330 114.005 118.080 114.175 ;
        RECT 117.330 113.715 117.585 114.005 ;
        RECT 117.755 113.455 118.085 113.835 ;
        RECT 118.255 113.715 118.425 115.835 ;
        RECT 118.595 115.035 118.920 115.820 ;
        RECT 119.090 115.545 119.340 116.005 ;
        RECT 119.510 115.505 119.760 115.835 ;
        RECT 119.975 115.505 120.655 115.835 ;
        RECT 119.510 115.375 119.680 115.505 ;
        RECT 119.285 115.205 119.680 115.375 ;
        RECT 118.655 113.985 119.115 115.035 ;
        RECT 119.285 113.845 119.455 115.205 ;
        RECT 119.850 114.945 120.315 115.335 ;
        RECT 119.625 114.135 119.975 114.755 ;
        RECT 120.145 114.355 120.315 114.945 ;
        RECT 120.485 114.725 120.655 115.505 ;
        RECT 120.825 115.405 120.995 115.745 ;
        RECT 121.230 115.575 121.560 116.005 ;
        RECT 121.730 115.405 121.900 115.745 ;
        RECT 122.195 115.545 122.565 116.005 ;
        RECT 120.825 115.235 121.900 115.405 ;
        RECT 122.735 115.375 122.905 115.835 ;
        RECT 123.140 115.495 124.010 115.835 ;
        RECT 124.180 115.545 124.430 116.005 ;
        RECT 122.345 115.205 122.905 115.375 ;
        RECT 122.345 115.065 122.515 115.205 ;
        RECT 121.015 114.895 122.515 115.065 ;
        RECT 123.210 115.035 123.670 115.325 ;
        RECT 120.485 114.555 122.175 114.725 ;
        RECT 120.145 114.135 120.500 114.355 ;
        RECT 120.670 113.845 120.840 114.555 ;
        RECT 121.045 114.135 121.835 114.385 ;
        RECT 122.005 114.375 122.175 114.555 ;
        RECT 122.345 114.205 122.515 114.895 ;
        RECT 118.785 113.455 119.115 113.815 ;
        RECT 119.285 113.675 119.780 113.845 ;
        RECT 119.985 113.675 120.840 113.845 ;
        RECT 121.715 113.455 122.045 113.915 ;
        RECT 122.255 113.815 122.515 114.205 ;
        RECT 122.705 115.025 123.670 115.035 ;
        RECT 123.840 115.115 124.010 115.495 ;
        RECT 124.600 115.455 124.770 115.745 ;
        RECT 124.950 115.625 125.280 116.005 ;
        RECT 124.600 115.285 125.400 115.455 ;
        RECT 122.705 114.865 123.380 115.025 ;
        RECT 123.840 114.945 125.060 115.115 ;
        RECT 122.705 114.075 122.915 114.865 ;
        RECT 123.840 114.855 124.010 114.945 ;
        RECT 123.085 114.075 123.435 114.695 ;
        RECT 123.605 114.685 124.010 114.855 ;
        RECT 123.605 113.905 123.775 114.685 ;
        RECT 123.945 114.235 124.165 114.515 ;
        RECT 124.345 114.405 124.885 114.775 ;
        RECT 125.230 114.695 125.400 115.285 ;
        RECT 125.620 114.865 125.925 116.005 ;
        RECT 126.095 114.815 126.350 115.695 ;
        RECT 125.230 114.665 125.970 114.695 ;
        RECT 123.945 114.065 124.475 114.235 ;
        RECT 122.255 113.645 122.605 113.815 ;
        RECT 122.825 113.625 123.775 113.905 ;
        RECT 123.945 113.455 124.135 113.895 ;
        RECT 124.305 113.835 124.475 114.065 ;
        RECT 124.645 114.005 124.885 114.405 ;
        RECT 125.055 114.365 125.970 114.665 ;
        RECT 125.055 114.190 125.380 114.365 ;
        RECT 125.055 113.835 125.375 114.190 ;
        RECT 126.140 114.165 126.350 114.815 ;
        RECT 126.525 114.915 127.735 116.005 ;
        RECT 126.525 114.375 127.045 114.915 ;
        RECT 127.215 114.205 127.735 114.745 ;
        RECT 124.305 113.665 125.375 113.835 ;
        RECT 125.620 113.455 125.925 113.915 ;
        RECT 126.095 113.635 126.350 114.165 ;
        RECT 126.525 113.455 127.735 114.205 ;
        RECT 20.640 113.285 127.820 113.455 ;
        RECT 20.725 112.535 21.935 113.285 ;
        RECT 20.725 111.995 21.245 112.535 ;
        RECT 22.105 112.515 23.775 113.285 ;
        RECT 21.415 111.825 21.935 112.365 ;
        RECT 20.725 110.735 21.935 111.825 ;
        RECT 22.105 111.825 22.855 112.345 ;
        RECT 23.025 111.995 23.775 112.515 ;
        RECT 24.005 112.465 24.215 113.285 ;
        RECT 24.385 112.485 24.715 113.115 ;
        RECT 24.385 111.885 24.635 112.485 ;
        RECT 24.885 112.465 25.115 113.285 ;
        RECT 25.365 112.465 25.595 113.285 ;
        RECT 25.765 112.485 26.095 113.115 ;
        RECT 24.805 112.045 25.135 112.295 ;
        RECT 25.345 112.045 25.675 112.295 ;
        RECT 25.845 111.885 26.095 112.485 ;
        RECT 26.265 112.465 26.475 113.285 ;
        RECT 26.745 112.465 26.975 113.285 ;
        RECT 27.145 112.485 27.475 113.115 ;
        RECT 26.725 112.045 27.055 112.295 ;
        RECT 27.225 111.885 27.475 112.485 ;
        RECT 27.645 112.465 27.855 113.285 ;
        RECT 28.090 112.575 28.345 113.105 ;
        RECT 28.515 112.825 28.820 113.285 ;
        RECT 29.065 112.905 30.135 113.075 ;
        RECT 22.105 110.735 23.775 111.825 ;
        RECT 24.005 110.735 24.215 111.875 ;
        RECT 24.385 110.905 24.715 111.885 ;
        RECT 24.885 110.735 25.115 111.875 ;
        RECT 25.365 110.735 25.595 111.875 ;
        RECT 25.765 110.905 26.095 111.885 ;
        RECT 26.265 110.735 26.475 111.875 ;
        RECT 26.745 110.735 26.975 111.875 ;
        RECT 27.145 110.905 27.475 111.885 ;
        RECT 28.090 111.925 28.300 112.575 ;
        RECT 29.065 112.550 29.385 112.905 ;
        RECT 29.060 112.375 29.385 112.550 ;
        RECT 28.470 112.075 29.385 112.375 ;
        RECT 29.555 112.335 29.795 112.735 ;
        RECT 29.965 112.675 30.135 112.905 ;
        RECT 30.305 112.845 30.495 113.285 ;
        RECT 30.665 112.835 31.615 113.115 ;
        RECT 31.835 112.925 32.185 113.095 ;
        RECT 29.965 112.505 30.495 112.675 ;
        RECT 28.470 112.045 29.210 112.075 ;
        RECT 27.645 110.735 27.855 111.875 ;
        RECT 28.090 111.045 28.345 111.925 ;
        RECT 28.515 110.735 28.820 111.875 ;
        RECT 29.040 111.455 29.210 112.045 ;
        RECT 29.555 111.965 30.095 112.335 ;
        RECT 30.275 112.225 30.495 112.505 ;
        RECT 30.665 112.055 30.835 112.835 ;
        RECT 30.430 111.885 30.835 112.055 ;
        RECT 31.005 112.045 31.355 112.665 ;
        RECT 30.430 111.795 30.600 111.885 ;
        RECT 31.525 111.875 31.735 112.665 ;
        RECT 29.380 111.625 30.600 111.795 ;
        RECT 31.060 111.715 31.735 111.875 ;
        RECT 29.040 111.285 29.840 111.455 ;
        RECT 29.160 110.735 29.490 111.115 ;
        RECT 29.670 110.995 29.840 111.285 ;
        RECT 30.430 111.245 30.600 111.625 ;
        RECT 30.770 111.705 31.735 111.715 ;
        RECT 31.925 112.535 32.185 112.925 ;
        RECT 32.395 112.825 32.725 113.285 ;
        RECT 33.600 112.895 34.455 113.065 ;
        RECT 34.660 112.895 35.155 113.065 ;
        RECT 35.325 112.925 35.655 113.285 ;
        RECT 31.925 111.845 32.095 112.535 ;
        RECT 32.265 112.185 32.435 112.365 ;
        RECT 32.605 112.355 33.395 112.605 ;
        RECT 33.600 112.185 33.770 112.895 ;
        RECT 33.940 112.385 34.295 112.605 ;
        RECT 32.265 112.015 33.955 112.185 ;
        RECT 30.770 111.415 31.230 111.705 ;
        RECT 31.925 111.675 33.425 111.845 ;
        RECT 31.925 111.535 32.095 111.675 ;
        RECT 31.535 111.365 32.095 111.535 ;
        RECT 30.010 110.735 30.260 111.195 ;
        RECT 30.430 110.905 31.300 111.245 ;
        RECT 31.535 110.905 31.705 111.365 ;
        RECT 32.540 111.335 33.615 111.505 ;
        RECT 31.875 110.735 32.245 111.195 ;
        RECT 32.540 110.995 32.710 111.335 ;
        RECT 32.880 110.735 33.210 111.165 ;
        RECT 33.445 110.995 33.615 111.335 ;
        RECT 33.785 111.235 33.955 112.015 ;
        RECT 34.125 111.795 34.295 112.385 ;
        RECT 34.465 111.985 34.815 112.605 ;
        RECT 34.125 111.405 34.590 111.795 ;
        RECT 34.985 111.535 35.155 112.895 ;
        RECT 35.325 111.705 35.785 112.755 ;
        RECT 34.760 111.365 35.155 111.535 ;
        RECT 34.760 111.235 34.930 111.365 ;
        RECT 33.785 110.905 34.465 111.235 ;
        RECT 34.680 110.905 34.930 111.235 ;
        RECT 35.100 110.735 35.350 111.195 ;
        RECT 35.520 110.920 35.845 111.705 ;
        RECT 36.015 110.905 36.185 113.025 ;
        RECT 36.355 112.905 36.685 113.285 ;
        RECT 36.855 112.735 37.110 113.025 ;
        RECT 36.360 112.565 37.110 112.735 ;
        RECT 36.360 111.575 36.590 112.565 ;
        RECT 37.285 112.560 37.575 113.285 ;
        RECT 37.835 112.735 38.005 113.115 ;
        RECT 38.185 112.905 38.515 113.285 ;
        RECT 37.835 112.565 38.500 112.735 ;
        RECT 38.695 112.610 38.955 113.115 ;
        RECT 36.760 111.745 37.110 112.395 ;
        RECT 37.765 112.015 38.095 112.385 ;
        RECT 38.330 112.310 38.500 112.565 ;
        RECT 38.330 111.980 38.615 112.310 ;
        RECT 36.360 111.405 37.110 111.575 ;
        RECT 36.355 110.735 36.685 111.235 ;
        RECT 36.855 110.905 37.110 111.405 ;
        RECT 37.285 110.735 37.575 111.900 ;
        RECT 38.330 111.835 38.500 111.980 ;
        RECT 37.835 111.665 38.500 111.835 ;
        RECT 38.785 111.810 38.955 112.610 ;
        RECT 39.165 112.465 39.395 113.285 ;
        RECT 39.565 112.485 39.895 113.115 ;
        RECT 39.145 112.045 39.475 112.295 ;
        RECT 39.645 111.885 39.895 112.485 ;
        RECT 40.065 112.465 40.275 113.285 ;
        RECT 40.510 112.575 40.765 113.105 ;
        RECT 40.935 112.825 41.240 113.285 ;
        RECT 41.485 112.905 42.555 113.075 ;
        RECT 37.835 110.905 38.005 111.665 ;
        RECT 38.185 110.735 38.515 111.495 ;
        RECT 38.685 110.905 38.955 111.810 ;
        RECT 39.165 110.735 39.395 111.875 ;
        RECT 39.565 110.905 39.895 111.885 ;
        RECT 40.510 111.925 40.720 112.575 ;
        RECT 41.485 112.550 41.805 112.905 ;
        RECT 41.480 112.375 41.805 112.550 ;
        RECT 40.890 112.075 41.805 112.375 ;
        RECT 41.975 112.335 42.215 112.735 ;
        RECT 42.385 112.675 42.555 112.905 ;
        RECT 42.725 112.845 42.915 113.285 ;
        RECT 43.085 112.835 44.035 113.115 ;
        RECT 44.255 112.925 44.605 113.095 ;
        RECT 42.385 112.505 42.915 112.675 ;
        RECT 40.890 112.045 41.630 112.075 ;
        RECT 40.065 110.735 40.275 111.875 ;
        RECT 40.510 111.045 40.765 111.925 ;
        RECT 40.935 110.735 41.240 111.875 ;
        RECT 41.460 111.455 41.630 112.045 ;
        RECT 41.975 111.965 42.515 112.335 ;
        RECT 42.695 112.225 42.915 112.505 ;
        RECT 43.085 112.055 43.255 112.835 ;
        RECT 42.850 111.885 43.255 112.055 ;
        RECT 43.425 112.045 43.775 112.665 ;
        RECT 42.850 111.795 43.020 111.885 ;
        RECT 43.945 111.875 44.155 112.665 ;
        RECT 41.800 111.625 43.020 111.795 ;
        RECT 43.480 111.715 44.155 111.875 ;
        RECT 41.460 111.285 42.260 111.455 ;
        RECT 41.580 110.735 41.910 111.115 ;
        RECT 42.090 110.995 42.260 111.285 ;
        RECT 42.850 111.245 43.020 111.625 ;
        RECT 43.190 111.705 44.155 111.715 ;
        RECT 44.345 112.535 44.605 112.925 ;
        RECT 44.815 112.825 45.145 113.285 ;
        RECT 46.020 112.895 46.875 113.065 ;
        RECT 47.080 112.895 47.575 113.065 ;
        RECT 47.745 112.925 48.075 113.285 ;
        RECT 44.345 111.845 44.515 112.535 ;
        RECT 44.685 112.185 44.855 112.365 ;
        RECT 45.025 112.355 45.815 112.605 ;
        RECT 46.020 112.185 46.190 112.895 ;
        RECT 46.360 112.385 46.715 112.605 ;
        RECT 44.685 112.015 46.375 112.185 ;
        RECT 43.190 111.415 43.650 111.705 ;
        RECT 44.345 111.675 45.845 111.845 ;
        RECT 44.345 111.535 44.515 111.675 ;
        RECT 43.955 111.365 44.515 111.535 ;
        RECT 42.430 110.735 42.680 111.195 ;
        RECT 42.850 110.905 43.720 111.245 ;
        RECT 43.955 110.905 44.125 111.365 ;
        RECT 44.960 111.335 46.035 111.505 ;
        RECT 44.295 110.735 44.665 111.195 ;
        RECT 44.960 110.995 45.130 111.335 ;
        RECT 45.300 110.735 45.630 111.165 ;
        RECT 45.865 110.995 46.035 111.335 ;
        RECT 46.205 111.235 46.375 112.015 ;
        RECT 46.545 111.795 46.715 112.385 ;
        RECT 46.885 111.985 47.235 112.605 ;
        RECT 46.545 111.405 47.010 111.795 ;
        RECT 47.405 111.535 47.575 112.895 ;
        RECT 47.745 111.705 48.205 112.755 ;
        RECT 47.180 111.365 47.575 111.535 ;
        RECT 47.180 111.235 47.350 111.365 ;
        RECT 46.205 110.905 46.885 111.235 ;
        RECT 47.100 110.905 47.350 111.235 ;
        RECT 47.520 110.735 47.770 111.195 ;
        RECT 47.940 110.920 48.265 111.705 ;
        RECT 48.435 110.905 48.605 113.025 ;
        RECT 48.775 112.905 49.105 113.285 ;
        RECT 49.275 112.735 49.530 113.025 ;
        RECT 48.780 112.565 49.530 112.735 ;
        RECT 49.705 112.610 49.965 113.115 ;
        RECT 50.145 112.905 50.475 113.285 ;
        RECT 50.655 112.735 50.825 113.115 ;
        RECT 48.780 111.575 49.010 112.565 ;
        RECT 49.180 111.745 49.530 112.395 ;
        RECT 49.705 111.810 49.875 112.610 ;
        RECT 50.160 112.565 50.825 112.735 ;
        RECT 51.550 112.575 51.805 113.105 ;
        RECT 51.975 112.825 52.280 113.285 ;
        RECT 52.525 112.905 53.595 113.075 ;
        RECT 50.160 112.310 50.330 112.565 ;
        RECT 50.045 111.980 50.330 112.310 ;
        RECT 50.565 112.015 50.895 112.385 ;
        RECT 50.160 111.835 50.330 111.980 ;
        RECT 51.550 111.925 51.760 112.575 ;
        RECT 52.525 112.550 52.845 112.905 ;
        RECT 52.520 112.375 52.845 112.550 ;
        RECT 51.930 112.075 52.845 112.375 ;
        RECT 53.015 112.335 53.255 112.735 ;
        RECT 53.425 112.675 53.595 112.905 ;
        RECT 53.765 112.845 53.955 113.285 ;
        RECT 54.125 112.835 55.075 113.115 ;
        RECT 55.295 112.925 55.645 113.095 ;
        RECT 53.425 112.505 53.955 112.675 ;
        RECT 51.930 112.045 52.670 112.075 ;
        RECT 48.780 111.405 49.530 111.575 ;
        RECT 48.775 110.735 49.105 111.235 ;
        RECT 49.275 110.905 49.530 111.405 ;
        RECT 49.705 110.905 49.975 111.810 ;
        RECT 50.160 111.665 50.825 111.835 ;
        RECT 50.145 110.735 50.475 111.495 ;
        RECT 50.655 110.905 50.825 111.665 ;
        RECT 51.550 111.045 51.805 111.925 ;
        RECT 51.975 110.735 52.280 111.875 ;
        RECT 52.500 111.455 52.670 112.045 ;
        RECT 53.015 111.965 53.555 112.335 ;
        RECT 53.735 112.225 53.955 112.505 ;
        RECT 54.125 112.055 54.295 112.835 ;
        RECT 53.890 111.885 54.295 112.055 ;
        RECT 54.465 112.045 54.815 112.665 ;
        RECT 53.890 111.795 54.060 111.885 ;
        RECT 54.985 111.875 55.195 112.665 ;
        RECT 52.840 111.625 54.060 111.795 ;
        RECT 54.520 111.715 55.195 111.875 ;
        RECT 52.500 111.285 53.300 111.455 ;
        RECT 52.620 110.735 52.950 111.115 ;
        RECT 53.130 110.995 53.300 111.285 ;
        RECT 53.890 111.245 54.060 111.625 ;
        RECT 54.230 111.705 55.195 111.715 ;
        RECT 55.385 112.535 55.645 112.925 ;
        RECT 55.855 112.825 56.185 113.285 ;
        RECT 57.060 112.895 57.915 113.065 ;
        RECT 58.120 112.895 58.615 113.065 ;
        RECT 58.785 112.925 59.115 113.285 ;
        RECT 55.385 111.845 55.555 112.535 ;
        RECT 55.725 112.185 55.895 112.365 ;
        RECT 56.065 112.355 56.855 112.605 ;
        RECT 57.060 112.185 57.230 112.895 ;
        RECT 57.400 112.385 57.755 112.605 ;
        RECT 55.725 112.015 57.415 112.185 ;
        RECT 54.230 111.415 54.690 111.705 ;
        RECT 55.385 111.675 56.885 111.845 ;
        RECT 55.385 111.535 55.555 111.675 ;
        RECT 54.995 111.365 55.555 111.535 ;
        RECT 53.470 110.735 53.720 111.195 ;
        RECT 53.890 110.905 54.760 111.245 ;
        RECT 54.995 110.905 55.165 111.365 ;
        RECT 56.000 111.335 57.075 111.505 ;
        RECT 55.335 110.735 55.705 111.195 ;
        RECT 56.000 110.995 56.170 111.335 ;
        RECT 56.340 110.735 56.670 111.165 ;
        RECT 56.905 110.995 57.075 111.335 ;
        RECT 57.245 111.235 57.415 112.015 ;
        RECT 57.585 111.795 57.755 112.385 ;
        RECT 57.925 111.985 58.275 112.605 ;
        RECT 57.585 111.405 58.050 111.795 ;
        RECT 58.445 111.535 58.615 112.895 ;
        RECT 58.785 111.705 59.245 112.755 ;
        RECT 58.220 111.365 58.615 111.535 ;
        RECT 58.220 111.235 58.390 111.365 ;
        RECT 57.245 110.905 57.925 111.235 ;
        RECT 58.140 110.905 58.390 111.235 ;
        RECT 58.560 110.735 58.810 111.195 ;
        RECT 58.980 110.920 59.305 111.705 ;
        RECT 59.475 110.905 59.645 113.025 ;
        RECT 59.815 112.905 60.145 113.285 ;
        RECT 60.315 112.735 60.570 113.025 ;
        RECT 59.820 112.565 60.570 112.735 ;
        RECT 60.835 112.735 61.005 113.115 ;
        RECT 61.185 112.905 61.515 113.285 ;
        RECT 60.835 112.565 61.500 112.735 ;
        RECT 61.695 112.610 61.955 113.115 ;
        RECT 59.820 111.575 60.050 112.565 ;
        RECT 60.220 111.745 60.570 112.395 ;
        RECT 60.765 112.015 61.095 112.385 ;
        RECT 61.330 112.310 61.500 112.565 ;
        RECT 61.330 111.980 61.615 112.310 ;
        RECT 61.330 111.835 61.500 111.980 ;
        RECT 60.835 111.665 61.500 111.835 ;
        RECT 61.785 111.810 61.955 112.610 ;
        RECT 63.045 112.560 63.335 113.285 ;
        RECT 63.505 112.535 64.715 113.285 ;
        RECT 64.975 112.735 65.145 113.115 ;
        RECT 65.325 112.905 65.655 113.285 ;
        RECT 64.975 112.565 65.640 112.735 ;
        RECT 65.835 112.610 66.095 113.115 ;
        RECT 59.820 111.405 60.570 111.575 ;
        RECT 59.815 110.735 60.145 111.235 ;
        RECT 60.315 110.905 60.570 111.405 ;
        RECT 60.835 110.905 61.005 111.665 ;
        RECT 61.185 110.735 61.515 111.495 ;
        RECT 61.685 110.905 61.955 111.810 ;
        RECT 63.045 110.735 63.335 111.900 ;
        RECT 63.505 111.825 64.025 112.365 ;
        RECT 64.195 111.995 64.715 112.535 ;
        RECT 64.905 112.015 65.235 112.385 ;
        RECT 65.470 112.310 65.640 112.565 ;
        RECT 65.470 111.980 65.755 112.310 ;
        RECT 65.470 111.835 65.640 111.980 ;
        RECT 63.505 110.735 64.715 111.825 ;
        RECT 64.975 111.665 65.640 111.835 ;
        RECT 65.925 111.810 66.095 112.610 ;
        RECT 64.975 110.905 65.145 111.665 ;
        RECT 65.325 110.735 65.655 111.495 ;
        RECT 65.825 110.905 66.095 111.810 ;
        RECT 66.270 112.575 66.525 113.105 ;
        RECT 66.695 112.825 67.000 113.285 ;
        RECT 67.245 112.905 68.315 113.075 ;
        RECT 66.270 111.925 66.480 112.575 ;
        RECT 67.245 112.550 67.565 112.905 ;
        RECT 67.240 112.375 67.565 112.550 ;
        RECT 66.650 112.075 67.565 112.375 ;
        RECT 67.735 112.335 67.975 112.735 ;
        RECT 68.145 112.675 68.315 112.905 ;
        RECT 68.485 112.845 68.675 113.285 ;
        RECT 68.845 112.835 69.795 113.115 ;
        RECT 70.015 112.925 70.365 113.095 ;
        RECT 68.145 112.505 68.675 112.675 ;
        RECT 66.650 112.045 67.390 112.075 ;
        RECT 66.270 111.045 66.525 111.925 ;
        RECT 66.695 110.735 67.000 111.875 ;
        RECT 67.220 111.455 67.390 112.045 ;
        RECT 67.735 111.965 68.275 112.335 ;
        RECT 68.455 112.225 68.675 112.505 ;
        RECT 68.845 112.055 69.015 112.835 ;
        RECT 68.610 111.885 69.015 112.055 ;
        RECT 69.185 112.045 69.535 112.665 ;
        RECT 68.610 111.795 68.780 111.885 ;
        RECT 69.705 111.875 69.915 112.665 ;
        RECT 67.560 111.625 68.780 111.795 ;
        RECT 69.240 111.715 69.915 111.875 ;
        RECT 67.220 111.285 68.020 111.455 ;
        RECT 67.340 110.735 67.670 111.115 ;
        RECT 67.850 110.995 68.020 111.285 ;
        RECT 68.610 111.245 68.780 111.625 ;
        RECT 68.950 111.705 69.915 111.715 ;
        RECT 70.105 112.535 70.365 112.925 ;
        RECT 70.575 112.825 70.905 113.285 ;
        RECT 71.780 112.895 72.635 113.065 ;
        RECT 72.840 112.895 73.335 113.065 ;
        RECT 73.505 112.925 73.835 113.285 ;
        RECT 70.105 111.845 70.275 112.535 ;
        RECT 70.445 112.185 70.615 112.365 ;
        RECT 70.785 112.355 71.575 112.605 ;
        RECT 71.780 112.185 71.950 112.895 ;
        RECT 72.120 112.385 72.475 112.605 ;
        RECT 70.445 112.015 72.135 112.185 ;
        RECT 68.950 111.415 69.410 111.705 ;
        RECT 70.105 111.675 71.605 111.845 ;
        RECT 70.105 111.535 70.275 111.675 ;
        RECT 69.715 111.365 70.275 111.535 ;
        RECT 68.190 110.735 68.440 111.195 ;
        RECT 68.610 110.905 69.480 111.245 ;
        RECT 69.715 110.905 69.885 111.365 ;
        RECT 70.720 111.335 71.795 111.505 ;
        RECT 70.055 110.735 70.425 111.195 ;
        RECT 70.720 110.995 70.890 111.335 ;
        RECT 71.060 110.735 71.390 111.165 ;
        RECT 71.625 110.995 71.795 111.335 ;
        RECT 71.965 111.235 72.135 112.015 ;
        RECT 72.305 111.795 72.475 112.385 ;
        RECT 72.645 111.985 72.995 112.605 ;
        RECT 72.305 111.405 72.770 111.795 ;
        RECT 73.165 111.535 73.335 112.895 ;
        RECT 73.505 111.705 73.965 112.755 ;
        RECT 72.940 111.365 73.335 111.535 ;
        RECT 72.940 111.235 73.110 111.365 ;
        RECT 71.965 110.905 72.645 111.235 ;
        RECT 72.860 110.905 73.110 111.235 ;
        RECT 73.280 110.735 73.530 111.195 ;
        RECT 73.700 110.920 74.025 111.705 ;
        RECT 74.195 110.905 74.365 113.025 ;
        RECT 74.535 112.905 74.865 113.285 ;
        RECT 75.035 112.735 75.290 113.025 ;
        RECT 74.540 112.565 75.290 112.735 ;
        RECT 74.540 111.575 74.770 112.565 ;
        RECT 75.465 112.535 76.675 113.285 ;
        RECT 74.940 111.745 75.290 112.395 ;
        RECT 75.465 111.825 75.985 112.365 ;
        RECT 76.155 111.995 76.675 112.535 ;
        RECT 76.905 112.465 77.115 113.285 ;
        RECT 77.285 112.485 77.615 113.115 ;
        RECT 77.285 111.885 77.535 112.485 ;
        RECT 77.785 112.465 78.015 113.285 ;
        RECT 78.230 112.575 78.485 113.105 ;
        RECT 78.655 112.825 78.960 113.285 ;
        RECT 79.205 112.905 80.275 113.075 ;
        RECT 77.705 112.045 78.035 112.295 ;
        RECT 78.230 111.925 78.440 112.575 ;
        RECT 79.205 112.550 79.525 112.905 ;
        RECT 79.200 112.375 79.525 112.550 ;
        RECT 78.610 112.075 79.525 112.375 ;
        RECT 79.695 112.335 79.935 112.735 ;
        RECT 80.105 112.675 80.275 112.905 ;
        RECT 80.445 112.845 80.635 113.285 ;
        RECT 80.805 112.835 81.755 113.115 ;
        RECT 81.975 112.925 82.325 113.095 ;
        RECT 80.105 112.505 80.635 112.675 ;
        RECT 78.610 112.045 79.350 112.075 ;
        RECT 74.540 111.405 75.290 111.575 ;
        RECT 74.535 110.735 74.865 111.235 ;
        RECT 75.035 110.905 75.290 111.405 ;
        RECT 75.465 110.735 76.675 111.825 ;
        RECT 76.905 110.735 77.115 111.875 ;
        RECT 77.285 110.905 77.615 111.885 ;
        RECT 77.785 110.735 78.015 111.875 ;
        RECT 78.230 111.045 78.485 111.925 ;
        RECT 78.655 110.735 78.960 111.875 ;
        RECT 79.180 111.455 79.350 112.045 ;
        RECT 79.695 111.965 80.235 112.335 ;
        RECT 80.415 112.225 80.635 112.505 ;
        RECT 80.805 112.055 80.975 112.835 ;
        RECT 80.570 111.885 80.975 112.055 ;
        RECT 81.145 112.045 81.495 112.665 ;
        RECT 80.570 111.795 80.740 111.885 ;
        RECT 81.665 111.875 81.875 112.665 ;
        RECT 79.520 111.625 80.740 111.795 ;
        RECT 81.200 111.715 81.875 111.875 ;
        RECT 79.180 111.285 79.980 111.455 ;
        RECT 79.300 110.735 79.630 111.115 ;
        RECT 79.810 110.995 79.980 111.285 ;
        RECT 80.570 111.245 80.740 111.625 ;
        RECT 80.910 111.705 81.875 111.715 ;
        RECT 82.065 112.535 82.325 112.925 ;
        RECT 82.535 112.825 82.865 113.285 ;
        RECT 83.740 112.895 84.595 113.065 ;
        RECT 84.800 112.895 85.295 113.065 ;
        RECT 85.465 112.925 85.795 113.285 ;
        RECT 82.065 111.845 82.235 112.535 ;
        RECT 82.405 112.185 82.575 112.365 ;
        RECT 82.745 112.355 83.535 112.605 ;
        RECT 83.740 112.185 83.910 112.895 ;
        RECT 84.080 112.385 84.435 112.605 ;
        RECT 82.405 112.015 84.095 112.185 ;
        RECT 80.910 111.415 81.370 111.705 ;
        RECT 82.065 111.675 83.565 111.845 ;
        RECT 82.065 111.535 82.235 111.675 ;
        RECT 81.675 111.365 82.235 111.535 ;
        RECT 80.150 110.735 80.400 111.195 ;
        RECT 80.570 110.905 81.440 111.245 ;
        RECT 81.675 110.905 81.845 111.365 ;
        RECT 82.680 111.335 83.755 111.505 ;
        RECT 82.015 110.735 82.385 111.195 ;
        RECT 82.680 110.995 82.850 111.335 ;
        RECT 83.020 110.735 83.350 111.165 ;
        RECT 83.585 110.995 83.755 111.335 ;
        RECT 83.925 111.235 84.095 112.015 ;
        RECT 84.265 111.795 84.435 112.385 ;
        RECT 84.605 111.985 84.955 112.605 ;
        RECT 84.265 111.405 84.730 111.795 ;
        RECT 85.125 111.535 85.295 112.895 ;
        RECT 85.465 111.705 85.925 112.755 ;
        RECT 84.900 111.365 85.295 111.535 ;
        RECT 84.900 111.235 85.070 111.365 ;
        RECT 83.925 110.905 84.605 111.235 ;
        RECT 84.820 110.905 85.070 111.235 ;
        RECT 85.240 110.735 85.490 111.195 ;
        RECT 85.660 110.920 85.985 111.705 ;
        RECT 86.155 110.905 86.325 113.025 ;
        RECT 86.495 112.905 86.825 113.285 ;
        RECT 86.995 112.735 87.250 113.025 ;
        RECT 86.500 112.565 87.250 112.735 ;
        RECT 87.425 112.610 87.685 113.115 ;
        RECT 87.865 112.905 88.195 113.285 ;
        RECT 88.375 112.735 88.545 113.115 ;
        RECT 86.500 111.575 86.730 112.565 ;
        RECT 86.900 111.745 87.250 112.395 ;
        RECT 87.425 111.810 87.595 112.610 ;
        RECT 87.880 112.565 88.545 112.735 ;
        RECT 87.880 112.310 88.050 112.565 ;
        RECT 88.805 112.560 89.095 113.285 ;
        RECT 89.325 112.465 89.535 113.285 ;
        RECT 89.705 112.485 90.035 113.115 ;
        RECT 87.765 111.980 88.050 112.310 ;
        RECT 88.285 112.015 88.615 112.385 ;
        RECT 87.880 111.835 88.050 111.980 ;
        RECT 86.500 111.405 87.250 111.575 ;
        RECT 86.495 110.735 86.825 111.235 ;
        RECT 86.995 110.905 87.250 111.405 ;
        RECT 87.425 110.905 87.695 111.810 ;
        RECT 87.880 111.665 88.545 111.835 ;
        RECT 87.865 110.735 88.195 111.495 ;
        RECT 88.375 110.905 88.545 111.665 ;
        RECT 88.805 110.735 89.095 111.900 ;
        RECT 89.705 111.885 89.955 112.485 ;
        RECT 90.205 112.465 90.435 113.285 ;
        RECT 90.650 112.575 90.905 113.105 ;
        RECT 91.075 112.825 91.380 113.285 ;
        RECT 91.625 112.905 92.695 113.075 ;
        RECT 90.125 112.045 90.455 112.295 ;
        RECT 90.650 111.925 90.860 112.575 ;
        RECT 91.625 112.550 91.945 112.905 ;
        RECT 91.620 112.375 91.945 112.550 ;
        RECT 91.030 112.075 91.945 112.375 ;
        RECT 92.115 112.335 92.355 112.735 ;
        RECT 92.525 112.675 92.695 112.905 ;
        RECT 92.865 112.845 93.055 113.285 ;
        RECT 93.225 112.835 94.175 113.115 ;
        RECT 94.395 112.925 94.745 113.095 ;
        RECT 92.525 112.505 93.055 112.675 ;
        RECT 91.030 112.045 91.770 112.075 ;
        RECT 89.325 110.735 89.535 111.875 ;
        RECT 89.705 110.905 90.035 111.885 ;
        RECT 90.205 110.735 90.435 111.875 ;
        RECT 90.650 111.045 90.905 111.925 ;
        RECT 91.075 110.735 91.380 111.875 ;
        RECT 91.600 111.455 91.770 112.045 ;
        RECT 92.115 111.965 92.655 112.335 ;
        RECT 92.835 112.225 93.055 112.505 ;
        RECT 93.225 112.055 93.395 112.835 ;
        RECT 92.990 111.885 93.395 112.055 ;
        RECT 93.565 112.045 93.915 112.665 ;
        RECT 92.990 111.795 93.160 111.885 ;
        RECT 94.085 111.875 94.295 112.665 ;
        RECT 91.940 111.625 93.160 111.795 ;
        RECT 93.620 111.715 94.295 111.875 ;
        RECT 91.600 111.285 92.400 111.455 ;
        RECT 91.720 110.735 92.050 111.115 ;
        RECT 92.230 110.995 92.400 111.285 ;
        RECT 92.990 111.245 93.160 111.625 ;
        RECT 93.330 111.705 94.295 111.715 ;
        RECT 94.485 112.535 94.745 112.925 ;
        RECT 94.955 112.825 95.285 113.285 ;
        RECT 96.160 112.895 97.015 113.065 ;
        RECT 97.220 112.895 97.715 113.065 ;
        RECT 97.885 112.925 98.215 113.285 ;
        RECT 94.485 111.845 94.655 112.535 ;
        RECT 94.825 112.185 94.995 112.365 ;
        RECT 95.165 112.355 95.955 112.605 ;
        RECT 96.160 112.185 96.330 112.895 ;
        RECT 96.500 112.385 96.855 112.605 ;
        RECT 94.825 112.015 96.515 112.185 ;
        RECT 93.330 111.415 93.790 111.705 ;
        RECT 94.485 111.675 95.985 111.845 ;
        RECT 94.485 111.535 94.655 111.675 ;
        RECT 94.095 111.365 94.655 111.535 ;
        RECT 92.570 110.735 92.820 111.195 ;
        RECT 92.990 110.905 93.860 111.245 ;
        RECT 94.095 110.905 94.265 111.365 ;
        RECT 95.100 111.335 96.175 111.505 ;
        RECT 94.435 110.735 94.805 111.195 ;
        RECT 95.100 110.995 95.270 111.335 ;
        RECT 95.440 110.735 95.770 111.165 ;
        RECT 96.005 110.995 96.175 111.335 ;
        RECT 96.345 111.235 96.515 112.015 ;
        RECT 96.685 111.795 96.855 112.385 ;
        RECT 97.025 111.985 97.375 112.605 ;
        RECT 96.685 111.405 97.150 111.795 ;
        RECT 97.545 111.535 97.715 112.895 ;
        RECT 97.885 111.705 98.345 112.755 ;
        RECT 97.320 111.365 97.715 111.535 ;
        RECT 97.320 111.235 97.490 111.365 ;
        RECT 96.345 110.905 97.025 111.235 ;
        RECT 97.240 110.905 97.490 111.235 ;
        RECT 97.660 110.735 97.910 111.195 ;
        RECT 98.080 110.920 98.405 111.705 ;
        RECT 98.575 110.905 98.745 113.025 ;
        RECT 98.915 112.905 99.245 113.285 ;
        RECT 99.415 112.735 99.670 113.025 ;
        RECT 98.920 112.565 99.670 112.735 ;
        RECT 99.845 112.610 100.105 113.115 ;
        RECT 100.285 112.905 100.615 113.285 ;
        RECT 100.795 112.735 100.965 113.115 ;
        RECT 98.920 111.575 99.150 112.565 ;
        RECT 99.320 111.745 99.670 112.395 ;
        RECT 99.845 111.810 100.015 112.610 ;
        RECT 100.300 112.565 100.965 112.735 ;
        RECT 101.690 112.575 101.945 113.105 ;
        RECT 102.115 112.825 102.420 113.285 ;
        RECT 102.665 112.905 103.735 113.075 ;
        RECT 100.300 112.310 100.470 112.565 ;
        RECT 100.185 111.980 100.470 112.310 ;
        RECT 100.705 112.015 101.035 112.385 ;
        RECT 100.300 111.835 100.470 111.980 ;
        RECT 101.690 111.925 101.900 112.575 ;
        RECT 102.665 112.550 102.985 112.905 ;
        RECT 102.660 112.375 102.985 112.550 ;
        RECT 102.070 112.075 102.985 112.375 ;
        RECT 103.155 112.335 103.395 112.735 ;
        RECT 103.565 112.675 103.735 112.905 ;
        RECT 103.905 112.845 104.095 113.285 ;
        RECT 104.265 112.835 105.215 113.115 ;
        RECT 105.435 112.925 105.785 113.095 ;
        RECT 103.565 112.505 104.095 112.675 ;
        RECT 102.070 112.045 102.810 112.075 ;
        RECT 98.920 111.405 99.670 111.575 ;
        RECT 98.915 110.735 99.245 111.235 ;
        RECT 99.415 110.905 99.670 111.405 ;
        RECT 99.845 110.905 100.115 111.810 ;
        RECT 100.300 111.665 100.965 111.835 ;
        RECT 100.285 110.735 100.615 111.495 ;
        RECT 100.795 110.905 100.965 111.665 ;
        RECT 101.690 111.045 101.945 111.925 ;
        RECT 102.115 110.735 102.420 111.875 ;
        RECT 102.640 111.455 102.810 112.045 ;
        RECT 103.155 111.965 103.695 112.335 ;
        RECT 103.875 112.225 104.095 112.505 ;
        RECT 104.265 112.055 104.435 112.835 ;
        RECT 104.030 111.885 104.435 112.055 ;
        RECT 104.605 112.045 104.955 112.665 ;
        RECT 104.030 111.795 104.200 111.885 ;
        RECT 105.125 111.875 105.335 112.665 ;
        RECT 102.980 111.625 104.200 111.795 ;
        RECT 104.660 111.715 105.335 111.875 ;
        RECT 102.640 111.285 103.440 111.455 ;
        RECT 102.760 110.735 103.090 111.115 ;
        RECT 103.270 110.995 103.440 111.285 ;
        RECT 104.030 111.245 104.200 111.625 ;
        RECT 104.370 111.705 105.335 111.715 ;
        RECT 105.525 112.535 105.785 112.925 ;
        RECT 105.995 112.825 106.325 113.285 ;
        RECT 107.200 112.895 108.055 113.065 ;
        RECT 108.260 112.895 108.755 113.065 ;
        RECT 108.925 112.925 109.255 113.285 ;
        RECT 105.525 111.845 105.695 112.535 ;
        RECT 105.865 112.185 106.035 112.365 ;
        RECT 106.205 112.355 106.995 112.605 ;
        RECT 107.200 112.185 107.370 112.895 ;
        RECT 107.540 112.385 107.895 112.605 ;
        RECT 105.865 112.015 107.555 112.185 ;
        RECT 104.370 111.415 104.830 111.705 ;
        RECT 105.525 111.675 107.025 111.845 ;
        RECT 105.525 111.535 105.695 111.675 ;
        RECT 105.135 111.365 105.695 111.535 ;
        RECT 103.610 110.735 103.860 111.195 ;
        RECT 104.030 110.905 104.900 111.245 ;
        RECT 105.135 110.905 105.305 111.365 ;
        RECT 106.140 111.335 107.215 111.505 ;
        RECT 105.475 110.735 105.845 111.195 ;
        RECT 106.140 110.995 106.310 111.335 ;
        RECT 106.480 110.735 106.810 111.165 ;
        RECT 107.045 110.995 107.215 111.335 ;
        RECT 107.385 111.235 107.555 112.015 ;
        RECT 107.725 111.795 107.895 112.385 ;
        RECT 108.065 111.985 108.415 112.605 ;
        RECT 107.725 111.405 108.190 111.795 ;
        RECT 108.585 111.535 108.755 112.895 ;
        RECT 108.925 111.705 109.385 112.755 ;
        RECT 108.360 111.365 108.755 111.535 ;
        RECT 108.360 111.235 108.530 111.365 ;
        RECT 107.385 110.905 108.065 111.235 ;
        RECT 108.280 110.905 108.530 111.235 ;
        RECT 108.700 110.735 108.950 111.195 ;
        RECT 109.120 110.920 109.445 111.705 ;
        RECT 109.615 110.905 109.785 113.025 ;
        RECT 109.955 112.905 110.285 113.285 ;
        RECT 110.455 112.735 110.710 113.025 ;
        RECT 109.960 112.565 110.710 112.735 ;
        RECT 110.975 112.735 111.145 113.115 ;
        RECT 111.325 112.905 111.655 113.285 ;
        RECT 110.975 112.565 111.640 112.735 ;
        RECT 111.835 112.610 112.095 113.115 ;
        RECT 109.960 111.575 110.190 112.565 ;
        RECT 110.360 111.745 110.710 112.395 ;
        RECT 110.905 112.015 111.235 112.385 ;
        RECT 111.470 112.310 111.640 112.565 ;
        RECT 111.470 111.980 111.755 112.310 ;
        RECT 111.470 111.835 111.640 111.980 ;
        RECT 110.975 111.665 111.640 111.835 ;
        RECT 111.925 111.810 112.095 112.610 ;
        RECT 113.275 112.735 113.445 113.115 ;
        RECT 113.625 112.905 113.955 113.285 ;
        RECT 113.275 112.565 113.940 112.735 ;
        RECT 114.135 112.610 114.395 113.115 ;
        RECT 113.205 112.015 113.535 112.385 ;
        RECT 113.770 112.310 113.940 112.565 ;
        RECT 113.770 111.980 114.055 112.310 ;
        RECT 113.770 111.835 113.940 111.980 ;
        RECT 109.960 111.405 110.710 111.575 ;
        RECT 109.955 110.735 110.285 111.235 ;
        RECT 110.455 110.905 110.710 111.405 ;
        RECT 110.975 110.905 111.145 111.665 ;
        RECT 111.325 110.735 111.655 111.495 ;
        RECT 111.825 110.905 112.095 111.810 ;
        RECT 113.275 111.665 113.940 111.835 ;
        RECT 114.225 111.810 114.395 112.610 ;
        RECT 114.565 112.560 114.855 113.285 ;
        RECT 115.525 112.465 115.755 113.285 ;
        RECT 115.925 112.485 116.255 113.115 ;
        RECT 115.505 112.045 115.835 112.295 ;
        RECT 113.275 110.905 113.445 111.665 ;
        RECT 113.625 110.735 113.955 111.495 ;
        RECT 114.125 110.905 114.395 111.810 ;
        RECT 114.565 110.735 114.855 111.900 ;
        RECT 116.005 111.885 116.255 112.485 ;
        RECT 116.425 112.465 116.635 113.285 ;
        RECT 117.330 112.575 117.585 113.105 ;
        RECT 117.755 112.825 118.060 113.285 ;
        RECT 118.305 112.905 119.375 113.075 ;
        RECT 115.525 110.735 115.755 111.875 ;
        RECT 115.925 110.905 116.255 111.885 ;
        RECT 117.330 111.925 117.540 112.575 ;
        RECT 118.305 112.550 118.625 112.905 ;
        RECT 118.300 112.375 118.625 112.550 ;
        RECT 117.710 112.075 118.625 112.375 ;
        RECT 118.795 112.335 119.035 112.735 ;
        RECT 119.205 112.675 119.375 112.905 ;
        RECT 119.545 112.845 119.735 113.285 ;
        RECT 119.905 112.835 120.855 113.115 ;
        RECT 121.075 112.925 121.425 113.095 ;
        RECT 119.205 112.505 119.735 112.675 ;
        RECT 117.710 112.045 118.450 112.075 ;
        RECT 116.425 110.735 116.635 111.875 ;
        RECT 117.330 111.045 117.585 111.925 ;
        RECT 117.755 110.735 118.060 111.875 ;
        RECT 118.280 111.455 118.450 112.045 ;
        RECT 118.795 111.965 119.335 112.335 ;
        RECT 119.515 112.225 119.735 112.505 ;
        RECT 119.905 112.055 120.075 112.835 ;
        RECT 119.670 111.885 120.075 112.055 ;
        RECT 120.245 112.045 120.595 112.665 ;
        RECT 119.670 111.795 119.840 111.885 ;
        RECT 120.765 111.875 120.975 112.665 ;
        RECT 118.620 111.625 119.840 111.795 ;
        RECT 120.300 111.715 120.975 111.875 ;
        RECT 118.280 111.285 119.080 111.455 ;
        RECT 118.400 110.735 118.730 111.115 ;
        RECT 118.910 110.995 119.080 111.285 ;
        RECT 119.670 111.245 119.840 111.625 ;
        RECT 120.010 111.705 120.975 111.715 ;
        RECT 121.165 112.535 121.425 112.925 ;
        RECT 121.635 112.825 121.965 113.285 ;
        RECT 122.840 112.895 123.695 113.065 ;
        RECT 123.900 112.895 124.395 113.065 ;
        RECT 124.565 112.925 124.895 113.285 ;
        RECT 121.165 111.845 121.335 112.535 ;
        RECT 121.505 112.185 121.675 112.365 ;
        RECT 121.845 112.355 122.635 112.605 ;
        RECT 122.840 112.185 123.010 112.895 ;
        RECT 123.180 112.385 123.535 112.605 ;
        RECT 121.505 112.015 123.195 112.185 ;
        RECT 120.010 111.415 120.470 111.705 ;
        RECT 121.165 111.675 122.665 111.845 ;
        RECT 121.165 111.535 121.335 111.675 ;
        RECT 120.775 111.365 121.335 111.535 ;
        RECT 119.250 110.735 119.500 111.195 ;
        RECT 119.670 110.905 120.540 111.245 ;
        RECT 120.775 110.905 120.945 111.365 ;
        RECT 121.780 111.335 122.855 111.505 ;
        RECT 121.115 110.735 121.485 111.195 ;
        RECT 121.780 110.995 121.950 111.335 ;
        RECT 122.120 110.735 122.450 111.165 ;
        RECT 122.685 110.995 122.855 111.335 ;
        RECT 123.025 111.235 123.195 112.015 ;
        RECT 123.365 111.795 123.535 112.385 ;
        RECT 123.705 111.985 124.055 112.605 ;
        RECT 123.365 111.405 123.830 111.795 ;
        RECT 124.225 111.535 124.395 112.895 ;
        RECT 124.565 111.705 125.025 112.755 ;
        RECT 124.000 111.365 124.395 111.535 ;
        RECT 124.000 111.235 124.170 111.365 ;
        RECT 123.025 110.905 123.705 111.235 ;
        RECT 123.920 110.905 124.170 111.235 ;
        RECT 124.340 110.735 124.590 111.195 ;
        RECT 124.760 110.920 125.085 111.705 ;
        RECT 125.255 110.905 125.425 113.025 ;
        RECT 125.595 112.905 125.925 113.285 ;
        RECT 126.095 112.735 126.350 113.025 ;
        RECT 125.600 112.565 126.350 112.735 ;
        RECT 125.600 111.575 125.830 112.565 ;
        RECT 126.525 112.535 127.735 113.285 ;
        RECT 126.000 111.745 126.350 112.395 ;
        RECT 126.525 111.825 127.045 112.365 ;
        RECT 127.215 111.995 127.735 112.535 ;
        RECT 125.600 111.405 126.350 111.575 ;
        RECT 125.595 110.735 125.925 111.235 ;
        RECT 126.095 110.905 126.350 111.405 ;
        RECT 126.525 110.735 127.735 111.825 ;
        RECT 20.640 110.565 127.820 110.735 ;
        RECT 20.725 109.475 21.935 110.565 ;
        RECT 20.725 108.765 21.245 109.305 ;
        RECT 21.415 108.935 21.935 109.475 ;
        RECT 22.565 109.475 24.235 110.565 ;
        RECT 22.565 108.955 23.315 109.475 ;
        RECT 24.405 109.400 24.695 110.565 ;
        RECT 24.870 110.130 30.215 110.565 ;
        RECT 23.485 108.785 24.235 109.305 ;
        RECT 26.460 108.880 26.810 110.130 ;
        RECT 30.475 109.635 30.645 110.395 ;
        RECT 30.825 109.805 31.155 110.565 ;
        RECT 30.475 109.465 31.140 109.635 ;
        RECT 31.325 109.490 31.595 110.395 ;
        RECT 31.770 109.895 32.025 110.395 ;
        RECT 32.195 110.065 32.525 110.565 ;
        RECT 31.770 109.725 32.520 109.895 ;
        RECT 20.725 108.015 21.935 108.765 ;
        RECT 22.565 108.015 24.235 108.785 ;
        RECT 24.405 108.015 24.695 108.740 ;
        RECT 28.290 108.560 28.630 109.390 ;
        RECT 30.970 109.320 31.140 109.465 ;
        RECT 30.405 108.915 30.735 109.285 ;
        RECT 30.970 108.990 31.255 109.320 ;
        RECT 30.970 108.735 31.140 108.990 ;
        RECT 30.475 108.565 31.140 108.735 ;
        RECT 31.425 108.690 31.595 109.490 ;
        RECT 31.770 108.905 32.120 109.555 ;
        RECT 32.290 108.735 32.520 109.725 ;
        RECT 24.870 108.015 30.215 108.560 ;
        RECT 30.475 108.185 30.645 108.565 ;
        RECT 30.825 108.015 31.155 108.395 ;
        RECT 31.335 108.185 31.595 108.690 ;
        RECT 31.770 108.565 32.520 108.735 ;
        RECT 31.770 108.275 32.025 108.565 ;
        RECT 32.195 108.015 32.525 108.395 ;
        RECT 32.695 108.275 32.865 110.395 ;
        RECT 33.035 109.595 33.360 110.380 ;
        RECT 33.530 110.105 33.780 110.565 ;
        RECT 33.950 110.065 34.200 110.395 ;
        RECT 34.415 110.065 35.095 110.395 ;
        RECT 33.950 109.935 34.120 110.065 ;
        RECT 33.725 109.765 34.120 109.935 ;
        RECT 33.095 108.545 33.555 109.595 ;
        RECT 33.725 108.405 33.895 109.765 ;
        RECT 34.290 109.505 34.755 109.895 ;
        RECT 34.065 108.695 34.415 109.315 ;
        RECT 34.585 108.915 34.755 109.505 ;
        RECT 34.925 109.285 35.095 110.065 ;
        RECT 35.265 109.965 35.435 110.305 ;
        RECT 35.670 110.135 36.000 110.565 ;
        RECT 36.170 109.965 36.340 110.305 ;
        RECT 36.635 110.105 37.005 110.565 ;
        RECT 35.265 109.795 36.340 109.965 ;
        RECT 37.175 109.935 37.345 110.395 ;
        RECT 37.580 110.055 38.450 110.395 ;
        RECT 38.620 110.105 38.870 110.565 ;
        RECT 36.785 109.765 37.345 109.935 ;
        RECT 36.785 109.625 36.955 109.765 ;
        RECT 35.455 109.455 36.955 109.625 ;
        RECT 37.650 109.595 38.110 109.885 ;
        RECT 34.925 109.115 36.615 109.285 ;
        RECT 34.585 108.695 34.940 108.915 ;
        RECT 35.110 108.405 35.280 109.115 ;
        RECT 35.485 108.695 36.275 108.945 ;
        RECT 36.445 108.935 36.615 109.115 ;
        RECT 36.785 108.765 36.955 109.455 ;
        RECT 33.225 108.015 33.555 108.375 ;
        RECT 33.725 108.235 34.220 108.405 ;
        RECT 34.425 108.235 35.280 108.405 ;
        RECT 36.155 108.015 36.485 108.475 ;
        RECT 36.695 108.375 36.955 108.765 ;
        RECT 37.145 109.585 38.110 109.595 ;
        RECT 38.280 109.675 38.450 110.055 ;
        RECT 39.040 110.015 39.210 110.305 ;
        RECT 39.390 110.185 39.720 110.565 ;
        RECT 39.040 109.845 39.840 110.015 ;
        RECT 37.145 109.425 37.820 109.585 ;
        RECT 38.280 109.505 39.500 109.675 ;
        RECT 37.145 108.635 37.355 109.425 ;
        RECT 38.280 109.415 38.450 109.505 ;
        RECT 37.525 108.635 37.875 109.255 ;
        RECT 38.045 109.245 38.450 109.415 ;
        RECT 38.045 108.465 38.215 109.245 ;
        RECT 38.385 108.795 38.605 109.075 ;
        RECT 38.785 108.965 39.325 109.335 ;
        RECT 39.670 109.255 39.840 109.845 ;
        RECT 40.060 109.425 40.365 110.565 ;
        RECT 40.535 109.375 40.790 110.255 ;
        RECT 40.970 109.895 41.225 110.395 ;
        RECT 41.395 110.065 41.725 110.565 ;
        RECT 40.970 109.725 41.720 109.895 ;
        RECT 39.670 109.225 40.410 109.255 ;
        RECT 38.385 108.625 38.915 108.795 ;
        RECT 36.695 108.205 37.045 108.375 ;
        RECT 37.265 108.185 38.215 108.465 ;
        RECT 38.385 108.015 38.575 108.455 ;
        RECT 38.745 108.395 38.915 108.625 ;
        RECT 39.085 108.565 39.325 108.965 ;
        RECT 39.495 108.925 40.410 109.225 ;
        RECT 39.495 108.750 39.820 108.925 ;
        RECT 39.495 108.395 39.815 108.750 ;
        RECT 40.580 108.725 40.790 109.375 ;
        RECT 40.970 108.905 41.320 109.555 ;
        RECT 41.490 108.735 41.720 109.725 ;
        RECT 38.745 108.225 39.815 108.395 ;
        RECT 40.060 108.015 40.365 108.475 ;
        RECT 40.535 108.195 40.790 108.725 ;
        RECT 40.970 108.565 41.720 108.735 ;
        RECT 40.970 108.275 41.225 108.565 ;
        RECT 41.395 108.015 41.725 108.395 ;
        RECT 41.895 108.275 42.065 110.395 ;
        RECT 42.235 109.595 42.560 110.380 ;
        RECT 42.730 110.105 42.980 110.565 ;
        RECT 43.150 110.065 43.400 110.395 ;
        RECT 43.615 110.065 44.295 110.395 ;
        RECT 43.150 109.935 43.320 110.065 ;
        RECT 42.925 109.765 43.320 109.935 ;
        RECT 42.295 108.545 42.755 109.595 ;
        RECT 42.925 108.405 43.095 109.765 ;
        RECT 43.490 109.505 43.955 109.895 ;
        RECT 43.265 108.695 43.615 109.315 ;
        RECT 43.785 108.915 43.955 109.505 ;
        RECT 44.125 109.285 44.295 110.065 ;
        RECT 44.465 109.965 44.635 110.305 ;
        RECT 44.870 110.135 45.200 110.565 ;
        RECT 45.370 109.965 45.540 110.305 ;
        RECT 45.835 110.105 46.205 110.565 ;
        RECT 44.465 109.795 45.540 109.965 ;
        RECT 46.375 109.935 46.545 110.395 ;
        RECT 46.780 110.055 47.650 110.395 ;
        RECT 47.820 110.105 48.070 110.565 ;
        RECT 45.985 109.765 46.545 109.935 ;
        RECT 45.985 109.625 46.155 109.765 ;
        RECT 44.655 109.455 46.155 109.625 ;
        RECT 46.850 109.595 47.310 109.885 ;
        RECT 44.125 109.115 45.815 109.285 ;
        RECT 43.785 108.695 44.140 108.915 ;
        RECT 44.310 108.405 44.480 109.115 ;
        RECT 44.685 108.695 45.475 108.945 ;
        RECT 45.645 108.935 45.815 109.115 ;
        RECT 45.985 108.765 46.155 109.455 ;
        RECT 42.425 108.015 42.755 108.375 ;
        RECT 42.925 108.235 43.420 108.405 ;
        RECT 43.625 108.235 44.480 108.405 ;
        RECT 45.355 108.015 45.685 108.475 ;
        RECT 45.895 108.375 46.155 108.765 ;
        RECT 46.345 109.585 47.310 109.595 ;
        RECT 47.480 109.675 47.650 110.055 ;
        RECT 48.240 110.015 48.410 110.305 ;
        RECT 48.590 110.185 48.920 110.565 ;
        RECT 48.240 109.845 49.040 110.015 ;
        RECT 46.345 109.425 47.020 109.585 ;
        RECT 47.480 109.505 48.700 109.675 ;
        RECT 46.345 108.635 46.555 109.425 ;
        RECT 47.480 109.415 47.650 109.505 ;
        RECT 46.725 108.635 47.075 109.255 ;
        RECT 47.245 109.245 47.650 109.415 ;
        RECT 47.245 108.465 47.415 109.245 ;
        RECT 47.585 108.795 47.805 109.075 ;
        RECT 47.985 108.965 48.525 109.335 ;
        RECT 48.870 109.255 49.040 109.845 ;
        RECT 49.260 109.425 49.565 110.565 ;
        RECT 49.735 109.375 49.990 110.255 ;
        RECT 50.165 109.400 50.455 110.565 ;
        RECT 51.085 109.475 53.675 110.565 ;
        RECT 48.870 109.225 49.610 109.255 ;
        RECT 47.585 108.625 48.115 108.795 ;
        RECT 45.895 108.205 46.245 108.375 ;
        RECT 46.465 108.185 47.415 108.465 ;
        RECT 47.585 108.015 47.775 108.455 ;
        RECT 47.945 108.395 48.115 108.625 ;
        RECT 48.285 108.565 48.525 108.965 ;
        RECT 48.695 108.925 49.610 109.225 ;
        RECT 48.695 108.750 49.020 108.925 ;
        RECT 48.695 108.395 49.015 108.750 ;
        RECT 49.780 108.725 49.990 109.375 ;
        RECT 51.085 108.955 52.295 109.475 ;
        RECT 53.885 109.425 54.115 110.565 ;
        RECT 54.285 109.415 54.615 110.395 ;
        RECT 54.785 109.425 54.995 110.565 ;
        RECT 55.265 109.425 55.495 110.565 ;
        RECT 55.665 109.415 55.995 110.395 ;
        RECT 56.165 109.425 56.375 110.565 ;
        RECT 52.465 108.785 53.675 109.305 ;
        RECT 53.865 109.005 54.195 109.255 ;
        RECT 47.945 108.225 49.015 108.395 ;
        RECT 49.260 108.015 49.565 108.475 ;
        RECT 49.735 108.195 49.990 108.725 ;
        RECT 50.165 108.015 50.455 108.740 ;
        RECT 51.085 108.015 53.675 108.785 ;
        RECT 53.885 108.015 54.115 108.835 ;
        RECT 54.365 108.815 54.615 109.415 ;
        RECT 55.245 109.005 55.575 109.255 ;
        RECT 54.285 108.185 54.615 108.815 ;
        RECT 54.785 108.015 54.995 108.835 ;
        RECT 55.265 108.015 55.495 108.835 ;
        RECT 55.745 108.815 55.995 109.415 ;
        RECT 56.610 109.375 56.865 110.255 ;
        RECT 57.035 109.425 57.340 110.565 ;
        RECT 57.680 110.185 58.010 110.565 ;
        RECT 58.190 110.015 58.360 110.305 ;
        RECT 58.530 110.105 58.780 110.565 ;
        RECT 57.560 109.845 58.360 110.015 ;
        RECT 58.950 110.055 59.820 110.395 ;
        RECT 55.665 108.185 55.995 108.815 ;
        RECT 56.165 108.015 56.375 108.835 ;
        RECT 56.610 108.725 56.820 109.375 ;
        RECT 57.560 109.255 57.730 109.845 ;
        RECT 58.950 109.675 59.120 110.055 ;
        RECT 60.055 109.935 60.225 110.395 ;
        RECT 60.395 110.105 60.765 110.565 ;
        RECT 61.060 109.965 61.230 110.305 ;
        RECT 61.400 110.135 61.730 110.565 ;
        RECT 61.965 109.965 62.135 110.305 ;
        RECT 57.900 109.505 59.120 109.675 ;
        RECT 59.290 109.595 59.750 109.885 ;
        RECT 60.055 109.765 60.615 109.935 ;
        RECT 61.060 109.795 62.135 109.965 ;
        RECT 62.305 110.065 62.985 110.395 ;
        RECT 63.200 110.065 63.450 110.395 ;
        RECT 63.620 110.105 63.870 110.565 ;
        RECT 60.445 109.625 60.615 109.765 ;
        RECT 59.290 109.585 60.255 109.595 ;
        RECT 58.950 109.415 59.120 109.505 ;
        RECT 59.580 109.425 60.255 109.585 ;
        RECT 56.990 109.225 57.730 109.255 ;
        RECT 56.990 108.925 57.905 109.225 ;
        RECT 57.580 108.750 57.905 108.925 ;
        RECT 56.610 108.195 56.865 108.725 ;
        RECT 57.035 108.015 57.340 108.475 ;
        RECT 57.585 108.395 57.905 108.750 ;
        RECT 58.075 108.965 58.615 109.335 ;
        RECT 58.950 109.245 59.355 109.415 ;
        RECT 58.075 108.565 58.315 108.965 ;
        RECT 58.795 108.795 59.015 109.075 ;
        RECT 58.485 108.625 59.015 108.795 ;
        RECT 58.485 108.395 58.655 108.625 ;
        RECT 59.185 108.465 59.355 109.245 ;
        RECT 59.525 108.635 59.875 109.255 ;
        RECT 60.045 108.635 60.255 109.425 ;
        RECT 60.445 109.455 61.945 109.625 ;
        RECT 60.445 108.765 60.615 109.455 ;
        RECT 62.305 109.285 62.475 110.065 ;
        RECT 63.280 109.935 63.450 110.065 ;
        RECT 60.785 109.115 62.475 109.285 ;
        RECT 62.645 109.505 63.110 109.895 ;
        RECT 63.280 109.765 63.675 109.935 ;
        RECT 60.785 108.935 60.955 109.115 ;
        RECT 57.585 108.225 58.655 108.395 ;
        RECT 58.825 108.015 59.015 108.455 ;
        RECT 59.185 108.185 60.135 108.465 ;
        RECT 60.445 108.375 60.705 108.765 ;
        RECT 61.125 108.695 61.915 108.945 ;
        RECT 60.355 108.205 60.705 108.375 ;
        RECT 60.915 108.015 61.245 108.475 ;
        RECT 62.120 108.405 62.290 109.115 ;
        RECT 62.645 108.915 62.815 109.505 ;
        RECT 62.460 108.695 62.815 108.915 ;
        RECT 62.985 108.695 63.335 109.315 ;
        RECT 63.505 108.405 63.675 109.765 ;
        RECT 64.040 109.595 64.365 110.380 ;
        RECT 63.845 108.545 64.305 109.595 ;
        RECT 62.120 108.235 62.975 108.405 ;
        RECT 63.180 108.235 63.675 108.405 ;
        RECT 63.845 108.015 64.175 108.375 ;
        RECT 64.535 108.275 64.705 110.395 ;
        RECT 64.875 110.065 65.205 110.565 ;
        RECT 65.375 109.895 65.630 110.395 ;
        RECT 64.880 109.725 65.630 109.895 ;
        RECT 64.880 108.735 65.110 109.725 ;
        RECT 65.280 108.905 65.630 109.555 ;
        RECT 65.810 109.375 66.065 110.255 ;
        RECT 66.235 109.425 66.540 110.565 ;
        RECT 66.880 110.185 67.210 110.565 ;
        RECT 67.390 110.015 67.560 110.305 ;
        RECT 67.730 110.105 67.980 110.565 ;
        RECT 66.760 109.845 67.560 110.015 ;
        RECT 68.150 110.055 69.020 110.395 ;
        RECT 64.880 108.565 65.630 108.735 ;
        RECT 64.875 108.015 65.205 108.395 ;
        RECT 65.375 108.275 65.630 108.565 ;
        RECT 65.810 108.725 66.020 109.375 ;
        RECT 66.760 109.255 66.930 109.845 ;
        RECT 68.150 109.675 68.320 110.055 ;
        RECT 69.255 109.935 69.425 110.395 ;
        RECT 69.595 110.105 69.965 110.565 ;
        RECT 70.260 109.965 70.430 110.305 ;
        RECT 70.600 110.135 70.930 110.565 ;
        RECT 71.165 109.965 71.335 110.305 ;
        RECT 67.100 109.505 68.320 109.675 ;
        RECT 68.490 109.595 68.950 109.885 ;
        RECT 69.255 109.765 69.815 109.935 ;
        RECT 70.260 109.795 71.335 109.965 ;
        RECT 71.505 110.065 72.185 110.395 ;
        RECT 72.400 110.065 72.650 110.395 ;
        RECT 72.820 110.105 73.070 110.565 ;
        RECT 69.645 109.625 69.815 109.765 ;
        RECT 68.490 109.585 69.455 109.595 ;
        RECT 68.150 109.415 68.320 109.505 ;
        RECT 68.780 109.425 69.455 109.585 ;
        RECT 66.190 109.225 66.930 109.255 ;
        RECT 66.190 108.925 67.105 109.225 ;
        RECT 66.780 108.750 67.105 108.925 ;
        RECT 65.810 108.195 66.065 108.725 ;
        RECT 66.235 108.015 66.540 108.475 ;
        RECT 66.785 108.395 67.105 108.750 ;
        RECT 67.275 108.965 67.815 109.335 ;
        RECT 68.150 109.245 68.555 109.415 ;
        RECT 67.275 108.565 67.515 108.965 ;
        RECT 67.995 108.795 68.215 109.075 ;
        RECT 67.685 108.625 68.215 108.795 ;
        RECT 67.685 108.395 67.855 108.625 ;
        RECT 68.385 108.465 68.555 109.245 ;
        RECT 68.725 108.635 69.075 109.255 ;
        RECT 69.245 108.635 69.455 109.425 ;
        RECT 69.645 109.455 71.145 109.625 ;
        RECT 69.645 108.765 69.815 109.455 ;
        RECT 71.505 109.285 71.675 110.065 ;
        RECT 72.480 109.935 72.650 110.065 ;
        RECT 69.985 109.115 71.675 109.285 ;
        RECT 71.845 109.505 72.310 109.895 ;
        RECT 72.480 109.765 72.875 109.935 ;
        RECT 69.985 108.935 70.155 109.115 ;
        RECT 66.785 108.225 67.855 108.395 ;
        RECT 68.025 108.015 68.215 108.455 ;
        RECT 68.385 108.185 69.335 108.465 ;
        RECT 69.645 108.375 69.905 108.765 ;
        RECT 70.325 108.695 71.115 108.945 ;
        RECT 69.555 108.205 69.905 108.375 ;
        RECT 70.115 108.015 70.445 108.475 ;
        RECT 71.320 108.405 71.490 109.115 ;
        RECT 71.845 108.915 72.015 109.505 ;
        RECT 71.660 108.695 72.015 108.915 ;
        RECT 72.185 108.695 72.535 109.315 ;
        RECT 72.705 108.405 72.875 109.765 ;
        RECT 73.240 109.595 73.565 110.380 ;
        RECT 73.045 108.545 73.505 109.595 ;
        RECT 71.320 108.235 72.175 108.405 ;
        RECT 72.380 108.235 72.875 108.405 ;
        RECT 73.045 108.015 73.375 108.375 ;
        RECT 73.735 108.275 73.905 110.395 ;
        RECT 74.075 110.065 74.405 110.565 ;
        RECT 74.575 109.895 74.830 110.395 ;
        RECT 74.080 109.725 74.830 109.895 ;
        RECT 74.080 108.735 74.310 109.725 ;
        RECT 74.480 108.905 74.830 109.555 ;
        RECT 75.925 109.400 76.215 110.565 ;
        RECT 76.390 109.375 76.645 110.255 ;
        RECT 76.815 109.425 77.120 110.565 ;
        RECT 77.460 110.185 77.790 110.565 ;
        RECT 77.970 110.015 78.140 110.305 ;
        RECT 78.310 110.105 78.560 110.565 ;
        RECT 77.340 109.845 78.140 110.015 ;
        RECT 78.730 110.055 79.600 110.395 ;
        RECT 74.080 108.565 74.830 108.735 ;
        RECT 74.075 108.015 74.405 108.395 ;
        RECT 74.575 108.275 74.830 108.565 ;
        RECT 75.925 108.015 76.215 108.740 ;
        RECT 76.390 108.725 76.600 109.375 ;
        RECT 77.340 109.255 77.510 109.845 ;
        RECT 78.730 109.675 78.900 110.055 ;
        RECT 79.835 109.935 80.005 110.395 ;
        RECT 80.175 110.105 80.545 110.565 ;
        RECT 80.840 109.965 81.010 110.305 ;
        RECT 81.180 110.135 81.510 110.565 ;
        RECT 81.745 109.965 81.915 110.305 ;
        RECT 77.680 109.505 78.900 109.675 ;
        RECT 79.070 109.595 79.530 109.885 ;
        RECT 79.835 109.765 80.395 109.935 ;
        RECT 80.840 109.795 81.915 109.965 ;
        RECT 82.085 110.065 82.765 110.395 ;
        RECT 82.980 110.065 83.230 110.395 ;
        RECT 83.400 110.105 83.650 110.565 ;
        RECT 80.225 109.625 80.395 109.765 ;
        RECT 79.070 109.585 80.035 109.595 ;
        RECT 78.730 109.415 78.900 109.505 ;
        RECT 79.360 109.425 80.035 109.585 ;
        RECT 76.770 109.225 77.510 109.255 ;
        RECT 76.770 108.925 77.685 109.225 ;
        RECT 77.360 108.750 77.685 108.925 ;
        RECT 76.390 108.195 76.645 108.725 ;
        RECT 76.815 108.015 77.120 108.475 ;
        RECT 77.365 108.395 77.685 108.750 ;
        RECT 77.855 108.965 78.395 109.335 ;
        RECT 78.730 109.245 79.135 109.415 ;
        RECT 77.855 108.565 78.095 108.965 ;
        RECT 78.575 108.795 78.795 109.075 ;
        RECT 78.265 108.625 78.795 108.795 ;
        RECT 78.265 108.395 78.435 108.625 ;
        RECT 78.965 108.465 79.135 109.245 ;
        RECT 79.305 108.635 79.655 109.255 ;
        RECT 79.825 108.635 80.035 109.425 ;
        RECT 80.225 109.455 81.725 109.625 ;
        RECT 80.225 108.765 80.395 109.455 ;
        RECT 82.085 109.285 82.255 110.065 ;
        RECT 83.060 109.935 83.230 110.065 ;
        RECT 80.565 109.115 82.255 109.285 ;
        RECT 82.425 109.505 82.890 109.895 ;
        RECT 83.060 109.765 83.455 109.935 ;
        RECT 80.565 108.935 80.735 109.115 ;
        RECT 77.365 108.225 78.435 108.395 ;
        RECT 78.605 108.015 78.795 108.455 ;
        RECT 78.965 108.185 79.915 108.465 ;
        RECT 80.225 108.375 80.485 108.765 ;
        RECT 80.905 108.695 81.695 108.945 ;
        RECT 80.135 108.205 80.485 108.375 ;
        RECT 80.695 108.015 81.025 108.475 ;
        RECT 81.900 108.405 82.070 109.115 ;
        RECT 82.425 108.915 82.595 109.505 ;
        RECT 82.240 108.695 82.595 108.915 ;
        RECT 82.765 108.695 83.115 109.315 ;
        RECT 83.285 108.405 83.455 109.765 ;
        RECT 83.820 109.595 84.145 110.380 ;
        RECT 83.625 108.545 84.085 109.595 ;
        RECT 81.900 108.235 82.755 108.405 ;
        RECT 82.960 108.235 83.455 108.405 ;
        RECT 83.625 108.015 83.955 108.375 ;
        RECT 84.315 108.275 84.485 110.395 ;
        RECT 84.655 110.065 84.985 110.565 ;
        RECT 85.155 109.895 85.410 110.395 ;
        RECT 84.660 109.725 85.410 109.895 ;
        RECT 85.590 109.895 85.845 110.395 ;
        RECT 86.015 110.065 86.345 110.565 ;
        RECT 85.590 109.725 86.340 109.895 ;
        RECT 84.660 108.735 84.890 109.725 ;
        RECT 85.060 108.905 85.410 109.555 ;
        RECT 85.590 108.905 85.940 109.555 ;
        RECT 86.110 108.735 86.340 109.725 ;
        RECT 84.660 108.565 85.410 108.735 ;
        RECT 84.655 108.015 84.985 108.395 ;
        RECT 85.155 108.275 85.410 108.565 ;
        RECT 85.590 108.565 86.340 108.735 ;
        RECT 85.590 108.275 85.845 108.565 ;
        RECT 86.015 108.015 86.345 108.395 ;
        RECT 86.515 108.275 86.685 110.395 ;
        RECT 86.855 109.595 87.180 110.380 ;
        RECT 87.350 110.105 87.600 110.565 ;
        RECT 87.770 110.065 88.020 110.395 ;
        RECT 88.235 110.065 88.915 110.395 ;
        RECT 87.770 109.935 87.940 110.065 ;
        RECT 87.545 109.765 87.940 109.935 ;
        RECT 86.915 108.545 87.375 109.595 ;
        RECT 87.545 108.405 87.715 109.765 ;
        RECT 88.110 109.505 88.575 109.895 ;
        RECT 87.885 108.695 88.235 109.315 ;
        RECT 88.405 108.915 88.575 109.505 ;
        RECT 88.745 109.285 88.915 110.065 ;
        RECT 89.085 109.965 89.255 110.305 ;
        RECT 89.490 110.135 89.820 110.565 ;
        RECT 89.990 109.965 90.160 110.305 ;
        RECT 90.455 110.105 90.825 110.565 ;
        RECT 89.085 109.795 90.160 109.965 ;
        RECT 90.995 109.935 91.165 110.395 ;
        RECT 91.400 110.055 92.270 110.395 ;
        RECT 92.440 110.105 92.690 110.565 ;
        RECT 90.605 109.765 91.165 109.935 ;
        RECT 90.605 109.625 90.775 109.765 ;
        RECT 89.275 109.455 90.775 109.625 ;
        RECT 91.470 109.595 91.930 109.885 ;
        RECT 88.745 109.115 90.435 109.285 ;
        RECT 88.405 108.695 88.760 108.915 ;
        RECT 88.930 108.405 89.100 109.115 ;
        RECT 89.305 108.695 90.095 108.945 ;
        RECT 90.265 108.935 90.435 109.115 ;
        RECT 90.605 108.765 90.775 109.455 ;
        RECT 87.045 108.015 87.375 108.375 ;
        RECT 87.545 108.235 88.040 108.405 ;
        RECT 88.245 108.235 89.100 108.405 ;
        RECT 89.975 108.015 90.305 108.475 ;
        RECT 90.515 108.375 90.775 108.765 ;
        RECT 90.965 109.585 91.930 109.595 ;
        RECT 92.100 109.675 92.270 110.055 ;
        RECT 92.860 110.015 93.030 110.305 ;
        RECT 93.210 110.185 93.540 110.565 ;
        RECT 92.860 109.845 93.660 110.015 ;
        RECT 90.965 109.425 91.640 109.585 ;
        RECT 92.100 109.505 93.320 109.675 ;
        RECT 90.965 108.635 91.175 109.425 ;
        RECT 92.100 109.415 92.270 109.505 ;
        RECT 91.345 108.635 91.695 109.255 ;
        RECT 91.865 109.245 92.270 109.415 ;
        RECT 91.865 108.465 92.035 109.245 ;
        RECT 92.205 108.795 92.425 109.075 ;
        RECT 92.605 108.965 93.145 109.335 ;
        RECT 93.490 109.255 93.660 109.845 ;
        RECT 93.880 109.425 94.185 110.565 ;
        RECT 94.355 109.375 94.610 110.255 ;
        RECT 93.490 109.225 94.230 109.255 ;
        RECT 92.205 108.625 92.735 108.795 ;
        RECT 90.515 108.205 90.865 108.375 ;
        RECT 91.085 108.185 92.035 108.465 ;
        RECT 92.205 108.015 92.395 108.455 ;
        RECT 92.565 108.395 92.735 108.625 ;
        RECT 92.905 108.565 93.145 108.965 ;
        RECT 93.315 108.925 94.230 109.225 ;
        RECT 93.315 108.750 93.640 108.925 ;
        RECT 93.315 108.395 93.635 108.750 ;
        RECT 94.400 108.725 94.610 109.375 ;
        RECT 94.785 109.475 95.995 110.565 ;
        RECT 96.170 110.130 101.515 110.565 ;
        RECT 94.785 108.935 95.305 109.475 ;
        RECT 95.475 108.765 95.995 109.305 ;
        RECT 97.760 108.880 98.110 110.130 ;
        RECT 101.685 109.400 101.975 110.565 ;
        RECT 102.605 109.475 105.195 110.565 ;
        RECT 92.565 108.225 93.635 108.395 ;
        RECT 93.880 108.015 94.185 108.475 ;
        RECT 94.355 108.195 94.610 108.725 ;
        RECT 94.785 108.015 95.995 108.765 ;
        RECT 99.590 108.560 99.930 109.390 ;
        RECT 102.605 108.955 103.815 109.475 ;
        RECT 105.370 109.375 105.625 110.255 ;
        RECT 105.795 109.425 106.100 110.565 ;
        RECT 106.440 110.185 106.770 110.565 ;
        RECT 106.950 110.015 107.120 110.305 ;
        RECT 107.290 110.105 107.540 110.565 ;
        RECT 106.320 109.845 107.120 110.015 ;
        RECT 107.710 110.055 108.580 110.395 ;
        RECT 103.985 108.785 105.195 109.305 ;
        RECT 96.170 108.015 101.515 108.560 ;
        RECT 101.685 108.015 101.975 108.740 ;
        RECT 102.605 108.015 105.195 108.785 ;
        RECT 105.370 108.725 105.580 109.375 ;
        RECT 106.320 109.255 106.490 109.845 ;
        RECT 107.710 109.675 107.880 110.055 ;
        RECT 108.815 109.935 108.985 110.395 ;
        RECT 109.155 110.105 109.525 110.565 ;
        RECT 109.820 109.965 109.990 110.305 ;
        RECT 110.160 110.135 110.490 110.565 ;
        RECT 110.725 109.965 110.895 110.305 ;
        RECT 106.660 109.505 107.880 109.675 ;
        RECT 108.050 109.595 108.510 109.885 ;
        RECT 108.815 109.765 109.375 109.935 ;
        RECT 109.820 109.795 110.895 109.965 ;
        RECT 111.065 110.065 111.745 110.395 ;
        RECT 111.960 110.065 112.210 110.395 ;
        RECT 112.380 110.105 112.630 110.565 ;
        RECT 109.205 109.625 109.375 109.765 ;
        RECT 108.050 109.585 109.015 109.595 ;
        RECT 107.710 109.415 107.880 109.505 ;
        RECT 108.340 109.425 109.015 109.585 ;
        RECT 105.750 109.225 106.490 109.255 ;
        RECT 105.750 108.925 106.665 109.225 ;
        RECT 106.340 108.750 106.665 108.925 ;
        RECT 105.370 108.195 105.625 108.725 ;
        RECT 105.795 108.015 106.100 108.475 ;
        RECT 106.345 108.395 106.665 108.750 ;
        RECT 106.835 108.965 107.375 109.335 ;
        RECT 107.710 109.245 108.115 109.415 ;
        RECT 106.835 108.565 107.075 108.965 ;
        RECT 107.555 108.795 107.775 109.075 ;
        RECT 107.245 108.625 107.775 108.795 ;
        RECT 107.245 108.395 107.415 108.625 ;
        RECT 107.945 108.465 108.115 109.245 ;
        RECT 108.285 108.635 108.635 109.255 ;
        RECT 108.805 108.635 109.015 109.425 ;
        RECT 109.205 109.455 110.705 109.625 ;
        RECT 109.205 108.765 109.375 109.455 ;
        RECT 111.065 109.285 111.235 110.065 ;
        RECT 112.040 109.935 112.210 110.065 ;
        RECT 109.545 109.115 111.235 109.285 ;
        RECT 111.405 109.505 111.870 109.895 ;
        RECT 112.040 109.765 112.435 109.935 ;
        RECT 109.545 108.935 109.715 109.115 ;
        RECT 106.345 108.225 107.415 108.395 ;
        RECT 107.585 108.015 107.775 108.455 ;
        RECT 107.945 108.185 108.895 108.465 ;
        RECT 109.205 108.375 109.465 108.765 ;
        RECT 109.885 108.695 110.675 108.945 ;
        RECT 109.115 108.205 109.465 108.375 ;
        RECT 109.675 108.015 110.005 108.475 ;
        RECT 110.880 108.405 111.050 109.115 ;
        RECT 111.405 108.915 111.575 109.505 ;
        RECT 111.220 108.695 111.575 108.915 ;
        RECT 111.745 108.695 112.095 109.315 ;
        RECT 112.265 108.405 112.435 109.765 ;
        RECT 112.800 109.595 113.125 110.380 ;
        RECT 112.605 108.545 113.065 109.595 ;
        RECT 110.880 108.235 111.735 108.405 ;
        RECT 111.940 108.235 112.435 108.405 ;
        RECT 112.605 108.015 112.935 108.375 ;
        RECT 113.295 108.275 113.465 110.395 ;
        RECT 113.635 110.065 113.965 110.565 ;
        RECT 114.135 109.895 114.390 110.395 ;
        RECT 113.640 109.725 114.390 109.895 ;
        RECT 113.640 108.735 113.870 109.725 ;
        RECT 114.040 108.905 114.390 109.555 ;
        RECT 114.570 109.375 114.825 110.255 ;
        RECT 114.995 109.425 115.300 110.565 ;
        RECT 115.640 110.185 115.970 110.565 ;
        RECT 116.150 110.015 116.320 110.305 ;
        RECT 116.490 110.105 116.740 110.565 ;
        RECT 115.520 109.845 116.320 110.015 ;
        RECT 116.910 110.055 117.780 110.395 ;
        RECT 113.640 108.565 114.390 108.735 ;
        RECT 113.635 108.015 113.965 108.395 ;
        RECT 114.135 108.275 114.390 108.565 ;
        RECT 114.570 108.725 114.780 109.375 ;
        RECT 115.520 109.255 115.690 109.845 ;
        RECT 116.910 109.675 117.080 110.055 ;
        RECT 118.015 109.935 118.185 110.395 ;
        RECT 118.355 110.105 118.725 110.565 ;
        RECT 119.020 109.965 119.190 110.305 ;
        RECT 119.360 110.135 119.690 110.565 ;
        RECT 119.925 109.965 120.095 110.305 ;
        RECT 115.860 109.505 117.080 109.675 ;
        RECT 117.250 109.595 117.710 109.885 ;
        RECT 118.015 109.765 118.575 109.935 ;
        RECT 119.020 109.795 120.095 109.965 ;
        RECT 120.265 110.065 120.945 110.395 ;
        RECT 121.160 110.065 121.410 110.395 ;
        RECT 121.580 110.105 121.830 110.565 ;
        RECT 118.405 109.625 118.575 109.765 ;
        RECT 117.250 109.585 118.215 109.595 ;
        RECT 116.910 109.415 117.080 109.505 ;
        RECT 117.540 109.425 118.215 109.585 ;
        RECT 114.950 109.225 115.690 109.255 ;
        RECT 114.950 108.925 115.865 109.225 ;
        RECT 115.540 108.750 115.865 108.925 ;
        RECT 114.570 108.195 114.825 108.725 ;
        RECT 114.995 108.015 115.300 108.475 ;
        RECT 115.545 108.395 115.865 108.750 ;
        RECT 116.035 108.965 116.575 109.335 ;
        RECT 116.910 109.245 117.315 109.415 ;
        RECT 116.035 108.565 116.275 108.965 ;
        RECT 116.755 108.795 116.975 109.075 ;
        RECT 116.445 108.625 116.975 108.795 ;
        RECT 116.445 108.395 116.615 108.625 ;
        RECT 117.145 108.465 117.315 109.245 ;
        RECT 117.485 108.635 117.835 109.255 ;
        RECT 118.005 108.635 118.215 109.425 ;
        RECT 118.405 109.455 119.905 109.625 ;
        RECT 118.405 108.765 118.575 109.455 ;
        RECT 120.265 109.285 120.435 110.065 ;
        RECT 121.240 109.935 121.410 110.065 ;
        RECT 118.745 109.115 120.435 109.285 ;
        RECT 120.605 109.505 121.070 109.895 ;
        RECT 121.240 109.765 121.635 109.935 ;
        RECT 118.745 108.935 118.915 109.115 ;
        RECT 115.545 108.225 116.615 108.395 ;
        RECT 116.785 108.015 116.975 108.455 ;
        RECT 117.145 108.185 118.095 108.465 ;
        RECT 118.405 108.375 118.665 108.765 ;
        RECT 119.085 108.695 119.875 108.945 ;
        RECT 118.315 108.205 118.665 108.375 ;
        RECT 118.875 108.015 119.205 108.475 ;
        RECT 120.080 108.405 120.250 109.115 ;
        RECT 120.605 108.915 120.775 109.505 ;
        RECT 120.420 108.695 120.775 108.915 ;
        RECT 120.945 108.695 121.295 109.315 ;
        RECT 121.465 108.405 121.635 109.765 ;
        RECT 122.000 109.595 122.325 110.380 ;
        RECT 121.805 108.545 122.265 109.595 ;
        RECT 120.080 108.235 120.935 108.405 ;
        RECT 121.140 108.235 121.635 108.405 ;
        RECT 121.805 108.015 122.135 108.375 ;
        RECT 122.495 108.275 122.665 110.395 ;
        RECT 122.835 110.065 123.165 110.565 ;
        RECT 123.335 109.895 123.590 110.395 ;
        RECT 122.840 109.725 123.590 109.895 ;
        RECT 122.840 108.735 123.070 109.725 ;
        RECT 123.240 108.905 123.590 109.555 ;
        RECT 123.765 109.475 124.975 110.565 ;
        RECT 125.145 109.490 125.415 110.395 ;
        RECT 125.585 109.805 125.915 110.565 ;
        RECT 126.095 109.635 126.275 110.395 ;
        RECT 123.765 108.935 124.285 109.475 ;
        RECT 124.455 108.765 124.975 109.305 ;
        RECT 122.840 108.565 123.590 108.735 ;
        RECT 122.835 108.015 123.165 108.395 ;
        RECT 123.335 108.275 123.590 108.565 ;
        RECT 123.765 108.015 124.975 108.765 ;
        RECT 125.145 108.690 125.325 109.490 ;
        RECT 125.600 109.465 126.275 109.635 ;
        RECT 126.525 109.475 127.735 110.565 ;
        RECT 125.600 109.320 125.770 109.465 ;
        RECT 125.495 108.990 125.770 109.320 ;
        RECT 125.600 108.735 125.770 108.990 ;
        RECT 125.995 108.915 126.335 109.285 ;
        RECT 126.525 108.935 127.045 109.475 ;
        RECT 127.215 108.765 127.735 109.305 ;
        RECT 125.145 108.185 125.405 108.690 ;
        RECT 125.600 108.565 126.265 108.735 ;
        RECT 125.585 108.015 125.915 108.395 ;
        RECT 126.095 108.185 126.265 108.565 ;
        RECT 126.525 108.015 127.735 108.765 ;
        RECT 20.640 107.845 127.820 108.015 ;
        RECT 20.725 107.095 21.935 107.845 ;
        RECT 20.725 106.555 21.245 107.095 ;
        RECT 22.565 107.075 24.235 107.845 ;
        RECT 24.405 107.120 24.695 107.845 ;
        RECT 24.870 107.135 25.125 107.665 ;
        RECT 25.295 107.385 25.600 107.845 ;
        RECT 25.845 107.465 26.915 107.635 ;
        RECT 21.415 106.385 21.935 106.925 ;
        RECT 20.725 105.295 21.935 106.385 ;
        RECT 22.565 106.385 23.315 106.905 ;
        RECT 23.485 106.555 24.235 107.075 ;
        RECT 24.870 106.485 25.080 107.135 ;
        RECT 25.845 107.110 26.165 107.465 ;
        RECT 25.840 106.935 26.165 107.110 ;
        RECT 25.250 106.635 26.165 106.935 ;
        RECT 26.335 106.895 26.575 107.295 ;
        RECT 26.745 107.235 26.915 107.465 ;
        RECT 27.085 107.405 27.275 107.845 ;
        RECT 27.445 107.395 28.395 107.675 ;
        RECT 28.615 107.485 28.965 107.655 ;
        RECT 26.745 107.065 27.275 107.235 ;
        RECT 25.250 106.605 25.990 106.635 ;
        RECT 22.565 105.295 24.235 106.385 ;
        RECT 24.405 105.295 24.695 106.460 ;
        RECT 24.870 105.605 25.125 106.485 ;
        RECT 25.295 105.295 25.600 106.435 ;
        RECT 25.820 106.015 25.990 106.605 ;
        RECT 26.335 106.525 26.875 106.895 ;
        RECT 27.055 106.785 27.275 107.065 ;
        RECT 27.445 106.615 27.615 107.395 ;
        RECT 27.210 106.445 27.615 106.615 ;
        RECT 27.785 106.605 28.135 107.225 ;
        RECT 27.210 106.355 27.380 106.445 ;
        RECT 28.305 106.435 28.515 107.225 ;
        RECT 26.160 106.185 27.380 106.355 ;
        RECT 27.840 106.275 28.515 106.435 ;
        RECT 25.820 105.845 26.620 106.015 ;
        RECT 25.940 105.295 26.270 105.675 ;
        RECT 26.450 105.555 26.620 105.845 ;
        RECT 27.210 105.805 27.380 106.185 ;
        RECT 27.550 106.265 28.515 106.275 ;
        RECT 28.705 107.095 28.965 107.485 ;
        RECT 29.175 107.385 29.505 107.845 ;
        RECT 30.380 107.455 31.235 107.625 ;
        RECT 31.440 107.455 31.935 107.625 ;
        RECT 32.105 107.485 32.435 107.845 ;
        RECT 28.705 106.405 28.875 107.095 ;
        RECT 29.045 106.745 29.215 106.925 ;
        RECT 29.385 106.915 30.175 107.165 ;
        RECT 30.380 106.745 30.550 107.455 ;
        RECT 30.720 106.945 31.075 107.165 ;
        RECT 29.045 106.575 30.735 106.745 ;
        RECT 27.550 105.975 28.010 106.265 ;
        RECT 28.705 106.235 30.205 106.405 ;
        RECT 28.705 106.095 28.875 106.235 ;
        RECT 28.315 105.925 28.875 106.095 ;
        RECT 26.790 105.295 27.040 105.755 ;
        RECT 27.210 105.465 28.080 105.805 ;
        RECT 28.315 105.465 28.485 105.925 ;
        RECT 29.320 105.895 30.395 106.065 ;
        RECT 28.655 105.295 29.025 105.755 ;
        RECT 29.320 105.555 29.490 105.895 ;
        RECT 29.660 105.295 29.990 105.725 ;
        RECT 30.225 105.555 30.395 105.895 ;
        RECT 30.565 105.795 30.735 106.575 ;
        RECT 30.905 106.355 31.075 106.945 ;
        RECT 31.245 106.545 31.595 107.165 ;
        RECT 30.905 105.965 31.370 106.355 ;
        RECT 31.765 106.095 31.935 107.455 ;
        RECT 32.105 106.265 32.565 107.315 ;
        RECT 31.540 105.925 31.935 106.095 ;
        RECT 31.540 105.795 31.710 105.925 ;
        RECT 30.565 105.465 31.245 105.795 ;
        RECT 31.460 105.465 31.710 105.795 ;
        RECT 31.880 105.295 32.130 105.755 ;
        RECT 32.300 105.480 32.625 106.265 ;
        RECT 32.795 105.465 32.965 107.585 ;
        RECT 33.135 107.465 33.465 107.845 ;
        RECT 33.635 107.295 33.890 107.585 ;
        RECT 33.140 107.125 33.890 107.295 ;
        RECT 33.140 106.135 33.370 107.125 ;
        RECT 34.525 107.075 37.115 107.845 ;
        RECT 37.285 107.120 37.575 107.845 ;
        RECT 37.745 107.095 38.955 107.845 ;
        RECT 39.130 107.300 44.475 107.845 ;
        RECT 44.650 107.300 49.995 107.845 ;
        RECT 33.540 106.305 33.890 106.955 ;
        RECT 34.525 106.385 35.735 106.905 ;
        RECT 35.905 106.555 37.115 107.075 ;
        RECT 33.140 105.965 33.890 106.135 ;
        RECT 33.135 105.295 33.465 105.795 ;
        RECT 33.635 105.465 33.890 105.965 ;
        RECT 34.525 105.295 37.115 106.385 ;
        RECT 37.285 105.295 37.575 106.460 ;
        RECT 37.745 106.385 38.265 106.925 ;
        RECT 38.435 106.555 38.955 107.095 ;
        RECT 37.745 105.295 38.955 106.385 ;
        RECT 40.720 105.730 41.070 106.980 ;
        RECT 42.550 106.470 42.890 107.300 ;
        RECT 46.240 105.730 46.590 106.980 ;
        RECT 48.070 106.470 48.410 107.300 ;
        RECT 50.165 107.120 50.455 107.845 ;
        RECT 50.625 107.095 51.835 107.845 ;
        RECT 52.010 107.300 57.355 107.845 ;
        RECT 57.530 107.300 62.875 107.845 ;
        RECT 39.130 105.295 44.475 105.730 ;
        RECT 44.650 105.295 49.995 105.730 ;
        RECT 50.165 105.295 50.455 106.460 ;
        RECT 50.625 106.385 51.145 106.925 ;
        RECT 51.315 106.555 51.835 107.095 ;
        RECT 50.625 105.295 51.835 106.385 ;
        RECT 53.600 105.730 53.950 106.980 ;
        RECT 55.430 106.470 55.770 107.300 ;
        RECT 59.120 105.730 59.470 106.980 ;
        RECT 60.950 106.470 61.290 107.300 ;
        RECT 63.045 107.120 63.335 107.845 ;
        RECT 63.505 107.075 65.175 107.845 ;
        RECT 52.010 105.295 57.355 105.730 ;
        RECT 57.530 105.295 62.875 105.730 ;
        RECT 63.045 105.295 63.335 106.460 ;
        RECT 63.505 106.385 64.255 106.905 ;
        RECT 64.425 106.555 65.175 107.075 ;
        RECT 65.385 107.025 65.615 107.845 ;
        RECT 65.785 107.045 66.115 107.675 ;
        RECT 65.365 106.605 65.695 106.855 ;
        RECT 65.865 106.445 66.115 107.045 ;
        RECT 66.285 107.025 66.495 107.845 ;
        RECT 67.225 107.025 67.455 107.845 ;
        RECT 67.625 107.045 67.955 107.675 ;
        RECT 67.205 106.605 67.535 106.855 ;
        RECT 67.705 106.445 67.955 107.045 ;
        RECT 68.125 107.025 68.335 107.845 ;
        RECT 68.565 107.075 70.235 107.845 ;
        RECT 70.410 107.300 75.755 107.845 ;
        RECT 63.505 105.295 65.175 106.385 ;
        RECT 65.385 105.295 65.615 106.435 ;
        RECT 65.785 105.465 66.115 106.445 ;
        RECT 66.285 105.295 66.495 106.435 ;
        RECT 67.225 105.295 67.455 106.435 ;
        RECT 67.625 105.465 67.955 106.445 ;
        RECT 68.125 105.295 68.335 106.435 ;
        RECT 68.565 106.385 69.315 106.905 ;
        RECT 69.485 106.555 70.235 107.075 ;
        RECT 68.565 105.295 70.235 106.385 ;
        RECT 72.000 105.730 72.350 106.980 ;
        RECT 73.830 106.470 74.170 107.300 ;
        RECT 75.925 107.120 76.215 107.845 ;
        RECT 76.385 107.095 77.595 107.845 ;
        RECT 77.770 107.300 83.115 107.845 ;
        RECT 83.290 107.300 88.635 107.845 ;
        RECT 70.410 105.295 75.755 105.730 ;
        RECT 75.925 105.295 76.215 106.460 ;
        RECT 76.385 106.385 76.905 106.925 ;
        RECT 77.075 106.555 77.595 107.095 ;
        RECT 76.385 105.295 77.595 106.385 ;
        RECT 79.360 105.730 79.710 106.980 ;
        RECT 81.190 106.470 81.530 107.300 ;
        RECT 84.880 105.730 85.230 106.980 ;
        RECT 86.710 106.470 87.050 107.300 ;
        RECT 88.805 107.120 89.095 107.845 ;
        RECT 89.725 107.075 92.315 107.845 ;
        RECT 92.490 107.295 92.745 107.585 ;
        RECT 92.915 107.465 93.245 107.845 ;
        RECT 92.490 107.125 93.240 107.295 ;
        RECT 77.770 105.295 83.115 105.730 ;
        RECT 83.290 105.295 88.635 105.730 ;
        RECT 88.805 105.295 89.095 106.460 ;
        RECT 89.725 106.385 90.935 106.905 ;
        RECT 91.105 106.555 92.315 107.075 ;
        RECT 89.725 105.295 92.315 106.385 ;
        RECT 92.490 106.305 92.840 106.955 ;
        RECT 93.010 106.135 93.240 107.125 ;
        RECT 92.490 105.965 93.240 106.135 ;
        RECT 92.490 105.465 92.745 105.965 ;
        RECT 92.915 105.295 93.245 105.795 ;
        RECT 93.415 105.465 93.585 107.585 ;
        RECT 93.945 107.485 94.275 107.845 ;
        RECT 94.445 107.455 94.940 107.625 ;
        RECT 95.145 107.455 96.000 107.625 ;
        RECT 93.815 106.265 94.275 107.315 ;
        RECT 93.755 105.480 94.080 106.265 ;
        RECT 94.445 106.095 94.615 107.455 ;
        RECT 94.785 106.545 95.135 107.165 ;
        RECT 95.305 106.945 95.660 107.165 ;
        RECT 95.305 106.355 95.475 106.945 ;
        RECT 95.830 106.745 96.000 107.455 ;
        RECT 96.875 107.385 97.205 107.845 ;
        RECT 97.415 107.485 97.765 107.655 ;
        RECT 96.205 106.915 96.995 107.165 ;
        RECT 97.415 107.095 97.675 107.485 ;
        RECT 97.985 107.395 98.935 107.675 ;
        RECT 99.105 107.405 99.295 107.845 ;
        RECT 99.465 107.465 100.535 107.635 ;
        RECT 97.165 106.745 97.335 106.925 ;
        RECT 94.445 105.925 94.840 106.095 ;
        RECT 95.010 105.965 95.475 106.355 ;
        RECT 95.645 106.575 97.335 106.745 ;
        RECT 94.670 105.795 94.840 105.925 ;
        RECT 95.645 105.795 95.815 106.575 ;
        RECT 97.505 106.405 97.675 107.095 ;
        RECT 96.175 106.235 97.675 106.405 ;
        RECT 97.865 106.435 98.075 107.225 ;
        RECT 98.245 106.605 98.595 107.225 ;
        RECT 98.765 106.615 98.935 107.395 ;
        RECT 99.465 107.235 99.635 107.465 ;
        RECT 99.105 107.065 99.635 107.235 ;
        RECT 99.105 106.785 99.325 107.065 ;
        RECT 99.805 106.895 100.045 107.295 ;
        RECT 98.765 106.445 99.170 106.615 ;
        RECT 99.505 106.525 100.045 106.895 ;
        RECT 100.215 107.110 100.535 107.465 ;
        RECT 100.780 107.385 101.085 107.845 ;
        RECT 101.255 107.135 101.510 107.665 ;
        RECT 100.215 106.935 100.540 107.110 ;
        RECT 100.215 106.635 101.130 106.935 ;
        RECT 100.390 106.605 101.130 106.635 ;
        RECT 97.865 106.275 98.540 106.435 ;
        RECT 99.000 106.355 99.170 106.445 ;
        RECT 97.865 106.265 98.830 106.275 ;
        RECT 97.505 106.095 97.675 106.235 ;
        RECT 94.250 105.295 94.500 105.755 ;
        RECT 94.670 105.465 94.920 105.795 ;
        RECT 95.135 105.465 95.815 105.795 ;
        RECT 95.985 105.895 97.060 106.065 ;
        RECT 97.505 105.925 98.065 106.095 ;
        RECT 98.370 105.975 98.830 106.265 ;
        RECT 99.000 106.185 100.220 106.355 ;
        RECT 95.985 105.555 96.155 105.895 ;
        RECT 96.390 105.295 96.720 105.725 ;
        RECT 96.890 105.555 97.060 105.895 ;
        RECT 97.355 105.295 97.725 105.755 ;
        RECT 97.895 105.465 98.065 105.925 ;
        RECT 99.000 105.805 99.170 106.185 ;
        RECT 100.390 106.015 100.560 106.605 ;
        RECT 101.300 106.485 101.510 107.135 ;
        RECT 101.685 107.120 101.975 107.845 ;
        RECT 102.145 107.095 103.355 107.845 ;
        RECT 103.530 107.300 108.875 107.845 ;
        RECT 109.050 107.300 114.395 107.845 ;
        RECT 98.300 105.465 99.170 105.805 ;
        RECT 99.760 105.845 100.560 106.015 ;
        RECT 99.340 105.295 99.590 105.755 ;
        RECT 99.760 105.555 99.930 105.845 ;
        RECT 100.110 105.295 100.440 105.675 ;
        RECT 100.780 105.295 101.085 106.435 ;
        RECT 101.255 105.605 101.510 106.485 ;
        RECT 101.685 105.295 101.975 106.460 ;
        RECT 102.145 106.385 102.665 106.925 ;
        RECT 102.835 106.555 103.355 107.095 ;
        RECT 102.145 105.295 103.355 106.385 ;
        RECT 105.120 105.730 105.470 106.980 ;
        RECT 106.950 106.470 107.290 107.300 ;
        RECT 110.640 105.730 110.990 106.980 ;
        RECT 112.470 106.470 112.810 107.300 ;
        RECT 114.565 107.120 114.855 107.845 ;
        RECT 115.490 107.300 120.835 107.845 ;
        RECT 121.010 107.300 126.355 107.845 ;
        RECT 103.530 105.295 108.875 105.730 ;
        RECT 109.050 105.295 114.395 105.730 ;
        RECT 114.565 105.295 114.855 106.460 ;
        RECT 117.080 105.730 117.430 106.980 ;
        RECT 118.910 106.470 119.250 107.300 ;
        RECT 122.600 105.730 122.950 106.980 ;
        RECT 124.430 106.470 124.770 107.300 ;
        RECT 126.525 107.095 127.735 107.845 ;
        RECT 126.525 106.385 127.045 106.925 ;
        RECT 127.215 106.555 127.735 107.095 ;
        RECT 115.490 105.295 120.835 105.730 ;
        RECT 121.010 105.295 126.355 105.730 ;
        RECT 126.525 105.295 127.735 106.385 ;
        RECT 20.640 105.125 127.820 105.295 ;
        RECT 19.165 66.070 30.165 66.940 ;
        RECT 19.165 54.930 20.835 66.070 ;
        RECT 21.465 65.555 26.465 65.725 ;
        RECT 21.235 55.300 21.405 65.340 ;
        RECT 26.525 55.300 26.695 65.340 ;
        RECT 27.095 54.930 27.265 66.070 ;
        RECT 27.895 65.555 28.895 65.725 ;
        RECT 27.665 55.300 27.835 65.340 ;
        RECT 28.955 55.300 29.125 65.340 ;
        RECT 29.525 54.930 30.165 66.070 ;
        RECT 19.165 52.860 30.165 54.930 ;
        RECT 19.165 49.370 21.005 52.860 ;
        RECT 22.765 52.780 30.165 52.860 ;
        RECT 21.635 52.350 22.135 52.520 ;
        RECT 21.405 50.095 21.575 52.135 ;
        RECT 22.195 50.095 22.365 52.135 ;
        RECT 21.635 49.710 22.135 49.880 ;
        RECT 22.765 49.370 25.085 52.780 ;
        RECT 25.715 52.270 26.215 52.440 ;
        RECT 19.165 48.650 25.085 49.370 ;
        RECT 19.135 48.040 23.045 48.260 ;
        RECT 19.135 45.640 20.855 48.040 ;
        RECT 21.485 47.530 21.985 47.700 ;
        RECT 21.255 46.320 21.425 47.360 ;
        RECT 22.045 46.320 22.215 47.360 ;
        RECT 21.485 45.980 21.985 46.150 ;
        RECT 22.615 45.640 23.045 48.040 ;
        RECT 24.025 46.290 25.085 48.650 ;
        RECT 25.485 47.015 25.655 52.055 ;
        RECT 26.275 47.015 26.445 52.055 ;
        RECT 25.715 46.630 26.215 46.800 ;
        RECT 26.845 46.290 27.015 52.780 ;
        RECT 27.645 52.270 28.145 52.440 ;
        RECT 27.415 47.015 27.585 52.055 ;
        RECT 28.205 47.015 28.375 52.055 ;
        RECT 27.645 46.630 28.145 46.800 ;
        RECT 28.775 46.290 30.165 52.780 ;
        RECT 30.365 66.080 41.365 66.950 ;
        RECT 30.365 54.940 32.035 66.080 ;
        RECT 32.665 65.565 37.665 65.735 ;
        RECT 32.435 55.310 32.605 65.350 ;
        RECT 37.725 55.310 37.895 65.350 ;
        RECT 38.295 54.940 38.465 66.080 ;
        RECT 39.095 65.565 40.095 65.735 ;
        RECT 38.865 55.310 39.035 65.350 ;
        RECT 40.155 55.310 40.325 65.350 ;
        RECT 40.725 54.940 41.365 66.080 ;
        RECT 30.365 52.870 41.365 54.940 ;
        RECT 30.365 49.380 32.205 52.870 ;
        RECT 33.965 52.790 41.365 52.870 ;
        RECT 32.835 52.360 33.335 52.530 ;
        RECT 32.605 50.105 32.775 52.145 ;
        RECT 33.395 50.105 33.565 52.145 ;
        RECT 32.835 49.720 33.335 49.890 ;
        RECT 33.965 49.380 36.285 52.790 ;
        RECT 36.915 52.280 37.415 52.450 ;
        RECT 30.365 48.660 36.285 49.380 ;
        RECT 24.025 45.800 30.165 46.290 ;
        RECT 30.335 48.050 34.245 48.270 ;
        RECT 19.135 45.370 23.045 45.640 ;
        RECT 30.335 45.650 32.055 48.050 ;
        RECT 32.685 47.540 33.185 47.710 ;
        RECT 32.455 46.330 32.625 47.370 ;
        RECT 33.245 46.330 33.415 47.370 ;
        RECT 32.685 45.990 33.185 46.160 ;
        RECT 33.815 45.650 34.245 48.050 ;
        RECT 35.225 46.300 36.285 48.660 ;
        RECT 36.685 47.025 36.855 52.065 ;
        RECT 37.475 47.025 37.645 52.065 ;
        RECT 36.915 46.640 37.415 46.810 ;
        RECT 38.045 46.300 38.215 52.790 ;
        RECT 38.845 52.280 39.345 52.450 ;
        RECT 38.615 47.025 38.785 52.065 ;
        RECT 39.405 47.025 39.575 52.065 ;
        RECT 38.845 46.640 39.345 46.810 ;
        RECT 39.975 46.300 41.365 52.790 ;
        RECT 41.585 66.050 52.585 66.920 ;
        RECT 41.585 54.910 43.255 66.050 ;
        RECT 43.885 65.535 48.885 65.705 ;
        RECT 43.655 55.280 43.825 65.320 ;
        RECT 48.945 55.280 49.115 65.320 ;
        RECT 49.515 54.910 49.685 66.050 ;
        RECT 50.315 65.535 51.315 65.705 ;
        RECT 50.085 55.280 50.255 65.320 ;
        RECT 51.375 55.280 51.545 65.320 ;
        RECT 51.945 54.910 52.585 66.050 ;
        RECT 41.585 52.840 52.585 54.910 ;
        RECT 41.585 49.350 43.425 52.840 ;
        RECT 45.185 52.760 52.585 52.840 ;
        RECT 44.055 52.330 44.555 52.500 ;
        RECT 43.825 50.075 43.995 52.115 ;
        RECT 44.615 50.075 44.785 52.115 ;
        RECT 44.055 49.690 44.555 49.860 ;
        RECT 45.185 49.350 47.505 52.760 ;
        RECT 48.135 52.250 48.635 52.420 ;
        RECT 41.585 48.630 47.505 49.350 ;
        RECT 35.225 45.810 41.365 46.300 ;
        RECT 41.555 48.020 45.465 48.240 ;
        RECT 30.335 45.380 34.245 45.650 ;
        RECT 41.555 45.620 43.275 48.020 ;
        RECT 43.905 47.510 44.405 47.680 ;
        RECT 43.675 46.300 43.845 47.340 ;
        RECT 44.465 46.300 44.635 47.340 ;
        RECT 43.905 45.960 44.405 46.130 ;
        RECT 45.035 45.620 45.465 48.020 ;
        RECT 46.445 46.270 47.505 48.630 ;
        RECT 47.905 46.995 48.075 52.035 ;
        RECT 48.695 46.995 48.865 52.035 ;
        RECT 48.135 46.610 48.635 46.780 ;
        RECT 49.265 46.270 49.435 52.760 ;
        RECT 50.065 52.250 50.565 52.420 ;
        RECT 49.835 46.995 50.005 52.035 ;
        RECT 50.625 46.995 50.795 52.035 ;
        RECT 50.065 46.610 50.565 46.780 ;
        RECT 51.195 46.270 52.585 52.760 ;
        RECT 52.835 66.030 63.835 66.900 ;
        RECT 52.835 54.890 54.505 66.030 ;
        RECT 55.135 65.515 60.135 65.685 ;
        RECT 54.905 55.260 55.075 65.300 ;
        RECT 60.195 55.260 60.365 65.300 ;
        RECT 60.765 54.890 60.935 66.030 ;
        RECT 61.565 65.515 62.565 65.685 ;
        RECT 61.335 55.260 61.505 65.300 ;
        RECT 62.625 55.260 62.795 65.300 ;
        RECT 63.195 54.890 63.835 66.030 ;
        RECT 52.835 52.820 63.835 54.890 ;
        RECT 52.835 49.330 54.675 52.820 ;
        RECT 56.435 52.740 63.835 52.820 ;
        RECT 55.305 52.310 55.805 52.480 ;
        RECT 55.075 50.055 55.245 52.095 ;
        RECT 55.865 50.055 56.035 52.095 ;
        RECT 55.305 49.670 55.805 49.840 ;
        RECT 56.435 49.330 58.755 52.740 ;
        RECT 59.385 52.230 59.885 52.400 ;
        RECT 52.835 48.610 58.755 49.330 ;
        RECT 46.445 45.780 52.585 46.270 ;
        RECT 52.805 48.000 56.715 48.220 ;
        RECT 41.555 45.350 45.465 45.620 ;
        RECT 52.805 45.600 54.525 48.000 ;
        RECT 55.155 47.490 55.655 47.660 ;
        RECT 54.925 46.280 55.095 47.320 ;
        RECT 55.715 46.280 55.885 47.320 ;
        RECT 55.155 45.940 55.655 46.110 ;
        RECT 56.285 45.600 56.715 48.000 ;
        RECT 57.695 46.250 58.755 48.610 ;
        RECT 59.155 46.975 59.325 52.015 ;
        RECT 59.945 46.975 60.115 52.015 ;
        RECT 59.385 46.590 59.885 46.760 ;
        RECT 60.515 46.250 60.685 52.740 ;
        RECT 61.315 52.230 61.815 52.400 ;
        RECT 61.085 46.975 61.255 52.015 ;
        RECT 61.875 46.975 62.045 52.015 ;
        RECT 61.315 46.590 61.815 46.760 ;
        RECT 62.445 46.250 63.835 52.740 ;
        RECT 64.055 66.020 75.055 66.890 ;
        RECT 64.055 54.880 65.725 66.020 ;
        RECT 66.355 65.505 71.355 65.675 ;
        RECT 66.125 55.250 66.295 65.290 ;
        RECT 71.415 55.250 71.585 65.290 ;
        RECT 71.985 54.880 72.155 66.020 ;
        RECT 72.785 65.505 73.785 65.675 ;
        RECT 72.555 55.250 72.725 65.290 ;
        RECT 73.845 55.250 74.015 65.290 ;
        RECT 74.415 54.880 75.055 66.020 ;
        RECT 64.055 52.810 75.055 54.880 ;
        RECT 64.055 49.320 65.895 52.810 ;
        RECT 67.655 52.730 75.055 52.810 ;
        RECT 66.525 52.300 67.025 52.470 ;
        RECT 66.295 50.045 66.465 52.085 ;
        RECT 67.085 50.045 67.255 52.085 ;
        RECT 66.525 49.660 67.025 49.830 ;
        RECT 67.655 49.320 69.975 52.730 ;
        RECT 70.605 52.220 71.105 52.390 ;
        RECT 64.055 48.600 69.975 49.320 ;
        RECT 57.695 45.760 63.835 46.250 ;
        RECT 64.025 47.990 67.935 48.210 ;
        RECT 52.805 45.330 56.715 45.600 ;
        RECT 64.025 45.590 65.745 47.990 ;
        RECT 66.375 47.480 66.875 47.650 ;
        RECT 66.145 46.270 66.315 47.310 ;
        RECT 66.935 46.270 67.105 47.310 ;
        RECT 66.375 45.930 66.875 46.100 ;
        RECT 67.505 45.590 67.935 47.990 ;
        RECT 68.915 46.240 69.975 48.600 ;
        RECT 70.375 46.965 70.545 52.005 ;
        RECT 71.165 46.965 71.335 52.005 ;
        RECT 70.605 46.580 71.105 46.750 ;
        RECT 71.735 46.240 71.905 52.730 ;
        RECT 72.535 52.220 73.035 52.390 ;
        RECT 72.305 46.965 72.475 52.005 ;
        RECT 73.095 46.965 73.265 52.005 ;
        RECT 72.535 46.580 73.035 46.750 ;
        RECT 73.665 46.240 75.055 52.730 ;
        RECT 75.295 66.010 86.295 66.880 ;
        RECT 75.295 54.870 76.965 66.010 ;
        RECT 77.595 65.495 82.595 65.665 ;
        RECT 77.365 55.240 77.535 65.280 ;
        RECT 82.655 55.240 82.825 65.280 ;
        RECT 83.225 54.870 83.395 66.010 ;
        RECT 84.025 65.495 85.025 65.665 ;
        RECT 83.795 55.240 83.965 65.280 ;
        RECT 85.085 55.240 85.255 65.280 ;
        RECT 85.655 54.870 86.295 66.010 ;
        RECT 75.295 52.800 86.295 54.870 ;
        RECT 75.295 49.310 77.135 52.800 ;
        RECT 78.895 52.720 86.295 52.800 ;
        RECT 77.765 52.290 78.265 52.460 ;
        RECT 77.535 50.035 77.705 52.075 ;
        RECT 78.325 50.035 78.495 52.075 ;
        RECT 77.765 49.650 78.265 49.820 ;
        RECT 78.895 49.310 81.215 52.720 ;
        RECT 81.845 52.210 82.345 52.380 ;
        RECT 75.295 48.590 81.215 49.310 ;
        RECT 68.915 45.750 75.055 46.240 ;
        RECT 75.265 47.980 79.175 48.200 ;
        RECT 64.025 45.320 67.935 45.590 ;
        RECT 75.265 45.580 76.985 47.980 ;
        RECT 77.615 47.470 78.115 47.640 ;
        RECT 77.385 46.260 77.555 47.300 ;
        RECT 78.175 46.260 78.345 47.300 ;
        RECT 77.615 45.920 78.115 46.090 ;
        RECT 78.745 45.580 79.175 47.980 ;
        RECT 80.155 46.230 81.215 48.590 ;
        RECT 81.615 46.955 81.785 51.995 ;
        RECT 82.405 46.955 82.575 51.995 ;
        RECT 81.845 46.570 82.345 46.740 ;
        RECT 82.975 46.230 83.145 52.720 ;
        RECT 83.775 52.210 84.275 52.380 ;
        RECT 83.545 46.955 83.715 51.995 ;
        RECT 84.335 46.955 84.505 51.995 ;
        RECT 83.775 46.570 84.275 46.740 ;
        RECT 84.905 46.230 86.295 52.720 ;
        RECT 86.545 66.020 97.545 66.890 ;
        RECT 131.125 66.880 140.025 66.890 ;
        RECT 86.545 54.880 88.215 66.020 ;
        RECT 88.845 65.505 93.845 65.675 ;
        RECT 88.615 55.250 88.785 65.290 ;
        RECT 93.905 55.250 94.075 65.290 ;
        RECT 94.475 54.880 94.645 66.020 ;
        RECT 95.275 65.505 96.275 65.675 ;
        RECT 95.045 55.250 95.215 65.290 ;
        RECT 96.335 55.250 96.505 65.290 ;
        RECT 96.905 54.880 97.545 66.020 ;
        RECT 86.545 52.810 97.545 54.880 ;
        RECT 86.545 49.320 88.385 52.810 ;
        RECT 90.145 52.730 97.545 52.810 ;
        RECT 89.015 52.300 89.515 52.470 ;
        RECT 88.785 50.045 88.955 52.085 ;
        RECT 89.575 50.045 89.745 52.085 ;
        RECT 89.015 49.660 89.515 49.830 ;
        RECT 90.145 49.320 92.465 52.730 ;
        RECT 93.095 52.220 93.595 52.390 ;
        RECT 86.545 48.600 92.465 49.320 ;
        RECT 80.155 45.740 86.295 46.230 ;
        RECT 86.515 47.990 90.425 48.210 ;
        RECT 75.265 45.310 79.175 45.580 ;
        RECT 86.515 45.590 88.235 47.990 ;
        RECT 88.865 47.480 89.365 47.650 ;
        RECT 88.635 46.270 88.805 47.310 ;
        RECT 89.425 46.270 89.595 47.310 ;
        RECT 88.865 45.930 89.365 46.100 ;
        RECT 89.995 45.590 90.425 47.990 ;
        RECT 91.405 46.240 92.465 48.600 ;
        RECT 92.865 46.965 93.035 52.005 ;
        RECT 93.655 46.965 93.825 52.005 ;
        RECT 93.095 46.580 93.595 46.750 ;
        RECT 94.225 46.240 94.395 52.730 ;
        RECT 95.025 52.220 95.525 52.390 ;
        RECT 94.795 46.965 94.965 52.005 ;
        RECT 95.585 46.965 95.755 52.005 ;
        RECT 95.025 46.580 95.525 46.750 ;
        RECT 96.155 46.240 97.545 52.730 ;
        RECT 97.825 66.010 108.825 66.880 ;
        RECT 97.825 54.870 99.495 66.010 ;
        RECT 100.125 65.495 105.125 65.665 ;
        RECT 99.895 55.240 100.065 65.280 ;
        RECT 105.185 55.240 105.355 65.280 ;
        RECT 105.755 54.870 105.925 66.010 ;
        RECT 106.555 65.495 107.555 65.665 ;
        RECT 106.325 55.240 106.495 65.280 ;
        RECT 107.615 55.240 107.785 65.280 ;
        RECT 108.185 54.870 108.825 66.010 ;
        RECT 97.825 52.800 108.825 54.870 ;
        RECT 97.825 49.310 99.665 52.800 ;
        RECT 101.425 52.720 108.825 52.800 ;
        RECT 100.295 52.290 100.795 52.460 ;
        RECT 100.065 50.035 100.235 52.075 ;
        RECT 100.855 50.035 101.025 52.075 ;
        RECT 100.295 49.650 100.795 49.820 ;
        RECT 101.425 49.310 103.745 52.720 ;
        RECT 104.375 52.210 104.875 52.380 ;
        RECT 97.825 48.590 103.745 49.310 ;
        RECT 91.405 45.750 97.545 46.240 ;
        RECT 97.795 47.980 101.705 48.200 ;
        RECT 86.515 45.320 90.425 45.590 ;
        RECT 97.795 45.580 99.515 47.980 ;
        RECT 100.145 47.470 100.645 47.640 ;
        RECT 99.915 46.260 100.085 47.300 ;
        RECT 100.705 46.260 100.875 47.300 ;
        RECT 100.145 45.920 100.645 46.090 ;
        RECT 101.275 45.580 101.705 47.980 ;
        RECT 102.685 46.230 103.745 48.590 ;
        RECT 104.145 46.955 104.315 51.995 ;
        RECT 104.935 46.955 105.105 51.995 ;
        RECT 104.375 46.570 104.875 46.740 ;
        RECT 105.505 46.230 105.675 52.720 ;
        RECT 106.305 52.210 106.805 52.380 ;
        RECT 106.075 46.955 106.245 51.995 ;
        RECT 106.865 46.955 107.035 51.995 ;
        RECT 106.305 46.570 106.805 46.740 ;
        RECT 107.435 46.230 108.825 52.720 ;
        RECT 109.095 66.010 120.095 66.880 ;
        RECT 109.095 54.870 110.765 66.010 ;
        RECT 111.395 65.495 116.395 65.665 ;
        RECT 111.165 55.240 111.335 65.280 ;
        RECT 116.455 55.240 116.625 65.280 ;
        RECT 117.025 54.870 117.195 66.010 ;
        RECT 117.825 65.495 118.825 65.665 ;
        RECT 117.595 55.240 117.765 65.280 ;
        RECT 118.885 55.240 119.055 65.280 ;
        RECT 119.455 54.870 120.095 66.010 ;
        RECT 109.095 52.800 120.095 54.870 ;
        RECT 109.095 49.310 110.935 52.800 ;
        RECT 112.695 52.720 120.095 52.800 ;
        RECT 111.565 52.290 112.065 52.460 ;
        RECT 111.335 50.035 111.505 52.075 ;
        RECT 112.125 50.035 112.295 52.075 ;
        RECT 111.565 49.650 112.065 49.820 ;
        RECT 112.695 49.310 115.015 52.720 ;
        RECT 115.645 52.210 116.145 52.380 ;
        RECT 109.095 48.590 115.015 49.310 ;
        RECT 102.685 45.740 108.825 46.230 ;
        RECT 109.065 47.980 112.975 48.200 ;
        RECT 97.795 45.310 101.705 45.580 ;
        RECT 109.065 45.580 110.785 47.980 ;
        RECT 111.415 47.470 111.915 47.640 ;
        RECT 111.185 46.260 111.355 47.300 ;
        RECT 111.975 46.260 112.145 47.300 ;
        RECT 111.415 45.920 111.915 46.090 ;
        RECT 112.545 45.580 112.975 47.980 ;
        RECT 113.955 46.230 115.015 48.590 ;
        RECT 115.415 46.955 115.585 51.995 ;
        RECT 116.205 46.955 116.375 51.995 ;
        RECT 115.645 46.570 116.145 46.740 ;
        RECT 116.775 46.230 116.945 52.720 ;
        RECT 117.575 52.210 118.075 52.380 ;
        RECT 117.345 46.955 117.515 51.995 ;
        RECT 118.135 46.955 118.305 51.995 ;
        RECT 117.575 46.570 118.075 46.740 ;
        RECT 118.705 46.230 120.095 52.720 ;
        RECT 120.345 66.010 140.025 66.880 ;
        RECT 120.345 54.870 122.015 66.010 ;
        RECT 122.645 65.495 127.645 65.665 ;
        RECT 122.415 55.240 122.585 65.280 ;
        RECT 127.705 55.240 127.875 65.280 ;
        RECT 128.275 54.870 128.445 66.010 ;
        RECT 130.705 65.980 140.025 66.010 ;
        RECT 129.075 65.495 130.075 65.665 ;
        RECT 128.845 55.240 129.015 65.280 ;
        RECT 130.135 55.240 130.305 65.280 ;
        RECT 130.705 54.870 132.765 65.980 ;
        RECT 133.395 65.465 138.395 65.635 ;
        RECT 133.165 55.210 133.335 65.250 ;
        RECT 138.455 55.210 138.625 65.250 ;
        RECT 120.345 54.840 132.765 54.870 ;
        RECT 139.025 54.840 140.025 65.980 ;
        RECT 120.345 54.720 140.025 54.840 ;
        RECT 120.345 53.550 140.035 54.720 ;
        RECT 120.345 52.800 131.345 53.550 ;
        RECT 120.345 49.310 122.185 52.800 ;
        RECT 123.945 52.720 131.345 52.800 ;
        RECT 122.815 52.290 123.315 52.460 ;
        RECT 122.585 50.035 122.755 52.075 ;
        RECT 123.375 50.035 123.545 52.075 ;
        RECT 122.815 49.650 123.315 49.820 ;
        RECT 123.945 49.310 126.265 52.720 ;
        RECT 126.895 52.210 127.395 52.380 ;
        RECT 120.345 48.590 126.265 49.310 ;
        RECT 113.955 45.740 120.095 46.230 ;
        RECT 120.315 47.980 124.225 48.200 ;
        RECT 109.065 45.310 112.975 45.580 ;
        RECT 120.315 45.580 122.035 47.980 ;
        RECT 122.665 47.470 123.165 47.640 ;
        RECT 122.435 46.260 122.605 47.300 ;
        RECT 123.225 46.260 123.395 47.300 ;
        RECT 122.665 45.920 123.165 46.090 ;
        RECT 123.795 45.580 124.225 47.980 ;
        RECT 125.205 46.230 126.265 48.590 ;
        RECT 126.665 46.955 126.835 51.995 ;
        RECT 127.455 46.955 127.625 51.995 ;
        RECT 126.895 46.570 127.395 46.740 ;
        RECT 128.025 46.230 128.195 52.720 ;
        RECT 128.825 52.210 129.325 52.380 ;
        RECT 128.595 46.955 128.765 51.995 ;
        RECT 129.385 46.955 129.555 51.995 ;
        RECT 128.825 46.570 129.325 46.740 ;
        RECT 129.955 46.230 131.345 52.720 ;
        RECT 125.205 45.740 131.345 46.230 ;
        RECT 120.315 45.310 124.225 45.580 ;
        RECT 25.695 39.770 29.605 40.040 ;
        RECT 18.575 39.120 24.715 39.610 ;
        RECT 18.575 32.630 19.965 39.120 ;
        RECT 20.595 38.610 21.095 38.780 ;
        RECT 20.365 33.355 20.535 38.395 ;
        RECT 21.155 33.355 21.325 38.395 ;
        RECT 20.595 32.970 21.095 33.140 ;
        RECT 21.725 32.630 21.895 39.120 ;
        RECT 22.525 38.610 23.025 38.780 ;
        RECT 22.295 33.355 22.465 38.395 ;
        RECT 23.085 33.355 23.255 38.395 ;
        RECT 23.655 36.760 24.715 39.120 ;
        RECT 25.695 37.370 26.125 39.770 ;
        RECT 26.755 39.260 27.255 39.430 ;
        RECT 26.525 38.050 26.695 39.090 ;
        RECT 27.315 38.050 27.485 39.090 ;
        RECT 26.755 37.710 27.255 37.880 ;
        RECT 27.885 37.370 29.605 39.770 ;
        RECT 36.975 39.770 40.885 40.040 ;
        RECT 25.695 37.150 29.605 37.370 ;
        RECT 29.855 39.120 35.995 39.610 ;
        RECT 23.655 36.040 29.575 36.760 ;
        RECT 22.525 32.970 23.025 33.140 ;
        RECT 23.655 32.630 25.975 36.040 ;
        RECT 26.605 35.530 27.105 35.700 ;
        RECT 26.375 33.275 26.545 35.315 ;
        RECT 27.165 33.275 27.335 35.315 ;
        RECT 26.605 32.890 27.105 33.060 ;
        RECT 18.575 32.550 25.975 32.630 ;
        RECT 27.735 32.550 29.575 36.040 ;
        RECT 18.575 30.480 29.575 32.550 ;
        RECT 18.575 19.340 19.215 30.480 ;
        RECT 19.615 20.070 19.785 30.110 ;
        RECT 20.905 20.070 21.075 30.110 ;
        RECT 19.845 19.685 20.845 19.855 ;
        RECT 21.475 19.340 21.645 30.480 ;
        RECT 22.045 20.070 22.215 30.110 ;
        RECT 27.335 20.070 27.505 30.110 ;
        RECT 22.275 19.685 27.275 19.855 ;
        RECT 27.905 19.340 29.575 30.480 ;
        RECT 18.575 18.470 29.575 19.340 ;
        RECT 29.855 32.630 31.245 39.120 ;
        RECT 31.875 38.610 32.375 38.780 ;
        RECT 31.645 33.355 31.815 38.395 ;
        RECT 32.435 33.355 32.605 38.395 ;
        RECT 31.875 32.970 32.375 33.140 ;
        RECT 33.005 32.630 33.175 39.120 ;
        RECT 33.805 38.610 34.305 38.780 ;
        RECT 33.575 33.355 33.745 38.395 ;
        RECT 34.365 33.355 34.535 38.395 ;
        RECT 34.935 36.760 35.995 39.120 ;
        RECT 36.975 37.370 37.405 39.770 ;
        RECT 38.035 39.260 38.535 39.430 ;
        RECT 37.805 38.050 37.975 39.090 ;
        RECT 38.595 38.050 38.765 39.090 ;
        RECT 38.035 37.710 38.535 37.880 ;
        RECT 39.165 37.370 40.885 39.770 ;
        RECT 48.265 39.750 52.175 40.020 ;
        RECT 36.975 37.150 40.885 37.370 ;
        RECT 41.145 39.100 47.285 39.590 ;
        RECT 34.935 36.040 40.855 36.760 ;
        RECT 33.805 32.970 34.305 33.140 ;
        RECT 34.935 32.630 37.255 36.040 ;
        RECT 37.885 35.530 38.385 35.700 ;
        RECT 37.655 33.275 37.825 35.315 ;
        RECT 38.445 33.275 38.615 35.315 ;
        RECT 37.885 32.890 38.385 33.060 ;
        RECT 29.855 32.550 37.255 32.630 ;
        RECT 39.015 32.550 40.855 36.040 ;
        RECT 29.855 30.480 40.855 32.550 ;
        RECT 29.855 19.340 30.495 30.480 ;
        RECT 30.895 20.070 31.065 30.110 ;
        RECT 32.185 20.070 32.355 30.110 ;
        RECT 31.125 19.685 32.125 19.855 ;
        RECT 32.755 19.340 32.925 30.480 ;
        RECT 33.325 20.070 33.495 30.110 ;
        RECT 38.615 20.070 38.785 30.110 ;
        RECT 33.555 19.685 38.555 19.855 ;
        RECT 39.185 19.340 40.855 30.480 ;
        RECT 29.855 18.470 40.855 19.340 ;
        RECT 41.145 32.610 42.535 39.100 ;
        RECT 43.165 38.590 43.665 38.760 ;
        RECT 42.935 33.335 43.105 38.375 ;
        RECT 43.725 33.335 43.895 38.375 ;
        RECT 43.165 32.950 43.665 33.120 ;
        RECT 44.295 32.610 44.465 39.100 ;
        RECT 45.095 38.590 45.595 38.760 ;
        RECT 44.865 33.335 45.035 38.375 ;
        RECT 45.655 33.335 45.825 38.375 ;
        RECT 46.225 36.740 47.285 39.100 ;
        RECT 48.265 37.350 48.695 39.750 ;
        RECT 49.325 39.240 49.825 39.410 ;
        RECT 49.095 38.030 49.265 39.070 ;
        RECT 49.885 38.030 50.055 39.070 ;
        RECT 49.325 37.690 49.825 37.860 ;
        RECT 50.455 37.350 52.175 39.750 ;
        RECT 59.485 39.750 63.395 40.020 ;
        RECT 48.265 37.130 52.175 37.350 ;
        RECT 52.365 39.100 58.505 39.590 ;
        RECT 46.225 36.020 52.145 36.740 ;
        RECT 45.095 32.950 45.595 33.120 ;
        RECT 46.225 32.610 48.545 36.020 ;
        RECT 49.175 35.510 49.675 35.680 ;
        RECT 48.945 33.255 49.115 35.295 ;
        RECT 49.735 33.255 49.905 35.295 ;
        RECT 49.175 32.870 49.675 33.040 ;
        RECT 41.145 32.530 48.545 32.610 ;
        RECT 50.305 32.530 52.145 36.020 ;
        RECT 41.145 30.460 52.145 32.530 ;
        RECT 41.145 19.320 41.785 30.460 ;
        RECT 42.185 20.050 42.355 30.090 ;
        RECT 43.475 20.050 43.645 30.090 ;
        RECT 42.415 19.665 43.415 19.835 ;
        RECT 44.045 19.320 44.215 30.460 ;
        RECT 44.615 20.050 44.785 30.090 ;
        RECT 49.905 20.050 50.075 30.090 ;
        RECT 44.845 19.665 49.845 19.835 ;
        RECT 50.475 19.320 52.145 30.460 ;
        RECT 41.145 18.450 52.145 19.320 ;
        RECT 52.365 32.610 53.755 39.100 ;
        RECT 54.385 38.590 54.885 38.760 ;
        RECT 54.155 33.335 54.325 38.375 ;
        RECT 54.945 33.335 55.115 38.375 ;
        RECT 54.385 32.950 54.885 33.120 ;
        RECT 55.515 32.610 55.685 39.100 ;
        RECT 56.315 38.590 56.815 38.760 ;
        RECT 56.085 33.335 56.255 38.375 ;
        RECT 56.875 33.335 57.045 38.375 ;
        RECT 57.445 36.740 58.505 39.100 ;
        RECT 59.485 37.350 59.915 39.750 ;
        RECT 60.545 39.240 61.045 39.410 ;
        RECT 60.315 38.030 60.485 39.070 ;
        RECT 61.105 38.030 61.275 39.070 ;
        RECT 60.545 37.690 61.045 37.860 ;
        RECT 61.675 37.350 63.395 39.750 ;
        RECT 70.685 39.750 74.595 40.020 ;
        RECT 59.485 37.130 63.395 37.350 ;
        RECT 63.565 39.100 69.705 39.590 ;
        RECT 57.445 36.020 63.365 36.740 ;
        RECT 56.315 32.950 56.815 33.120 ;
        RECT 57.445 32.610 59.765 36.020 ;
        RECT 60.395 35.510 60.895 35.680 ;
        RECT 60.165 33.255 60.335 35.295 ;
        RECT 60.955 33.255 61.125 35.295 ;
        RECT 60.395 32.870 60.895 33.040 ;
        RECT 52.365 32.530 59.765 32.610 ;
        RECT 61.525 32.530 63.365 36.020 ;
        RECT 52.365 30.460 63.365 32.530 ;
        RECT 52.365 19.320 53.005 30.460 ;
        RECT 53.405 20.050 53.575 30.090 ;
        RECT 54.695 20.050 54.865 30.090 ;
        RECT 53.635 19.665 54.635 19.835 ;
        RECT 55.265 19.320 55.435 30.460 ;
        RECT 55.835 20.050 56.005 30.090 ;
        RECT 61.125 20.050 61.295 30.090 ;
        RECT 56.065 19.665 61.065 19.835 ;
        RECT 61.695 19.320 63.365 30.460 ;
        RECT 52.365 18.450 63.365 19.320 ;
        RECT 63.565 32.610 64.955 39.100 ;
        RECT 65.585 38.590 66.085 38.760 ;
        RECT 65.355 33.335 65.525 38.375 ;
        RECT 66.145 33.335 66.315 38.375 ;
        RECT 65.585 32.950 66.085 33.120 ;
        RECT 66.715 32.610 66.885 39.100 ;
        RECT 67.515 38.590 68.015 38.760 ;
        RECT 67.285 33.335 67.455 38.375 ;
        RECT 68.075 33.335 68.245 38.375 ;
        RECT 68.645 36.740 69.705 39.100 ;
        RECT 70.685 37.350 71.115 39.750 ;
        RECT 71.745 39.240 72.245 39.410 ;
        RECT 71.515 38.030 71.685 39.070 ;
        RECT 72.305 38.030 72.475 39.070 ;
        RECT 71.745 37.690 72.245 37.860 ;
        RECT 72.875 37.350 74.595 39.750 ;
        RECT 81.975 39.740 85.885 40.010 ;
        RECT 70.685 37.130 74.595 37.350 ;
        RECT 74.855 39.090 80.995 39.580 ;
        RECT 68.645 36.020 74.565 36.740 ;
        RECT 67.515 32.950 68.015 33.120 ;
        RECT 68.645 32.610 70.965 36.020 ;
        RECT 71.595 35.510 72.095 35.680 ;
        RECT 71.365 33.255 71.535 35.295 ;
        RECT 72.155 33.255 72.325 35.295 ;
        RECT 71.595 32.870 72.095 33.040 ;
        RECT 63.565 32.530 70.965 32.610 ;
        RECT 72.725 32.530 74.565 36.020 ;
        RECT 63.565 30.460 74.565 32.530 ;
        RECT 63.565 19.320 64.205 30.460 ;
        RECT 64.605 20.050 64.775 30.090 ;
        RECT 65.895 20.050 66.065 30.090 ;
        RECT 64.835 19.665 65.835 19.835 ;
        RECT 66.465 19.320 66.635 30.460 ;
        RECT 67.035 20.050 67.205 30.090 ;
        RECT 72.325 20.050 72.495 30.090 ;
        RECT 67.265 19.665 72.265 19.835 ;
        RECT 72.895 19.320 74.565 30.460 ;
        RECT 63.565 18.450 74.565 19.320 ;
        RECT 74.855 32.600 76.245 39.090 ;
        RECT 76.875 38.580 77.375 38.750 ;
        RECT 76.645 33.325 76.815 38.365 ;
        RECT 77.435 33.325 77.605 38.365 ;
        RECT 76.875 32.940 77.375 33.110 ;
        RECT 78.005 32.600 78.175 39.090 ;
        RECT 78.805 38.580 79.305 38.750 ;
        RECT 78.575 33.325 78.745 38.365 ;
        RECT 79.365 33.325 79.535 38.365 ;
        RECT 79.935 36.730 80.995 39.090 ;
        RECT 81.975 37.340 82.405 39.740 ;
        RECT 83.035 39.230 83.535 39.400 ;
        RECT 82.805 38.020 82.975 39.060 ;
        RECT 83.595 38.020 83.765 39.060 ;
        RECT 83.035 37.680 83.535 37.850 ;
        RECT 84.165 37.340 85.885 39.740 ;
        RECT 93.215 39.760 97.125 40.030 ;
        RECT 81.975 37.120 85.885 37.340 ;
        RECT 86.095 39.110 92.235 39.600 ;
        RECT 79.935 36.010 85.855 36.730 ;
        RECT 78.805 32.940 79.305 33.110 ;
        RECT 79.935 32.600 82.255 36.010 ;
        RECT 82.885 35.500 83.385 35.670 ;
        RECT 82.655 33.245 82.825 35.285 ;
        RECT 83.445 33.245 83.615 35.285 ;
        RECT 82.885 32.860 83.385 33.030 ;
        RECT 74.855 32.520 82.255 32.600 ;
        RECT 84.015 32.520 85.855 36.010 ;
        RECT 74.855 30.450 85.855 32.520 ;
        RECT 74.855 19.310 75.495 30.450 ;
        RECT 75.895 20.040 76.065 30.080 ;
        RECT 77.185 20.040 77.355 30.080 ;
        RECT 76.125 19.655 77.125 19.825 ;
        RECT 77.755 19.310 77.925 30.450 ;
        RECT 78.325 20.040 78.495 30.080 ;
        RECT 83.615 20.040 83.785 30.080 ;
        RECT 78.555 19.655 83.555 19.825 ;
        RECT 84.185 19.310 85.855 30.450 ;
        RECT 74.855 18.440 85.855 19.310 ;
        RECT 86.095 32.620 87.485 39.110 ;
        RECT 88.115 38.600 88.615 38.770 ;
        RECT 87.885 33.345 88.055 38.385 ;
        RECT 88.675 33.345 88.845 38.385 ;
        RECT 88.115 32.960 88.615 33.130 ;
        RECT 89.245 32.620 89.415 39.110 ;
        RECT 90.045 38.600 90.545 38.770 ;
        RECT 89.815 33.345 89.985 38.385 ;
        RECT 90.605 33.345 90.775 38.385 ;
        RECT 91.175 36.750 92.235 39.110 ;
        RECT 93.215 37.360 93.645 39.760 ;
        RECT 94.275 39.250 94.775 39.420 ;
        RECT 94.045 38.040 94.215 39.080 ;
        RECT 94.835 38.040 95.005 39.080 ;
        RECT 94.275 37.700 94.775 37.870 ;
        RECT 95.405 37.360 97.125 39.760 ;
        RECT 104.425 39.780 108.335 40.050 ;
        RECT 93.215 37.140 97.125 37.360 ;
        RECT 97.305 39.130 103.445 39.620 ;
        RECT 91.175 36.030 97.095 36.750 ;
        RECT 90.045 32.960 90.545 33.130 ;
        RECT 91.175 32.620 93.495 36.030 ;
        RECT 94.125 35.520 94.625 35.690 ;
        RECT 93.895 33.265 94.065 35.305 ;
        RECT 94.685 33.265 94.855 35.305 ;
        RECT 94.125 32.880 94.625 33.050 ;
        RECT 86.095 32.540 93.495 32.620 ;
        RECT 95.255 32.540 97.095 36.030 ;
        RECT 86.095 30.470 97.095 32.540 ;
        RECT 86.095 19.330 86.735 30.470 ;
        RECT 87.135 20.060 87.305 30.100 ;
        RECT 88.425 20.060 88.595 30.100 ;
        RECT 87.365 19.675 88.365 19.845 ;
        RECT 88.995 19.330 89.165 30.470 ;
        RECT 89.565 20.060 89.735 30.100 ;
        RECT 94.855 20.060 95.025 30.100 ;
        RECT 89.795 19.675 94.795 19.845 ;
        RECT 95.425 19.330 97.095 30.470 ;
        RECT 86.095 18.460 97.095 19.330 ;
        RECT 97.305 32.640 98.695 39.130 ;
        RECT 99.325 38.620 99.825 38.790 ;
        RECT 99.095 33.365 99.265 38.405 ;
        RECT 99.885 33.365 100.055 38.405 ;
        RECT 99.325 32.980 99.825 33.150 ;
        RECT 100.455 32.640 100.625 39.130 ;
        RECT 101.255 38.620 101.755 38.790 ;
        RECT 101.025 33.365 101.195 38.405 ;
        RECT 101.815 33.365 101.985 38.405 ;
        RECT 102.385 36.770 103.445 39.130 ;
        RECT 104.425 37.380 104.855 39.780 ;
        RECT 105.485 39.270 105.985 39.440 ;
        RECT 105.255 38.060 105.425 39.100 ;
        RECT 106.045 38.060 106.215 39.100 ;
        RECT 105.485 37.720 105.985 37.890 ;
        RECT 106.615 37.380 108.335 39.780 ;
        RECT 115.625 39.820 119.535 40.090 ;
        RECT 104.425 37.160 108.335 37.380 ;
        RECT 108.505 39.170 114.645 39.660 ;
        RECT 102.385 36.050 108.305 36.770 ;
        RECT 101.255 32.980 101.755 33.150 ;
        RECT 102.385 32.640 104.705 36.050 ;
        RECT 105.335 35.540 105.835 35.710 ;
        RECT 105.105 33.285 105.275 35.325 ;
        RECT 105.895 33.285 106.065 35.325 ;
        RECT 105.335 32.900 105.835 33.070 ;
        RECT 97.305 32.560 104.705 32.640 ;
        RECT 106.465 32.560 108.305 36.050 ;
        RECT 97.305 30.490 108.305 32.560 ;
        RECT 97.305 19.350 97.945 30.490 ;
        RECT 98.345 20.080 98.515 30.120 ;
        RECT 99.635 20.080 99.805 30.120 ;
        RECT 98.575 19.695 99.575 19.865 ;
        RECT 100.205 19.350 100.375 30.490 ;
        RECT 100.775 20.080 100.945 30.120 ;
        RECT 106.065 20.080 106.235 30.120 ;
        RECT 101.005 19.695 106.005 19.865 ;
        RECT 106.635 19.350 108.305 30.490 ;
        RECT 97.305 18.480 108.305 19.350 ;
        RECT 108.505 32.680 109.895 39.170 ;
        RECT 110.525 38.660 111.025 38.830 ;
        RECT 110.295 33.405 110.465 38.445 ;
        RECT 111.085 33.405 111.255 38.445 ;
        RECT 110.525 33.020 111.025 33.190 ;
        RECT 111.655 32.680 111.825 39.170 ;
        RECT 112.455 38.660 112.955 38.830 ;
        RECT 112.225 33.405 112.395 38.445 ;
        RECT 113.015 33.405 113.185 38.445 ;
        RECT 113.585 36.810 114.645 39.170 ;
        RECT 115.625 37.420 116.055 39.820 ;
        RECT 116.685 39.310 117.185 39.480 ;
        RECT 116.455 38.100 116.625 39.140 ;
        RECT 117.245 38.100 117.415 39.140 ;
        RECT 116.685 37.760 117.185 37.930 ;
        RECT 117.815 37.420 119.535 39.820 ;
        RECT 126.835 39.840 130.745 40.110 ;
        RECT 115.625 37.200 119.535 37.420 ;
        RECT 119.715 39.190 125.855 39.680 ;
        RECT 113.585 36.090 119.505 36.810 ;
        RECT 112.455 33.020 112.955 33.190 ;
        RECT 113.585 32.680 115.905 36.090 ;
        RECT 116.535 35.580 117.035 35.750 ;
        RECT 116.305 33.325 116.475 35.365 ;
        RECT 117.095 33.325 117.265 35.365 ;
        RECT 116.535 32.940 117.035 33.110 ;
        RECT 108.505 32.600 115.905 32.680 ;
        RECT 117.665 32.600 119.505 36.090 ;
        RECT 108.505 30.530 119.505 32.600 ;
        RECT 108.505 19.390 109.145 30.530 ;
        RECT 109.545 20.120 109.715 30.160 ;
        RECT 110.835 20.120 111.005 30.160 ;
        RECT 109.775 19.735 110.775 19.905 ;
        RECT 111.405 19.390 111.575 30.530 ;
        RECT 111.975 20.120 112.145 30.160 ;
        RECT 117.265 20.120 117.435 30.160 ;
        RECT 112.205 19.735 117.205 19.905 ;
        RECT 117.835 19.390 119.505 30.530 ;
        RECT 108.505 18.520 119.505 19.390 ;
        RECT 119.715 32.700 121.105 39.190 ;
        RECT 121.735 38.680 122.235 38.850 ;
        RECT 121.505 33.425 121.675 38.465 ;
        RECT 122.295 33.425 122.465 38.465 ;
        RECT 121.735 33.040 122.235 33.210 ;
        RECT 122.865 32.700 123.035 39.190 ;
        RECT 123.665 38.680 124.165 38.850 ;
        RECT 123.435 33.425 123.605 38.465 ;
        RECT 124.225 33.425 124.395 38.465 ;
        RECT 124.795 36.830 125.855 39.190 ;
        RECT 126.835 37.440 127.265 39.840 ;
        RECT 127.895 39.330 128.395 39.500 ;
        RECT 127.665 38.120 127.835 39.160 ;
        RECT 128.455 38.120 128.625 39.160 ;
        RECT 127.895 37.780 128.395 37.950 ;
        RECT 129.025 37.440 130.745 39.840 ;
        RECT 126.835 37.220 130.745 37.440 ;
        RECT 124.795 36.110 130.715 36.830 ;
        RECT 123.665 33.040 124.165 33.210 ;
        RECT 124.795 32.700 127.115 36.110 ;
        RECT 127.745 35.600 128.245 35.770 ;
        RECT 127.515 33.345 127.685 35.385 ;
        RECT 128.305 33.345 128.475 35.385 ;
        RECT 127.745 32.960 128.245 33.130 ;
        RECT 119.715 32.620 127.115 32.700 ;
        RECT 128.875 32.620 130.715 36.110 ;
        RECT 119.715 31.140 130.715 32.620 ;
        RECT 119.715 30.550 139.465 31.140 ;
        RECT 119.715 19.410 120.355 30.550 ;
        RECT 120.755 20.140 120.925 30.180 ;
        RECT 122.045 20.140 122.215 30.180 ;
        RECT 120.985 19.755 121.985 19.925 ;
        RECT 122.615 19.410 122.785 30.550 ;
        RECT 129.045 30.520 139.465 30.550 ;
        RECT 123.185 20.140 123.355 30.180 ;
        RECT 128.475 20.140 128.645 30.180 ;
        RECT 123.415 19.755 128.415 19.925 ;
        RECT 129.045 19.410 132.075 30.520 ;
        RECT 132.475 20.110 132.645 30.150 ;
        RECT 137.765 20.110 137.935 30.150 ;
        RECT 132.705 19.725 137.705 19.895 ;
        RECT 119.715 19.380 132.075 19.410 ;
        RECT 138.335 19.380 139.465 30.520 ;
        RECT 119.715 18.540 139.465 19.380 ;
        RECT 131.925 18.520 139.465 18.540 ;
      LAYER met1 ;
        RECT 135.340 223.880 136.790 225.180 ;
        RECT 20.640 211.050 127.820 211.530 ;
        RECT 20.640 208.330 127.820 208.810 ;
        RECT 20.640 205.610 127.820 206.090 ;
        RECT 20.640 202.890 127.820 203.370 ;
        RECT 72.690 201.810 73.010 202.070 ;
        RECT 72.230 201.470 72.550 201.730 ;
        RECT 64.870 200.990 65.190 201.050 ;
        RECT 70.405 200.990 70.695 201.035 ;
        RECT 64.870 200.850 70.695 200.990 ;
        RECT 64.870 200.790 65.190 200.850 ;
        RECT 70.405 200.805 70.695 200.850 ;
        RECT 20.640 200.170 127.820 200.650 ;
        RECT 62.125 199.970 62.415 200.015 ;
        RECT 62.125 199.830 66.940 199.970 ;
        RECT 62.125 199.785 62.415 199.830 ;
        RECT 49.685 199.630 50.335 199.675 ;
        RECT 52.450 199.630 52.770 199.690 ;
        RECT 53.285 199.630 53.575 199.675 ;
        RECT 49.685 199.490 53.575 199.630 ;
        RECT 49.685 199.445 50.335 199.490 ;
        RECT 52.450 199.430 52.770 199.490 ;
        RECT 52.985 199.445 53.575 199.490 ;
        RECT 46.490 199.290 46.780 199.335 ;
        RECT 48.325 199.290 48.615 199.335 ;
        RECT 51.905 199.290 52.195 199.335 ;
        RECT 46.490 199.150 52.195 199.290 ;
        RECT 46.490 199.105 46.780 199.150 ;
        RECT 48.325 199.105 48.615 199.150 ;
        RECT 51.905 199.105 52.195 199.150 ;
        RECT 52.985 199.130 53.275 199.445 ;
        RECT 64.870 199.430 65.190 199.690 ;
        RECT 66.800 199.630 66.940 199.830 ;
        RECT 67.165 199.630 67.815 199.675 ;
        RECT 70.765 199.630 71.055 199.675 ;
        RECT 66.800 199.490 71.055 199.630 ;
        RECT 67.165 199.445 67.815 199.490 ;
        RECT 70.465 199.445 71.055 199.490 ;
        RECT 71.310 199.630 71.630 199.690 ;
        RECT 77.750 199.630 78.070 199.690 ;
        RECT 99.945 199.630 100.235 199.675 ;
        RECT 100.750 199.630 101.070 199.690 ;
        RECT 103.185 199.630 103.835 199.675 ;
        RECT 71.310 199.490 78.900 199.630 ;
        RECT 62.585 199.105 62.875 199.335 ;
        RECT 63.970 199.290 64.260 199.335 ;
        RECT 65.805 199.290 66.095 199.335 ;
        RECT 69.385 199.290 69.675 199.335 ;
        RECT 63.970 199.150 69.675 199.290 ;
        RECT 63.970 199.105 64.260 199.150 ;
        RECT 65.805 199.105 66.095 199.150 ;
        RECT 69.385 199.105 69.675 199.150 ;
        RECT 70.465 199.130 70.755 199.445 ;
        RECT 71.310 199.430 71.630 199.490 ;
        RECT 77.750 199.430 78.070 199.490 ;
        RECT 46.010 198.750 46.330 199.010 ;
        RECT 47.405 198.950 47.695 198.995 ;
        RECT 49.230 198.950 49.550 199.010 ;
        RECT 47.405 198.810 49.550 198.950 ;
        RECT 47.405 198.765 47.695 198.810 ;
        RECT 49.230 198.750 49.550 198.810 ;
        RECT 46.895 198.610 47.185 198.655 ;
        RECT 48.785 198.610 49.075 198.655 ;
        RECT 51.905 198.610 52.195 198.655 ;
        RECT 46.895 198.470 52.195 198.610 ;
        RECT 46.895 198.425 47.185 198.470 ;
        RECT 48.785 198.425 49.075 198.470 ;
        RECT 51.905 198.425 52.195 198.470 ;
        RECT 54.750 198.070 55.070 198.330 ;
        RECT 62.660 198.270 62.800 199.105 ;
        RECT 74.070 199.090 74.390 199.350 ;
        RECT 74.990 199.290 75.310 199.350 ;
        RECT 78.760 199.335 78.900 199.490 ;
        RECT 99.945 199.490 103.835 199.630 ;
        RECT 99.945 199.445 100.535 199.490 ;
        RECT 75.925 199.290 76.215 199.335 ;
        RECT 74.990 199.150 76.215 199.290 ;
        RECT 74.990 199.090 75.310 199.150 ;
        RECT 75.925 199.105 76.215 199.150 ;
        RECT 78.685 199.105 78.975 199.335 ;
        RECT 80.970 199.090 81.290 199.350 ;
        RECT 100.245 199.130 100.535 199.445 ;
        RECT 100.750 199.430 101.070 199.490 ;
        RECT 103.185 199.445 103.835 199.490 ;
        RECT 111.330 199.630 111.650 199.690 ;
        RECT 112.265 199.630 112.555 199.675 ;
        RECT 111.330 199.490 112.555 199.630 ;
        RECT 111.330 199.430 111.650 199.490 ;
        RECT 112.265 199.445 112.555 199.490 ;
        RECT 116.505 199.630 116.795 199.675 ;
        RECT 119.745 199.630 120.395 199.675 ;
        RECT 116.505 199.490 120.395 199.630 ;
        RECT 116.505 199.445 117.095 199.490 ;
        RECT 119.745 199.445 120.395 199.490 ;
        RECT 120.990 199.630 121.310 199.690 ;
        RECT 122.385 199.630 122.675 199.675 ;
        RECT 120.990 199.490 122.675 199.630 ;
        RECT 116.805 199.350 117.095 199.445 ;
        RECT 120.990 199.430 121.310 199.490 ;
        RECT 122.385 199.445 122.675 199.490 ;
        RECT 101.325 199.290 101.615 199.335 ;
        RECT 104.905 199.290 105.195 199.335 ;
        RECT 106.740 199.290 107.030 199.335 ;
        RECT 101.325 199.150 107.030 199.290 ;
        RECT 101.325 199.105 101.615 199.150 ;
        RECT 104.905 199.105 105.195 199.150 ;
        RECT 106.740 199.105 107.030 199.150 ;
        RECT 110.410 199.290 110.730 199.350 ;
        RECT 111.805 199.290 112.095 199.335 ;
        RECT 110.410 199.150 112.095 199.290 ;
        RECT 110.410 199.090 110.730 199.150 ;
        RECT 111.805 199.105 112.095 199.150 ;
        RECT 116.805 199.130 117.170 199.350 ;
        RECT 116.850 199.090 117.170 199.130 ;
        RECT 117.885 199.290 118.175 199.335 ;
        RECT 121.465 199.290 121.755 199.335 ;
        RECT 123.300 199.290 123.590 199.335 ;
        RECT 117.885 199.150 123.590 199.290 ;
        RECT 117.885 199.105 118.175 199.150 ;
        RECT 121.465 199.105 121.755 199.150 ;
        RECT 123.300 199.105 123.590 199.150 ;
        RECT 63.490 198.750 63.810 199.010 ;
        RECT 72.230 198.950 72.550 199.010 ;
        RECT 75.450 198.950 75.770 199.010 ;
        RECT 72.230 198.810 75.770 198.950 ;
        RECT 72.230 198.750 72.550 198.810 ;
        RECT 75.450 198.750 75.770 198.810 ;
        RECT 81.445 198.950 81.735 198.995 ;
        RECT 81.890 198.950 82.210 199.010 ;
        RECT 81.445 198.810 82.210 198.950 ;
        RECT 81.445 198.765 81.735 198.810 ;
        RECT 81.890 198.750 82.210 198.810 ;
        RECT 105.810 198.750 106.130 199.010 ;
        RECT 107.205 198.950 107.495 198.995 ;
        RECT 109.030 198.950 109.350 199.010 ;
        RECT 107.205 198.810 109.350 198.950 ;
        RECT 107.205 198.765 107.495 198.810 ;
        RECT 109.030 198.750 109.350 198.810 ;
        RECT 110.870 198.750 111.190 199.010 ;
        RECT 118.690 198.950 119.010 199.010 ;
        RECT 123.765 198.950 124.055 198.995 ;
        RECT 118.690 198.810 124.055 198.950 ;
        RECT 118.690 198.750 119.010 198.810 ;
        RECT 123.765 198.765 124.055 198.810 ;
        RECT 64.375 198.610 64.665 198.655 ;
        RECT 66.265 198.610 66.555 198.655 ;
        RECT 69.385 198.610 69.675 198.655 ;
        RECT 64.375 198.470 69.675 198.610 ;
        RECT 64.375 198.425 64.665 198.470 ;
        RECT 66.265 198.425 66.555 198.470 ;
        RECT 69.385 198.425 69.675 198.470 ;
        RECT 73.165 198.610 73.455 198.655 ;
        RECT 75.910 198.610 76.230 198.670 ;
        RECT 80.970 198.610 81.290 198.670 ;
        RECT 73.165 198.470 76.230 198.610 ;
        RECT 73.165 198.425 73.455 198.470 ;
        RECT 75.910 198.410 76.230 198.470 ;
        RECT 76.460 198.470 81.290 198.610 ;
        RECT 71.310 198.270 71.630 198.330 ;
        RECT 62.660 198.130 71.630 198.270 ;
        RECT 71.310 198.070 71.630 198.130 ;
        RECT 72.230 198.270 72.550 198.330 ;
        RECT 75.465 198.270 75.755 198.315 ;
        RECT 76.460 198.270 76.600 198.470 ;
        RECT 80.970 198.410 81.290 198.470 ;
        RECT 101.325 198.610 101.615 198.655 ;
        RECT 104.445 198.610 104.735 198.655 ;
        RECT 106.335 198.610 106.625 198.655 ;
        RECT 101.325 198.470 106.625 198.610 ;
        RECT 101.325 198.425 101.615 198.470 ;
        RECT 104.445 198.425 104.735 198.470 ;
        RECT 106.335 198.425 106.625 198.470 ;
        RECT 111.790 198.610 112.110 198.670 ;
        RECT 115.025 198.610 115.315 198.655 ;
        RECT 111.790 198.470 115.315 198.610 ;
        RECT 111.790 198.410 112.110 198.470 ;
        RECT 115.025 198.425 115.315 198.470 ;
        RECT 117.885 198.610 118.175 198.655 ;
        RECT 121.005 198.610 121.295 198.655 ;
        RECT 122.895 198.610 123.185 198.655 ;
        RECT 117.885 198.470 123.185 198.610 ;
        RECT 117.885 198.425 118.175 198.470 ;
        RECT 121.005 198.425 121.295 198.470 ;
        RECT 122.895 198.425 123.185 198.470 ;
        RECT 72.230 198.130 76.600 198.270 ;
        RECT 72.230 198.070 72.550 198.130 ;
        RECT 75.465 198.085 75.755 198.130 ;
        RECT 79.130 198.070 79.450 198.330 ;
        RECT 82.350 198.070 82.670 198.330 ;
        RECT 98.450 198.070 98.770 198.330 ;
        RECT 114.105 198.270 114.395 198.315 ;
        RECT 119.610 198.270 119.930 198.330 ;
        RECT 114.105 198.130 119.930 198.270 ;
        RECT 114.105 198.085 114.395 198.130 ;
        RECT 119.610 198.070 119.930 198.130 ;
        RECT 20.640 197.450 127.820 197.930 ;
        RECT 69.945 197.250 70.235 197.295 ;
        RECT 72.690 197.250 73.010 197.310 ;
        RECT 69.945 197.110 73.010 197.250 ;
        RECT 69.945 197.065 70.235 197.110 ;
        RECT 72.690 197.050 73.010 197.110 ;
        RECT 77.750 197.250 78.070 197.310 ;
        RECT 77.750 197.110 100.520 197.250 ;
        RECT 77.750 197.050 78.070 197.110 ;
        RECT 58.905 196.725 59.195 196.955 ;
        RECT 76.370 196.910 76.690 196.970 ;
        RECT 72.780 196.770 76.690 196.910 ;
        RECT 46.470 196.570 46.790 196.630 ;
        RECT 55.685 196.570 55.975 196.615 ;
        RECT 46.470 196.430 55.975 196.570 ;
        RECT 46.470 196.370 46.790 196.430 ;
        RECT 55.685 196.385 55.975 196.430 ;
        RECT 31.290 196.230 31.610 196.290 ;
        RECT 34.525 196.230 34.815 196.275 ;
        RECT 42.345 196.230 42.635 196.275 ;
        RECT 31.290 196.090 42.635 196.230 ;
        RECT 58.980 196.230 59.120 196.725 ;
        RECT 71.310 196.570 71.630 196.630 ;
        RECT 66.800 196.430 71.630 196.570 ;
        RECT 66.800 196.275 66.940 196.430 ;
        RECT 71.310 196.370 71.630 196.430 ;
        RECT 72.230 196.370 72.550 196.630 ;
        RECT 72.780 196.615 72.920 196.770 ;
        RECT 76.370 196.710 76.690 196.770 ;
        RECT 80.165 196.910 80.455 196.955 ;
        RECT 83.285 196.910 83.575 196.955 ;
        RECT 85.175 196.910 85.465 196.955 ;
        RECT 80.165 196.770 85.465 196.910 ;
        RECT 80.165 196.725 80.455 196.770 ;
        RECT 83.285 196.725 83.575 196.770 ;
        RECT 85.175 196.725 85.465 196.770 ;
        RECT 87.430 196.910 87.720 196.955 ;
        RECT 89.290 196.910 89.580 196.955 ;
        RECT 92.070 196.910 92.360 196.955 ;
        RECT 87.430 196.770 92.360 196.910 ;
        RECT 87.430 196.725 87.720 196.770 ;
        RECT 89.290 196.725 89.580 196.770 ;
        RECT 92.070 196.725 92.360 196.770 ;
        RECT 72.705 196.385 72.995 196.615 ;
        RECT 73.610 196.570 73.930 196.630 ;
        RECT 74.990 196.570 75.310 196.630 ;
        RECT 73.610 196.430 75.310 196.570 ;
        RECT 73.610 196.370 73.930 196.430 ;
        RECT 74.990 196.370 75.310 196.430 ;
        RECT 82.350 196.570 82.670 196.630 ;
        RECT 84.665 196.570 84.955 196.615 ;
        RECT 82.350 196.430 84.955 196.570 ;
        RECT 82.350 196.370 82.670 196.430 ;
        RECT 84.665 196.385 84.955 196.430 ;
        RECT 86.490 196.570 86.810 196.630 ;
        RECT 88.805 196.570 89.095 196.615 ;
        RECT 86.490 196.430 89.095 196.570 ;
        RECT 86.490 196.370 86.810 196.430 ;
        RECT 88.805 196.385 89.095 196.430 ;
        RECT 100.380 196.570 100.520 197.110 ;
        RECT 100.750 197.050 101.070 197.310 ;
        RECT 103.985 197.250 104.275 197.295 ;
        RECT 105.810 197.250 106.130 197.310 ;
        RECT 103.985 197.110 106.130 197.250 ;
        RECT 103.985 197.065 104.275 197.110 ;
        RECT 105.810 197.050 106.130 197.110 ;
        RECT 112.365 196.910 112.655 196.955 ;
        RECT 115.485 196.910 115.775 196.955 ;
        RECT 117.375 196.910 117.665 196.955 ;
        RECT 112.365 196.770 117.665 196.910 ;
        RECT 112.365 196.725 112.655 196.770 ;
        RECT 115.485 196.725 115.775 196.770 ;
        RECT 117.375 196.725 117.665 196.770 ;
        RECT 118.705 196.725 118.995 196.955 ;
        RECT 109.505 196.570 109.795 196.615 ;
        RECT 110.410 196.570 110.730 196.630 ;
        RECT 100.380 196.430 108.340 196.570 ;
        RECT 59.825 196.230 60.115 196.275 ;
        RECT 58.980 196.090 60.115 196.230 ;
        RECT 31.290 196.030 31.610 196.090 ;
        RECT 34.525 196.045 34.815 196.090 ;
        RECT 42.345 196.045 42.635 196.090 ;
        RECT 59.825 196.045 60.115 196.090 ;
        RECT 66.725 196.045 67.015 196.275 ;
        RECT 73.165 196.230 73.455 196.275 ;
        RECT 74.530 196.230 74.850 196.290 ;
        RECT 79.130 196.250 79.450 196.290 ;
        RECT 69.100 196.090 72.920 196.230 ;
        RECT 46.945 195.890 47.235 195.935 ;
        RECT 51.070 195.890 51.390 195.950 ;
        RECT 54.750 195.890 55.070 195.950 ;
        RECT 69.100 195.935 69.240 196.090 ;
        RECT 57.065 195.890 57.355 195.935 ;
        RECT 46.945 195.750 57.355 195.890 ;
        RECT 46.945 195.705 47.235 195.750 ;
        RECT 51.070 195.690 51.390 195.750 ;
        RECT 54.750 195.690 55.070 195.750 ;
        RECT 57.065 195.705 57.355 195.750 ;
        RECT 69.025 195.705 69.315 195.935 ;
        RECT 70.105 195.890 70.395 195.935 ;
        RECT 72.780 195.890 72.920 196.090 ;
        RECT 73.165 196.090 74.850 196.230 ;
        RECT 73.165 196.045 73.455 196.090 ;
        RECT 74.530 196.030 74.850 196.090 ;
        RECT 79.085 196.030 79.450 196.250 ;
        RECT 80.165 196.230 80.455 196.275 ;
        RECT 83.745 196.230 84.035 196.275 ;
        RECT 85.580 196.230 85.870 196.275 ;
        RECT 80.165 196.090 85.870 196.230 ;
        RECT 80.165 196.045 80.455 196.090 ;
        RECT 83.745 196.045 84.035 196.090 ;
        RECT 85.580 196.045 85.870 196.090 ;
        RECT 86.045 196.230 86.335 196.275 ;
        RECT 86.965 196.230 87.255 196.275 ;
        RECT 88.330 196.230 88.650 196.290 ;
        RECT 100.380 196.275 100.520 196.430 ;
        RECT 92.070 196.230 92.360 196.275 ;
        RECT 86.045 196.090 88.650 196.230 ;
        RECT 86.045 196.045 86.335 196.090 ;
        RECT 86.965 196.045 87.255 196.090 ;
        RECT 88.330 196.030 88.650 196.090 ;
        RECT 89.825 196.090 92.360 196.230 ;
        RECT 75.910 195.890 76.230 195.950 ;
        RECT 79.085 195.935 79.375 196.030 ;
        RECT 89.825 195.935 90.040 196.090 ;
        RECT 92.070 196.045 92.360 196.090 ;
        RECT 100.305 196.045 100.595 196.275 ;
        RECT 103.050 196.030 103.370 196.290 ;
        RECT 108.200 196.275 108.340 196.430 ;
        RECT 109.505 196.430 110.730 196.570 ;
        RECT 109.505 196.385 109.795 196.430 ;
        RECT 110.410 196.370 110.730 196.430 ;
        RECT 116.865 196.570 117.155 196.615 ;
        RECT 118.780 196.570 118.920 196.725 ;
        RECT 116.865 196.430 118.920 196.570 ;
        RECT 116.865 196.385 117.155 196.430 ;
        RECT 108.125 196.230 108.415 196.275 ;
        RECT 109.950 196.230 110.270 196.290 ;
        RECT 108.125 196.090 110.270 196.230 ;
        RECT 108.125 196.045 108.415 196.090 ;
        RECT 109.950 196.030 110.270 196.090 ;
        RECT 111.285 195.935 111.575 196.250 ;
        RECT 112.365 196.230 112.655 196.275 ;
        RECT 115.945 196.230 116.235 196.275 ;
        RECT 117.780 196.230 118.070 196.275 ;
        RECT 112.365 196.090 118.070 196.230 ;
        RECT 112.365 196.045 112.655 196.090 ;
        RECT 115.945 196.045 116.235 196.090 ;
        RECT 117.780 196.045 118.070 196.090 ;
        RECT 118.230 196.030 118.550 196.290 ;
        RECT 119.610 196.030 119.930 196.290 ;
        RECT 70.105 195.750 71.540 195.890 ;
        RECT 72.780 195.750 76.230 195.890 ;
        RECT 70.105 195.705 70.395 195.750 ;
        RECT 34.065 195.550 34.355 195.595 ;
        RECT 34.510 195.550 34.830 195.610 ;
        RECT 34.065 195.410 34.830 195.550 ;
        RECT 34.065 195.365 34.355 195.410 ;
        RECT 34.510 195.350 34.830 195.410 ;
        RECT 42.790 195.350 43.110 195.610 ;
        RECT 43.710 195.550 44.030 195.610 ;
        RECT 47.405 195.550 47.695 195.595 ;
        RECT 43.710 195.410 47.695 195.550 ;
        RECT 43.710 195.350 44.030 195.410 ;
        RECT 47.405 195.365 47.695 195.410 ;
        RECT 49.245 195.550 49.535 195.595 ;
        RECT 50.150 195.550 50.470 195.610 ;
        RECT 49.245 195.410 50.470 195.550 ;
        RECT 49.245 195.365 49.535 195.410 ;
        RECT 50.150 195.350 50.470 195.410 ;
        RECT 56.130 195.550 56.450 195.610 ;
        RECT 56.605 195.550 56.895 195.595 ;
        RECT 56.130 195.410 56.895 195.550 ;
        RECT 56.130 195.350 56.450 195.410 ;
        RECT 56.605 195.365 56.895 195.410 ;
        RECT 60.745 195.550 61.035 195.595 ;
        RECT 61.190 195.550 61.510 195.610 ;
        RECT 60.745 195.410 61.510 195.550 ;
        RECT 60.745 195.365 61.035 195.410 ;
        RECT 61.190 195.350 61.510 195.410 ;
        RECT 67.170 195.350 67.490 195.610 ;
        RECT 70.850 195.350 71.170 195.610 ;
        RECT 71.400 195.595 71.540 195.750 ;
        RECT 75.910 195.690 76.230 195.750 ;
        RECT 78.785 195.890 79.375 195.935 ;
        RECT 82.025 195.890 82.675 195.935 ;
        RECT 78.785 195.750 82.675 195.890 ;
        RECT 78.785 195.705 79.075 195.750 ;
        RECT 82.025 195.705 82.675 195.750 ;
        RECT 87.890 195.890 88.180 195.935 ;
        RECT 89.750 195.890 90.040 195.935 ;
        RECT 90.670 195.890 90.960 195.935 ;
        RECT 93.930 195.890 94.220 195.935 ;
        RECT 87.890 195.750 90.040 195.890 ;
        RECT 87.890 195.705 88.180 195.750 ;
        RECT 89.750 195.705 90.040 195.750 ;
        RECT 90.260 195.750 94.220 195.890 ;
        RECT 71.325 195.365 71.615 195.595 ;
        RECT 74.990 195.550 75.310 195.610 ;
        RECT 77.305 195.550 77.595 195.595 ;
        RECT 74.990 195.410 77.595 195.550 ;
        RECT 74.990 195.350 75.310 195.410 ;
        RECT 77.305 195.365 77.595 195.410 ;
        RECT 86.490 195.550 86.810 195.610 ;
        RECT 90.260 195.550 90.400 195.750 ;
        RECT 90.670 195.705 90.960 195.750 ;
        RECT 93.930 195.705 94.220 195.750 ;
        RECT 108.585 195.890 108.875 195.935 ;
        RECT 110.985 195.890 111.575 195.935 ;
        RECT 114.225 195.890 114.875 195.935 ;
        RECT 108.585 195.750 114.875 195.890 ;
        RECT 108.585 195.705 108.875 195.750 ;
        RECT 110.985 195.705 111.275 195.750 ;
        RECT 114.225 195.705 114.875 195.750 ;
        RECT 86.490 195.410 90.400 195.550 ;
        RECT 95.935 195.550 96.225 195.595 ;
        RECT 97.990 195.550 98.310 195.610 ;
        RECT 95.935 195.410 98.310 195.550 ;
        RECT 86.490 195.350 86.810 195.410 ;
        RECT 95.935 195.365 96.225 195.410 ;
        RECT 97.990 195.350 98.310 195.410 ;
        RECT 20.640 194.730 127.820 195.210 ;
        RECT 48.785 194.345 49.075 194.575 ;
        RECT 49.230 194.530 49.550 194.590 ;
        RECT 50.165 194.530 50.455 194.575 ;
        RECT 49.230 194.390 50.455 194.530 ;
        RECT 29.450 193.990 29.770 194.250 ;
        RECT 31.745 194.190 32.395 194.235 ;
        RECT 34.510 194.190 34.830 194.250 ;
        RECT 35.345 194.190 35.635 194.235 ;
        RECT 31.745 194.050 35.635 194.190 ;
        RECT 31.745 194.005 32.395 194.050 ;
        RECT 34.510 193.990 34.830 194.050 ;
        RECT 35.045 194.005 35.635 194.050 ;
        RECT 41.360 194.190 41.650 194.235 ;
        RECT 42.790 194.190 43.110 194.250 ;
        RECT 44.620 194.190 44.910 194.235 ;
        RECT 41.360 194.050 44.910 194.190 ;
        RECT 41.360 194.005 41.650 194.050 ;
        RECT 28.550 193.850 28.840 193.895 ;
        RECT 30.385 193.850 30.675 193.895 ;
        RECT 33.965 193.850 34.255 193.895 ;
        RECT 28.550 193.710 34.255 193.850 ;
        RECT 28.550 193.665 28.840 193.710 ;
        RECT 30.385 193.665 30.675 193.710 ;
        RECT 33.965 193.665 34.255 193.710 ;
        RECT 35.045 193.690 35.335 194.005 ;
        RECT 42.790 193.990 43.110 194.050 ;
        RECT 44.620 194.005 44.910 194.050 ;
        RECT 45.540 194.190 45.830 194.235 ;
        RECT 47.400 194.190 47.690 194.235 ;
        RECT 45.540 194.050 47.690 194.190 ;
        RECT 45.540 194.005 45.830 194.050 ;
        RECT 47.400 194.005 47.690 194.050 ;
        RECT 43.220 193.850 43.510 193.895 ;
        RECT 45.540 193.850 45.755 194.005 ;
        RECT 43.220 193.710 45.755 193.850 ;
        RECT 43.220 193.665 43.510 193.710 ;
        RECT 46.010 193.650 46.330 193.910 ;
        RECT 46.485 193.850 46.775 193.895 ;
        RECT 48.860 193.850 49.000 194.345 ;
        RECT 49.230 194.330 49.550 194.390 ;
        RECT 50.165 194.345 50.455 194.390 ;
        RECT 52.005 194.530 52.295 194.575 ;
        RECT 52.450 194.530 52.770 194.590 ;
        RECT 73.610 194.530 73.930 194.590 ;
        RECT 52.005 194.390 52.770 194.530 ;
        RECT 52.005 194.345 52.295 194.390 ;
        RECT 52.450 194.330 52.770 194.390 ;
        RECT 63.580 194.390 73.930 194.530 ;
        RECT 55.325 194.190 55.615 194.235 ;
        RECT 57.510 194.190 57.830 194.250 ;
        RECT 58.565 194.190 59.215 194.235 ;
        RECT 55.325 194.050 59.215 194.190 ;
        RECT 55.325 194.005 55.915 194.050 ;
        RECT 46.485 193.710 49.000 193.850 ;
        RECT 46.485 193.665 46.775 193.710 ;
        RECT 49.690 193.650 50.010 193.910 ;
        RECT 50.150 193.850 50.470 193.910 ;
        RECT 51.085 193.850 51.375 193.895 ;
        RECT 50.150 193.710 51.375 193.850 ;
        RECT 50.150 193.650 50.470 193.710 ;
        RECT 51.085 193.665 51.375 193.710 ;
        RECT 52.465 193.665 52.755 193.895 ;
        RECT 55.625 193.690 55.915 194.005 ;
        RECT 57.510 193.990 57.830 194.050 ;
        RECT 58.565 194.005 59.215 194.050 ;
        RECT 61.190 193.990 61.510 194.250 ;
        RECT 63.580 194.235 63.720 194.390 ;
        RECT 73.610 194.330 73.930 194.390 ;
        RECT 74.070 194.330 74.390 194.590 ;
        RECT 80.050 194.530 80.370 194.590 ;
        RECT 78.300 194.390 80.370 194.530 ;
        RECT 63.505 194.005 63.795 194.235 ;
        RECT 66.365 194.190 66.655 194.235 ;
        RECT 67.170 194.190 67.490 194.250 ;
        RECT 69.605 194.190 70.255 194.235 ;
        RECT 66.365 194.050 70.255 194.190 ;
        RECT 66.365 194.005 66.955 194.050 ;
        RECT 56.705 193.850 56.995 193.895 ;
        RECT 60.285 193.850 60.575 193.895 ;
        RECT 62.120 193.850 62.410 193.895 ;
        RECT 56.705 193.710 62.410 193.850 ;
        RECT 56.705 193.665 56.995 193.710 ;
        RECT 60.285 193.665 60.575 193.710 ;
        RECT 62.120 193.665 62.410 193.710 ;
        RECT 66.665 193.690 66.955 194.005 ;
        RECT 67.170 193.990 67.490 194.050 ;
        RECT 69.605 194.005 70.255 194.050 ;
        RECT 72.230 193.990 72.550 194.250 ;
        RECT 78.300 194.235 78.440 194.390 ;
        RECT 80.050 194.330 80.370 194.390 ;
        RECT 80.525 194.530 80.815 194.575 ;
        RECT 80.970 194.530 81.290 194.590 ;
        RECT 80.525 194.390 81.290 194.530 ;
        RECT 80.525 194.345 80.815 194.390 ;
        RECT 80.970 194.330 81.290 194.390 ;
        RECT 85.585 194.530 85.875 194.575 ;
        RECT 86.030 194.530 86.350 194.590 ;
        RECT 85.585 194.390 86.350 194.530 ;
        RECT 85.585 194.345 85.875 194.390 ;
        RECT 86.030 194.330 86.350 194.390 ;
        RECT 86.490 194.330 86.810 194.590 ;
        RECT 102.605 194.530 102.895 194.575 ;
        RECT 103.050 194.530 103.370 194.590 ;
        RECT 111.330 194.530 111.650 194.590 ;
        RECT 102.605 194.390 103.370 194.530 ;
        RECT 102.605 194.345 102.895 194.390 ;
        RECT 103.050 194.330 103.370 194.390 ;
        RECT 105.440 194.390 111.650 194.530 ;
        RECT 78.225 194.190 78.515 194.235 ;
        RECT 87.885 194.190 88.175 194.235 ;
        RECT 91.500 194.190 91.790 194.235 ;
        RECT 94.760 194.190 95.050 194.235 ;
        RECT 75.540 194.050 78.515 194.190 ;
        RECT 67.745 193.850 68.035 193.895 ;
        RECT 71.325 193.850 71.615 193.895 ;
        RECT 73.160 193.850 73.450 193.895 ;
        RECT 67.745 193.710 73.450 193.850 ;
        RECT 67.745 193.665 68.035 193.710 ;
        RECT 71.325 193.665 71.615 193.710 ;
        RECT 73.160 193.665 73.450 193.710 ;
        RECT 74.530 193.850 74.850 193.910 ;
        RECT 75.540 193.895 75.680 194.050 ;
        RECT 78.225 194.005 78.515 194.050 ;
        RECT 79.220 194.050 82.580 194.190 ;
        RECT 75.465 193.850 75.755 193.895 ;
        RECT 74.530 193.710 75.755 193.850 ;
        RECT 28.070 193.510 28.390 193.570 ;
        RECT 46.100 193.510 46.240 193.650 ;
        RECT 48.325 193.510 48.615 193.555 ;
        RECT 49.230 193.510 49.550 193.570 ;
        RECT 28.070 193.370 49.550 193.510 ;
        RECT 52.540 193.510 52.680 193.665 ;
        RECT 74.530 193.650 74.850 193.710 ;
        RECT 75.465 193.665 75.755 193.710 ;
        RECT 76.370 193.850 76.690 193.910 ;
        RECT 79.220 193.895 79.360 194.050 ;
        RECT 76.845 193.850 77.135 193.895 ;
        RECT 79.145 193.850 79.435 193.895 ;
        RECT 76.370 193.710 79.435 193.850 ;
        RECT 76.370 193.650 76.690 193.710 ;
        RECT 76.845 193.665 77.135 193.710 ;
        RECT 79.145 193.665 79.435 193.710 ;
        RECT 79.605 193.665 79.895 193.895 ;
        RECT 80.050 193.850 80.370 193.910 ;
        RECT 82.440 193.895 82.580 194.050 ;
        RECT 87.885 194.050 95.050 194.190 ;
        RECT 87.885 194.005 88.175 194.050 ;
        RECT 91.500 194.005 91.790 194.050 ;
        RECT 94.760 194.005 95.050 194.050 ;
        RECT 95.680 194.190 95.970 194.235 ;
        RECT 97.540 194.190 97.830 194.235 ;
        RECT 95.680 194.050 97.830 194.190 ;
        RECT 95.680 194.005 95.970 194.050 ;
        RECT 97.540 194.005 97.830 194.050 ;
        RECT 98.450 194.190 98.770 194.250 ;
        RECT 100.305 194.190 100.595 194.235 ;
        RECT 105.440 194.190 105.580 194.390 ;
        RECT 111.330 194.330 111.650 194.390 ;
        RECT 111.790 194.330 112.110 194.590 ;
        RECT 116.405 194.530 116.695 194.575 ;
        RECT 116.850 194.530 117.170 194.590 ;
        RECT 116.405 194.390 117.170 194.530 ;
        RECT 116.405 194.345 116.695 194.390 ;
        RECT 116.850 194.330 117.170 194.390 ;
        RECT 120.085 194.530 120.375 194.575 ;
        RECT 120.990 194.530 121.310 194.590 ;
        RECT 120.085 194.390 121.310 194.530 ;
        RECT 120.085 194.345 120.375 194.390 ;
        RECT 120.990 194.330 121.310 194.390 ;
        RECT 98.450 194.050 105.580 194.190 ;
        RECT 109.950 194.190 110.270 194.250 ;
        RECT 109.950 194.050 116.160 194.190 ;
        RECT 81.445 193.850 81.735 193.895 ;
        RECT 80.050 193.710 81.735 193.850 ;
        RECT 57.970 193.510 58.290 193.570 ;
        RECT 52.540 193.370 58.290 193.510 ;
        RECT 28.070 193.310 28.390 193.370 ;
        RECT 48.325 193.325 48.615 193.370 ;
        RECT 49.230 193.310 49.550 193.370 ;
        RECT 57.970 193.310 58.290 193.370 ;
        RECT 62.585 193.510 62.875 193.555 ;
        RECT 63.950 193.510 64.270 193.570 ;
        RECT 73.625 193.510 73.915 193.555 ;
        RECT 62.585 193.370 73.915 193.510 ;
        RECT 62.585 193.325 62.875 193.370 ;
        RECT 63.950 193.310 64.270 193.370 ;
        RECT 73.625 193.325 73.915 193.370 ;
        RECT 74.990 193.510 75.310 193.570 ;
        RECT 79.680 193.510 79.820 193.665 ;
        RECT 80.050 193.650 80.370 193.710 ;
        RECT 81.445 193.665 81.735 193.710 ;
        RECT 82.365 193.665 82.655 193.895 ;
        RECT 84.650 193.650 84.970 193.910 ;
        RECT 86.965 193.850 87.255 193.895 ;
        RECT 87.425 193.850 87.715 193.895 ;
        RECT 90.630 193.850 90.950 193.910 ;
        RECT 86.965 193.710 90.950 193.850 ;
        RECT 86.965 193.665 87.255 193.710 ;
        RECT 87.425 193.665 87.715 193.710 ;
        RECT 90.630 193.650 90.950 193.710 ;
        RECT 93.360 193.850 93.650 193.895 ;
        RECT 95.680 193.850 95.895 194.005 ;
        RECT 98.450 193.990 98.770 194.050 ;
        RECT 100.305 194.005 100.595 194.050 ;
        RECT 109.950 193.990 110.270 194.050 ;
        RECT 93.360 193.710 95.895 193.850 ;
        RECT 93.360 193.665 93.650 193.710 ;
        RECT 96.610 193.650 96.930 193.910 ;
        RECT 97.990 193.850 98.310 193.910 ;
        RECT 100.765 193.850 101.055 193.895 ;
        RECT 97.990 193.710 101.055 193.850 ;
        RECT 97.990 193.650 98.310 193.710 ;
        RECT 100.765 193.665 101.055 193.710 ;
        RECT 110.410 193.850 110.730 193.910 ;
        RECT 116.020 193.895 116.160 194.050 ;
        RECT 112.265 193.850 112.555 193.895 ;
        RECT 110.410 193.710 112.555 193.850 ;
        RECT 110.410 193.650 110.730 193.710 ;
        RECT 112.265 193.665 112.555 193.710 ;
        RECT 115.945 193.665 116.235 193.895 ;
        RECT 119.165 193.665 119.455 193.895 ;
        RECT 74.990 193.370 79.820 193.510 ;
        RECT 88.790 193.510 89.110 193.570 ;
        RECT 98.465 193.510 98.755 193.555 ;
        RECT 88.790 193.370 98.755 193.510 ;
        RECT 74.990 193.310 75.310 193.370 ;
        RECT 88.790 193.310 89.110 193.370 ;
        RECT 98.465 193.325 98.755 193.370 ;
        RECT 99.845 193.325 100.135 193.555 ;
        RECT 28.955 193.170 29.245 193.215 ;
        RECT 30.845 193.170 31.135 193.215 ;
        RECT 33.965 193.170 34.255 193.215 ;
        RECT 28.955 193.030 34.255 193.170 ;
        RECT 28.955 192.985 29.245 193.030 ;
        RECT 30.845 192.985 31.135 193.030 ;
        RECT 33.965 192.985 34.255 193.030 ;
        RECT 43.220 193.170 43.510 193.215 ;
        RECT 46.000 193.170 46.290 193.215 ;
        RECT 47.860 193.170 48.150 193.215 ;
        RECT 43.220 193.030 48.150 193.170 ;
        RECT 43.220 192.985 43.510 193.030 ;
        RECT 46.000 192.985 46.290 193.030 ;
        RECT 47.860 192.985 48.150 193.030 ;
        RECT 56.705 193.170 56.995 193.215 ;
        RECT 59.825 193.170 60.115 193.215 ;
        RECT 61.715 193.170 62.005 193.215 ;
        RECT 56.705 193.030 62.005 193.170 ;
        RECT 56.705 192.985 56.995 193.030 ;
        RECT 59.825 192.985 60.115 193.030 ;
        RECT 61.715 192.985 62.005 193.030 ;
        RECT 67.745 193.170 68.035 193.215 ;
        RECT 70.865 193.170 71.155 193.215 ;
        RECT 72.755 193.170 73.045 193.215 ;
        RECT 67.745 193.030 73.045 193.170 ;
        RECT 67.745 192.985 68.035 193.030 ;
        RECT 70.865 192.985 71.155 193.030 ;
        RECT 72.755 192.985 73.045 193.030 ;
        RECT 93.360 193.170 93.650 193.215 ;
        RECT 96.140 193.170 96.430 193.215 ;
        RECT 98.000 193.170 98.290 193.215 ;
        RECT 93.360 193.030 98.290 193.170 ;
        RECT 99.920 193.170 100.060 193.325 ;
        RECT 110.870 193.310 111.190 193.570 ;
        RECT 119.240 193.510 119.380 193.665 ;
        RECT 114.180 193.370 119.380 193.510 ;
        RECT 106.270 193.170 106.590 193.230 ;
        RECT 110.960 193.170 111.100 193.310 ;
        RECT 114.180 193.215 114.320 193.370 ;
        RECT 99.920 193.030 111.100 193.170 ;
        RECT 93.360 192.985 93.650 193.030 ;
        RECT 96.140 192.985 96.430 193.030 ;
        RECT 98.000 192.985 98.290 193.030 ;
        RECT 106.270 192.970 106.590 193.030 ;
        RECT 114.105 192.985 114.395 193.215 ;
        RECT 36.825 192.830 37.115 192.875 ;
        RECT 37.730 192.830 38.050 192.890 ;
        RECT 36.825 192.690 38.050 192.830 ;
        RECT 36.825 192.645 37.115 192.690 ;
        RECT 37.730 192.630 38.050 192.690 ;
        RECT 39.355 192.830 39.645 192.875 ;
        RECT 40.030 192.830 40.350 192.890 ;
        RECT 39.355 192.690 40.350 192.830 ;
        RECT 39.355 192.645 39.645 192.690 ;
        RECT 40.030 192.630 40.350 192.690 ;
        RECT 53.845 192.830 54.135 192.875 ;
        RECT 56.130 192.830 56.450 192.890 ;
        RECT 53.845 192.690 56.450 192.830 ;
        RECT 53.845 192.645 54.135 192.690 ;
        RECT 56.130 192.630 56.450 192.690 ;
        RECT 75.450 192.630 75.770 192.890 ;
        RECT 77.290 192.630 77.610 192.890 ;
        RECT 81.890 192.630 82.210 192.890 ;
        RECT 89.250 192.875 89.570 192.890 ;
        RECT 89.250 192.645 89.785 192.875 ;
        RECT 89.250 192.630 89.570 192.645 ;
        RECT 20.640 192.010 127.820 192.490 ;
        RECT 46.025 191.810 46.315 191.855 ;
        RECT 49.690 191.810 50.010 191.870 ;
        RECT 46.025 191.670 50.010 191.810 ;
        RECT 46.025 191.625 46.315 191.670 ;
        RECT 49.690 191.610 50.010 191.670 ;
        RECT 57.510 191.610 57.830 191.870 ;
        RECT 71.785 191.810 72.075 191.855 ;
        RECT 72.230 191.810 72.550 191.870 ;
        RECT 71.785 191.670 72.550 191.810 ;
        RECT 71.785 191.625 72.075 191.670 ;
        RECT 72.230 191.610 72.550 191.670 ;
        RECT 72.690 191.810 73.010 191.870 ;
        RECT 74.085 191.810 74.375 191.855 ;
        RECT 72.690 191.670 74.375 191.810 ;
        RECT 72.690 191.610 73.010 191.670 ;
        RECT 74.085 191.625 74.375 191.670 ;
        RECT 77.290 191.810 77.610 191.870 ;
        RECT 77.765 191.810 78.055 191.855 ;
        RECT 77.290 191.670 78.055 191.810 ;
        RECT 77.290 191.610 77.610 191.670 ;
        RECT 77.765 191.625 78.055 191.670 ;
        RECT 84.650 191.810 84.970 191.870 ;
        RECT 89.265 191.810 89.555 191.855 ;
        RECT 84.650 191.670 89.555 191.810 ;
        RECT 84.650 191.610 84.970 191.670 ;
        RECT 89.265 191.625 89.555 191.670 ;
        RECT 94.325 191.810 94.615 191.855 ;
        RECT 96.610 191.810 96.930 191.870 ;
        RECT 94.325 191.670 96.930 191.810 ;
        RECT 94.325 191.625 94.615 191.670 ;
        RECT 96.610 191.610 96.930 191.670 ;
        RECT 29.450 191.470 29.770 191.530 ;
        RECT 34.065 191.470 34.355 191.515 ;
        RECT 29.450 191.330 34.355 191.470 ;
        RECT 29.450 191.270 29.770 191.330 ;
        RECT 34.065 191.285 34.355 191.330 ;
        RECT 35.445 191.285 35.735 191.515 ;
        RECT 73.150 191.470 73.470 191.530 ;
        RECT 111.445 191.470 111.735 191.515 ;
        RECT 114.565 191.470 114.855 191.515 ;
        RECT 116.455 191.470 116.745 191.515 ;
        RECT 73.150 191.330 75.680 191.470 ;
        RECT 31.290 190.790 31.610 190.850 ;
        RECT 31.765 190.790 32.055 190.835 ;
        RECT 31.290 190.650 32.055 190.790 ;
        RECT 31.290 190.590 31.610 190.650 ;
        RECT 31.765 190.605 32.055 190.650 ;
        RECT 34.985 190.790 35.275 190.835 ;
        RECT 35.520 190.790 35.660 191.285 ;
        RECT 73.150 191.270 73.470 191.330 ;
        RECT 38.665 191.130 38.955 191.175 ;
        RECT 43.250 191.130 43.570 191.190 ;
        RECT 46.470 191.130 46.790 191.190 ;
        RECT 38.665 190.990 46.790 191.130 ;
        RECT 38.665 190.945 38.955 190.990 ;
        RECT 43.250 190.930 43.570 190.990 ;
        RECT 46.470 190.930 46.790 190.990 ;
        RECT 69.470 191.130 69.790 191.190 ;
        RECT 73.625 191.130 73.915 191.175 ;
        RECT 74.530 191.130 74.850 191.190 ;
        RECT 69.470 190.990 74.850 191.130 ;
        RECT 69.470 190.930 69.790 190.990 ;
        RECT 73.625 190.945 73.915 190.990 ;
        RECT 74.530 190.930 74.850 190.990 ;
        RECT 34.985 190.650 35.660 190.790 ;
        RECT 34.985 190.605 35.275 190.650 ;
        RECT 53.845 190.605 54.135 190.835 ;
        RECT 54.750 190.790 55.070 190.850 ;
        RECT 55.685 190.790 55.975 190.835 ;
        RECT 54.750 190.650 55.975 190.790 ;
        RECT 37.730 190.450 38.050 190.510 ;
        RECT 53.920 190.450 54.060 190.605 ;
        RECT 54.750 190.590 55.070 190.650 ;
        RECT 55.685 190.605 55.975 190.650 ;
        RECT 57.970 190.790 58.290 190.850 ;
        RECT 61.190 190.790 61.510 190.850 ;
        RECT 57.970 190.650 61.510 190.790 ;
        RECT 57.970 190.590 58.290 190.650 ;
        RECT 61.190 190.590 61.510 190.650 ;
        RECT 70.850 190.590 71.170 190.850 ;
        RECT 71.770 190.790 72.090 190.850 ;
        RECT 74.070 190.790 74.390 190.850 ;
        RECT 75.540 190.835 75.680 191.330 ;
        RECT 111.445 191.330 116.745 191.470 ;
        RECT 111.445 191.285 111.735 191.330 ;
        RECT 114.565 191.285 114.855 191.330 ;
        RECT 116.455 191.285 116.745 191.330 ;
        RECT 81.890 191.130 82.210 191.190 ;
        RECT 76.920 190.990 82.210 191.130 ;
        RECT 75.005 190.790 75.295 190.835 ;
        RECT 71.770 190.650 75.295 190.790 ;
        RECT 71.770 190.590 72.090 190.650 ;
        RECT 74.070 190.590 74.390 190.650 ;
        RECT 75.005 190.605 75.295 190.650 ;
        RECT 75.465 190.605 75.755 190.835 ;
        RECT 58.060 190.450 58.200 190.590 ;
        RECT 76.370 190.450 76.690 190.510 ;
        RECT 76.920 190.495 77.060 190.990 ;
        RECT 81.890 190.930 82.210 190.990 ;
        RECT 91.550 191.130 91.870 191.190 ;
        RECT 92.025 191.130 92.315 191.175 ;
        RECT 91.550 190.990 92.315 191.130 ;
        RECT 91.550 190.930 91.870 190.990 ;
        RECT 92.025 190.945 92.315 190.990 ;
        RECT 109.030 191.130 109.350 191.190 ;
        RECT 117.325 191.130 117.615 191.175 ;
        RECT 118.230 191.130 118.550 191.190 ;
        RECT 109.030 190.990 118.550 191.130 ;
        RECT 109.030 190.930 109.350 190.990 ;
        RECT 117.325 190.945 117.615 190.990 ;
        RECT 118.230 190.930 118.550 190.990 ;
        RECT 79.145 190.790 79.435 190.835 ;
        RECT 78.760 190.650 79.435 190.790 ;
        RECT 37.730 190.310 44.400 190.450 ;
        RECT 53.920 190.310 58.200 190.450 ;
        RECT 74.620 190.310 76.690 190.450 ;
        RECT 37.730 190.250 38.050 190.310 ;
        RECT 32.210 189.910 32.530 190.170 ;
        RECT 36.810 190.110 37.130 190.170 ;
        RECT 37.285 190.110 37.575 190.155 ;
        RECT 36.810 189.970 37.575 190.110 ;
        RECT 36.810 189.910 37.130 189.970 ;
        RECT 37.285 189.925 37.575 189.970 ;
        RECT 40.030 190.110 40.350 190.170 ;
        RECT 43.710 190.110 44.030 190.170 ;
        RECT 44.260 190.155 44.400 190.310 ;
        RECT 40.030 189.970 44.030 190.110 ;
        RECT 40.030 189.910 40.350 189.970 ;
        RECT 43.710 189.910 44.030 189.970 ;
        RECT 44.185 190.110 44.475 190.155 ;
        RECT 46.010 190.110 46.330 190.170 ;
        RECT 44.185 189.970 46.330 190.110 ;
        RECT 44.185 189.925 44.475 189.970 ;
        RECT 46.010 189.910 46.330 189.970 ;
        RECT 53.370 189.910 53.690 190.170 ;
        RECT 56.590 189.910 56.910 190.170 ;
        RECT 70.390 190.110 70.710 190.170 ;
        RECT 74.620 190.155 74.760 190.310 ;
        RECT 76.370 190.250 76.690 190.310 ;
        RECT 76.845 190.265 77.135 190.495 ;
        RECT 74.545 190.110 74.835 190.155 ;
        RECT 70.390 189.970 74.835 190.110 ;
        RECT 70.390 189.910 70.710 189.970 ;
        RECT 74.545 189.925 74.835 189.970 ;
        RECT 75.910 190.110 76.230 190.170 ;
        RECT 78.760 190.155 78.900 190.650 ;
        RECT 79.145 190.605 79.435 190.650 ;
        RECT 93.390 190.590 93.710 190.850 ;
        RECT 90.170 190.450 90.490 190.510 ;
        RECT 91.565 190.450 91.855 190.495 ;
        RECT 97.990 190.450 98.310 190.510 ;
        RECT 110.365 190.495 110.655 190.810 ;
        RECT 111.445 190.790 111.735 190.835 ;
        RECT 115.025 190.790 115.315 190.835 ;
        RECT 116.860 190.790 117.150 190.835 ;
        RECT 111.445 190.650 117.150 190.790 ;
        RECT 111.445 190.605 111.735 190.650 ;
        RECT 115.025 190.605 115.315 190.650 ;
        RECT 116.860 190.605 117.150 190.650 ;
        RECT 119.150 190.790 119.470 190.850 ;
        RECT 120.545 190.790 120.835 190.835 ;
        RECT 119.150 190.650 120.835 190.790 ;
        RECT 119.150 190.590 119.470 190.650 ;
        RECT 120.545 190.605 120.835 190.650 ;
        RECT 90.170 190.310 98.310 190.450 ;
        RECT 90.170 190.250 90.490 190.310 ;
        RECT 91.565 190.265 91.855 190.310 ;
        RECT 97.990 190.250 98.310 190.310 ;
        RECT 110.065 190.450 110.655 190.495 ;
        RECT 112.250 190.450 112.570 190.510 ;
        RECT 113.305 190.450 113.955 190.495 ;
        RECT 110.065 190.310 113.955 190.450 ;
        RECT 110.065 190.265 110.355 190.310 ;
        RECT 112.250 190.250 112.570 190.310 ;
        RECT 113.305 190.265 113.955 190.310 ;
        RECT 115.930 190.250 116.250 190.510 ;
        RECT 77.845 190.110 78.135 190.155 ;
        RECT 75.910 189.970 78.135 190.110 ;
        RECT 75.910 189.910 76.230 189.970 ;
        RECT 77.845 189.925 78.135 189.970 ;
        RECT 78.685 189.925 78.975 190.155 ;
        RECT 80.065 190.110 80.355 190.155 ;
        RECT 80.970 190.110 81.290 190.170 ;
        RECT 80.065 189.970 81.290 190.110 ;
        RECT 80.065 189.925 80.355 189.970 ;
        RECT 80.970 189.910 81.290 189.970 ;
        RECT 86.030 190.110 86.350 190.170 ;
        RECT 89.250 190.110 89.570 190.170 ;
        RECT 91.105 190.110 91.395 190.155 ;
        RECT 86.030 189.970 91.395 190.110 ;
        RECT 86.030 189.910 86.350 189.970 ;
        RECT 89.250 189.910 89.570 189.970 ;
        RECT 91.105 189.925 91.395 189.970 ;
        RECT 105.810 190.110 106.130 190.170 ;
        RECT 108.585 190.110 108.875 190.155 ;
        RECT 105.810 189.970 108.875 190.110 ;
        RECT 105.810 189.910 106.130 189.970 ;
        RECT 108.585 189.925 108.875 189.970 ;
        RECT 121.465 190.110 121.755 190.155 ;
        RECT 123.290 190.110 123.610 190.170 ;
        RECT 121.465 189.970 123.610 190.110 ;
        RECT 121.465 189.925 121.755 189.970 ;
        RECT 123.290 189.910 123.610 189.970 ;
        RECT 20.640 189.290 127.820 189.770 ;
        RECT 88.345 189.090 88.635 189.135 ;
        RECT 93.390 189.090 93.710 189.150 ;
        RECT 109.045 189.090 109.335 189.135 ;
        RECT 88.345 188.950 93.710 189.090 ;
        RECT 88.345 188.905 88.635 188.950 ;
        RECT 93.390 188.890 93.710 188.950 ;
        RECT 107.280 188.950 109.335 189.090 ;
        RECT 32.210 188.795 32.530 188.810 ;
        RECT 31.745 188.750 32.530 188.795 ;
        RECT 35.345 188.750 35.635 188.795 ;
        RECT 31.745 188.610 35.635 188.750 ;
        RECT 31.745 188.565 32.530 188.610 ;
        RECT 32.210 188.550 32.530 188.565 ;
        RECT 35.045 188.565 35.635 188.610 ;
        RECT 50.725 188.750 51.015 188.795 ;
        RECT 53.370 188.750 53.690 188.810 ;
        RECT 53.965 188.750 54.615 188.795 ;
        RECT 50.725 188.610 54.615 188.750 ;
        RECT 50.725 188.565 51.315 188.610 ;
        RECT 28.070 188.210 28.390 188.470 ;
        RECT 28.550 188.410 28.840 188.455 ;
        RECT 30.385 188.410 30.675 188.455 ;
        RECT 33.965 188.410 34.255 188.455 ;
        RECT 28.550 188.270 34.255 188.410 ;
        RECT 28.550 188.225 28.840 188.270 ;
        RECT 30.385 188.225 30.675 188.270 ;
        RECT 33.965 188.225 34.255 188.270 ;
        RECT 35.045 188.250 35.335 188.565 ;
        RECT 51.025 188.250 51.315 188.565 ;
        RECT 53.370 188.550 53.690 188.610 ;
        RECT 53.965 188.565 54.615 188.610 ;
        RECT 56.590 188.550 56.910 188.810 ;
        RECT 57.050 188.750 57.370 188.810 ;
        RECT 58.905 188.750 59.195 188.795 ;
        RECT 57.050 188.610 59.195 188.750 ;
        RECT 57.050 188.550 57.370 188.610 ;
        RECT 58.905 188.565 59.195 188.610 ;
        RECT 72.705 188.750 72.995 188.795 ;
        RECT 75.105 188.750 75.395 188.795 ;
        RECT 78.345 188.750 78.995 188.795 ;
        RECT 72.705 188.610 78.995 188.750 ;
        RECT 72.705 188.565 72.995 188.610 ;
        RECT 75.105 188.565 75.695 188.610 ;
        RECT 78.345 188.565 78.995 188.610 ;
        RECT 52.105 188.410 52.395 188.455 ;
        RECT 55.685 188.410 55.975 188.455 ;
        RECT 57.520 188.410 57.810 188.455 ;
        RECT 52.105 188.270 57.810 188.410 ;
        RECT 52.105 188.225 52.395 188.270 ;
        RECT 55.685 188.225 55.975 188.270 ;
        RECT 57.520 188.225 57.810 188.270 ;
        RECT 59.365 188.410 59.655 188.455 ;
        RECT 61.190 188.410 61.510 188.470 ;
        RECT 59.365 188.270 61.510 188.410 ;
        RECT 59.365 188.225 59.655 188.270 ;
        RECT 61.190 188.210 61.510 188.270 ;
        RECT 71.310 188.410 71.630 188.470 ;
        RECT 72.245 188.410 72.535 188.455 ;
        RECT 71.310 188.270 72.535 188.410 ;
        RECT 71.310 188.210 71.630 188.270 ;
        RECT 72.245 188.225 72.535 188.270 ;
        RECT 75.405 188.250 75.695 188.565 ;
        RECT 80.970 188.550 81.290 188.810 ;
        RECT 85.570 188.750 85.890 188.810 ;
        RECT 107.280 188.795 107.420 188.950 ;
        RECT 109.045 188.905 109.335 188.950 ;
        RECT 109.950 188.890 110.270 189.150 ;
        RECT 111.805 189.090 112.095 189.135 ;
        RECT 112.250 189.090 112.570 189.150 ;
        RECT 111.805 188.950 112.570 189.090 ;
        RECT 111.805 188.905 112.095 188.950 ;
        RECT 112.250 188.890 112.570 188.950 ;
        RECT 86.505 188.750 86.795 188.795 ;
        RECT 85.570 188.610 86.795 188.750 ;
        RECT 85.570 188.550 85.890 188.610 ;
        RECT 86.505 188.565 86.795 188.610 ;
        RECT 98.925 188.750 99.215 188.795 ;
        RECT 101.325 188.750 101.615 188.795 ;
        RECT 104.565 188.750 105.215 188.795 ;
        RECT 98.925 188.610 105.215 188.750 ;
        RECT 98.925 188.565 99.215 188.610 ;
        RECT 101.325 188.565 101.915 188.610 ;
        RECT 104.565 188.565 105.215 188.610 ;
        RECT 107.205 188.565 107.495 188.795 ;
        RECT 110.040 188.750 110.180 188.890 ;
        RECT 113.645 188.750 113.935 188.795 ;
        RECT 117.425 188.750 117.715 188.795 ;
        RECT 120.665 188.750 121.315 188.795 ;
        RECT 110.040 188.610 112.480 188.750 ;
        RECT 76.485 188.410 76.775 188.455 ;
        RECT 80.065 188.410 80.355 188.455 ;
        RECT 81.900 188.410 82.190 188.455 ;
        RECT 76.485 188.270 82.190 188.410 ;
        RECT 76.485 188.225 76.775 188.270 ;
        RECT 80.065 188.225 80.355 188.270 ;
        RECT 81.900 188.225 82.190 188.270 ;
        RECT 90.630 188.410 90.950 188.470 ;
        RECT 91.565 188.410 91.855 188.455 ;
        RECT 98.465 188.410 98.755 188.455 ;
        RECT 90.630 188.270 98.755 188.410 ;
        RECT 90.630 188.210 90.950 188.270 ;
        RECT 91.565 188.225 91.855 188.270 ;
        RECT 98.465 188.225 98.755 188.270 ;
        RECT 101.625 188.250 101.915 188.565 ;
        RECT 102.705 188.410 102.995 188.455 ;
        RECT 106.285 188.410 106.575 188.455 ;
        RECT 108.120 188.410 108.410 188.455 ;
        RECT 102.705 188.270 108.410 188.410 ;
        RECT 102.705 188.225 102.995 188.270 ;
        RECT 106.285 188.225 106.575 188.270 ;
        RECT 108.120 188.225 108.410 188.270 ;
        RECT 109.950 188.210 110.270 188.470 ;
        RECT 112.340 188.455 112.480 188.610 ;
        RECT 113.645 188.610 121.315 188.750 ;
        RECT 113.645 188.565 113.935 188.610 ;
        RECT 117.425 188.565 118.015 188.610 ;
        RECT 120.665 188.565 121.315 188.610 ;
        RECT 112.265 188.410 112.555 188.455 ;
        RECT 113.185 188.410 113.475 188.455 ;
        RECT 112.265 188.270 113.475 188.410 ;
        RECT 112.265 188.225 112.555 188.270 ;
        RECT 113.185 188.225 113.475 188.270 ;
        RECT 117.725 188.250 118.015 188.565 ;
        RECT 123.290 188.550 123.610 188.810 ;
        RECT 118.805 188.410 119.095 188.455 ;
        RECT 122.385 188.410 122.675 188.455 ;
        RECT 124.220 188.410 124.510 188.455 ;
        RECT 118.805 188.270 124.510 188.410 ;
        RECT 118.805 188.225 119.095 188.270 ;
        RECT 122.385 188.225 122.675 188.270 ;
        RECT 124.220 188.225 124.510 188.270 ;
        RECT 36.810 187.870 37.130 188.130 ;
        RECT 57.985 188.070 58.275 188.115 ;
        RECT 63.950 188.070 64.270 188.130 ;
        RECT 57.985 187.930 64.270 188.070 ;
        RECT 57.985 187.885 58.275 187.930 ;
        RECT 63.950 187.870 64.270 187.930 ;
        RECT 82.365 188.070 82.655 188.115 ;
        RECT 85.110 188.070 85.430 188.130 ;
        RECT 82.365 187.930 85.430 188.070 ;
        RECT 82.365 187.885 82.655 187.930 ;
        RECT 85.110 187.870 85.430 187.930 ;
        RECT 85.585 187.885 85.875 188.115 ;
        RECT 28.955 187.730 29.245 187.775 ;
        RECT 30.845 187.730 31.135 187.775 ;
        RECT 33.965 187.730 34.255 187.775 ;
        RECT 28.955 187.590 34.255 187.730 ;
        RECT 28.955 187.545 29.245 187.590 ;
        RECT 30.845 187.545 31.135 187.590 ;
        RECT 33.965 187.545 34.255 187.590 ;
        RECT 52.105 187.730 52.395 187.775 ;
        RECT 55.225 187.730 55.515 187.775 ;
        RECT 57.115 187.730 57.405 187.775 ;
        RECT 52.105 187.590 57.405 187.730 ;
        RECT 52.105 187.545 52.395 187.590 ;
        RECT 55.225 187.545 55.515 187.590 ;
        RECT 57.115 187.545 57.405 187.590 ;
        RECT 76.485 187.730 76.775 187.775 ;
        RECT 79.605 187.730 79.895 187.775 ;
        RECT 81.495 187.730 81.785 187.775 ;
        RECT 76.485 187.590 81.785 187.730 ;
        RECT 85.660 187.730 85.800 187.885 ;
        RECT 86.030 187.870 86.350 188.130 ;
        RECT 91.090 187.870 91.410 188.130 ;
        RECT 108.585 188.070 108.875 188.115 ;
        RECT 109.030 188.070 109.350 188.130 ;
        RECT 108.585 187.930 109.350 188.070 ;
        RECT 108.585 187.885 108.875 187.930 ;
        RECT 109.030 187.870 109.350 187.930 ;
        RECT 118.230 188.070 118.550 188.130 ;
        RECT 124.670 188.070 124.990 188.130 ;
        RECT 118.230 187.930 124.990 188.070 ;
        RECT 118.230 187.870 118.550 187.930 ;
        RECT 124.670 187.870 124.990 187.930 ;
        RECT 89.710 187.730 90.030 187.790 ;
        RECT 91.550 187.730 91.870 187.790 ;
        RECT 85.660 187.590 91.870 187.730 ;
        RECT 76.485 187.545 76.775 187.590 ;
        RECT 79.605 187.545 79.895 187.590 ;
        RECT 81.495 187.545 81.785 187.590 ;
        RECT 89.710 187.530 90.030 187.590 ;
        RECT 91.550 187.530 91.870 187.590 ;
        RECT 102.705 187.730 102.995 187.775 ;
        RECT 105.825 187.730 106.115 187.775 ;
        RECT 107.715 187.730 108.005 187.775 ;
        RECT 102.705 187.590 108.005 187.730 ;
        RECT 102.705 187.545 102.995 187.590 ;
        RECT 105.825 187.545 106.115 187.590 ;
        RECT 107.715 187.545 108.005 187.590 ;
        RECT 118.805 187.730 119.095 187.775 ;
        RECT 121.925 187.730 122.215 187.775 ;
        RECT 123.815 187.730 124.105 187.775 ;
        RECT 118.805 187.590 124.105 187.730 ;
        RECT 118.805 187.545 119.095 187.590 ;
        RECT 121.925 187.545 122.215 187.590 ;
        RECT 123.815 187.545 124.105 187.590 ;
        RECT 29.450 187.435 29.770 187.450 ;
        RECT 29.405 187.205 29.770 187.435 ;
        RECT 29.450 187.190 29.770 187.205 ;
        RECT 46.470 187.390 46.790 187.450 ;
        RECT 49.245 187.390 49.535 187.435 ;
        RECT 46.470 187.250 49.535 187.390 ;
        RECT 46.470 187.190 46.790 187.250 ;
        RECT 49.245 187.205 49.535 187.250 ;
        RECT 73.150 187.390 73.470 187.450 ;
        RECT 73.625 187.390 73.915 187.435 ;
        RECT 73.150 187.250 73.915 187.390 ;
        RECT 73.150 187.190 73.470 187.250 ;
        RECT 73.625 187.205 73.915 187.250 ;
        RECT 98.910 187.390 99.230 187.450 ;
        RECT 99.845 187.390 100.135 187.435 ;
        RECT 98.910 187.250 100.135 187.390 ;
        RECT 98.910 187.190 99.230 187.250 ;
        RECT 99.845 187.205 100.135 187.250 ;
        RECT 115.470 187.390 115.790 187.450 ;
        RECT 115.945 187.390 116.235 187.435 ;
        RECT 115.470 187.250 116.235 187.390 ;
        RECT 115.470 187.190 115.790 187.250 ;
        RECT 115.945 187.205 116.235 187.250 ;
        RECT 20.640 186.570 127.820 187.050 ;
        RECT 54.750 186.170 55.070 186.430 ;
        RECT 107.665 186.370 107.955 186.415 ;
        RECT 109.950 186.370 110.270 186.430 ;
        RECT 107.665 186.230 110.270 186.370 ;
        RECT 107.665 186.185 107.955 186.230 ;
        RECT 109.950 186.170 110.270 186.230 ;
        RECT 111.420 186.230 116.160 186.370 ;
        RECT 29.450 186.030 29.770 186.090 ;
        RECT 33.145 186.030 33.435 186.075 ;
        RECT 29.450 185.890 33.435 186.030 ;
        RECT 29.450 185.830 29.770 185.890 ;
        RECT 33.145 185.845 33.435 185.890 ;
        RECT 58.085 186.030 58.375 186.075 ;
        RECT 61.205 186.030 61.495 186.075 ;
        RECT 63.095 186.030 63.385 186.075 ;
        RECT 76.385 186.030 76.675 186.075 ;
        RECT 58.085 185.890 63.385 186.030 ;
        RECT 58.085 185.845 58.375 185.890 ;
        RECT 61.205 185.845 61.495 185.890 ;
        RECT 63.095 185.845 63.385 185.890 ;
        RECT 73.700 185.890 76.675 186.030 ;
        RECT 37.745 185.690 38.035 185.735 ;
        RECT 43.250 185.690 43.570 185.750 ;
        RECT 46.945 185.690 47.235 185.735 ;
        RECT 51.990 185.690 52.310 185.750 ;
        RECT 73.150 185.735 73.470 185.750 ;
        RECT 73.700 185.735 73.840 185.890 ;
        RECT 76.385 185.845 76.675 185.890 ;
        RECT 79.245 186.030 79.535 186.075 ;
        RECT 82.365 186.030 82.655 186.075 ;
        RECT 84.255 186.030 84.545 186.075 ;
        RECT 79.245 185.890 84.545 186.030 ;
        RECT 79.245 185.845 79.535 185.890 ;
        RECT 82.365 185.845 82.655 185.890 ;
        RECT 84.255 185.845 84.545 185.890 ;
        RECT 90.285 186.030 90.575 186.075 ;
        RECT 93.405 186.030 93.695 186.075 ;
        RECT 95.295 186.030 95.585 186.075 ;
        RECT 90.285 185.890 95.585 186.030 ;
        RECT 90.285 185.845 90.575 185.890 ;
        RECT 93.405 185.845 93.695 185.890 ;
        RECT 95.295 185.845 95.585 185.890 ;
        RECT 73.040 185.690 73.470 185.735 ;
        RECT 33.680 185.550 36.120 185.690 ;
        RECT 31.290 185.350 31.610 185.410 ;
        RECT 33.680 185.350 33.820 185.550 ;
        RECT 35.980 185.410 36.120 185.550 ;
        RECT 37.745 185.550 52.310 185.690 ;
        RECT 37.745 185.505 38.035 185.550 ;
        RECT 43.250 185.490 43.570 185.550 ;
        RECT 46.945 185.505 47.235 185.550 ;
        RECT 51.990 185.490 52.310 185.550 ;
        RECT 71.170 185.550 73.470 185.690 ;
        RECT 31.290 185.210 33.820 185.350 ;
        RECT 34.065 185.350 34.355 185.395 ;
        RECT 35.890 185.350 36.210 185.410 ;
        RECT 44.645 185.350 44.935 185.395 ;
        RECT 57.050 185.370 57.370 185.410 ;
        RECT 34.065 185.210 34.740 185.350 ;
        RECT 31.290 185.150 31.610 185.210 ;
        RECT 34.065 185.165 34.355 185.210 ;
        RECT 31.750 184.470 32.070 184.730 ;
        RECT 34.600 184.715 34.740 185.210 ;
        RECT 35.890 185.210 44.935 185.350 ;
        RECT 35.890 185.150 36.210 185.210 ;
        RECT 44.645 185.165 44.935 185.210 ;
        RECT 57.005 185.150 57.370 185.370 ;
        RECT 58.085 185.350 58.375 185.395 ;
        RECT 61.665 185.350 61.955 185.395 ;
        RECT 63.500 185.350 63.790 185.395 ;
        RECT 58.085 185.210 63.790 185.350 ;
        RECT 58.085 185.165 58.375 185.210 ;
        RECT 61.665 185.165 61.955 185.210 ;
        RECT 63.500 185.165 63.790 185.210 ;
        RECT 63.950 185.150 64.270 185.410 ;
        RECT 69.025 185.350 69.315 185.395 ;
        RECT 71.170 185.350 71.310 185.550 ;
        RECT 73.040 185.505 73.470 185.550 ;
        RECT 73.625 185.505 73.915 185.735 ;
        RECT 74.085 185.690 74.375 185.735 ;
        RECT 74.990 185.690 75.310 185.750 ;
        RECT 74.085 185.550 75.310 185.690 ;
        RECT 74.085 185.505 74.375 185.550 ;
        RECT 73.150 185.490 73.470 185.505 ;
        RECT 69.025 185.210 71.310 185.350 ;
        RECT 71.785 185.350 72.075 185.395 ;
        RECT 73.700 185.350 73.840 185.505 ;
        RECT 74.990 185.490 75.310 185.550 ;
        RECT 85.110 185.690 85.430 185.750 ;
        RECT 88.790 185.690 89.110 185.750 ;
        RECT 85.110 185.550 89.110 185.690 ;
        RECT 85.110 185.490 85.430 185.550 ;
        RECT 88.790 185.490 89.110 185.550 ;
        RECT 89.710 185.690 90.030 185.750 ;
        RECT 97.545 185.690 97.835 185.735 ;
        RECT 104.445 185.690 104.735 185.735 ;
        RECT 106.270 185.690 106.590 185.750 ;
        RECT 111.420 185.690 111.560 186.230 ;
        RECT 111.790 186.030 112.110 186.090 ;
        RECT 111.790 185.890 114.320 186.030 ;
        RECT 111.790 185.830 112.110 185.890 ;
        RECT 112.265 185.690 112.555 185.735 ;
        RECT 89.710 185.550 112.555 185.690 ;
        RECT 89.710 185.490 90.030 185.550 ;
        RECT 97.545 185.505 97.835 185.550 ;
        RECT 104.445 185.505 104.735 185.550 ;
        RECT 106.270 185.490 106.590 185.550 ;
        RECT 112.265 185.505 112.555 185.550 ;
        RECT 71.785 185.210 73.840 185.350 ;
        RECT 69.025 185.165 69.315 185.210 ;
        RECT 71.785 185.165 72.075 185.210 ;
        RECT 36.365 185.010 36.655 185.055 ;
        RECT 37.270 185.010 37.590 185.070 ;
        RECT 36.365 184.870 37.590 185.010 ;
        RECT 36.365 184.825 36.655 184.870 ;
        RECT 37.270 184.810 37.590 184.870 ;
        RECT 40.490 185.010 40.810 185.070 ;
        RECT 57.005 185.055 57.295 185.150 ;
        RECT 72.780 185.070 72.920 185.210 ;
        RECT 75.465 185.165 75.755 185.395 ;
        RECT 47.405 185.010 47.695 185.055 ;
        RECT 52.465 185.010 52.755 185.055 ;
        RECT 40.490 184.870 47.695 185.010 ;
        RECT 40.490 184.810 40.810 184.870 ;
        RECT 47.405 184.825 47.695 184.870 ;
        RECT 47.940 184.870 52.755 185.010 ;
        RECT 34.525 184.485 34.815 184.715 ;
        RECT 36.810 184.670 37.130 184.730 ;
        RECT 38.650 184.670 38.970 184.730 ;
        RECT 36.810 184.530 38.970 184.670 ;
        RECT 36.810 184.470 37.130 184.530 ;
        RECT 38.650 184.470 38.970 184.530 ;
        RECT 44.170 184.470 44.490 184.730 ;
        RECT 46.470 184.670 46.790 184.730 ;
        RECT 47.940 184.715 48.080 184.870 ;
        RECT 52.465 184.825 52.755 184.870 ;
        RECT 56.705 185.010 57.295 185.055 ;
        RECT 59.945 185.010 60.595 185.055 ;
        RECT 56.705 184.870 60.595 185.010 ;
        RECT 56.705 184.825 56.995 184.870 ;
        RECT 59.945 184.825 60.595 184.870 ;
        RECT 62.570 184.810 62.890 185.070 ;
        RECT 72.690 184.810 73.010 185.070 ;
        RECT 73.610 185.010 73.930 185.070 ;
        RECT 75.540 185.010 75.680 185.165 ;
        RECT 73.610 184.870 75.680 185.010 ;
        RECT 76.370 185.010 76.690 185.070 ;
        RECT 78.165 185.055 78.455 185.370 ;
        RECT 79.245 185.350 79.535 185.395 ;
        RECT 82.825 185.350 83.115 185.395 ;
        RECT 84.660 185.350 84.950 185.395 ;
        RECT 79.245 185.210 84.950 185.350 ;
        RECT 79.245 185.165 79.535 185.210 ;
        RECT 82.825 185.165 83.115 185.210 ;
        RECT 84.660 185.165 84.950 185.210 ;
        RECT 77.865 185.010 78.455 185.055 ;
        RECT 81.105 185.010 81.755 185.055 ;
        RECT 76.370 184.870 81.755 185.010 ;
        RECT 73.610 184.810 73.930 184.870 ;
        RECT 76.370 184.810 76.690 184.870 ;
        RECT 77.865 184.825 78.155 184.870 ;
        RECT 81.105 184.825 81.755 184.870 ;
        RECT 83.730 184.810 84.050 185.070 ;
        RECT 89.205 185.055 89.495 185.370 ;
        RECT 90.285 185.350 90.575 185.395 ;
        RECT 93.865 185.350 94.155 185.395 ;
        RECT 95.700 185.350 95.990 185.395 ;
        RECT 90.285 185.210 95.990 185.350 ;
        RECT 90.285 185.165 90.575 185.210 ;
        RECT 93.865 185.165 94.155 185.210 ;
        RECT 95.700 185.165 95.990 185.210 ;
        RECT 96.150 185.150 96.470 185.410 ;
        RECT 105.810 185.350 106.130 185.410 ;
        RECT 109.490 185.350 109.810 185.410 ;
        RECT 112.725 185.350 113.015 185.395 ;
        RECT 105.810 185.210 113.015 185.350 ;
        RECT 114.180 185.350 114.320 185.890 ;
        RECT 116.020 185.735 116.160 186.230 ;
        RECT 119.150 186.170 119.470 186.430 ;
        RECT 115.945 185.505 116.235 185.735 ;
        RECT 117.325 185.350 117.615 185.395 ;
        RECT 114.180 185.210 117.615 185.350 ;
        RECT 105.810 185.150 106.130 185.210 ;
        RECT 109.490 185.150 109.810 185.210 ;
        RECT 112.725 185.165 113.015 185.210 ;
        RECT 117.325 185.165 117.615 185.210 ;
        RECT 88.905 185.010 89.495 185.055 ;
        RECT 91.090 185.010 91.410 185.070 ;
        RECT 92.145 185.010 92.795 185.055 ;
        RECT 88.905 184.870 92.795 185.010 ;
        RECT 88.905 184.825 89.195 184.870 ;
        RECT 91.090 184.810 91.410 184.870 ;
        RECT 92.145 184.825 92.795 184.870 ;
        RECT 94.310 185.010 94.630 185.070 ;
        RECT 94.785 185.010 95.075 185.055 ;
        RECT 105.365 185.010 105.655 185.055 ;
        RECT 115.470 185.010 115.790 185.070 ;
        RECT 116.865 185.010 117.155 185.055 ;
        RECT 94.310 184.870 95.075 185.010 ;
        RECT 94.310 184.810 94.630 184.870 ;
        RECT 94.785 184.825 95.075 184.870 ;
        RECT 99.000 184.870 105.655 185.010 ;
        RECT 99.000 184.730 99.140 184.870 ;
        RECT 105.365 184.825 105.655 184.870 ;
        RECT 113.260 184.870 117.155 185.010 ;
        RECT 113.260 184.730 113.400 184.870 ;
        RECT 115.470 184.810 115.790 184.870 ;
        RECT 116.865 184.825 117.155 184.870 ;
        RECT 47.865 184.670 48.155 184.715 ;
        RECT 46.470 184.530 48.155 184.670 ;
        RECT 46.470 184.470 46.790 184.530 ;
        RECT 47.865 184.485 48.155 184.530 ;
        RECT 49.690 184.470 50.010 184.730 ;
        RECT 52.925 184.670 53.215 184.715 ;
        RECT 54.290 184.670 54.610 184.730 ;
        RECT 55.225 184.670 55.515 184.715 ;
        RECT 52.925 184.530 55.515 184.670 ;
        RECT 52.925 184.485 53.215 184.530 ;
        RECT 54.290 184.470 54.610 184.530 ;
        RECT 55.225 184.485 55.515 184.530 ;
        RECT 69.470 184.470 69.790 184.730 ;
        RECT 70.390 184.670 70.710 184.730 ;
        RECT 70.865 184.670 71.155 184.715 ;
        RECT 70.390 184.530 71.155 184.670 ;
        RECT 70.390 184.470 70.710 184.530 ;
        RECT 70.865 184.485 71.155 184.530 ;
        RECT 72.245 184.670 72.535 184.715 ;
        RECT 74.070 184.670 74.390 184.730 ;
        RECT 72.245 184.530 74.390 184.670 ;
        RECT 72.245 184.485 72.535 184.530 ;
        RECT 74.070 184.470 74.390 184.530 ;
        RECT 85.570 184.670 85.890 184.730 ;
        RECT 87.425 184.670 87.715 184.715 ;
        RECT 85.570 184.530 87.715 184.670 ;
        RECT 85.570 184.470 85.890 184.530 ;
        RECT 87.425 184.485 87.715 184.530 ;
        RECT 93.850 184.670 94.170 184.730 ;
        RECT 98.465 184.670 98.755 184.715 ;
        RECT 93.850 184.530 98.755 184.670 ;
        RECT 93.850 184.470 94.170 184.530 ;
        RECT 98.465 184.485 98.755 184.530 ;
        RECT 98.910 184.470 99.230 184.730 ;
        RECT 100.290 184.670 100.610 184.730 ;
        RECT 100.765 184.670 101.055 184.715 ;
        RECT 100.290 184.530 101.055 184.670 ;
        RECT 100.290 184.470 100.610 184.530 ;
        RECT 100.765 184.485 101.055 184.530 ;
        RECT 113.170 184.470 113.490 184.730 ;
        RECT 115.010 184.470 115.330 184.730 ;
        RECT 20.640 183.850 127.820 184.330 ;
        RECT 40.490 183.450 40.810 183.710 ;
        RECT 49.705 183.650 49.995 183.695 ;
        RECT 47.940 183.510 49.995 183.650 ;
        RECT 31.750 183.355 32.070 183.370 ;
        RECT 31.745 183.310 32.395 183.355 ;
        RECT 35.345 183.310 35.635 183.355 ;
        RECT 31.745 183.170 35.635 183.310 ;
        RECT 31.745 183.125 32.395 183.170 ;
        RECT 35.045 183.125 35.635 183.170 ;
        RECT 41.985 183.310 42.275 183.355 ;
        RECT 44.170 183.310 44.490 183.370 ;
        RECT 47.940 183.355 48.080 183.510 ;
        RECT 49.705 183.465 49.995 183.510 ;
        RECT 61.665 183.650 61.955 183.695 ;
        RECT 62.570 183.650 62.890 183.710 ;
        RECT 61.665 183.510 62.890 183.650 ;
        RECT 61.665 183.465 61.955 183.510 ;
        RECT 62.570 183.450 62.890 183.510 ;
        RECT 72.690 183.450 73.010 183.710 ;
        RECT 73.150 183.450 73.470 183.710 ;
        RECT 76.370 183.650 76.690 183.710 ;
        RECT 77.305 183.650 77.595 183.695 ;
        RECT 76.370 183.510 77.595 183.650 ;
        RECT 76.370 183.450 76.690 183.510 ;
        RECT 77.305 183.465 77.595 183.510 ;
        RECT 79.605 183.650 79.895 183.695 ;
        RECT 83.730 183.650 84.050 183.710 ;
        RECT 79.605 183.510 84.050 183.650 ;
        RECT 79.605 183.465 79.895 183.510 ;
        RECT 83.730 183.450 84.050 183.510 ;
        RECT 84.190 183.650 84.510 183.710 ;
        RECT 91.565 183.650 91.855 183.695 ;
        RECT 93.850 183.650 94.170 183.710 ;
        RECT 84.190 183.510 94.170 183.650 ;
        RECT 84.190 183.450 84.510 183.510 ;
        RECT 91.565 183.465 91.855 183.510 ;
        RECT 93.850 183.450 94.170 183.510 ;
        RECT 115.930 183.450 116.250 183.710 ;
        RECT 45.225 183.310 45.875 183.355 ;
        RECT 41.985 183.170 45.875 183.310 ;
        RECT 41.985 183.125 42.575 183.170 ;
        RECT 31.750 183.110 32.070 183.125 ;
        RECT 28.070 182.770 28.390 183.030 ;
        RECT 28.550 182.970 28.840 183.015 ;
        RECT 30.385 182.970 30.675 183.015 ;
        RECT 33.965 182.970 34.255 183.015 ;
        RECT 28.550 182.830 34.255 182.970 ;
        RECT 28.550 182.785 28.840 182.830 ;
        RECT 30.385 182.785 30.675 182.830 ;
        RECT 33.965 182.785 34.255 182.830 ;
        RECT 35.045 182.810 35.335 183.125 ;
        RECT 42.285 182.810 42.575 183.125 ;
        RECT 44.170 183.110 44.490 183.170 ;
        RECT 45.225 183.125 45.875 183.170 ;
        RECT 47.865 183.125 48.155 183.355 ;
        RECT 73.610 183.310 73.930 183.370 ;
        RECT 74.990 183.310 75.310 183.370 ;
        RECT 75.465 183.310 75.755 183.355 ;
        RECT 85.585 183.310 85.875 183.355 ;
        RECT 73.610 183.170 75.755 183.310 ;
        RECT 73.610 183.110 73.930 183.170 ;
        RECT 74.990 183.110 75.310 183.170 ;
        RECT 75.465 183.125 75.755 183.170 ;
        RECT 76.920 183.170 85.875 183.310 ;
        RECT 43.365 182.970 43.655 183.015 ;
        RECT 46.945 182.970 47.235 183.015 ;
        RECT 48.780 182.970 49.070 183.015 ;
        RECT 43.365 182.830 49.070 182.970 ;
        RECT 43.365 182.785 43.655 182.830 ;
        RECT 46.945 182.785 47.235 182.830 ;
        RECT 48.780 182.785 49.070 182.830 ;
        RECT 49.230 182.770 49.550 183.030 ;
        RECT 49.690 182.970 50.010 183.030 ;
        RECT 50.625 182.970 50.915 183.015 ;
        RECT 49.690 182.830 50.915 182.970 ;
        RECT 49.690 182.770 50.010 182.830 ;
        RECT 50.625 182.785 50.915 182.830 ;
        RECT 56.590 182.970 56.910 183.030 ;
        RECT 60.745 182.970 61.035 183.015 ;
        RECT 56.590 182.830 61.035 182.970 ;
        RECT 56.590 182.770 56.910 182.830 ;
        RECT 60.745 182.785 61.035 182.830 ;
        RECT 71.310 182.970 71.630 183.030 ;
        RECT 76.920 183.015 77.060 183.170 ;
        RECT 85.585 183.125 85.875 183.170 ;
        RECT 95.345 183.310 95.635 183.355 ;
        RECT 97.530 183.310 97.850 183.370 ;
        RECT 98.585 183.310 99.235 183.355 ;
        RECT 95.345 183.170 99.235 183.310 ;
        RECT 95.345 183.125 95.935 183.170 ;
        RECT 76.845 182.970 77.135 183.015 ;
        RECT 71.310 182.830 77.135 182.970 ;
        RECT 71.310 182.770 71.630 182.830 ;
        RECT 76.845 182.785 77.135 182.830 ;
        RECT 79.130 182.770 79.450 183.030 ;
        RECT 84.205 182.785 84.495 183.015 ;
        RECT 91.105 182.970 91.395 183.015 ;
        RECT 85.660 182.830 91.395 182.970 ;
        RECT 29.450 182.430 29.770 182.690 ;
        RECT 28.955 182.290 29.245 182.335 ;
        RECT 30.845 182.290 31.135 182.335 ;
        RECT 33.965 182.290 34.255 182.335 ;
        RECT 28.955 182.150 34.255 182.290 ;
        RECT 28.955 182.105 29.245 182.150 ;
        RECT 30.845 182.105 31.135 182.150 ;
        RECT 33.965 182.105 34.255 182.150 ;
        RECT 43.365 182.290 43.655 182.335 ;
        RECT 46.485 182.290 46.775 182.335 ;
        RECT 48.375 182.290 48.665 182.335 ;
        RECT 43.365 182.150 48.665 182.290 ;
        RECT 43.365 182.105 43.655 182.150 ;
        RECT 46.485 182.105 46.775 182.150 ;
        RECT 48.375 182.105 48.665 182.150 ;
        RECT 74.530 182.290 74.850 182.350 ;
        RECT 75.465 182.290 75.755 182.335 ;
        RECT 74.530 182.150 75.755 182.290 ;
        RECT 74.530 182.090 74.850 182.150 ;
        RECT 75.465 182.105 75.755 182.150 ;
        RECT 76.370 182.290 76.690 182.350 ;
        RECT 84.280 182.290 84.420 182.785 ;
        RECT 85.660 182.690 85.800 182.830 ;
        RECT 91.105 182.785 91.395 182.830 ;
        RECT 95.645 182.810 95.935 183.125 ;
        RECT 97.530 183.110 97.850 183.170 ;
        RECT 98.585 183.125 99.235 183.170 ;
        RECT 101.210 183.110 101.530 183.370 ;
        RECT 112.710 183.310 113.030 183.370 ;
        RECT 111.420 183.170 113.030 183.310 ;
        RECT 96.725 182.970 97.015 183.015 ;
        RECT 100.305 182.970 100.595 183.015 ;
        RECT 102.140 182.970 102.430 183.015 ;
        RECT 96.725 182.830 102.430 182.970 ;
        RECT 96.725 182.785 97.015 182.830 ;
        RECT 100.305 182.785 100.595 182.830 ;
        RECT 102.140 182.785 102.430 182.830 ;
        RECT 106.270 182.970 106.590 183.030 ;
        RECT 109.950 182.970 110.270 183.030 ;
        RECT 111.420 183.015 111.560 183.170 ;
        RECT 112.710 183.110 113.030 183.170 ;
        RECT 111.345 182.970 111.635 183.015 ;
        RECT 106.270 182.830 111.635 182.970 ;
        RECT 106.270 182.770 106.590 182.830 ;
        RECT 109.950 182.770 110.270 182.830 ;
        RECT 111.345 182.785 111.635 182.830 ;
        RECT 111.790 182.770 112.110 183.030 ;
        RECT 112.250 182.770 112.570 183.030 ;
        RECT 113.185 182.785 113.475 183.015 ;
        RECT 85.570 182.430 85.890 182.690 ;
        RECT 89.710 182.630 90.030 182.690 ;
        RECT 90.185 182.630 90.475 182.675 ;
        RECT 96.150 182.630 96.470 182.690 ;
        RECT 102.605 182.630 102.895 182.675 ;
        RECT 89.710 182.490 90.475 182.630 ;
        RECT 89.710 182.430 90.030 182.490 ;
        RECT 90.185 182.445 90.475 182.490 ;
        RECT 92.560 182.490 102.895 182.630 ;
        RECT 86.950 182.290 87.270 182.350 ;
        RECT 76.370 182.150 87.270 182.290 ;
        RECT 76.370 182.090 76.690 182.150 ;
        RECT 86.950 182.090 87.270 182.150 ;
        RECT 89.250 182.290 89.570 182.350 ;
        RECT 92.560 182.290 92.700 182.490 ;
        RECT 96.150 182.430 96.470 182.490 ;
        RECT 102.605 182.445 102.895 182.490 ;
        RECT 110.870 182.630 111.190 182.690 ;
        RECT 113.260 182.630 113.400 182.785 ;
        RECT 115.010 182.770 115.330 183.030 ;
        RECT 110.870 182.490 113.400 182.630 ;
        RECT 110.870 182.430 111.190 182.490 ;
        RECT 89.250 182.150 92.700 182.290 ;
        RECT 96.725 182.290 97.015 182.335 ;
        RECT 99.845 182.290 100.135 182.335 ;
        RECT 101.735 182.290 102.025 182.335 ;
        RECT 96.725 182.150 102.025 182.290 ;
        RECT 89.250 182.090 89.570 182.150 ;
        RECT 96.725 182.105 97.015 182.150 ;
        RECT 99.845 182.105 100.135 182.150 ;
        RECT 101.735 182.105 102.025 182.150 ;
        RECT 36.825 181.950 37.115 181.995 ;
        RECT 37.270 181.950 37.590 182.010 ;
        RECT 40.950 181.950 41.270 182.010 ;
        RECT 36.825 181.810 41.270 181.950 ;
        RECT 36.825 181.765 37.115 181.810 ;
        RECT 37.270 181.750 37.590 181.810 ;
        RECT 40.950 181.750 41.270 181.810 ;
        RECT 71.785 181.950 72.075 181.995 ;
        RECT 72.690 181.950 73.010 182.010 ;
        RECT 71.785 181.810 73.010 181.950 ;
        RECT 71.785 181.765 72.075 181.810 ;
        RECT 72.690 181.750 73.010 181.810 ;
        RECT 93.405 181.950 93.695 181.995 ;
        RECT 93.850 181.950 94.170 182.010 ;
        RECT 93.405 181.810 94.170 181.950 ;
        RECT 93.405 181.765 93.695 181.810 ;
        RECT 93.850 181.750 94.170 181.810 ;
        RECT 109.965 181.950 110.255 181.995 ;
        RECT 112.250 181.950 112.570 182.010 ;
        RECT 109.965 181.810 112.570 181.950 ;
        RECT 109.965 181.765 110.255 181.810 ;
        RECT 112.250 181.750 112.570 181.810 ;
        RECT 20.640 181.130 127.820 181.610 ;
        RECT 51.990 180.930 52.310 180.990 ;
        RECT 43.340 180.790 52.310 180.930 ;
        RECT 29.450 180.590 29.770 180.650 ;
        RECT 35.445 180.590 35.735 180.635 ;
        RECT 29.450 180.450 35.735 180.590 ;
        RECT 29.450 180.390 29.770 180.450 ;
        RECT 35.445 180.405 35.735 180.450 ;
        RECT 40.045 180.250 40.335 180.295 ;
        RECT 43.340 180.250 43.480 180.790 ;
        RECT 51.990 180.730 52.310 180.790 ;
        RECT 56.590 180.730 56.910 180.990 ;
        RECT 70.405 180.930 70.695 180.975 ;
        RECT 81.430 180.930 81.750 180.990 ;
        RECT 64.500 180.790 81.750 180.930 ;
        RECT 51.530 180.590 51.850 180.650 ;
        RECT 64.500 180.590 64.640 180.790 ;
        RECT 70.405 180.745 70.695 180.790 ;
        RECT 81.430 180.730 81.750 180.790 ;
        RECT 82.365 180.930 82.655 180.975 ;
        RECT 89.710 180.930 90.030 180.990 ;
        RECT 82.365 180.790 90.030 180.930 ;
        RECT 82.365 180.745 82.655 180.790 ;
        RECT 89.710 180.730 90.030 180.790 ;
        RECT 94.310 180.730 94.630 180.990 ;
        RECT 101.210 180.730 101.530 180.990 ;
        RECT 51.530 180.450 64.640 180.590 ;
        RECT 51.530 180.390 51.850 180.450 ;
        RECT 68.105 180.405 68.395 180.635 ;
        RECT 96.610 180.590 96.930 180.650 ;
        RECT 81.060 180.450 96.930 180.590 ;
        RECT 40.045 180.110 43.480 180.250 ;
        RECT 46.470 180.250 46.790 180.310 ;
        RECT 51.990 180.250 52.310 180.310 ;
        RECT 53.845 180.250 54.135 180.295 ;
        RECT 57.985 180.250 58.275 180.295 ;
        RECT 61.665 180.250 61.955 180.295 ;
        RECT 46.470 180.110 49.000 180.250 ;
        RECT 40.045 180.065 40.335 180.110 ;
        RECT 46.470 180.050 46.790 180.110 ;
        RECT 36.365 179.910 36.655 179.955 ;
        RECT 38.665 179.910 38.955 179.955 ;
        RECT 40.490 179.910 40.810 179.970 ;
        RECT 36.365 179.770 37.040 179.910 ;
        RECT 36.365 179.725 36.655 179.770 ;
        RECT 36.900 179.275 37.040 179.770 ;
        RECT 38.665 179.770 40.810 179.910 ;
        RECT 38.665 179.725 38.955 179.770 ;
        RECT 40.490 179.710 40.810 179.770 ;
        RECT 45.090 179.910 45.410 179.970 ;
        RECT 47.865 179.910 48.155 179.955 ;
        RECT 45.090 179.770 48.155 179.910 ;
        RECT 45.090 179.710 45.410 179.770 ;
        RECT 47.865 179.725 48.155 179.770 ;
        RECT 48.310 179.710 48.630 179.970 ;
        RECT 48.860 179.955 49.000 180.110 ;
        RECT 51.990 180.110 61.955 180.250 ;
        RECT 51.990 180.050 52.310 180.110 ;
        RECT 53.845 180.065 54.135 180.110 ;
        RECT 57.985 180.065 58.275 180.110 ;
        RECT 61.665 180.065 61.955 180.110 ;
        RECT 68.180 180.250 68.320 180.405 ;
        RECT 81.060 180.250 81.200 180.450 ;
        RECT 96.610 180.390 96.930 180.450 ;
        RECT 97.085 180.590 97.375 180.635 ;
        RECT 97.530 180.590 97.850 180.650 ;
        RECT 120.185 180.590 120.475 180.635 ;
        RECT 123.305 180.590 123.595 180.635 ;
        RECT 125.195 180.590 125.485 180.635 ;
        RECT 97.085 180.450 97.850 180.590 ;
        RECT 97.085 180.405 97.375 180.450 ;
        RECT 97.530 180.390 97.850 180.450 ;
        RECT 104.060 180.450 116.160 180.590 ;
        RECT 68.180 180.110 81.200 180.250 ;
        RECT 81.430 180.250 81.750 180.310 ;
        RECT 96.700 180.250 96.840 180.390 ;
        RECT 103.510 180.250 103.830 180.310 ;
        RECT 81.430 180.110 85.340 180.250 ;
        RECT 96.700 180.110 103.830 180.250 ;
        RECT 48.785 179.725 49.075 179.955 ;
        RECT 49.705 179.910 49.995 179.955 ;
        RECT 50.150 179.910 50.470 179.970 ;
        RECT 68.180 179.910 68.320 180.110 ;
        RECT 81.430 180.050 81.750 180.110 ;
        RECT 49.705 179.770 50.470 179.910 ;
        RECT 49.705 179.725 49.995 179.770 ;
        RECT 50.150 179.710 50.470 179.770 ;
        RECT 50.700 179.770 68.320 179.910 ;
        RECT 69.025 179.910 69.315 179.955 ;
        RECT 69.485 179.910 69.775 179.955 ;
        RECT 71.310 179.910 71.630 179.970 ;
        RECT 69.025 179.770 71.630 179.910 ;
        RECT 44.630 179.570 44.950 179.630 ;
        RECT 50.700 179.570 50.840 179.770 ;
        RECT 69.025 179.725 69.315 179.770 ;
        RECT 69.485 179.725 69.775 179.770 ;
        RECT 71.310 179.710 71.630 179.770 ;
        RECT 80.510 179.910 80.830 179.970 ;
        RECT 85.200 179.955 85.340 180.110 ;
        RECT 103.510 180.050 103.830 180.110 ;
        RECT 84.665 179.910 84.955 179.955 ;
        RECT 80.510 179.770 84.955 179.910 ;
        RECT 80.510 179.710 80.830 179.770 ;
        RECT 84.665 179.725 84.955 179.770 ;
        RECT 85.125 179.725 85.415 179.955 ;
        RECT 85.570 179.710 85.890 179.970 ;
        RECT 86.490 179.710 86.810 179.970 ;
        RECT 93.405 179.910 93.695 179.955 ;
        RECT 93.850 179.910 94.170 179.970 ;
        RECT 93.405 179.770 94.170 179.910 ;
        RECT 93.405 179.725 93.695 179.770 ;
        RECT 93.850 179.710 94.170 179.770 ;
        RECT 97.545 179.725 97.835 179.955 ;
        RECT 44.630 179.430 50.840 179.570 ;
        RECT 44.630 179.370 44.950 179.430 ;
        RECT 54.290 179.370 54.610 179.630 ;
        RECT 56.130 179.570 56.450 179.630 ;
        RECT 58.905 179.570 59.195 179.615 ;
        RECT 59.810 179.570 60.130 179.630 ;
        RECT 56.130 179.430 60.130 179.570 ;
        RECT 56.130 179.370 56.450 179.430 ;
        RECT 58.905 179.385 59.195 179.430 ;
        RECT 59.810 179.370 60.130 179.430 ;
        RECT 63.045 179.570 63.335 179.615 ;
        RECT 73.610 179.570 73.930 179.630 ;
        RECT 80.985 179.570 81.275 179.615 ;
        RECT 63.045 179.430 81.275 179.570 ;
        RECT 63.045 179.385 63.335 179.430 ;
        RECT 73.610 179.370 73.930 179.430 ;
        RECT 80.985 179.385 81.275 179.430 ;
        RECT 90.630 179.570 90.950 179.630 ;
        RECT 97.620 179.570 97.760 179.725 ;
        RECT 100.290 179.710 100.610 179.970 ;
        RECT 103.065 179.910 103.355 179.955 ;
        RECT 104.060 179.910 104.200 180.450 ;
        RECT 113.170 180.250 113.490 180.310 ;
        RECT 111.420 180.110 113.490 180.250 ;
        RECT 103.065 179.770 104.200 179.910 ;
        RECT 106.270 179.910 106.590 179.970 ;
        RECT 108.125 179.910 108.415 179.955 ;
        RECT 106.270 179.770 108.415 179.910 ;
        RECT 103.065 179.725 103.355 179.770 ;
        RECT 103.140 179.570 103.280 179.725 ;
        RECT 106.270 179.710 106.590 179.770 ;
        RECT 108.125 179.725 108.415 179.770 ;
        RECT 108.585 179.725 108.875 179.955 ;
        RECT 109.045 179.910 109.335 179.955 ;
        RECT 109.490 179.910 109.810 179.970 ;
        RECT 109.045 179.770 109.810 179.910 ;
        RECT 109.045 179.725 109.335 179.770 ;
        RECT 90.630 179.430 103.280 179.570 ;
        RECT 103.510 179.570 103.830 179.630 ;
        RECT 108.660 179.570 108.800 179.725 ;
        RECT 109.490 179.710 109.810 179.770 ;
        RECT 109.965 179.910 110.255 179.955 ;
        RECT 110.425 179.910 110.715 179.955 ;
        RECT 110.870 179.910 111.190 179.970 ;
        RECT 111.420 179.955 111.560 180.110 ;
        RECT 113.170 180.050 113.490 180.110 ;
        RECT 109.965 179.770 111.190 179.910 ;
        RECT 109.965 179.725 110.255 179.770 ;
        RECT 110.425 179.725 110.715 179.770 ;
        RECT 110.870 179.710 111.190 179.770 ;
        RECT 111.345 179.725 111.635 179.955 ;
        RECT 111.790 179.710 112.110 179.970 ;
        RECT 112.265 179.910 112.555 179.955 ;
        RECT 112.710 179.910 113.030 179.970 ;
        RECT 116.020 179.955 116.160 180.450 ;
        RECT 120.185 180.450 125.485 180.590 ;
        RECT 120.185 180.405 120.475 180.450 ;
        RECT 123.305 180.405 123.595 180.450 ;
        RECT 125.195 180.405 125.485 180.450 ;
        RECT 124.210 180.250 124.530 180.310 ;
        RECT 124.685 180.250 124.975 180.295 ;
        RECT 124.210 180.110 124.975 180.250 ;
        RECT 124.210 180.050 124.530 180.110 ;
        RECT 124.685 180.065 124.975 180.110 ;
        RECT 112.265 179.770 113.030 179.910 ;
        RECT 112.265 179.725 112.555 179.770 ;
        RECT 112.710 179.710 113.030 179.770 ;
        RECT 115.945 179.910 116.235 179.955 ;
        RECT 116.850 179.910 117.170 179.970 ;
        RECT 115.945 179.770 117.170 179.910 ;
        RECT 115.945 179.725 116.235 179.770 ;
        RECT 116.850 179.710 117.170 179.770 ;
        RECT 111.880 179.570 112.020 179.710 ;
        RECT 119.105 179.615 119.395 179.930 ;
        RECT 120.185 179.910 120.475 179.955 ;
        RECT 123.765 179.910 124.055 179.955 ;
        RECT 125.600 179.910 125.890 179.955 ;
        RECT 120.185 179.770 125.890 179.910 ;
        RECT 120.185 179.725 120.475 179.770 ;
        RECT 123.765 179.725 124.055 179.770 ;
        RECT 125.600 179.725 125.890 179.770 ;
        RECT 126.065 179.725 126.355 179.955 ;
        RECT 103.510 179.430 112.020 179.570 ;
        RECT 116.405 179.570 116.695 179.615 ;
        RECT 118.805 179.570 119.395 179.615 ;
        RECT 122.045 179.570 122.695 179.615 ;
        RECT 116.405 179.430 122.695 179.570 ;
        RECT 90.630 179.370 90.950 179.430 ;
        RECT 103.510 179.370 103.830 179.430 ;
        RECT 116.405 179.385 116.695 179.430 ;
        RECT 118.805 179.385 119.095 179.430 ;
        RECT 122.045 179.385 122.695 179.430 ;
        RECT 124.670 179.570 124.990 179.630 ;
        RECT 126.140 179.570 126.280 179.725 ;
        RECT 124.670 179.430 126.280 179.570 ;
        RECT 124.670 179.370 124.990 179.430 ;
        RECT 36.825 179.045 37.115 179.275 ;
        RECT 39.125 179.230 39.415 179.275 ;
        RECT 40.950 179.230 41.270 179.290 ;
        RECT 39.125 179.090 41.270 179.230 ;
        RECT 39.125 179.045 39.415 179.090 ;
        RECT 40.950 179.030 41.270 179.090 ;
        RECT 45.550 179.230 45.870 179.290 ;
        RECT 46.485 179.230 46.775 179.275 ;
        RECT 45.550 179.090 46.775 179.230 ;
        RECT 45.550 179.030 45.870 179.090 ;
        RECT 46.485 179.045 46.775 179.090 ;
        RECT 48.310 179.230 48.630 179.290 ;
        RECT 51.530 179.230 51.850 179.290 ;
        RECT 48.310 179.090 51.850 179.230 ;
        RECT 48.310 179.030 48.630 179.090 ;
        RECT 51.530 179.030 51.850 179.090 ;
        RECT 53.830 179.230 54.150 179.290 ;
        RECT 54.765 179.230 55.055 179.275 ;
        RECT 58.445 179.230 58.735 179.275 ;
        RECT 53.830 179.090 58.735 179.230 ;
        RECT 53.830 179.030 54.150 179.090 ;
        RECT 54.765 179.045 55.055 179.090 ;
        RECT 58.445 179.045 58.735 179.090 ;
        RECT 60.745 179.230 61.035 179.275 ;
        RECT 64.410 179.230 64.730 179.290 ;
        RECT 60.745 179.090 64.730 179.230 ;
        RECT 60.745 179.045 61.035 179.090 ;
        RECT 64.410 179.030 64.730 179.090 ;
        RECT 69.010 179.230 69.330 179.290 ;
        RECT 71.770 179.230 72.090 179.290 ;
        RECT 74.990 179.230 75.310 179.290 ;
        RECT 69.010 179.090 75.310 179.230 ;
        RECT 69.010 179.030 69.330 179.090 ;
        RECT 71.770 179.030 72.090 179.090 ;
        RECT 74.990 179.030 75.310 179.090 ;
        RECT 82.350 179.230 82.670 179.290 ;
        RECT 83.285 179.230 83.575 179.275 ;
        RECT 82.350 179.090 83.575 179.230 ;
        RECT 82.350 179.030 82.670 179.090 ;
        RECT 83.285 179.045 83.575 179.090 ;
        RECT 102.605 179.230 102.895 179.275 ;
        RECT 103.050 179.230 103.370 179.290 ;
        RECT 102.605 179.090 103.370 179.230 ;
        RECT 102.605 179.045 102.895 179.090 ;
        RECT 103.050 179.030 103.370 179.090 ;
        RECT 106.745 179.230 107.035 179.275 ;
        RECT 109.490 179.230 109.810 179.290 ;
        RECT 106.745 179.090 109.810 179.230 ;
        RECT 106.745 179.045 107.035 179.090 ;
        RECT 109.490 179.030 109.810 179.090 ;
        RECT 113.645 179.230 113.935 179.275 ;
        RECT 114.550 179.230 114.870 179.290 ;
        RECT 113.645 179.090 114.870 179.230 ;
        RECT 113.645 179.045 113.935 179.090 ;
        RECT 114.550 179.030 114.870 179.090 ;
        RECT 117.310 179.030 117.630 179.290 ;
        RECT 20.640 178.410 127.820 178.890 ;
        RECT 40.490 178.010 40.810 178.270 ;
        RECT 50.150 178.210 50.470 178.270 ;
        RECT 47.020 178.070 50.470 178.210 ;
        RECT 40.580 177.870 40.720 178.010 ;
        RECT 40.580 177.730 45.320 177.870 ;
        RECT 39.125 177.530 39.415 177.575 ;
        RECT 39.570 177.530 39.890 177.590 ;
        RECT 39.125 177.390 39.890 177.530 ;
        RECT 39.125 177.345 39.415 177.390 ;
        RECT 39.570 177.330 39.890 177.390 ;
        RECT 40.030 177.330 40.350 177.590 ;
        RECT 40.505 177.345 40.795 177.575 ;
        RECT 40.965 177.530 41.255 177.575 ;
        RECT 41.870 177.530 42.190 177.590 ;
        RECT 44.185 177.530 44.475 177.575 ;
        RECT 40.965 177.390 44.475 177.530 ;
        RECT 40.965 177.345 41.255 177.390 ;
        RECT 40.580 176.850 40.720 177.345 ;
        RECT 41.870 177.330 42.190 177.390 ;
        RECT 44.185 177.345 44.475 177.390 ;
        RECT 41.410 177.190 41.730 177.250 ;
        RECT 42.345 177.190 42.635 177.235 ;
        RECT 41.410 177.050 42.635 177.190 ;
        RECT 44.260 177.190 44.400 177.345 ;
        RECT 44.630 177.330 44.950 177.590 ;
        RECT 45.180 177.575 45.320 177.730 ;
        RECT 45.105 177.345 45.395 177.575 ;
        RECT 46.025 177.530 46.315 177.575 ;
        RECT 46.485 177.530 46.775 177.575 ;
        RECT 47.020 177.530 47.160 178.070 ;
        RECT 50.150 178.010 50.470 178.070 ;
        RECT 53.830 178.010 54.150 178.270 ;
        RECT 63.505 178.210 63.795 178.255 ;
        RECT 73.150 178.210 73.470 178.270 ;
        RECT 74.530 178.210 74.850 178.270 ;
        RECT 61.280 178.070 63.795 178.210 ;
        RECT 54.290 177.870 54.610 177.930 ;
        RECT 58.890 177.915 59.210 177.930 ;
        RECT 61.280 177.915 61.420 178.070 ;
        RECT 63.505 178.025 63.795 178.070 ;
        RECT 68.180 178.070 74.850 178.210 ;
        RECT 47.480 177.730 54.610 177.870 ;
        RECT 47.480 177.575 47.620 177.730 ;
        RECT 54.290 177.670 54.610 177.730 ;
        RECT 55.325 177.870 55.615 177.915 ;
        RECT 58.565 177.870 59.215 177.915 ;
        RECT 55.325 177.730 59.215 177.870 ;
        RECT 55.325 177.685 55.915 177.730 ;
        RECT 58.565 177.685 59.215 177.730 ;
        RECT 61.205 177.685 61.495 177.915 ;
        RECT 46.025 177.390 47.160 177.530 ;
        RECT 46.025 177.345 46.315 177.390 ;
        RECT 46.485 177.345 46.775 177.390 ;
        RECT 47.405 177.345 47.695 177.575 ;
        RECT 47.850 177.330 48.170 177.590 ;
        RECT 48.310 177.330 48.630 177.590 ;
        RECT 50.150 177.330 50.470 177.590 ;
        RECT 51.070 177.330 51.390 177.590 ;
        RECT 51.530 177.330 51.850 177.590 ;
        RECT 51.990 177.330 52.310 177.590 ;
        RECT 55.625 177.370 55.915 177.685 ;
        RECT 58.890 177.670 59.210 177.685 ;
        RECT 56.705 177.530 56.995 177.575 ;
        RECT 60.285 177.530 60.575 177.575 ;
        RECT 62.120 177.530 62.410 177.575 ;
        RECT 56.705 177.390 62.410 177.530 ;
        RECT 56.705 177.345 56.995 177.390 ;
        RECT 60.285 177.345 60.575 177.390 ;
        RECT 62.120 177.345 62.410 177.390 ;
        RECT 64.410 177.330 64.730 177.590 ;
        RECT 67.185 177.530 67.475 177.575 ;
        RECT 68.180 177.530 68.320 178.070 ;
        RECT 69.025 177.530 69.315 177.575 ;
        RECT 67.185 177.390 67.860 177.530 ;
        RECT 68.180 177.390 69.315 177.530 ;
        RECT 67.185 177.345 67.475 177.390 ;
        RECT 58.430 177.190 58.750 177.250 ;
        RECT 62.585 177.190 62.875 177.235 ;
        RECT 63.950 177.190 64.270 177.250 ;
        RECT 44.260 177.050 54.060 177.190 ;
        RECT 41.410 176.990 41.730 177.050 ;
        RECT 42.345 177.005 42.635 177.050 ;
        RECT 44.170 176.850 44.490 176.910 ;
        RECT 40.580 176.710 44.490 176.850 ;
        RECT 44.170 176.650 44.490 176.710 ;
        RECT 44.630 176.850 44.950 176.910 ;
        RECT 47.850 176.850 48.170 176.910 ;
        RECT 51.530 176.850 51.850 176.910 ;
        RECT 44.630 176.710 51.850 176.850 ;
        RECT 44.630 176.650 44.950 176.710 ;
        RECT 47.850 176.650 48.170 176.710 ;
        RECT 51.530 176.650 51.850 176.710 ;
        RECT 42.330 176.510 42.650 176.570 ;
        RECT 42.805 176.510 43.095 176.555 ;
        RECT 42.330 176.370 43.095 176.510 ;
        RECT 42.330 176.310 42.650 176.370 ;
        RECT 42.805 176.325 43.095 176.370 ;
        RECT 46.470 176.510 46.790 176.570 ;
        RECT 49.705 176.510 49.995 176.555 ;
        RECT 46.470 176.370 49.995 176.510 ;
        RECT 46.470 176.310 46.790 176.370 ;
        RECT 49.705 176.325 49.995 176.370 ;
        RECT 52.910 176.510 53.230 176.570 ;
        RECT 53.385 176.510 53.675 176.555 ;
        RECT 52.910 176.370 53.675 176.510 ;
        RECT 53.920 176.510 54.060 177.050 ;
        RECT 58.430 177.050 64.270 177.190 ;
        RECT 58.430 176.990 58.750 177.050 ;
        RECT 62.585 177.005 62.875 177.050 ;
        RECT 63.950 176.990 64.270 177.050 ;
        RECT 56.705 176.850 56.995 176.895 ;
        RECT 59.825 176.850 60.115 176.895 ;
        RECT 61.715 176.850 62.005 176.895 ;
        RECT 56.705 176.710 62.005 176.850 ;
        RECT 56.705 176.665 56.995 176.710 ;
        RECT 59.825 176.665 60.115 176.710 ;
        RECT 61.715 176.665 62.005 176.710 ;
        RECT 67.720 176.570 67.860 177.390 ;
        RECT 69.025 177.345 69.315 177.390 ;
        RECT 69.945 177.530 70.235 177.575 ;
        RECT 70.390 177.530 70.710 177.590 ;
        RECT 69.945 177.390 70.710 177.530 ;
        RECT 69.945 177.345 70.235 177.390 ;
        RECT 70.390 177.330 70.710 177.390 ;
        RECT 71.785 177.530 72.075 177.575 ;
        RECT 72.780 177.530 72.920 178.070 ;
        RECT 73.150 178.010 73.470 178.070 ;
        RECT 74.530 178.010 74.850 178.070 ;
        RECT 74.990 178.010 75.310 178.270 ;
        RECT 81.430 178.210 81.750 178.270 ;
        RECT 111.790 178.210 112.110 178.270 ;
        RECT 81.430 178.070 85.340 178.210 ;
        RECT 81.430 178.010 81.750 178.070 ;
        RECT 75.080 177.870 75.220 178.010 ;
        RECT 71.785 177.390 72.920 177.530 ;
        RECT 73.240 177.730 75.220 177.870 ;
        RECT 81.060 177.730 84.880 177.870 ;
        RECT 71.785 177.345 72.075 177.390 ;
        RECT 68.550 176.990 68.870 177.250 ;
        RECT 69.470 176.990 69.790 177.250 ;
        RECT 72.230 176.990 72.550 177.250 ;
        RECT 73.240 177.235 73.380 177.730 ;
        RECT 81.060 177.590 81.200 177.730 ;
        RECT 74.085 177.530 74.375 177.575 ;
        RECT 74.990 177.530 75.310 177.590 ;
        RECT 74.085 177.390 75.310 177.530 ;
        RECT 74.085 177.345 74.375 177.390 ;
        RECT 74.990 177.330 75.310 177.390 ;
        RECT 80.970 177.330 81.290 177.590 ;
        RECT 81.430 177.330 81.750 177.590 ;
        RECT 81.890 177.330 82.210 177.590 ;
        RECT 84.740 177.575 84.880 177.730 ;
        RECT 85.200 177.575 85.340 178.070 ;
        RECT 110.500 178.070 112.110 178.210 ;
        RECT 90.170 177.870 90.490 177.930 ;
        RECT 85.660 177.730 90.490 177.870 ;
        RECT 85.660 177.575 85.800 177.730 ;
        RECT 90.170 177.670 90.490 177.730 ;
        RECT 90.630 177.670 90.950 177.930 ;
        RECT 98.910 177.870 99.230 177.930 ;
        RECT 96.700 177.730 99.230 177.870 ;
        RECT 82.825 177.530 83.115 177.575 ;
        RECT 82.715 177.390 83.115 177.530 ;
        RECT 82.825 177.345 83.115 177.390 ;
        RECT 84.665 177.345 84.955 177.575 ;
        RECT 85.125 177.345 85.415 177.575 ;
        RECT 85.585 177.345 85.875 177.575 ;
        RECT 72.705 177.005 72.995 177.235 ;
        RECT 73.165 177.005 73.455 177.235 ;
        RECT 82.900 177.190 83.040 177.345 ;
        RECT 86.490 177.330 86.810 177.590 ;
        RECT 86.950 177.530 87.270 177.590 ;
        RECT 89.265 177.530 89.555 177.575 ;
        RECT 86.950 177.390 89.555 177.530 ;
        RECT 86.950 177.330 87.270 177.390 ;
        RECT 89.265 177.345 89.555 177.390 ;
        RECT 94.770 177.530 95.090 177.590 ;
        RECT 96.700 177.575 96.840 177.730 ;
        RECT 98.910 177.670 99.230 177.730 ;
        RECT 100.865 177.870 101.155 177.915 ;
        RECT 103.050 177.870 103.370 177.930 ;
        RECT 104.105 177.870 104.755 177.915 ;
        RECT 100.865 177.730 104.755 177.870 ;
        RECT 100.865 177.685 101.455 177.730 ;
        RECT 95.705 177.530 95.995 177.575 ;
        RECT 94.770 177.390 95.995 177.530 ;
        RECT 94.770 177.330 95.090 177.390 ;
        RECT 95.705 177.345 95.995 177.390 ;
        RECT 96.625 177.345 96.915 177.575 ;
        RECT 97.070 177.330 97.390 177.590 ;
        RECT 97.545 177.345 97.835 177.575 ;
        RECT 101.165 177.370 101.455 177.685 ;
        RECT 103.050 177.670 103.370 177.730 ;
        RECT 104.105 177.685 104.755 177.730 ;
        RECT 110.500 177.605 110.640 178.070 ;
        RECT 111.790 178.010 112.110 178.070 ;
        RECT 123.305 178.210 123.595 178.255 ;
        RECT 124.210 178.210 124.530 178.270 ;
        RECT 123.305 178.070 124.530 178.210 ;
        RECT 123.305 178.025 123.595 178.070 ;
        RECT 124.210 178.010 124.530 178.070 ;
        RECT 102.245 177.530 102.535 177.575 ;
        RECT 105.825 177.530 106.115 177.575 ;
        RECT 107.660 177.530 107.950 177.575 ;
        RECT 102.245 177.390 107.950 177.530 ;
        RECT 102.245 177.345 102.535 177.390 ;
        RECT 105.825 177.345 106.115 177.390 ;
        RECT 107.660 177.345 107.950 177.390 ;
        RECT 108.125 177.530 108.415 177.575 ;
        RECT 109.030 177.530 109.350 177.590 ;
        RECT 108.125 177.390 109.350 177.530 ;
        RECT 108.125 177.345 108.415 177.390 ;
        RECT 86.580 177.190 86.720 177.330 ;
        RECT 97.620 177.190 97.760 177.345 ;
        RECT 109.030 177.330 109.350 177.390 ;
        RECT 109.950 177.330 110.270 177.590 ;
        RECT 110.425 177.375 110.715 177.605 ;
        RECT 110.885 177.530 111.175 177.575 ;
        RECT 111.330 177.530 111.650 177.590 ;
        RECT 110.885 177.390 111.650 177.530 ;
        RECT 110.885 177.345 111.175 177.390 ;
        RECT 111.330 177.330 111.650 177.390 ;
        RECT 111.805 177.345 112.095 177.575 ;
        RECT 116.850 177.530 117.170 177.590 ;
        RECT 118.705 177.530 118.995 177.575 ;
        RECT 116.850 177.390 118.995 177.530 ;
        RECT 106.270 177.190 106.590 177.250 ;
        RECT 82.900 177.050 86.720 177.190 ;
        RECT 97.160 177.050 106.590 177.190 ;
        RECT 69.560 176.850 69.700 176.990 ;
        RECT 72.780 176.850 72.920 177.005 ;
        RECT 82.900 176.910 83.040 177.050 ;
        RECT 75.005 176.850 75.295 176.895 ;
        RECT 75.910 176.850 76.230 176.910 ;
        RECT 82.810 176.850 83.130 176.910 ;
        RECT 69.560 176.710 74.760 176.850 ;
        RECT 63.950 176.510 64.270 176.570 ;
        RECT 53.920 176.370 64.270 176.510 ;
        RECT 52.910 176.310 53.230 176.370 ;
        RECT 53.385 176.325 53.675 176.370 ;
        RECT 63.950 176.310 64.270 176.370 ;
        RECT 66.250 176.310 66.570 176.570 ;
        RECT 67.630 176.310 67.950 176.570 ;
        RECT 70.865 176.510 71.155 176.555 ;
        RECT 71.310 176.510 71.630 176.570 ;
        RECT 70.865 176.370 71.630 176.510 ;
        RECT 74.620 176.510 74.760 176.710 ;
        RECT 75.005 176.710 83.130 176.850 ;
        RECT 75.005 176.665 75.295 176.710 ;
        RECT 75.910 176.650 76.230 176.710 ;
        RECT 82.810 176.650 83.130 176.710 ;
        RECT 83.270 176.650 83.590 176.910 ;
        RECT 83.730 176.850 84.050 176.910 ;
        RECT 97.160 176.850 97.300 177.050 ;
        RECT 106.270 176.990 106.590 177.050 ;
        RECT 106.730 176.990 107.050 177.250 ;
        RECT 83.730 176.710 97.300 176.850 ;
        RECT 83.730 176.650 84.050 176.710 ;
        RECT 99.370 176.650 99.690 176.910 ;
        RECT 102.245 176.850 102.535 176.895 ;
        RECT 105.365 176.850 105.655 176.895 ;
        RECT 107.255 176.850 107.545 176.895 ;
        RECT 102.245 176.710 107.545 176.850 ;
        RECT 102.245 176.665 102.535 176.710 ;
        RECT 105.365 176.665 105.655 176.710 ;
        RECT 107.255 176.665 107.545 176.710 ;
        RECT 108.110 176.850 108.430 176.910 ;
        RECT 110.870 176.850 111.190 176.910 ;
        RECT 111.880 176.850 112.020 177.345 ;
        RECT 116.850 177.330 117.170 177.390 ;
        RECT 118.705 177.345 118.995 177.390 ;
        RECT 122.385 177.345 122.675 177.575 ;
        RECT 115.470 177.190 115.790 177.250 ;
        RECT 122.460 177.190 122.600 177.345 ;
        RECT 115.470 177.050 122.600 177.190 ;
        RECT 115.470 176.990 115.790 177.050 ;
        RECT 108.110 176.710 112.020 176.850 ;
        RECT 108.110 176.650 108.430 176.710 ;
        RECT 110.870 176.650 111.190 176.710 ;
        RECT 78.670 176.510 78.990 176.570 ;
        RECT 74.620 176.370 78.990 176.510 ;
        RECT 70.865 176.325 71.155 176.370 ;
        RECT 71.310 176.310 71.630 176.370 ;
        RECT 78.670 176.310 78.990 176.370 ;
        RECT 79.590 176.310 79.910 176.570 ;
        RECT 98.925 176.510 99.215 176.555 ;
        RECT 99.830 176.510 100.150 176.570 ;
        RECT 98.925 176.370 100.150 176.510 ;
        RECT 98.925 176.325 99.215 176.370 ;
        RECT 99.830 176.310 100.150 176.370 ;
        RECT 103.970 176.510 104.290 176.570 ;
        RECT 108.585 176.510 108.875 176.555 ;
        RECT 103.970 176.370 108.875 176.510 ;
        RECT 103.970 176.310 104.290 176.370 ;
        RECT 108.585 176.325 108.875 176.370 ;
        RECT 118.230 176.510 118.550 176.570 ;
        RECT 119.165 176.510 119.455 176.555 ;
        RECT 118.230 176.370 119.455 176.510 ;
        RECT 118.230 176.310 118.550 176.370 ;
        RECT 119.165 176.325 119.455 176.370 ;
        RECT 20.640 175.690 127.820 176.170 ;
        RECT 45.090 175.490 45.410 175.550 ;
        RECT 48.310 175.490 48.630 175.550 ;
        RECT 45.090 175.350 48.630 175.490 ;
        RECT 45.090 175.290 45.410 175.350 ;
        RECT 48.310 175.290 48.630 175.350 ;
        RECT 50.150 175.490 50.470 175.550 ;
        RECT 56.590 175.490 56.910 175.550 ;
        RECT 50.150 175.350 56.910 175.490 ;
        RECT 50.150 175.290 50.470 175.350 ;
        RECT 56.590 175.290 56.910 175.350 ;
        RECT 58.890 175.490 59.210 175.550 ;
        RECT 61.205 175.490 61.495 175.535 ;
        RECT 58.890 175.350 61.495 175.490 ;
        RECT 58.890 175.290 59.210 175.350 ;
        RECT 61.205 175.305 61.495 175.350 ;
        RECT 63.950 175.490 64.270 175.550 ;
        RECT 68.550 175.490 68.870 175.550 ;
        RECT 63.950 175.350 68.870 175.490 ;
        RECT 63.950 175.290 64.270 175.350 ;
        RECT 68.550 175.290 68.870 175.350 ;
        RECT 70.390 175.490 70.710 175.550 ;
        RECT 72.230 175.490 72.550 175.550 ;
        RECT 70.390 175.350 72.550 175.490 ;
        RECT 70.390 175.290 70.710 175.350 ;
        RECT 72.230 175.290 72.550 175.350 ;
        RECT 73.610 175.290 73.930 175.550 ;
        RECT 74.530 175.490 74.850 175.550 ;
        RECT 81.890 175.490 82.210 175.550 ;
        RECT 85.570 175.490 85.890 175.550 ;
        RECT 74.530 175.350 77.980 175.490 ;
        RECT 74.530 175.290 74.850 175.350 ;
        RECT 25.735 175.150 26.025 175.195 ;
        RECT 27.625 175.150 27.915 175.195 ;
        RECT 30.745 175.150 31.035 175.195 ;
        RECT 25.735 175.010 31.035 175.150 ;
        RECT 25.735 174.965 26.025 175.010 ;
        RECT 27.625 174.965 27.915 175.010 ;
        RECT 30.745 174.965 31.035 175.010 ;
        RECT 37.730 175.150 38.050 175.210 ;
        RECT 43.265 175.150 43.555 175.195 ;
        RECT 37.730 175.010 43.555 175.150 ;
        RECT 37.730 174.950 38.050 175.010 ;
        RECT 43.265 174.965 43.555 175.010 ;
        RECT 51.990 175.150 52.310 175.210 ;
        RECT 57.065 175.150 57.355 175.195 ;
        RECT 51.990 175.010 57.355 175.150 ;
        RECT 51.990 174.950 52.310 175.010 ;
        RECT 57.065 174.965 57.355 175.010 ;
        RECT 71.770 175.150 72.090 175.210 ;
        RECT 71.770 175.010 77.520 175.150 ;
        RECT 71.770 174.950 72.090 175.010 ;
        RECT 26.230 174.610 26.550 174.870 ;
        RECT 53.830 174.810 54.150 174.870 ;
        RECT 66.250 174.810 66.570 174.870 ;
        RECT 37.820 174.670 42.100 174.810 ;
        RECT 24.850 174.270 25.170 174.530 ;
        RECT 37.820 174.515 37.960 174.670 ;
        RECT 41.960 174.530 42.100 174.670 ;
        RECT 53.830 174.670 55.900 174.810 ;
        RECT 53.830 174.610 54.150 174.670 ;
        RECT 25.330 174.470 25.620 174.515 ;
        RECT 27.165 174.470 27.455 174.515 ;
        RECT 30.745 174.470 31.035 174.515 ;
        RECT 25.330 174.330 31.035 174.470 ;
        RECT 25.330 174.285 25.620 174.330 ;
        RECT 27.165 174.285 27.455 174.330 ;
        RECT 30.745 174.285 31.035 174.330 ;
        RECT 24.390 174.130 24.710 174.190 ;
        RECT 31.825 174.175 32.115 174.490 ;
        RECT 37.745 174.285 38.035 174.515 ;
        RECT 38.205 174.285 38.495 174.515 ;
        RECT 28.525 174.130 29.175 174.175 ;
        RECT 31.825 174.130 32.415 174.175 ;
        RECT 24.390 173.990 32.415 174.130 ;
        RECT 24.390 173.930 24.710 173.990 ;
        RECT 28.525 173.945 29.175 173.990 ;
        RECT 32.125 173.945 32.415 173.990 ;
        RECT 36.350 173.930 36.670 174.190 ;
        RECT 38.280 174.130 38.420 174.285 ;
        RECT 38.650 174.270 38.970 174.530 ;
        RECT 39.570 174.470 39.890 174.530 ;
        RECT 40.045 174.470 40.335 174.515 ;
        RECT 39.570 174.330 40.335 174.470 ;
        RECT 39.570 174.270 39.890 174.330 ;
        RECT 40.045 174.285 40.335 174.330 ;
        RECT 40.950 174.270 41.270 174.530 ;
        RECT 41.425 174.285 41.715 174.515 ;
        RECT 41.500 174.130 41.640 174.285 ;
        RECT 41.870 174.270 42.190 174.530 ;
        RECT 52.450 174.470 52.770 174.530 ;
        RECT 54.765 174.470 55.055 174.515 ;
        RECT 52.450 174.330 55.055 174.470 ;
        RECT 52.450 174.270 52.770 174.330 ;
        RECT 54.765 174.285 55.055 174.330 ;
        RECT 44.170 174.130 44.490 174.190 ;
        RECT 38.280 173.990 44.490 174.130 ;
        RECT 44.170 173.930 44.490 173.990 ;
        RECT 51.070 174.130 51.390 174.190 ;
        RECT 53.385 174.130 53.675 174.175 ;
        RECT 51.070 173.990 53.675 174.130 ;
        RECT 54.840 174.130 54.980 174.285 ;
        RECT 55.210 174.270 55.530 174.530 ;
        RECT 55.760 174.515 55.900 174.670 ;
        RECT 57.140 174.670 66.570 174.810 ;
        RECT 55.685 174.285 55.975 174.515 ;
        RECT 56.590 174.270 56.910 174.530 ;
        RECT 57.140 174.130 57.280 174.670 ;
        RECT 58.520 174.515 58.660 174.670 ;
        RECT 66.250 174.610 66.570 174.670 ;
        RECT 72.230 174.810 72.550 174.870 ;
        RECT 77.380 174.855 77.520 175.010 ;
        RECT 77.840 174.855 77.980 175.350 ;
        RECT 81.890 175.350 85.890 175.490 ;
        RECT 81.890 175.290 82.210 175.350 ;
        RECT 85.570 175.290 85.890 175.350 ;
        RECT 86.950 175.490 87.270 175.550 ;
        RECT 105.365 175.490 105.655 175.535 ;
        RECT 106.730 175.490 107.050 175.550 ;
        RECT 111.790 175.490 112.110 175.550 ;
        RECT 86.950 175.350 94.080 175.490 ;
        RECT 86.950 175.290 87.270 175.350 ;
        RECT 86.050 175.150 86.340 175.195 ;
        RECT 87.910 175.150 88.200 175.195 ;
        RECT 90.690 175.150 90.980 175.195 ;
        RECT 86.050 175.010 90.980 175.150 ;
        RECT 86.050 174.965 86.340 175.010 ;
        RECT 87.910 174.965 88.200 175.010 ;
        RECT 90.690 174.965 90.980 175.010 ;
        RECT 72.230 174.670 76.140 174.810 ;
        RECT 72.230 174.610 72.550 174.670 ;
        RECT 58.445 174.285 58.735 174.515 ;
        RECT 58.890 174.270 59.210 174.530 ;
        RECT 59.365 174.470 59.655 174.515 ;
        RECT 59.810 174.470 60.130 174.530 ;
        RECT 59.365 174.330 60.130 174.470 ;
        RECT 59.365 174.285 59.655 174.330 ;
        RECT 59.810 174.270 60.130 174.330 ;
        RECT 60.270 174.270 60.590 174.530 ;
        RECT 61.190 174.470 61.510 174.530 ;
        RECT 61.665 174.470 61.955 174.515 ;
        RECT 61.190 174.330 61.955 174.470 ;
        RECT 61.190 174.270 61.510 174.330 ;
        RECT 61.665 174.285 61.955 174.330 ;
        RECT 67.630 174.470 67.950 174.530 ;
        RECT 69.485 174.470 69.775 174.515 ;
        RECT 69.945 174.470 70.235 174.515 ;
        RECT 67.630 174.330 70.235 174.470 ;
        RECT 67.630 174.270 67.950 174.330 ;
        RECT 69.485 174.285 69.775 174.330 ;
        RECT 69.945 174.285 70.235 174.330 ;
        RECT 71.310 174.270 71.630 174.530 ;
        RECT 73.150 174.270 73.470 174.530 ;
        RECT 74.085 174.285 74.375 174.515 ;
        RECT 54.840 173.990 57.280 174.130 ;
        RECT 57.600 173.990 58.660 174.130 ;
        RECT 51.070 173.930 51.390 173.990 ;
        RECT 53.385 173.945 53.675 173.990 ;
        RECT 29.910 173.790 30.230 173.850 ;
        RECT 33.605 173.790 33.895 173.835 ;
        RECT 29.910 173.650 33.895 173.790 ;
        RECT 29.910 173.590 30.230 173.650 ;
        RECT 33.605 173.605 33.895 173.650 ;
        RECT 55.210 173.790 55.530 173.850 ;
        RECT 57.600 173.790 57.740 173.990 ;
        RECT 58.520 173.940 58.660 173.990 ;
        RECT 58.890 173.940 59.210 174.000 ;
        RECT 58.520 173.800 59.210 173.940 ;
        RECT 55.210 173.650 57.740 173.790 ;
        RECT 58.890 173.740 59.210 173.800 ;
        RECT 74.160 173.790 74.300 174.285 ;
        RECT 75.450 174.270 75.770 174.530 ;
        RECT 76.000 174.470 76.140 174.670 ;
        RECT 77.305 174.625 77.595 174.855 ;
        RECT 77.765 174.625 78.055 174.855 ;
        RECT 78.670 174.610 78.990 174.870 ;
        RECT 81.430 174.810 81.750 174.870 ;
        RECT 84.650 174.810 84.970 174.870 ;
        RECT 87.425 174.810 87.715 174.855 ;
        RECT 89.250 174.810 89.570 174.870 ;
        RECT 81.430 174.670 83.960 174.810 ;
        RECT 81.430 174.610 81.750 174.670 ;
        RECT 78.225 174.470 78.515 174.515 ;
        RECT 79.130 174.470 79.450 174.530 ;
        RECT 76.000 174.330 79.450 174.470 ;
        RECT 78.225 174.285 78.515 174.330 ;
        RECT 79.130 174.270 79.450 174.330 ;
        RECT 80.970 174.470 81.290 174.530 ;
        RECT 83.820 174.515 83.960 174.670 ;
        RECT 84.650 174.670 87.715 174.810 ;
        RECT 84.650 174.610 84.970 174.670 ;
        RECT 87.425 174.625 87.715 174.670 ;
        RECT 87.960 174.670 89.570 174.810 ;
        RECT 83.285 174.470 83.575 174.515 ;
        RECT 80.970 174.330 83.575 174.470 ;
        RECT 80.970 174.270 81.290 174.330 ;
        RECT 83.285 174.285 83.575 174.330 ;
        RECT 83.745 174.285 84.035 174.515 ;
        RECT 84.190 174.270 84.510 174.530 ;
        RECT 85.125 174.285 85.415 174.515 ;
        RECT 85.585 174.470 85.875 174.515 ;
        RECT 87.960 174.470 88.100 174.670 ;
        RECT 89.250 174.610 89.570 174.670 ;
        RECT 90.690 174.470 90.980 174.515 ;
        RECT 85.585 174.330 88.100 174.470 ;
        RECT 88.445 174.330 90.980 174.470 ;
        RECT 85.585 174.285 85.875 174.330 ;
        RECT 74.530 174.130 74.850 174.190 ;
        RECT 76.385 174.130 76.675 174.175 ;
        RECT 74.530 173.990 76.675 174.130 ;
        RECT 74.530 173.930 74.850 173.990 ;
        RECT 76.385 173.945 76.675 173.990 ;
        RECT 81.890 173.930 82.210 174.190 ;
        RECT 82.810 174.130 83.130 174.190 ;
        RECT 85.200 174.130 85.340 174.285 ;
        RECT 88.445 174.175 88.660 174.330 ;
        RECT 90.690 174.285 90.980 174.330 ;
        RECT 93.940 174.470 94.080 175.350 ;
        RECT 100.840 175.350 105.120 175.490 ;
        RECT 100.840 175.150 100.980 175.350 ;
        RECT 94.860 175.010 100.980 175.150 ;
        RECT 94.860 174.870 95.000 175.010 ;
        RECT 101.225 174.965 101.515 175.195 ;
        RECT 94.770 174.610 95.090 174.870 ;
        RECT 98.465 174.810 98.755 174.855 ;
        RECT 100.750 174.810 101.070 174.870 ;
        RECT 98.465 174.670 101.070 174.810 ;
        RECT 98.465 174.625 98.755 174.670 ;
        RECT 100.750 174.610 101.070 174.670 ;
        RECT 99.385 174.470 99.675 174.515 ;
        RECT 93.940 174.330 99.675 174.470 ;
        RECT 101.300 174.470 101.440 174.965 ;
        RECT 104.445 174.470 104.735 174.515 ;
        RECT 101.300 174.330 104.735 174.470 ;
        RECT 104.980 174.470 105.120 175.350 ;
        RECT 105.365 175.350 107.050 175.490 ;
        RECT 105.365 175.305 105.655 175.350 ;
        RECT 106.730 175.290 107.050 175.350 ;
        RECT 110.040 175.350 112.110 175.490 ;
        RECT 108.570 174.950 108.890 175.210 ;
        RECT 108.110 174.470 108.430 174.530 ;
        RECT 104.980 174.330 108.430 174.470 ;
        RECT 82.810 173.990 85.340 174.130 ;
        RECT 86.510 174.130 86.800 174.175 ;
        RECT 88.370 174.130 88.660 174.175 ;
        RECT 86.510 173.990 88.660 174.130 ;
        RECT 82.810 173.930 83.130 173.990 ;
        RECT 86.510 173.945 86.800 173.990 ;
        RECT 88.370 173.945 88.660 173.990 ;
        RECT 89.290 174.130 89.580 174.175 ;
        RECT 91.090 174.130 91.410 174.190 ;
        RECT 92.550 174.130 92.840 174.175 ;
        RECT 89.290 173.990 92.840 174.130 ;
        RECT 93.940 174.130 94.080 174.330 ;
        RECT 99.385 174.285 99.675 174.330 ;
        RECT 104.445 174.285 104.735 174.330 ;
        RECT 108.110 174.270 108.430 174.330 ;
        RECT 108.660 174.455 108.800 174.950 ;
        RECT 110.040 174.810 110.180 175.350 ;
        RECT 111.790 175.290 112.110 175.350 ;
        RECT 115.470 175.290 115.790 175.550 ;
        RECT 115.945 175.150 116.235 175.195 ;
        RECT 117.770 175.150 118.090 175.210 ;
        RECT 115.945 175.010 118.090 175.150 ;
        RECT 115.945 174.965 116.235 175.010 ;
        RECT 117.770 174.950 118.090 175.010 ;
        RECT 118.805 175.150 119.095 175.195 ;
        RECT 121.925 175.150 122.215 175.195 ;
        RECT 123.815 175.150 124.105 175.195 ;
        RECT 118.805 175.010 124.105 175.150 ;
        RECT 118.805 174.965 119.095 175.010 ;
        RECT 121.925 174.965 122.215 175.010 ;
        RECT 123.815 174.965 124.105 175.010 ;
        RECT 109.580 174.670 110.180 174.810 ;
        RECT 109.580 174.515 109.720 174.670 ;
        RECT 110.410 174.610 110.730 174.870 ;
        RECT 111.330 174.610 111.650 174.870 ;
        RECT 112.710 174.610 113.030 174.870 ;
        RECT 124.670 174.610 124.990 174.870 ;
        RECT 108.940 174.455 109.230 174.500 ;
        RECT 108.660 174.315 109.230 174.455 ;
        RECT 108.940 174.270 109.230 174.315 ;
        RECT 109.505 174.285 109.795 174.515 ;
        RECT 109.965 174.440 110.255 174.515 ;
        RECT 110.500 174.440 110.640 174.610 ;
        RECT 109.965 174.300 110.640 174.440 ;
        RECT 111.420 174.470 111.560 174.610 ;
        RECT 135.635 174.550 136.775 223.880 ;
        RECT 138.130 223.810 139.580 225.110 ;
        RECT 143.180 223.840 144.630 225.140 ;
        RECT 113.645 174.470 113.935 174.515 ;
        RECT 111.420 174.330 113.935 174.470 ;
        RECT 109.965 174.285 110.255 174.300 ;
        RECT 113.645 174.285 113.935 174.330 ;
        RECT 94.555 174.130 94.845 174.175 ;
        RECT 93.940 173.990 94.845 174.130 ;
        RECT 89.290 173.945 89.580 173.990 ;
        RECT 91.090 173.930 91.410 173.990 ;
        RECT 92.550 173.945 92.840 173.990 ;
        RECT 94.555 173.945 94.845 173.990 ;
        RECT 98.910 174.130 99.230 174.190 ;
        RECT 110.870 174.130 111.190 174.190 ;
        RECT 98.910 173.990 111.190 174.130 ;
        RECT 98.910 173.930 99.230 173.990 ;
        RECT 110.870 173.930 111.190 173.990 ;
        RECT 111.330 173.930 111.650 174.190 ;
        RECT 117.725 174.175 118.015 174.490 ;
        RECT 118.805 174.470 119.095 174.515 ;
        RECT 122.385 174.470 122.675 174.515 ;
        RECT 124.220 174.470 124.510 174.515 ;
        RECT 118.805 174.330 124.510 174.470 ;
        RECT 118.805 174.285 119.095 174.330 ;
        RECT 122.385 174.285 122.675 174.330 ;
        RECT 124.220 174.285 124.510 174.330 ;
        RECT 117.425 174.130 118.015 174.175 ;
        RECT 118.230 174.130 118.550 174.190 ;
        RECT 120.665 174.130 121.315 174.175 ;
        RECT 117.425 173.990 121.315 174.130 ;
        RECT 117.425 173.945 117.715 173.990 ;
        RECT 118.230 173.930 118.550 173.990 ;
        RECT 120.665 173.945 121.315 173.990 ;
        RECT 121.910 174.130 122.230 174.190 ;
        RECT 123.305 174.130 123.595 174.175 ;
        RECT 121.910 173.990 123.595 174.130 ;
        RECT 121.910 173.930 122.230 173.990 ;
        RECT 123.305 173.945 123.595 173.990 ;
        RECT 74.990 173.790 75.310 173.850 ;
        RECT 74.160 173.650 75.310 173.790 ;
        RECT 55.210 173.590 55.530 173.650 ;
        RECT 74.990 173.590 75.310 173.650 ;
        RECT 113.170 173.590 113.490 173.850 ;
        RECT 20.640 172.970 127.820 173.450 ;
        RECT 135.580 173.430 136.830 174.550 ;
        RECT 135.635 173.420 136.775 173.430 ;
        RECT 24.390 172.570 24.710 172.830 ;
        RECT 73.610 172.770 73.930 172.830 ;
        RECT 75.465 172.770 75.755 172.815 ;
        RECT 70.020 172.630 75.755 172.770 ;
        RECT 25.785 172.430 26.075 172.475 ;
        RECT 28.185 172.430 28.475 172.475 ;
        RECT 31.425 172.430 32.075 172.475 ;
        RECT 25.785 172.290 32.075 172.430 ;
        RECT 25.785 172.245 26.075 172.290 ;
        RECT 28.185 172.245 28.775 172.290 ;
        RECT 31.425 172.245 32.075 172.290 ;
        RECT 34.065 172.430 34.355 172.475 ;
        RECT 34.510 172.430 34.830 172.490 ;
        RECT 34.065 172.290 34.830 172.430 ;
        RECT 34.065 172.245 34.355 172.290 ;
        RECT 24.865 172.090 25.155 172.135 ;
        RECT 25.325 172.090 25.615 172.135 ;
        RECT 24.865 171.950 28.300 172.090 ;
        RECT 24.865 171.905 25.155 171.950 ;
        RECT 25.325 171.905 25.615 171.950 ;
        RECT 26.690 170.870 27.010 171.130 ;
        RECT 28.160 171.070 28.300 171.950 ;
        RECT 28.485 171.930 28.775 172.245 ;
        RECT 34.510 172.230 34.830 172.290 ;
        RECT 44.630 172.430 44.950 172.490 ;
        RECT 44.630 172.290 45.780 172.430 ;
        RECT 44.630 172.230 44.950 172.290 ;
        RECT 29.565 172.090 29.855 172.135 ;
        RECT 33.145 172.090 33.435 172.135 ;
        RECT 34.980 172.090 35.270 172.135 ;
        RECT 29.565 171.950 35.270 172.090 ;
        RECT 29.565 171.905 29.855 171.950 ;
        RECT 33.145 171.905 33.435 171.950 ;
        RECT 34.980 171.905 35.270 171.950 ;
        RECT 42.345 172.090 42.635 172.135 ;
        RECT 42.345 171.950 44.400 172.090 ;
        RECT 42.345 171.905 42.635 171.950 ;
        RECT 35.430 171.750 35.750 171.810 ;
        RECT 43.710 171.750 44.030 171.810 ;
        RECT 35.430 171.610 44.030 171.750 ;
        RECT 35.430 171.550 35.750 171.610 ;
        RECT 43.710 171.550 44.030 171.610 ;
        RECT 29.565 171.410 29.855 171.455 ;
        RECT 32.685 171.410 32.975 171.455 ;
        RECT 34.575 171.410 34.865 171.455 ;
        RECT 35.890 171.410 36.210 171.470 ;
        RECT 44.260 171.410 44.400 171.950 ;
        RECT 45.090 171.890 45.410 172.150 ;
        RECT 45.640 172.135 45.780 172.290 ;
        RECT 45.565 171.905 45.855 172.135 ;
        RECT 46.010 171.890 46.330 172.150 ;
        RECT 46.945 171.905 47.235 172.135 ;
        RECT 47.020 171.750 47.160 171.905 ;
        RECT 47.390 171.890 47.710 172.150 ;
        RECT 70.020 172.135 70.160 172.630 ;
        RECT 73.610 172.570 73.930 172.630 ;
        RECT 75.465 172.585 75.755 172.630 ;
        RECT 84.205 172.770 84.495 172.815 ;
        RECT 84.650 172.770 84.970 172.830 ;
        RECT 84.205 172.630 84.970 172.770 ;
        RECT 84.205 172.585 84.495 172.630 ;
        RECT 84.650 172.570 84.970 172.630 ;
        RECT 90.645 172.770 90.935 172.815 ;
        RECT 91.090 172.770 91.410 172.830 ;
        RECT 90.645 172.630 91.410 172.770 ;
        RECT 90.645 172.585 90.935 172.630 ;
        RECT 91.090 172.570 91.410 172.630 ;
        RECT 119.625 172.585 119.915 172.815 ;
        RECT 121.465 172.770 121.755 172.815 ;
        RECT 121.910 172.770 122.230 172.830 ;
        RECT 121.465 172.630 122.230 172.770 ;
        RECT 121.465 172.585 121.755 172.630 ;
        RECT 71.770 172.430 72.090 172.490 ;
        RECT 73.165 172.430 73.455 172.475 ;
        RECT 70.940 172.290 73.455 172.430 ;
        RECT 70.940 172.135 71.080 172.290 ;
        RECT 71.770 172.230 72.090 172.290 ;
        RECT 73.165 172.245 73.455 172.290 ;
        RECT 83.730 172.430 84.050 172.490 ;
        RECT 86.505 172.430 86.795 172.475 ;
        RECT 83.730 172.290 86.795 172.430 ;
        RECT 83.730 172.230 84.050 172.290 ;
        RECT 86.505 172.245 86.795 172.290 ;
        RECT 107.665 172.430 107.955 172.475 ;
        RECT 109.030 172.430 109.350 172.490 ;
        RECT 107.665 172.290 109.350 172.430 ;
        RECT 107.665 172.245 107.955 172.290 ;
        RECT 109.030 172.230 109.350 172.290 ;
        RECT 113.170 172.430 113.490 172.490 ;
        RECT 117.310 172.430 117.630 172.490 ;
        RECT 117.785 172.430 118.075 172.475 ;
        RECT 113.170 172.290 118.075 172.430 ;
        RECT 113.170 172.230 113.490 172.290 ;
        RECT 117.310 172.230 117.630 172.290 ;
        RECT 117.785 172.245 118.075 172.290 ;
        RECT 69.945 171.905 70.235 172.135 ;
        RECT 70.405 171.905 70.695 172.135 ;
        RECT 70.865 171.905 71.155 172.135 ;
        RECT 71.325 172.090 71.615 172.135 ;
        RECT 75.450 172.090 75.770 172.150 ;
        RECT 71.325 171.950 75.770 172.090 ;
        RECT 71.325 171.905 71.615 171.950 ;
        RECT 55.670 171.750 55.990 171.810 ;
        RECT 47.020 171.610 55.990 171.750 ;
        RECT 55.670 171.550 55.990 171.610 ;
        RECT 56.145 171.750 56.435 171.795 ;
        RECT 58.430 171.750 58.750 171.810 ;
        RECT 56.145 171.610 58.750 171.750 ;
        RECT 56.145 171.565 56.435 171.610 ;
        RECT 58.430 171.550 58.750 171.610 ;
        RECT 69.470 171.750 69.790 171.810 ;
        RECT 70.480 171.750 70.620 171.905 ;
        RECT 75.450 171.890 75.770 171.950 ;
        RECT 83.285 172.090 83.575 172.135 ;
        RECT 91.105 172.090 91.395 172.135 ;
        RECT 94.310 172.090 94.630 172.150 ;
        RECT 83.285 171.950 84.880 172.090 ;
        RECT 83.285 171.905 83.575 171.950 ;
        RECT 75.925 171.750 76.215 171.795 ;
        RECT 69.470 171.610 76.215 171.750 ;
        RECT 69.470 171.550 69.790 171.610 ;
        RECT 75.925 171.565 76.215 171.610 ;
        RECT 53.830 171.410 54.150 171.470 ;
        RECT 29.565 171.270 34.865 171.410 ;
        RECT 29.565 171.225 29.855 171.270 ;
        RECT 32.685 171.225 32.975 171.270 ;
        RECT 34.575 171.225 34.865 171.270 ;
        RECT 35.060 171.270 54.150 171.410 ;
        RECT 30.830 171.070 31.150 171.130 ;
        RECT 35.060 171.070 35.200 171.270 ;
        RECT 35.890 171.210 36.210 171.270 ;
        RECT 53.830 171.210 54.150 171.270 ;
        RECT 70.390 171.410 70.710 171.470 ;
        RECT 84.740 171.455 84.880 171.950 ;
        RECT 91.105 171.950 94.630 172.090 ;
        RECT 91.105 171.905 91.395 171.950 ;
        RECT 94.310 171.890 94.630 171.950 ;
        RECT 98.910 171.890 99.230 172.150 ;
        RECT 119.700 172.090 119.840 172.585 ;
        RECT 121.910 172.570 122.230 172.630 ;
        RECT 122.830 172.230 123.150 172.490 ;
        RECT 120.545 172.090 120.835 172.135 ;
        RECT 119.700 171.950 120.835 172.090 ;
        RECT 133.500 172.050 136.690 172.190 ;
        RECT 120.545 171.905 120.835 171.950 ;
        RECT 129.260 171.930 136.690 172.050 ;
        RECT 138.330 171.930 139.470 223.810 ;
        RECT 86.950 171.550 87.270 171.810 ;
        RECT 87.425 171.565 87.715 171.795 ;
        RECT 112.710 171.750 113.030 171.810 ;
        RECT 116.405 171.750 116.695 171.795 ;
        RECT 112.710 171.610 116.695 171.750 ;
        RECT 73.165 171.410 73.455 171.455 ;
        RECT 70.390 171.270 73.455 171.410 ;
        RECT 70.390 171.210 70.710 171.270 ;
        RECT 73.165 171.225 73.455 171.270 ;
        RECT 84.665 171.225 84.955 171.455 ;
        RECT 87.500 171.410 87.640 171.565 ;
        RECT 112.710 171.550 113.030 171.610 ;
        RECT 116.405 171.565 116.695 171.610 ;
        RECT 117.325 171.750 117.615 171.795 ;
        RECT 117.770 171.750 118.090 171.810 ;
        RECT 117.325 171.610 118.090 171.750 ;
        RECT 117.325 171.565 117.615 171.610 ;
        RECT 87.040 171.270 87.640 171.410 ;
        RECT 28.160 170.930 35.200 171.070 ;
        RECT 30.830 170.870 31.150 170.930 ;
        RECT 42.790 170.870 43.110 171.130 ;
        RECT 43.725 171.070 44.015 171.115 ;
        RECT 44.630 171.070 44.950 171.130 ;
        RECT 43.725 170.930 44.950 171.070 ;
        RECT 43.725 170.885 44.015 170.930 ;
        RECT 44.630 170.870 44.950 170.930 ;
        RECT 72.230 170.870 72.550 171.130 ;
        RECT 73.610 171.070 73.930 171.130 ;
        RECT 76.845 171.070 77.135 171.115 ;
        RECT 73.610 170.930 77.135 171.070 ;
        RECT 73.610 170.870 73.930 170.930 ;
        RECT 76.845 170.885 77.135 170.930 ;
        RECT 82.810 171.070 83.130 171.130 ;
        RECT 87.040 171.070 87.180 171.270 ;
        RECT 82.810 170.930 87.180 171.070 ;
        RECT 88.790 171.070 89.110 171.130 ;
        RECT 93.865 171.070 94.155 171.115 ;
        RECT 88.790 170.930 94.155 171.070 ;
        RECT 82.810 170.870 83.130 170.930 ;
        RECT 88.790 170.870 89.110 170.930 ;
        RECT 93.865 170.885 94.155 170.930 ;
        RECT 116.390 171.070 116.710 171.130 ;
        RECT 117.400 171.070 117.540 171.565 ;
        RECT 117.770 171.550 118.090 171.610 ;
        RECT 118.690 171.410 119.010 171.470 ;
        RECT 121.925 171.410 122.215 171.455 ;
        RECT 118.690 171.270 122.215 171.410 ;
        RECT 118.690 171.210 119.010 171.270 ;
        RECT 121.925 171.225 122.215 171.270 ;
        RECT 116.390 170.930 117.540 171.070 ;
        RECT 116.390 170.870 116.710 170.930 ;
        RECT 129.260 170.790 139.470 171.930 ;
        RECT 20.640 170.250 127.820 170.730 ;
        RECT 133.500 170.600 136.690 170.790 ;
        RECT 23.945 170.050 24.235 170.095 ;
        RECT 26.230 170.050 26.550 170.110 ;
        RECT 23.945 169.910 26.550 170.050 ;
        RECT 23.945 169.865 24.235 169.910 ;
        RECT 26.230 169.850 26.550 169.910 ;
        RECT 55.670 170.050 55.990 170.110 ;
        RECT 69.470 170.050 69.790 170.110 ;
        RECT 74.085 170.050 74.375 170.095 ;
        RECT 55.670 169.910 74.375 170.050 ;
        RECT 55.670 169.850 55.990 169.910 ;
        RECT 69.470 169.850 69.790 169.910 ;
        RECT 74.085 169.865 74.375 169.910 ;
        RECT 24.850 169.710 25.170 169.770 ;
        RECT 27.165 169.710 27.455 169.755 ;
        RECT 35.430 169.710 35.750 169.770 ;
        RECT 24.850 169.570 35.750 169.710 ;
        RECT 24.850 169.510 25.170 169.570 ;
        RECT 27.165 169.525 27.455 169.570 ;
        RECT 35.430 169.510 35.750 169.570 ;
        RECT 36.925 169.710 37.215 169.755 ;
        RECT 40.045 169.710 40.335 169.755 ;
        RECT 41.935 169.710 42.225 169.755 ;
        RECT 50.610 169.710 50.930 169.770 ;
        RECT 51.085 169.710 51.375 169.755 ;
        RECT 36.925 169.570 42.225 169.710 ;
        RECT 36.925 169.525 37.215 169.570 ;
        RECT 40.045 169.525 40.335 169.570 ;
        RECT 41.935 169.525 42.225 169.570 ;
        RECT 47.020 169.570 51.375 169.710 ;
        RECT 34.065 169.370 34.355 169.415 ;
        RECT 34.970 169.370 35.290 169.430 ;
        RECT 47.020 169.415 47.160 169.570 ;
        RECT 50.610 169.510 50.930 169.570 ;
        RECT 51.085 169.525 51.375 169.570 ;
        RECT 80.065 169.710 80.355 169.755 ;
        RECT 82.810 169.710 83.130 169.770 ;
        RECT 87.425 169.710 87.715 169.755 ;
        RECT 90.170 169.710 90.490 169.770 ;
        RECT 115.930 169.710 116.250 169.770 ;
        RECT 80.065 169.570 84.420 169.710 ;
        RECT 80.065 169.525 80.355 169.570 ;
        RECT 82.810 169.510 83.130 169.570 ;
        RECT 34.065 169.230 35.290 169.370 ;
        RECT 34.065 169.185 34.355 169.230 ;
        RECT 34.970 169.170 35.290 169.230 ;
        RECT 46.945 169.185 47.235 169.415 ;
        RECT 47.405 169.370 47.695 169.415 ;
        RECT 51.530 169.370 51.850 169.430 ;
        RECT 47.405 169.230 51.850 169.370 ;
        RECT 47.405 169.185 47.695 169.230 ;
        RECT 23.010 168.830 23.330 169.090 ;
        RECT 33.590 168.830 33.910 169.090 ;
        RECT 34.050 168.690 34.370 168.750 ;
        RECT 35.845 168.735 36.135 169.050 ;
        RECT 36.925 169.030 37.215 169.075 ;
        RECT 40.505 169.030 40.795 169.075 ;
        RECT 42.340 169.030 42.630 169.075 ;
        RECT 36.925 168.890 42.630 169.030 ;
        RECT 36.925 168.845 37.215 168.890 ;
        RECT 40.505 168.845 40.795 168.890 ;
        RECT 42.340 168.845 42.630 168.890 ;
        RECT 42.805 169.030 43.095 169.075 ;
        RECT 43.710 169.030 44.030 169.090 ;
        RECT 44.645 169.030 44.935 169.075 ;
        RECT 42.805 168.890 44.935 169.030 ;
        RECT 42.805 168.845 43.095 168.890 ;
        RECT 43.710 168.830 44.030 168.890 ;
        RECT 44.645 168.845 44.935 168.890 ;
        RECT 45.090 169.030 45.410 169.090 ;
        RECT 47.480 169.030 47.620 169.185 ;
        RECT 51.530 169.170 51.850 169.230 ;
        RECT 53.830 169.370 54.150 169.430 ;
        RECT 58.905 169.370 59.195 169.415 ;
        RECT 53.830 169.230 59.195 169.370 ;
        RECT 53.830 169.170 54.150 169.230 ;
        RECT 58.905 169.185 59.195 169.230 ;
        RECT 61.190 169.370 61.510 169.430 ;
        RECT 61.665 169.370 61.955 169.415 ;
        RECT 72.230 169.370 72.550 169.430 ;
        RECT 84.280 169.415 84.420 169.570 ;
        RECT 87.425 169.570 90.490 169.710 ;
        RECT 87.425 169.525 87.715 169.570 ;
        RECT 90.170 169.510 90.490 169.570 ;
        RECT 103.600 169.570 116.250 169.710 ;
        RECT 61.190 169.230 72.550 169.370 ;
        RECT 61.190 169.170 61.510 169.230 ;
        RECT 61.665 169.185 61.955 169.230 ;
        RECT 72.230 169.170 72.550 169.230 ;
        RECT 84.205 169.185 84.495 169.415 ;
        RECT 91.550 169.370 91.870 169.430 ;
        RECT 94.310 169.370 94.630 169.430 ;
        RECT 103.600 169.370 103.740 169.570 ;
        RECT 115.930 169.510 116.250 169.570 ;
        RECT 91.550 169.230 103.740 169.370 ;
        RECT 91.550 169.170 91.870 169.230 ;
        RECT 94.310 169.170 94.630 169.230 ;
        RECT 45.090 168.890 47.620 169.030 ;
        RECT 47.865 169.030 48.155 169.075 ;
        RECT 50.150 169.030 50.470 169.090 ;
        RECT 47.865 168.890 50.470 169.030 ;
        RECT 35.545 168.690 36.135 168.735 ;
        RECT 38.785 168.690 39.435 168.735 ;
        RECT 34.050 168.550 39.435 168.690 ;
        RECT 34.050 168.490 34.370 168.550 ;
        RECT 35.545 168.505 35.835 168.550 ;
        RECT 38.785 168.505 39.435 168.550 ;
        RECT 40.030 168.690 40.350 168.750 ;
        RECT 41.425 168.690 41.715 168.735 ;
        RECT 40.030 168.550 41.715 168.690 ;
        RECT 44.720 168.690 44.860 168.845 ;
        RECT 45.090 168.830 45.410 168.890 ;
        RECT 47.865 168.845 48.155 168.890 ;
        RECT 50.150 168.830 50.470 168.890 ;
        RECT 55.685 169.030 55.975 169.075 ;
        RECT 58.430 169.030 58.750 169.090 ;
        RECT 55.685 168.890 58.750 169.030 ;
        RECT 55.685 168.845 55.975 168.890 ;
        RECT 58.430 168.830 58.750 168.890 ;
        RECT 59.825 169.030 60.115 169.075 ;
        RECT 60.270 169.030 60.590 169.090 ;
        RECT 62.585 169.030 62.875 169.075 ;
        RECT 64.885 169.030 65.175 169.075 ;
        RECT 71.770 169.030 72.090 169.090 ;
        RECT 59.825 168.890 72.090 169.030 ;
        RECT 59.825 168.845 60.115 168.890 ;
        RECT 60.270 168.830 60.590 168.890 ;
        RECT 62.585 168.845 62.875 168.890 ;
        RECT 64.885 168.845 65.175 168.890 ;
        RECT 71.770 168.830 72.090 168.890 ;
        RECT 74.990 168.830 75.310 169.090 ;
        RECT 80.050 169.030 80.370 169.090 ;
        RECT 83.730 169.030 84.050 169.090 ;
        RECT 85.125 169.030 85.415 169.075 ;
        RECT 80.050 168.890 85.415 169.030 ;
        RECT 80.050 168.830 80.370 168.890 ;
        RECT 83.730 168.830 84.050 168.890 ;
        RECT 85.125 168.845 85.415 168.890 ;
        RECT 96.610 168.830 96.930 169.090 ;
        RECT 99.000 169.075 99.140 169.230 ;
        RECT 98.925 168.845 99.215 169.075 ;
        RECT 101.210 169.030 101.530 169.090 ;
        RECT 103.600 169.075 103.740 169.230 ;
        RECT 112.265 169.370 112.555 169.415 ;
        RECT 112.710 169.370 113.030 169.430 ;
        RECT 112.265 169.230 113.030 169.370 ;
        RECT 112.265 169.185 112.555 169.230 ;
        RECT 112.710 169.170 113.030 169.230 ;
        RECT 102.145 169.030 102.435 169.075 ;
        RECT 101.210 168.890 102.435 169.030 ;
        RECT 101.210 168.830 101.530 168.890 ;
        RECT 102.145 168.845 102.435 168.890 ;
        RECT 103.525 168.845 103.815 169.075 ;
        RECT 107.205 169.030 107.495 169.075 ;
        RECT 109.030 169.030 109.350 169.090 ;
        RECT 107.205 168.890 109.350 169.030 ;
        RECT 107.205 168.845 107.495 168.890 ;
        RECT 109.030 168.830 109.350 168.890 ;
        RECT 110.885 169.030 111.175 169.075 ;
        RECT 116.850 169.030 117.170 169.090 ;
        RECT 110.885 168.890 117.170 169.030 ;
        RECT 110.885 168.845 111.175 168.890 ;
        RECT 116.850 168.830 117.170 168.890 ;
        RECT 118.690 169.030 119.010 169.090 ;
        RECT 120.545 169.030 120.835 169.075 ;
        RECT 118.690 168.890 120.835 169.030 ;
        RECT 118.690 168.830 119.010 168.890 ;
        RECT 120.545 168.845 120.835 168.890 ;
        RECT 49.230 168.690 49.550 168.750 ;
        RECT 44.720 168.550 49.550 168.690 ;
        RECT 40.030 168.490 40.350 168.550 ;
        RECT 41.425 168.505 41.715 168.550 ;
        RECT 49.230 168.490 49.550 168.550 ;
        RECT 52.465 168.690 52.755 168.735 ;
        RECT 75.450 168.690 75.770 168.750 ;
        RECT 78.685 168.690 78.975 168.735 ;
        RECT 52.465 168.550 78.975 168.690 ;
        RECT 52.465 168.505 52.755 168.550 ;
        RECT 75.450 168.490 75.770 168.550 ;
        RECT 78.685 168.505 78.975 168.550 ;
        RECT 106.270 168.690 106.590 168.750 ;
        RECT 112.725 168.690 113.015 168.735 ;
        RECT 106.270 168.550 113.015 168.690 ;
        RECT 106.270 168.490 106.590 168.550 ;
        RECT 112.725 168.505 113.015 168.550 ;
        RECT 113.185 168.690 113.475 168.735 ;
        RECT 115.470 168.690 115.790 168.750 ;
        RECT 113.185 168.550 115.790 168.690 ;
        RECT 113.185 168.505 113.475 168.550 ;
        RECT 115.470 168.490 115.790 168.550 ;
        RECT 115.930 168.690 116.250 168.750 ;
        RECT 119.165 168.690 119.455 168.735 ;
        RECT 115.930 168.550 119.455 168.690 ;
        RECT 115.930 168.490 116.250 168.550 ;
        RECT 119.165 168.505 119.455 168.550 ;
        RECT 49.690 168.150 50.010 168.410 ;
        RECT 64.425 168.350 64.715 168.395 ;
        RECT 76.370 168.350 76.690 168.410 ;
        RECT 64.425 168.210 76.690 168.350 ;
        RECT 64.425 168.165 64.715 168.210 ;
        RECT 76.370 168.150 76.690 168.210 ;
        RECT 85.110 168.350 85.430 168.410 ;
        RECT 85.585 168.350 85.875 168.395 ;
        RECT 85.110 168.210 85.875 168.350 ;
        RECT 85.110 168.150 85.430 168.210 ;
        RECT 85.585 168.165 85.875 168.210 ;
        RECT 89.250 168.150 89.570 168.410 ;
        RECT 99.370 168.150 99.690 168.410 ;
        RECT 103.050 168.150 103.370 168.410 ;
        RECT 103.985 168.350 104.275 168.395 ;
        RECT 105.810 168.350 106.130 168.410 ;
        RECT 103.985 168.210 106.130 168.350 ;
        RECT 103.985 168.165 104.275 168.210 ;
        RECT 105.810 168.150 106.130 168.210 ;
        RECT 110.410 168.150 110.730 168.410 ;
        RECT 115.010 168.150 115.330 168.410 ;
        RECT 117.310 168.150 117.630 168.410 ;
        RECT 20.640 167.530 127.820 168.010 ;
        RECT 23.010 167.330 23.330 167.390 ;
        RECT 27.625 167.330 27.915 167.375 ;
        RECT 23.010 167.190 27.915 167.330 ;
        RECT 23.010 167.130 23.330 167.190 ;
        RECT 27.625 167.145 27.915 167.190 ;
        RECT 34.985 167.145 35.275 167.375 ;
        RECT 26.690 166.990 27.010 167.050 ;
        RECT 29.465 166.990 29.755 167.035 ;
        RECT 35.060 166.990 35.200 167.145 ;
        RECT 40.030 167.130 40.350 167.390 ;
        RECT 88.790 167.330 89.110 167.390 ;
        RECT 85.200 167.190 89.110 167.330 ;
        RECT 35.890 166.990 36.210 167.050 ;
        RECT 26.690 166.850 36.210 166.990 ;
        RECT 26.690 166.790 27.010 166.850 ;
        RECT 29.465 166.805 29.755 166.850 ;
        RECT 35.890 166.790 36.210 166.850 ;
        RECT 41.985 166.990 42.275 167.035 ;
        RECT 42.790 166.990 43.110 167.050 ;
        RECT 45.225 166.990 45.875 167.035 ;
        RECT 41.985 166.850 45.875 166.990 ;
        RECT 41.985 166.805 42.575 166.850 ;
        RECT 34.525 166.650 34.815 166.695 ;
        RECT 34.970 166.650 35.290 166.710 ;
        RECT 34.525 166.510 38.420 166.650 ;
        RECT 34.525 166.465 34.815 166.510 ;
        RECT 34.970 166.450 35.290 166.510 ;
        RECT 29.910 166.110 30.230 166.370 ;
        RECT 30.370 166.310 30.690 166.370 ;
        RECT 30.845 166.310 31.135 166.355 ;
        RECT 35.445 166.310 35.735 166.355 ;
        RECT 30.370 166.170 35.735 166.310 ;
        RECT 38.280 166.310 38.420 166.510 ;
        RECT 39.110 166.450 39.430 166.710 ;
        RECT 42.285 166.490 42.575 166.805 ;
        RECT 42.790 166.790 43.110 166.850 ;
        RECT 45.225 166.805 45.875 166.850 ;
        RECT 51.185 166.990 51.475 167.035 ;
        RECT 53.370 166.990 53.690 167.050 ;
        RECT 54.425 166.990 55.075 167.035 ;
        RECT 51.185 166.850 55.075 166.990 ;
        RECT 51.185 166.805 51.775 166.850 ;
        RECT 43.365 166.650 43.655 166.695 ;
        RECT 46.945 166.650 47.235 166.695 ;
        RECT 48.780 166.650 49.070 166.695 ;
        RECT 43.365 166.510 49.070 166.650 ;
        RECT 43.365 166.465 43.655 166.510 ;
        RECT 46.945 166.465 47.235 166.510 ;
        RECT 48.780 166.465 49.070 166.510 ;
        RECT 49.230 166.450 49.550 166.710 ;
        RECT 51.485 166.490 51.775 166.805 ;
        RECT 53.370 166.790 53.690 166.850 ;
        RECT 54.425 166.805 55.075 166.850 ;
        RECT 74.070 166.990 74.390 167.050 ;
        RECT 81.380 166.990 81.670 167.035 ;
        RECT 84.640 166.990 84.930 167.035 ;
        RECT 85.200 166.990 85.340 167.190 ;
        RECT 88.790 167.130 89.110 167.190 ;
        RECT 89.265 167.145 89.555 167.375 ;
        RECT 74.070 166.850 75.220 166.990 ;
        RECT 74.070 166.790 74.390 166.850 ;
        RECT 52.565 166.650 52.855 166.695 ;
        RECT 56.145 166.650 56.435 166.695 ;
        RECT 57.980 166.650 58.270 166.695 ;
        RECT 52.565 166.510 58.270 166.650 ;
        RECT 52.565 166.465 52.855 166.510 ;
        RECT 56.145 166.465 56.435 166.510 ;
        RECT 57.980 166.465 58.270 166.510 ;
        RECT 60.270 166.450 60.590 166.710 ;
        RECT 64.410 166.450 64.730 166.710 ;
        RECT 74.530 166.450 74.850 166.710 ;
        RECT 75.080 166.695 75.220 166.850 ;
        RECT 81.380 166.850 85.340 166.990 ;
        RECT 85.560 166.990 85.850 167.035 ;
        RECT 87.420 166.990 87.710 167.035 ;
        RECT 85.560 166.850 87.710 166.990 ;
        RECT 81.380 166.805 81.670 166.850 ;
        RECT 84.640 166.805 84.930 166.850 ;
        RECT 85.560 166.805 85.850 166.850 ;
        RECT 87.420 166.805 87.710 166.850 ;
        RECT 75.005 166.465 75.295 166.695 ;
        RECT 83.240 166.650 83.530 166.695 ;
        RECT 85.560 166.650 85.775 166.805 ;
        RECT 83.240 166.510 85.775 166.650 ;
        RECT 86.505 166.650 86.795 166.695 ;
        RECT 89.340 166.650 89.480 167.145 ;
        RECT 89.710 166.990 90.030 167.050 ;
        RECT 97.940 166.990 98.230 167.035 ;
        RECT 99.370 166.990 99.690 167.050 ;
        RECT 110.410 167.035 110.730 167.050 ;
        RECT 101.200 166.990 101.490 167.035 ;
        RECT 89.710 166.850 92.240 166.990 ;
        RECT 89.710 166.790 90.030 166.850 ;
        RECT 86.505 166.510 89.480 166.650 ;
        RECT 83.240 166.465 83.530 166.510 ;
        RECT 86.505 166.465 86.795 166.510 ;
        RECT 90.170 166.450 90.490 166.710 ;
        RECT 91.550 166.450 91.870 166.710 ;
        RECT 92.100 166.695 92.240 166.850 ;
        RECT 97.940 166.850 101.490 166.990 ;
        RECT 97.940 166.805 98.230 166.850 ;
        RECT 99.370 166.790 99.690 166.850 ;
        RECT 101.200 166.805 101.490 166.850 ;
        RECT 102.120 166.990 102.410 167.035 ;
        RECT 103.980 166.990 104.270 167.035 ;
        RECT 102.120 166.850 104.270 166.990 ;
        RECT 102.120 166.805 102.410 166.850 ;
        RECT 103.980 166.805 104.270 166.850 ;
        RECT 106.845 166.990 107.135 167.035 ;
        RECT 110.085 166.990 110.735 167.035 ;
        RECT 106.845 166.850 110.735 166.990 ;
        RECT 106.845 166.805 107.435 166.850 ;
        RECT 110.085 166.805 110.735 166.850 ;
        RECT 116.965 166.990 117.255 167.035 ;
        RECT 120.205 166.990 120.855 167.035 ;
        RECT 116.965 166.850 120.855 166.990 ;
        RECT 116.965 166.805 117.555 166.850 ;
        RECT 120.205 166.805 120.855 166.850 ;
        RECT 121.450 166.990 121.770 167.050 ;
        RECT 122.845 166.990 123.135 167.035 ;
        RECT 121.450 166.850 123.135 166.990 ;
        RECT 92.025 166.465 92.315 166.695 ;
        RECT 95.245 166.465 95.535 166.695 ;
        RECT 99.800 166.650 100.090 166.695 ;
        RECT 102.120 166.650 102.335 166.805 ;
        RECT 99.800 166.510 102.335 166.650 ;
        RECT 99.800 166.465 100.090 166.510 ;
        RECT 42.790 166.310 43.110 166.370 ;
        RECT 38.280 166.170 43.110 166.310 ;
        RECT 30.370 166.110 30.690 166.170 ;
        RECT 30.845 166.125 31.135 166.170 ;
        RECT 35.445 166.125 35.735 166.170 ;
        RECT 34.970 165.970 35.290 166.030 ;
        RECT 35.520 165.970 35.660 166.125 ;
        RECT 42.790 166.110 43.110 166.170 ;
        RECT 47.850 166.110 48.170 166.370 ;
        RECT 57.050 166.110 57.370 166.370 ;
        RECT 58.430 166.110 58.750 166.370 ;
        RECT 61.205 166.125 61.495 166.355 ;
        RECT 73.150 166.310 73.470 166.370 ;
        RECT 75.910 166.310 76.230 166.370 ;
        RECT 73.150 166.170 76.230 166.310 ;
        RECT 34.970 165.830 35.660 165.970 ;
        RECT 43.365 165.970 43.655 166.015 ;
        RECT 46.485 165.970 46.775 166.015 ;
        RECT 48.375 165.970 48.665 166.015 ;
        RECT 43.365 165.830 48.665 165.970 ;
        RECT 34.970 165.770 35.290 165.830 ;
        RECT 43.365 165.785 43.655 165.830 ;
        RECT 46.485 165.785 46.775 165.830 ;
        RECT 48.375 165.785 48.665 165.830 ;
        RECT 52.565 165.970 52.855 166.015 ;
        RECT 55.685 165.970 55.975 166.015 ;
        RECT 57.575 165.970 57.865 166.015 ;
        RECT 61.280 165.970 61.420 166.125 ;
        RECT 73.150 166.110 73.470 166.170 ;
        RECT 75.910 166.110 76.230 166.170 ;
        RECT 76.385 166.125 76.675 166.355 ;
        RECT 88.345 166.310 88.635 166.355 ;
        RECT 89.250 166.310 89.570 166.370 ;
        RECT 95.320 166.310 95.460 166.465 ;
        RECT 103.050 166.450 103.370 166.710 ;
        RECT 107.145 166.490 107.435 166.805 ;
        RECT 110.410 166.790 110.730 166.805 ;
        RECT 117.265 166.710 117.555 166.805 ;
        RECT 121.450 166.790 121.770 166.850 ;
        RECT 122.845 166.805 123.135 166.850 ;
        RECT 108.225 166.650 108.515 166.695 ;
        RECT 111.805 166.650 112.095 166.695 ;
        RECT 113.640 166.650 113.930 166.695 ;
        RECT 108.225 166.510 113.930 166.650 ;
        RECT 108.225 166.465 108.515 166.510 ;
        RECT 111.805 166.465 112.095 166.510 ;
        RECT 113.640 166.465 113.930 166.510 ;
        RECT 117.265 166.490 117.630 166.710 ;
        RECT 117.310 166.450 117.630 166.490 ;
        RECT 118.345 166.650 118.635 166.695 ;
        RECT 121.925 166.650 122.215 166.695 ;
        RECT 123.760 166.650 124.050 166.695 ;
        RECT 118.345 166.510 124.050 166.650 ;
        RECT 118.345 166.465 118.635 166.510 ;
        RECT 121.925 166.465 122.215 166.510 ;
        RECT 123.760 166.465 124.050 166.510 ;
        RECT 95.690 166.310 96.010 166.370 ;
        RECT 104.905 166.310 105.195 166.355 ;
        RECT 88.345 166.170 105.195 166.310 ;
        RECT 88.345 166.125 88.635 166.170 ;
        RECT 52.565 165.830 57.865 165.970 ;
        RECT 52.565 165.785 52.855 165.830 ;
        RECT 55.685 165.785 55.975 165.830 ;
        RECT 57.575 165.785 57.865 165.830 ;
        RECT 58.060 165.830 61.420 165.970 ;
        RECT 58.060 165.690 58.200 165.830 ;
        RECT 75.450 165.770 75.770 166.030 ;
        RECT 76.460 165.970 76.600 166.125 ;
        RECT 89.250 166.110 89.570 166.170 ;
        RECT 95.690 166.110 96.010 166.170 ;
        RECT 104.905 166.125 105.195 166.170 ;
        RECT 105.365 166.310 105.655 166.355 ;
        RECT 106.270 166.310 106.590 166.370 ;
        RECT 105.365 166.170 106.590 166.310 ;
        RECT 105.365 166.125 105.655 166.170 ;
        RECT 106.270 166.110 106.590 166.170 ;
        RECT 109.030 166.310 109.350 166.370 ;
        RECT 114.105 166.310 114.395 166.355 ;
        RECT 124.225 166.310 124.515 166.355 ;
        RECT 126.050 166.310 126.370 166.370 ;
        RECT 109.030 166.170 126.370 166.310 ;
        RECT 109.030 166.110 109.350 166.170 ;
        RECT 114.105 166.125 114.395 166.170 ;
        RECT 124.225 166.125 124.515 166.170 ;
        RECT 126.050 166.110 126.370 166.170 ;
        RECT 76.000 165.830 76.600 165.970 ;
        RECT 83.240 165.970 83.530 166.015 ;
        RECT 86.020 165.970 86.310 166.015 ;
        RECT 87.880 165.970 88.170 166.015 ;
        RECT 99.800 165.970 100.090 166.015 ;
        RECT 102.580 165.970 102.870 166.015 ;
        RECT 104.440 165.970 104.730 166.015 ;
        RECT 83.240 165.830 88.170 165.970 ;
        RECT 31.290 165.630 31.610 165.690 ;
        RECT 32.685 165.630 32.975 165.675 ;
        RECT 31.290 165.490 32.975 165.630 ;
        RECT 31.290 165.430 31.610 165.490 ;
        RECT 32.685 165.445 32.975 165.490 ;
        RECT 40.505 165.630 40.795 165.675 ;
        RECT 45.090 165.630 45.410 165.690 ;
        RECT 40.505 165.490 45.410 165.630 ;
        RECT 40.505 165.445 40.795 165.490 ;
        RECT 45.090 165.430 45.410 165.490 ;
        RECT 49.230 165.630 49.550 165.690 ;
        RECT 49.705 165.630 49.995 165.675 ;
        RECT 50.150 165.630 50.470 165.690 ;
        RECT 49.230 165.490 50.470 165.630 ;
        RECT 49.230 165.430 49.550 165.490 ;
        RECT 49.705 165.445 49.995 165.490 ;
        RECT 50.150 165.430 50.470 165.490 ;
        RECT 57.970 165.430 58.290 165.690 ;
        RECT 65.345 165.630 65.635 165.675 ;
        RECT 65.790 165.630 66.110 165.690 ;
        RECT 65.345 165.490 66.110 165.630 ;
        RECT 65.345 165.445 65.635 165.490 ;
        RECT 65.790 165.430 66.110 165.490 ;
        RECT 74.990 165.630 75.310 165.690 ;
        RECT 76.000 165.630 76.140 165.830 ;
        RECT 83.240 165.785 83.530 165.830 ;
        RECT 86.020 165.785 86.310 165.830 ;
        RECT 87.880 165.785 88.170 165.830 ;
        RECT 90.720 165.830 94.540 165.970 ;
        RECT 74.990 165.490 76.140 165.630 ;
        RECT 79.375 165.630 79.665 165.675 ;
        RECT 80.050 165.630 80.370 165.690 ;
        RECT 79.375 165.490 80.370 165.630 ;
        RECT 74.990 165.430 75.310 165.490 ;
        RECT 79.375 165.445 79.665 165.490 ;
        RECT 80.050 165.430 80.370 165.490 ;
        RECT 84.190 165.630 84.510 165.690 ;
        RECT 90.720 165.630 90.860 165.830 ;
        RECT 84.190 165.490 90.860 165.630 ;
        RECT 84.190 165.430 84.510 165.490 ;
        RECT 91.090 165.430 91.410 165.690 ;
        RECT 92.945 165.630 93.235 165.675 ;
        RECT 93.850 165.630 94.170 165.690 ;
        RECT 92.945 165.490 94.170 165.630 ;
        RECT 94.400 165.630 94.540 165.830 ;
        RECT 99.800 165.830 104.730 165.970 ;
        RECT 99.800 165.785 100.090 165.830 ;
        RECT 102.580 165.785 102.870 165.830 ;
        RECT 104.440 165.785 104.730 165.830 ;
        RECT 108.225 165.970 108.515 166.015 ;
        RECT 111.345 165.970 111.635 166.015 ;
        RECT 113.235 165.970 113.525 166.015 ;
        RECT 108.225 165.830 113.525 165.970 ;
        RECT 108.225 165.785 108.515 165.830 ;
        RECT 111.345 165.785 111.635 165.830 ;
        RECT 113.235 165.785 113.525 165.830 ;
        RECT 118.345 165.970 118.635 166.015 ;
        RECT 121.465 165.970 121.755 166.015 ;
        RECT 123.355 165.970 123.645 166.015 ;
        RECT 118.345 165.830 123.645 165.970 ;
        RECT 118.345 165.785 118.635 165.830 ;
        RECT 121.465 165.785 121.755 165.830 ;
        RECT 123.355 165.785 123.645 165.830 ;
        RECT 95.935 165.630 96.225 165.675 ;
        RECT 97.990 165.630 98.310 165.690 ;
        RECT 94.400 165.490 98.310 165.630 ;
        RECT 92.945 165.445 93.235 165.490 ;
        RECT 93.850 165.430 94.170 165.490 ;
        RECT 95.935 165.445 96.225 165.490 ;
        RECT 97.990 165.430 98.310 165.490 ;
        RECT 112.820 165.630 113.110 165.675 ;
        RECT 114.090 165.630 114.410 165.690 ;
        RECT 112.820 165.490 114.410 165.630 ;
        RECT 112.820 165.445 113.110 165.490 ;
        RECT 114.090 165.430 114.410 165.490 ;
        RECT 115.470 165.630 115.790 165.690 ;
        RECT 116.850 165.630 117.170 165.690 ;
        RECT 115.470 165.490 117.170 165.630 ;
        RECT 115.470 165.430 115.790 165.490 ;
        RECT 116.850 165.430 117.170 165.490 ;
        RECT 135.580 165.470 136.830 166.590 ;
        RECT 20.640 164.810 127.820 165.290 ;
        RECT 33.145 164.610 33.435 164.655 ;
        RECT 34.050 164.610 34.370 164.670 ;
        RECT 33.145 164.470 34.370 164.610 ;
        RECT 33.145 164.425 33.435 164.470 ;
        RECT 34.050 164.410 34.370 164.470 ;
        RECT 39.110 164.610 39.430 164.670 ;
        RECT 39.585 164.610 39.875 164.655 ;
        RECT 39.110 164.470 39.875 164.610 ;
        RECT 39.110 164.410 39.430 164.470 ;
        RECT 39.585 164.425 39.875 164.470 ;
        RECT 40.030 164.610 40.350 164.670 ;
        RECT 47.850 164.610 48.170 164.670 ;
        RECT 48.785 164.610 49.075 164.655 ;
        RECT 40.030 164.470 46.700 164.610 ;
        RECT 40.030 164.410 40.350 164.470 ;
        RECT 32.225 164.270 32.515 164.315 ;
        RECT 34.510 164.270 34.830 164.330 ;
        RECT 32.225 164.130 34.830 164.270 ;
        RECT 32.225 164.085 32.515 164.130 ;
        RECT 34.510 164.070 34.830 164.130 ;
        RECT 35.890 164.270 36.210 164.330 ;
        RECT 46.010 164.270 46.330 164.330 ;
        RECT 35.890 164.130 46.330 164.270 ;
        RECT 46.560 164.270 46.700 164.470 ;
        RECT 47.850 164.470 49.075 164.610 ;
        RECT 47.850 164.410 48.170 164.470 ;
        RECT 48.785 164.425 49.075 164.470 ;
        RECT 53.370 164.410 53.690 164.670 ;
        RECT 55.225 164.610 55.515 164.655 ;
        RECT 57.050 164.610 57.370 164.670 ;
        RECT 71.325 164.610 71.615 164.655 ;
        RECT 94.770 164.610 95.090 164.670 ;
        RECT 55.225 164.470 57.370 164.610 ;
        RECT 55.225 164.425 55.515 164.470 ;
        RECT 57.050 164.410 57.370 164.470 ;
        RECT 57.600 164.470 95.090 164.610 ;
        RECT 57.600 164.270 57.740 164.470 ;
        RECT 71.325 164.425 71.615 164.470 ;
        RECT 94.770 164.410 95.090 164.470 ;
        RECT 101.210 164.410 101.530 164.670 ;
        RECT 114.090 164.410 114.410 164.670 ;
        RECT 121.450 164.410 121.770 164.670 ;
        RECT 46.560 164.130 57.740 164.270 ;
        RECT 62.540 164.270 62.830 164.315 ;
        RECT 65.320 164.270 65.610 164.315 ;
        RECT 67.180 164.270 67.470 164.315 ;
        RECT 62.540 164.130 67.470 164.270 ;
        RECT 35.890 164.070 36.210 164.130 ;
        RECT 46.010 164.070 46.330 164.130 ;
        RECT 62.540 164.085 62.830 164.130 ;
        RECT 65.320 164.085 65.610 164.130 ;
        RECT 67.180 164.085 67.470 164.130 ;
        RECT 86.045 164.270 86.335 164.315 ;
        RECT 89.710 164.270 90.030 164.330 ;
        RECT 86.045 164.130 90.030 164.270 ;
        RECT 86.045 164.085 86.335 164.130 ;
        RECT 89.710 164.070 90.030 164.130 ;
        RECT 90.600 164.270 90.890 164.315 ;
        RECT 93.380 164.270 93.670 164.315 ;
        RECT 95.240 164.270 95.530 164.315 ;
        RECT 90.600 164.130 95.530 164.270 ;
        RECT 90.600 164.085 90.890 164.130 ;
        RECT 93.380 164.085 93.670 164.130 ;
        RECT 95.240 164.085 95.530 164.130 ;
        RECT 97.990 164.270 98.310 164.330 ;
        RECT 106.240 164.270 106.530 164.315 ;
        RECT 109.020 164.270 109.310 164.315 ;
        RECT 110.880 164.270 111.170 164.315 ;
        RECT 97.990 164.130 99.140 164.270 ;
        RECT 97.990 164.070 98.310 164.130 ;
        RECT 27.625 163.930 27.915 163.975 ;
        RECT 30.370 163.930 30.690 163.990 ;
        RECT 27.625 163.790 30.690 163.930 ;
        RECT 27.625 163.745 27.915 163.790 ;
        RECT 30.370 163.730 30.690 163.790 ;
        RECT 30.830 163.930 31.150 163.990 ;
        RECT 34.970 163.930 35.290 163.990 ;
        RECT 42.805 163.930 43.095 163.975 ;
        RECT 50.610 163.930 50.930 163.990 ;
        RECT 30.830 163.790 32.900 163.930 ;
        RECT 30.830 163.730 31.150 163.790 ;
        RECT 26.245 163.590 26.535 163.635 ;
        RECT 29.450 163.590 29.770 163.650 ;
        RECT 26.245 163.450 29.770 163.590 ;
        RECT 26.245 163.405 26.535 163.450 ;
        RECT 29.450 163.390 29.770 163.450 ;
        RECT 31.290 163.390 31.610 163.650 ;
        RECT 32.760 163.635 32.900 163.790 ;
        RECT 34.970 163.790 50.930 163.930 ;
        RECT 34.970 163.730 35.290 163.790 ;
        RECT 35.980 163.650 36.120 163.790 ;
        RECT 42.805 163.745 43.095 163.790 ;
        RECT 50.610 163.730 50.930 163.790 ;
        RECT 58.430 163.930 58.750 163.990 ;
        RECT 58.430 163.790 65.560 163.930 ;
        RECT 58.430 163.730 58.750 163.790 ;
        RECT 32.685 163.405 32.975 163.635 ;
        RECT 35.890 163.390 36.210 163.650 ;
        RECT 37.270 163.590 37.590 163.650 ;
        RECT 37.270 163.450 49.460 163.590 ;
        RECT 37.270 163.390 37.590 163.450 ;
        RECT 28.545 163.250 28.835 163.295 ;
        RECT 29.910 163.250 30.230 163.310 ;
        RECT 40.490 163.250 40.810 163.310 ;
        RECT 28.545 163.110 40.810 163.250 ;
        RECT 28.545 163.065 28.835 163.110 ;
        RECT 29.910 163.050 30.230 163.110 ;
        RECT 40.490 163.050 40.810 163.110 ;
        RECT 41.425 163.250 41.715 163.295 ;
        RECT 45.090 163.250 45.410 163.310 ;
        RECT 41.425 163.110 45.410 163.250 ;
        RECT 41.425 163.065 41.715 163.110 ;
        RECT 45.090 163.050 45.410 163.110 ;
        RECT 25.770 162.710 26.090 162.970 ;
        RECT 28.070 162.710 28.390 162.970 ;
        RECT 30.385 162.910 30.675 162.955 ;
        RECT 33.590 162.910 33.910 162.970 ;
        RECT 30.385 162.770 33.910 162.910 ;
        RECT 30.385 162.725 30.675 162.770 ;
        RECT 33.590 162.710 33.910 162.770 ;
        RECT 41.885 162.910 42.175 162.955 ;
        RECT 42.790 162.910 43.110 162.970 ;
        RECT 41.885 162.770 43.110 162.910 ;
        RECT 49.320 162.910 49.460 163.450 ;
        RECT 49.690 163.390 50.010 163.650 ;
        RECT 53.830 163.390 54.150 163.650 ;
        RECT 54.290 163.390 54.610 163.650 ;
        RECT 57.065 163.405 57.355 163.635 ;
        RECT 62.540 163.590 62.830 163.635 ;
        RECT 65.420 163.590 65.560 163.790 ;
        RECT 65.790 163.730 66.110 163.990 ;
        RECT 82.810 163.930 83.130 163.990 ;
        RECT 82.810 163.790 93.620 163.930 ;
        RECT 82.810 163.730 83.130 163.790 ;
        RECT 67.645 163.590 67.935 163.635 ;
        RECT 70.850 163.590 71.170 163.650 ;
        RECT 62.540 163.450 65.075 163.590 ;
        RECT 65.420 163.450 71.170 163.590 ;
        RECT 62.540 163.405 62.830 163.450 ;
        RECT 57.140 162.910 57.280 163.405 ;
        RECT 64.860 163.295 65.075 163.450 ;
        RECT 67.645 163.405 67.935 163.450 ;
        RECT 70.850 163.390 71.170 163.450 ;
        RECT 72.245 163.405 72.535 163.635 ;
        RECT 72.705 163.590 72.995 163.635 ;
        RECT 74.530 163.590 74.850 163.650 ;
        RECT 72.705 163.450 74.850 163.590 ;
        RECT 72.705 163.405 72.995 163.450 ;
        RECT 57.525 163.250 57.815 163.295 ;
        RECT 60.680 163.250 60.970 163.295 ;
        RECT 63.940 163.250 64.230 163.295 ;
        RECT 57.525 163.110 64.230 163.250 ;
        RECT 57.525 163.065 57.815 163.110 ;
        RECT 60.680 163.065 60.970 163.110 ;
        RECT 63.940 163.065 64.230 163.110 ;
        RECT 64.860 163.250 65.150 163.295 ;
        RECT 66.720 163.250 67.010 163.295 ;
        RECT 64.860 163.110 67.010 163.250 ;
        RECT 72.320 163.250 72.460 163.405 ;
        RECT 74.530 163.390 74.850 163.450 ;
        RECT 90.600 163.590 90.890 163.635 ;
        RECT 93.480 163.590 93.620 163.790 ;
        RECT 93.850 163.730 94.170 163.990 ;
        RECT 95.690 163.730 96.010 163.990 ;
        RECT 99.000 163.975 99.140 164.130 ;
        RECT 106.240 164.130 111.170 164.270 ;
        RECT 106.240 164.085 106.530 164.130 ;
        RECT 109.020 164.085 109.310 164.130 ;
        RECT 110.880 164.085 111.170 164.130 ;
        RECT 119.165 164.085 119.455 164.315 ;
        RECT 98.465 163.745 98.755 163.975 ;
        RECT 98.925 163.745 99.215 163.975 ;
        RECT 103.510 163.930 103.830 163.990 ;
        RECT 109.505 163.930 109.795 163.975 ;
        RECT 103.510 163.790 109.795 163.930 ;
        RECT 98.540 163.590 98.680 163.745 ;
        RECT 103.510 163.730 103.830 163.790 ;
        RECT 109.505 163.745 109.795 163.790 ;
        RECT 112.710 163.930 113.030 163.990 ;
        RECT 115.945 163.930 116.235 163.975 ;
        RECT 112.710 163.790 116.235 163.930 ;
        RECT 112.710 163.730 113.030 163.790 ;
        RECT 115.945 163.745 116.235 163.790 ;
        RECT 100.750 163.590 101.070 163.650 ;
        RECT 90.600 163.450 93.135 163.590 ;
        RECT 93.480 163.450 101.070 163.590 ;
        RECT 90.600 163.405 90.890 163.450 ;
        RECT 74.990 163.250 75.310 163.310 ;
        RECT 72.320 163.110 75.310 163.250 ;
        RECT 64.860 163.065 65.150 163.110 ;
        RECT 66.720 163.065 67.010 163.110 ;
        RECT 74.990 163.050 75.310 163.110 ;
        RECT 84.190 163.050 84.510 163.310 ;
        RECT 88.740 163.250 89.030 163.295 ;
        RECT 91.090 163.250 91.410 163.310 ;
        RECT 92.920 163.295 93.135 163.450 ;
        RECT 100.750 163.390 101.070 163.450 ;
        RECT 106.240 163.590 106.530 163.635 ;
        RECT 109.030 163.590 109.350 163.650 ;
        RECT 111.345 163.590 111.635 163.635 ;
        RECT 106.240 163.450 108.775 163.590 ;
        RECT 106.240 163.405 106.530 163.450 ;
        RECT 92.000 163.250 92.290 163.295 ;
        RECT 88.740 163.110 92.290 163.250 ;
        RECT 88.740 163.065 89.030 163.110 ;
        RECT 91.090 163.050 91.410 163.110 ;
        RECT 92.000 163.065 92.290 163.110 ;
        RECT 92.920 163.250 93.210 163.295 ;
        RECT 94.780 163.250 95.070 163.295 ;
        RECT 92.920 163.110 95.070 163.250 ;
        RECT 92.920 163.065 93.210 163.110 ;
        RECT 94.780 163.065 95.070 163.110 ;
        RECT 104.380 163.250 104.670 163.295 ;
        RECT 105.810 163.250 106.130 163.310 ;
        RECT 108.560 163.295 108.775 163.450 ;
        RECT 109.030 163.450 111.635 163.590 ;
        RECT 109.030 163.390 109.350 163.450 ;
        RECT 111.345 163.405 111.635 163.450 ;
        RECT 115.010 163.390 115.330 163.650 ;
        RECT 119.240 163.590 119.380 164.085 ;
        RECT 120.545 163.590 120.835 163.635 ;
        RECT 119.240 163.450 120.835 163.590 ;
        RECT 120.545 163.405 120.835 163.450 ;
        RECT 107.640 163.250 107.930 163.295 ;
        RECT 104.380 163.110 107.930 163.250 ;
        RECT 104.380 163.065 104.670 163.110 ;
        RECT 105.810 163.050 106.130 163.110 ;
        RECT 107.640 163.065 107.930 163.110 ;
        RECT 108.560 163.250 108.850 163.295 ;
        RECT 110.420 163.250 110.710 163.295 ;
        RECT 108.560 163.110 110.710 163.250 ;
        RECT 108.560 163.065 108.850 163.110 ;
        RECT 110.420 163.065 110.710 163.110 ;
        RECT 116.390 163.250 116.710 163.310 ;
        RECT 117.325 163.250 117.615 163.295 ;
        RECT 116.390 163.110 117.615 163.250 ;
        RECT 116.390 163.050 116.710 163.110 ;
        RECT 117.325 163.065 117.615 163.110 ;
        RECT 57.970 162.910 58.290 162.970 ;
        RECT 49.320 162.770 58.290 162.910 ;
        RECT 41.885 162.725 42.175 162.770 ;
        RECT 42.790 162.710 43.110 162.770 ;
        RECT 57.970 162.710 58.290 162.770 ;
        RECT 58.675 162.910 58.965 162.955 ;
        RECT 59.810 162.910 60.130 162.970 ;
        RECT 58.675 162.770 60.130 162.910 ;
        RECT 58.675 162.725 58.965 162.770 ;
        RECT 59.810 162.710 60.130 162.770 ;
        RECT 62.110 162.910 62.430 162.970 ;
        RECT 73.625 162.910 73.915 162.955 ;
        RECT 79.130 162.910 79.450 162.970 ;
        RECT 62.110 162.770 79.450 162.910 ;
        RECT 62.110 162.710 62.430 162.770 ;
        RECT 73.625 162.725 73.915 162.770 ;
        RECT 79.130 162.710 79.450 162.770 ;
        RECT 83.745 162.910 84.035 162.955 ;
        RECT 85.110 162.910 85.430 162.970 ;
        RECT 86.735 162.910 87.025 162.955 ;
        RECT 83.745 162.770 87.025 162.910 ;
        RECT 83.745 162.725 84.035 162.770 ;
        RECT 85.110 162.710 85.430 162.770 ;
        RECT 86.735 162.725 87.025 162.770 ;
        RECT 99.385 162.910 99.675 162.955 ;
        RECT 101.670 162.910 101.990 162.970 ;
        RECT 102.375 162.910 102.665 162.955 ;
        RECT 104.890 162.910 105.210 162.970 ;
        RECT 99.385 162.770 105.210 162.910 ;
        RECT 99.385 162.725 99.675 162.770 ;
        RECT 101.670 162.710 101.990 162.770 ;
        RECT 102.375 162.725 102.665 162.770 ;
        RECT 104.890 162.710 105.210 162.770 ;
        RECT 116.850 162.710 117.170 162.970 ;
        RECT 20.640 162.090 127.820 162.570 ;
        RECT 23.255 161.890 23.545 161.935 ;
        RECT 28.070 161.890 28.390 161.950 ;
        RECT 23.255 161.750 28.390 161.890 ;
        RECT 23.255 161.705 23.545 161.750 ;
        RECT 28.070 161.690 28.390 161.750 ;
        RECT 32.685 161.705 32.975 161.935 ;
        RECT 48.310 161.890 48.630 161.950 ;
        RECT 52.465 161.890 52.755 161.935 ;
        RECT 54.290 161.890 54.610 161.950 ;
        RECT 62.110 161.890 62.430 161.950 ;
        RECT 39.200 161.750 43.020 161.890 ;
        RECT 25.260 161.550 25.550 161.595 ;
        RECT 25.770 161.550 26.090 161.610 ;
        RECT 28.520 161.550 28.810 161.595 ;
        RECT 25.260 161.410 28.810 161.550 ;
        RECT 25.260 161.365 25.550 161.410 ;
        RECT 25.770 161.350 26.090 161.410 ;
        RECT 28.520 161.365 28.810 161.410 ;
        RECT 29.440 161.550 29.730 161.595 ;
        RECT 31.300 161.550 31.590 161.595 ;
        RECT 29.440 161.410 31.590 161.550 ;
        RECT 29.440 161.365 29.730 161.410 ;
        RECT 31.300 161.365 31.590 161.410 ;
        RECT 27.120 161.210 27.410 161.255 ;
        RECT 29.440 161.210 29.655 161.365 ;
        RECT 27.120 161.070 29.655 161.210 ;
        RECT 30.385 161.210 30.675 161.255 ;
        RECT 32.760 161.210 32.900 161.705 ;
        RECT 39.200 161.270 39.340 161.750 ;
        RECT 40.490 161.550 40.810 161.610 ;
        RECT 40.490 161.410 42.100 161.550 ;
        RECT 40.490 161.350 40.810 161.410 ;
        RECT 30.385 161.070 32.900 161.210 ;
        RECT 27.120 161.025 27.410 161.070 ;
        RECT 30.385 161.025 30.675 161.070 ;
        RECT 33.590 161.010 33.910 161.270 ;
        RECT 35.905 161.210 36.195 161.255 ;
        RECT 37.270 161.210 37.590 161.270 ;
        RECT 35.905 161.070 37.590 161.210 ;
        RECT 35.905 161.025 36.195 161.070 ;
        RECT 31.290 160.870 31.610 160.930 ;
        RECT 32.225 160.870 32.515 160.915 ;
        RECT 35.430 160.870 35.750 160.930 ;
        RECT 31.290 160.730 35.750 160.870 ;
        RECT 31.290 160.670 31.610 160.730 ;
        RECT 32.225 160.685 32.515 160.730 ;
        RECT 35.430 160.670 35.750 160.730 ;
        RECT 27.120 160.530 27.410 160.575 ;
        RECT 29.900 160.530 30.190 160.575 ;
        RECT 31.760 160.530 32.050 160.575 ;
        RECT 35.980 160.530 36.120 161.025 ;
        RECT 37.270 161.010 37.590 161.070 ;
        RECT 37.745 161.210 38.035 161.255 ;
        RECT 38.190 161.210 38.510 161.270 ;
        RECT 37.745 161.070 38.510 161.210 ;
        RECT 37.745 161.025 38.035 161.070 ;
        RECT 38.190 161.010 38.510 161.070 ;
        RECT 38.650 161.010 38.970 161.270 ;
        RECT 39.110 161.010 39.430 161.270 ;
        RECT 39.570 161.010 39.890 161.270 ;
        RECT 41.365 161.025 41.655 161.255 ;
        RECT 41.960 161.230 42.100 161.410 ;
        RECT 42.345 161.230 42.635 161.285 ;
        RECT 42.880 161.255 43.020 161.750 ;
        RECT 47.020 161.750 52.220 161.890 ;
        RECT 47.020 161.550 47.160 161.750 ;
        RECT 48.310 161.690 48.630 161.750 ;
        RECT 44.720 161.410 47.160 161.550 ;
        RECT 41.960 161.090 42.635 161.230 ;
        RECT 42.345 161.055 42.635 161.090 ;
        RECT 42.805 161.025 43.095 161.255 ;
        RECT 43.365 161.210 43.655 161.255 ;
        RECT 44.160 161.210 44.400 161.230 ;
        RECT 44.720 161.210 44.860 161.410 ;
        RECT 47.020 161.270 47.160 161.410 ;
        RECT 49.230 161.550 49.550 161.610 ;
        RECT 50.165 161.550 50.455 161.595 ;
        RECT 49.230 161.410 50.455 161.550 ;
        RECT 52.080 161.550 52.220 161.750 ;
        RECT 52.465 161.750 54.610 161.890 ;
        RECT 52.465 161.705 52.755 161.750 ;
        RECT 54.290 161.690 54.610 161.750 ;
        RECT 57.600 161.750 62.430 161.890 ;
        RECT 57.600 161.550 57.740 161.750 ;
        RECT 62.110 161.690 62.430 161.750 ;
        RECT 62.585 161.890 62.875 161.935 ;
        RECT 64.410 161.890 64.730 161.950 ;
        RECT 62.585 161.750 64.730 161.890 ;
        RECT 62.585 161.705 62.875 161.750 ;
        RECT 64.410 161.690 64.730 161.750 ;
        RECT 71.770 161.890 72.090 161.950 ;
        RECT 71.770 161.750 100.520 161.890 ;
        RECT 71.770 161.690 72.090 161.750 ;
        RECT 52.080 161.410 57.740 161.550 ;
        RECT 57.970 161.550 58.290 161.610 ;
        RECT 74.530 161.550 74.850 161.610 ;
        RECT 85.110 161.550 85.430 161.610 ;
        RECT 57.970 161.410 66.020 161.550 ;
        RECT 49.230 161.350 49.550 161.410 ;
        RECT 50.165 161.365 50.455 161.410 ;
        RECT 57.970 161.350 58.290 161.410 ;
        RECT 46.010 161.255 46.330 161.270 ;
        RECT 43.340 161.200 43.655 161.210 ;
        RECT 43.800 161.200 44.860 161.210 ;
        RECT 43.340 161.070 44.860 161.200 ;
        RECT 43.340 161.060 43.940 161.070 ;
        RECT 43.365 161.025 43.655 161.060 ;
        RECT 45.105 161.025 45.395 161.255 ;
        RECT 45.920 161.025 46.330 161.255 ;
        RECT 46.485 161.025 46.775 161.255 ;
        RECT 40.030 160.870 40.350 160.930 ;
        RECT 40.965 160.870 41.255 160.915 ;
        RECT 40.030 160.730 41.255 160.870 ;
        RECT 40.030 160.670 40.350 160.730 ;
        RECT 40.965 160.685 41.255 160.730 ;
        RECT 27.120 160.390 32.050 160.530 ;
        RECT 27.120 160.345 27.410 160.390 ;
        RECT 29.900 160.345 30.190 160.390 ;
        RECT 31.760 160.345 32.050 160.390 ;
        RECT 35.060 160.390 36.120 160.530 ;
        RECT 41.500 160.530 41.640 161.025 ;
        RECT 45.180 160.530 45.320 161.025 ;
        RECT 46.010 161.010 46.330 161.025 ;
        RECT 46.560 160.870 46.700 161.025 ;
        RECT 46.930 161.010 47.250 161.270 ;
        RECT 50.625 161.210 50.915 161.255 ;
        RECT 53.370 161.210 53.690 161.270 ;
        RECT 50.625 161.070 53.690 161.210 ;
        RECT 50.625 161.025 50.915 161.070 ;
        RECT 53.370 161.010 53.690 161.070 ;
        RECT 60.745 161.210 61.035 161.255 ;
        RECT 61.190 161.210 61.510 161.270 ;
        RECT 65.880 161.255 66.020 161.410 ;
        RECT 72.320 161.410 74.850 161.550 ;
        RECT 60.745 161.070 61.510 161.210 ;
        RECT 60.745 161.025 61.035 161.070 ;
        RECT 61.190 161.010 61.510 161.070 ;
        RECT 65.805 161.025 66.095 161.255 ;
        RECT 70.390 161.010 70.710 161.270 ;
        RECT 72.320 161.255 72.460 161.410 ;
        RECT 74.530 161.350 74.850 161.410 ;
        RECT 83.360 161.410 85.430 161.550 ;
        RECT 72.245 161.025 72.535 161.255 ;
        RECT 72.705 161.210 72.995 161.255 ;
        RECT 74.070 161.210 74.390 161.270 ;
        RECT 72.705 161.070 74.390 161.210 ;
        RECT 72.705 161.025 72.995 161.070 ;
        RECT 74.070 161.010 74.390 161.070 ;
        RECT 74.990 161.210 75.310 161.270 ;
        RECT 75.925 161.210 76.215 161.255 ;
        RECT 74.990 161.070 76.215 161.210 ;
        RECT 74.990 161.010 75.310 161.070 ;
        RECT 75.925 161.025 76.215 161.070 ;
        RECT 79.130 161.210 79.450 161.270 ;
        RECT 82.365 161.210 82.655 161.255 ;
        RECT 79.130 161.070 82.655 161.210 ;
        RECT 79.130 161.010 79.450 161.070 ;
        RECT 82.365 161.025 82.655 161.070 ;
        RECT 82.810 161.010 83.130 161.270 ;
        RECT 83.360 161.255 83.500 161.410 ;
        RECT 85.110 161.350 85.430 161.410 ;
        RECT 83.285 161.025 83.575 161.255 ;
        RECT 84.205 161.210 84.495 161.255 ;
        RECT 84.650 161.210 84.970 161.270 ;
        RECT 84.205 161.070 84.970 161.210 ;
        RECT 84.205 161.025 84.495 161.070 ;
        RECT 84.650 161.010 84.970 161.070 ;
        RECT 47.390 160.870 47.710 160.930 ;
        RECT 46.560 160.730 47.710 160.870 ;
        RECT 47.390 160.670 47.710 160.730 ;
        RECT 49.705 160.870 49.995 160.915 ;
        RECT 49.705 160.730 50.840 160.870 ;
        RECT 49.705 160.685 49.995 160.730 ;
        RECT 50.700 160.590 50.840 160.730 ;
        RECT 59.810 160.670 60.130 160.930 ;
        RECT 60.270 160.670 60.590 160.930 ;
        RECT 41.500 160.390 45.780 160.530 ;
        RECT 29.450 160.190 29.770 160.250 ;
        RECT 35.060 160.190 35.200 160.390 ;
        RECT 29.450 160.050 35.200 160.190 ;
        RECT 35.430 160.190 35.750 160.250 ;
        RECT 36.365 160.190 36.655 160.235 ;
        RECT 35.430 160.050 36.655 160.190 ;
        RECT 29.450 159.990 29.770 160.050 ;
        RECT 35.430 159.990 35.750 160.050 ;
        RECT 36.365 160.005 36.655 160.050 ;
        RECT 44.645 160.190 44.935 160.235 ;
        RECT 45.090 160.190 45.410 160.250 ;
        RECT 44.645 160.050 45.410 160.190 ;
        RECT 45.640 160.190 45.780 160.390 ;
        RECT 50.610 160.330 50.930 160.590 ;
        RECT 52.450 160.530 52.770 160.590 ;
        RECT 69.485 160.530 69.775 160.575 ;
        RECT 79.130 160.530 79.450 160.590 ;
        RECT 52.450 160.390 79.450 160.530 ;
        RECT 100.380 160.530 100.520 161.750 ;
        RECT 103.510 161.690 103.830 161.950 ;
        RECT 103.985 161.705 104.275 161.935 ;
        RECT 102.605 161.210 102.895 161.255 ;
        RECT 104.060 161.210 104.200 161.705 ;
        RECT 105.810 161.690 106.130 161.950 ;
        RECT 104.890 161.550 105.210 161.610 ;
        RECT 106.285 161.550 106.575 161.595 ;
        RECT 104.890 161.410 106.575 161.550 ;
        RECT 104.890 161.350 105.210 161.410 ;
        RECT 106.285 161.365 106.575 161.410 ;
        RECT 102.605 161.070 104.200 161.210 ;
        RECT 116.405 161.210 116.695 161.255 ;
        RECT 118.690 161.210 119.010 161.270 ;
        RECT 116.405 161.070 119.010 161.210 ;
        RECT 102.605 161.025 102.895 161.070 ;
        RECT 116.405 161.025 116.695 161.070 ;
        RECT 100.750 160.870 101.070 160.930 ;
        RECT 106.745 160.870 107.035 160.915 ;
        RECT 112.710 160.870 113.030 160.930 ;
        RECT 100.750 160.730 113.030 160.870 ;
        RECT 100.750 160.670 101.070 160.730 ;
        RECT 106.745 160.685 107.035 160.730 ;
        RECT 112.710 160.670 113.030 160.730 ;
        RECT 116.480 160.530 116.620 161.025 ;
        RECT 118.690 161.010 119.010 161.070 ;
        RECT 117.310 160.670 117.630 160.930 ;
        RECT 100.380 160.390 116.620 160.530 ;
        RECT 52.450 160.330 52.770 160.390 ;
        RECT 69.485 160.345 69.775 160.390 ;
        RECT 79.130 160.330 79.450 160.390 ;
        RECT 46.010 160.190 46.330 160.250 ;
        RECT 45.640 160.050 46.330 160.190 ;
        RECT 44.645 160.005 44.935 160.050 ;
        RECT 45.090 159.990 45.410 160.050 ;
        RECT 46.010 159.990 46.330 160.050 ;
        RECT 48.325 160.190 48.615 160.235 ;
        RECT 49.230 160.190 49.550 160.250 ;
        RECT 48.325 160.050 49.550 160.190 ;
        RECT 48.325 160.005 48.615 160.050 ;
        RECT 49.230 159.990 49.550 160.050 ;
        RECT 66.250 159.990 66.570 160.250 ;
        RECT 71.310 159.990 71.630 160.250 ;
        RECT 71.770 160.190 72.090 160.250 ;
        RECT 73.625 160.190 73.915 160.235 ;
        RECT 71.770 160.050 73.915 160.190 ;
        RECT 71.770 159.990 72.090 160.050 ;
        RECT 73.625 160.005 73.915 160.050 ;
        RECT 75.005 160.190 75.295 160.235 ;
        RECT 76.830 160.190 77.150 160.250 ;
        RECT 75.005 160.050 77.150 160.190 ;
        RECT 75.005 160.005 75.295 160.050 ;
        RECT 76.830 159.990 77.150 160.050 ;
        RECT 80.985 160.190 81.275 160.235 ;
        RECT 81.890 160.190 82.210 160.250 ;
        RECT 80.985 160.050 82.210 160.190 ;
        RECT 80.985 160.005 81.275 160.050 ;
        RECT 81.890 159.990 82.210 160.050 ;
        RECT 20.640 159.370 127.820 159.850 ;
        RECT 34.295 159.170 34.585 159.215 ;
        RECT 39.110 159.170 39.430 159.230 ;
        RECT 34.295 159.030 39.430 159.170 ;
        RECT 34.295 158.985 34.585 159.030 ;
        RECT 39.110 158.970 39.430 159.030 ;
        RECT 53.920 159.030 72.460 159.170 ;
        RECT 29.450 158.830 29.770 158.890 ;
        RECT 26.780 158.690 29.770 158.830 ;
        RECT 26.780 158.210 26.920 158.690 ;
        RECT 29.450 158.630 29.770 158.690 ;
        RECT 38.160 158.830 38.450 158.875 ;
        RECT 40.940 158.830 41.230 158.875 ;
        RECT 42.800 158.830 43.090 158.875 ;
        RECT 53.920 158.830 54.060 159.030 ;
        RECT 38.160 158.690 43.090 158.830 ;
        RECT 38.160 158.645 38.450 158.690 ;
        RECT 40.940 158.645 41.230 158.690 ;
        RECT 42.800 158.645 43.090 158.690 ;
        RECT 46.100 158.690 54.060 158.830 ;
        RECT 46.100 158.550 46.240 158.690 ;
        RECT 28.085 158.305 28.375 158.535 ;
        RECT 26.690 157.950 27.010 158.210 ;
        RECT 28.160 157.810 28.300 158.305 ;
        RECT 43.250 158.290 43.570 158.550 ;
        RECT 46.010 158.290 46.330 158.550 ;
        RECT 48.770 158.490 49.090 158.550 ;
        RECT 47.480 158.350 49.090 158.490 ;
        RECT 38.160 158.150 38.450 158.195 ;
        RECT 41.425 158.150 41.715 158.195 ;
        RECT 41.870 158.150 42.190 158.210 ;
        RECT 38.160 158.010 40.695 158.150 ;
        RECT 38.160 157.965 38.450 158.010 ;
        RECT 30.370 157.810 30.690 157.870 ;
        RECT 28.160 157.670 30.690 157.810 ;
        RECT 30.370 157.610 30.690 157.670 ;
        RECT 35.430 157.810 35.750 157.870 ;
        RECT 40.480 157.855 40.695 158.010 ;
        RECT 41.425 158.010 42.190 158.150 ;
        RECT 41.425 157.965 41.715 158.010 ;
        RECT 41.870 157.950 42.190 158.010 ;
        RECT 44.170 158.150 44.490 158.210 ;
        RECT 46.100 158.150 46.240 158.290 ;
        RECT 47.480 158.195 47.620 158.350 ;
        RECT 48.770 158.290 49.090 158.350 ;
        RECT 51.530 158.490 51.850 158.550 ;
        RECT 51.530 158.350 53.140 158.490 ;
        RECT 51.530 158.290 51.850 158.350 ;
        RECT 46.485 158.150 46.775 158.195 ;
        RECT 44.170 158.010 46.775 158.150 ;
        RECT 44.170 157.950 44.490 158.010 ;
        RECT 46.485 157.965 46.775 158.010 ;
        RECT 47.405 157.965 47.695 158.195 ;
        RECT 47.850 157.950 48.170 158.210 ;
        RECT 48.310 158.150 48.630 158.210 ;
        RECT 49.690 158.150 50.010 158.210 ;
        RECT 52.005 158.150 52.295 158.195 ;
        RECT 48.310 158.010 52.295 158.150 ;
        RECT 48.310 157.950 48.630 158.010 ;
        RECT 49.690 157.950 50.010 158.010 ;
        RECT 52.005 157.965 52.295 158.010 ;
        RECT 52.450 157.950 52.770 158.210 ;
        RECT 53.000 158.195 53.140 158.350 ;
        RECT 53.920 158.195 54.060 158.690 ;
        RECT 57.050 158.830 57.370 158.890 ;
        RECT 57.985 158.830 58.275 158.875 ;
        RECT 57.050 158.690 58.275 158.830 ;
        RECT 57.050 158.630 57.370 158.690 ;
        RECT 57.985 158.645 58.275 158.690 ;
        RECT 58.430 158.830 58.750 158.890 ;
        RECT 67.140 158.830 67.430 158.875 ;
        RECT 69.920 158.830 70.210 158.875 ;
        RECT 71.780 158.830 72.070 158.875 ;
        RECT 58.430 158.690 60.500 158.830 ;
        RECT 58.430 158.630 58.750 158.690 ;
        RECT 59.810 158.290 60.130 158.550 ;
        RECT 60.360 158.535 60.500 158.690 ;
        RECT 67.140 158.690 72.070 158.830 ;
        RECT 72.320 158.830 72.460 159.030 ;
        RECT 73.610 158.970 73.930 159.230 ;
        RECT 79.130 159.170 79.450 159.230 ;
        RECT 82.810 159.170 83.130 159.230 ;
        RECT 117.310 159.170 117.630 159.230 ;
        RECT 79.130 159.030 83.130 159.170 ;
        RECT 79.130 158.970 79.450 159.030 ;
        RECT 82.810 158.970 83.130 159.030 ;
        RECT 93.940 159.030 117.630 159.170 ;
        RECT 76.830 158.830 77.150 158.890 ;
        RECT 84.650 158.830 84.970 158.890 ;
        RECT 72.320 158.690 84.970 158.830 ;
        RECT 67.140 158.645 67.430 158.690 ;
        RECT 69.920 158.645 70.210 158.690 ;
        RECT 71.780 158.645 72.070 158.690 ;
        RECT 76.830 158.630 77.150 158.690 ;
        RECT 60.285 158.305 60.575 158.535 ;
        RECT 62.570 158.490 62.890 158.550 ;
        RECT 62.570 158.350 70.160 158.490 ;
        RECT 62.570 158.290 62.890 158.350 ;
        RECT 52.925 157.965 53.215 158.195 ;
        RECT 53.845 157.965 54.135 158.195 ;
        RECT 57.970 158.150 58.290 158.210 ;
        RECT 58.445 158.150 58.735 158.195 ;
        RECT 59.350 158.150 59.670 158.210 ;
        RECT 57.970 158.010 59.670 158.150 ;
        RECT 57.970 157.950 58.290 158.010 ;
        RECT 58.445 157.965 58.735 158.010 ;
        RECT 59.350 157.950 59.670 158.010 ;
        RECT 67.140 158.150 67.430 158.195 ;
        RECT 70.020 158.150 70.160 158.350 ;
        RECT 70.390 158.290 70.710 158.550 ;
        RECT 70.850 158.490 71.170 158.550 ;
        RECT 72.245 158.490 72.535 158.535 ;
        RECT 70.850 158.350 72.535 158.490 ;
        RECT 70.850 158.290 71.310 158.350 ;
        RECT 72.245 158.305 72.535 158.350 ;
        RECT 74.545 158.490 74.835 158.535 ;
        RECT 75.450 158.490 75.770 158.550 ;
        RECT 74.545 158.350 75.770 158.490 ;
        RECT 74.545 158.305 74.835 158.350 ;
        RECT 75.450 158.290 75.770 158.350 ;
        RECT 71.170 158.150 71.310 158.290 ;
        RECT 67.140 158.010 69.675 158.150 ;
        RECT 70.020 158.010 71.310 158.150 ;
        RECT 73.165 158.150 73.455 158.195 ;
        RECT 73.610 158.150 73.930 158.210 ;
        RECT 73.165 158.010 73.930 158.150 ;
        RECT 67.140 157.965 67.430 158.010 ;
        RECT 36.300 157.810 36.590 157.855 ;
        RECT 39.560 157.810 39.850 157.855 ;
        RECT 35.430 157.670 39.850 157.810 ;
        RECT 35.430 157.610 35.750 157.670 ;
        RECT 36.300 157.625 36.590 157.670 ;
        RECT 39.560 157.625 39.850 157.670 ;
        RECT 40.480 157.810 40.770 157.855 ;
        RECT 42.340 157.810 42.630 157.855 ;
        RECT 40.480 157.670 42.630 157.810 ;
        RECT 47.940 157.810 48.080 157.950 ;
        RECT 52.540 157.810 52.680 157.950 ;
        RECT 47.940 157.670 52.680 157.810 ;
        RECT 57.510 157.810 57.830 157.870 ;
        RECT 60.270 157.810 60.590 157.870 ;
        RECT 60.745 157.810 61.035 157.855 ;
        RECT 57.510 157.670 61.035 157.810 ;
        RECT 40.480 157.625 40.770 157.670 ;
        RECT 42.340 157.625 42.630 157.670 ;
        RECT 57.510 157.610 57.830 157.670 ;
        RECT 60.270 157.610 60.590 157.670 ;
        RECT 60.745 157.625 61.035 157.670 ;
        RECT 61.190 157.810 61.510 157.870 ;
        RECT 63.275 157.810 63.565 157.855 ;
        RECT 63.950 157.810 64.270 157.870 ;
        RECT 61.190 157.670 64.270 157.810 ;
        RECT 61.190 157.610 61.510 157.670 ;
        RECT 63.275 157.625 63.565 157.670 ;
        RECT 63.950 157.610 64.270 157.670 ;
        RECT 65.280 157.810 65.570 157.855 ;
        RECT 66.250 157.810 66.570 157.870 ;
        RECT 69.460 157.855 69.675 158.010 ;
        RECT 73.165 157.965 73.455 158.010 ;
        RECT 73.610 157.950 73.930 158.010 ;
        RECT 74.990 157.950 75.310 158.210 ;
        RECT 78.670 157.950 78.990 158.210 ;
        RECT 79.130 157.950 79.450 158.210 ;
        RECT 79.605 158.150 79.895 158.195 ;
        RECT 80.050 158.150 80.370 158.210 ;
        RECT 79.605 158.010 80.370 158.150 ;
        RECT 79.605 157.965 79.895 158.010 ;
        RECT 80.050 157.950 80.370 158.010 ;
        RECT 80.525 158.150 80.815 158.195 ;
        RECT 81.060 158.150 81.200 158.690 ;
        RECT 84.650 158.630 84.970 158.690 ;
        RECT 86.950 158.490 87.270 158.550 ;
        RECT 83.360 158.350 87.270 158.490 ;
        RECT 80.525 158.010 81.200 158.150 ;
        RECT 80.525 157.965 80.815 158.010 ;
        RECT 82.365 157.965 82.655 158.195 ;
        RECT 68.540 157.810 68.830 157.855 ;
        RECT 65.280 157.670 68.830 157.810 ;
        RECT 65.280 157.625 65.570 157.670 ;
        RECT 66.250 157.610 66.570 157.670 ;
        RECT 68.540 157.625 68.830 157.670 ;
        RECT 69.460 157.810 69.750 157.855 ;
        RECT 71.320 157.810 71.610 157.855 ;
        RECT 69.460 157.670 71.610 157.810 ;
        RECT 78.760 157.810 78.900 157.950 ;
        RECT 82.440 157.810 82.580 157.965 ;
        RECT 82.810 157.950 83.130 158.210 ;
        RECT 83.360 158.195 83.500 158.350 ;
        RECT 86.950 158.290 87.270 158.350 ;
        RECT 83.285 157.965 83.575 158.195 ;
        RECT 84.205 158.150 84.495 158.195 ;
        RECT 84.650 158.150 84.970 158.210 ;
        RECT 93.940 158.195 94.080 159.030 ;
        RECT 117.310 158.970 117.630 159.030 ;
        RECT 116.850 158.490 117.170 158.550 ;
        RECT 108.200 158.350 117.170 158.490 ;
        RECT 84.205 158.010 84.970 158.150 ;
        RECT 84.205 157.965 84.495 158.010 ;
        RECT 84.650 157.950 84.970 158.010 ;
        RECT 93.865 158.150 94.155 158.195 ;
        RECT 94.310 158.150 94.630 158.210 ;
        RECT 93.865 158.010 94.630 158.150 ;
        RECT 93.865 157.965 94.155 158.010 ;
        RECT 94.310 157.950 94.630 158.010 ;
        RECT 105.350 158.150 105.670 158.210 ;
        RECT 108.200 158.195 108.340 158.350 ;
        RECT 116.850 158.290 117.170 158.350 ;
        RECT 107.205 158.150 107.495 158.195 ;
        RECT 105.350 158.010 107.495 158.150 ;
        RECT 105.350 157.950 105.670 158.010 ;
        RECT 107.205 157.965 107.495 158.010 ;
        RECT 108.125 157.965 108.415 158.195 ;
        RECT 108.585 157.965 108.875 158.195 ;
        RECT 109.045 158.150 109.335 158.195 ;
        RECT 109.490 158.150 109.810 158.210 ;
        RECT 112.265 158.150 112.555 158.195 ;
        RECT 109.045 158.010 112.555 158.150 ;
        RECT 109.045 157.965 109.335 158.010 ;
        RECT 78.760 157.670 82.580 157.810 ;
        RECT 82.900 157.810 83.040 157.950 ;
        RECT 83.730 157.810 84.050 157.870 ;
        RECT 82.900 157.670 84.050 157.810 ;
        RECT 69.460 157.625 69.750 157.670 ;
        RECT 71.320 157.625 71.610 157.670 ;
        RECT 26.230 157.270 26.550 157.530 ;
        RECT 28.070 157.470 28.390 157.530 ;
        RECT 28.545 157.470 28.835 157.515 ;
        RECT 28.070 157.330 28.835 157.470 ;
        RECT 28.070 157.270 28.390 157.330 ;
        RECT 28.545 157.285 28.835 157.330 ;
        RECT 29.005 157.470 29.295 157.515 ;
        RECT 29.450 157.470 29.770 157.530 ;
        RECT 29.005 157.330 29.770 157.470 ;
        RECT 29.005 157.285 29.295 157.330 ;
        RECT 29.450 157.270 29.770 157.330 ;
        RECT 30.845 157.470 31.135 157.515 ;
        RECT 33.590 157.470 33.910 157.530 ;
        RECT 30.845 157.330 33.910 157.470 ;
        RECT 30.845 157.285 31.135 157.330 ;
        RECT 33.590 157.270 33.910 157.330 ;
        RECT 49.705 157.470 49.995 157.515 ;
        RECT 50.150 157.470 50.470 157.530 ;
        RECT 49.705 157.330 50.470 157.470 ;
        RECT 49.705 157.285 49.995 157.330 ;
        RECT 50.150 157.270 50.470 157.330 ;
        RECT 50.625 157.470 50.915 157.515 ;
        RECT 51.530 157.470 51.850 157.530 ;
        RECT 50.625 157.330 51.850 157.470 ;
        RECT 50.625 157.285 50.915 157.330 ;
        RECT 51.530 157.270 51.850 157.330 ;
        RECT 62.585 157.470 62.875 157.515 ;
        RECT 64.410 157.470 64.730 157.530 ;
        RECT 62.585 157.330 64.730 157.470 ;
        RECT 62.585 157.285 62.875 157.330 ;
        RECT 64.410 157.270 64.730 157.330 ;
        RECT 74.530 157.470 74.850 157.530 ;
        RECT 75.005 157.470 75.295 157.515 ;
        RECT 74.530 157.330 75.295 157.470 ;
        RECT 74.530 157.270 74.850 157.330 ;
        RECT 75.005 157.285 75.295 157.330 ;
        RECT 76.370 157.470 76.690 157.530 ;
        RECT 77.305 157.470 77.595 157.515 ;
        RECT 76.370 157.330 77.595 157.470 ;
        RECT 76.370 157.270 76.690 157.330 ;
        RECT 77.305 157.285 77.595 157.330 ;
        RECT 80.970 157.270 81.290 157.530 ;
        RECT 82.440 157.470 82.580 157.670 ;
        RECT 83.730 157.610 84.050 157.670 ;
        RECT 82.810 157.470 83.130 157.530 ;
        RECT 82.440 157.330 83.130 157.470 ;
        RECT 82.810 157.270 83.130 157.330 ;
        RECT 93.405 157.470 93.695 157.515 ;
        RECT 93.850 157.470 94.170 157.530 ;
        RECT 93.405 157.330 94.170 157.470 ;
        RECT 107.280 157.470 107.420 157.965 ;
        RECT 108.660 157.810 108.800 157.965 ;
        RECT 109.490 157.950 109.810 158.010 ;
        RECT 112.265 157.965 112.555 158.010 ;
        RECT 112.710 157.950 113.030 158.210 ;
        RECT 113.170 157.950 113.490 158.210 ;
        RECT 114.090 158.195 114.410 158.210 ;
        RECT 114.075 158.150 114.410 158.195 ;
        RECT 113.895 158.010 114.410 158.150 ;
        RECT 114.075 157.965 114.410 158.010 ;
        RECT 114.090 157.950 114.410 157.965 ;
        RECT 112.800 157.810 112.940 157.950 ;
        RECT 108.660 157.670 112.940 157.810 ;
        RECT 109.950 157.470 110.270 157.530 ;
        RECT 107.280 157.330 110.270 157.470 ;
        RECT 93.405 157.285 93.695 157.330 ;
        RECT 93.850 157.270 94.170 157.330 ;
        RECT 109.950 157.270 110.270 157.330 ;
        RECT 110.410 157.270 110.730 157.530 ;
        RECT 110.885 157.470 111.175 157.515 ;
        RECT 111.790 157.470 112.110 157.530 ;
        RECT 110.885 157.330 112.110 157.470 ;
        RECT 110.885 157.285 111.175 157.330 ;
        RECT 111.790 157.270 112.110 157.330 ;
        RECT 20.640 156.650 127.820 157.130 ;
        RECT 23.255 156.450 23.545 156.495 ;
        RECT 28.070 156.450 28.390 156.510 ;
        RECT 23.255 156.310 32.440 156.450 ;
        RECT 23.255 156.265 23.545 156.310 ;
        RECT 28.070 156.250 28.390 156.310 ;
        RECT 25.260 156.110 25.550 156.155 ;
        RECT 26.230 156.110 26.550 156.170 ;
        RECT 28.520 156.110 28.810 156.155 ;
        RECT 25.260 155.970 28.810 156.110 ;
        RECT 25.260 155.925 25.550 155.970 ;
        RECT 26.230 155.910 26.550 155.970 ;
        RECT 28.520 155.925 28.810 155.970 ;
        RECT 29.440 156.110 29.730 156.155 ;
        RECT 31.300 156.110 31.590 156.155 ;
        RECT 29.440 155.970 31.590 156.110 ;
        RECT 32.300 156.110 32.440 156.310 ;
        RECT 41.870 156.250 42.190 156.510 ;
        RECT 42.790 156.450 43.110 156.510 ;
        RECT 83.730 156.450 84.050 156.510 ;
        RECT 42.790 156.310 46.240 156.450 ;
        RECT 42.790 156.250 43.110 156.310 ;
        RECT 38.650 156.110 38.970 156.170 ;
        RECT 39.585 156.110 39.875 156.155 ;
        RECT 32.300 155.970 39.875 156.110 ;
        RECT 29.440 155.925 29.730 155.970 ;
        RECT 31.300 155.925 31.590 155.970 ;
        RECT 27.120 155.770 27.410 155.815 ;
        RECT 29.440 155.770 29.655 155.925 ;
        RECT 38.650 155.910 38.970 155.970 ;
        RECT 39.585 155.925 39.875 155.970 ;
        RECT 27.120 155.630 29.655 155.770 ;
        RECT 30.385 155.770 30.675 155.815 ;
        RECT 30.385 155.630 32.900 155.770 ;
        RECT 27.120 155.585 27.410 155.630 ;
        RECT 30.385 155.585 30.675 155.630 ;
        RECT 31.290 155.430 31.610 155.490 ;
        RECT 32.225 155.430 32.515 155.475 ;
        RECT 31.290 155.290 32.515 155.430 ;
        RECT 31.290 155.230 31.610 155.290 ;
        RECT 32.225 155.245 32.515 155.290 ;
        RECT 32.760 155.135 32.900 155.630 ;
        RECT 33.590 155.570 33.910 155.830 ;
        RECT 42.805 155.770 43.095 155.815 ;
        RECT 41.500 155.630 43.095 155.770 ;
        RECT 35.890 155.430 36.210 155.490 ;
        RECT 38.205 155.430 38.495 155.475 ;
        RECT 35.890 155.290 38.495 155.430 ;
        RECT 35.890 155.230 36.210 155.290 ;
        RECT 38.205 155.245 38.495 155.290 ;
        RECT 39.110 155.230 39.430 155.490 ;
        RECT 41.500 155.135 41.640 155.630 ;
        RECT 42.805 155.585 43.095 155.630 ;
        RECT 44.170 155.770 44.490 155.830 ;
        RECT 46.100 155.815 46.240 156.310 ;
        RECT 83.360 156.310 84.050 156.450 ;
        RECT 55.620 156.110 55.910 156.155 ;
        RECT 57.050 156.110 57.370 156.170 ;
        RECT 58.880 156.110 59.170 156.155 ;
        RECT 55.620 155.970 59.170 156.110 ;
        RECT 55.620 155.925 55.910 155.970 ;
        RECT 57.050 155.910 57.370 155.970 ;
        RECT 58.880 155.925 59.170 155.970 ;
        RECT 59.800 156.110 60.090 156.155 ;
        RECT 61.660 156.110 61.950 156.155 ;
        RECT 59.800 155.970 61.950 156.110 ;
        RECT 59.800 155.925 60.090 155.970 ;
        RECT 61.660 155.925 61.950 155.970 ;
        RECT 68.090 156.110 68.410 156.170 ;
        RECT 70.390 156.110 70.710 156.170 ;
        RECT 68.090 155.970 70.710 156.110 ;
        RECT 45.105 155.770 45.395 155.815 ;
        RECT 44.170 155.630 45.395 155.770 ;
        RECT 44.170 155.570 44.490 155.630 ;
        RECT 45.105 155.585 45.395 155.630 ;
        RECT 46.025 155.585 46.315 155.815 ;
        RECT 46.470 155.570 46.790 155.830 ;
        RECT 46.945 155.770 47.235 155.815 ;
        RECT 49.690 155.770 50.010 155.830 ;
        RECT 46.945 155.630 50.010 155.770 ;
        RECT 46.945 155.585 47.235 155.630 ;
        RECT 49.690 155.570 50.010 155.630 ;
        RECT 57.480 155.770 57.770 155.815 ;
        RECT 59.800 155.770 60.015 155.925 ;
        RECT 68.090 155.910 68.410 155.970 ;
        RECT 70.390 155.910 70.710 155.970 ;
        RECT 74.530 156.110 74.850 156.170 ;
        RECT 79.145 156.110 79.435 156.155 ;
        RECT 74.530 155.970 79.435 156.110 ;
        RECT 74.530 155.910 74.850 155.970 ;
        RECT 79.145 155.925 79.435 155.970 ;
        RECT 81.430 155.910 81.750 156.170 ;
        RECT 57.480 155.630 60.015 155.770 ;
        RECT 57.480 155.585 57.770 155.630 ;
        RECT 62.570 155.570 62.890 155.830 ;
        RECT 64.410 155.570 64.730 155.830 ;
        RECT 66.710 155.570 67.030 155.830 ;
        RECT 69.485 155.585 69.775 155.815 ;
        RECT 71.325 155.770 71.615 155.815 ;
        RECT 73.610 155.770 73.930 155.830 ;
        RECT 71.325 155.630 73.930 155.770 ;
        RECT 71.325 155.585 71.615 155.630 ;
        RECT 60.745 155.430 61.035 155.475 ;
        RECT 69.560 155.430 69.700 155.585 ;
        RECT 73.610 155.570 73.930 155.630 ;
        RECT 74.990 155.770 75.310 155.830 ;
        RECT 75.465 155.770 75.755 155.815 ;
        RECT 74.990 155.630 75.755 155.770 ;
        RECT 74.990 155.570 75.310 155.630 ;
        RECT 75.465 155.585 75.755 155.630 ;
        RECT 82.810 155.570 83.130 155.830 ;
        RECT 83.360 155.815 83.500 156.310 ;
        RECT 83.730 156.250 84.050 156.310 ;
        RECT 86.950 156.450 87.270 156.510 ;
        RECT 97.990 156.450 98.310 156.510 ;
        RECT 86.950 156.310 98.310 156.450 ;
        RECT 86.950 156.250 87.270 156.310 ;
        RECT 97.990 156.250 98.310 156.310 ;
        RECT 107.190 156.450 107.510 156.510 ;
        RECT 109.490 156.450 109.810 156.510 ;
        RECT 107.190 156.310 109.810 156.450 ;
        RECT 107.190 156.250 107.510 156.310 ;
        RECT 109.490 156.250 109.810 156.310 ;
        RECT 109.950 156.450 110.270 156.510 ;
        RECT 114.090 156.450 114.410 156.510 ;
        RECT 109.950 156.310 114.410 156.450 ;
        RECT 109.950 156.250 110.270 156.310 ;
        RECT 91.500 156.110 91.790 156.155 ;
        RECT 93.850 156.110 94.170 156.170 ;
        RECT 94.760 156.110 95.050 156.155 ;
        RECT 91.500 155.970 95.050 156.110 ;
        RECT 91.500 155.925 91.790 155.970 ;
        RECT 93.850 155.910 94.170 155.970 ;
        RECT 94.760 155.925 95.050 155.970 ;
        RECT 95.680 156.110 95.970 156.155 ;
        RECT 97.540 156.110 97.830 156.155 ;
        RECT 95.680 155.970 97.830 156.110 ;
        RECT 95.680 155.925 95.970 155.970 ;
        RECT 97.540 155.925 97.830 155.970 ;
        RECT 106.270 156.110 106.590 156.170 ;
        RECT 109.580 156.110 109.720 156.250 ;
        RECT 110.870 156.110 111.190 156.170 ;
        RECT 106.270 155.970 108.800 156.110 ;
        RECT 109.580 155.970 110.180 156.110 ;
        RECT 83.285 155.585 83.575 155.815 ;
        RECT 83.745 155.770 84.035 155.815 ;
        RECT 84.190 155.770 84.510 155.830 ;
        RECT 83.745 155.630 84.510 155.770 ;
        RECT 83.745 155.585 84.035 155.630 ;
        RECT 84.190 155.570 84.510 155.630 ;
        RECT 84.650 155.570 84.970 155.830 ;
        RECT 93.360 155.770 93.650 155.815 ;
        RECT 95.680 155.770 95.895 155.925 ;
        RECT 106.270 155.910 106.590 155.970 ;
        RECT 93.360 155.630 95.895 155.770 ;
        RECT 93.360 155.585 93.650 155.630 ;
        RECT 96.610 155.570 96.930 155.830 ;
        RECT 100.750 155.570 101.070 155.830 ;
        RECT 101.210 155.570 101.530 155.830 ;
        RECT 101.670 155.570 101.990 155.830 ;
        RECT 102.605 155.585 102.895 155.815 ;
        RECT 107.190 155.770 107.510 155.830 ;
        RECT 108.660 155.815 108.800 155.970 ;
        RECT 107.665 155.770 107.955 155.815 ;
        RECT 107.190 155.630 107.955 155.770 ;
        RECT 75.080 155.430 75.220 155.570 ;
        RECT 60.745 155.290 63.720 155.430 ;
        RECT 60.745 155.245 61.035 155.290 ;
        RECT 63.580 155.135 63.720 155.290 ;
        RECT 67.260 155.290 69.240 155.430 ;
        RECT 69.560 155.290 75.220 155.430 ;
        RECT 95.690 155.430 96.010 155.490 ;
        RECT 98.465 155.430 98.755 155.475 ;
        RECT 102.680 155.430 102.820 155.585 ;
        RECT 107.190 155.570 107.510 155.630 ;
        RECT 107.665 155.585 107.955 155.630 ;
        RECT 108.125 155.585 108.415 155.815 ;
        RECT 108.585 155.585 108.875 155.815 ;
        RECT 105.350 155.430 105.670 155.490 ;
        RECT 95.690 155.290 98.755 155.430 ;
        RECT 27.120 155.090 27.410 155.135 ;
        RECT 29.900 155.090 30.190 155.135 ;
        RECT 31.760 155.090 32.050 155.135 ;
        RECT 27.120 154.950 32.050 155.090 ;
        RECT 27.120 154.905 27.410 154.950 ;
        RECT 29.900 154.905 30.190 154.950 ;
        RECT 31.760 154.905 32.050 154.950 ;
        RECT 32.685 154.905 32.975 155.135 ;
        RECT 41.425 154.905 41.715 155.135 ;
        RECT 57.480 155.090 57.770 155.135 ;
        RECT 60.260 155.090 60.550 155.135 ;
        RECT 62.120 155.090 62.410 155.135 ;
        RECT 57.480 154.950 62.410 155.090 ;
        RECT 57.480 154.905 57.770 154.950 ;
        RECT 60.260 154.905 60.550 154.950 ;
        RECT 62.120 154.905 62.410 154.950 ;
        RECT 63.505 154.905 63.795 155.135 ;
        RECT 48.310 154.550 48.630 154.810 ;
        RECT 53.615 154.750 53.905 154.795 ;
        RECT 57.970 154.750 58.290 154.810 ;
        RECT 53.615 154.610 58.290 154.750 ;
        RECT 53.615 154.565 53.905 154.610 ;
        RECT 57.970 154.550 58.290 154.610 ;
        RECT 59.810 154.750 60.130 154.810 ;
        RECT 67.260 154.750 67.400 155.290 ;
        RECT 67.645 155.090 67.935 155.135 ;
        RECT 68.090 155.090 68.410 155.150 ;
        RECT 67.645 154.950 68.410 155.090 ;
        RECT 67.645 154.905 67.935 154.950 ;
        RECT 68.090 154.890 68.410 154.950 ;
        RECT 59.810 154.610 67.400 154.750 ;
        RECT 59.810 154.550 60.130 154.610 ;
        RECT 68.550 154.550 68.870 154.810 ;
        RECT 69.100 154.750 69.240 155.290 ;
        RECT 95.690 155.230 96.010 155.290 ;
        RECT 98.465 155.245 98.755 155.290 ;
        RECT 99.000 155.290 105.670 155.430 ;
        RECT 70.405 155.090 70.695 155.135 ;
        RECT 70.850 155.090 71.170 155.150 ;
        RECT 70.405 154.950 71.170 155.090 ;
        RECT 70.405 154.905 70.695 154.950 ;
        RECT 70.850 154.890 71.170 154.950 ;
        RECT 72.690 155.090 73.010 155.150 ;
        RECT 76.385 155.090 76.675 155.135 ;
        RECT 93.360 155.090 93.650 155.135 ;
        RECT 96.140 155.090 96.430 155.135 ;
        RECT 98.000 155.090 98.290 155.135 ;
        RECT 72.690 154.950 93.160 155.090 ;
        RECT 72.690 154.890 73.010 154.950 ;
        RECT 76.385 154.905 76.675 154.950 ;
        RECT 73.165 154.750 73.455 154.795 ;
        RECT 69.100 154.610 73.455 154.750 ;
        RECT 73.165 154.565 73.455 154.610 ;
        RECT 80.525 154.750 80.815 154.795 ;
        RECT 86.950 154.750 87.270 154.810 ;
        RECT 80.525 154.610 87.270 154.750 ;
        RECT 80.525 154.565 80.815 154.610 ;
        RECT 86.950 154.550 87.270 154.610 ;
        RECT 89.495 154.750 89.785 154.795 ;
        RECT 90.630 154.750 90.950 154.810 ;
        RECT 89.495 154.610 90.950 154.750 ;
        RECT 93.020 154.750 93.160 154.950 ;
        RECT 93.360 154.950 98.290 155.090 ;
        RECT 93.360 154.905 93.650 154.950 ;
        RECT 96.140 154.905 96.430 154.950 ;
        RECT 98.000 154.905 98.290 154.950 ;
        RECT 99.000 154.750 99.140 155.290 ;
        RECT 105.350 155.230 105.670 155.290 ;
        RECT 93.020 154.610 99.140 154.750 ;
        RECT 89.495 154.565 89.785 154.610 ;
        RECT 90.630 154.550 90.950 154.610 ;
        RECT 99.370 154.550 99.690 154.810 ;
        RECT 106.270 154.550 106.590 154.810 ;
        RECT 106.730 154.750 107.050 154.810 ;
        RECT 108.200 154.750 108.340 155.585 ;
        RECT 109.490 155.570 109.810 155.830 ;
        RECT 110.040 155.770 110.180 155.970 ;
        RECT 110.870 155.970 112.480 156.110 ;
        RECT 110.870 155.910 111.190 155.970 ;
        RECT 112.340 155.815 112.480 155.970 ;
        RECT 113.260 155.815 113.400 156.310 ;
        RECT 114.090 156.250 114.410 156.310 ;
        RECT 116.405 156.110 116.695 156.155 ;
        RECT 118.805 156.110 119.095 156.155 ;
        RECT 122.045 156.110 122.695 156.155 ;
        RECT 116.405 155.970 122.695 156.110 ;
        RECT 116.405 155.925 116.695 155.970 ;
        RECT 118.805 155.925 119.395 155.970 ;
        RECT 122.045 155.925 122.695 155.970 ;
        RECT 124.210 156.110 124.530 156.170 ;
        RECT 124.685 156.110 124.975 156.155 ;
        RECT 124.210 155.970 124.975 156.110 ;
        RECT 111.345 155.770 111.635 155.815 ;
        RECT 110.040 155.630 111.635 155.770 ;
        RECT 111.345 155.585 111.635 155.630 ;
        RECT 111.805 155.585 112.095 155.815 ;
        RECT 112.265 155.585 112.555 155.815 ;
        RECT 113.185 155.585 113.475 155.815 ;
        RECT 111.880 155.430 112.020 155.585 ;
        RECT 115.930 155.570 116.250 155.830 ;
        RECT 119.105 155.610 119.395 155.925 ;
        RECT 124.210 155.910 124.530 155.970 ;
        RECT 124.685 155.925 124.975 155.970 ;
        RECT 120.185 155.770 120.475 155.815 ;
        RECT 123.765 155.770 124.055 155.815 ;
        RECT 125.600 155.770 125.890 155.815 ;
        RECT 120.185 155.630 125.890 155.770 ;
        RECT 120.185 155.585 120.475 155.630 ;
        RECT 123.765 155.585 124.055 155.630 ;
        RECT 125.600 155.585 125.890 155.630 ;
        RECT 112.710 155.430 113.030 155.490 ;
        RECT 111.880 155.290 113.030 155.430 ;
        RECT 108.570 155.090 108.890 155.150 ;
        RECT 109.965 155.090 110.255 155.135 ;
        RECT 108.570 154.950 110.255 155.090 ;
        RECT 108.570 154.890 108.890 154.950 ;
        RECT 109.965 154.905 110.255 154.950 ;
        RECT 111.880 154.750 112.020 155.290 ;
        RECT 112.710 155.230 113.030 155.290 ;
        RECT 126.050 155.230 126.370 155.490 ;
        RECT 120.185 155.090 120.475 155.135 ;
        RECT 123.305 155.090 123.595 155.135 ;
        RECT 125.195 155.090 125.485 155.135 ;
        RECT 120.185 154.950 125.485 155.090 ;
        RECT 120.185 154.905 120.475 154.950 ;
        RECT 123.305 154.905 123.595 154.950 ;
        RECT 125.195 154.905 125.485 154.950 ;
        RECT 106.730 154.610 112.020 154.750 ;
        RECT 106.730 154.550 107.050 154.610 ;
        RECT 117.310 154.550 117.630 154.810 ;
        RECT 20.640 153.930 127.820 154.410 ;
        RECT 49.690 153.530 50.010 153.790 ;
        RECT 52.450 153.530 52.770 153.790 ;
        RECT 64.885 153.730 65.175 153.775 ;
        RECT 66.710 153.730 67.030 153.790 ;
        RECT 64.885 153.590 67.030 153.730 ;
        RECT 64.885 153.545 65.175 153.590 ;
        RECT 66.710 153.530 67.030 153.590 ;
        RECT 71.310 153.730 71.630 153.790 ;
        RECT 79.130 153.730 79.450 153.790 ;
        RECT 80.985 153.730 81.275 153.775 ;
        RECT 100.750 153.730 101.070 153.790 ;
        RECT 107.190 153.730 107.510 153.790 ;
        RECT 117.310 153.730 117.630 153.790 ;
        RECT 71.310 153.590 75.220 153.730 ;
        RECT 71.310 153.530 71.630 153.590 ;
        RECT 44.170 153.390 44.490 153.450 ;
        RECT 44.170 153.250 46.240 153.390 ;
        RECT 44.170 153.190 44.490 153.250 ;
        RECT 30.370 153.050 30.690 153.110 ;
        RECT 32.210 153.050 32.530 153.110 ;
        RECT 30.370 152.910 32.530 153.050 ;
        RECT 30.370 152.850 30.690 152.910 ;
        RECT 32.210 152.850 32.530 152.910 ;
        RECT 36.670 152.910 45.320 153.050 ;
        RECT 25.785 152.710 26.075 152.755 ;
        RECT 28.530 152.710 28.850 152.770 ;
        RECT 36.670 152.710 36.810 152.910 ;
        RECT 44.170 152.755 44.490 152.770 ;
        RECT 45.180 152.755 45.320 152.910 ;
        RECT 46.100 152.755 46.240 153.250 ;
        RECT 50.610 153.190 50.930 153.450 ;
        RECT 59.810 153.390 60.130 153.450 ;
        RECT 75.080 153.390 75.220 153.590 ;
        RECT 79.130 153.590 81.275 153.730 ;
        RECT 79.130 153.530 79.450 153.590 ;
        RECT 80.985 153.545 81.275 153.590 ;
        RECT 81.520 153.590 107.510 153.730 ;
        RECT 81.520 153.390 81.660 153.590 ;
        RECT 100.750 153.530 101.070 153.590 ;
        RECT 107.190 153.530 107.510 153.590 ;
        RECT 109.580 153.590 117.630 153.730 ;
        RECT 85.570 153.390 85.890 153.450 ;
        RECT 59.810 153.250 61.880 153.390 ;
        RECT 59.810 153.190 60.130 153.250 ;
        RECT 49.245 153.050 49.535 153.095 ;
        RECT 51.070 153.050 51.390 153.110 ;
        RECT 49.245 152.910 51.390 153.050 ;
        RECT 49.245 152.865 49.535 152.910 ;
        RECT 51.070 152.850 51.390 152.910 ;
        RECT 51.990 152.850 52.310 153.110 ;
        RECT 61.740 153.095 61.880 153.250 ;
        RECT 73.700 153.250 74.760 153.390 ;
        RECT 75.080 153.250 81.660 153.390 ;
        RECT 84.740 153.250 85.890 153.390 ;
        RECT 57.065 153.050 57.355 153.095 ;
        RECT 53.000 152.910 57.355 153.050 ;
        RECT 25.785 152.570 27.380 152.710 ;
        RECT 25.785 152.525 26.075 152.570 ;
        RECT 26.690 151.830 27.010 152.090 ;
        RECT 27.240 152.075 27.380 152.570 ;
        RECT 28.530 152.570 36.810 152.710 ;
        RECT 28.530 152.510 28.850 152.570 ;
        RECT 44.085 152.525 44.490 152.755 ;
        RECT 44.645 152.525 44.935 152.755 ;
        RECT 45.105 152.525 45.395 152.755 ;
        RECT 46.025 152.525 46.315 152.755 ;
        RECT 44.170 152.510 44.490 152.525 ;
        RECT 29.450 152.370 29.770 152.430 ;
        RECT 41.870 152.370 42.190 152.430 ;
        RECT 29.450 152.230 42.190 152.370 ;
        RECT 29.450 152.170 29.770 152.230 ;
        RECT 41.870 152.170 42.190 152.230 ;
        RECT 27.165 151.845 27.455 152.075 ;
        RECT 29.005 152.030 29.295 152.075 ;
        RECT 33.130 152.030 33.450 152.090 ;
        RECT 29.005 151.890 33.450 152.030 ;
        RECT 29.005 151.845 29.295 151.890 ;
        RECT 33.130 151.830 33.450 151.890 ;
        RECT 42.805 152.030 43.095 152.075 ;
        RECT 43.250 152.030 43.570 152.090 ;
        RECT 42.805 151.890 43.570 152.030 ;
        RECT 42.805 151.845 43.095 151.890 ;
        RECT 43.250 151.830 43.570 151.890 ;
        RECT 44.170 152.030 44.490 152.090 ;
        RECT 44.720 152.030 44.860 152.525 ;
        RECT 48.310 152.510 48.630 152.770 ;
        RECT 51.530 152.510 51.850 152.770 ;
        RECT 53.000 152.755 53.140 152.910 ;
        RECT 57.065 152.865 57.355 152.910 ;
        RECT 58.060 152.910 60.500 153.050 ;
        RECT 52.925 152.525 53.215 152.755 ;
        RECT 54.750 152.510 55.070 152.770 ;
        RECT 55.225 152.525 55.515 152.755 ;
        RECT 55.685 152.525 55.975 152.755 ;
        RECT 56.590 152.710 56.910 152.770 ;
        RECT 58.060 152.710 58.200 152.910 ;
        RECT 56.590 152.570 58.200 152.710 ;
        RECT 49.705 152.370 49.995 152.415 ;
        RECT 53.385 152.370 53.675 152.415 ;
        RECT 49.705 152.230 53.675 152.370 ;
        RECT 49.705 152.185 49.995 152.230 ;
        RECT 53.385 152.185 53.675 152.230 ;
        RECT 44.170 151.890 44.860 152.030 ;
        RECT 47.405 152.030 47.695 152.075 ;
        RECT 50.610 152.030 50.930 152.090 ;
        RECT 47.405 151.890 50.930 152.030 ;
        RECT 55.300 152.030 55.440 152.525 ;
        RECT 55.760 152.370 55.900 152.525 ;
        RECT 56.590 152.510 56.910 152.570 ;
        RECT 58.430 152.510 58.750 152.770 ;
        RECT 60.360 152.755 60.500 152.910 ;
        RECT 61.665 152.865 61.955 153.095 ;
        RECT 62.110 153.050 62.430 153.110 ;
        RECT 62.585 153.050 62.875 153.095 ;
        RECT 63.950 153.050 64.270 153.110 ;
        RECT 62.110 152.910 64.270 153.050 ;
        RECT 62.110 152.850 62.430 152.910 ;
        RECT 62.585 152.865 62.875 152.910 ;
        RECT 63.950 152.850 64.270 152.910 ;
        RECT 65.330 152.850 65.650 153.110 ;
        RECT 68.550 153.050 68.870 153.110 ;
        RECT 73.700 153.050 73.840 153.250 ;
        RECT 68.550 152.910 73.840 153.050 ;
        RECT 68.550 152.850 68.870 152.910 ;
        RECT 74.070 152.850 74.390 153.110 ;
        RECT 74.620 153.050 74.760 153.250 ;
        RECT 81.905 153.050 82.195 153.095 ;
        RECT 83.270 153.050 83.590 153.110 ;
        RECT 84.740 153.050 84.880 153.250 ;
        RECT 85.570 153.190 85.890 153.250 ;
        RECT 91.980 153.390 92.270 153.435 ;
        RECT 94.760 153.390 95.050 153.435 ;
        RECT 96.620 153.390 96.910 153.435 ;
        RECT 91.980 153.250 96.910 153.390 ;
        RECT 91.980 153.205 92.270 153.250 ;
        RECT 94.760 153.205 95.050 153.250 ;
        RECT 96.620 153.205 96.910 153.250 ;
        RECT 97.990 153.390 98.310 153.450 ;
        RECT 97.990 153.250 98.680 153.390 ;
        RECT 97.990 153.190 98.310 153.250 ;
        RECT 90.630 153.050 90.950 153.110 ;
        RECT 94.310 153.050 94.630 153.110 ;
        RECT 74.620 152.910 81.660 153.050 ;
        RECT 58.905 152.525 59.195 152.755 ;
        RECT 59.365 152.525 59.655 152.755 ;
        RECT 60.285 152.710 60.575 152.755 ;
        RECT 68.640 152.710 68.780 152.850 ;
        RECT 60.285 152.570 68.780 152.710 ;
        RECT 73.150 152.710 73.470 152.770 ;
        RECT 74.160 152.710 74.300 152.850 ;
        RECT 76.385 152.710 76.675 152.755 ;
        RECT 73.150 152.570 76.675 152.710 ;
        RECT 60.285 152.525 60.575 152.570 ;
        RECT 57.510 152.370 57.830 152.430 ;
        RECT 55.760 152.230 57.830 152.370 ;
        RECT 57.510 152.170 57.830 152.230 ;
        RECT 55.670 152.030 55.990 152.090 ;
        RECT 58.980 152.030 59.120 152.525 ;
        RECT 59.440 152.370 59.580 152.525 ;
        RECT 73.150 152.510 73.470 152.570 ;
        RECT 76.385 152.525 76.675 152.570 ;
        RECT 80.970 152.510 81.290 152.770 ;
        RECT 81.520 152.710 81.660 152.910 ;
        RECT 81.905 152.910 83.590 153.050 ;
        RECT 81.905 152.865 82.195 152.910 ;
        RECT 83.270 152.850 83.590 152.910 ;
        RECT 83.820 152.910 84.880 153.050 ;
        RECT 85.200 152.910 90.950 153.050 ;
        RECT 83.820 152.710 83.960 152.910 ;
        RECT 81.520 152.570 83.960 152.710 ;
        RECT 84.190 152.510 84.510 152.770 ;
        RECT 85.200 152.755 85.340 152.910 ;
        RECT 90.630 152.850 90.950 152.910 ;
        RECT 91.640 152.910 94.630 153.050 ;
        RECT 84.665 152.525 84.955 152.755 ;
        RECT 85.125 152.525 85.415 152.755 ;
        RECT 85.570 152.710 85.890 152.770 ;
        RECT 86.045 152.710 86.335 152.755 ;
        RECT 85.570 152.570 86.335 152.710 ;
        RECT 62.110 152.370 62.430 152.430 ;
        RECT 59.440 152.230 62.430 152.370 ;
        RECT 62.110 152.170 62.430 152.230 ;
        RECT 62.660 152.230 71.310 152.370 ;
        RECT 62.660 152.030 62.800 152.230 ;
        RECT 55.300 151.890 62.800 152.030 ;
        RECT 63.045 152.030 63.335 152.075 ;
        RECT 65.330 152.030 65.650 152.090 ;
        RECT 63.045 151.890 65.650 152.030 ;
        RECT 71.170 152.030 71.310 152.230 ;
        RECT 74.070 152.170 74.390 152.430 ;
        RECT 80.510 152.370 80.830 152.430 ;
        RECT 77.380 152.230 80.830 152.370 ;
        RECT 77.380 152.075 77.520 152.230 ;
        RECT 80.510 152.170 80.830 152.230 ;
        RECT 82.365 152.370 82.655 152.415 ;
        RECT 82.825 152.370 83.115 152.415 ;
        RECT 84.740 152.370 84.880 152.525 ;
        RECT 85.570 152.510 85.890 152.570 ;
        RECT 86.045 152.525 86.335 152.570 ;
        RECT 87.410 152.710 87.730 152.770 ;
        RECT 91.640 152.710 91.780 152.910 ;
        RECT 94.310 152.850 94.630 152.910 ;
        RECT 95.690 153.050 96.010 153.110 ;
        RECT 98.540 153.095 98.680 153.250 ;
        RECT 97.085 153.050 97.375 153.095 ;
        RECT 95.690 152.910 97.375 153.050 ;
        RECT 95.690 152.850 96.010 152.910 ;
        RECT 97.085 152.865 97.375 152.910 ;
        RECT 98.465 152.865 98.755 153.095 ;
        RECT 107.650 153.050 107.970 153.110 ;
        RECT 106.360 152.910 107.970 153.050 ;
        RECT 87.410 152.570 91.780 152.710 ;
        RECT 91.980 152.710 92.270 152.755 ;
        RECT 91.980 152.570 94.515 152.710 ;
        RECT 87.410 152.510 87.730 152.570 ;
        RECT 91.980 152.525 92.270 152.570 ;
        RECT 94.300 152.415 94.515 152.570 ;
        RECT 95.230 152.510 95.550 152.770 ;
        RECT 103.050 152.510 103.370 152.770 ;
        RECT 103.525 152.525 103.815 152.755 ;
        RECT 82.365 152.230 83.115 152.370 ;
        RECT 82.365 152.185 82.655 152.230 ;
        RECT 82.825 152.185 83.115 152.230 ;
        RECT 84.280 152.230 84.880 152.370 ;
        RECT 86.965 152.370 87.255 152.415 ;
        RECT 90.120 152.370 90.410 152.415 ;
        RECT 93.380 152.370 93.670 152.415 ;
        RECT 86.965 152.230 93.670 152.370 ;
        RECT 77.305 152.030 77.595 152.075 ;
        RECT 71.170 151.890 77.595 152.030 ;
        RECT 44.170 151.830 44.490 151.890 ;
        RECT 47.405 151.845 47.695 151.890 ;
        RECT 50.610 151.830 50.930 151.890 ;
        RECT 55.670 151.830 55.990 151.890 ;
        RECT 63.045 151.845 63.335 151.890 ;
        RECT 65.330 151.830 65.650 151.890 ;
        RECT 77.305 151.845 77.595 151.890 ;
        RECT 80.050 151.830 80.370 152.090 ;
        RECT 80.600 152.030 80.740 152.170 ;
        RECT 84.280 152.030 84.420 152.230 ;
        RECT 86.965 152.185 87.255 152.230 ;
        RECT 90.120 152.185 90.410 152.230 ;
        RECT 93.380 152.185 93.670 152.230 ;
        RECT 94.300 152.370 94.590 152.415 ;
        RECT 96.160 152.370 96.450 152.415 ;
        RECT 99.385 152.370 99.675 152.415 ;
        RECT 103.600 152.370 103.740 152.525 ;
        RECT 105.350 152.510 105.670 152.770 ;
        RECT 106.360 152.755 106.500 152.910 ;
        RECT 107.650 152.850 107.970 152.910 ;
        RECT 106.285 152.525 106.575 152.755 ;
        RECT 106.730 152.510 107.050 152.770 ;
        RECT 107.190 152.510 107.510 152.770 ;
        RECT 108.570 152.710 108.890 152.770 ;
        RECT 109.045 152.710 109.335 152.755 ;
        RECT 108.570 152.570 109.335 152.710 ;
        RECT 109.580 152.710 109.720 153.590 ;
        RECT 109.950 153.390 110.270 153.450 ;
        RECT 109.950 153.250 111.560 153.390 ;
        RECT 109.950 153.190 110.270 153.250 ;
        RECT 109.860 152.710 110.150 152.755 ;
        RECT 109.580 152.570 110.150 152.710 ;
        RECT 108.570 152.510 108.890 152.570 ;
        RECT 109.045 152.525 109.335 152.570 ;
        RECT 109.860 152.525 110.150 152.570 ;
        RECT 110.440 152.525 110.730 152.755 ;
        RECT 110.885 152.720 111.175 152.755 ;
        RECT 111.420 152.720 111.560 153.250 ;
        RECT 110.885 152.580 111.560 152.720 ;
        RECT 110.885 152.525 111.175 152.580 ;
        RECT 94.300 152.230 96.450 152.370 ;
        RECT 94.300 152.185 94.590 152.230 ;
        RECT 96.160 152.185 96.450 152.230 ;
        RECT 96.700 152.230 99.675 152.370 ;
        RECT 80.600 151.890 84.420 152.030 ;
        RECT 87.870 152.075 88.190 152.090 ;
        RECT 87.870 151.845 88.405 152.075 ;
        RECT 90.630 152.030 90.950 152.090 ;
        RECT 96.700 152.030 96.840 152.230 ;
        RECT 99.385 152.185 99.675 152.230 ;
        RECT 101.300 152.230 103.740 152.370 ;
        RECT 105.810 152.370 106.130 152.430 ;
        RECT 108.110 152.370 108.430 152.430 ;
        RECT 110.500 152.370 110.640 152.525 ;
        RECT 105.810 152.230 108.430 152.370 ;
        RECT 90.630 151.890 96.840 152.030 ;
        RECT 98.450 152.030 98.770 152.090 ;
        RECT 101.300 152.075 101.440 152.230 ;
        RECT 105.810 152.170 106.130 152.230 ;
        RECT 108.110 152.170 108.430 152.230 ;
        RECT 109.580 152.230 110.640 152.370 ;
        RECT 113.260 152.370 113.400 153.590 ;
        RECT 117.310 153.530 117.630 153.590 ;
        RECT 121.925 153.730 122.215 153.775 ;
        RECT 124.210 153.730 124.530 153.790 ;
        RECT 121.925 153.590 124.530 153.730 ;
        RECT 121.925 153.545 122.215 153.590 ;
        RECT 124.210 153.530 124.530 153.590 ;
        RECT 113.645 153.050 113.935 153.095 ;
        RECT 114.090 153.050 114.410 153.110 ;
        RECT 117.785 153.050 118.075 153.095 ;
        RECT 113.645 152.910 118.075 153.050 ;
        RECT 113.645 152.865 113.935 152.910 ;
        RECT 114.090 152.850 114.410 152.910 ;
        RECT 117.785 152.865 118.075 152.910 ;
        RECT 117.310 152.710 117.630 152.770 ;
        RECT 118.705 152.710 118.995 152.755 ;
        RECT 121.005 152.710 121.295 152.755 ;
        RECT 117.310 152.570 118.995 152.710 ;
        RECT 117.310 152.510 117.630 152.570 ;
        RECT 118.705 152.525 118.995 152.570 ;
        RECT 119.470 152.570 121.295 152.710 ;
        RECT 114.105 152.370 114.395 152.415 ;
        RECT 113.260 152.230 114.395 152.370 ;
        RECT 98.925 152.030 99.215 152.075 ;
        RECT 98.450 151.890 99.215 152.030 ;
        RECT 87.870 151.830 88.190 151.845 ;
        RECT 90.630 151.830 90.950 151.890 ;
        RECT 98.450 151.830 98.770 151.890 ;
        RECT 98.925 151.845 99.215 151.890 ;
        RECT 101.225 151.845 101.515 152.075 ;
        RECT 102.590 151.830 102.910 152.090 ;
        RECT 104.430 151.830 104.750 152.090 ;
        RECT 108.570 151.830 108.890 152.090 ;
        RECT 109.580 152.030 109.720 152.230 ;
        RECT 114.105 152.185 114.395 152.230 ;
        RECT 118.230 152.170 118.550 152.430 ;
        RECT 109.950 152.030 110.270 152.090 ;
        RECT 109.580 151.890 110.270 152.030 ;
        RECT 109.950 151.830 110.270 151.890 ;
        RECT 112.265 152.030 112.555 152.075 ;
        RECT 113.170 152.030 113.490 152.090 ;
        RECT 112.265 151.890 113.490 152.030 ;
        RECT 112.265 151.845 112.555 151.890 ;
        RECT 113.170 151.830 113.490 151.890 ;
        RECT 113.630 152.030 113.950 152.090 ;
        RECT 114.565 152.030 114.855 152.075 ;
        RECT 113.630 151.890 114.855 152.030 ;
        RECT 113.630 151.830 113.950 151.890 ;
        RECT 114.565 151.845 114.855 151.890 ;
        RECT 116.405 152.030 116.695 152.075 ;
        RECT 119.470 152.030 119.610 152.570 ;
        RECT 121.005 152.525 121.295 152.570 ;
        RECT 122.385 152.525 122.675 152.755 ;
        RECT 122.460 152.370 122.600 152.525 ;
        RECT 120.620 152.230 122.600 152.370 ;
        RECT 120.620 152.075 120.760 152.230 ;
        RECT 116.405 151.890 119.610 152.030 ;
        RECT 116.405 151.845 116.695 151.890 ;
        RECT 120.545 151.845 120.835 152.075 ;
        RECT 123.305 152.030 123.595 152.075 ;
        RECT 124.210 152.030 124.530 152.090 ;
        RECT 123.305 151.890 124.530 152.030 ;
        RECT 123.305 151.845 123.595 151.890 ;
        RECT 124.210 151.830 124.530 151.890 ;
        RECT 20.640 151.210 127.820 151.690 ;
        RECT 22.335 151.010 22.625 151.055 ;
        RECT 29.450 151.010 29.770 151.070 ;
        RECT 22.335 150.870 29.770 151.010 ;
        RECT 22.335 150.825 22.625 150.870 ;
        RECT 29.450 150.810 29.770 150.870 ;
        RECT 35.445 150.825 35.735 151.055 ;
        RECT 39.110 151.010 39.430 151.070 ;
        RECT 67.630 151.010 67.950 151.070 ;
        RECT 72.690 151.010 73.010 151.070 ;
        RECT 84.190 151.010 84.510 151.070 ;
        RECT 39.110 150.870 45.780 151.010 ;
        RECT 24.340 150.670 24.630 150.715 ;
        RECT 25.770 150.670 26.090 150.730 ;
        RECT 27.600 150.670 27.890 150.715 ;
        RECT 24.340 150.530 27.890 150.670 ;
        RECT 24.340 150.485 24.630 150.530 ;
        RECT 25.770 150.470 26.090 150.530 ;
        RECT 27.600 150.485 27.890 150.530 ;
        RECT 28.520 150.670 28.810 150.715 ;
        RECT 30.380 150.670 30.670 150.715 ;
        RECT 33.605 150.670 33.895 150.715 ;
        RECT 28.520 150.530 30.670 150.670 ;
        RECT 28.520 150.485 28.810 150.530 ;
        RECT 30.380 150.485 30.670 150.530 ;
        RECT 30.920 150.530 33.895 150.670 ;
        RECT 35.520 150.670 35.660 150.825 ;
        RECT 39.110 150.810 39.430 150.870 ;
        RECT 35.520 150.530 37.040 150.670 ;
        RECT 26.200 150.330 26.490 150.375 ;
        RECT 28.520 150.330 28.735 150.485 ;
        RECT 26.200 150.190 28.735 150.330 ;
        RECT 28.990 150.330 29.310 150.390 ;
        RECT 30.920 150.330 31.060 150.530 ;
        RECT 33.605 150.485 33.895 150.530 ;
        RECT 28.990 150.190 31.060 150.330 ;
        RECT 31.305 150.330 31.595 150.375 ;
        RECT 35.890 150.330 36.210 150.390 ;
        RECT 36.900 150.375 37.040 150.530 ;
        RECT 41.040 150.530 43.940 150.670 ;
        RECT 41.040 150.390 41.180 150.530 ;
        RECT 43.800 150.390 43.940 150.530 ;
        RECT 31.305 150.190 36.210 150.330 ;
        RECT 26.200 150.145 26.490 150.190 ;
        RECT 28.990 150.130 29.310 150.190 ;
        RECT 31.305 150.145 31.595 150.190 ;
        RECT 35.890 150.130 36.210 150.190 ;
        RECT 36.825 150.145 37.115 150.375 ;
        RECT 40.950 150.130 41.270 150.390 ;
        RECT 41.425 150.145 41.715 150.375 ;
        RECT 26.690 149.990 27.010 150.050 ;
        RECT 29.465 149.990 29.755 150.035 ;
        RECT 26.690 149.850 29.755 149.990 ;
        RECT 26.690 149.790 27.010 149.850 ;
        RECT 29.465 149.805 29.755 149.850 ;
        RECT 32.210 149.790 32.530 150.050 ;
        RECT 33.130 149.790 33.450 150.050 ;
        RECT 41.500 149.990 41.640 150.145 ;
        RECT 41.870 150.130 42.190 150.390 ;
        RECT 42.790 150.130 43.110 150.390 ;
        RECT 43.710 150.330 44.030 150.390 ;
        RECT 45.640 150.375 45.780 150.870 ;
        RECT 46.560 150.870 73.010 151.010 ;
        RECT 46.560 150.390 46.700 150.870 ;
        RECT 67.630 150.810 67.950 150.870 ;
        RECT 72.690 150.810 73.010 150.870 ;
        RECT 82.440 150.870 84.510 151.010 ;
        RECT 58.430 150.670 58.750 150.730 ;
        RECT 70.850 150.670 71.170 150.730 ;
        RECT 80.525 150.670 80.815 150.715 ;
        RECT 80.985 150.670 81.275 150.715 ;
        RECT 58.430 150.530 80.280 150.670 ;
        RECT 58.430 150.470 58.750 150.530 ;
        RECT 70.850 150.470 71.170 150.530 ;
        RECT 44.645 150.330 44.935 150.375 ;
        RECT 43.710 150.190 44.935 150.330 ;
        RECT 43.710 150.130 44.030 150.190 ;
        RECT 44.645 150.145 44.935 150.190 ;
        RECT 45.105 150.145 45.395 150.375 ;
        RECT 45.565 150.145 45.855 150.375 ;
        RECT 44.170 149.990 44.490 150.050 ;
        RECT 45.180 149.990 45.320 150.145 ;
        RECT 41.500 149.850 45.320 149.990 ;
        RECT 45.640 149.990 45.780 150.145 ;
        RECT 46.470 150.130 46.790 150.390 ;
        RECT 50.610 150.330 50.930 150.390 ;
        RECT 58.890 150.330 59.210 150.390 ;
        RECT 50.610 150.190 59.210 150.330 ;
        RECT 50.610 150.130 50.930 150.190 ;
        RECT 58.890 150.130 59.210 150.190 ;
        RECT 61.190 150.330 61.510 150.390 ;
        RECT 66.725 150.330 67.015 150.375 ;
        RECT 61.190 150.190 67.015 150.330 ;
        RECT 61.190 150.130 61.510 150.190 ;
        RECT 66.725 150.145 67.015 150.190 ;
        RECT 70.390 150.130 70.710 150.390 ;
        RECT 73.150 150.130 73.470 150.390 ;
        RECT 73.610 150.130 73.930 150.390 ;
        RECT 76.370 150.330 76.690 150.390 ;
        RECT 79.145 150.330 79.435 150.375 ;
        RECT 76.370 150.190 79.435 150.330 ;
        RECT 76.370 150.130 76.690 150.190 ;
        RECT 79.145 150.145 79.435 150.190 ;
        RECT 79.590 150.130 79.910 150.390 ;
        RECT 80.140 150.330 80.280 150.530 ;
        RECT 80.525 150.530 81.275 150.670 ;
        RECT 80.525 150.485 80.815 150.530 ;
        RECT 80.985 150.485 81.275 150.530 ;
        RECT 82.440 150.375 82.580 150.870 ;
        RECT 84.190 150.810 84.510 150.870 ;
        RECT 90.630 150.810 90.950 151.070 ;
        RECT 94.325 151.010 94.615 151.055 ;
        RECT 95.230 151.010 95.550 151.070 ;
        RECT 94.325 150.870 95.550 151.010 ;
        RECT 94.325 150.825 94.615 150.870 ;
        RECT 95.230 150.810 95.550 150.870 ;
        RECT 95.705 151.010 95.995 151.055 ;
        RECT 96.610 151.010 96.930 151.070 ;
        RECT 95.705 150.870 96.930 151.010 ;
        RECT 95.705 150.825 95.995 150.870 ;
        RECT 96.610 150.810 96.930 150.870 ;
        RECT 98.450 151.010 98.770 151.070 ;
        RECT 113.630 151.010 113.950 151.070 ;
        RECT 98.450 150.870 113.950 151.010 ;
        RECT 98.450 150.810 98.770 150.870 ;
        RECT 86.045 150.670 86.335 150.715 ;
        RECT 87.870 150.670 88.190 150.730 ;
        RECT 91.105 150.670 91.395 150.715 ;
        RECT 83.360 150.530 91.395 150.670 ;
        RECT 83.360 150.375 83.500 150.530 ;
        RECT 86.045 150.485 86.335 150.530 ;
        RECT 87.870 150.470 88.190 150.530 ;
        RECT 91.105 150.485 91.395 150.530 ;
        RECT 99.945 150.670 100.235 150.715 ;
        RECT 102.590 150.670 102.910 150.730 ;
        RECT 103.185 150.670 103.835 150.715 ;
        RECT 99.945 150.530 103.835 150.670 ;
        RECT 99.945 150.485 100.535 150.530 ;
        RECT 82.365 150.330 82.655 150.375 ;
        RECT 80.140 150.190 82.655 150.330 ;
        RECT 82.365 150.145 82.655 150.190 ;
        RECT 82.825 150.145 83.115 150.375 ;
        RECT 83.285 150.145 83.575 150.375 ;
        RECT 84.205 150.330 84.495 150.375 ;
        RECT 84.650 150.330 84.970 150.390 ;
        RECT 84.205 150.190 84.970 150.330 ;
        RECT 84.205 150.145 84.495 150.190 ;
        RECT 80.510 149.990 80.830 150.050 ;
        RECT 82.900 149.990 83.040 150.145 ;
        RECT 84.650 150.130 84.970 150.190 ;
        RECT 85.110 150.330 85.430 150.390 ;
        RECT 86.505 150.330 86.795 150.375 ;
        RECT 93.405 150.330 93.695 150.375 ;
        RECT 85.110 150.190 86.795 150.330 ;
        RECT 85.110 150.130 85.430 150.190 ;
        RECT 86.505 150.145 86.795 150.190 ;
        RECT 88.420 150.190 93.695 150.330 ;
        RECT 83.730 149.990 84.050 150.050 ;
        RECT 45.640 149.850 46.240 149.990 ;
        RECT 44.170 149.790 44.490 149.850 ;
        RECT 26.200 149.650 26.490 149.695 ;
        RECT 28.980 149.650 29.270 149.695 ;
        RECT 30.840 149.650 31.130 149.695 ;
        RECT 26.200 149.510 31.130 149.650 ;
        RECT 26.200 149.465 26.490 149.510 ;
        RECT 28.980 149.465 29.270 149.510 ;
        RECT 30.840 149.465 31.130 149.510 ;
        RECT 31.290 149.650 31.610 149.710 ;
        RECT 33.220 149.650 33.360 149.790 ;
        RECT 46.100 149.650 46.240 149.850 ;
        RECT 80.510 149.850 84.050 149.990 ;
        RECT 80.510 149.790 80.830 149.850 ;
        RECT 83.730 149.790 84.050 149.850 ;
        RECT 85.585 149.990 85.875 150.035 ;
        RECT 86.950 149.990 87.270 150.050 ;
        RECT 85.585 149.850 87.270 149.990 ;
        RECT 85.585 149.805 85.875 149.850 ;
        RECT 86.950 149.790 87.270 149.850 ;
        RECT 53.370 149.650 53.690 149.710 ;
        RECT 31.290 149.510 40.260 149.650 ;
        RECT 46.100 149.510 53.690 149.650 ;
        RECT 31.290 149.450 31.610 149.510 ;
        RECT 34.050 149.310 34.370 149.370 ;
        RECT 35.905 149.310 36.195 149.355 ;
        RECT 34.050 149.170 36.195 149.310 ;
        RECT 34.050 149.110 34.370 149.170 ;
        RECT 35.905 149.125 36.195 149.170 ;
        RECT 39.110 149.310 39.430 149.370 ;
        RECT 39.585 149.310 39.875 149.355 ;
        RECT 39.110 149.170 39.875 149.310 ;
        RECT 40.120 149.310 40.260 149.510 ;
        RECT 53.370 149.450 53.690 149.510 ;
        RECT 72.245 149.650 72.535 149.695 ;
        RECT 73.610 149.650 73.930 149.710 ;
        RECT 72.245 149.510 73.930 149.650 ;
        RECT 72.245 149.465 72.535 149.510 ;
        RECT 73.610 149.450 73.930 149.510 ;
        RECT 78.225 149.650 78.515 149.695 ;
        RECT 87.870 149.650 88.190 149.710 ;
        RECT 88.420 149.695 88.560 150.190 ;
        RECT 93.405 150.145 93.695 150.190 ;
        RECT 94.785 150.145 95.075 150.375 ;
        RECT 100.245 150.170 100.535 150.485 ;
        RECT 102.590 150.470 102.910 150.530 ;
        RECT 103.185 150.485 103.835 150.530 ;
        RECT 104.430 150.670 104.750 150.730 ;
        RECT 105.825 150.670 106.115 150.715 ;
        RECT 104.430 150.530 106.115 150.670 ;
        RECT 104.430 150.470 104.750 150.530 ;
        RECT 105.825 150.485 106.115 150.530 ;
        RECT 109.950 150.670 110.270 150.730 ;
        RECT 109.950 150.530 111.100 150.670 ;
        RECT 109.950 150.470 110.270 150.530 ;
        RECT 101.325 150.330 101.615 150.375 ;
        RECT 104.905 150.330 105.195 150.375 ;
        RECT 106.740 150.330 107.030 150.375 ;
        RECT 101.325 150.190 107.030 150.330 ;
        RECT 101.325 150.145 101.615 150.190 ;
        RECT 104.905 150.145 105.195 150.190 ;
        RECT 106.740 150.145 107.030 150.190 ;
        RECT 108.110 150.330 108.430 150.390 ;
        RECT 110.410 150.330 110.730 150.390 ;
        RECT 110.960 150.375 111.100 150.530 ;
        RECT 111.420 150.375 111.560 150.870 ;
        RECT 113.630 150.810 113.950 150.870 ;
        RECT 119.100 150.670 119.390 150.715 ;
        RECT 120.530 150.670 120.850 150.730 ;
        RECT 122.360 150.670 122.650 150.715 ;
        RECT 119.100 150.530 122.650 150.670 ;
        RECT 119.100 150.485 119.390 150.530 ;
        RECT 120.530 150.470 120.850 150.530 ;
        RECT 122.360 150.485 122.650 150.530 ;
        RECT 123.280 150.670 123.570 150.715 ;
        RECT 125.140 150.670 125.430 150.715 ;
        RECT 123.280 150.530 125.430 150.670 ;
        RECT 123.280 150.485 123.570 150.530 ;
        RECT 125.140 150.485 125.430 150.530 ;
        RECT 108.110 150.190 110.730 150.330 ;
        RECT 89.725 149.805 90.015 150.035 ;
        RECT 94.860 149.990 95.000 150.145 ;
        RECT 108.110 150.130 108.430 150.190 ;
        RECT 110.410 150.130 110.730 150.190 ;
        RECT 110.885 150.145 111.175 150.375 ;
        RECT 111.345 150.145 111.635 150.375 ;
        RECT 112.265 150.330 112.555 150.375 ;
        RECT 112.710 150.330 113.030 150.390 ;
        RECT 115.470 150.330 115.790 150.390 ;
        RECT 112.265 150.190 115.790 150.330 ;
        RECT 112.265 150.145 112.555 150.190 ;
        RECT 112.710 150.130 113.030 150.190 ;
        RECT 115.470 150.130 115.790 150.190 ;
        RECT 120.960 150.330 121.250 150.375 ;
        RECT 123.280 150.330 123.495 150.485 ;
        RECT 120.960 150.190 123.495 150.330 ;
        RECT 120.960 150.145 121.250 150.190 ;
        RECT 124.210 150.130 124.530 150.390 ;
        RECT 126.050 150.130 126.370 150.390 ;
        RECT 93.020 149.850 95.000 149.990 ;
        RECT 107.205 149.990 107.495 150.035 ;
        RECT 126.140 149.990 126.280 150.130 ;
        RECT 107.205 149.850 126.280 149.990 ;
        RECT 78.225 149.510 88.190 149.650 ;
        RECT 78.225 149.465 78.515 149.510 ;
        RECT 87.870 149.450 88.190 149.510 ;
        RECT 88.345 149.465 88.635 149.695 ;
        RECT 41.870 149.310 42.190 149.370 ;
        RECT 40.120 149.170 42.190 149.310 ;
        RECT 39.110 149.110 39.430 149.170 ;
        RECT 39.585 149.125 39.875 149.170 ;
        RECT 41.870 149.110 42.190 149.170 ;
        RECT 42.790 149.310 43.110 149.370 ;
        RECT 43.265 149.310 43.555 149.355 ;
        RECT 42.790 149.170 43.555 149.310 ;
        RECT 42.790 149.110 43.110 149.170 ;
        RECT 43.265 149.125 43.555 149.170 ;
        RECT 59.350 149.310 59.670 149.370 ;
        RECT 61.190 149.310 61.510 149.370 ;
        RECT 59.350 149.170 61.510 149.310 ;
        RECT 59.350 149.110 59.670 149.170 ;
        RECT 61.190 149.110 61.510 149.170 ;
        RECT 67.170 149.110 67.490 149.370 ;
        RECT 71.325 149.310 71.615 149.355 ;
        RECT 72.690 149.310 73.010 149.370 ;
        RECT 71.325 149.170 73.010 149.310 ;
        RECT 71.325 149.125 71.615 149.170 ;
        RECT 72.690 149.110 73.010 149.170 ;
        RECT 74.530 149.110 74.850 149.370 ;
        RECT 80.510 149.110 80.830 149.370 ;
        RECT 86.950 149.310 87.270 149.370 ;
        RECT 89.800 149.310 89.940 149.805 ;
        RECT 93.020 149.695 93.160 149.850 ;
        RECT 107.205 149.805 107.495 149.850 ;
        RECT 92.945 149.465 93.235 149.695 ;
        RECT 101.325 149.650 101.615 149.695 ;
        RECT 104.445 149.650 104.735 149.695 ;
        RECT 106.335 149.650 106.625 149.695 ;
        RECT 101.325 149.510 106.625 149.650 ;
        RECT 101.325 149.465 101.615 149.510 ;
        RECT 104.445 149.465 104.735 149.510 ;
        RECT 106.335 149.465 106.625 149.510 ;
        RECT 110.410 149.650 110.730 149.710 ;
        RECT 113.170 149.650 113.490 149.710 ;
        RECT 110.410 149.510 113.490 149.650 ;
        RECT 110.410 149.450 110.730 149.510 ;
        RECT 113.170 149.450 113.490 149.510 ;
        RECT 120.960 149.650 121.250 149.695 ;
        RECT 123.740 149.650 124.030 149.695 ;
        RECT 125.600 149.650 125.890 149.695 ;
        RECT 120.960 149.510 125.890 149.650 ;
        RECT 120.960 149.465 121.250 149.510 ;
        RECT 123.740 149.465 124.030 149.510 ;
        RECT 125.600 149.465 125.890 149.510 ;
        RECT 86.950 149.170 89.940 149.310 ;
        RECT 86.950 149.110 87.270 149.170 ;
        RECT 109.030 149.110 109.350 149.370 ;
        RECT 110.870 149.310 111.190 149.370 ;
        RECT 112.710 149.310 113.030 149.370 ;
        RECT 110.870 149.170 113.030 149.310 ;
        RECT 110.870 149.110 111.190 149.170 ;
        RECT 112.710 149.110 113.030 149.170 ;
        RECT 114.090 149.310 114.410 149.370 ;
        RECT 117.095 149.310 117.385 149.355 ;
        RECT 118.230 149.310 118.550 149.370 ;
        RECT 114.090 149.170 118.550 149.310 ;
        RECT 114.090 149.110 114.410 149.170 ;
        RECT 117.095 149.125 117.385 149.170 ;
        RECT 118.230 149.110 118.550 149.170 ;
        RECT 20.640 148.490 127.820 148.970 ;
        RECT 25.770 148.090 26.090 148.350 ;
        RECT 26.935 148.290 27.225 148.335 ;
        RECT 31.290 148.290 31.610 148.350 ;
        RECT 26.935 148.150 31.610 148.290 ;
        RECT 26.935 148.105 27.225 148.150 ;
        RECT 31.290 148.090 31.610 148.150 ;
        RECT 51.990 148.090 52.310 148.350 ;
        RECT 53.370 148.290 53.690 148.350 ;
        RECT 55.670 148.290 55.990 148.350 ;
        RECT 53.370 148.150 55.990 148.290 ;
        RECT 53.370 148.090 53.690 148.150 ;
        RECT 55.670 148.090 55.990 148.150 ;
        RECT 71.770 148.290 72.090 148.350 ;
        RECT 71.770 148.150 74.300 148.290 ;
        RECT 71.770 148.090 72.090 148.150 ;
        RECT 30.800 147.950 31.090 147.995 ;
        RECT 33.580 147.950 33.870 147.995 ;
        RECT 35.440 147.950 35.730 147.995 ;
        RECT 30.800 147.810 35.730 147.950 ;
        RECT 30.800 147.765 31.090 147.810 ;
        RECT 33.580 147.765 33.870 147.810 ;
        RECT 35.440 147.765 35.730 147.810 ;
        RECT 51.085 147.950 51.375 147.995 ;
        RECT 54.290 147.950 54.610 148.010 ;
        RECT 51.085 147.810 54.610 147.950 ;
        RECT 51.085 147.765 51.375 147.810 ;
        RECT 54.290 147.750 54.610 147.810 ;
        RECT 54.750 147.950 55.070 148.010 ;
        RECT 58.430 147.950 58.750 148.010 ;
        RECT 54.750 147.810 58.750 147.950 ;
        RECT 54.750 147.750 55.070 147.810 ;
        RECT 34.050 147.410 34.370 147.670 ;
        RECT 35.890 147.410 36.210 147.670 ;
        RECT 44.170 147.610 44.490 147.670 ;
        RECT 41.500 147.470 44.490 147.610 ;
        RECT 26.230 147.070 26.550 147.330 ;
        RECT 30.800 147.270 31.090 147.315 ;
        RECT 30.800 147.130 33.335 147.270 ;
        RECT 30.800 147.085 31.090 147.130 ;
        RECT 28.940 146.930 29.230 146.975 ;
        RECT 30.370 146.930 30.690 146.990 ;
        RECT 33.120 146.975 33.335 147.130 ;
        RECT 40.950 147.070 41.270 147.330 ;
        RECT 41.500 147.315 41.640 147.470 ;
        RECT 44.170 147.410 44.490 147.470 ;
        RECT 52.910 147.410 53.230 147.670 ;
        RECT 41.425 147.085 41.715 147.315 ;
        RECT 41.870 147.070 42.190 147.330 ;
        RECT 42.805 147.270 43.095 147.315 ;
        RECT 46.470 147.270 46.790 147.330 ;
        RECT 42.805 147.130 46.790 147.270 ;
        RECT 42.805 147.085 43.095 147.130 ;
        RECT 46.470 147.070 46.790 147.130 ;
        RECT 50.150 147.270 50.470 147.330 ;
        RECT 55.300 147.315 55.440 147.810 ;
        RECT 58.430 147.750 58.750 147.810 ;
        RECT 68.205 147.950 68.495 147.995 ;
        RECT 71.325 147.950 71.615 147.995 ;
        RECT 73.215 147.950 73.505 147.995 ;
        RECT 68.205 147.810 73.505 147.950 ;
        RECT 74.160 147.950 74.300 148.150 ;
        RECT 82.810 148.090 83.130 148.350 ;
        RECT 108.125 148.105 108.415 148.335 ;
        RECT 108.585 148.290 108.875 148.335 ;
        RECT 108.585 148.150 110.640 148.290 ;
        RECT 108.585 148.105 108.875 148.150 ;
        RECT 101.210 147.950 101.530 148.010 ;
        RECT 74.160 147.810 101.530 147.950 ;
        RECT 108.200 147.950 108.340 148.105 ;
        RECT 109.950 147.950 110.270 148.010 ;
        RECT 108.200 147.810 110.270 147.950 ;
        RECT 110.500 147.950 110.640 148.150 ;
        RECT 110.870 148.090 111.190 148.350 ;
        RECT 120.530 148.090 120.850 148.350 ;
        RECT 115.010 147.950 115.330 148.010 ;
        RECT 110.500 147.810 115.330 147.950 ;
        RECT 68.205 147.765 68.495 147.810 ;
        RECT 71.325 147.765 71.615 147.810 ;
        RECT 73.215 147.765 73.505 147.810 ;
        RECT 101.210 147.750 101.530 147.810 ;
        RECT 109.950 147.750 110.270 147.810 ;
        RECT 115.010 147.750 115.330 147.810 ;
        RECT 57.510 147.610 57.830 147.670 ;
        RECT 56.220 147.470 57.830 147.610 ;
        RECT 52.005 147.270 52.295 147.315 ;
        RECT 50.150 147.130 52.295 147.270 ;
        RECT 50.150 147.070 50.470 147.130 ;
        RECT 52.005 147.085 52.295 147.130 ;
        RECT 55.225 147.085 55.515 147.315 ;
        RECT 55.670 147.070 55.990 147.330 ;
        RECT 56.220 147.315 56.360 147.470 ;
        RECT 57.510 147.410 57.830 147.470 ;
        RECT 58.060 147.470 60.960 147.610 ;
        RECT 56.145 147.085 56.435 147.315 ;
        RECT 56.590 147.270 56.910 147.330 ;
        RECT 57.065 147.270 57.355 147.315 ;
        RECT 58.060 147.270 58.200 147.470 ;
        RECT 56.590 147.130 58.200 147.270 ;
        RECT 58.430 147.270 58.750 147.330 ;
        RECT 60.820 147.315 60.960 147.470 ;
        RECT 72.690 147.410 73.010 147.670 ;
        RECT 82.350 147.410 82.670 147.670 ;
        RECT 103.970 147.610 104.290 147.670 ;
        RECT 107.205 147.610 107.495 147.655 ;
        RECT 103.970 147.470 107.495 147.610 ;
        RECT 103.970 147.410 104.290 147.470 ;
        RECT 107.205 147.425 107.495 147.470 ;
        RECT 109.030 147.410 109.350 147.670 ;
        RECT 110.425 147.610 110.715 147.655 ;
        RECT 112.250 147.610 112.570 147.670 ;
        RECT 110.425 147.470 112.570 147.610 ;
        RECT 110.425 147.425 110.715 147.470 ;
        RECT 112.250 147.410 112.570 147.470 ;
        RECT 58.905 147.270 59.195 147.315 ;
        RECT 58.430 147.130 59.195 147.270 ;
        RECT 56.590 147.070 56.910 147.130 ;
        RECT 57.065 147.085 57.355 147.130 ;
        RECT 58.430 147.070 58.750 147.130 ;
        RECT 58.905 147.085 59.195 147.130 ;
        RECT 59.365 147.085 59.655 147.315 ;
        RECT 59.825 147.085 60.115 147.315 ;
        RECT 60.745 147.085 61.035 147.315 ;
        RECT 61.190 147.270 61.510 147.330 ;
        RECT 62.125 147.270 62.415 147.315 ;
        RECT 67.170 147.290 67.490 147.330 ;
        RECT 61.190 147.130 62.415 147.270 ;
        RECT 32.200 146.930 32.490 146.975 ;
        RECT 28.940 146.790 32.490 146.930 ;
        RECT 28.940 146.745 29.230 146.790 ;
        RECT 30.370 146.730 30.690 146.790 ;
        RECT 32.200 146.745 32.490 146.790 ;
        RECT 33.120 146.930 33.410 146.975 ;
        RECT 34.980 146.930 35.270 146.975 ;
        RECT 33.120 146.790 35.270 146.930 ;
        RECT 33.120 146.745 33.410 146.790 ;
        RECT 34.980 146.745 35.270 146.790 ;
        RECT 53.385 146.930 53.675 146.975 ;
        RECT 57.525 146.930 57.815 146.975 ;
        RECT 53.385 146.790 57.815 146.930 ;
        RECT 53.385 146.745 53.675 146.790 ;
        RECT 57.525 146.745 57.815 146.790 ;
        RECT 39.585 146.590 39.875 146.635 ;
        RECT 40.490 146.590 40.810 146.650 ;
        RECT 39.585 146.450 40.810 146.590 ;
        RECT 39.585 146.405 39.875 146.450 ;
        RECT 40.490 146.390 40.810 146.450 ;
        RECT 50.150 146.590 50.470 146.650 ;
        RECT 53.845 146.590 54.135 146.635 ;
        RECT 50.150 146.450 54.135 146.590 ;
        RECT 50.150 146.390 50.470 146.450 ;
        RECT 53.845 146.405 54.135 146.450 ;
        RECT 55.670 146.590 55.990 146.650 ;
        RECT 59.440 146.590 59.580 147.085 ;
        RECT 59.900 146.930 60.040 147.085 ;
        RECT 61.190 147.070 61.510 147.130 ;
        RECT 62.125 147.085 62.415 147.130 ;
        RECT 67.125 147.070 67.490 147.290 ;
        RECT 68.205 147.270 68.495 147.315 ;
        RECT 71.785 147.270 72.075 147.315 ;
        RECT 73.620 147.270 73.910 147.315 ;
        RECT 68.205 147.130 73.910 147.270 ;
        RECT 68.205 147.085 68.495 147.130 ;
        RECT 71.785 147.085 72.075 147.130 ;
        RECT 73.620 147.085 73.910 147.130 ;
        RECT 74.085 147.270 74.375 147.315 ;
        RECT 75.450 147.270 75.770 147.330 ;
        RECT 74.085 147.130 75.770 147.270 ;
        RECT 74.085 147.085 74.375 147.130 ;
        RECT 75.450 147.070 75.770 147.130 ;
        RECT 81.890 147.270 82.210 147.330 ;
        RECT 82.825 147.270 83.115 147.315 ;
        RECT 81.890 147.130 83.115 147.270 ;
        RECT 81.890 147.070 82.210 147.130 ;
        RECT 82.825 147.085 83.115 147.130 ;
        RECT 105.810 147.270 106.130 147.330 ;
        RECT 106.745 147.270 107.035 147.315 ;
        RECT 105.810 147.130 107.035 147.270 ;
        RECT 105.810 147.070 106.130 147.130 ;
        RECT 106.745 147.085 107.035 147.130 ;
        RECT 108.125 147.270 108.415 147.315 ;
        RECT 109.120 147.270 109.260 147.410 ;
        RECT 108.125 147.130 109.260 147.270 ;
        RECT 108.125 147.085 108.415 147.130 ;
        RECT 109.490 147.070 109.810 147.330 ;
        RECT 112.725 147.270 113.015 147.315 ;
        RECT 110.040 147.130 113.015 147.270 ;
        RECT 67.125 146.975 67.415 147.070 ;
        RECT 66.825 146.930 67.415 146.975 ;
        RECT 70.065 146.930 70.715 146.975 ;
        RECT 59.900 146.790 65.560 146.930 ;
        RECT 65.420 146.650 65.560 146.790 ;
        RECT 66.825 146.790 70.715 146.930 ;
        RECT 66.825 146.745 67.115 146.790 ;
        RECT 70.065 146.745 70.715 146.790 ;
        RECT 81.445 146.930 81.735 146.975 ;
        RECT 82.350 146.930 82.670 146.990 ;
        RECT 81.445 146.790 82.670 146.930 ;
        RECT 81.445 146.745 81.735 146.790 ;
        RECT 82.350 146.730 82.670 146.790 ;
        RECT 109.030 146.930 109.350 146.990 ;
        RECT 110.040 146.930 110.180 147.130 ;
        RECT 112.725 147.085 113.015 147.130 ;
        RECT 113.170 147.070 113.490 147.330 ;
        RECT 113.645 147.270 113.935 147.315 ;
        RECT 114.090 147.270 114.410 147.330 ;
        RECT 113.645 147.130 114.410 147.270 ;
        RECT 113.645 147.085 113.935 147.130 ;
        RECT 114.090 147.070 114.410 147.130 ;
        RECT 114.565 147.270 114.855 147.315 ;
        RECT 115.470 147.270 115.790 147.330 ;
        RECT 114.565 147.130 115.790 147.270 ;
        RECT 114.565 147.085 114.855 147.130 ;
        RECT 115.470 147.070 115.790 147.130 ;
        RECT 115.930 147.270 116.250 147.330 ;
        RECT 120.070 147.270 120.390 147.330 ;
        RECT 115.930 147.130 120.390 147.270 ;
        RECT 115.930 147.070 116.250 147.130 ;
        RECT 120.070 147.070 120.390 147.130 ;
        RECT 109.030 146.790 110.180 146.930 ;
        RECT 110.885 146.930 111.175 146.975 ;
        RECT 111.345 146.930 111.635 146.975 ;
        RECT 119.610 146.930 119.930 146.990 ;
        RECT 110.885 146.790 111.635 146.930 ;
        RECT 109.030 146.730 109.350 146.790 ;
        RECT 110.885 146.745 111.175 146.790 ;
        RECT 111.345 146.745 111.635 146.790 ;
        RECT 119.470 146.730 119.930 146.930 ;
        RECT 55.670 146.450 59.580 146.590 ;
        RECT 60.730 146.590 61.050 146.650 ;
        RECT 61.665 146.590 61.955 146.635 ;
        RECT 60.730 146.450 61.955 146.590 ;
        RECT 55.670 146.390 55.990 146.450 ;
        RECT 60.730 146.390 61.050 146.450 ;
        RECT 61.665 146.405 61.955 146.450 ;
        RECT 65.330 146.390 65.650 146.650 ;
        RECT 83.745 146.590 84.035 146.635 ;
        RECT 85.570 146.590 85.890 146.650 ;
        RECT 83.745 146.450 85.890 146.590 ;
        RECT 83.745 146.405 84.035 146.450 ;
        RECT 85.570 146.390 85.890 146.450 ;
        RECT 105.825 146.590 106.115 146.635 ;
        RECT 119.470 146.590 119.610 146.730 ;
        RECT 105.825 146.450 119.610 146.590 ;
        RECT 105.825 146.405 106.115 146.450 ;
        RECT 20.640 145.770 127.820 146.250 ;
        RECT 30.370 145.370 30.690 145.630 ;
        RECT 50.625 145.570 50.915 145.615 ;
        RECT 54.750 145.570 55.070 145.630 ;
        RECT 48.400 145.430 50.915 145.570 ;
        RECT 41.870 145.030 42.190 145.290 ;
        RECT 44.645 145.230 44.935 145.275 ;
        RECT 48.400 145.230 48.540 145.430 ;
        RECT 50.625 145.385 50.915 145.430 ;
        RECT 52.080 145.430 55.070 145.570 ;
        RECT 44.645 145.090 48.540 145.230 ;
        RECT 44.645 145.045 44.935 145.090 ;
        RECT 50.150 145.030 50.470 145.290 ;
        RECT 26.230 144.890 26.550 144.950 ;
        RECT 29.925 144.890 30.215 144.935 ;
        RECT 26.230 144.750 30.215 144.890 ;
        RECT 26.230 144.690 26.550 144.750 ;
        RECT 29.925 144.705 30.215 144.750 ;
        RECT 40.505 144.890 40.795 144.935 ;
        RECT 42.790 144.890 43.110 144.950 ;
        RECT 40.505 144.750 43.110 144.890 ;
        RECT 40.505 144.705 40.795 144.750 ;
        RECT 42.790 144.690 43.110 144.750 ;
        RECT 43.250 144.690 43.570 144.950 ;
        RECT 45.090 144.890 45.410 144.950 ;
        RECT 46.025 144.890 46.315 144.935 ;
        RECT 45.090 144.750 46.315 144.890 ;
        RECT 45.090 144.690 45.410 144.750 ;
        RECT 46.025 144.705 46.315 144.750 ;
        RECT 47.405 144.705 47.695 144.935 ;
        RECT 48.785 144.890 49.075 144.935 ;
        RECT 49.230 144.890 49.550 144.950 ;
        RECT 52.080 144.935 52.220 145.430 ;
        RECT 54.750 145.370 55.070 145.430 ;
        RECT 57.510 145.570 57.830 145.630 ;
        RECT 60.745 145.570 61.035 145.615 ;
        RECT 57.510 145.430 61.035 145.570 ;
        RECT 57.510 145.370 57.830 145.430 ;
        RECT 60.745 145.385 61.035 145.430 ;
        RECT 65.330 145.570 65.650 145.630 ;
        RECT 69.485 145.570 69.775 145.615 ;
        RECT 65.330 145.430 69.775 145.570 ;
        RECT 65.330 145.370 65.650 145.430 ;
        RECT 69.485 145.385 69.775 145.430 ;
        RECT 70.390 145.570 70.710 145.630 ;
        RECT 71.785 145.570 72.075 145.615 ;
        RECT 70.390 145.430 72.075 145.570 ;
        RECT 70.390 145.370 70.710 145.430 ;
        RECT 71.785 145.385 72.075 145.430 ;
        RECT 82.350 145.370 82.670 145.630 ;
        RECT 83.730 145.370 84.050 145.630 ;
        RECT 53.370 145.230 53.690 145.290 ;
        RECT 52.540 145.090 53.690 145.230 ;
        RECT 54.840 145.230 54.980 145.370 ;
        RECT 67.170 145.230 67.490 145.290 ;
        RECT 74.530 145.230 74.850 145.290 ;
        RECT 83.820 145.230 83.960 145.370 ;
        RECT 54.840 145.090 55.900 145.230 ;
        RECT 52.540 144.935 52.680 145.090 ;
        RECT 53.370 145.030 53.690 145.090 ;
        RECT 48.785 144.750 49.550 144.890 ;
        RECT 48.785 144.705 49.075 144.750 ;
        RECT 41.410 144.350 41.730 144.610 ;
        RECT 42.330 144.550 42.650 144.610 ;
        RECT 43.725 144.550 44.015 144.595 ;
        RECT 42.330 144.410 44.015 144.550 ;
        RECT 42.330 144.350 42.650 144.410 ;
        RECT 43.725 144.365 44.015 144.410 ;
        RECT 45.550 144.550 45.870 144.610 ;
        RECT 46.485 144.550 46.775 144.595 ;
        RECT 45.550 144.410 46.775 144.550 ;
        RECT 45.550 144.350 45.870 144.410 ;
        RECT 46.485 144.365 46.775 144.410 ;
        RECT 30.830 144.210 31.150 144.270 ;
        RECT 39.585 144.210 39.875 144.255 ;
        RECT 30.830 144.070 39.875 144.210 ;
        RECT 47.480 144.210 47.620 144.705 ;
        RECT 49.230 144.690 49.550 144.750 ;
        RECT 52.005 144.705 52.295 144.935 ;
        RECT 52.465 144.705 52.755 144.935 ;
        RECT 52.925 144.705 53.215 144.935 ;
        RECT 53.845 144.890 54.135 144.935 ;
        RECT 55.210 144.890 55.530 144.950 ;
        RECT 55.760 144.935 55.900 145.090 ;
        RECT 56.680 145.090 60.500 145.230 ;
        RECT 53.845 144.750 55.530 144.890 ;
        RECT 53.845 144.705 54.135 144.750 ;
        RECT 47.850 144.550 48.170 144.610 ;
        RECT 49.705 144.550 49.995 144.595 ;
        RECT 47.850 144.410 49.995 144.550 ;
        RECT 53.000 144.550 53.140 144.705 ;
        RECT 55.210 144.690 55.530 144.750 ;
        RECT 55.685 144.705 55.975 144.935 ;
        RECT 56.130 144.690 56.450 144.950 ;
        RECT 56.680 144.935 56.820 145.090 ;
        RECT 56.605 144.705 56.895 144.935 ;
        RECT 57.050 144.890 57.370 144.950 ;
        RECT 57.525 144.890 57.815 144.935 ;
        RECT 57.050 144.750 57.815 144.890 ;
        RECT 57.050 144.690 57.370 144.750 ;
        RECT 57.525 144.705 57.815 144.750 ;
        RECT 60.360 144.610 60.500 145.090 ;
        RECT 65.880 145.090 74.850 145.230 ;
        RECT 65.880 144.935 66.020 145.090 ;
        RECT 67.170 145.030 67.490 145.090 ;
        RECT 74.530 145.030 74.850 145.090 ;
        RECT 80.140 145.090 84.420 145.230 ;
        RECT 65.805 144.705 66.095 144.935 ;
        RECT 66.265 144.705 66.555 144.935 ;
        RECT 53.000 144.410 57.740 144.550 ;
        RECT 47.850 144.350 48.170 144.410 ;
        RECT 49.705 144.365 49.995 144.410 ;
        RECT 57.600 144.270 57.740 144.410 ;
        RECT 59.810 144.350 60.130 144.610 ;
        RECT 60.270 144.350 60.590 144.610 ;
        RECT 66.340 144.550 66.480 144.705 ;
        RECT 66.710 144.690 67.030 144.950 ;
        RECT 67.630 144.690 67.950 144.950 ;
        RECT 69.930 144.690 70.250 144.950 ;
        RECT 72.230 144.890 72.550 144.950 ;
        RECT 73.165 144.890 73.455 144.935 ;
        RECT 75.910 144.890 76.230 144.950 ;
        RECT 80.140 144.935 80.280 145.090 ;
        RECT 72.230 144.750 76.230 144.890 ;
        RECT 72.230 144.690 72.550 144.750 ;
        RECT 73.165 144.705 73.455 144.750 ;
        RECT 75.910 144.690 76.230 144.750 ;
        RECT 78.685 144.890 78.975 144.935 ;
        RECT 78.685 144.750 79.360 144.890 ;
        RECT 78.685 144.705 78.975 144.750 ;
        RECT 68.090 144.550 68.410 144.610 ;
        RECT 66.340 144.410 68.410 144.550 ;
        RECT 68.090 144.350 68.410 144.410 ;
        RECT 68.565 144.365 68.855 144.595 ;
        RECT 69.470 144.550 69.790 144.610 ;
        RECT 76.370 144.550 76.690 144.610 ;
        RECT 69.470 144.410 76.690 144.550 ;
        RECT 54.305 144.210 54.595 144.255 ;
        RECT 47.480 144.070 54.595 144.210 ;
        RECT 30.830 144.010 31.150 144.070 ;
        RECT 39.585 144.025 39.875 144.070 ;
        RECT 54.305 144.025 54.595 144.070 ;
        RECT 57.510 144.010 57.830 144.270 ;
        RECT 59.900 144.210 60.040 144.350 ;
        RECT 68.640 144.210 68.780 144.365 ;
        RECT 69.470 144.350 69.790 144.410 ;
        RECT 76.370 144.350 76.690 144.410 ;
        RECT 70.850 144.210 71.170 144.270 ;
        RECT 59.900 144.070 71.170 144.210 ;
        RECT 79.220 144.210 79.360 144.750 ;
        RECT 79.605 144.705 79.895 144.935 ;
        RECT 80.065 144.705 80.355 144.935 ;
        RECT 80.525 144.890 80.815 144.935 ;
        RECT 83.730 144.890 84.050 144.950 ;
        RECT 84.280 144.935 84.420 145.090 ;
        RECT 110.410 145.030 110.730 145.290 ;
        RECT 80.525 144.750 84.050 144.890 ;
        RECT 80.525 144.705 80.815 144.750 ;
        RECT 79.680 144.550 79.820 144.705 ;
        RECT 83.730 144.690 84.050 144.750 ;
        RECT 84.205 144.705 84.495 144.935 ;
        RECT 84.665 144.890 84.955 144.935 ;
        RECT 85.110 144.890 85.430 144.950 ;
        RECT 84.665 144.750 85.430 144.890 ;
        RECT 84.665 144.705 84.955 144.750 ;
        RECT 85.110 144.690 85.430 144.750 ;
        RECT 85.585 144.890 85.875 144.935 ;
        RECT 86.030 144.890 86.350 144.950 ;
        RECT 85.585 144.750 86.350 144.890 ;
        RECT 85.585 144.705 85.875 144.750 ;
        RECT 79.680 144.410 84.880 144.550 ;
        RECT 84.740 144.270 84.880 144.410 ;
        RECT 79.220 144.070 82.580 144.210 ;
        RECT 70.850 144.010 71.170 144.070 ;
        RECT 36.810 143.870 37.130 143.930 ;
        RECT 40.505 143.870 40.795 143.915 ;
        RECT 36.810 143.730 40.795 143.870 ;
        RECT 36.810 143.670 37.130 143.730 ;
        RECT 40.505 143.685 40.795 143.730 ;
        RECT 42.345 143.870 42.635 143.915 ;
        RECT 42.790 143.870 43.110 143.930 ;
        RECT 42.345 143.730 43.110 143.870 ;
        RECT 42.345 143.685 42.635 143.730 ;
        RECT 42.790 143.670 43.110 143.730 ;
        RECT 44.170 143.670 44.490 143.930 ;
        RECT 45.105 143.870 45.395 143.915 ;
        RECT 45.550 143.870 45.870 143.930 ;
        RECT 45.105 143.730 45.870 143.870 ;
        RECT 45.105 143.685 45.395 143.730 ;
        RECT 45.550 143.670 45.870 143.730 ;
        RECT 46.470 143.670 46.790 143.930 ;
        RECT 47.865 143.870 48.155 143.915 ;
        RECT 48.310 143.870 48.630 143.930 ;
        RECT 47.865 143.730 48.630 143.870 ;
        RECT 47.865 143.685 48.155 143.730 ;
        RECT 48.310 143.670 48.630 143.730 ;
        RECT 48.770 143.670 49.090 143.930 ;
        RECT 61.190 143.870 61.510 143.930 ;
        RECT 62.585 143.870 62.875 143.915 ;
        RECT 61.190 143.730 62.875 143.870 ;
        RECT 61.190 143.670 61.510 143.730 ;
        RECT 62.585 143.685 62.875 143.730 ;
        RECT 64.410 143.670 64.730 143.930 ;
        RECT 71.770 143.870 72.090 143.930 ;
        RECT 72.705 143.870 72.995 143.915 ;
        RECT 71.770 143.730 72.995 143.870 ;
        RECT 71.770 143.670 72.090 143.730 ;
        RECT 72.705 143.685 72.995 143.730 ;
        RECT 81.890 143.670 82.210 143.930 ;
        RECT 82.440 143.870 82.580 144.070 ;
        RECT 84.650 144.010 84.970 144.270 ;
        RECT 85.660 143.870 85.800 144.705 ;
        RECT 86.030 144.690 86.350 144.750 ;
        RECT 111.330 144.690 111.650 144.950 ;
        RECT 111.790 144.690 112.110 144.950 ;
        RECT 117.785 144.890 118.075 144.935 ;
        RECT 119.625 144.890 119.915 144.935 ;
        RECT 120.070 144.890 120.390 144.950 ;
        RECT 117.785 144.750 120.390 144.890 ;
        RECT 117.785 144.705 118.075 144.750 ;
        RECT 119.625 144.705 119.915 144.750 ;
        RECT 120.070 144.690 120.390 144.750 ;
        RECT 108.110 144.550 108.430 144.610 ;
        RECT 115.470 144.550 115.790 144.610 ;
        RECT 108.110 144.410 115.790 144.550 ;
        RECT 108.110 144.350 108.430 144.410 ;
        RECT 115.470 144.350 115.790 144.410 ;
        RECT 109.030 144.210 109.350 144.270 ;
        RECT 110.410 144.210 110.730 144.270 ;
        RECT 109.030 144.070 110.730 144.210 ;
        RECT 109.030 144.010 109.350 144.070 ;
        RECT 110.410 144.010 110.730 144.070 ;
        RECT 82.440 143.730 85.800 143.870 ;
        RECT 94.310 143.870 94.630 143.930 ;
        RECT 102.130 143.870 102.450 143.930 ;
        RECT 94.310 143.730 102.450 143.870 ;
        RECT 94.310 143.670 94.630 143.730 ;
        RECT 102.130 143.670 102.450 143.730 ;
        RECT 111.790 143.670 112.110 143.930 ;
        RECT 112.725 143.870 113.015 143.915 ;
        RECT 115.930 143.870 116.250 143.930 ;
        RECT 112.725 143.730 116.250 143.870 ;
        RECT 112.725 143.685 113.015 143.730 ;
        RECT 115.930 143.670 116.250 143.730 ;
        RECT 118.230 143.670 118.550 143.930 ;
        RECT 120.070 143.670 120.390 143.930 ;
        RECT 20.640 143.050 127.820 143.530 ;
        RECT 43.710 142.650 44.030 142.910 ;
        RECT 46.485 142.850 46.775 142.895 ;
        RECT 48.770 142.850 49.090 142.910 ;
        RECT 46.485 142.710 49.090 142.850 ;
        RECT 46.485 142.665 46.775 142.710 ;
        RECT 48.770 142.650 49.090 142.710 ;
        RECT 68.090 142.850 68.410 142.910 ;
        RECT 73.610 142.850 73.930 142.910 ;
        RECT 81.905 142.850 82.195 142.895 ;
        RECT 82.350 142.850 82.670 142.910 ;
        RECT 68.090 142.710 81.660 142.850 ;
        RECT 68.090 142.650 68.410 142.710 ;
        RECT 73.610 142.650 73.930 142.710 ;
        RECT 60.240 142.510 60.530 142.555 ;
        RECT 63.020 142.510 63.310 142.555 ;
        RECT 64.880 142.510 65.170 142.555 ;
        RECT 60.240 142.370 65.170 142.510 ;
        RECT 60.240 142.325 60.530 142.370 ;
        RECT 63.020 142.325 63.310 142.370 ;
        RECT 64.880 142.325 65.170 142.370 ;
        RECT 70.360 142.510 70.650 142.555 ;
        RECT 73.140 142.510 73.430 142.555 ;
        RECT 75.000 142.510 75.290 142.555 ;
        RECT 70.360 142.370 75.290 142.510 ;
        RECT 81.520 142.510 81.660 142.710 ;
        RECT 81.905 142.710 82.670 142.850 ;
        RECT 81.905 142.665 82.195 142.710 ;
        RECT 82.350 142.650 82.670 142.710 ;
        RECT 85.110 142.850 85.430 142.910 ;
        RECT 86.030 142.850 86.350 142.910 ;
        RECT 86.735 142.850 87.025 142.895 ;
        RECT 111.330 142.850 111.650 142.910 ;
        RECT 112.710 142.850 113.030 142.910 ;
        RECT 85.110 142.710 87.025 142.850 ;
        RECT 85.110 142.650 85.430 142.710 ;
        RECT 86.030 142.650 86.350 142.710 ;
        RECT 86.735 142.665 87.025 142.710 ;
        RECT 87.500 142.710 99.600 142.850 ;
        RECT 81.520 142.370 83.040 142.510 ;
        RECT 70.360 142.325 70.650 142.370 ;
        RECT 73.140 142.325 73.430 142.370 ;
        RECT 75.000 142.325 75.290 142.370 ;
        RECT 40.030 142.170 40.350 142.230 ;
        RECT 43.265 142.170 43.555 142.215 ;
        RECT 64.410 142.170 64.730 142.230 ;
        RECT 40.030 142.030 43.555 142.170 ;
        RECT 40.030 141.970 40.350 142.030 ;
        RECT 43.265 141.985 43.555 142.030 ;
        RECT 44.720 142.030 64.730 142.170 ;
        RECT 42.805 141.830 43.095 141.875 ;
        RECT 44.720 141.830 44.860 142.030 ;
        RECT 64.410 141.970 64.730 142.030 ;
        RECT 66.495 142.170 66.785 142.215 ;
        RECT 69.930 142.170 70.250 142.230 ;
        RECT 66.495 142.030 70.250 142.170 ;
        RECT 66.495 141.985 66.785 142.030 ;
        RECT 69.930 141.970 70.250 142.030 ;
        RECT 74.530 141.970 74.850 142.230 ;
        RECT 75.450 141.970 75.770 142.230 ;
        RECT 81.430 141.970 81.750 142.230 ;
        RECT 42.805 141.690 44.860 141.830 ;
        RECT 42.805 141.645 43.095 141.690 ;
        RECT 45.090 141.630 45.410 141.890 ;
        RECT 45.565 141.830 45.855 141.875 ;
        RECT 46.010 141.830 46.330 141.890 ;
        RECT 45.565 141.690 46.330 141.830 ;
        RECT 45.565 141.645 45.855 141.690 ;
        RECT 46.010 141.630 46.330 141.690 ;
        RECT 60.240 141.830 60.530 141.875 ;
        RECT 60.240 141.690 62.775 141.830 ;
        RECT 60.240 141.645 60.530 141.690 ;
        RECT 44.185 141.490 44.475 141.535 ;
        RECT 44.630 141.490 44.950 141.550 ;
        RECT 44.185 141.350 44.950 141.490 ;
        RECT 44.185 141.305 44.475 141.350 ;
        RECT 44.630 141.290 44.950 141.350 ;
        RECT 58.380 141.490 58.670 141.535 ;
        RECT 60.730 141.490 61.050 141.550 ;
        RECT 62.560 141.535 62.775 141.690 ;
        RECT 63.490 141.630 63.810 141.890 ;
        RECT 63.950 141.830 64.270 141.890 ;
        RECT 65.345 141.830 65.635 141.875 ;
        RECT 63.950 141.690 65.635 141.830 ;
        RECT 63.950 141.630 64.270 141.690 ;
        RECT 65.345 141.645 65.635 141.690 ;
        RECT 70.360 141.830 70.650 141.875 ;
        RECT 70.360 141.690 72.895 141.830 ;
        RECT 70.360 141.645 70.650 141.690 ;
        RECT 71.770 141.535 72.090 141.550 ;
        RECT 61.640 141.490 61.930 141.535 ;
        RECT 58.380 141.350 61.930 141.490 ;
        RECT 58.380 141.305 58.670 141.350 ;
        RECT 60.730 141.290 61.050 141.350 ;
        RECT 61.640 141.305 61.930 141.350 ;
        RECT 62.560 141.490 62.850 141.535 ;
        RECT 64.420 141.490 64.710 141.535 ;
        RECT 62.560 141.350 64.710 141.490 ;
        RECT 62.560 141.305 62.850 141.350 ;
        RECT 64.420 141.305 64.710 141.350 ;
        RECT 68.500 141.490 68.790 141.535 ;
        RECT 71.760 141.490 72.090 141.535 ;
        RECT 68.500 141.350 72.090 141.490 ;
        RECT 68.500 141.305 68.790 141.350 ;
        RECT 71.760 141.305 72.090 141.350 ;
        RECT 72.680 141.535 72.895 141.690 ;
        RECT 73.610 141.630 73.930 141.890 ;
        RECT 74.620 141.830 74.760 141.970 ;
        RECT 80.525 141.830 80.815 141.875 ;
        RECT 80.970 141.830 81.290 141.890 ;
        RECT 74.620 141.690 80.280 141.830 ;
        RECT 72.680 141.490 72.970 141.535 ;
        RECT 74.540 141.490 74.830 141.535 ;
        RECT 72.680 141.350 74.830 141.490 ;
        RECT 80.140 141.490 80.280 141.690 ;
        RECT 80.525 141.690 81.290 141.830 ;
        RECT 80.525 141.645 80.815 141.690 ;
        RECT 80.970 141.630 81.290 141.690 ;
        RECT 81.890 141.630 82.210 141.890 ;
        RECT 82.900 141.830 83.040 142.370 ;
        RECT 83.360 142.370 87.180 142.510 ;
        RECT 83.360 142.215 83.500 142.370 ;
        RECT 87.040 142.230 87.180 142.370 ;
        RECT 83.285 141.985 83.575 142.215 ;
        RECT 83.745 142.170 84.035 142.215 ;
        RECT 86.030 142.170 86.350 142.230 ;
        RECT 83.745 142.030 86.350 142.170 ;
        RECT 83.745 141.985 84.035 142.030 ;
        RECT 86.030 141.970 86.350 142.030 ;
        RECT 86.950 141.970 87.270 142.230 ;
        RECT 87.500 141.830 87.640 142.710 ;
        RECT 90.600 142.510 90.890 142.555 ;
        RECT 93.380 142.510 93.670 142.555 ;
        RECT 95.240 142.510 95.530 142.555 ;
        RECT 90.600 142.370 95.530 142.510 ;
        RECT 90.600 142.325 90.890 142.370 ;
        RECT 93.380 142.325 93.670 142.370 ;
        RECT 95.240 142.325 95.530 142.370 ;
        RECT 99.460 142.510 99.600 142.710 ;
        RECT 110.095 142.710 113.030 142.850 ;
        RECT 110.095 142.510 110.235 142.710 ;
        RECT 111.330 142.650 111.650 142.710 ;
        RECT 112.710 142.650 113.030 142.710 ;
        RECT 99.460 142.370 110.235 142.510 ;
        RECT 87.870 142.170 88.190 142.230 ;
        RECT 87.870 142.030 93.620 142.170 ;
        RECT 87.870 141.970 88.190 142.030 ;
        RECT 82.900 141.690 87.640 141.830 ;
        RECT 90.600 141.830 90.890 141.875 ;
        RECT 93.480 141.830 93.620 142.030 ;
        RECT 93.850 141.970 94.170 142.230 ;
        RECT 96.150 142.170 96.470 142.230 ;
        RECT 96.150 142.030 99.140 142.170 ;
        RECT 96.150 141.970 96.470 142.030 ;
        RECT 95.705 141.830 95.995 141.875 ;
        RECT 90.600 141.690 93.135 141.830 ;
        RECT 93.480 141.690 95.995 141.830 ;
        RECT 90.600 141.645 90.890 141.690 ;
        RECT 86.490 141.490 86.810 141.550 ;
        RECT 88.790 141.535 89.110 141.550 ;
        RECT 92.920 141.535 93.135 141.690 ;
        RECT 95.705 141.645 95.995 141.690 ;
        RECT 97.530 141.630 97.850 141.890 ;
        RECT 98.005 141.830 98.295 141.875 ;
        RECT 98.450 141.830 98.770 141.890 ;
        RECT 99.000 141.875 99.140 142.030 ;
        RECT 99.460 141.875 99.600 142.370 ;
        RECT 104.905 142.170 105.195 142.215 ;
        RECT 105.810 142.170 106.130 142.230 ;
        RECT 104.905 142.030 106.130 142.170 ;
        RECT 110.095 142.170 110.235 142.370 ;
        RECT 110.410 142.510 110.730 142.570 ;
        RECT 120.960 142.510 121.250 142.555 ;
        RECT 123.740 142.510 124.030 142.555 ;
        RECT 125.600 142.510 125.890 142.555 ;
        RECT 110.410 142.370 111.100 142.510 ;
        RECT 110.410 142.310 110.730 142.370 ;
        RECT 110.095 142.030 110.640 142.170 ;
        RECT 104.905 141.985 105.195 142.030 ;
        RECT 105.810 141.970 106.130 142.030 ;
        RECT 98.005 141.690 98.770 141.830 ;
        RECT 98.005 141.645 98.295 141.690 ;
        RECT 98.450 141.630 98.770 141.690 ;
        RECT 98.925 141.645 99.215 141.875 ;
        RECT 99.385 141.645 99.675 141.875 ;
        RECT 99.845 141.830 100.135 141.875 ;
        RECT 100.290 141.830 100.610 141.890 ;
        RECT 99.845 141.690 100.610 141.830 ;
        RECT 99.845 141.645 100.135 141.690 ;
        RECT 100.290 141.630 100.610 141.690 ;
        RECT 102.130 141.630 102.450 141.890 ;
        RECT 104.430 141.830 104.750 141.890 ;
        RECT 108.110 141.830 108.430 141.890 ;
        RECT 110.500 141.875 110.640 142.030 ;
        RECT 110.960 141.875 111.100 142.370 ;
        RECT 120.960 142.370 125.890 142.510 ;
        RECT 120.960 142.325 121.250 142.370 ;
        RECT 123.740 142.325 124.030 142.370 ;
        RECT 125.600 142.325 125.890 142.370 ;
        RECT 113.170 141.970 113.490 142.230 ;
        RECT 114.090 142.170 114.410 142.230 ;
        RECT 123.290 142.170 123.610 142.230 ;
        RECT 124.225 142.170 124.515 142.215 ;
        RECT 114.090 142.030 114.780 142.170 ;
        RECT 114.090 141.970 114.410 142.030 ;
        RECT 114.640 141.875 114.780 142.030 ;
        RECT 123.290 142.030 124.515 142.170 ;
        RECT 123.290 141.970 123.610 142.030 ;
        RECT 124.225 141.985 124.515 142.030 ;
        RECT 109.045 141.830 109.335 141.875 ;
        RECT 104.430 141.690 109.335 141.830 ;
        RECT 104.430 141.630 104.750 141.690 ;
        RECT 108.110 141.630 108.430 141.690 ;
        RECT 109.045 141.645 109.335 141.690 ;
        RECT 109.965 141.645 110.255 141.875 ;
        RECT 110.425 141.645 110.715 141.875 ;
        RECT 110.885 141.645 111.175 141.875 ;
        RECT 114.565 141.645 114.855 141.875 ;
        RECT 120.960 141.830 121.250 141.875 ;
        RECT 124.670 141.830 124.990 141.890 ;
        RECT 126.065 141.830 126.355 141.875 ;
        RECT 120.960 141.690 123.495 141.830 ;
        RECT 120.960 141.645 121.250 141.690 ;
        RECT 80.140 141.350 86.810 141.490 ;
        RECT 72.680 141.305 72.970 141.350 ;
        RECT 74.540 141.305 74.830 141.350 ;
        RECT 71.770 141.290 72.090 141.305 ;
        RECT 86.490 141.290 86.810 141.350 ;
        RECT 88.740 141.490 89.110 141.535 ;
        RECT 92.000 141.490 92.290 141.535 ;
        RECT 88.740 141.350 92.290 141.490 ;
        RECT 88.740 141.305 89.110 141.350 ;
        RECT 92.000 141.305 92.290 141.350 ;
        RECT 92.920 141.490 93.210 141.535 ;
        RECT 94.780 141.490 95.070 141.535 ;
        RECT 92.920 141.350 95.070 141.490 ;
        RECT 92.920 141.305 93.210 141.350 ;
        RECT 94.780 141.305 95.070 141.350 ;
        RECT 104.890 141.490 105.210 141.550 ;
        RECT 105.365 141.490 105.655 141.535 ;
        RECT 104.890 141.350 105.655 141.490 ;
        RECT 88.790 141.290 89.110 141.305 ;
        RECT 104.890 141.290 105.210 141.350 ;
        RECT 105.365 141.305 105.655 141.350 ;
        RECT 105.825 141.490 106.115 141.535 ;
        RECT 108.570 141.490 108.890 141.550 ;
        RECT 105.825 141.350 108.890 141.490 ;
        RECT 110.040 141.490 110.180 141.645 ;
        RECT 112.710 141.490 113.030 141.550 ;
        RECT 114.105 141.490 114.395 141.535 ;
        RECT 117.095 141.490 117.385 141.535 ;
        RECT 110.040 141.350 117.385 141.490 ;
        RECT 105.825 141.305 106.115 141.350 ;
        RECT 108.570 141.290 108.890 141.350 ;
        RECT 112.710 141.290 113.030 141.350 ;
        RECT 114.105 141.305 114.395 141.350 ;
        RECT 117.095 141.305 117.385 141.350 ;
        RECT 119.100 141.490 119.390 141.535 ;
        RECT 120.070 141.490 120.390 141.550 ;
        RECT 123.280 141.535 123.495 141.690 ;
        RECT 124.670 141.690 126.355 141.830 ;
        RECT 124.670 141.630 124.990 141.690 ;
        RECT 126.065 141.645 126.355 141.690 ;
        RECT 122.360 141.490 122.650 141.535 ;
        RECT 119.100 141.350 122.650 141.490 ;
        RECT 119.100 141.305 119.390 141.350 ;
        RECT 120.070 141.290 120.390 141.350 ;
        RECT 122.360 141.305 122.650 141.350 ;
        RECT 123.280 141.490 123.570 141.535 ;
        RECT 125.140 141.490 125.430 141.535 ;
        RECT 123.280 141.350 125.430 141.490 ;
        RECT 123.280 141.305 123.570 141.350 ;
        RECT 125.140 141.305 125.430 141.350 ;
        RECT 135.635 141.220 136.775 165.470 ;
        RECT 38.190 141.150 38.510 141.210 ;
        RECT 41.885 141.150 42.175 141.195 ;
        RECT 38.190 141.010 42.175 141.150 ;
        RECT 38.190 140.950 38.510 141.010 ;
        RECT 41.885 140.965 42.175 141.010 ;
        RECT 56.375 141.150 56.665 141.195 ;
        RECT 60.270 141.150 60.590 141.210 ;
        RECT 56.375 141.010 60.590 141.150 ;
        RECT 56.375 140.965 56.665 141.010 ;
        RECT 60.270 140.950 60.590 141.010 ;
        RECT 79.605 141.150 79.895 141.195 ;
        RECT 81.430 141.150 81.750 141.210 ;
        RECT 79.605 141.010 81.750 141.150 ;
        RECT 79.605 140.965 79.895 141.010 ;
        RECT 81.430 140.950 81.750 141.010 ;
        RECT 84.205 141.150 84.495 141.195 ;
        RECT 85.110 141.150 85.430 141.210 ;
        RECT 84.205 141.010 85.430 141.150 ;
        RECT 84.205 140.965 84.495 141.010 ;
        RECT 85.110 140.950 85.430 141.010 ;
        RECT 86.030 140.950 86.350 141.210 ;
        RECT 96.625 141.150 96.915 141.195 ;
        RECT 97.070 141.150 97.390 141.210 ;
        RECT 96.625 141.010 97.390 141.150 ;
        RECT 96.625 140.965 96.915 141.010 ;
        RECT 97.070 140.950 97.390 141.010 ;
        RECT 100.750 141.150 101.070 141.210 ;
        RECT 101.225 141.150 101.515 141.195 ;
        RECT 100.750 141.010 101.515 141.150 ;
        RECT 100.750 140.950 101.070 141.010 ;
        RECT 101.225 140.965 101.515 141.010 ;
        RECT 102.590 140.950 102.910 141.210 ;
        RECT 107.665 141.150 107.955 141.195 ;
        RECT 109.950 141.150 110.270 141.210 ;
        RECT 107.665 141.010 110.270 141.150 ;
        RECT 107.665 140.965 107.955 141.010 ;
        RECT 109.950 140.950 110.270 141.010 ;
        RECT 112.265 141.150 112.555 141.195 ;
        RECT 113.630 141.150 113.950 141.210 ;
        RECT 112.265 141.010 113.950 141.150 ;
        RECT 112.265 140.965 112.555 141.010 ;
        RECT 113.630 140.950 113.950 141.010 ;
        RECT 116.390 140.950 116.710 141.210 ;
        RECT 20.640 140.330 127.820 140.810 ;
        RECT 135.580 140.230 136.830 141.220 ;
        RECT 32.685 139.945 32.975 140.175 ;
        RECT 25.260 139.790 25.550 139.835 ;
        RECT 27.610 139.790 27.930 139.850 ;
        RECT 28.520 139.790 28.810 139.835 ;
        RECT 25.260 139.650 28.810 139.790 ;
        RECT 25.260 139.605 25.550 139.650 ;
        RECT 27.610 139.590 27.930 139.650 ;
        RECT 28.520 139.605 28.810 139.650 ;
        RECT 29.440 139.790 29.730 139.835 ;
        RECT 31.300 139.790 31.590 139.835 ;
        RECT 29.440 139.650 31.590 139.790 ;
        RECT 29.440 139.605 29.730 139.650 ;
        RECT 31.300 139.605 31.590 139.650 ;
        RECT 27.120 139.450 27.410 139.495 ;
        RECT 29.440 139.450 29.655 139.605 ;
        RECT 27.120 139.310 29.655 139.450 ;
        RECT 30.385 139.450 30.675 139.495 ;
        RECT 32.760 139.450 32.900 139.945 ;
        RECT 41.870 139.930 42.190 140.190 ;
        RECT 44.170 139.930 44.490 140.190 ;
        RECT 46.470 139.930 46.790 140.190 ;
        RECT 62.585 140.130 62.875 140.175 ;
        RECT 63.490 140.130 63.810 140.190 ;
        RECT 62.585 139.990 63.810 140.130 ;
        RECT 62.585 139.945 62.875 139.990 ;
        RECT 63.490 139.930 63.810 139.990 ;
        RECT 64.410 140.130 64.730 140.190 ;
        RECT 72.705 140.130 72.995 140.175 ;
        RECT 73.610 140.130 73.930 140.190 ;
        RECT 64.410 139.990 72.000 140.130 ;
        RECT 64.410 139.930 64.730 139.990 ;
        RECT 41.960 139.790 42.100 139.930 ;
        RECT 66.265 139.790 66.555 139.835 ;
        RECT 41.960 139.650 66.555 139.790 ;
        RECT 66.265 139.605 66.555 139.650 ;
        RECT 68.640 139.650 70.160 139.790 ;
        RECT 30.385 139.310 32.900 139.450 ;
        RECT 33.605 139.450 33.895 139.495 ;
        RECT 34.050 139.450 34.370 139.510 ;
        RECT 33.605 139.310 34.370 139.450 ;
        RECT 27.120 139.265 27.410 139.310 ;
        RECT 30.385 139.265 30.675 139.310 ;
        RECT 33.605 139.265 33.895 139.310 ;
        RECT 34.050 139.250 34.370 139.310 ;
        RECT 34.970 139.450 35.290 139.510 ;
        RECT 35.445 139.450 35.735 139.495 ;
        RECT 38.650 139.450 38.970 139.510 ;
        RECT 34.970 139.310 38.970 139.450 ;
        RECT 34.970 139.250 35.290 139.310 ;
        RECT 35.445 139.265 35.735 139.310 ;
        RECT 38.650 139.250 38.970 139.310 ;
        RECT 41.870 139.250 42.190 139.510 ;
        RECT 43.265 139.450 43.555 139.495 ;
        RECT 45.565 139.450 45.855 139.495 ;
        RECT 46.010 139.450 46.330 139.510 ;
        RECT 50.625 139.450 50.915 139.495 ;
        RECT 52.925 139.450 53.215 139.495 ;
        RECT 53.370 139.450 53.690 139.510 ;
        RECT 43.265 139.310 53.690 139.450 ;
        RECT 43.265 139.265 43.555 139.310 ;
        RECT 45.565 139.265 45.855 139.310 ;
        RECT 46.010 139.250 46.330 139.310 ;
        RECT 50.625 139.265 50.915 139.310 ;
        RECT 52.925 139.265 53.215 139.310 ;
        RECT 53.370 139.250 53.690 139.310 ;
        RECT 61.190 139.450 61.510 139.510 ;
        RECT 61.665 139.450 61.955 139.495 ;
        RECT 61.190 139.310 61.955 139.450 ;
        RECT 61.190 139.250 61.510 139.310 ;
        RECT 61.665 139.265 61.955 139.310 ;
        RECT 67.170 139.450 67.490 139.510 ;
        RECT 67.645 139.450 67.935 139.495 ;
        RECT 67.170 139.310 67.935 139.450 ;
        RECT 67.170 139.250 67.490 139.310 ;
        RECT 67.645 139.265 67.935 139.310 ;
        RECT 68.090 139.250 68.410 139.510 ;
        RECT 68.640 139.495 68.780 139.650 ;
        RECT 70.020 139.510 70.160 139.650 ;
        RECT 70.850 139.590 71.170 139.850 ;
        RECT 68.565 139.265 68.855 139.495 ;
        RECT 69.470 139.250 69.790 139.510 ;
        RECT 69.930 139.250 70.250 139.510 ;
        RECT 71.860 139.495 72.000 139.990 ;
        RECT 72.705 139.990 73.930 140.130 ;
        RECT 72.705 139.945 72.995 139.990 ;
        RECT 73.610 139.930 73.930 139.990 ;
        RECT 87.885 140.130 88.175 140.175 ;
        RECT 88.790 140.130 89.110 140.190 ;
        RECT 98.450 140.130 98.770 140.190 ;
        RECT 104.430 140.130 104.750 140.190 ;
        RECT 108.110 140.130 108.430 140.190 ;
        RECT 87.885 139.990 89.110 140.130 ;
        RECT 87.885 139.945 88.175 139.990 ;
        RECT 88.790 139.930 89.110 139.990 ;
        RECT 89.800 139.990 108.430 140.130 ;
        RECT 76.370 139.790 76.690 139.850 ;
        RECT 89.800 139.790 89.940 139.990 ;
        RECT 98.450 139.930 98.770 139.990 ;
        RECT 104.430 139.930 104.750 139.990 ;
        RECT 108.110 139.930 108.430 139.990 ;
        RECT 109.030 140.130 109.350 140.190 ;
        RECT 111.805 140.130 112.095 140.175 ;
        RECT 109.030 139.990 112.095 140.130 ;
        RECT 109.030 139.930 109.350 139.990 ;
        RECT 111.805 139.945 112.095 139.990 ;
        RECT 112.265 140.130 112.555 140.175 ;
        RECT 112.710 140.130 113.030 140.190 ;
        RECT 135.635 140.155 136.775 140.230 ;
        RECT 112.265 139.990 113.030 140.130 ;
        RECT 112.265 139.945 112.555 139.990 ;
        RECT 76.370 139.650 89.940 139.790 ;
        RECT 91.090 139.790 91.410 139.850 ;
        RECT 91.960 139.790 92.250 139.835 ;
        RECT 95.220 139.790 95.510 139.835 ;
        RECT 91.090 139.650 95.510 139.790 ;
        RECT 76.370 139.590 76.690 139.650 ;
        RECT 91.090 139.590 91.410 139.650 ;
        RECT 91.960 139.605 92.250 139.650 ;
        RECT 95.220 139.605 95.510 139.650 ;
        RECT 96.140 139.790 96.430 139.835 ;
        RECT 98.000 139.790 98.290 139.835 ;
        RECT 96.140 139.650 98.290 139.790 ;
        RECT 96.140 139.605 96.430 139.650 ;
        RECT 98.000 139.605 98.290 139.650 ;
        RECT 101.620 139.790 101.910 139.835 ;
        RECT 102.590 139.790 102.910 139.850 ;
        RECT 104.880 139.790 105.170 139.835 ;
        RECT 101.620 139.650 105.170 139.790 ;
        RECT 101.620 139.605 101.910 139.650 ;
        RECT 71.325 139.265 71.615 139.495 ;
        RECT 71.785 139.265 72.075 139.495 ;
        RECT 81.890 139.450 82.210 139.510 ;
        RECT 81.890 139.310 82.405 139.450 ;
        RECT 31.290 139.110 31.610 139.170 ;
        RECT 32.225 139.110 32.515 139.155 ;
        RECT 35.890 139.110 36.210 139.170 ;
        RECT 31.290 138.970 36.210 139.110 ;
        RECT 31.290 138.910 31.610 138.970 ;
        RECT 32.225 138.925 32.515 138.970 ;
        RECT 35.890 138.910 36.210 138.970 ;
        RECT 37.270 139.110 37.590 139.170 ;
        RECT 42.345 139.110 42.635 139.155 ;
        RECT 37.270 138.970 42.635 139.110 ;
        RECT 37.270 138.910 37.590 138.970 ;
        RECT 42.345 138.925 42.635 138.970 ;
        RECT 44.645 138.925 44.935 139.155 ;
        RECT 27.120 138.770 27.410 138.815 ;
        RECT 29.900 138.770 30.190 138.815 ;
        RECT 31.760 138.770 32.050 138.815 ;
        RECT 44.720 138.770 44.860 138.925 ;
        RECT 49.690 138.910 50.010 139.170 ;
        RECT 50.150 139.110 50.470 139.170 ;
        RECT 51.545 139.110 51.835 139.155 ;
        RECT 50.150 138.970 51.835 139.110 ;
        RECT 50.150 138.910 50.470 138.970 ;
        RECT 51.545 138.925 51.835 138.970 ;
        RECT 51.990 138.910 52.310 139.170 ;
        RECT 53.830 138.910 54.150 139.170 ;
        RECT 71.400 139.110 71.540 139.265 ;
        RECT 81.890 139.250 82.210 139.310 ;
        RECT 87.410 139.250 87.730 139.510 ;
        RECT 93.820 139.450 94.110 139.495 ;
        RECT 96.140 139.450 96.355 139.605 ;
        RECT 102.590 139.590 102.910 139.650 ;
        RECT 104.880 139.605 105.170 139.650 ;
        RECT 105.800 139.790 106.090 139.835 ;
        RECT 107.660 139.790 107.950 139.835 ;
        RECT 105.800 139.650 107.950 139.790 ;
        RECT 105.800 139.605 106.090 139.650 ;
        RECT 107.660 139.605 107.950 139.650 ;
        RECT 93.820 139.310 96.355 139.450 ;
        RECT 93.820 139.265 94.110 139.310 ;
        RECT 97.070 139.250 97.390 139.510 ;
        RECT 103.480 139.450 103.770 139.495 ;
        RECT 105.800 139.450 106.015 139.605 ;
        RECT 103.480 139.310 106.015 139.450 ;
        RECT 106.745 139.450 107.035 139.495 ;
        RECT 106.745 139.310 109.260 139.450 ;
        RECT 103.480 139.265 103.770 139.310 ;
        RECT 106.745 139.265 107.035 139.310 ;
        RECT 74.990 139.110 75.310 139.170 ;
        RECT 71.400 138.970 75.310 139.110 ;
        RECT 74.990 138.910 75.310 138.970 ;
        RECT 80.970 138.910 81.290 139.170 ;
        RECT 82.810 138.910 83.130 139.170 ;
        RECT 98.925 139.110 99.215 139.155 ;
        RECT 105.810 139.110 106.130 139.170 ;
        RECT 108.585 139.110 108.875 139.155 ;
        RECT 98.925 138.970 108.875 139.110 ;
        RECT 98.925 138.925 99.215 138.970 ;
        RECT 105.810 138.910 106.130 138.970 ;
        RECT 108.585 138.925 108.875 138.970 ;
        RECT 109.120 138.815 109.260 139.310 ;
        RECT 109.950 139.250 110.270 139.510 ;
        RECT 110.885 139.110 111.175 139.155 ;
        RECT 109.580 138.970 111.175 139.110 ;
        RECT 111.880 139.110 112.020 139.945 ;
        RECT 112.710 139.930 113.030 139.990 ;
        RECT 117.260 139.790 117.550 139.835 ;
        RECT 118.230 139.790 118.550 139.850 ;
        RECT 120.520 139.790 120.810 139.835 ;
        RECT 117.260 139.650 120.810 139.790 ;
        RECT 117.260 139.605 117.550 139.650 ;
        RECT 118.230 139.590 118.550 139.650 ;
        RECT 120.520 139.605 120.810 139.650 ;
        RECT 121.440 139.790 121.730 139.835 ;
        RECT 123.300 139.790 123.590 139.835 ;
        RECT 121.440 139.650 123.590 139.790 ;
        RECT 121.440 139.605 121.730 139.650 ;
        RECT 123.300 139.605 123.590 139.650 ;
        RECT 119.120 139.450 119.410 139.495 ;
        RECT 121.440 139.450 121.655 139.605 ;
        RECT 119.120 139.310 121.655 139.450 ;
        RECT 121.910 139.450 122.230 139.510 ;
        RECT 122.385 139.450 122.675 139.495 ;
        RECT 121.910 139.310 122.675 139.450 ;
        RECT 119.120 139.265 119.410 139.310 ;
        RECT 121.910 139.250 122.230 139.310 ;
        RECT 122.385 139.265 122.675 139.310 ;
        RECT 129.090 139.190 134.150 139.405 ;
        RECT 143.370 139.390 144.510 223.840 ;
        RECT 137.240 139.380 144.510 139.390 ;
        RECT 136.210 139.190 144.510 139.380 ;
        RECT 115.255 139.110 115.545 139.155 ;
        RECT 111.880 138.970 115.545 139.110 ;
        RECT 27.120 138.630 32.050 138.770 ;
        RECT 27.120 138.585 27.410 138.630 ;
        RECT 29.900 138.585 30.190 138.630 ;
        RECT 31.760 138.585 32.050 138.630 ;
        RECT 32.300 138.630 44.860 138.770 ;
        RECT 93.820 138.770 94.110 138.815 ;
        RECT 96.600 138.770 96.890 138.815 ;
        RECT 98.460 138.770 98.750 138.815 ;
        RECT 93.820 138.630 98.750 138.770 ;
        RECT 23.255 138.430 23.545 138.475 ;
        RECT 29.450 138.430 29.770 138.490 ;
        RECT 32.300 138.430 32.440 138.630 ;
        RECT 93.820 138.585 94.110 138.630 ;
        RECT 96.600 138.585 96.890 138.630 ;
        RECT 98.460 138.585 98.750 138.630 ;
        RECT 103.480 138.770 103.770 138.815 ;
        RECT 106.260 138.770 106.550 138.815 ;
        RECT 108.120 138.770 108.410 138.815 ;
        RECT 103.480 138.630 108.410 138.770 ;
        RECT 103.480 138.585 103.770 138.630 ;
        RECT 106.260 138.585 106.550 138.630 ;
        RECT 108.120 138.585 108.410 138.630 ;
        RECT 109.045 138.585 109.335 138.815 ;
        RECT 23.255 138.290 32.440 138.430 ;
        RECT 35.430 138.430 35.750 138.490 ;
        RECT 35.905 138.430 36.195 138.475 ;
        RECT 35.430 138.290 36.195 138.430 ;
        RECT 23.255 138.245 23.545 138.290 ;
        RECT 29.450 138.230 29.770 138.290 ;
        RECT 35.430 138.230 35.750 138.290 ;
        RECT 35.905 138.245 36.195 138.290 ;
        RECT 39.570 138.430 39.890 138.490 ;
        RECT 90.170 138.475 90.490 138.490 ;
        RECT 40.965 138.430 41.255 138.475 ;
        RECT 39.570 138.290 41.255 138.430 ;
        RECT 39.570 138.230 39.890 138.290 ;
        RECT 40.965 138.245 41.255 138.290 ;
        RECT 89.955 138.245 90.490 138.475 ;
        RECT 90.170 138.230 90.490 138.245 ;
        RECT 96.150 138.430 96.470 138.490 ;
        RECT 99.615 138.430 99.905 138.475 ;
        RECT 104.890 138.430 105.210 138.490 ;
        RECT 96.150 138.290 105.210 138.430 ;
        RECT 96.150 138.230 96.470 138.290 ;
        RECT 99.615 138.245 99.905 138.290 ;
        RECT 104.890 138.230 105.210 138.290 ;
        RECT 105.350 138.430 105.670 138.490 ;
        RECT 109.580 138.430 109.720 138.970 ;
        RECT 110.885 138.925 111.175 138.970 ;
        RECT 115.255 138.925 115.545 138.970 ;
        RECT 124.225 139.110 124.515 139.155 ;
        RECT 124.670 139.110 124.990 139.170 ;
        RECT 124.225 138.970 124.990 139.110 ;
        RECT 124.225 138.925 124.515 138.970 ;
        RECT 110.960 138.770 111.100 138.925 ;
        RECT 124.670 138.910 124.990 138.970 ;
        RECT 113.170 138.770 113.490 138.830 ;
        RECT 110.960 138.630 113.490 138.770 ;
        RECT 113.170 138.570 113.490 138.630 ;
        RECT 119.120 138.770 119.410 138.815 ;
        RECT 121.900 138.770 122.190 138.815 ;
        RECT 123.760 138.770 124.050 138.815 ;
        RECT 119.120 138.630 124.050 138.770 ;
        RECT 119.120 138.585 119.410 138.630 ;
        RECT 121.900 138.585 122.190 138.630 ;
        RECT 123.760 138.585 124.050 138.630 ;
        RECT 129.090 138.530 144.510 139.190 ;
        RECT 105.350 138.290 109.720 138.430 ;
        RECT 105.350 138.230 105.670 138.290 ;
        RECT 114.090 138.230 114.410 138.490 ;
        RECT 123.290 138.430 123.610 138.490 ;
        RECT 124.670 138.430 124.990 138.490 ;
        RECT 123.290 138.290 124.990 138.430 ;
        RECT 123.290 138.230 123.610 138.290 ;
        RECT 124.670 138.230 124.990 138.290 ;
        RECT 129.090 138.225 134.150 138.530 ;
        RECT 136.210 138.250 144.510 138.530 ;
        RECT 136.210 138.240 138.350 138.250 ;
        RECT 20.640 137.610 127.820 138.090 ;
        RECT 27.165 137.410 27.455 137.455 ;
        RECT 27.610 137.410 27.930 137.470 ;
        RECT 27.165 137.270 27.930 137.410 ;
        RECT 27.165 137.225 27.455 137.270 ;
        RECT 27.610 137.210 27.930 137.270 ;
        RECT 28.990 137.410 29.310 137.470 ;
        RECT 37.270 137.410 37.590 137.470 ;
        RECT 28.990 137.270 37.590 137.410 ;
        RECT 28.990 137.210 29.310 137.270 ;
        RECT 37.270 137.210 37.590 137.270 ;
        RECT 38.650 137.410 38.970 137.470 ;
        RECT 38.650 137.270 41.640 137.410 ;
        RECT 38.650 137.210 38.970 137.270 ;
        RECT 29.910 136.870 30.230 137.130 ;
        RECT 31.765 137.070 32.055 137.115 ;
        RECT 34.050 137.070 34.370 137.130 ;
        RECT 31.765 136.930 34.370 137.070 ;
        RECT 31.765 136.885 32.055 136.930 ;
        RECT 34.050 136.870 34.370 136.930 ;
        RECT 36.320 137.070 36.610 137.115 ;
        RECT 39.100 137.070 39.390 137.115 ;
        RECT 40.960 137.070 41.250 137.115 ;
        RECT 36.320 136.930 41.250 137.070 ;
        RECT 41.500 137.070 41.640 137.270 ;
        RECT 41.870 137.210 42.190 137.470 ;
        RECT 52.450 137.210 52.770 137.470 ;
        RECT 53.370 137.410 53.690 137.470 ;
        RECT 79.130 137.410 79.450 137.470 ;
        RECT 80.065 137.410 80.355 137.455 ;
        RECT 53.370 137.270 72.920 137.410 ;
        RECT 53.370 137.210 53.690 137.270 ;
        RECT 67.170 137.070 67.490 137.130 ;
        RECT 41.500 136.930 49.460 137.070 ;
        RECT 36.320 136.885 36.610 136.930 ;
        RECT 39.100 136.885 39.390 136.930 ;
        RECT 40.960 136.885 41.250 136.930 ;
        RECT 29.005 136.730 29.295 136.775 ;
        RECT 30.000 136.730 30.140 136.870 ;
        RECT 29.005 136.590 30.140 136.730 ;
        RECT 35.890 136.730 36.210 136.790 ;
        RECT 35.890 136.590 39.340 136.730 ;
        RECT 29.005 136.545 29.295 136.590 ;
        RECT 35.890 136.530 36.210 136.590 ;
        RECT 27.610 136.400 27.930 136.450 ;
        RECT 27.425 136.390 27.930 136.400 ;
        RECT 29.450 136.390 29.770 136.450 ;
        RECT 29.925 136.390 30.215 136.435 ;
        RECT 34.970 136.390 35.290 136.450 ;
        RECT 27.425 136.260 29.220 136.390 ;
        RECT 27.610 136.250 29.220 136.260 ;
        RECT 27.610 136.190 27.930 136.250 ;
        RECT 29.080 136.050 29.220 136.250 ;
        RECT 29.450 136.250 30.215 136.390 ;
        RECT 29.450 136.190 29.770 136.250 ;
        RECT 29.925 136.205 30.215 136.250 ;
        RECT 34.140 136.250 35.290 136.390 ;
        RECT 34.140 136.050 34.280 136.250 ;
        RECT 34.970 136.190 35.290 136.250 ;
        RECT 36.320 136.390 36.610 136.435 ;
        RECT 39.200 136.390 39.340 136.590 ;
        RECT 39.570 136.530 39.890 136.790 ;
        RECT 45.105 136.730 45.395 136.775 ;
        RECT 45.105 136.590 45.780 136.730 ;
        RECT 45.105 136.545 45.395 136.590 ;
        RECT 41.425 136.390 41.715 136.435 ;
        RECT 36.320 136.250 38.855 136.390 ;
        RECT 39.200 136.250 41.715 136.390 ;
        RECT 36.320 136.205 36.610 136.250 ;
        RECT 29.080 135.910 34.280 136.050 ;
        RECT 34.460 136.050 34.750 136.095 ;
        RECT 35.430 136.050 35.750 136.110 ;
        RECT 38.640 136.095 38.855 136.250 ;
        RECT 41.425 136.205 41.715 136.250 ;
        RECT 37.720 136.050 38.010 136.095 ;
        RECT 34.460 135.910 38.010 136.050 ;
        RECT 34.460 135.865 34.750 135.910 ;
        RECT 35.430 135.850 35.750 135.910 ;
        RECT 37.720 135.865 38.010 135.910 ;
        RECT 38.640 136.050 38.930 136.095 ;
        RECT 40.500 136.050 40.790 136.095 ;
        RECT 38.640 135.910 40.790 136.050 ;
        RECT 38.640 135.865 38.930 135.910 ;
        RECT 40.500 135.865 40.790 135.910 ;
        RECT 43.725 136.050 44.015 136.095 ;
        RECT 45.090 136.050 45.410 136.110 ;
        RECT 43.725 135.910 45.410 136.050 ;
        RECT 45.640 136.050 45.780 136.590 ;
        RECT 49.320 136.435 49.460 136.930 ;
        RECT 65.880 136.930 67.490 137.070 ;
        RECT 51.530 136.730 51.850 136.790 ;
        RECT 64.425 136.730 64.715 136.775 ;
        RECT 51.530 136.590 64.715 136.730 ;
        RECT 51.530 136.530 51.850 136.590 ;
        RECT 64.425 136.545 64.715 136.590 ;
        RECT 65.880 136.450 66.020 136.930 ;
        RECT 67.170 136.870 67.490 136.930 ;
        RECT 68.090 136.730 68.410 136.790 ;
        RECT 72.780 136.775 72.920 137.270 ;
        RECT 79.130 137.270 80.355 137.410 ;
        RECT 79.130 137.210 79.450 137.270 ;
        RECT 80.065 137.225 80.355 137.270 ;
        RECT 80.510 137.210 80.830 137.470 ;
        RECT 82.350 137.410 82.670 137.470 ;
        RECT 82.825 137.410 83.115 137.455 ;
        RECT 82.350 137.270 83.115 137.410 ;
        RECT 82.350 137.210 82.670 137.270 ;
        RECT 82.825 137.225 83.115 137.270 ;
        RECT 91.090 137.210 91.410 137.470 ;
        RECT 92.945 137.410 93.235 137.455 ;
        RECT 93.850 137.410 94.170 137.470 ;
        RECT 92.945 137.270 94.170 137.410 ;
        RECT 92.945 137.225 93.235 137.270 ;
        RECT 93.850 137.210 94.170 137.270 ;
        RECT 97.530 137.410 97.850 137.470 ;
        RECT 98.005 137.410 98.295 137.455 ;
        RECT 97.530 137.270 98.295 137.410 ;
        RECT 97.530 137.210 97.850 137.270 ;
        RECT 98.005 137.225 98.295 137.270 ;
        RECT 100.765 137.410 101.055 137.455 ;
        RECT 102.130 137.410 102.450 137.470 ;
        RECT 100.765 137.270 102.450 137.410 ;
        RECT 100.765 137.225 101.055 137.270 ;
        RECT 102.130 137.210 102.450 137.270 ;
        RECT 106.270 137.210 106.590 137.470 ;
        RECT 109.030 137.410 109.350 137.470 ;
        RECT 109.950 137.410 110.270 137.470 ;
        RECT 109.030 137.270 110.270 137.410 ;
        RECT 109.030 137.210 109.350 137.270 ;
        RECT 109.950 137.210 110.270 137.270 ;
        RECT 113.170 137.210 113.490 137.470 ;
        RECT 120.545 137.410 120.835 137.455 ;
        RECT 121.450 137.410 121.770 137.470 ;
        RECT 120.545 137.270 121.770 137.410 ;
        RECT 120.545 137.225 120.835 137.270 ;
        RECT 121.450 137.210 121.770 137.270 ;
        RECT 122.845 137.410 123.135 137.455 ;
        RECT 124.670 137.410 124.990 137.470 ;
        RECT 122.845 137.270 124.990 137.410 ;
        RECT 122.845 137.225 123.135 137.270 ;
        RECT 124.670 137.210 124.990 137.270 ;
        RECT 85.110 137.070 85.430 137.130 ;
        RECT 90.170 137.070 90.490 137.130 ;
        RECT 105.350 137.070 105.670 137.130 ;
        RECT 85.110 136.930 95.920 137.070 ;
        RECT 85.110 136.870 85.430 136.930 ;
        RECT 90.170 136.870 90.490 136.930 ;
        RECT 66.340 136.590 68.410 136.730 ;
        RECT 49.245 136.390 49.535 136.435 ;
        RECT 51.070 136.390 51.390 136.450 ;
        RECT 49.245 136.250 51.390 136.390 ;
        RECT 49.245 136.205 49.535 136.250 ;
        RECT 51.070 136.190 51.390 136.250 ;
        RECT 51.990 136.190 52.310 136.450 ;
        RECT 53.370 136.190 53.690 136.450 ;
        RECT 53.845 136.205 54.135 136.435 ;
        RECT 52.910 136.050 53.230 136.110 ;
        RECT 53.920 136.050 54.060 136.205 ;
        RECT 65.790 136.190 66.110 136.450 ;
        RECT 66.340 136.435 66.480 136.590 ;
        RECT 68.090 136.530 68.410 136.590 ;
        RECT 72.705 136.730 72.995 136.775 ;
        RECT 72.705 136.590 79.360 136.730 ;
        RECT 72.705 136.545 72.995 136.590 ;
        RECT 66.265 136.205 66.555 136.435 ;
        RECT 66.725 136.205 67.015 136.435 ;
        RECT 67.645 136.390 67.935 136.435 ;
        RECT 69.470 136.390 69.790 136.450 ;
        RECT 67.645 136.250 69.790 136.390 ;
        RECT 67.645 136.205 67.935 136.250 ;
        RECT 45.640 135.910 51.760 136.050 ;
        RECT 43.725 135.865 44.015 135.910 ;
        RECT 29.465 135.710 29.755 135.755 ;
        RECT 32.455 135.710 32.745 135.755 ;
        RECT 43.800 135.710 43.940 135.865 ;
        RECT 45.090 135.850 45.410 135.910 ;
        RECT 29.465 135.570 43.940 135.710 ;
        RECT 29.465 135.525 29.755 135.570 ;
        RECT 32.455 135.525 32.745 135.570 ;
        RECT 44.170 135.510 44.490 135.770 ;
        RECT 46.010 135.710 46.330 135.770 ;
        RECT 48.785 135.710 49.075 135.755 ;
        RECT 46.010 135.570 49.075 135.710 ;
        RECT 46.010 135.510 46.330 135.570 ;
        RECT 48.785 135.525 49.075 135.570 ;
        RECT 50.150 135.710 50.470 135.770 ;
        RECT 51.085 135.710 51.375 135.755 ;
        RECT 50.150 135.570 51.375 135.710 ;
        RECT 51.620 135.710 51.760 135.910 ;
        RECT 52.910 135.910 54.060 136.050 ;
        RECT 52.910 135.850 53.230 135.910 ;
        RECT 57.065 135.865 57.355 136.095 ;
        RECT 66.800 136.050 66.940 136.205 ;
        RECT 69.470 136.190 69.790 136.250 ;
        RECT 73.610 136.190 73.930 136.450 ;
        RECT 78.670 136.190 78.990 136.450 ;
        RECT 79.220 136.435 79.360 136.590 ;
        RECT 82.350 136.530 82.670 136.790 ;
        RECT 86.030 136.730 86.350 136.790 ;
        RECT 95.780 136.775 95.920 136.930 ;
        RECT 99.000 136.930 105.670 137.070 ;
        RECT 86.030 136.590 92.240 136.730 ;
        RECT 86.030 136.530 86.350 136.590 ;
        RECT 79.145 136.390 79.435 136.435 ;
        RECT 81.445 136.390 81.735 136.435 ;
        RECT 81.890 136.390 82.210 136.450 ;
        RECT 83.745 136.390 84.035 136.435 ;
        RECT 79.145 136.250 84.035 136.390 ;
        RECT 79.145 136.205 79.435 136.250 ;
        RECT 81.445 136.205 81.735 136.250 ;
        RECT 81.890 136.190 82.210 136.250 ;
        RECT 83.745 136.205 84.035 136.250 ;
        RECT 84.650 136.190 84.970 136.450 ;
        RECT 85.110 136.190 85.430 136.450 ;
        RECT 87.410 136.390 87.730 136.450 ;
        RECT 90.630 136.390 90.950 136.450 ;
        RECT 92.100 136.435 92.240 136.590 ;
        RECT 94.785 136.545 95.075 136.775 ;
        RECT 95.705 136.545 95.995 136.775 ;
        RECT 87.410 136.250 90.950 136.390 ;
        RECT 87.410 136.190 87.730 136.250 ;
        RECT 90.630 136.190 90.950 136.250 ;
        RECT 92.025 136.205 92.315 136.435 ;
        RECT 94.860 136.390 95.000 136.545 ;
        RECT 99.000 136.390 99.140 136.930 ;
        RECT 105.350 136.870 105.670 136.930 ;
        RECT 99.830 136.530 100.150 136.790 ;
        RECT 106.745 136.730 107.035 136.775 ;
        RECT 108.570 136.730 108.890 136.790 ;
        RECT 111.330 136.730 111.650 136.790 ;
        RECT 106.745 136.590 108.890 136.730 ;
        RECT 106.745 136.545 107.035 136.590 ;
        RECT 108.570 136.530 108.890 136.590 ;
        RECT 109.580 136.590 111.650 136.730 ;
        RECT 94.860 136.250 99.140 136.390 ;
        RECT 68.550 136.050 68.870 136.110 ;
        RECT 66.800 135.910 68.870 136.050 ;
        RECT 55.670 135.710 55.990 135.770 ;
        RECT 51.620 135.570 55.990 135.710 ;
        RECT 57.140 135.710 57.280 135.865 ;
        RECT 68.550 135.850 68.870 135.910 ;
        RECT 86.950 136.050 87.270 136.110 ;
        RECT 94.860 136.050 95.000 136.250 ;
        RECT 99.370 136.190 99.690 136.450 ;
        RECT 100.750 136.190 101.070 136.450 ;
        RECT 109.580 136.435 109.720 136.590 ;
        RECT 111.330 136.530 111.650 136.590 ;
        RECT 113.185 136.730 113.475 136.775 ;
        RECT 114.550 136.730 114.870 136.790 ;
        RECT 113.185 136.590 114.870 136.730 ;
        RECT 113.185 136.545 113.475 136.590 ;
        RECT 114.550 136.530 114.870 136.590 ;
        RECT 116.390 136.730 116.710 136.790 ;
        RECT 116.390 136.590 122.140 136.730 ;
        RECT 116.390 136.530 116.710 136.590 ;
        RECT 105.825 136.205 106.115 136.435 ;
        RECT 109.045 136.205 109.335 136.435 ;
        RECT 109.505 136.205 109.795 136.435 ;
        RECT 86.950 135.910 95.000 136.050 ;
        RECT 86.950 135.850 87.270 135.910 ;
        RECT 96.150 135.850 96.470 136.110 ;
        RECT 105.900 136.050 106.040 136.205 ;
        RECT 106.730 136.050 107.050 136.110 ;
        RECT 105.900 135.910 107.050 136.050 ;
        RECT 106.730 135.850 107.050 135.910 ;
        RECT 107.205 136.050 107.495 136.095 ;
        RECT 107.665 136.050 107.955 136.095 ;
        RECT 107.205 135.910 107.955 136.050 ;
        RECT 109.120 136.050 109.260 136.205 ;
        RECT 109.950 136.190 110.270 136.450 ;
        RECT 110.885 136.205 111.175 136.435 ;
        RECT 110.410 136.050 110.730 136.110 ;
        RECT 109.120 135.910 110.730 136.050 ;
        RECT 107.205 135.865 107.495 135.910 ;
        RECT 107.665 135.865 107.955 135.910 ;
        RECT 110.410 135.850 110.730 135.910 ;
        RECT 73.610 135.710 73.930 135.770 ;
        RECT 57.140 135.570 73.930 135.710 ;
        RECT 50.150 135.510 50.470 135.570 ;
        RECT 51.085 135.525 51.375 135.570 ;
        RECT 55.670 135.510 55.990 135.570 ;
        RECT 73.610 135.510 73.930 135.570 ;
        RECT 86.030 135.510 86.350 135.770 ;
        RECT 98.450 135.510 98.770 135.770 ;
        RECT 104.905 135.710 105.195 135.755 ;
        RECT 105.350 135.710 105.670 135.770 ;
        RECT 104.905 135.570 105.670 135.710 ;
        RECT 104.905 135.525 105.195 135.570 ;
        RECT 105.350 135.510 105.670 135.570 ;
        RECT 108.110 135.710 108.430 135.770 ;
        RECT 110.960 135.710 111.100 136.205 ;
        RECT 112.250 136.190 112.570 136.450 ;
        RECT 113.630 136.190 113.950 136.450 ;
        RECT 114.090 136.390 114.410 136.450 ;
        RECT 122.000 136.435 122.140 136.590 ;
        RECT 119.625 136.390 119.915 136.435 ;
        RECT 114.090 136.250 119.915 136.390 ;
        RECT 114.090 136.190 114.410 136.250 ;
        RECT 119.625 136.205 119.915 136.250 ;
        RECT 121.925 136.205 122.215 136.435 ;
        RECT 108.110 135.570 111.100 135.710 ;
        RECT 108.110 135.510 108.430 135.570 ;
        RECT 111.330 135.510 111.650 135.770 ;
        RECT 20.640 134.890 127.820 135.370 ;
        RECT 22.335 134.690 22.625 134.735 ;
        RECT 28.990 134.690 29.310 134.750 ;
        RECT 22.335 134.550 29.310 134.690 ;
        RECT 22.335 134.505 22.625 134.550 ;
        RECT 28.990 134.490 29.310 134.550 ;
        RECT 34.525 134.690 34.815 134.735 ;
        RECT 34.970 134.690 35.290 134.750 ;
        RECT 39.110 134.690 39.430 134.750 ;
        RECT 51.530 134.690 51.850 134.750 ;
        RECT 34.525 134.550 35.290 134.690 ;
        RECT 34.525 134.505 34.815 134.550 ;
        RECT 34.970 134.490 35.290 134.550 ;
        RECT 35.520 134.550 39.430 134.690 ;
        RECT 24.340 134.350 24.630 134.395 ;
        RECT 26.690 134.350 27.010 134.410 ;
        RECT 27.600 134.350 27.890 134.395 ;
        RECT 24.340 134.210 27.890 134.350 ;
        RECT 24.340 134.165 24.630 134.210 ;
        RECT 26.690 134.150 27.010 134.210 ;
        RECT 27.600 134.165 27.890 134.210 ;
        RECT 28.520 134.350 28.810 134.395 ;
        RECT 30.380 134.350 30.670 134.395 ;
        RECT 28.520 134.210 30.670 134.350 ;
        RECT 28.520 134.165 28.810 134.210 ;
        RECT 30.380 134.165 30.670 134.210 ;
        RECT 26.200 134.010 26.490 134.055 ;
        RECT 28.520 134.010 28.735 134.165 ;
        RECT 26.200 133.870 28.735 134.010 ;
        RECT 31.290 134.010 31.610 134.070 ;
        RECT 32.685 134.010 32.975 134.055 ;
        RECT 34.050 134.010 34.370 134.070 ;
        RECT 35.520 134.055 35.660 134.550 ;
        RECT 39.110 134.490 39.430 134.550 ;
        RECT 41.960 134.550 51.850 134.690 ;
        RECT 41.960 134.395 42.100 134.550 ;
        RECT 51.530 134.490 51.850 134.550 ;
        RECT 51.990 134.690 52.310 134.750 ;
        RECT 52.465 134.690 52.755 134.735 ;
        RECT 51.990 134.550 52.755 134.690 ;
        RECT 51.990 134.490 52.310 134.550 ;
        RECT 52.465 134.505 52.755 134.550 ;
        RECT 57.510 134.690 57.830 134.750 ;
        RECT 60.285 134.690 60.575 134.735 ;
        RECT 57.510 134.550 60.575 134.690 ;
        RECT 57.510 134.490 57.830 134.550 ;
        RECT 60.285 134.505 60.575 134.550 ;
        RECT 68.090 134.490 68.410 134.750 ;
        RECT 109.045 134.690 109.335 134.735 ;
        RECT 109.490 134.690 109.810 134.750 ;
        RECT 71.400 134.550 107.880 134.690 ;
        RECT 36.825 134.350 37.115 134.395 ;
        RECT 36.825 134.210 41.640 134.350 ;
        RECT 36.825 134.165 37.115 134.210 ;
        RECT 31.290 133.870 32.440 134.010 ;
        RECT 26.200 133.825 26.490 133.870 ;
        RECT 31.290 133.810 31.610 133.870 ;
        RECT 29.465 133.670 29.755 133.715 ;
        RECT 32.300 133.670 32.440 133.870 ;
        RECT 32.685 133.870 34.370 134.010 ;
        RECT 32.685 133.825 32.975 133.870 ;
        RECT 34.050 133.810 34.370 133.870 ;
        RECT 35.445 133.825 35.735 134.055 ;
        RECT 38.205 134.010 38.495 134.055 ;
        RECT 35.980 133.870 38.495 134.010 ;
        RECT 35.980 133.730 36.120 133.870 ;
        RECT 38.205 133.825 38.495 133.870 ;
        RECT 40.490 133.810 40.810 134.070 ;
        RECT 41.500 134.010 41.640 134.210 ;
        RECT 41.885 134.165 42.175 134.395 ;
        RECT 43.250 134.150 43.570 134.410 ;
        RECT 64.885 134.350 65.175 134.395 ;
        RECT 68.180 134.350 68.320 134.490 ;
        RECT 71.400 134.395 71.540 134.550 ;
        RECT 71.325 134.350 71.615 134.395 ;
        RECT 50.700 134.210 65.175 134.350 ;
        RECT 50.700 134.010 50.840 134.210 ;
        RECT 64.885 134.165 65.175 134.210 ;
        RECT 66.800 134.210 68.320 134.350 ;
        RECT 70.020 134.210 71.615 134.350 ;
        RECT 54.305 134.010 54.595 134.055 ;
        RECT 41.500 133.870 50.840 134.010 ;
        RECT 51.160 133.870 54.595 134.010 ;
        RECT 35.890 133.670 36.210 133.730 ;
        RECT 29.465 133.530 31.980 133.670 ;
        RECT 32.300 133.530 36.210 133.670 ;
        RECT 29.465 133.485 29.755 133.530 ;
        RECT 31.840 133.375 31.980 133.530 ;
        RECT 35.890 133.470 36.210 133.530 ;
        RECT 36.350 133.470 36.670 133.730 ;
        RECT 37.730 133.670 38.050 133.730 ;
        RECT 40.965 133.670 41.255 133.715 ;
        RECT 37.730 133.530 41.255 133.670 ;
        RECT 37.730 133.470 38.050 133.530 ;
        RECT 40.965 133.485 41.255 133.530 ;
        RECT 44.170 133.670 44.490 133.730 ;
        RECT 49.690 133.670 50.010 133.730 ;
        RECT 51.160 133.670 51.300 133.870 ;
        RECT 54.305 133.825 54.595 133.870 ;
        RECT 56.130 134.010 56.450 134.070 ;
        RECT 57.525 134.010 57.815 134.055 ;
        RECT 56.130 133.870 57.815 134.010 ;
        RECT 56.130 133.810 56.450 133.870 ;
        RECT 57.525 133.825 57.815 133.870 ;
        RECT 60.270 134.010 60.590 134.070 ;
        RECT 60.745 134.010 61.035 134.055 ;
        RECT 60.270 133.870 61.035 134.010 ;
        RECT 60.270 133.810 60.590 133.870 ;
        RECT 60.745 133.825 61.035 133.870 ;
        RECT 65.790 134.010 66.110 134.070 ;
        RECT 66.800 134.055 66.940 134.210 ;
        RECT 66.265 134.010 66.555 134.055 ;
        RECT 65.790 133.870 66.555 134.010 ;
        RECT 65.790 133.810 66.110 133.870 ;
        RECT 66.265 133.825 66.555 133.870 ;
        RECT 66.725 133.825 67.015 134.055 ;
        RECT 67.170 133.810 67.490 134.070 ;
        RECT 68.105 134.010 68.395 134.055 ;
        RECT 69.470 134.010 69.790 134.070 ;
        RECT 68.105 133.870 69.790 134.010 ;
        RECT 68.105 133.825 68.395 133.870 ;
        RECT 69.470 133.810 69.790 133.870 ;
        RECT 44.170 133.530 51.300 133.670 ;
        RECT 52.910 133.670 53.230 133.730 ;
        RECT 54.765 133.670 55.055 133.715 ;
        RECT 52.910 133.530 55.055 133.670 ;
        RECT 44.170 133.470 44.490 133.530 ;
        RECT 49.690 133.470 50.010 133.530 ;
        RECT 52.910 133.470 53.230 133.530 ;
        RECT 54.765 133.485 55.055 133.530 ;
        RECT 55.670 133.470 55.990 133.730 ;
        RECT 59.810 133.470 60.130 133.730 ;
        RECT 26.200 133.330 26.490 133.375 ;
        RECT 28.980 133.330 29.270 133.375 ;
        RECT 30.840 133.330 31.130 133.375 ;
        RECT 26.200 133.190 31.130 133.330 ;
        RECT 26.200 133.145 26.490 133.190 ;
        RECT 28.980 133.145 29.270 133.190 ;
        RECT 30.840 133.145 31.130 133.190 ;
        RECT 31.765 133.145 32.055 133.375 ;
        RECT 34.510 133.330 34.830 133.390 ;
        RECT 42.330 133.330 42.650 133.390 ;
        RECT 70.020 133.330 70.160 134.210 ;
        RECT 71.325 134.165 71.615 134.210 ;
        RECT 72.245 134.350 72.535 134.395 ;
        RECT 73.150 134.350 73.470 134.410 ;
        RECT 76.830 134.350 77.150 134.410 ;
        RECT 80.920 134.350 81.210 134.395 ;
        RECT 84.180 134.350 84.470 134.395 ;
        RECT 72.245 134.210 74.300 134.350 ;
        RECT 72.245 134.165 72.535 134.210 ;
        RECT 73.150 134.150 73.470 134.210 ;
        RECT 74.160 134.055 74.300 134.210 ;
        RECT 76.830 134.210 84.470 134.350 ;
        RECT 76.830 134.150 77.150 134.210 ;
        RECT 80.920 134.165 81.210 134.210 ;
        RECT 84.180 134.165 84.470 134.210 ;
        RECT 85.100 134.350 85.390 134.395 ;
        RECT 86.960 134.350 87.250 134.395 ;
        RECT 85.100 134.210 87.250 134.350 ;
        RECT 85.100 134.165 85.390 134.210 ;
        RECT 86.960 134.165 87.250 134.210 ;
        RECT 74.085 133.825 74.375 134.055 ;
        RECT 82.780 134.010 83.070 134.055 ;
        RECT 85.100 134.010 85.315 134.165 ;
        RECT 82.780 133.870 85.315 134.010 ;
        RECT 82.780 133.825 83.070 133.870 ;
        RECT 86.030 133.810 86.350 134.070 ;
        RECT 107.190 134.010 107.510 134.070 ;
        RECT 107.740 134.055 107.880 134.550 ;
        RECT 109.045 134.550 109.810 134.690 ;
        RECT 109.045 134.505 109.335 134.550 ;
        RECT 109.490 134.490 109.810 134.550 ;
        RECT 111.790 134.490 112.110 134.750 ;
        RECT 135.660 134.480 136.800 134.510 ;
        RECT 108.585 134.350 108.875 134.395 ;
        RECT 110.870 134.350 111.190 134.410 ;
        RECT 108.585 134.210 111.190 134.350 ;
        RECT 108.585 134.165 108.875 134.210 ;
        RECT 110.870 134.150 111.190 134.210 ;
        RECT 107.665 134.010 107.955 134.055 ;
        RECT 109.965 134.010 110.255 134.055 ;
        RECT 112.250 134.010 112.570 134.070 ;
        RECT 112.725 134.010 113.015 134.055 ;
        RECT 107.190 133.870 113.015 134.010 ;
        RECT 107.190 133.810 107.510 133.870 ;
        RECT 107.665 133.825 107.955 133.870 ;
        RECT 109.965 133.825 110.255 133.870 ;
        RECT 112.250 133.810 112.570 133.870 ;
        RECT 112.725 133.825 113.015 133.870 ;
        RECT 74.990 133.470 75.310 133.730 ;
        RECT 87.870 133.470 88.190 133.730 ;
        RECT 106.745 133.670 107.035 133.715 ;
        RECT 110.410 133.670 110.730 133.730 ;
        RECT 106.745 133.530 110.730 133.670 ;
        RECT 106.745 133.485 107.035 133.530 ;
        RECT 110.410 133.470 110.730 133.530 ;
        RECT 110.870 133.470 111.190 133.730 ;
        RECT 113.645 133.670 113.935 133.715 ;
        RECT 112.800 133.530 113.935 133.670 ;
        RECT 112.800 133.390 112.940 133.530 ;
        RECT 113.645 133.485 113.935 133.530 ;
        RECT 135.590 133.400 136.850 134.480 ;
        RECT 34.510 133.190 40.720 133.330 ;
        RECT 34.510 133.130 34.830 133.190 ;
        RECT 36.350 132.790 36.670 133.050 ;
        RECT 37.730 132.990 38.050 133.050 ;
        RECT 40.580 133.035 40.720 133.190 ;
        RECT 42.330 133.190 70.160 133.330 ;
        RECT 82.780 133.330 83.070 133.375 ;
        RECT 85.560 133.330 85.850 133.375 ;
        RECT 87.420 133.330 87.710 133.375 ;
        RECT 82.780 133.190 87.710 133.330 ;
        RECT 42.330 133.130 42.650 133.190 ;
        RECT 82.780 133.145 83.070 133.190 ;
        RECT 85.560 133.145 85.850 133.190 ;
        RECT 87.420 133.145 87.710 133.190 ;
        RECT 112.710 133.130 113.030 133.390 ;
        RECT 39.585 132.990 39.875 133.035 ;
        RECT 37.730 132.850 39.875 132.990 ;
        RECT 37.730 132.790 38.050 132.850 ;
        RECT 39.585 132.805 39.875 132.850 ;
        RECT 40.505 132.805 40.795 133.035 ;
        RECT 49.690 132.790 50.010 133.050 ;
        RECT 51.070 132.990 51.390 133.050 ;
        RECT 56.605 132.990 56.895 133.035 ;
        RECT 51.070 132.850 56.895 132.990 ;
        RECT 51.070 132.790 51.390 132.850 ;
        RECT 56.605 132.805 56.895 132.850 ;
        RECT 61.190 132.990 61.510 133.050 ;
        RECT 62.585 132.990 62.875 133.035 ;
        RECT 61.190 132.850 62.875 132.990 ;
        RECT 61.190 132.790 61.510 132.850 ;
        RECT 62.585 132.805 62.875 132.850 ;
        RECT 73.165 132.990 73.455 133.035 ;
        RECT 73.610 132.990 73.930 133.050 ;
        RECT 79.130 133.035 79.450 133.050 ;
        RECT 73.165 132.850 73.930 132.990 ;
        RECT 73.165 132.805 73.455 132.850 ;
        RECT 73.610 132.790 73.930 132.850 ;
        RECT 78.915 132.990 79.450 133.035 ;
        RECT 84.190 132.990 84.510 133.050 ;
        RECT 78.915 132.850 84.510 132.990 ;
        RECT 78.915 132.805 79.450 132.850 ;
        RECT 79.130 132.790 79.450 132.805 ;
        RECT 84.190 132.790 84.510 132.850 ;
        RECT 20.640 132.170 127.820 132.650 ;
        RECT 26.245 131.970 26.535 132.015 ;
        RECT 26.690 131.970 27.010 132.030 ;
        RECT 26.245 131.830 27.010 131.970 ;
        RECT 26.245 131.785 26.535 131.830 ;
        RECT 26.690 131.770 27.010 131.830 ;
        RECT 30.845 131.970 31.135 132.015 ;
        RECT 34.050 131.970 34.370 132.030 ;
        RECT 30.845 131.830 34.370 131.970 ;
        RECT 30.845 131.785 31.135 131.830 ;
        RECT 34.050 131.770 34.370 131.830 ;
        RECT 40.735 131.970 41.025 132.015 ;
        RECT 44.170 131.970 44.490 132.030 ;
        RECT 40.735 131.830 44.490 131.970 ;
        RECT 40.735 131.785 41.025 131.830 ;
        RECT 44.170 131.770 44.490 131.830 ;
        RECT 56.130 131.770 56.450 132.030 ;
        RECT 76.830 131.770 77.150 132.030 ;
        RECT 85.110 131.970 85.430 132.030 ;
        RECT 85.585 131.970 85.875 132.015 ;
        RECT 85.110 131.830 85.875 131.970 ;
        RECT 85.110 131.770 85.430 131.830 ;
        RECT 85.585 131.785 85.875 131.830 ;
        RECT 106.270 131.770 106.590 132.030 ;
        RECT 44.600 131.630 44.890 131.675 ;
        RECT 47.380 131.630 47.670 131.675 ;
        RECT 49.240 131.630 49.530 131.675 ;
        RECT 44.600 131.490 49.530 131.630 ;
        RECT 44.600 131.445 44.890 131.490 ;
        RECT 47.380 131.445 47.670 131.490 ;
        RECT 49.240 131.445 49.530 131.490 ;
        RECT 49.690 131.630 50.010 131.690 ;
        RECT 59.810 131.630 60.130 131.690 ;
        RECT 63.490 131.630 63.810 131.690 ;
        RECT 84.190 131.630 84.510 131.690 ;
        RECT 49.690 131.490 59.120 131.630 ;
        RECT 49.690 131.430 50.010 131.490 ;
        RECT 28.085 131.105 28.375 131.335 ;
        RECT 28.545 131.290 28.835 131.335 ;
        RECT 29.450 131.290 29.770 131.350 ;
        RECT 28.545 131.150 29.770 131.290 ;
        RECT 28.545 131.105 28.835 131.150 ;
        RECT 26.690 130.750 27.010 131.010 ;
        RECT 28.160 130.610 28.300 131.105 ;
        RECT 29.450 131.090 29.770 131.150 ;
        RECT 31.290 131.090 31.610 131.350 ;
        RECT 47.865 131.290 48.155 131.335 ;
        RECT 50.150 131.290 50.470 131.350 ;
        RECT 47.865 131.150 50.470 131.290 ;
        RECT 47.865 131.105 48.155 131.150 ;
        RECT 50.150 131.090 50.470 131.150 ;
        RECT 28.990 130.750 29.310 131.010 ;
        RECT 40.045 130.950 40.335 130.995 ;
        RECT 43.250 130.950 43.570 131.010 ;
        RECT 40.045 130.810 43.570 130.950 ;
        RECT 40.045 130.765 40.335 130.810 ;
        RECT 43.250 130.750 43.570 130.810 ;
        RECT 44.600 130.950 44.890 130.995 ;
        RECT 49.705 130.950 49.995 130.995 ;
        RECT 50.700 130.950 50.840 131.490 ;
        RECT 51.530 131.290 51.850 131.350 ;
        RECT 53.385 131.290 53.675 131.335 ;
        RECT 55.670 131.290 55.990 131.350 ;
        RECT 51.530 131.150 55.990 131.290 ;
        RECT 51.530 131.090 51.850 131.150 ;
        RECT 53.385 131.105 53.675 131.150 ;
        RECT 55.670 131.090 55.990 131.150 ;
        RECT 44.600 130.810 47.135 130.950 ;
        RECT 44.600 130.765 44.890 130.810 ;
        RECT 29.910 130.610 30.230 130.670 ;
        RECT 46.010 130.655 46.330 130.670 ;
        RECT 28.160 130.470 30.230 130.610 ;
        RECT 29.910 130.410 30.230 130.470 ;
        RECT 42.740 130.610 43.030 130.655 ;
        RECT 46.000 130.610 46.330 130.655 ;
        RECT 42.740 130.470 46.330 130.610 ;
        RECT 42.740 130.425 43.030 130.470 ;
        RECT 46.000 130.425 46.330 130.470 ;
        RECT 46.920 130.655 47.135 130.810 ;
        RECT 49.705 130.810 50.840 130.950 ;
        RECT 49.705 130.765 49.995 130.810 ;
        RECT 51.990 130.750 52.310 131.010 ;
        RECT 58.980 130.995 59.120 131.490 ;
        RECT 59.810 131.490 68.780 131.630 ;
        RECT 59.810 131.430 60.130 131.490 ;
        RECT 63.490 131.430 63.810 131.490 ;
        RECT 61.190 131.290 61.510 131.350 ;
        RECT 68.640 131.335 68.780 131.490 ;
        RECT 84.190 131.490 96.380 131.630 ;
        RECT 84.190 131.430 84.510 131.490 ;
        RECT 61.190 131.150 64.640 131.290 ;
        RECT 61.190 131.090 61.510 131.150 ;
        RECT 58.905 130.950 59.195 130.995 ;
        RECT 63.950 130.950 64.270 131.010 ;
        RECT 64.500 130.995 64.640 131.150 ;
        RECT 68.565 131.105 68.855 131.335 ;
        RECT 72.690 131.290 73.010 131.350 ;
        RECT 75.005 131.290 75.295 131.335 ;
        RECT 80.985 131.290 81.275 131.335 ;
        RECT 82.825 131.290 83.115 131.335 ;
        RECT 72.690 131.150 74.760 131.290 ;
        RECT 72.690 131.090 73.010 131.150 ;
        RECT 58.905 130.810 64.270 130.950 ;
        RECT 58.905 130.765 59.195 130.810 ;
        RECT 63.950 130.750 64.270 130.810 ;
        RECT 64.425 130.765 64.715 130.995 ;
        RECT 66.710 130.950 67.030 131.010 ;
        RECT 69.485 130.950 69.775 130.995 ;
        RECT 66.710 130.810 69.775 130.950 ;
        RECT 66.710 130.750 67.030 130.810 ;
        RECT 69.485 130.765 69.775 130.810 ;
        RECT 73.610 130.750 73.930 131.010 ;
        RECT 74.620 130.950 74.760 131.150 ;
        RECT 75.005 131.150 83.115 131.290 ;
        RECT 75.005 131.105 75.295 131.150 ;
        RECT 80.985 131.105 81.275 131.150 ;
        RECT 82.825 131.105 83.115 131.150 ;
        RECT 76.370 130.950 76.690 131.010 ;
        RECT 74.620 130.810 76.690 130.950 ;
        RECT 76.370 130.750 76.690 130.810 ;
        RECT 82.900 130.670 83.040 131.105 ;
        RECT 83.745 130.950 84.035 130.995 ;
        RECT 84.280 130.950 84.420 131.430 ;
        RECT 95.690 131.290 96.010 131.350 ;
        RECT 96.240 131.335 96.380 131.490 ;
        RECT 98.465 131.445 98.755 131.675 ;
        RECT 114.105 131.630 114.395 131.675 ;
        RECT 114.105 131.490 119.610 131.630 ;
        RECT 114.105 131.445 114.395 131.490 ;
        RECT 83.745 130.810 84.420 130.950 ;
        RECT 84.740 131.150 96.010 131.290 ;
        RECT 83.745 130.765 84.035 130.810 ;
        RECT 46.920 130.610 47.210 130.655 ;
        RECT 48.780 130.610 49.070 130.655 ;
        RECT 46.920 130.470 49.070 130.610 ;
        RECT 46.920 130.425 47.210 130.470 ;
        RECT 48.780 130.425 49.070 130.470 ;
        RECT 52.450 130.610 52.770 130.670 ;
        RECT 53.830 130.610 54.150 130.670 ;
        RECT 52.450 130.470 54.150 130.610 ;
        RECT 46.010 130.410 46.330 130.425 ;
        RECT 52.450 130.410 52.770 130.470 ;
        RECT 53.830 130.410 54.150 130.470 ;
        RECT 80.065 130.610 80.355 130.655 ;
        RECT 80.510 130.610 80.830 130.670 ;
        RECT 80.065 130.470 80.830 130.610 ;
        RECT 80.065 130.425 80.355 130.470 ;
        RECT 80.510 130.410 80.830 130.470 ;
        RECT 82.810 130.610 83.130 130.670 ;
        RECT 84.740 130.610 84.880 131.150 ;
        RECT 95.690 131.090 96.010 131.150 ;
        RECT 96.165 131.105 96.455 131.335 ;
        RECT 90.630 130.950 90.950 131.010 ;
        RECT 93.405 130.950 93.695 130.995 ;
        RECT 90.630 130.810 93.695 130.950 ;
        RECT 98.540 130.950 98.680 131.445 ;
        RECT 103.050 131.290 103.370 131.350 ;
        RECT 111.345 131.290 111.635 131.335 ;
        RECT 113.630 131.290 113.950 131.350 ;
        RECT 103.050 131.150 107.420 131.290 ;
        RECT 103.050 131.090 103.370 131.150 ;
        RECT 107.280 131.010 107.420 131.150 ;
        RECT 111.345 131.150 113.950 131.290 ;
        RECT 119.470 131.290 119.610 131.490 ;
        RECT 119.470 131.150 120.760 131.290 ;
        RECT 111.345 131.105 111.635 131.150 ;
        RECT 113.630 131.090 113.950 131.150 ;
        RECT 99.845 130.950 100.135 130.995 ;
        RECT 98.540 130.810 100.135 130.950 ;
        RECT 90.630 130.750 90.950 130.810 ;
        RECT 93.405 130.765 93.695 130.810 ;
        RECT 99.845 130.765 100.135 130.810 ;
        RECT 105.365 130.950 105.655 130.995 ;
        RECT 105.810 130.950 106.130 131.010 ;
        RECT 105.365 130.810 106.130 130.950 ;
        RECT 105.365 130.765 105.655 130.810 ;
        RECT 105.810 130.750 106.130 130.810 ;
        RECT 107.190 130.750 107.510 131.010 ;
        RECT 108.125 130.950 108.415 130.995 ;
        RECT 109.490 130.950 109.810 131.010 ;
        RECT 108.125 130.810 109.810 130.950 ;
        RECT 108.125 130.765 108.415 130.810 ;
        RECT 109.490 130.750 109.810 130.810 ;
        RECT 116.850 130.950 117.170 131.010 ;
        RECT 120.620 130.995 120.760 131.150 ;
        RECT 118.245 130.950 118.535 130.995 ;
        RECT 116.850 130.810 118.535 130.950 ;
        RECT 116.850 130.750 117.170 130.810 ;
        RECT 118.245 130.765 118.535 130.810 ;
        RECT 120.545 130.765 120.835 130.995 ;
        RECT 82.810 130.470 84.880 130.610 ;
        RECT 93.865 130.610 94.155 130.655 ;
        RECT 96.150 130.610 96.470 130.670 ;
        RECT 93.865 130.470 96.470 130.610 ;
        RECT 82.810 130.410 83.130 130.470 ;
        RECT 93.865 130.425 94.155 130.470 ;
        RECT 96.150 130.410 96.470 130.470 ;
        RECT 96.610 130.610 96.930 130.670 ;
        RECT 110.870 130.610 111.190 130.670 ;
        RECT 111.805 130.610 112.095 130.655 ;
        RECT 96.610 130.470 112.095 130.610 ;
        RECT 96.610 130.410 96.930 130.470 ;
        RECT 110.870 130.410 111.190 130.470 ;
        RECT 111.805 130.425 112.095 130.470 ;
        RECT 49.230 130.270 49.550 130.330 ;
        RECT 51.545 130.270 51.835 130.315 ;
        RECT 49.230 130.130 51.835 130.270 ;
        RECT 49.230 130.070 49.550 130.130 ;
        RECT 51.545 130.085 51.835 130.130 ;
        RECT 52.910 130.270 53.230 130.330 ;
        RECT 54.305 130.270 54.595 130.315 ;
        RECT 52.910 130.130 54.595 130.270 ;
        RECT 52.910 130.070 53.230 130.130 ;
        RECT 54.305 130.085 54.595 130.130 ;
        RECT 60.730 130.270 61.050 130.330 ;
        RECT 63.505 130.270 63.795 130.315 ;
        RECT 60.730 130.130 63.795 130.270 ;
        RECT 60.730 130.070 61.050 130.130 ;
        RECT 63.505 130.085 63.795 130.130 ;
        RECT 67.170 130.270 67.490 130.330 ;
        RECT 69.945 130.270 70.235 130.315 ;
        RECT 67.170 130.130 70.235 130.270 ;
        RECT 67.170 130.070 67.490 130.130 ;
        RECT 69.945 130.085 70.235 130.130 ;
        RECT 71.785 130.270 72.075 130.315 ;
        RECT 72.690 130.270 73.010 130.330 ;
        RECT 71.785 130.130 73.010 130.270 ;
        RECT 71.785 130.085 72.075 130.130 ;
        RECT 72.690 130.070 73.010 130.130 ;
        RECT 74.530 130.270 74.850 130.330 ;
        RECT 77.765 130.270 78.055 130.315 ;
        RECT 74.530 130.130 78.055 130.270 ;
        RECT 74.530 130.070 74.850 130.130 ;
        RECT 77.765 130.085 78.055 130.130 ;
        RECT 79.605 130.270 79.895 130.315 ;
        RECT 82.350 130.270 82.670 130.330 ;
        RECT 83.285 130.270 83.575 130.315 ;
        RECT 83.730 130.270 84.050 130.330 ;
        RECT 79.605 130.130 84.050 130.270 ;
        RECT 79.605 130.085 79.895 130.130 ;
        RECT 82.350 130.070 82.670 130.130 ;
        RECT 83.285 130.085 83.575 130.130 ;
        RECT 83.730 130.070 84.050 130.130 ;
        RECT 94.310 130.270 94.630 130.330 ;
        RECT 98.925 130.270 99.215 130.315 ;
        RECT 94.310 130.130 99.215 130.270 ;
        RECT 94.310 130.070 94.630 130.130 ;
        RECT 98.925 130.085 99.215 130.130 ;
        RECT 112.265 130.270 112.555 130.315 ;
        RECT 112.710 130.270 113.030 130.330 ;
        RECT 112.265 130.130 113.030 130.270 ;
        RECT 112.265 130.085 112.555 130.130 ;
        RECT 112.710 130.070 113.030 130.130 ;
        RECT 118.690 130.070 119.010 130.330 ;
        RECT 121.465 130.270 121.755 130.315 ;
        RECT 122.830 130.270 123.150 130.330 ;
        RECT 121.465 130.130 123.150 130.270 ;
        RECT 121.465 130.085 121.755 130.130 ;
        RECT 122.830 130.070 123.150 130.130 ;
        RECT 20.640 129.450 127.820 129.930 ;
        RECT 34.510 129.050 34.830 129.310 ;
        RECT 36.810 129.050 37.130 129.310 ;
        RECT 43.955 129.250 44.245 129.295 ;
        RECT 52.910 129.250 53.230 129.310 ;
        RECT 43.955 129.110 53.230 129.250 ;
        RECT 43.955 129.065 44.245 129.110 ;
        RECT 52.910 129.050 53.230 129.110 ;
        RECT 53.615 129.250 53.905 129.295 ;
        RECT 57.510 129.250 57.830 129.310 ;
        RECT 63.965 129.250 64.255 129.295 ;
        RECT 53.615 129.110 57.830 129.250 ;
        RECT 53.615 129.065 53.905 129.110 ;
        RECT 57.510 129.050 57.830 129.110 ;
        RECT 59.440 129.110 64.255 129.250 ;
        RECT 36.350 128.910 36.670 128.970 ;
        RECT 49.230 128.955 49.550 128.970 ;
        RECT 38.205 128.910 38.495 128.955 ;
        RECT 36.350 128.770 38.495 128.910 ;
        RECT 36.350 128.710 36.670 128.770 ;
        RECT 38.205 128.725 38.495 128.770 ;
        RECT 45.960 128.910 46.250 128.955 ;
        RECT 49.220 128.910 49.550 128.955 ;
        RECT 45.960 128.770 49.550 128.910 ;
        RECT 45.960 128.725 46.250 128.770 ;
        RECT 49.220 128.725 49.550 128.770 ;
        RECT 49.230 128.710 49.550 128.725 ;
        RECT 50.140 128.910 50.430 128.955 ;
        RECT 52.000 128.910 52.290 128.955 ;
        RECT 50.140 128.770 52.290 128.910 ;
        RECT 50.140 128.725 50.430 128.770 ;
        RECT 52.000 128.725 52.290 128.770 ;
        RECT 55.620 128.910 55.910 128.955 ;
        RECT 58.880 128.910 59.170 128.955 ;
        RECT 59.440 128.910 59.580 129.110 ;
        RECT 63.965 129.065 64.255 129.110 ;
        RECT 66.710 129.250 67.030 129.310 ;
        RECT 67.415 129.250 67.705 129.295 ;
        RECT 66.710 129.110 67.705 129.250 ;
        RECT 66.710 129.050 67.030 129.110 ;
        RECT 67.415 129.065 67.705 129.110 ;
        RECT 96.610 129.250 96.930 129.310 ;
        RECT 101.455 129.250 101.745 129.295 ;
        RECT 96.610 129.110 101.745 129.250 ;
        RECT 96.610 129.050 96.930 129.110 ;
        RECT 101.455 129.065 101.745 129.110 ;
        RECT 105.810 129.250 106.130 129.310 ;
        RECT 108.585 129.250 108.875 129.295 ;
        RECT 105.810 129.110 108.875 129.250 ;
        RECT 105.810 129.050 106.130 129.110 ;
        RECT 108.585 129.065 108.875 129.110 ;
        RECT 113.170 129.050 113.490 129.310 ;
        RECT 55.620 128.770 59.580 128.910 ;
        RECT 59.800 128.910 60.090 128.955 ;
        RECT 61.660 128.910 61.950 128.955 ;
        RECT 59.800 128.770 61.950 128.910 ;
        RECT 55.620 128.725 55.910 128.770 ;
        RECT 58.880 128.725 59.170 128.770 ;
        RECT 59.800 128.725 60.090 128.770 ;
        RECT 61.660 128.725 61.950 128.770 ;
        RECT 69.420 128.910 69.710 128.955 ;
        RECT 70.850 128.910 71.170 128.970 ;
        RECT 72.680 128.910 72.970 128.955 ;
        RECT 69.420 128.770 72.970 128.910 ;
        RECT 69.420 128.725 69.710 128.770 ;
        RECT 29.925 128.570 30.215 128.615 ;
        RECT 30.370 128.570 30.690 128.630 ;
        RECT 29.925 128.430 30.690 128.570 ;
        RECT 29.925 128.385 30.215 128.430 ;
        RECT 30.370 128.370 30.690 128.430 ;
        RECT 33.605 128.570 33.895 128.615 ;
        RECT 35.905 128.570 36.195 128.615 ;
        RECT 39.125 128.570 39.415 128.615 ;
        RECT 42.330 128.570 42.650 128.630 ;
        RECT 33.605 128.430 42.650 128.570 ;
        RECT 33.605 128.385 33.895 128.430 ;
        RECT 35.905 128.385 36.195 128.430 ;
        RECT 39.125 128.385 39.415 128.430 ;
        RECT 42.330 128.370 42.650 128.430 ;
        RECT 43.265 128.570 43.555 128.615 ;
        RECT 43.710 128.570 44.030 128.630 ;
        RECT 43.265 128.430 44.030 128.570 ;
        RECT 43.265 128.385 43.555 128.430 ;
        RECT 43.710 128.370 44.030 128.430 ;
        RECT 47.820 128.570 48.110 128.615 ;
        RECT 50.140 128.570 50.355 128.725 ;
        RECT 47.820 128.430 50.355 128.570 ;
        RECT 47.820 128.385 48.110 128.430 ;
        RECT 51.070 128.370 51.390 128.630 ;
        RECT 57.480 128.570 57.770 128.615 ;
        RECT 59.800 128.570 60.015 128.725 ;
        RECT 70.850 128.710 71.170 128.770 ;
        RECT 72.680 128.725 72.970 128.770 ;
        RECT 73.600 128.910 73.890 128.955 ;
        RECT 75.460 128.910 75.750 128.955 ;
        RECT 73.600 128.770 75.750 128.910 ;
        RECT 73.600 128.725 73.890 128.770 ;
        RECT 75.460 128.725 75.750 128.770 ;
        RECT 57.480 128.430 60.015 128.570 ;
        RECT 57.480 128.385 57.770 128.430 ;
        RECT 60.730 128.370 61.050 128.630 ;
        RECT 62.585 128.570 62.875 128.615 ;
        RECT 63.950 128.570 64.270 128.630 ;
        RECT 62.585 128.430 64.270 128.570 ;
        RECT 62.585 128.385 62.875 128.430 ;
        RECT 29.005 128.045 29.295 128.275 ;
        RECT 29.450 128.230 29.770 128.290 ;
        RECT 32.685 128.230 32.975 128.275 ;
        RECT 29.450 128.090 32.975 128.230 ;
        RECT 29.080 127.890 29.220 128.045 ;
        RECT 29.450 128.030 29.770 128.090 ;
        RECT 32.685 128.045 32.975 128.090 ;
        RECT 34.050 128.230 34.370 128.290 ;
        RECT 34.985 128.230 35.275 128.275 ;
        RECT 34.050 128.090 35.275 128.230 ;
        RECT 34.050 128.030 34.370 128.090 ;
        RECT 34.985 128.045 35.275 128.090 ;
        RECT 40.045 128.045 40.335 128.275 ;
        RECT 41.425 128.230 41.715 128.275 ;
        RECT 42.790 128.230 43.110 128.290 ;
        RECT 41.425 128.090 43.110 128.230 ;
        RECT 41.425 128.045 41.715 128.090 ;
        RECT 29.910 127.890 30.230 127.950 ;
        RECT 29.080 127.750 30.230 127.890 ;
        RECT 29.910 127.690 30.230 127.750 ;
        RECT 30.370 127.890 30.690 127.950 ;
        RECT 40.120 127.890 40.260 128.045 ;
        RECT 42.790 128.030 43.110 128.090 ;
        RECT 49.230 128.230 49.550 128.290 ;
        RECT 52.925 128.230 53.215 128.275 ;
        RECT 57.970 128.230 58.290 128.290 ;
        RECT 62.660 128.230 62.800 128.385 ;
        RECT 63.950 128.370 64.270 128.430 ;
        RECT 64.425 128.570 64.715 128.615 ;
        RECT 70.390 128.570 70.710 128.630 ;
        RECT 64.425 128.430 70.710 128.570 ;
        RECT 64.425 128.385 64.715 128.430 ;
        RECT 70.390 128.370 70.710 128.430 ;
        RECT 71.280 128.570 71.570 128.615 ;
        RECT 73.600 128.570 73.815 128.725 ;
        RECT 79.590 128.710 79.910 128.970 ;
        RECT 96.150 128.955 96.470 128.970 ;
        RECT 93.410 128.910 93.700 128.955 ;
        RECT 95.270 128.910 95.560 128.955 ;
        RECT 93.410 128.770 95.560 128.910 ;
        RECT 93.410 128.725 93.700 128.770 ;
        RECT 95.270 128.725 95.560 128.770 ;
        RECT 71.280 128.430 73.815 128.570 ;
        RECT 71.280 128.385 71.570 128.430 ;
        RECT 94.310 128.370 94.630 128.630 ;
        RECT 95.345 128.570 95.560 128.725 ;
        RECT 96.150 128.910 96.480 128.955 ;
        RECT 99.450 128.910 99.740 128.955 ;
        RECT 96.150 128.770 99.740 128.910 ;
        RECT 96.150 128.725 96.480 128.770 ;
        RECT 99.450 128.725 99.740 128.770 ;
        RECT 112.710 128.910 113.030 128.970 ;
        RECT 115.715 128.910 116.005 128.955 ;
        RECT 112.710 128.770 116.005 128.910 ;
        RECT 96.150 128.710 96.470 128.725 ;
        RECT 112.710 128.710 113.030 128.770 ;
        RECT 115.715 128.725 116.005 128.770 ;
        RECT 117.720 128.910 118.010 128.955 ;
        RECT 118.690 128.910 119.010 128.970 ;
        RECT 120.980 128.910 121.270 128.955 ;
        RECT 117.720 128.770 121.270 128.910 ;
        RECT 117.720 128.725 118.010 128.770 ;
        RECT 118.690 128.710 119.010 128.770 ;
        RECT 120.980 128.725 121.270 128.770 ;
        RECT 121.900 128.910 122.190 128.955 ;
        RECT 123.760 128.910 124.050 128.955 ;
        RECT 121.900 128.770 124.050 128.910 ;
        RECT 121.900 128.725 122.190 128.770 ;
        RECT 123.760 128.725 124.050 128.770 ;
        RECT 97.590 128.570 97.880 128.615 ;
        RECT 95.345 128.430 97.880 128.570 ;
        RECT 97.590 128.385 97.880 128.430 ;
        RECT 98.910 128.570 99.230 128.630 ;
        RECT 102.145 128.570 102.435 128.615 ;
        RECT 98.910 128.430 102.435 128.570 ;
        RECT 98.910 128.370 99.230 128.430 ;
        RECT 102.145 128.385 102.435 128.430 ;
        RECT 112.250 128.370 112.570 128.630 ;
        RECT 119.580 128.570 119.870 128.615 ;
        RECT 121.900 128.570 122.115 128.725 ;
        RECT 119.580 128.430 122.115 128.570 ;
        RECT 119.580 128.385 119.870 128.430 ;
        RECT 122.830 128.370 123.150 128.630 ;
        RECT 124.210 128.570 124.530 128.630 ;
        RECT 124.685 128.570 124.975 128.615 ;
        RECT 124.210 128.430 124.975 128.570 ;
        RECT 124.210 128.370 124.530 128.430 ;
        RECT 124.685 128.385 124.975 128.430 ;
        RECT 49.230 128.090 62.800 128.230 ;
        RECT 73.610 128.230 73.930 128.290 ;
        RECT 74.545 128.230 74.835 128.275 ;
        RECT 73.610 128.090 74.835 128.230 ;
        RECT 49.230 128.030 49.550 128.090 ;
        RECT 52.925 128.045 53.215 128.090 ;
        RECT 57.970 128.030 58.290 128.090 ;
        RECT 73.610 128.030 73.930 128.090 ;
        RECT 74.545 128.045 74.835 128.090 ;
        RECT 75.450 128.230 75.770 128.290 ;
        RECT 76.385 128.230 76.675 128.275 ;
        RECT 75.450 128.090 76.675 128.230 ;
        RECT 75.450 128.030 75.770 128.090 ;
        RECT 76.385 128.045 76.675 128.090 ;
        RECT 92.485 128.045 92.775 128.275 ;
        RECT 109.030 128.230 109.350 128.290 ;
        RECT 111.345 128.230 111.635 128.275 ;
        RECT 109.030 128.090 111.635 128.230 ;
        RECT 30.370 127.750 40.260 127.890 ;
        RECT 47.820 127.890 48.110 127.935 ;
        RECT 50.600 127.890 50.890 127.935 ;
        RECT 52.460 127.890 52.750 127.935 ;
        RECT 47.820 127.750 52.750 127.890 ;
        RECT 30.370 127.690 30.690 127.750 ;
        RECT 47.820 127.705 48.110 127.750 ;
        RECT 50.600 127.705 50.890 127.750 ;
        RECT 52.460 127.705 52.750 127.750 ;
        RECT 57.480 127.890 57.770 127.935 ;
        RECT 60.260 127.890 60.550 127.935 ;
        RECT 62.120 127.890 62.410 127.935 ;
        RECT 57.480 127.750 62.410 127.890 ;
        RECT 57.480 127.705 57.770 127.750 ;
        RECT 60.260 127.705 60.550 127.750 ;
        RECT 62.120 127.705 62.410 127.750 ;
        RECT 71.280 127.890 71.570 127.935 ;
        RECT 74.060 127.890 74.350 127.935 ;
        RECT 75.920 127.890 76.210 127.935 ;
        RECT 71.280 127.750 76.210 127.890 ;
        RECT 76.460 127.890 76.600 128.045 ;
        RECT 86.045 127.890 86.335 127.935 ;
        RECT 87.870 127.890 88.190 127.950 ;
        RECT 92.560 127.890 92.700 128.045 ;
        RECT 109.030 128.030 109.350 128.090 ;
        RECT 111.345 128.045 111.635 128.090 ;
        RECT 76.460 127.750 92.700 127.890 ;
        RECT 92.950 127.890 93.240 127.935 ;
        RECT 94.810 127.890 95.100 127.935 ;
        RECT 97.590 127.890 97.880 127.935 ;
        RECT 92.950 127.750 97.880 127.890 ;
        RECT 71.280 127.705 71.570 127.750 ;
        RECT 74.060 127.705 74.350 127.750 ;
        RECT 75.920 127.705 76.210 127.750 ;
        RECT 86.045 127.705 86.335 127.750 ;
        RECT 87.870 127.690 88.190 127.750 ;
        RECT 92.950 127.705 93.240 127.750 ;
        RECT 94.810 127.705 95.100 127.750 ;
        RECT 97.590 127.705 97.880 127.750 ;
        RECT 119.580 127.890 119.870 127.935 ;
        RECT 122.360 127.890 122.650 127.935 ;
        RECT 124.220 127.890 124.510 127.935 ;
        RECT 119.580 127.750 124.510 127.890 ;
        RECT 119.580 127.705 119.870 127.750 ;
        RECT 122.360 127.705 122.650 127.750 ;
        RECT 124.220 127.705 124.510 127.750 ;
        RECT 31.290 127.550 31.610 127.610 ;
        RECT 31.765 127.550 32.055 127.595 ;
        RECT 31.290 127.410 32.055 127.550 ;
        RECT 31.290 127.350 31.610 127.410 ;
        RECT 31.765 127.365 32.055 127.410 ;
        RECT 20.640 126.730 127.820 127.210 ;
        RECT 29.910 126.530 30.230 126.590 ;
        RECT 32.915 126.530 33.205 126.575 ;
        RECT 42.790 126.530 43.110 126.590 ;
        RECT 29.910 126.390 31.060 126.530 ;
        RECT 29.910 126.330 30.230 126.390 ;
        RECT 26.690 125.850 27.010 125.910 ;
        RECT 24.940 125.710 27.010 125.850 ;
        RECT 24.940 125.555 25.080 125.710 ;
        RECT 26.690 125.650 27.010 125.710 ;
        RECT 28.990 125.850 29.310 125.910 ;
        RECT 30.920 125.895 31.060 126.390 ;
        RECT 32.915 126.390 43.110 126.530 ;
        RECT 32.915 126.345 33.205 126.390 ;
        RECT 42.790 126.330 43.110 126.390 ;
        RECT 73.610 126.330 73.930 126.590 ;
        RECT 78.915 126.530 79.205 126.575 ;
        RECT 80.510 126.530 80.830 126.590 ;
        RECT 113.630 126.530 113.950 126.590 ;
        RECT 117.770 126.530 118.090 126.590 ;
        RECT 78.915 126.390 80.830 126.530 ;
        RECT 78.915 126.345 79.205 126.390 ;
        RECT 80.510 126.330 80.830 126.390 ;
        RECT 111.880 126.390 118.090 126.530 ;
        RECT 36.780 126.190 37.070 126.235 ;
        RECT 39.560 126.190 39.850 126.235 ;
        RECT 41.420 126.190 41.710 126.235 ;
        RECT 36.780 126.050 41.710 126.190 ;
        RECT 36.780 126.005 37.070 126.050 ;
        RECT 39.560 126.005 39.850 126.050 ;
        RECT 41.420 126.005 41.710 126.050 ;
        RECT 82.780 126.190 83.070 126.235 ;
        RECT 85.560 126.190 85.850 126.235 ;
        RECT 87.420 126.190 87.710 126.235 ;
        RECT 82.780 126.050 87.710 126.190 ;
        RECT 82.780 126.005 83.070 126.050 ;
        RECT 85.560 126.005 85.850 126.050 ;
        RECT 87.420 126.005 87.710 126.050 ;
        RECT 98.540 126.050 107.420 126.190 ;
        RECT 29.925 125.850 30.215 125.895 ;
        RECT 28.990 125.710 30.215 125.850 ;
        RECT 28.990 125.650 29.310 125.710 ;
        RECT 29.925 125.665 30.215 125.710 ;
        RECT 30.845 125.850 31.135 125.895 ;
        RECT 33.590 125.850 33.910 125.910 ;
        RECT 43.725 125.850 44.015 125.895 ;
        RECT 51.530 125.850 51.850 125.910 ;
        RECT 30.845 125.710 51.850 125.850 ;
        RECT 30.845 125.665 31.135 125.710 ;
        RECT 33.590 125.650 33.910 125.710 ;
        RECT 43.725 125.665 44.015 125.710 ;
        RECT 51.530 125.650 51.850 125.710 ;
        RECT 62.125 125.850 62.415 125.895 ;
        RECT 63.950 125.850 64.270 125.910 ;
        RECT 67.185 125.850 67.475 125.895 ;
        RECT 62.125 125.710 67.475 125.850 ;
        RECT 62.125 125.665 62.415 125.710 ;
        RECT 63.950 125.650 64.270 125.710 ;
        RECT 67.185 125.665 67.475 125.710 ;
        RECT 70.390 125.850 70.710 125.910 ;
        RECT 84.650 125.850 84.970 125.910 ;
        RECT 70.390 125.710 72.000 125.850 ;
        RECT 70.390 125.650 70.710 125.710 ;
        RECT 23.945 125.510 24.235 125.555 ;
        RECT 24.865 125.510 25.155 125.555 ;
        RECT 23.945 125.370 25.155 125.510 ;
        RECT 23.945 125.325 24.235 125.370 ;
        RECT 24.865 125.325 25.155 125.370 ;
        RECT 26.245 125.510 26.535 125.555 ;
        RECT 36.780 125.510 37.070 125.555 ;
        RECT 26.245 125.370 27.840 125.510 ;
        RECT 26.245 125.325 26.535 125.370 ;
        RECT 23.470 124.630 23.790 124.890 ;
        RECT 25.310 124.630 25.630 124.890 ;
        RECT 27.150 124.630 27.470 124.890 ;
        RECT 27.700 124.875 27.840 125.370 ;
        RECT 36.780 125.370 39.315 125.510 ;
        RECT 36.780 125.325 37.070 125.370 ;
        RECT 34.920 125.170 35.210 125.215 ;
        RECT 36.350 125.170 36.670 125.230 ;
        RECT 39.100 125.215 39.315 125.370 ;
        RECT 40.030 125.310 40.350 125.570 ;
        RECT 41.885 125.325 42.175 125.555 ;
        RECT 42.790 125.510 43.110 125.570 ;
        RECT 44.185 125.510 44.475 125.555 ;
        RECT 42.790 125.370 44.475 125.510 ;
        RECT 38.180 125.170 38.470 125.215 ;
        RECT 34.920 125.030 38.470 125.170 ;
        RECT 34.920 124.985 35.210 125.030 ;
        RECT 36.350 124.970 36.670 125.030 ;
        RECT 38.180 124.985 38.470 125.030 ;
        RECT 39.100 125.170 39.390 125.215 ;
        RECT 40.960 125.170 41.250 125.215 ;
        RECT 39.100 125.030 41.250 125.170 ;
        RECT 39.100 124.985 39.390 125.030 ;
        RECT 40.960 124.985 41.250 125.030 ;
        RECT 27.625 124.645 27.915 124.875 ;
        RECT 29.450 124.630 29.770 124.890 ;
        RECT 35.890 124.830 36.210 124.890 ;
        RECT 41.960 124.830 42.100 125.325 ;
        RECT 42.790 125.310 43.110 125.370 ;
        RECT 44.185 125.325 44.475 125.370 ;
        RECT 57.510 125.510 57.830 125.570 ;
        RECT 63.045 125.510 63.335 125.555 ;
        RECT 57.510 125.370 63.335 125.510 ;
        RECT 57.510 125.310 57.830 125.370 ;
        RECT 63.045 125.325 63.335 125.370 ;
        RECT 70.850 125.510 71.170 125.570 ;
        RECT 71.860 125.555 72.000 125.710 ;
        RECT 84.650 125.710 87.180 125.850 ;
        RECT 84.650 125.650 84.970 125.710 ;
        RECT 71.325 125.510 71.615 125.555 ;
        RECT 70.850 125.370 71.615 125.510 ;
        RECT 70.850 125.310 71.170 125.370 ;
        RECT 71.325 125.325 71.615 125.370 ;
        RECT 71.785 125.510 72.075 125.555 ;
        RECT 72.230 125.510 72.550 125.570 ;
        RECT 71.785 125.370 72.550 125.510 ;
        RECT 71.785 125.325 72.075 125.370 ;
        RECT 72.230 125.310 72.550 125.370 ;
        RECT 72.690 125.310 73.010 125.570 ;
        RECT 74.530 125.310 74.850 125.570 ;
        RECT 76.370 125.510 76.690 125.570 ;
        RECT 77.305 125.510 77.595 125.555 ;
        RECT 76.370 125.370 77.595 125.510 ;
        RECT 76.370 125.310 76.690 125.370 ;
        RECT 77.305 125.325 77.595 125.370 ;
        RECT 82.780 125.510 83.070 125.555 ;
        RECT 86.045 125.510 86.335 125.555 ;
        RECT 86.490 125.510 86.810 125.570 ;
        RECT 82.780 125.370 85.315 125.510 ;
        RECT 82.780 125.325 83.070 125.370 ;
        RECT 85.100 125.215 85.315 125.370 ;
        RECT 86.045 125.370 86.810 125.510 ;
        RECT 87.040 125.510 87.180 125.710 ;
        RECT 87.870 125.650 88.190 125.910 ;
        RECT 93.865 125.850 94.155 125.895 ;
        RECT 95.690 125.850 96.010 125.910 ;
        RECT 98.540 125.895 98.680 126.050 ;
        RECT 107.280 125.895 107.420 126.050 ;
        RECT 111.880 125.895 112.020 126.390 ;
        RECT 113.630 126.330 113.950 126.390 ;
        RECT 117.770 126.330 118.090 126.390 ;
        RECT 112.710 126.190 113.030 126.250 ;
        RECT 112.340 126.050 113.030 126.190 ;
        RECT 112.340 125.895 112.480 126.050 ;
        RECT 112.710 125.990 113.030 126.050 ;
        RECT 119.120 126.190 119.410 126.235 ;
        RECT 121.900 126.190 122.190 126.235 ;
        RECT 123.760 126.190 124.050 126.235 ;
        RECT 119.120 126.050 124.050 126.190 ;
        RECT 119.120 126.005 119.410 126.050 ;
        RECT 121.900 126.005 122.190 126.050 ;
        RECT 123.760 126.005 124.050 126.050 ;
        RECT 124.685 126.005 124.975 126.235 ;
        RECT 98.465 125.850 98.755 125.895 ;
        RECT 107.205 125.850 107.495 125.895 ;
        RECT 111.805 125.850 112.095 125.895 ;
        RECT 93.865 125.710 98.755 125.850 ;
        RECT 93.865 125.665 94.155 125.710 ;
        RECT 95.690 125.650 96.010 125.710 ;
        RECT 98.465 125.665 98.755 125.710 ;
        RECT 101.760 125.710 105.120 125.850 ;
        RECT 87.040 125.370 87.640 125.510 ;
        RECT 86.045 125.325 86.335 125.370 ;
        RECT 86.490 125.310 86.810 125.370 ;
        RECT 52.005 125.170 52.295 125.215 ;
        RECT 44.720 125.030 52.295 125.170 ;
        RECT 44.720 124.890 44.860 125.030 ;
        RECT 52.005 124.985 52.295 125.030 ;
        RECT 62.585 125.170 62.875 125.215 ;
        RECT 80.920 125.170 81.210 125.215 ;
        RECT 84.180 125.170 84.470 125.215 ;
        RECT 85.100 125.170 85.390 125.215 ;
        RECT 86.960 125.170 87.250 125.215 ;
        RECT 62.585 125.030 68.780 125.170 ;
        RECT 62.585 124.985 62.875 125.030 ;
        RECT 68.640 124.890 68.780 125.030 ;
        RECT 80.920 125.030 84.880 125.170 ;
        RECT 80.920 124.985 81.210 125.030 ;
        RECT 84.180 124.985 84.470 125.030 ;
        RECT 35.890 124.690 42.100 124.830 ;
        RECT 35.890 124.630 36.210 124.690 ;
        RECT 44.630 124.630 44.950 124.890 ;
        RECT 46.010 124.830 46.330 124.890 ;
        RECT 46.485 124.830 46.775 124.875 ;
        RECT 46.010 124.690 46.775 124.830 ;
        RECT 46.010 124.630 46.330 124.690 ;
        RECT 46.485 124.645 46.775 124.690 ;
        RECT 52.450 124.630 52.770 124.890 ;
        RECT 54.290 124.630 54.610 124.890 ;
        RECT 64.870 124.630 65.190 124.890 ;
        RECT 67.170 124.830 67.490 124.890 ;
        RECT 68.105 124.830 68.395 124.875 ;
        RECT 67.170 124.690 68.395 124.830 ;
        RECT 67.170 124.630 67.490 124.690 ;
        RECT 68.105 124.645 68.395 124.690 ;
        RECT 68.550 124.630 68.870 124.890 ;
        RECT 70.405 124.830 70.695 124.875 ;
        RECT 71.310 124.830 71.630 124.890 ;
        RECT 70.405 124.690 71.630 124.830 ;
        RECT 70.405 124.645 70.695 124.690 ;
        RECT 71.310 124.630 71.630 124.690 ;
        RECT 75.465 124.830 75.755 124.875 ;
        RECT 76.370 124.830 76.690 124.890 ;
        RECT 75.465 124.690 76.690 124.830 ;
        RECT 75.465 124.645 75.755 124.690 ;
        RECT 76.370 124.630 76.690 124.690 ;
        RECT 77.765 124.830 78.055 124.875 ;
        RECT 79.590 124.830 79.910 124.890 ;
        RECT 77.765 124.690 79.910 124.830 ;
        RECT 84.740 124.830 84.880 125.030 ;
        RECT 85.100 125.030 87.250 125.170 ;
        RECT 87.500 125.170 87.640 125.370 ;
        RECT 89.250 125.310 89.570 125.570 ;
        RECT 98.925 125.510 99.215 125.555 ;
        RECT 101.760 125.510 101.900 125.710 ;
        RECT 98.925 125.370 101.900 125.510 ;
        RECT 98.925 125.325 99.215 125.370 ;
        RECT 102.130 125.310 102.450 125.570 ;
        RECT 103.050 125.310 103.370 125.570 ;
        RECT 103.525 125.325 103.815 125.555 ;
        RECT 104.445 125.325 104.735 125.555 ;
        RECT 104.980 125.510 105.120 125.710 ;
        RECT 107.205 125.710 112.095 125.850 ;
        RECT 107.205 125.665 107.495 125.710 ;
        RECT 111.805 125.665 112.095 125.710 ;
        RECT 112.265 125.665 112.555 125.895 ;
        RECT 124.760 125.850 124.900 126.005 ;
        RECT 123.840 125.710 124.900 125.850 ;
        RECT 106.270 125.510 106.590 125.570 ;
        RECT 108.125 125.510 108.415 125.555 ;
        RECT 109.490 125.510 109.810 125.570 ;
        RECT 104.980 125.370 109.810 125.510 ;
        RECT 92.485 125.170 92.775 125.215 ;
        RECT 103.600 125.170 103.740 125.325 ;
        RECT 87.500 125.030 92.775 125.170 ;
        RECT 85.100 124.985 85.390 125.030 ;
        RECT 86.960 124.985 87.250 125.030 ;
        RECT 92.485 124.985 92.775 125.030 ;
        RECT 99.460 125.030 103.740 125.170 ;
        RECT 104.520 125.170 104.660 125.325 ;
        RECT 106.270 125.310 106.590 125.370 ;
        RECT 108.125 125.325 108.415 125.370 ;
        RECT 109.490 125.310 109.810 125.370 ;
        RECT 110.410 125.510 110.730 125.570 ;
        RECT 112.725 125.510 113.015 125.555 ;
        RECT 115.255 125.510 115.545 125.555 ;
        RECT 116.390 125.510 116.710 125.570 ;
        RECT 110.410 125.370 116.710 125.510 ;
        RECT 110.410 125.310 110.730 125.370 ;
        RECT 112.725 125.325 113.015 125.370 ;
        RECT 115.255 125.325 115.545 125.370 ;
        RECT 116.390 125.310 116.710 125.370 ;
        RECT 119.120 125.510 119.410 125.555 ;
        RECT 122.385 125.510 122.675 125.555 ;
        RECT 123.840 125.510 123.980 125.710 ;
        RECT 119.120 125.370 121.655 125.510 ;
        RECT 119.120 125.325 119.410 125.370 ;
        RECT 113.630 125.170 113.950 125.230 ;
        RECT 104.520 125.030 113.950 125.170 ;
        RECT 86.030 124.830 86.350 124.890 ;
        RECT 84.740 124.690 86.350 124.830 ;
        RECT 77.765 124.645 78.055 124.690 ;
        RECT 79.590 124.630 79.910 124.690 ;
        RECT 86.030 124.630 86.350 124.690 ;
        RECT 89.710 124.630 90.030 124.890 ;
        RECT 90.630 124.630 90.950 124.890 ;
        RECT 92.930 124.830 93.250 124.890 ;
        RECT 99.460 124.875 99.600 125.030 ;
        RECT 113.630 124.970 113.950 125.030 ;
        RECT 117.260 125.170 117.550 125.215 ;
        RECT 119.610 125.170 119.930 125.230 ;
        RECT 121.440 125.215 121.655 125.370 ;
        RECT 122.385 125.370 123.980 125.510 ;
        RECT 122.385 125.325 122.675 125.370 ;
        RECT 124.210 125.310 124.530 125.570 ;
        RECT 125.605 125.325 125.895 125.555 ;
        RECT 120.520 125.170 120.810 125.215 ;
        RECT 117.260 125.030 120.810 125.170 ;
        RECT 117.260 124.985 117.550 125.030 ;
        RECT 119.610 124.970 119.930 125.030 ;
        RECT 120.520 124.985 120.810 125.030 ;
        RECT 121.440 125.170 121.730 125.215 ;
        RECT 123.300 125.170 123.590 125.215 ;
        RECT 125.680 125.170 125.820 125.325 ;
        RECT 121.440 125.030 123.590 125.170 ;
        RECT 121.440 124.985 121.730 125.030 ;
        RECT 123.300 124.985 123.590 125.030 ;
        RECT 123.840 125.030 125.820 125.170 ;
        RECT 99.385 124.830 99.675 124.875 ;
        RECT 92.930 124.690 99.675 124.830 ;
        RECT 92.930 124.630 93.250 124.690 ;
        RECT 99.385 124.645 99.675 124.690 ;
        RECT 101.210 124.630 101.530 124.890 ;
        RECT 104.890 124.630 105.210 124.890 ;
        RECT 107.665 124.830 107.955 124.875 ;
        RECT 109.030 124.830 109.350 124.890 ;
        RECT 107.665 124.690 109.350 124.830 ;
        RECT 107.665 124.645 107.955 124.690 ;
        RECT 109.030 124.630 109.350 124.690 ;
        RECT 109.965 124.830 110.255 124.875 ;
        RECT 112.250 124.830 112.570 124.890 ;
        RECT 109.965 124.690 112.570 124.830 ;
        RECT 109.965 124.645 110.255 124.690 ;
        RECT 112.250 124.630 112.570 124.690 ;
        RECT 114.565 124.830 114.855 124.875 ;
        RECT 123.840 124.830 123.980 125.030 ;
        RECT 114.565 124.690 123.980 124.830 ;
        RECT 114.565 124.645 114.855 124.690 ;
        RECT 20.640 124.010 127.820 124.490 ;
        RECT 22.795 123.810 23.085 123.855 ;
        RECT 29.450 123.810 29.770 123.870 ;
        RECT 22.795 123.670 29.770 123.810 ;
        RECT 22.795 123.625 23.085 123.670 ;
        RECT 29.450 123.610 29.770 123.670 ;
        RECT 30.370 123.810 30.690 123.870 ;
        RECT 34.525 123.810 34.815 123.855 ;
        RECT 30.370 123.670 34.815 123.810 ;
        RECT 30.370 123.610 30.690 123.670 ;
        RECT 34.525 123.625 34.815 123.670 ;
        RECT 36.825 123.625 37.115 123.855 ;
        RECT 38.665 123.625 38.955 123.855 ;
        RECT 49.015 123.810 49.305 123.855 ;
        RECT 52.450 123.810 52.770 123.870 ;
        RECT 49.015 123.670 52.770 123.810 ;
        RECT 49.015 123.625 49.305 123.670 ;
        RECT 23.470 123.470 23.790 123.530 ;
        RECT 24.800 123.470 25.090 123.515 ;
        RECT 28.060 123.470 28.350 123.515 ;
        RECT 23.470 123.330 28.350 123.470 ;
        RECT 23.470 123.270 23.790 123.330 ;
        RECT 24.800 123.285 25.090 123.330 ;
        RECT 28.060 123.285 28.350 123.330 ;
        RECT 28.980 123.470 29.270 123.515 ;
        RECT 30.840 123.470 31.130 123.515 ;
        RECT 28.980 123.330 31.130 123.470 ;
        RECT 28.980 123.285 29.270 123.330 ;
        RECT 30.840 123.285 31.130 123.330 ;
        RECT 34.985 123.470 35.275 123.515 ;
        RECT 34.985 123.330 36.580 123.470 ;
        RECT 34.985 123.285 35.275 123.330 ;
        RECT 26.660 123.130 26.950 123.175 ;
        RECT 28.980 123.130 29.195 123.285 ;
        RECT 26.660 122.990 29.195 123.130 ;
        RECT 31.765 123.130 32.055 123.175 ;
        RECT 34.510 123.130 34.830 123.190 ;
        RECT 35.890 123.130 36.210 123.190 ;
        RECT 31.765 122.990 36.210 123.130 ;
        RECT 26.660 122.945 26.950 122.990 ;
        RECT 31.765 122.945 32.055 122.990 ;
        RECT 34.510 122.930 34.830 122.990 ;
        RECT 35.890 122.930 36.210 122.990 ;
        RECT 27.150 122.790 27.470 122.850 ;
        RECT 29.925 122.790 30.215 122.835 ;
        RECT 27.150 122.650 30.215 122.790 ;
        RECT 27.150 122.590 27.470 122.650 ;
        RECT 29.925 122.605 30.215 122.650 ;
        RECT 33.590 122.590 33.910 122.850 ;
        RECT 36.440 122.790 36.580 123.330 ;
        RECT 36.900 123.130 37.040 123.625 ;
        RECT 38.740 123.470 38.880 123.625 ;
        RECT 52.450 123.610 52.770 123.670 ;
        RECT 66.035 123.810 66.325 123.855 ;
        RECT 67.170 123.810 67.490 123.870 ;
        RECT 66.035 123.670 67.490 123.810 ;
        RECT 66.035 123.625 66.325 123.670 ;
        RECT 67.170 123.610 67.490 123.670 ;
        RECT 75.910 123.810 76.230 123.870 ;
        RECT 83.730 123.810 84.050 123.870 ;
        RECT 84.895 123.810 85.185 123.855 ;
        RECT 75.910 123.670 83.500 123.810 ;
        RECT 75.910 123.610 76.230 123.670 ;
        RECT 40.030 123.470 40.350 123.530 ;
        RECT 38.740 123.330 40.350 123.470 ;
        RECT 40.030 123.270 40.350 123.330 ;
        RECT 41.360 123.470 41.650 123.515 ;
        RECT 42.790 123.470 43.110 123.530 ;
        RECT 44.620 123.470 44.910 123.515 ;
        RECT 41.360 123.330 44.910 123.470 ;
        RECT 41.360 123.285 41.650 123.330 ;
        RECT 42.790 123.270 43.110 123.330 ;
        RECT 44.620 123.285 44.910 123.330 ;
        RECT 45.540 123.470 45.830 123.515 ;
        RECT 47.400 123.470 47.690 123.515 ;
        RECT 45.540 123.330 47.690 123.470 ;
        RECT 45.540 123.285 45.830 123.330 ;
        RECT 47.400 123.285 47.690 123.330 ;
        RECT 51.020 123.470 51.310 123.515 ;
        RECT 53.370 123.470 53.690 123.530 ;
        RECT 54.280 123.470 54.570 123.515 ;
        RECT 51.020 123.330 54.570 123.470 ;
        RECT 51.020 123.285 51.310 123.330 ;
        RECT 37.745 123.130 38.035 123.175 ;
        RECT 36.900 122.990 38.035 123.130 ;
        RECT 37.745 122.945 38.035 122.990 ;
        RECT 43.220 123.130 43.510 123.175 ;
        RECT 45.540 123.130 45.755 123.285 ;
        RECT 53.370 123.270 53.690 123.330 ;
        RECT 54.280 123.285 54.570 123.330 ;
        RECT 55.200 123.470 55.490 123.515 ;
        RECT 57.060 123.470 57.350 123.515 ;
        RECT 55.200 123.330 57.350 123.470 ;
        RECT 55.200 123.285 55.490 123.330 ;
        RECT 57.060 123.285 57.350 123.330 ;
        RECT 68.040 123.470 68.330 123.515 ;
        RECT 69.470 123.470 69.790 123.530 ;
        RECT 79.590 123.515 79.910 123.530 ;
        RECT 71.300 123.470 71.590 123.515 ;
        RECT 68.040 123.330 71.590 123.470 ;
        RECT 68.040 123.285 68.330 123.330 ;
        RECT 43.220 122.990 45.755 123.130 ;
        RECT 48.325 123.130 48.615 123.175 ;
        RECT 49.230 123.130 49.550 123.190 ;
        RECT 48.325 122.990 49.550 123.130 ;
        RECT 43.220 122.945 43.510 122.990 ;
        RECT 48.325 122.945 48.615 122.990 ;
        RECT 49.230 122.930 49.550 122.990 ;
        RECT 52.880 123.130 53.170 123.175 ;
        RECT 55.200 123.130 55.415 123.285 ;
        RECT 69.470 123.270 69.790 123.330 ;
        RECT 71.300 123.285 71.590 123.330 ;
        RECT 72.220 123.470 72.510 123.515 ;
        RECT 74.080 123.470 74.370 123.515 ;
        RECT 72.220 123.330 74.370 123.470 ;
        RECT 72.220 123.285 72.510 123.330 ;
        RECT 74.080 123.285 74.370 123.330 ;
        RECT 76.850 123.470 77.140 123.515 ;
        RECT 78.710 123.470 79.000 123.515 ;
        RECT 76.850 123.330 79.000 123.470 ;
        RECT 76.850 123.285 77.140 123.330 ;
        RECT 78.710 123.285 79.000 123.330 ;
        RECT 52.880 122.990 55.415 123.130 ;
        RECT 52.880 122.945 53.170 122.990 ;
        RECT 57.970 122.930 58.290 123.190 ;
        RECT 61.665 122.945 61.955 123.175 ;
        RECT 64.870 123.130 65.190 123.190 ;
        RECT 65.345 123.130 65.635 123.175 ;
        RECT 64.870 122.990 65.635 123.130 ;
        RECT 42.330 122.790 42.650 122.850 ;
        RECT 36.440 122.650 42.650 122.790 ;
        RECT 42.330 122.590 42.650 122.650 ;
        RECT 46.470 122.590 46.790 122.850 ;
        RECT 56.130 122.590 56.450 122.850 ;
        RECT 58.890 122.790 59.210 122.850 ;
        RECT 61.740 122.790 61.880 122.945 ;
        RECT 64.870 122.930 65.190 122.990 ;
        RECT 65.345 122.945 65.635 122.990 ;
        RECT 69.900 123.130 70.190 123.175 ;
        RECT 72.220 123.130 72.435 123.285 ;
        RECT 69.900 122.990 72.435 123.130 ;
        RECT 75.005 123.130 75.295 123.175 ;
        RECT 75.450 123.130 75.770 123.190 ;
        RECT 75.925 123.130 76.215 123.175 ;
        RECT 75.005 122.990 76.215 123.130 ;
        RECT 69.900 122.945 70.190 122.990 ;
        RECT 75.005 122.945 75.295 122.990 ;
        RECT 75.450 122.930 75.770 122.990 ;
        RECT 75.925 122.945 76.215 122.990 ;
        RECT 76.370 123.130 76.690 123.190 ;
        RECT 77.765 123.130 78.055 123.175 ;
        RECT 76.370 122.990 78.055 123.130 ;
        RECT 78.785 123.130 79.000 123.285 ;
        RECT 79.590 123.470 79.920 123.515 ;
        RECT 82.890 123.470 83.180 123.515 ;
        RECT 79.590 123.330 83.180 123.470 ;
        RECT 79.590 123.285 79.920 123.330 ;
        RECT 82.890 123.285 83.180 123.330 ;
        RECT 79.590 123.270 79.910 123.285 ;
        RECT 81.030 123.130 81.320 123.175 ;
        RECT 78.785 122.990 81.320 123.130 ;
        RECT 83.360 123.130 83.500 123.670 ;
        RECT 83.730 123.670 85.185 123.810 ;
        RECT 83.730 123.610 84.050 123.670 ;
        RECT 84.895 123.625 85.185 123.670 ;
        RECT 86.030 123.610 86.350 123.870 ;
        RECT 86.490 123.810 86.810 123.870 ;
        RECT 86.965 123.810 87.255 123.855 ;
        RECT 86.490 123.670 87.255 123.810 ;
        RECT 86.490 123.610 86.810 123.670 ;
        RECT 86.965 123.625 87.255 123.670 ;
        RECT 92.255 123.810 92.545 123.855 ;
        RECT 92.930 123.810 93.250 123.870 ;
        RECT 105.810 123.810 106.130 123.870 ;
        RECT 116.390 123.810 116.710 123.870 ;
        RECT 117.325 123.810 117.615 123.855 ;
        RECT 92.255 123.670 93.250 123.810 ;
        RECT 92.255 123.625 92.545 123.670 ;
        RECT 92.930 123.610 93.250 123.670 ;
        RECT 103.600 123.670 110.640 123.810 ;
        RECT 89.710 123.470 90.030 123.530 ;
        RECT 94.260 123.470 94.550 123.515 ;
        RECT 97.520 123.470 97.810 123.515 ;
        RECT 86.580 123.330 88.560 123.470 ;
        RECT 86.580 123.175 86.720 123.330 ;
        RECT 86.505 123.130 86.795 123.175 ;
        RECT 83.360 122.990 86.795 123.130 ;
        RECT 76.370 122.930 76.690 122.990 ;
        RECT 77.765 122.945 78.055 122.990 ;
        RECT 81.030 122.945 81.320 122.990 ;
        RECT 86.505 122.945 86.795 122.990 ;
        RECT 87.885 122.945 88.175 123.175 ;
        RECT 88.420 123.130 88.560 123.330 ;
        RECT 89.710 123.330 97.810 123.470 ;
        RECT 89.710 123.270 90.030 123.330 ;
        RECT 94.260 123.285 94.550 123.330 ;
        RECT 97.520 123.285 97.810 123.330 ;
        RECT 98.440 123.470 98.730 123.515 ;
        RECT 100.300 123.470 100.590 123.515 ;
        RECT 98.440 123.330 100.590 123.470 ;
        RECT 98.440 123.285 98.730 123.330 ;
        RECT 100.300 123.285 100.590 123.330 ;
        RECT 89.250 123.130 89.570 123.190 ;
        RECT 88.420 122.990 89.570 123.130 ;
        RECT 70.390 122.790 70.710 122.850 ;
        RECT 58.890 122.650 70.710 122.790 ;
        RECT 58.890 122.590 59.210 122.650 ;
        RECT 70.390 122.590 70.710 122.650 ;
        RECT 73.150 122.590 73.470 122.850 ;
        RECT 85.570 122.790 85.890 122.850 ;
        RECT 87.960 122.790 88.100 122.945 ;
        RECT 89.250 122.930 89.570 122.990 ;
        RECT 90.630 122.930 90.950 123.190 ;
        RECT 96.120 123.130 96.410 123.175 ;
        RECT 98.440 123.130 98.655 123.285 ;
        RECT 96.120 122.990 98.655 123.130 ;
        RECT 101.225 123.130 101.515 123.175 ;
        RECT 103.600 123.130 103.740 123.670 ;
        RECT 105.810 123.610 106.130 123.670 ;
        RECT 103.920 123.470 104.210 123.515 ;
        RECT 104.890 123.470 105.210 123.530 ;
        RECT 107.180 123.470 107.470 123.515 ;
        RECT 103.920 123.330 107.470 123.470 ;
        RECT 103.920 123.285 104.210 123.330 ;
        RECT 104.890 123.270 105.210 123.330 ;
        RECT 107.180 123.285 107.470 123.330 ;
        RECT 108.100 123.470 108.390 123.515 ;
        RECT 109.960 123.470 110.250 123.515 ;
        RECT 108.100 123.330 110.250 123.470 ;
        RECT 108.100 123.285 108.390 123.330 ;
        RECT 109.960 123.285 110.250 123.330 ;
        RECT 101.225 122.990 103.740 123.130 ;
        RECT 105.780 123.130 106.070 123.175 ;
        RECT 108.100 123.130 108.315 123.285 ;
        RECT 105.780 122.990 108.315 123.130 ;
        RECT 110.500 123.130 110.640 123.670 ;
        RECT 116.390 123.670 117.615 123.810 ;
        RECT 116.390 123.610 116.710 123.670 ;
        RECT 117.325 123.625 117.615 123.670 ;
        RECT 119.610 123.610 119.930 123.870 ;
        RECT 116.480 123.330 119.380 123.470 ;
        RECT 116.480 123.190 116.620 123.330 ;
        RECT 110.870 123.130 111.190 123.190 ;
        RECT 110.500 122.990 111.190 123.130 ;
        RECT 96.120 122.945 96.410 122.990 ;
        RECT 101.225 122.945 101.515 122.990 ;
        RECT 105.780 122.945 106.070 122.990 ;
        RECT 110.870 122.930 111.190 122.990 ;
        RECT 112.250 122.930 112.570 123.190 ;
        RECT 113.630 123.130 113.950 123.190 ;
        RECT 116.390 123.130 116.710 123.190 ;
        RECT 119.240 123.175 119.380 123.330 ;
        RECT 113.630 122.990 116.710 123.130 ;
        RECT 113.630 122.930 113.950 122.990 ;
        RECT 116.390 122.930 116.710 122.990 ;
        RECT 116.865 122.945 117.155 123.175 ;
        RECT 119.165 122.945 119.455 123.175 ;
        RECT 85.570 122.650 88.100 122.790 ;
        RECT 85.570 122.590 85.890 122.650 ;
        RECT 99.370 122.590 99.690 122.850 ;
        RECT 101.915 122.790 102.205 122.835 ;
        RECT 106.270 122.790 106.590 122.850 ;
        RECT 101.915 122.650 106.590 122.790 ;
        RECT 101.915 122.605 102.205 122.650 ;
        RECT 106.270 122.590 106.590 122.650 ;
        RECT 109.045 122.790 109.335 122.835 ;
        RECT 116.940 122.790 117.080 122.945 ;
        RECT 109.045 122.650 111.560 122.790 ;
        RECT 109.045 122.605 109.335 122.650 ;
        RECT 111.420 122.495 111.560 122.650 ;
        RECT 112.800 122.650 117.080 122.790 ;
        RECT 26.660 122.450 26.950 122.495 ;
        RECT 29.440 122.450 29.730 122.495 ;
        RECT 31.300 122.450 31.590 122.495 ;
        RECT 26.660 122.310 31.590 122.450 ;
        RECT 26.660 122.265 26.950 122.310 ;
        RECT 29.440 122.265 29.730 122.310 ;
        RECT 31.300 122.265 31.590 122.310 ;
        RECT 43.220 122.450 43.510 122.495 ;
        RECT 46.000 122.450 46.290 122.495 ;
        RECT 47.860 122.450 48.150 122.495 ;
        RECT 43.220 122.310 48.150 122.450 ;
        RECT 43.220 122.265 43.510 122.310 ;
        RECT 46.000 122.265 46.290 122.310 ;
        RECT 47.860 122.265 48.150 122.310 ;
        RECT 52.880 122.450 53.170 122.495 ;
        RECT 55.660 122.450 55.950 122.495 ;
        RECT 57.520 122.450 57.810 122.495 ;
        RECT 52.880 122.310 57.810 122.450 ;
        RECT 52.880 122.265 53.170 122.310 ;
        RECT 55.660 122.265 55.950 122.310 ;
        RECT 57.520 122.265 57.810 122.310 ;
        RECT 69.900 122.450 70.190 122.495 ;
        RECT 72.680 122.450 72.970 122.495 ;
        RECT 74.540 122.450 74.830 122.495 ;
        RECT 69.900 122.310 74.830 122.450 ;
        RECT 69.900 122.265 70.190 122.310 ;
        RECT 72.680 122.265 72.970 122.310 ;
        RECT 74.540 122.265 74.830 122.310 ;
        RECT 76.390 122.450 76.680 122.495 ;
        RECT 78.250 122.450 78.540 122.495 ;
        RECT 81.030 122.450 81.320 122.495 ;
        RECT 76.390 122.310 81.320 122.450 ;
        RECT 76.390 122.265 76.680 122.310 ;
        RECT 78.250 122.265 78.540 122.310 ;
        RECT 81.030 122.265 81.320 122.310 ;
        RECT 96.120 122.450 96.410 122.495 ;
        RECT 98.900 122.450 99.190 122.495 ;
        RECT 100.760 122.450 101.050 122.495 ;
        RECT 96.120 122.310 101.050 122.450 ;
        RECT 96.120 122.265 96.410 122.310 ;
        RECT 98.900 122.265 99.190 122.310 ;
        RECT 100.760 122.265 101.050 122.310 ;
        RECT 105.780 122.450 106.070 122.495 ;
        RECT 108.560 122.450 108.850 122.495 ;
        RECT 110.420 122.450 110.710 122.495 ;
        RECT 105.780 122.310 110.710 122.450 ;
        RECT 105.780 122.265 106.070 122.310 ;
        RECT 108.560 122.265 108.850 122.310 ;
        RECT 110.420 122.265 110.710 122.310 ;
        RECT 111.345 122.265 111.635 122.495 ;
        RECT 34.050 122.110 34.370 122.170 ;
        RECT 39.355 122.110 39.645 122.155 ;
        RECT 44.630 122.110 44.950 122.170 ;
        RECT 34.050 121.970 44.950 122.110 ;
        RECT 34.050 121.910 34.370 121.970 ;
        RECT 39.355 121.925 39.645 121.970 ;
        RECT 44.630 121.910 44.950 121.970 ;
        RECT 62.125 122.110 62.415 122.155 ;
        RECT 63.950 122.110 64.270 122.170 ;
        RECT 62.125 121.970 64.270 122.110 ;
        RECT 62.125 121.925 62.415 121.970 ;
        RECT 63.950 121.910 64.270 121.970 ;
        RECT 64.410 121.910 64.730 122.170 ;
        RECT 89.710 121.910 90.030 122.170 ;
        RECT 91.565 122.110 91.855 122.155 ;
        RECT 93.850 122.110 94.170 122.170 ;
        RECT 91.565 121.970 94.170 122.110 ;
        RECT 91.565 121.925 91.855 121.970 ;
        RECT 93.850 121.910 94.170 121.970 ;
        RECT 109.030 122.110 109.350 122.170 ;
        RECT 112.800 122.110 112.940 122.650 ;
        RECT 117.770 122.590 118.090 122.850 ;
        RECT 109.030 121.970 112.940 122.110 ;
        RECT 113.185 122.110 113.475 122.155 ;
        RECT 113.630 122.110 113.950 122.170 ;
        RECT 113.185 121.970 113.950 122.110 ;
        RECT 109.030 121.910 109.350 121.970 ;
        RECT 113.185 121.925 113.475 121.970 ;
        RECT 113.630 121.910 113.950 121.970 ;
        RECT 115.010 121.910 115.330 122.170 ;
        RECT 20.640 121.290 127.820 121.770 ;
        RECT 25.095 121.090 25.385 121.135 ;
        RECT 30.370 121.090 30.690 121.150 ;
        RECT 25.095 120.950 30.690 121.090 ;
        RECT 25.095 120.905 25.385 120.950 ;
        RECT 30.370 120.890 30.690 120.950 ;
        RECT 36.350 120.890 36.670 121.150 ;
        RECT 42.790 121.090 43.110 121.150 ;
        RECT 43.265 121.090 43.555 121.135 ;
        RECT 42.790 120.950 43.555 121.090 ;
        RECT 42.790 120.890 43.110 120.950 ;
        RECT 43.265 120.905 43.555 120.950 ;
        RECT 46.470 121.090 46.790 121.150 ;
        RECT 46.945 121.090 47.235 121.135 ;
        RECT 46.470 120.950 47.235 121.090 ;
        RECT 46.470 120.890 46.790 120.950 ;
        RECT 46.945 120.905 47.235 120.950 ;
        RECT 52.925 121.090 53.215 121.135 ;
        RECT 53.370 121.090 53.690 121.150 ;
        RECT 52.925 120.950 53.690 121.090 ;
        RECT 52.925 120.905 53.215 120.950 ;
        RECT 53.370 120.890 53.690 120.950 ;
        RECT 55.685 121.090 55.975 121.135 ;
        RECT 56.130 121.090 56.450 121.150 ;
        RECT 55.685 120.950 56.450 121.090 ;
        RECT 55.685 120.905 55.975 120.950 ;
        RECT 56.130 120.890 56.450 120.950 ;
        RECT 68.550 121.135 68.870 121.150 ;
        RECT 68.550 120.905 69.085 121.135 ;
        RECT 69.470 121.090 69.790 121.150 ;
        RECT 69.945 121.090 70.235 121.135 ;
        RECT 69.470 120.950 70.235 121.090 ;
        RECT 68.550 120.890 68.870 120.905 ;
        RECT 69.470 120.890 69.790 120.950 ;
        RECT 69.945 120.905 70.235 120.950 ;
        RECT 72.245 121.090 72.535 121.135 ;
        RECT 73.150 121.090 73.470 121.150 ;
        RECT 72.245 120.950 73.470 121.090 ;
        RECT 72.245 120.905 72.535 120.950 ;
        RECT 73.150 120.890 73.470 120.950 ;
        RECT 85.570 120.890 85.890 121.150 ;
        RECT 99.370 121.090 99.690 121.150 ;
        RECT 100.305 121.090 100.595 121.135 ;
        RECT 99.370 120.950 100.595 121.090 ;
        RECT 99.370 120.890 99.690 120.950 ;
        RECT 100.305 120.905 100.595 120.950 ;
        RECT 108.355 121.090 108.645 121.135 ;
        RECT 109.030 121.090 109.350 121.150 ;
        RECT 108.355 120.950 109.350 121.090 ;
        RECT 108.355 120.905 108.645 120.950 ;
        RECT 109.030 120.890 109.350 120.950 ;
        RECT 28.960 120.750 29.250 120.795 ;
        RECT 31.740 120.750 32.030 120.795 ;
        RECT 33.600 120.750 33.890 120.795 ;
        RECT 28.960 120.610 33.890 120.750 ;
        RECT 28.960 120.565 29.250 120.610 ;
        RECT 31.740 120.565 32.030 120.610 ;
        RECT 33.600 120.565 33.890 120.610 ;
        RECT 60.290 120.750 60.580 120.795 ;
        RECT 62.150 120.750 62.440 120.795 ;
        RECT 64.930 120.750 65.220 120.795 ;
        RECT 60.290 120.610 65.220 120.750 ;
        RECT 60.290 120.565 60.580 120.610 ;
        RECT 62.150 120.565 62.440 120.610 ;
        RECT 64.930 120.565 65.220 120.610 ;
        RECT 90.140 120.750 90.430 120.795 ;
        RECT 92.920 120.750 93.210 120.795 ;
        RECT 94.780 120.750 95.070 120.795 ;
        RECT 90.140 120.610 95.070 120.750 ;
        RECT 90.140 120.565 90.430 120.610 ;
        RECT 92.920 120.565 93.210 120.610 ;
        RECT 94.780 120.565 95.070 120.610 ;
        RECT 112.220 120.750 112.510 120.795 ;
        RECT 115.000 120.750 115.290 120.795 ;
        RECT 116.860 120.750 117.150 120.795 ;
        RECT 112.220 120.610 117.150 120.750 ;
        RECT 112.220 120.565 112.510 120.610 ;
        RECT 115.000 120.565 115.290 120.610 ;
        RECT 116.860 120.565 117.150 120.610 ;
        RECT 34.065 120.410 34.355 120.455 ;
        RECT 34.510 120.410 34.830 120.470 ;
        RECT 51.990 120.410 52.310 120.470 ;
        RECT 57.525 120.410 57.815 120.455 ;
        RECT 34.065 120.270 34.830 120.410 ;
        RECT 34.065 120.225 34.355 120.270 ;
        RECT 34.510 120.210 34.830 120.270 ;
        RECT 43.800 120.270 57.815 120.410 ;
        RECT 28.960 120.070 29.250 120.115 ;
        RECT 28.960 119.930 31.495 120.070 ;
        RECT 28.960 119.885 29.250 119.930 ;
        RECT 25.310 119.730 25.630 119.790 ;
        RECT 31.280 119.775 31.495 119.930 ;
        RECT 32.210 119.870 32.530 120.130 ;
        RECT 43.800 120.115 43.940 120.270 ;
        RECT 51.990 120.210 52.310 120.270 ;
        RECT 35.905 120.070 36.195 120.115 ;
        RECT 43.725 120.070 44.015 120.115 ;
        RECT 35.905 119.930 44.015 120.070 ;
        RECT 35.905 119.885 36.195 119.930 ;
        RECT 43.725 119.885 44.015 119.930 ;
        RECT 46.010 119.870 46.330 120.130 ;
        RECT 53.460 120.115 53.600 120.270 ;
        RECT 57.525 120.225 57.815 120.270 ;
        RECT 57.970 120.410 58.290 120.470 ;
        RECT 59.825 120.410 60.115 120.455 ;
        RECT 61.665 120.410 61.955 120.455 ;
        RECT 64.410 120.410 64.730 120.470 ;
        RECT 57.970 120.270 60.500 120.410 ;
        RECT 57.970 120.210 58.290 120.270 ;
        RECT 59.825 120.225 60.115 120.270 ;
        RECT 60.360 120.130 60.500 120.270 ;
        RECT 61.665 120.270 64.730 120.410 ;
        RECT 61.665 120.225 61.955 120.270 ;
        RECT 64.410 120.210 64.730 120.270 ;
        RECT 82.810 120.210 83.130 120.470 ;
        RECT 83.285 120.410 83.575 120.455 ;
        RECT 84.650 120.410 84.970 120.470 ;
        RECT 86.275 120.410 86.565 120.455 ;
        RECT 83.285 120.270 86.565 120.410 ;
        RECT 83.285 120.225 83.575 120.270 ;
        RECT 84.650 120.210 84.970 120.270 ;
        RECT 86.275 120.225 86.565 120.270 ;
        RECT 87.870 120.410 88.190 120.470 ;
        RECT 93.405 120.410 93.695 120.455 ;
        RECT 93.850 120.410 94.170 120.470 ;
        RECT 87.870 120.270 93.160 120.410 ;
        RECT 87.870 120.210 88.190 120.270 ;
        RECT 53.385 119.885 53.675 120.115 ;
        RECT 54.290 120.070 54.610 120.130 ;
        RECT 54.765 120.070 55.055 120.115 ;
        RECT 54.290 119.930 55.055 120.070 ;
        RECT 54.290 119.870 54.610 119.930 ;
        RECT 54.765 119.885 55.055 119.930 ;
        RECT 58.890 119.870 59.210 120.130 ;
        RECT 60.270 119.870 60.590 120.130 ;
        RECT 64.930 120.070 65.220 120.115 ;
        RECT 62.685 119.930 65.220 120.070 ;
        RECT 62.685 119.775 62.900 119.930 ;
        RECT 64.930 119.885 65.220 119.930 ;
        RECT 70.390 119.870 70.710 120.130 ;
        RECT 71.310 119.870 71.630 120.130 ;
        RECT 80.510 120.070 80.830 120.130 ;
        RECT 83.745 120.070 84.035 120.115 ;
        RECT 80.510 119.930 84.035 120.070 ;
        RECT 80.510 119.870 80.830 119.930 ;
        RECT 83.745 119.885 84.035 119.930 ;
        RECT 90.140 120.070 90.430 120.115 ;
        RECT 93.020 120.070 93.160 120.270 ;
        RECT 93.405 120.270 94.170 120.410 ;
        RECT 93.405 120.225 93.695 120.270 ;
        RECT 93.850 120.210 94.170 120.270 ;
        RECT 110.870 120.410 111.190 120.470 ;
        RECT 110.870 120.270 115.240 120.410 ;
        RECT 110.870 120.210 111.190 120.270 ;
        RECT 95.245 120.070 95.535 120.115 ;
        RECT 90.140 119.930 92.675 120.070 ;
        RECT 93.020 119.930 95.535 120.070 ;
        RECT 90.140 119.885 90.430 119.930 ;
        RECT 27.100 119.730 27.390 119.775 ;
        RECT 30.360 119.730 30.650 119.775 ;
        RECT 25.310 119.590 30.650 119.730 ;
        RECT 25.310 119.530 25.630 119.590 ;
        RECT 27.100 119.545 27.390 119.590 ;
        RECT 30.360 119.545 30.650 119.590 ;
        RECT 31.280 119.730 31.570 119.775 ;
        RECT 33.140 119.730 33.430 119.775 ;
        RECT 31.280 119.590 33.430 119.730 ;
        RECT 31.280 119.545 31.570 119.590 ;
        RECT 33.140 119.545 33.430 119.590 ;
        RECT 60.750 119.730 61.040 119.775 ;
        RECT 62.610 119.730 62.900 119.775 ;
        RECT 60.750 119.590 62.900 119.730 ;
        RECT 60.750 119.545 61.040 119.590 ;
        RECT 62.610 119.545 62.900 119.590 ;
        RECT 63.490 119.775 63.810 119.790 ;
        RECT 63.490 119.730 63.820 119.775 ;
        RECT 66.790 119.730 67.080 119.775 ;
        RECT 63.490 119.590 67.080 119.730 ;
        RECT 63.490 119.545 63.820 119.590 ;
        RECT 66.790 119.545 67.080 119.590 ;
        RECT 88.280 119.730 88.570 119.775 ;
        RECT 89.710 119.730 90.030 119.790 ;
        RECT 92.460 119.775 92.675 119.930 ;
        RECT 95.245 119.885 95.535 119.930 ;
        RECT 101.210 119.870 101.530 120.130 ;
        RECT 112.220 120.070 112.510 120.115 ;
        RECT 115.100 120.070 115.240 120.270 ;
        RECT 115.470 120.210 115.790 120.470 ;
        RECT 117.325 120.070 117.615 120.115 ;
        RECT 124.210 120.070 124.530 120.130 ;
        RECT 112.220 119.930 114.755 120.070 ;
        RECT 115.100 119.930 124.530 120.070 ;
        RECT 112.220 119.885 112.510 119.930 ;
        RECT 113.630 119.775 113.950 119.790 ;
        RECT 91.540 119.730 91.830 119.775 ;
        RECT 88.280 119.590 91.830 119.730 ;
        RECT 88.280 119.545 88.570 119.590 ;
        RECT 63.490 119.530 63.810 119.545 ;
        RECT 89.710 119.530 90.030 119.590 ;
        RECT 91.540 119.545 91.830 119.590 ;
        RECT 92.460 119.730 92.750 119.775 ;
        RECT 94.320 119.730 94.610 119.775 ;
        RECT 92.460 119.590 94.610 119.730 ;
        RECT 92.460 119.545 92.750 119.590 ;
        RECT 94.320 119.545 94.610 119.590 ;
        RECT 110.360 119.730 110.650 119.775 ;
        RECT 113.620 119.730 113.950 119.775 ;
        RECT 110.360 119.590 113.950 119.730 ;
        RECT 110.360 119.545 110.650 119.590 ;
        RECT 113.620 119.545 113.950 119.590 ;
        RECT 114.540 119.775 114.755 119.930 ;
        RECT 117.325 119.885 117.615 119.930 ;
        RECT 124.210 119.870 124.530 119.930 ;
        RECT 114.540 119.730 114.830 119.775 ;
        RECT 116.400 119.730 116.690 119.775 ;
        RECT 114.540 119.590 116.690 119.730 ;
        RECT 114.540 119.545 114.830 119.590 ;
        RECT 116.400 119.545 116.690 119.590 ;
        RECT 113.630 119.530 113.950 119.545 ;
        RECT 20.640 118.570 127.820 119.050 ;
        RECT 32.210 118.170 32.530 118.430 ;
        RECT 115.470 118.370 115.790 118.430 ;
        RECT 115.945 118.370 116.235 118.415 ;
        RECT 115.470 118.230 116.235 118.370 ;
        RECT 115.470 118.170 115.790 118.230 ;
        RECT 115.945 118.185 116.235 118.230 ;
        RECT 120.070 118.030 120.390 118.090 ;
        RECT 120.070 117.890 123.520 118.030 ;
        RECT 120.070 117.830 120.390 117.890 ;
        RECT 31.290 117.490 31.610 117.750 ;
        RECT 115.010 117.490 115.330 117.750 ;
        RECT 116.850 117.690 117.170 117.750 ;
        RECT 123.380 117.735 123.520 117.890 ;
        RECT 119.625 117.690 119.915 117.735 ;
        RECT 116.850 117.550 119.915 117.690 ;
        RECT 116.850 117.490 117.170 117.550 ;
        RECT 119.625 117.505 119.915 117.550 ;
        RECT 121.005 117.505 121.295 117.735 ;
        RECT 123.305 117.505 123.595 117.735 ;
        RECT 115.930 117.350 116.250 117.410 ;
        RECT 121.080 117.350 121.220 117.505 ;
        RECT 115.930 117.210 121.220 117.350 ;
        RECT 115.930 117.150 116.250 117.210 ;
        RECT 121.925 117.010 122.215 117.055 ;
        RECT 124.670 117.010 124.990 117.070 ;
        RECT 121.925 116.870 124.990 117.010 ;
        RECT 121.925 116.825 122.215 116.870 ;
        RECT 124.670 116.810 124.990 116.870 ;
        RECT 119.610 116.670 119.930 116.730 ;
        RECT 120.085 116.670 120.375 116.715 ;
        RECT 119.610 116.530 120.375 116.670 ;
        RECT 119.610 116.470 119.930 116.530 ;
        RECT 120.085 116.485 120.375 116.530 ;
        RECT 121.450 116.670 121.770 116.730 ;
        RECT 122.385 116.670 122.675 116.715 ;
        RECT 121.450 116.530 122.675 116.670 ;
        RECT 121.450 116.470 121.770 116.530 ;
        RECT 122.385 116.485 122.675 116.530 ;
        RECT 20.640 115.850 127.820 116.330 ;
        RECT 70.390 115.650 70.710 115.710 ;
        RECT 81.430 115.650 81.750 115.710 ;
        RECT 70.390 115.510 77.520 115.650 ;
        RECT 70.390 115.450 70.710 115.510 ;
        RECT 29.565 115.310 29.855 115.355 ;
        RECT 32.685 115.310 32.975 115.355 ;
        RECT 34.575 115.310 34.865 115.355 ;
        RECT 29.565 115.170 34.865 115.310 ;
        RECT 29.565 115.125 29.855 115.170 ;
        RECT 32.685 115.125 32.975 115.170 ;
        RECT 34.575 115.125 34.865 115.170 ;
        RECT 37.285 115.125 37.575 115.355 ;
        RECT 54.750 115.310 55.070 115.370 ;
        RECT 77.380 115.310 77.520 115.510 ;
        RECT 81.430 115.510 95.000 115.650 ;
        RECT 81.430 115.450 81.750 115.510 ;
        RECT 54.750 115.170 71.080 115.310 ;
        RECT 77.380 115.170 83.500 115.310 ;
        RECT 34.065 114.970 34.355 115.015 ;
        RECT 37.360 114.970 37.500 115.125 ;
        RECT 54.750 115.110 55.070 115.170 ;
        RECT 34.065 114.830 37.500 114.970 ;
        RECT 50.610 114.970 50.930 115.030 ;
        RECT 64.870 114.970 65.190 115.030 ;
        RECT 50.610 114.830 65.190 114.970 ;
        RECT 34.065 114.785 34.355 114.830 ;
        RECT 50.610 114.770 50.930 114.830 ;
        RECT 64.870 114.770 65.190 114.830 ;
        RECT 25.770 114.290 26.090 114.350 ;
        RECT 28.485 114.335 28.775 114.650 ;
        RECT 29.565 114.630 29.855 114.675 ;
        RECT 33.145 114.630 33.435 114.675 ;
        RECT 34.980 114.630 35.270 114.675 ;
        RECT 29.565 114.490 35.270 114.630 ;
        RECT 29.565 114.445 29.855 114.490 ;
        RECT 33.145 114.445 33.435 114.490 ;
        RECT 34.980 114.445 35.270 114.490 ;
        RECT 35.430 114.430 35.750 114.690 ;
        RECT 35.890 114.630 36.210 114.690 ;
        RECT 36.825 114.630 37.115 114.675 ;
        RECT 35.890 114.490 37.115 114.630 ;
        RECT 35.890 114.430 36.210 114.490 ;
        RECT 36.825 114.445 37.115 114.490 ;
        RECT 38.190 114.430 38.510 114.690 ;
        RECT 39.585 114.445 39.875 114.675 ;
        RECT 43.250 114.630 43.570 114.690 ;
        RECT 45.565 114.630 45.855 114.675 ;
        RECT 43.250 114.490 45.855 114.630 ;
        RECT 28.185 114.290 28.775 114.335 ;
        RECT 31.425 114.290 32.075 114.335 ;
        RECT 39.660 114.290 39.800 114.445 ;
        RECT 43.250 114.430 43.570 114.490 ;
        RECT 45.565 114.445 45.855 114.490 ;
        RECT 49.245 114.445 49.535 114.675 ;
        RECT 50.150 114.630 50.470 114.690 ;
        RECT 53.845 114.630 54.135 114.675 ;
        RECT 50.150 114.490 54.135 114.630 ;
        RECT 40.030 114.290 40.350 114.350 ;
        RECT 49.320 114.290 49.460 114.445 ;
        RECT 50.150 114.430 50.470 114.490 ;
        RECT 53.845 114.445 54.135 114.490 ;
        RECT 62.585 114.630 62.875 114.675 ;
        RECT 70.390 114.630 70.710 114.690 ;
        RECT 70.940 114.675 71.080 115.170 ;
        RECT 74.990 114.970 75.310 115.030 ;
        RECT 79.145 114.970 79.435 115.015 ;
        RECT 74.990 114.830 79.435 114.970 ;
        RECT 74.990 114.770 75.310 114.830 ;
        RECT 79.145 114.785 79.435 114.830 ;
        RECT 62.585 114.490 70.710 114.630 ;
        RECT 62.585 114.445 62.875 114.490 ;
        RECT 70.390 114.430 70.710 114.490 ;
        RECT 70.865 114.445 71.155 114.675 ;
        RECT 79.590 114.430 79.910 114.690 ;
        RECT 80.065 114.445 80.355 114.675 ;
        RECT 80.510 114.630 80.830 114.690 ;
        RECT 83.360 114.675 83.500 115.170 ;
        RECT 81.445 114.630 81.735 114.675 ;
        RECT 80.510 114.490 81.735 114.630 ;
        RECT 57.510 114.290 57.830 114.350 ;
        RECT 63.965 114.290 64.255 114.335 ;
        RECT 25.770 114.150 32.075 114.290 ;
        RECT 25.770 114.090 26.090 114.150 ;
        RECT 28.185 114.105 28.475 114.150 ;
        RECT 31.425 114.105 32.075 114.150 ;
        RECT 35.520 114.150 64.255 114.290 ;
        RECT 26.705 113.950 26.995 113.995 ;
        RECT 27.150 113.950 27.470 114.010 ;
        RECT 26.705 113.810 27.470 113.950 ;
        RECT 26.705 113.765 26.995 113.810 ;
        RECT 27.150 113.750 27.470 113.810 ;
        RECT 27.610 113.950 27.930 114.010 ;
        RECT 35.520 113.950 35.660 114.150 ;
        RECT 40.030 114.090 40.350 114.150 ;
        RECT 57.510 114.090 57.830 114.150 ;
        RECT 63.965 114.105 64.255 114.150 ;
        RECT 79.130 114.290 79.450 114.350 ;
        RECT 80.140 114.290 80.280 114.445 ;
        RECT 80.510 114.430 80.830 114.490 ;
        RECT 81.445 114.445 81.735 114.490 ;
        RECT 83.285 114.445 83.575 114.675 ;
        RECT 86.030 114.430 86.350 114.690 ;
        RECT 94.860 114.675 95.000 115.510 ;
        RECT 105.350 115.310 105.670 115.370 ;
        RECT 107.665 115.310 107.955 115.355 ;
        RECT 109.490 115.310 109.810 115.370 ;
        RECT 105.350 115.170 106.960 115.310 ;
        RECT 105.350 115.110 105.670 115.170 ;
        RECT 106.820 114.675 106.960 115.170 ;
        RECT 107.665 115.170 109.810 115.310 ;
        RECT 107.665 115.125 107.955 115.170 ;
        RECT 109.490 115.110 109.810 115.170 ;
        RECT 118.195 115.310 118.485 115.355 ;
        RECT 120.085 115.310 120.375 115.355 ;
        RECT 123.205 115.310 123.495 115.355 ;
        RECT 118.195 115.170 123.495 115.310 ;
        RECT 118.195 115.125 118.485 115.170 ;
        RECT 120.085 115.125 120.375 115.170 ;
        RECT 123.205 115.125 123.495 115.170 ;
        RECT 110.870 114.970 111.190 115.030 ;
        RECT 117.325 114.970 117.615 115.015 ;
        RECT 110.870 114.830 117.615 114.970 ;
        RECT 110.870 114.770 111.190 114.830 ;
        RECT 117.325 114.785 117.615 114.830 ;
        RECT 118.705 114.970 118.995 115.015 ;
        RECT 121.450 114.970 121.770 115.030 ;
        RECT 118.705 114.830 121.770 114.970 ;
        RECT 118.705 114.785 118.995 114.830 ;
        RECT 121.450 114.770 121.770 114.830 ;
        RECT 94.325 114.445 94.615 114.675 ;
        RECT 94.785 114.445 95.075 114.675 ;
        RECT 97.545 114.630 97.835 114.675 ;
        RECT 105.365 114.630 105.655 114.675 ;
        RECT 97.545 114.490 105.655 114.630 ;
        RECT 97.545 114.445 97.835 114.490 ;
        RECT 105.365 114.445 105.655 114.490 ;
        RECT 106.745 114.445 107.035 114.675 ;
        RECT 109.045 114.630 109.335 114.675 ;
        RECT 115.945 114.630 116.235 114.675 ;
        RECT 116.850 114.630 117.170 114.690 ;
        RECT 109.045 114.490 117.170 114.630 ;
        RECT 109.045 114.445 109.335 114.490 ;
        RECT 115.945 114.445 116.235 114.490 ;
        RECT 84.665 114.290 84.955 114.335 ;
        RECT 90.170 114.290 90.490 114.350 ;
        RECT 94.400 114.290 94.540 114.445 ;
        RECT 97.620 114.290 97.760 114.445 ;
        RECT 79.130 114.150 97.760 114.290 ;
        RECT 105.440 114.290 105.580 114.445 ;
        RECT 109.120 114.290 109.260 114.445 ;
        RECT 116.850 114.430 117.170 114.490 ;
        RECT 117.790 114.630 118.080 114.675 ;
        RECT 119.625 114.630 119.915 114.675 ;
        RECT 123.205 114.630 123.495 114.675 ;
        RECT 117.790 114.490 123.495 114.630 ;
        RECT 117.790 114.445 118.080 114.490 ;
        RECT 119.625 114.445 119.915 114.490 ;
        RECT 123.205 114.445 123.495 114.490 ;
        RECT 124.285 114.335 124.575 114.650 ;
        RECT 105.440 114.150 109.260 114.290 ;
        RECT 116.405 114.290 116.695 114.335 ;
        RECT 120.985 114.290 121.635 114.335 ;
        RECT 124.285 114.290 124.875 114.335 ;
        RECT 116.405 114.150 124.875 114.290 ;
        RECT 79.130 114.090 79.450 114.150 ;
        RECT 84.665 114.105 84.955 114.150 ;
        RECT 90.170 114.090 90.490 114.150 ;
        RECT 116.405 114.105 116.695 114.150 ;
        RECT 120.985 114.105 121.635 114.150 ;
        RECT 124.585 114.105 124.875 114.150 ;
        RECT 27.610 113.810 35.660 113.950 ;
        RECT 27.610 113.750 27.930 113.810 ;
        RECT 35.890 113.750 36.210 114.010 ;
        RECT 38.650 113.950 38.970 114.010 ;
        RECT 39.125 113.950 39.415 113.995 ;
        RECT 38.650 113.810 39.415 113.950 ;
        RECT 38.650 113.750 38.970 113.810 ;
        RECT 39.125 113.765 39.415 113.810 ;
        RECT 46.470 113.750 46.790 114.010 ;
        RECT 48.785 113.950 49.075 113.995 ;
        RECT 49.230 113.950 49.550 114.010 ;
        RECT 48.785 113.810 49.550 113.950 ;
        RECT 48.785 113.765 49.075 113.810 ;
        RECT 49.230 113.750 49.550 113.810 ;
        RECT 54.765 113.950 55.055 113.995 ;
        RECT 57.050 113.950 57.370 114.010 ;
        RECT 54.765 113.810 57.370 113.950 ;
        RECT 54.765 113.765 55.055 113.810 ;
        RECT 57.050 113.750 57.370 113.810 ;
        RECT 71.785 113.950 72.075 113.995 ;
        RECT 73.610 113.950 73.930 114.010 ;
        RECT 71.785 113.810 73.930 113.950 ;
        RECT 71.785 113.765 72.075 113.810 ;
        RECT 73.610 113.750 73.930 113.810 ;
        RECT 80.510 113.750 80.830 114.010 ;
        RECT 82.365 113.950 82.655 113.995 ;
        RECT 83.730 113.950 84.050 114.010 ;
        RECT 82.365 113.810 84.050 113.950 ;
        RECT 82.365 113.765 82.655 113.810 ;
        RECT 83.730 113.750 84.050 113.810 ;
        RECT 86.950 113.750 87.270 114.010 ;
        RECT 93.865 113.950 94.155 113.995 ;
        RECT 94.310 113.950 94.630 114.010 ;
        RECT 93.865 113.810 94.630 113.950 ;
        RECT 93.865 113.765 94.155 113.810 ;
        RECT 94.310 113.750 94.630 113.810 ;
        RECT 95.705 113.950 95.995 113.995 ;
        RECT 96.610 113.950 96.930 114.010 ;
        RECT 95.705 113.810 96.930 113.950 ;
        RECT 95.705 113.765 95.995 113.810 ;
        RECT 96.610 113.750 96.930 113.810 ;
        RECT 98.005 113.950 98.295 113.995 ;
        RECT 98.910 113.950 99.230 114.010 ;
        RECT 98.005 113.810 99.230 113.950 ;
        RECT 98.005 113.765 98.295 113.810 ;
        RECT 98.910 113.750 99.230 113.810 ;
        RECT 104.905 113.950 105.195 113.995 ;
        RECT 105.350 113.950 105.670 114.010 ;
        RECT 104.905 113.810 105.670 113.950 ;
        RECT 104.905 113.765 105.195 113.810 ;
        RECT 105.350 113.750 105.670 113.810 ;
        RECT 108.585 113.950 108.875 113.995 ;
        RECT 109.030 113.950 109.350 114.010 ;
        RECT 108.585 113.810 109.350 113.950 ;
        RECT 108.585 113.765 108.875 113.810 ;
        RECT 109.030 113.750 109.350 113.810 ;
        RECT 126.065 113.950 126.355 113.995 ;
        RECT 126.510 113.950 126.830 114.010 ;
        RECT 126.065 113.810 126.830 113.950 ;
        RECT 126.065 113.765 126.355 113.810 ;
        RECT 126.510 113.750 126.830 113.810 ;
        RECT 20.640 113.130 127.820 113.610 ;
        RECT 25.770 112.730 26.090 112.990 ;
        RECT 28.085 112.930 28.375 112.975 ;
        RECT 31.290 112.930 31.610 112.990 ;
        RECT 35.890 112.930 36.210 112.990 ;
        RECT 28.085 112.790 31.610 112.930 ;
        RECT 28.085 112.745 28.375 112.790 ;
        RECT 31.290 112.730 31.610 112.790 ;
        RECT 35.520 112.790 36.210 112.930 ;
        RECT 35.520 112.635 35.660 112.790 ;
        RECT 35.890 112.730 36.210 112.790 ;
        RECT 36.810 112.930 37.130 112.990 ;
        RECT 38.665 112.930 38.955 112.975 ;
        RECT 36.810 112.790 38.955 112.930 ;
        RECT 36.810 112.730 37.130 112.790 ;
        RECT 38.665 112.745 38.955 112.790 ;
        RECT 40.505 112.930 40.795 112.975 ;
        RECT 43.710 112.930 44.030 112.990 ;
        RECT 40.505 112.790 44.030 112.930 ;
        RECT 40.505 112.745 40.795 112.790 ;
        RECT 43.710 112.730 44.030 112.790 ;
        RECT 46.010 112.930 46.330 112.990 ;
        RECT 51.545 112.930 51.835 112.975 ;
        RECT 54.750 112.930 55.070 112.990 ;
        RECT 46.010 112.790 50.840 112.930 ;
        RECT 46.010 112.730 46.330 112.790 ;
        RECT 27.165 112.590 27.455 112.635 ;
        RECT 29.565 112.590 29.855 112.635 ;
        RECT 32.805 112.590 33.455 112.635 ;
        RECT 27.165 112.450 33.455 112.590 ;
        RECT 27.165 112.405 27.455 112.450 ;
        RECT 29.565 112.405 30.155 112.450 ;
        RECT 32.805 112.405 33.455 112.450 ;
        RECT 35.445 112.405 35.735 112.635 ;
        RECT 39.585 112.590 39.875 112.635 ;
        RECT 41.985 112.590 42.275 112.635 ;
        RECT 45.225 112.590 45.875 112.635 ;
        RECT 39.585 112.450 45.875 112.590 ;
        RECT 39.585 112.405 39.875 112.450 ;
        RECT 41.985 112.405 42.575 112.450 ;
        RECT 45.225 112.405 45.875 112.450 ;
        RECT 46.470 112.590 46.790 112.650 ;
        RECT 47.865 112.590 48.155 112.635 ;
        RECT 46.470 112.450 48.155 112.590 ;
        RECT 24.865 112.250 25.155 112.295 ;
        RECT 25.325 112.250 25.615 112.295 ;
        RECT 26.705 112.250 26.995 112.295 ;
        RECT 27.610 112.250 27.930 112.310 ;
        RECT 24.865 112.110 27.930 112.250 ;
        RECT 24.865 112.065 25.155 112.110 ;
        RECT 25.325 112.065 25.615 112.110 ;
        RECT 26.705 112.065 26.995 112.110 ;
        RECT 27.610 112.050 27.930 112.110 ;
        RECT 29.865 112.090 30.155 112.405 ;
        RECT 30.945 112.250 31.235 112.295 ;
        RECT 34.525 112.250 34.815 112.295 ;
        RECT 36.360 112.250 36.650 112.295 ;
        RECT 30.945 112.110 36.650 112.250 ;
        RECT 30.945 112.065 31.235 112.110 ;
        RECT 34.525 112.065 34.815 112.110 ;
        RECT 36.360 112.065 36.650 112.110 ;
        RECT 37.730 112.050 38.050 112.310 ;
        RECT 39.125 112.250 39.415 112.295 ;
        RECT 40.030 112.250 40.350 112.310 ;
        RECT 39.125 112.110 40.350 112.250 ;
        RECT 39.125 112.065 39.415 112.110 ;
        RECT 40.030 112.050 40.350 112.110 ;
        RECT 42.285 112.090 42.575 112.405 ;
        RECT 46.470 112.390 46.790 112.450 ;
        RECT 47.865 112.405 48.155 112.450 ;
        RECT 43.365 112.250 43.655 112.295 ;
        RECT 46.945 112.250 47.235 112.295 ;
        RECT 48.780 112.250 49.070 112.295 ;
        RECT 43.365 112.110 49.070 112.250 ;
        RECT 43.365 112.065 43.655 112.110 ;
        RECT 46.945 112.065 47.235 112.110 ;
        RECT 48.780 112.065 49.070 112.110 ;
        RECT 49.245 112.250 49.535 112.295 ;
        RECT 49.690 112.250 50.010 112.310 ;
        RECT 50.700 112.295 50.840 112.790 ;
        RECT 51.545 112.790 55.070 112.930 ;
        RECT 51.545 112.745 51.835 112.790 ;
        RECT 54.750 112.730 55.070 112.790 ;
        RECT 57.050 112.730 57.370 112.990 ;
        RECT 78.225 112.930 78.515 112.975 ;
        RECT 82.350 112.930 82.670 112.990 ;
        RECT 78.225 112.790 82.670 112.930 ;
        RECT 78.225 112.745 78.515 112.790 ;
        RECT 82.350 112.730 82.670 112.790 ;
        RECT 87.425 112.745 87.715 112.975 ;
        RECT 90.645 112.930 90.935 112.975 ;
        RECT 93.850 112.930 94.170 112.990 ;
        RECT 90.645 112.790 94.170 112.930 ;
        RECT 90.645 112.745 90.935 112.790 ;
        RECT 53.025 112.590 53.315 112.635 ;
        RECT 53.830 112.590 54.150 112.650 ;
        RECT 56.265 112.590 56.915 112.635 ;
        RECT 53.025 112.450 56.915 112.590 ;
        RECT 57.140 112.590 57.280 112.730 ;
        RECT 58.905 112.590 59.195 112.635 ;
        RECT 57.140 112.450 59.195 112.590 ;
        RECT 53.025 112.405 53.615 112.450 ;
        RECT 49.245 112.110 50.010 112.250 ;
        RECT 49.245 112.065 49.535 112.110 ;
        RECT 49.690 112.050 50.010 112.110 ;
        RECT 50.625 112.065 50.915 112.295 ;
        RECT 53.325 112.090 53.615 112.405 ;
        RECT 53.830 112.390 54.150 112.450 ;
        RECT 56.265 112.405 56.915 112.450 ;
        RECT 58.905 112.405 59.195 112.450 ;
        RECT 59.350 112.590 59.670 112.650 ;
        RECT 67.745 112.590 68.035 112.635 ;
        RECT 70.985 112.590 71.635 112.635 ;
        RECT 59.350 112.450 60.960 112.590 ;
        RECT 59.350 112.390 59.670 112.450 ;
        RECT 60.820 112.295 60.960 112.450 ;
        RECT 67.745 112.450 71.635 112.590 ;
        RECT 67.745 112.405 68.335 112.450 ;
        RECT 70.985 112.405 71.635 112.450 ;
        RECT 68.045 112.310 68.335 112.405 ;
        RECT 73.610 112.390 73.930 112.650 ;
        RECT 79.705 112.590 79.995 112.635 ;
        RECT 80.510 112.590 80.830 112.650 ;
        RECT 82.945 112.590 83.595 112.635 ;
        RECT 79.705 112.450 83.595 112.590 ;
        RECT 79.705 112.405 80.295 112.450 ;
        RECT 54.405 112.250 54.695 112.295 ;
        RECT 57.985 112.250 58.275 112.295 ;
        RECT 59.820 112.250 60.110 112.295 ;
        RECT 54.405 112.110 60.110 112.250 ;
        RECT 54.405 112.065 54.695 112.110 ;
        RECT 57.985 112.065 58.275 112.110 ;
        RECT 59.820 112.065 60.110 112.110 ;
        RECT 60.745 112.065 61.035 112.295 ;
        RECT 64.870 112.050 65.190 112.310 ;
        RECT 68.045 112.090 68.410 112.310 ;
        RECT 68.090 112.050 68.410 112.090 ;
        RECT 69.125 112.250 69.415 112.295 ;
        RECT 72.705 112.250 72.995 112.295 ;
        RECT 74.540 112.250 74.830 112.295 ;
        RECT 69.125 112.110 74.830 112.250 ;
        RECT 69.125 112.065 69.415 112.110 ;
        RECT 72.705 112.065 72.995 112.110 ;
        RECT 74.540 112.065 74.830 112.110 ;
        RECT 75.005 112.250 75.295 112.295 ;
        RECT 75.450 112.250 75.770 112.310 ;
        RECT 75.005 112.110 75.770 112.250 ;
        RECT 75.005 112.065 75.295 112.110 ;
        RECT 75.450 112.050 75.770 112.110 ;
        RECT 77.765 112.250 78.055 112.295 ;
        RECT 79.130 112.250 79.450 112.310 ;
        RECT 77.765 112.110 79.450 112.250 ;
        RECT 77.765 112.065 78.055 112.110 ;
        RECT 79.130 112.050 79.450 112.110 ;
        RECT 80.005 112.090 80.295 112.405 ;
        RECT 80.510 112.390 80.830 112.450 ;
        RECT 82.945 112.405 83.595 112.450 ;
        RECT 85.585 112.590 85.875 112.635 ;
        RECT 87.500 112.590 87.640 112.745 ;
        RECT 93.850 112.730 94.170 112.790 ;
        RECT 96.150 112.930 96.470 112.990 ;
        RECT 99.845 112.930 100.135 112.975 ;
        RECT 96.150 112.790 100.135 112.930 ;
        RECT 96.150 112.730 96.470 112.790 ;
        RECT 99.845 112.745 100.135 112.790 ;
        RECT 101.685 112.930 101.975 112.975 ;
        RECT 104.430 112.930 104.750 112.990 ;
        RECT 101.685 112.790 104.750 112.930 ;
        RECT 101.685 112.745 101.975 112.790 ;
        RECT 104.430 112.730 104.750 112.790 ;
        RECT 114.105 112.930 114.395 112.975 ;
        RECT 118.230 112.930 118.550 112.990 ;
        RECT 114.105 112.790 118.550 112.930 ;
        RECT 114.105 112.745 114.395 112.790 ;
        RECT 118.230 112.730 118.550 112.790 ;
        RECT 85.585 112.450 87.640 112.590 ;
        RECT 92.125 112.590 92.415 112.635 ;
        RECT 94.310 112.590 94.630 112.650 ;
        RECT 95.365 112.590 96.015 112.635 ;
        RECT 92.125 112.450 96.015 112.590 ;
        RECT 85.585 112.405 85.875 112.450 ;
        RECT 92.125 112.405 92.715 112.450 ;
        RECT 81.085 112.250 81.375 112.295 ;
        RECT 84.665 112.250 84.955 112.295 ;
        RECT 86.500 112.250 86.790 112.295 ;
        RECT 81.085 112.110 86.790 112.250 ;
        RECT 81.085 112.065 81.375 112.110 ;
        RECT 84.665 112.065 84.955 112.110 ;
        RECT 86.500 112.065 86.790 112.110 ;
        RECT 86.965 112.250 87.255 112.295 ;
        RECT 87.870 112.250 88.190 112.310 ;
        RECT 86.965 112.110 88.190 112.250 ;
        RECT 86.965 112.065 87.255 112.110 ;
        RECT 87.870 112.050 88.190 112.110 ;
        RECT 88.330 112.050 88.650 112.310 ;
        RECT 90.170 112.050 90.490 112.310 ;
        RECT 92.425 112.090 92.715 112.405 ;
        RECT 94.310 112.390 94.630 112.450 ;
        RECT 95.365 112.405 96.015 112.450 ;
        RECT 96.610 112.590 96.930 112.650 ;
        RECT 98.005 112.590 98.295 112.635 ;
        RECT 96.610 112.450 98.295 112.590 ;
        RECT 96.610 112.390 96.930 112.450 ;
        RECT 98.005 112.405 98.295 112.450 ;
        RECT 98.450 112.590 98.770 112.650 ;
        RECT 103.165 112.590 103.455 112.635 ;
        RECT 105.350 112.590 105.670 112.650 ;
        RECT 106.405 112.590 107.055 112.635 ;
        RECT 98.450 112.450 100.980 112.590 ;
        RECT 98.450 112.390 98.770 112.450 ;
        RECT 100.840 112.295 100.980 112.450 ;
        RECT 103.165 112.450 107.055 112.590 ;
        RECT 103.165 112.405 103.755 112.450 ;
        RECT 93.505 112.250 93.795 112.295 ;
        RECT 97.085 112.250 97.375 112.295 ;
        RECT 98.920 112.250 99.210 112.295 ;
        RECT 93.505 112.110 99.210 112.250 ;
        RECT 93.505 112.065 93.795 112.110 ;
        RECT 97.085 112.065 97.375 112.110 ;
        RECT 98.920 112.065 99.210 112.110 ;
        RECT 100.765 112.065 101.055 112.295 ;
        RECT 103.465 112.090 103.755 112.405 ;
        RECT 105.350 112.390 105.670 112.450 ;
        RECT 106.405 112.405 107.055 112.450 ;
        RECT 109.045 112.590 109.335 112.635 ;
        RECT 109.490 112.590 109.810 112.650 ;
        RECT 109.045 112.450 109.810 112.590 ;
        RECT 109.045 112.405 109.335 112.450 ;
        RECT 109.490 112.390 109.810 112.450 ;
        RECT 118.805 112.590 119.095 112.635 ;
        RECT 119.610 112.590 119.930 112.650 ;
        RECT 122.045 112.590 122.695 112.635 ;
        RECT 118.805 112.450 122.695 112.590 ;
        RECT 118.805 112.405 119.395 112.450 ;
        RECT 104.545 112.250 104.835 112.295 ;
        RECT 108.125 112.250 108.415 112.295 ;
        RECT 109.960 112.250 110.250 112.295 ;
        RECT 104.545 112.110 110.250 112.250 ;
        RECT 104.545 112.065 104.835 112.110 ;
        RECT 108.125 112.065 108.415 112.110 ;
        RECT 109.960 112.065 110.250 112.110 ;
        RECT 110.410 112.050 110.730 112.310 ;
        RECT 110.885 112.250 111.175 112.295 ;
        RECT 111.330 112.250 111.650 112.310 ;
        RECT 110.885 112.110 111.650 112.250 ;
        RECT 110.885 112.065 111.175 112.110 ;
        RECT 111.330 112.050 111.650 112.110 ;
        RECT 113.185 112.250 113.475 112.295 ;
        RECT 114.550 112.250 114.870 112.310 ;
        RECT 113.185 112.110 114.870 112.250 ;
        RECT 113.185 112.065 113.475 112.110 ;
        RECT 114.550 112.050 114.870 112.110 ;
        RECT 115.485 112.250 115.775 112.295 ;
        RECT 116.850 112.250 117.170 112.310 ;
        RECT 115.485 112.110 117.170 112.250 ;
        RECT 115.485 112.065 115.775 112.110 ;
        RECT 116.850 112.050 117.170 112.110 ;
        RECT 119.105 112.090 119.395 112.405 ;
        RECT 119.610 112.390 119.930 112.450 ;
        RECT 122.045 112.405 122.695 112.450 ;
        RECT 124.670 112.390 124.990 112.650 ;
        RECT 120.185 112.250 120.475 112.295 ;
        RECT 123.765 112.250 124.055 112.295 ;
        RECT 125.600 112.250 125.890 112.295 ;
        RECT 120.185 112.110 125.890 112.250 ;
        RECT 120.185 112.065 120.475 112.110 ;
        RECT 123.765 112.065 124.055 112.110 ;
        RECT 125.600 112.065 125.890 112.110 ;
        RECT 24.390 111.710 24.710 111.970 ;
        RECT 35.430 111.910 35.750 111.970 ;
        RECT 36.825 111.910 37.115 111.955 ;
        RECT 35.430 111.770 37.115 111.910 ;
        RECT 35.430 111.710 35.750 111.770 ;
        RECT 36.825 111.725 37.115 111.770 ;
        RECT 42.790 111.910 43.110 111.970 ;
        RECT 42.790 111.770 49.920 111.910 ;
        RECT 42.790 111.710 43.110 111.770 ;
        RECT 49.780 111.615 49.920 111.770 ;
        RECT 60.270 111.710 60.590 111.970 ;
        RECT 66.265 111.910 66.555 111.955 ;
        RECT 71.310 111.910 71.630 111.970 ;
        RECT 66.265 111.770 71.630 111.910 ;
        RECT 66.265 111.725 66.555 111.770 ;
        RECT 71.310 111.710 71.630 111.770 ;
        RECT 77.305 111.910 77.595 111.955 ;
        RECT 78.210 111.910 78.530 111.970 ;
        RECT 77.305 111.770 78.530 111.910 ;
        RECT 77.305 111.725 77.595 111.770 ;
        RECT 78.210 111.710 78.530 111.770 ;
        RECT 89.710 111.710 90.030 111.970 ;
        RECT 99.385 111.910 99.675 111.955 ;
        RECT 110.500 111.910 110.640 112.050 ;
        RECT 114.090 111.910 114.410 111.970 ;
        RECT 99.385 111.770 114.410 111.910 ;
        RECT 99.385 111.725 99.675 111.770 ;
        RECT 114.090 111.710 114.410 111.770 ;
        RECT 115.945 111.910 116.235 111.955 ;
        RECT 116.390 111.910 116.710 111.970 ;
        RECT 115.945 111.770 116.710 111.910 ;
        RECT 115.945 111.725 116.235 111.770 ;
        RECT 116.390 111.710 116.710 111.770 ;
        RECT 117.325 111.910 117.615 111.955 ;
        RECT 120.990 111.910 121.310 111.970 ;
        RECT 117.325 111.770 121.310 111.910 ;
        RECT 117.325 111.725 117.615 111.770 ;
        RECT 120.990 111.710 121.310 111.770 ;
        RECT 124.670 111.910 124.990 111.970 ;
        RECT 126.065 111.910 126.355 111.955 ;
        RECT 124.670 111.770 126.355 111.910 ;
        RECT 124.670 111.710 124.990 111.770 ;
        RECT 126.065 111.725 126.355 111.770 ;
        RECT 30.945 111.570 31.235 111.615 ;
        RECT 34.065 111.570 34.355 111.615 ;
        RECT 35.955 111.570 36.245 111.615 ;
        RECT 30.945 111.430 36.245 111.570 ;
        RECT 30.945 111.385 31.235 111.430 ;
        RECT 34.065 111.385 34.355 111.430 ;
        RECT 35.955 111.385 36.245 111.430 ;
        RECT 43.365 111.570 43.655 111.615 ;
        RECT 46.485 111.570 46.775 111.615 ;
        RECT 48.375 111.570 48.665 111.615 ;
        RECT 43.365 111.430 48.665 111.570 ;
        RECT 43.365 111.385 43.655 111.430 ;
        RECT 46.485 111.385 46.775 111.430 ;
        RECT 48.375 111.385 48.665 111.430 ;
        RECT 49.705 111.570 49.995 111.615 ;
        RECT 54.405 111.570 54.695 111.615 ;
        RECT 57.525 111.570 57.815 111.615 ;
        RECT 59.415 111.570 59.705 111.615 ;
        RECT 49.705 111.430 50.105 111.570 ;
        RECT 54.405 111.430 59.705 111.570 ;
        RECT 49.705 111.385 49.995 111.430 ;
        RECT 54.405 111.385 54.695 111.430 ;
        RECT 57.525 111.385 57.815 111.430 ;
        RECT 59.415 111.385 59.705 111.430 ;
        RECT 69.125 111.570 69.415 111.615 ;
        RECT 72.245 111.570 72.535 111.615 ;
        RECT 74.135 111.570 74.425 111.615 ;
        RECT 69.125 111.430 74.425 111.570 ;
        RECT 69.125 111.385 69.415 111.430 ;
        RECT 72.245 111.385 72.535 111.430 ;
        RECT 74.135 111.385 74.425 111.430 ;
        RECT 81.085 111.570 81.375 111.615 ;
        RECT 84.205 111.570 84.495 111.615 ;
        RECT 86.095 111.570 86.385 111.615 ;
        RECT 81.085 111.430 86.385 111.570 ;
        RECT 81.085 111.385 81.375 111.430 ;
        RECT 84.205 111.385 84.495 111.430 ;
        RECT 86.095 111.385 86.385 111.430 ;
        RECT 93.505 111.570 93.795 111.615 ;
        RECT 96.625 111.570 96.915 111.615 ;
        RECT 98.515 111.570 98.805 111.615 ;
        RECT 93.505 111.430 98.805 111.570 ;
        RECT 93.505 111.385 93.795 111.430 ;
        RECT 96.625 111.385 96.915 111.430 ;
        RECT 98.515 111.385 98.805 111.430 ;
        RECT 104.545 111.570 104.835 111.615 ;
        RECT 107.665 111.570 107.955 111.615 ;
        RECT 109.555 111.570 109.845 111.615 ;
        RECT 120.185 111.570 120.475 111.615 ;
        RECT 123.305 111.570 123.595 111.615 ;
        RECT 125.195 111.570 125.485 111.615 ;
        RECT 104.545 111.430 109.845 111.570 ;
        RECT 104.545 111.385 104.835 111.430 ;
        RECT 107.665 111.385 107.955 111.430 ;
        RECT 109.555 111.385 109.845 111.430 ;
        RECT 111.420 111.430 112.940 111.570 ;
        RECT 61.665 111.230 61.955 111.275 ;
        RECT 63.950 111.230 64.270 111.290 ;
        RECT 61.665 111.090 64.270 111.230 ;
        RECT 61.665 111.045 61.955 111.090 ;
        RECT 63.950 111.030 64.270 111.090 ;
        RECT 65.790 111.030 66.110 111.290 ;
        RECT 79.590 111.230 79.910 111.290 ;
        RECT 111.420 111.230 111.560 111.430 ;
        RECT 79.590 111.090 111.560 111.230 ;
        RECT 111.805 111.230 112.095 111.275 ;
        RECT 112.250 111.230 112.570 111.290 ;
        RECT 111.805 111.090 112.570 111.230 ;
        RECT 112.800 111.230 112.940 111.430 ;
        RECT 120.185 111.430 125.485 111.570 ;
        RECT 120.185 111.385 120.475 111.430 ;
        RECT 123.305 111.385 123.595 111.430 ;
        RECT 125.195 111.385 125.485 111.430 ;
        RECT 124.210 111.230 124.530 111.290 ;
        RECT 112.800 111.090 124.530 111.230 ;
        RECT 79.590 111.030 79.910 111.090 ;
        RECT 111.805 111.045 112.095 111.090 ;
        RECT 112.250 111.030 112.570 111.090 ;
        RECT 124.210 111.030 124.530 111.090 ;
        RECT 20.640 110.410 127.820 110.890 ;
        RECT 33.590 110.210 33.910 110.270 ;
        RECT 35.430 110.210 35.750 110.270 ;
        RECT 53.830 110.210 54.150 110.270 ;
        RECT 54.305 110.210 54.595 110.255 ;
        RECT 31.840 110.070 41.180 110.210 ;
        RECT 31.840 109.575 31.980 110.070 ;
        RECT 33.590 110.010 33.910 110.070 ;
        RECT 35.430 110.010 35.750 110.070 ;
        RECT 32.635 109.870 32.925 109.915 ;
        RECT 34.525 109.870 34.815 109.915 ;
        RECT 37.645 109.870 37.935 109.915 ;
        RECT 32.635 109.730 37.935 109.870 ;
        RECT 32.635 109.685 32.925 109.730 ;
        RECT 34.525 109.685 34.815 109.730 ;
        RECT 37.645 109.685 37.935 109.730 ;
        RECT 31.765 109.345 32.055 109.575 ;
        RECT 33.145 109.530 33.435 109.575 ;
        RECT 35.890 109.530 36.210 109.590 ;
        RECT 41.040 109.575 41.180 110.070 ;
        RECT 53.830 110.070 54.595 110.210 ;
        RECT 53.830 110.010 54.150 110.070 ;
        RECT 54.305 110.025 54.595 110.070 ;
        RECT 60.270 110.210 60.590 110.270 ;
        RECT 87.870 110.210 88.190 110.270 ;
        RECT 124.670 110.210 124.990 110.270 ;
        RECT 60.270 110.070 65.560 110.210 ;
        RECT 60.270 110.010 60.590 110.070 ;
        RECT 41.835 109.870 42.125 109.915 ;
        RECT 43.725 109.870 44.015 109.915 ;
        RECT 46.845 109.870 47.135 109.915 ;
        RECT 41.835 109.730 47.135 109.870 ;
        RECT 41.835 109.685 42.125 109.730 ;
        RECT 43.725 109.685 44.015 109.730 ;
        RECT 46.845 109.685 47.135 109.730 ;
        RECT 59.465 109.870 59.755 109.915 ;
        RECT 62.585 109.870 62.875 109.915 ;
        RECT 64.475 109.870 64.765 109.915 ;
        RECT 59.465 109.730 64.765 109.870 ;
        RECT 59.465 109.685 59.755 109.730 ;
        RECT 62.585 109.685 62.875 109.730 ;
        RECT 64.475 109.685 64.765 109.730 ;
        RECT 33.145 109.390 36.210 109.530 ;
        RECT 33.145 109.345 33.435 109.390 ;
        RECT 35.890 109.330 36.210 109.390 ;
        RECT 40.965 109.345 41.255 109.575 ;
        RECT 42.345 109.530 42.635 109.575 ;
        RECT 42.790 109.530 43.110 109.590 ;
        RECT 42.345 109.390 43.110 109.530 ;
        RECT 42.345 109.345 42.635 109.390 ;
        RECT 42.790 109.330 43.110 109.390 ;
        RECT 63.950 109.330 64.270 109.590 ;
        RECT 65.420 109.575 65.560 110.070 ;
        RECT 85.660 110.070 88.190 110.210 ;
        RECT 68.665 109.870 68.955 109.915 ;
        RECT 71.785 109.870 72.075 109.915 ;
        RECT 73.675 109.870 73.965 109.915 ;
        RECT 68.665 109.730 73.965 109.870 ;
        RECT 68.665 109.685 68.955 109.730 ;
        RECT 71.785 109.685 72.075 109.730 ;
        RECT 73.675 109.685 73.965 109.730 ;
        RECT 79.245 109.870 79.535 109.915 ;
        RECT 82.365 109.870 82.655 109.915 ;
        RECT 84.255 109.870 84.545 109.915 ;
        RECT 79.245 109.730 84.545 109.870 ;
        RECT 79.245 109.685 79.535 109.730 ;
        RECT 82.365 109.685 82.655 109.730 ;
        RECT 84.255 109.685 84.545 109.730 ;
        RECT 65.345 109.345 65.635 109.575 ;
        RECT 65.790 109.530 66.110 109.590 ;
        RECT 73.165 109.530 73.455 109.575 ;
        RECT 65.790 109.390 73.455 109.530 ;
        RECT 65.790 109.330 66.110 109.390 ;
        RECT 73.165 109.345 73.455 109.390 ;
        RECT 74.545 109.530 74.835 109.575 ;
        RECT 76.370 109.530 76.690 109.590 ;
        RECT 74.545 109.390 76.690 109.530 ;
        RECT 74.545 109.345 74.835 109.390 ;
        RECT 76.370 109.330 76.690 109.390 ;
        RECT 83.730 109.330 84.050 109.590 ;
        RECT 85.660 109.575 85.800 110.070 ;
        RECT 87.870 110.010 88.190 110.070 ;
        RECT 116.940 110.070 124.990 110.210 ;
        RECT 86.455 109.870 86.745 109.915 ;
        RECT 88.345 109.870 88.635 109.915 ;
        RECT 91.465 109.870 91.755 109.915 ;
        RECT 86.455 109.730 91.755 109.870 ;
        RECT 86.455 109.685 86.745 109.730 ;
        RECT 88.345 109.685 88.635 109.730 ;
        RECT 91.465 109.685 91.755 109.730 ;
        RECT 108.225 109.870 108.515 109.915 ;
        RECT 111.345 109.870 111.635 109.915 ;
        RECT 113.235 109.870 113.525 109.915 ;
        RECT 108.225 109.730 113.525 109.870 ;
        RECT 108.225 109.685 108.515 109.730 ;
        RECT 111.345 109.685 111.635 109.730 ;
        RECT 113.235 109.685 113.525 109.730 ;
        RECT 85.125 109.530 85.415 109.575 ;
        RECT 85.585 109.530 85.875 109.575 ;
        RECT 85.125 109.390 85.875 109.530 ;
        RECT 85.125 109.345 85.415 109.390 ;
        RECT 85.585 109.345 85.875 109.390 ;
        RECT 86.950 109.330 87.270 109.590 ;
        RECT 112.250 109.530 112.570 109.590 ;
        RECT 112.725 109.530 113.015 109.575 ;
        RECT 112.250 109.390 113.015 109.530 ;
        RECT 112.250 109.330 112.570 109.390 ;
        RECT 112.725 109.345 113.015 109.390 ;
        RECT 114.090 109.530 114.410 109.590 ;
        RECT 116.940 109.530 117.080 110.070 ;
        RECT 117.425 109.870 117.715 109.915 ;
        RECT 120.545 109.870 120.835 109.915 ;
        RECT 122.435 109.870 122.725 109.915 ;
        RECT 117.425 109.730 122.725 109.870 ;
        RECT 117.425 109.685 117.715 109.730 ;
        RECT 120.545 109.685 120.835 109.730 ;
        RECT 122.435 109.685 122.725 109.730 ;
        RECT 114.090 109.390 117.080 109.530 ;
        RECT 118.230 109.530 118.550 109.590 ;
        RECT 123.380 109.575 123.520 110.070 ;
        RECT 124.670 110.010 124.990 110.070 ;
        RECT 124.210 109.870 124.530 109.930 ;
        RECT 125.145 109.870 125.435 109.915 ;
        RECT 124.210 109.730 125.435 109.870 ;
        RECT 124.210 109.670 124.530 109.730 ;
        RECT 125.145 109.685 125.435 109.730 ;
        RECT 121.925 109.530 122.215 109.575 ;
        RECT 118.230 109.390 122.215 109.530 ;
        RECT 114.090 109.330 114.410 109.390 ;
        RECT 118.230 109.330 118.550 109.390 ;
        RECT 121.925 109.345 122.215 109.390 ;
        RECT 123.305 109.345 123.595 109.575 ;
        RECT 30.385 109.190 30.675 109.235 ;
        RECT 30.830 109.190 31.150 109.250 ;
        RECT 30.385 109.050 31.150 109.190 ;
        RECT 30.385 109.005 30.675 109.050 ;
        RECT 30.830 108.990 31.150 109.050 ;
        RECT 32.230 109.190 32.520 109.235 ;
        RECT 34.065 109.190 34.355 109.235 ;
        RECT 37.645 109.190 37.935 109.235 ;
        RECT 32.230 109.050 37.935 109.190 ;
        RECT 32.230 109.005 32.520 109.050 ;
        RECT 34.065 109.005 34.355 109.050 ;
        RECT 37.645 109.005 37.935 109.050 ;
        RECT 38.650 109.210 38.970 109.250 ;
        RECT 38.650 108.990 39.015 109.210 ;
        RECT 41.430 109.190 41.720 109.235 ;
        RECT 43.265 109.190 43.555 109.235 ;
        RECT 46.845 109.190 47.135 109.235 ;
        RECT 41.430 109.050 47.135 109.190 ;
        RECT 41.430 109.005 41.720 109.050 ;
        RECT 43.265 109.005 43.555 109.050 ;
        RECT 46.845 109.005 47.135 109.050 ;
        RECT 38.725 108.895 39.015 108.990 ;
        RECT 47.925 108.895 48.215 109.210 ;
        RECT 53.845 109.190 54.135 109.235 ;
        RECT 55.225 109.190 55.515 109.235 ;
        RECT 57.510 109.190 57.830 109.250 ;
        RECT 53.845 109.050 57.830 109.190 ;
        RECT 53.845 109.005 54.135 109.050 ;
        RECT 55.225 109.005 55.515 109.050 ;
        RECT 57.510 108.990 57.830 109.050 ;
        RECT 35.425 108.850 36.075 108.895 ;
        RECT 38.725 108.850 39.315 108.895 ;
        RECT 35.425 108.710 39.315 108.850 ;
        RECT 35.425 108.665 36.075 108.710 ;
        RECT 39.025 108.665 39.315 108.710 ;
        RECT 44.625 108.850 45.275 108.895 ;
        RECT 47.925 108.850 48.515 108.895 ;
        RECT 49.230 108.850 49.550 108.910 ;
        RECT 58.385 108.895 58.675 109.210 ;
        RECT 59.465 109.190 59.755 109.235 ;
        RECT 63.045 109.190 63.335 109.235 ;
        RECT 64.880 109.190 65.170 109.235 ;
        RECT 59.465 109.050 65.170 109.190 ;
        RECT 59.465 109.005 59.755 109.050 ;
        RECT 63.045 109.005 63.335 109.050 ;
        RECT 64.880 109.005 65.170 109.050 ;
        RECT 44.625 108.710 49.550 108.850 ;
        RECT 44.625 108.665 45.275 108.710 ;
        RECT 48.225 108.665 48.515 108.710 ;
        RECT 49.230 108.650 49.550 108.710 ;
        RECT 55.685 108.850 55.975 108.895 ;
        RECT 58.085 108.850 58.675 108.895 ;
        RECT 61.325 108.850 61.975 108.895 ;
        RECT 55.685 108.710 61.975 108.850 ;
        RECT 55.685 108.665 55.975 108.710 ;
        RECT 58.085 108.665 58.375 108.710 ;
        RECT 61.325 108.665 61.975 108.710 ;
        RECT 66.250 108.850 66.570 108.910 ;
        RECT 67.585 108.895 67.875 109.210 ;
        RECT 68.665 109.190 68.955 109.235 ;
        RECT 72.245 109.190 72.535 109.235 ;
        RECT 74.080 109.190 74.370 109.235 ;
        RECT 78.210 109.210 78.530 109.250 ;
        RECT 68.665 109.050 74.370 109.190 ;
        RECT 68.665 109.005 68.955 109.050 ;
        RECT 72.245 109.005 72.535 109.050 ;
        RECT 74.080 109.005 74.370 109.050 ;
        RECT 78.165 108.990 78.530 109.210 ;
        RECT 79.245 109.190 79.535 109.235 ;
        RECT 82.825 109.190 83.115 109.235 ;
        RECT 84.660 109.190 84.950 109.235 ;
        RECT 79.245 109.050 84.950 109.190 ;
        RECT 79.245 109.005 79.535 109.050 ;
        RECT 82.825 109.005 83.115 109.050 ;
        RECT 84.660 109.005 84.950 109.050 ;
        RECT 86.050 109.190 86.340 109.235 ;
        RECT 87.885 109.190 88.175 109.235 ;
        RECT 91.465 109.190 91.755 109.235 ;
        RECT 86.050 109.050 91.755 109.190 ;
        RECT 86.050 109.005 86.340 109.050 ;
        RECT 87.885 109.005 88.175 109.050 ;
        RECT 91.465 109.005 91.755 109.050 ;
        RECT 78.165 108.895 78.455 108.990 ;
        RECT 89.710 108.895 90.030 108.910 ;
        RECT 67.285 108.850 67.875 108.895 ;
        RECT 70.525 108.850 71.175 108.895 ;
        RECT 66.250 108.710 71.175 108.850 ;
        RECT 66.250 108.650 66.570 108.710 ;
        RECT 67.285 108.665 67.575 108.710 ;
        RECT 70.525 108.665 71.175 108.710 ;
        RECT 77.865 108.850 78.455 108.895 ;
        RECT 81.105 108.850 81.755 108.895 ;
        RECT 77.865 108.710 81.755 108.850 ;
        RECT 77.865 108.665 78.155 108.710 ;
        RECT 81.105 108.665 81.755 108.710 ;
        RECT 89.245 108.850 90.030 108.895 ;
        RECT 92.545 108.895 92.835 109.210 ;
        RECT 107.145 108.895 107.435 109.210 ;
        RECT 108.225 109.190 108.515 109.235 ;
        RECT 111.805 109.190 112.095 109.235 ;
        RECT 113.640 109.190 113.930 109.235 ;
        RECT 116.390 109.210 116.710 109.250 ;
        RECT 108.225 109.050 113.930 109.190 ;
        RECT 108.225 109.005 108.515 109.050 ;
        RECT 111.805 109.005 112.095 109.050 ;
        RECT 113.640 109.005 113.930 109.050 ;
        RECT 116.345 108.990 116.710 109.210 ;
        RECT 117.425 109.190 117.715 109.235 ;
        RECT 121.005 109.190 121.295 109.235 ;
        RECT 122.840 109.190 123.130 109.235 ;
        RECT 117.425 109.050 123.130 109.190 ;
        RECT 117.425 109.005 117.715 109.050 ;
        RECT 121.005 109.005 121.295 109.050 ;
        RECT 122.840 109.005 123.130 109.050 ;
        RECT 126.065 109.190 126.355 109.235 ;
        RECT 131.110 109.190 131.430 109.250 ;
        RECT 126.065 109.050 131.430 109.190 ;
        RECT 126.065 109.005 126.355 109.050 ;
        RECT 131.110 108.990 131.430 109.050 ;
        RECT 92.545 108.850 93.135 108.895 ;
        RECT 89.245 108.710 93.135 108.850 ;
        RECT 89.245 108.665 90.030 108.710 ;
        RECT 92.845 108.665 93.135 108.710 ;
        RECT 106.845 108.850 107.435 108.895 ;
        RECT 109.030 108.850 109.350 108.910 ;
        RECT 116.345 108.895 116.635 108.990 ;
        RECT 110.085 108.850 110.735 108.895 ;
        RECT 106.845 108.710 110.735 108.850 ;
        RECT 106.845 108.665 107.135 108.710 ;
        RECT 89.710 108.650 90.030 108.665 ;
        RECT 109.030 108.650 109.350 108.710 ;
        RECT 110.085 108.665 110.735 108.710 ;
        RECT 116.045 108.850 116.635 108.895 ;
        RECT 119.285 108.850 119.935 108.895 ;
        RECT 116.045 108.710 119.935 108.850 ;
        RECT 116.045 108.665 116.335 108.710 ;
        RECT 119.285 108.665 119.935 108.710 ;
        RECT 31.305 108.510 31.595 108.555 ;
        RECT 32.210 108.510 32.530 108.570 ;
        RECT 31.305 108.370 32.530 108.510 ;
        RECT 31.305 108.325 31.595 108.370 ;
        RECT 32.210 108.310 32.530 108.370 ;
        RECT 38.190 108.510 38.510 108.570 ;
        RECT 40.505 108.510 40.795 108.555 ;
        RECT 38.190 108.370 40.795 108.510 ;
        RECT 38.190 108.310 38.510 108.370 ;
        RECT 40.505 108.325 40.795 108.370 ;
        RECT 49.690 108.310 50.010 108.570 ;
        RECT 56.605 108.510 56.895 108.555 ;
        RECT 60.270 108.510 60.590 108.570 ;
        RECT 56.605 108.370 60.590 108.510 ;
        RECT 56.605 108.325 56.895 108.370 ;
        RECT 60.270 108.310 60.590 108.370 ;
        RECT 65.790 108.310 66.110 108.570 ;
        RECT 76.370 108.310 76.690 108.570 ;
        RECT 88.330 108.510 88.650 108.570 ;
        RECT 94.325 108.510 94.615 108.555 ;
        RECT 88.330 108.370 94.615 108.510 ;
        RECT 88.330 108.310 88.650 108.370 ;
        RECT 94.325 108.325 94.615 108.370 ;
        RECT 105.365 108.510 105.655 108.555 ;
        RECT 109.490 108.510 109.810 108.570 ;
        RECT 105.365 108.370 109.810 108.510 ;
        RECT 105.365 108.325 105.655 108.370 ;
        RECT 109.490 108.310 109.810 108.370 ;
        RECT 114.565 108.510 114.855 108.555 ;
        RECT 115.470 108.510 115.790 108.570 ;
        RECT 114.565 108.370 115.790 108.510 ;
        RECT 114.565 108.325 114.855 108.370 ;
        RECT 115.470 108.310 115.790 108.370 ;
        RECT 20.640 107.690 127.820 108.170 ;
        RECT 65.805 107.490 66.095 107.535 ;
        RECT 66.250 107.490 66.570 107.550 ;
        RECT 65.805 107.350 66.570 107.490 ;
        RECT 65.805 107.305 66.095 107.350 ;
        RECT 66.250 107.290 66.570 107.350 ;
        RECT 67.645 107.490 67.935 107.535 ;
        RECT 68.090 107.490 68.410 107.550 ;
        RECT 67.645 107.350 68.410 107.490 ;
        RECT 67.645 107.305 67.935 107.350 ;
        RECT 68.090 107.290 68.410 107.350 ;
        RECT 24.390 107.150 24.710 107.210 ;
        RECT 26.345 107.150 26.635 107.195 ;
        RECT 29.585 107.150 30.235 107.195 ;
        RECT 24.390 107.010 30.235 107.150 ;
        RECT 24.390 106.950 24.710 107.010 ;
        RECT 26.345 106.965 26.935 107.010 ;
        RECT 29.585 106.965 30.235 107.010 ;
        RECT 26.645 106.650 26.935 106.965 ;
        RECT 32.210 106.950 32.530 107.210 ;
        RECT 96.145 107.150 96.795 107.195 ;
        RECT 98.910 107.150 99.230 107.210 ;
        RECT 99.745 107.150 100.035 107.195 ;
        RECT 96.145 107.010 100.035 107.150 ;
        RECT 96.145 106.965 96.795 107.010 ;
        RECT 98.910 106.950 99.230 107.010 ;
        RECT 99.445 106.965 100.035 107.010 ;
        RECT 27.725 106.810 28.015 106.855 ;
        RECT 31.305 106.810 31.595 106.855 ;
        RECT 33.140 106.810 33.430 106.855 ;
        RECT 27.725 106.670 33.430 106.810 ;
        RECT 27.725 106.625 28.015 106.670 ;
        RECT 31.305 106.625 31.595 106.670 ;
        RECT 33.140 106.625 33.430 106.670 ;
        RECT 33.590 106.610 33.910 106.870 ;
        RECT 57.510 106.810 57.830 106.870 ;
        RECT 65.345 106.810 65.635 106.855 ;
        RECT 67.185 106.810 67.475 106.855 ;
        RECT 57.510 106.670 67.475 106.810 ;
        RECT 57.510 106.610 57.830 106.670 ;
        RECT 65.345 106.625 65.635 106.670 ;
        RECT 67.185 106.625 67.475 106.670 ;
        RECT 87.870 106.810 88.190 106.870 ;
        RECT 92.485 106.810 92.775 106.855 ;
        RECT 87.870 106.670 92.775 106.810 ;
        RECT 87.870 106.610 88.190 106.670 ;
        RECT 92.485 106.625 92.775 106.670 ;
        RECT 92.950 106.810 93.240 106.855 ;
        RECT 94.785 106.810 95.075 106.855 ;
        RECT 98.365 106.810 98.655 106.855 ;
        RECT 92.950 106.670 98.655 106.810 ;
        RECT 92.950 106.625 93.240 106.670 ;
        RECT 94.785 106.625 95.075 106.670 ;
        RECT 98.365 106.625 98.655 106.670 ;
        RECT 99.445 106.650 99.735 106.965 ;
        RECT 135.660 106.690 136.800 133.400 ;
        RECT 133.100 106.600 136.850 106.690 ;
        RECT 93.865 106.470 94.155 106.515 ;
        RECT 96.150 106.470 96.470 106.530 ;
        RECT 93.865 106.330 96.470 106.470 ;
        RECT 93.865 106.285 94.155 106.330 ;
        RECT 96.150 106.270 96.470 106.330 ;
        RECT 27.725 106.130 28.015 106.175 ;
        RECT 30.845 106.130 31.135 106.175 ;
        RECT 32.735 106.130 33.025 106.175 ;
        RECT 27.725 105.990 33.025 106.130 ;
        RECT 27.725 105.945 28.015 105.990 ;
        RECT 30.845 105.945 31.135 105.990 ;
        RECT 32.735 105.945 33.025 105.990 ;
        RECT 93.355 106.130 93.645 106.175 ;
        RECT 95.245 106.130 95.535 106.175 ;
        RECT 98.365 106.130 98.655 106.175 ;
        RECT 93.355 105.990 98.655 106.130 ;
        RECT 93.355 105.945 93.645 105.990 ;
        RECT 95.245 105.945 95.535 105.990 ;
        RECT 98.365 105.945 98.655 105.990 ;
        RECT 21.630 105.790 21.950 105.850 ;
        RECT 24.865 105.790 25.155 105.835 ;
        RECT 21.630 105.650 25.155 105.790 ;
        RECT 21.630 105.590 21.950 105.650 ;
        RECT 24.865 105.605 25.155 105.650 ;
        RECT 98.910 105.790 99.230 105.850 ;
        RECT 101.225 105.790 101.515 105.835 ;
        RECT 98.910 105.650 101.515 105.790 ;
        RECT 98.910 105.590 99.230 105.650 ;
        RECT 101.225 105.605 101.515 105.650 ;
        RECT 129.700 105.630 136.850 106.600 ;
        RECT 133.100 105.500 136.850 105.630 ;
        RECT 20.640 104.970 127.820 105.450 ;
        RECT 133.330 76.630 136.060 77.830 ;
        RECT 137.920 77.810 143.450 77.960 ;
        RECT 21.115 74.380 23.065 74.390 ;
        RECT 19.415 73.240 23.065 74.380 ;
        RECT 19.415 73.230 21.125 73.240 ;
        RECT 28.135 73.230 30.305 74.410 ;
        RECT 32.315 74.390 34.265 74.400 ;
        RECT 30.615 73.250 34.265 74.390 ;
        RECT 30.615 73.240 32.325 73.250 ;
        RECT 39.425 73.200 41.595 74.380 ;
        RECT 43.535 74.360 45.485 74.370 ;
        RECT 41.835 73.220 45.485 74.360 ;
        RECT 54.785 74.340 56.735 74.350 ;
        RECT 41.835 73.210 43.545 73.220 ;
        RECT 3.910 73.080 6.100 73.190 ;
        RECT 50.005 73.140 52.175 74.320 ;
        RECT 53.085 73.200 56.735 74.340 ;
        RECT 53.085 73.190 54.795 73.200 ;
        RECT 61.425 73.170 63.595 74.350 ;
        RECT 66.005 74.330 67.955 74.340 ;
        RECT 64.305 73.190 67.955 74.330 ;
        RECT 64.305 73.180 66.015 73.190 ;
        RECT 72.535 73.180 74.705 74.360 ;
        RECT 77.245 74.320 79.195 74.330 ;
        RECT 75.545 73.180 79.195 74.320 ;
        RECT 75.545 73.170 77.255 73.180 ;
        RECT 83.805 73.170 85.975 74.350 ;
        RECT 88.495 74.330 90.445 74.340 ;
        RECT 86.795 73.190 90.445 74.330 ;
        RECT 99.775 74.320 101.725 74.330 ;
        RECT 86.795 73.180 88.505 73.190 ;
        RECT 94.995 73.110 97.165 74.290 ;
        RECT 98.075 73.180 101.725 74.320 ;
        RECT 98.075 73.170 99.785 73.180 ;
        RECT 106.405 73.160 108.575 74.340 ;
        RECT 111.045 74.320 112.995 74.330 ;
        RECT 109.345 73.180 112.995 74.320 ;
        RECT 109.345 73.170 111.055 73.180 ;
        RECT 117.605 73.160 119.775 74.340 ;
        RECT 122.295 74.320 124.245 74.330 ;
        RECT 120.595 73.180 124.245 74.320 ;
        RECT 129.455 73.240 131.625 74.420 ;
        RECT 120.595 73.170 122.305 73.180 ;
        RECT 3.910 72.820 12.240 73.080 ;
        RECT 29.635 72.840 43.235 72.850 ;
        RECT 18.435 72.820 43.235 72.840 ;
        RECT 3.910 72.800 54.455 72.820 ;
        RECT 3.910 72.790 65.705 72.800 ;
        RECT 133.960 72.790 135.640 76.630 ;
        RECT 137.190 76.610 143.450 77.810 ;
        RECT 137.920 75.460 143.450 76.610 ;
        RECT 3.910 72.780 76.925 72.790 ;
        RECT 85.815 72.780 99.415 72.790 ;
        RECT 132.085 72.780 140.600 72.790 ;
        RECT 3.910 71.700 140.600 72.780 ;
        RECT 3.910 71.690 32.035 71.700 ;
        RECT 3.910 71.670 19.135 71.690 ;
        RECT 40.855 71.670 140.600 71.700 ;
        RECT 3.910 71.500 12.240 71.670 ;
        RECT 52.105 71.650 140.600 71.670 ;
        RECT 63.325 71.640 140.600 71.650 ;
        RECT 74.565 71.630 88.165 71.640 ;
        RECT 97.095 71.630 133.215 71.640 ;
        RECT 3.910 71.370 6.100 71.500 ;
        RECT 10.800 71.180 11.950 71.500 ;
        RECT 10.800 69.480 11.915 71.180 ;
        RECT 29.635 71.170 43.285 71.180 ;
        RECT 15.510 71.155 17.040 71.160 ;
        RECT 18.435 71.155 43.285 71.170 ;
        RECT 12.285 71.150 43.285 71.155 ;
        RECT 12.285 71.130 54.505 71.150 ;
        RECT 141.810 71.140 143.230 75.460 ;
        RECT 12.285 71.120 65.755 71.130 ;
        RECT 12.285 71.110 76.975 71.120 ;
        RECT 85.815 71.110 99.465 71.120 ;
        RECT 140.220 71.110 143.240 71.140 ;
        RECT 12.285 70.030 143.240 71.110 ;
        RECT 12.285 70.020 32.085 70.030 ;
        RECT 12.285 70.005 19.375 70.020 ;
        RECT 10.800 13.800 11.950 69.480 ;
        RECT 12.320 15.450 13.470 70.005 ;
        RECT 15.510 68.660 17.040 70.005 ;
        RECT 40.855 70.000 143.240 70.030 ;
        RECT 52.105 69.980 143.240 70.000 ;
        RECT 63.325 69.970 143.240 69.980 ;
        RECT 74.565 69.960 88.215 69.970 ;
        RECT 97.095 69.960 143.240 69.970 ;
        RECT 140.220 69.910 143.240 69.960 ;
        RECT 29.645 69.670 43.315 69.680 ;
        RECT 18.445 69.650 43.315 69.670 ;
        RECT 18.445 69.630 54.535 69.650 ;
        RECT 18.445 69.620 65.785 69.630 ;
        RECT 139.590 69.620 150.610 69.640 ;
        RECT 18.445 69.610 77.005 69.620 ;
        RECT 85.825 69.610 99.495 69.620 ;
        RECT 132.155 69.610 150.610 69.620 ;
        RECT 18.445 69.570 150.610 69.610 ;
        RECT 18.445 68.530 150.740 69.570 ;
        RECT 18.445 68.520 32.115 68.530 ;
        RECT 40.865 68.500 150.740 68.530 ;
        RECT 52.115 68.490 143.320 68.500 ;
        RECT 52.115 68.480 140.670 68.490 ;
        RECT 63.335 68.470 140.670 68.480 ;
        RECT 74.575 68.460 88.245 68.470 ;
        RECT 97.105 68.460 133.295 68.470 ;
        RECT 141.080 68.450 142.300 68.490 ;
        RECT 149.360 68.470 150.740 68.500 ;
        RECT 29.655 68.100 43.325 68.110 ;
        RECT 13.950 68.080 43.325 68.100 ;
        RECT 13.950 68.060 54.545 68.080 ;
        RECT 13.950 68.050 65.795 68.060 ;
        RECT 13.950 68.040 77.015 68.050 ;
        RECT 85.835 68.040 99.505 68.050 ;
        RECT 139.530 68.040 143.320 68.060 ;
        RECT 13.950 66.960 152.870 68.040 ;
        RECT 13.950 66.950 32.125 66.960 ;
        RECT 13.950 18.530 15.100 66.950 ;
        RECT 40.875 66.930 152.870 66.960 ;
        RECT 52.125 66.910 152.870 66.930 ;
        RECT 63.345 66.900 152.870 66.910 ;
        RECT 74.585 66.890 88.255 66.900 ;
        RECT 97.115 66.890 143.320 66.900 ;
        RECT 141.030 66.770 142.490 66.890 ;
        RECT 21.405 65.510 26.555 65.790 ;
        RECT 27.815 65.490 28.965 65.800 ;
        RECT 32.605 65.520 37.755 65.800 ;
        RECT 39.015 65.500 40.165 65.810 ;
        RECT 43.825 65.490 48.975 65.770 ;
        RECT 50.235 65.470 51.385 65.780 ;
        RECT 149.460 65.760 150.600 65.780 ;
        RECT 55.075 65.470 60.225 65.750 ;
        RECT 61.485 65.450 62.635 65.760 ;
        RECT 66.295 65.460 71.445 65.740 ;
        RECT 72.705 65.440 73.855 65.750 ;
        RECT 77.535 65.450 82.685 65.730 ;
        RECT 83.945 65.430 85.095 65.740 ;
        RECT 88.785 65.460 93.935 65.740 ;
        RECT 95.195 65.440 96.345 65.750 ;
        RECT 100.065 65.450 105.215 65.730 ;
        RECT 106.475 65.430 107.625 65.740 ;
        RECT 111.335 65.450 116.485 65.730 ;
        RECT 117.745 65.430 118.895 65.740 ;
        RECT 122.585 65.450 127.735 65.730 ;
        RECT 128.995 65.430 130.145 65.740 ;
        RECT 133.315 65.430 138.455 65.690 ;
        RECT 21.205 65.140 21.435 65.320 ;
        RECT 26.495 65.190 26.725 65.320 ;
        RECT 21.125 55.220 21.485 65.140 ;
        RECT 26.435 55.240 26.805 65.190 ;
        RECT 27.635 65.150 27.865 65.320 ;
        RECT 27.565 55.200 27.935 65.150 ;
        RECT 28.925 65.140 29.155 65.320 ;
        RECT 32.405 65.150 32.635 65.330 ;
        RECT 37.695 65.200 37.925 65.330 ;
        RECT 28.835 55.250 29.255 65.140 ;
        RECT 32.325 55.230 32.685 65.150 ;
        RECT 37.635 55.250 38.005 65.200 ;
        RECT 38.835 65.160 39.065 65.330 ;
        RECT 38.765 55.210 39.135 65.160 ;
        RECT 40.125 65.150 40.355 65.330 ;
        RECT 40.035 55.260 40.455 65.150 ;
        RECT 43.625 65.120 43.855 65.300 ;
        RECT 48.915 65.170 49.145 65.300 ;
        RECT 43.545 55.200 43.905 65.120 ;
        RECT 48.855 55.220 49.225 65.170 ;
        RECT 50.055 65.130 50.285 65.300 ;
        RECT 49.985 55.180 50.355 65.130 ;
        RECT 51.345 65.120 51.575 65.300 ;
        RECT 51.255 55.230 51.675 65.120 ;
        RECT 54.875 65.100 55.105 65.280 ;
        RECT 60.165 65.150 60.395 65.280 ;
        RECT 54.795 55.180 55.155 65.100 ;
        RECT 60.105 55.200 60.475 65.150 ;
        RECT 61.305 65.110 61.535 65.280 ;
        RECT 61.235 55.160 61.605 65.110 ;
        RECT 62.595 65.100 62.825 65.280 ;
        RECT 62.505 55.210 62.925 65.100 ;
        RECT 66.095 65.090 66.325 65.270 ;
        RECT 71.385 65.140 71.615 65.270 ;
        RECT 66.015 55.170 66.375 65.090 ;
        RECT 71.325 55.190 71.695 65.140 ;
        RECT 72.525 65.100 72.755 65.270 ;
        RECT 72.455 55.150 72.825 65.100 ;
        RECT 73.815 65.090 74.045 65.270 ;
        RECT 73.725 55.200 74.145 65.090 ;
        RECT 77.335 65.080 77.565 65.260 ;
        RECT 82.625 65.130 82.855 65.260 ;
        RECT 77.255 55.160 77.615 65.080 ;
        RECT 82.565 55.180 82.935 65.130 ;
        RECT 83.765 65.090 83.995 65.260 ;
        RECT 83.695 55.140 84.065 65.090 ;
        RECT 85.055 65.080 85.285 65.260 ;
        RECT 88.585 65.090 88.815 65.270 ;
        RECT 93.875 65.140 94.105 65.270 ;
        RECT 84.965 55.190 85.385 65.080 ;
        RECT 88.505 55.170 88.865 65.090 ;
        RECT 93.815 55.190 94.185 65.140 ;
        RECT 95.015 65.100 95.245 65.270 ;
        RECT 94.945 55.150 95.315 65.100 ;
        RECT 96.305 65.090 96.535 65.270 ;
        RECT 96.215 55.200 96.635 65.090 ;
        RECT 99.865 65.080 100.095 65.260 ;
        RECT 105.155 65.130 105.385 65.260 ;
        RECT 99.785 55.160 100.145 65.080 ;
        RECT 105.095 55.180 105.465 65.130 ;
        RECT 106.295 65.090 106.525 65.260 ;
        RECT 106.225 55.140 106.595 65.090 ;
        RECT 107.585 65.080 107.815 65.260 ;
        RECT 111.135 65.080 111.365 65.260 ;
        RECT 116.425 65.130 116.655 65.260 ;
        RECT 107.495 55.190 107.915 65.080 ;
        RECT 111.055 55.160 111.415 65.080 ;
        RECT 116.365 55.180 116.735 65.130 ;
        RECT 117.565 65.090 117.795 65.260 ;
        RECT 117.495 55.140 117.865 65.090 ;
        RECT 118.855 65.080 119.085 65.260 ;
        RECT 122.385 65.080 122.615 65.260 ;
        RECT 127.675 65.130 127.905 65.260 ;
        RECT 118.765 55.190 119.185 65.080 ;
        RECT 122.305 55.160 122.665 65.080 ;
        RECT 127.615 55.180 127.985 65.130 ;
        RECT 128.815 65.090 129.045 65.260 ;
        RECT 128.745 55.140 129.115 65.090 ;
        RECT 130.105 65.080 130.335 65.260 ;
        RECT 133.135 65.130 133.365 65.230 ;
        RECT 130.015 55.190 130.435 65.080 ;
        RECT 133.005 55.240 133.405 65.130 ;
        RECT 138.425 65.100 138.655 65.230 ;
        RECT 133.135 55.230 133.365 55.240 ;
        RECT 138.345 55.130 138.725 65.100 ;
        RECT 149.340 64.660 150.720 65.760 ;
        RECT 20.815 54.230 25.555 54.530 ;
        RECT 32.015 54.240 36.755 54.540 ;
        RECT 43.235 54.210 47.975 54.510 ;
        RECT 54.485 54.190 59.225 54.490 ;
        RECT 65.705 54.180 70.445 54.480 ;
        RECT 76.945 54.170 81.685 54.470 ;
        RECT 88.195 54.180 92.935 54.480 ;
        RECT 99.475 54.170 104.215 54.470 ;
        RECT 110.745 54.170 115.485 54.470 ;
        RECT 121.995 54.170 126.735 54.470 ;
        RECT 21.655 52.320 22.115 52.550 ;
        RECT 25.625 52.280 26.255 52.560 ;
        RECT 25.735 52.240 26.195 52.280 ;
        RECT 27.665 52.240 28.125 52.470 ;
        RECT 32.855 52.330 33.315 52.560 ;
        RECT 36.825 52.290 37.455 52.570 ;
        RECT 36.935 52.250 37.395 52.290 ;
        RECT 38.865 52.250 39.325 52.480 ;
        RECT 44.075 52.300 44.535 52.530 ;
        RECT 48.045 52.260 48.675 52.540 ;
        RECT 48.155 52.220 48.615 52.260 ;
        RECT 50.085 52.220 50.545 52.450 ;
        RECT 55.325 52.280 55.785 52.510 ;
        RECT 59.295 52.240 59.925 52.520 ;
        RECT 59.405 52.200 59.865 52.240 ;
        RECT 61.335 52.200 61.795 52.430 ;
        RECT 66.545 52.270 67.005 52.500 ;
        RECT 70.515 52.230 71.145 52.510 ;
        RECT 70.625 52.190 71.085 52.230 ;
        RECT 72.555 52.190 73.015 52.420 ;
        RECT 77.785 52.260 78.245 52.490 ;
        RECT 81.755 52.220 82.385 52.500 ;
        RECT 81.865 52.180 82.325 52.220 ;
        RECT 83.795 52.180 84.255 52.410 ;
        RECT 89.035 52.270 89.495 52.500 ;
        RECT 93.005 52.230 93.635 52.510 ;
        RECT 93.115 52.190 93.575 52.230 ;
        RECT 95.045 52.190 95.505 52.420 ;
        RECT 100.315 52.260 100.775 52.490 ;
        RECT 104.285 52.220 104.915 52.500 ;
        RECT 104.395 52.180 104.855 52.220 ;
        RECT 106.325 52.180 106.785 52.410 ;
        RECT 111.585 52.260 112.045 52.490 ;
        RECT 115.555 52.220 116.185 52.500 ;
        RECT 115.665 52.180 116.125 52.220 ;
        RECT 117.595 52.180 118.055 52.410 ;
        RECT 122.835 52.260 123.295 52.490 ;
        RECT 126.805 52.220 127.435 52.500 ;
        RECT 126.915 52.180 127.375 52.220 ;
        RECT 128.845 52.180 129.305 52.410 ;
        RECT 21.375 52.010 21.605 52.115 ;
        RECT 21.245 50.290 21.615 52.010 ;
        RECT 22.165 51.890 22.395 52.115 ;
        RECT 25.455 51.980 25.685 52.035 ;
        RECT 21.375 50.115 21.605 50.290 ;
        RECT 22.155 50.210 22.525 51.890 ;
        RECT 22.165 50.115 22.395 50.210 ;
        RECT 21.525 49.670 22.245 49.930 ;
        RECT 19.295 46.650 20.065 47.720 ;
        RECT 21.385 47.490 22.105 47.750 ;
        RECT 21.225 47.200 21.455 47.340 ;
        RECT 21.085 46.430 21.475 47.200 ;
        RECT 22.015 47.190 22.245 47.340 ;
        RECT 22.005 46.450 22.375 47.190 ;
        RECT 25.305 47.010 25.735 51.980 ;
        RECT 26.245 51.970 26.475 52.035 ;
        RECT 27.385 51.970 27.615 52.035 ;
        RECT 26.185 46.970 26.585 51.970 ;
        RECT 27.265 46.970 27.665 51.970 ;
        RECT 28.175 51.940 28.405 52.035 ;
        RECT 32.575 52.020 32.805 52.125 ;
        RECT 28.115 46.970 28.545 51.940 ;
        RECT 32.445 50.300 32.815 52.020 ;
        RECT 33.365 51.900 33.595 52.125 ;
        RECT 36.655 51.990 36.885 52.045 ;
        RECT 32.575 50.125 32.805 50.300 ;
        RECT 33.355 50.220 33.725 51.900 ;
        RECT 33.365 50.125 33.595 50.220 ;
        RECT 32.725 49.680 33.445 49.940 ;
        RECT 25.735 46.600 26.195 46.830 ;
        RECT 27.665 46.710 28.125 46.830 ;
        RECT 27.515 46.600 28.125 46.710 ;
        RECT 30.495 46.660 31.265 47.730 ;
        RECT 32.585 47.500 33.305 47.760 ;
        RECT 32.425 47.210 32.655 47.350 ;
        RECT 21.225 46.340 21.455 46.430 ;
        RECT 22.015 46.340 22.245 46.450 ;
        RECT 27.515 46.430 28.095 46.600 ;
        RECT 32.285 46.440 32.675 47.210 ;
        RECT 33.215 47.200 33.445 47.350 ;
        RECT 33.205 46.460 33.575 47.200 ;
        RECT 36.505 47.020 36.935 51.990 ;
        RECT 37.445 51.980 37.675 52.045 ;
        RECT 38.585 51.980 38.815 52.045 ;
        RECT 37.385 46.980 37.785 51.980 ;
        RECT 38.465 46.980 38.865 51.980 ;
        RECT 39.375 51.950 39.605 52.045 ;
        RECT 43.795 51.990 44.025 52.095 ;
        RECT 39.315 46.980 39.745 51.950 ;
        RECT 43.665 50.270 44.035 51.990 ;
        RECT 44.585 51.870 44.815 52.095 ;
        RECT 47.875 51.960 48.105 52.015 ;
        RECT 43.795 50.095 44.025 50.270 ;
        RECT 44.575 50.190 44.945 51.870 ;
        RECT 44.585 50.095 44.815 50.190 ;
        RECT 43.945 49.650 44.665 49.910 ;
        RECT 36.935 46.610 37.395 46.840 ;
        RECT 38.865 46.720 39.325 46.840 ;
        RECT 38.715 46.610 39.325 46.720 ;
        RECT 41.715 46.630 42.485 47.700 ;
        RECT 43.805 47.470 44.525 47.730 ;
        RECT 43.645 47.180 43.875 47.320 ;
        RECT 32.425 46.350 32.655 46.440 ;
        RECT 33.215 46.350 33.445 46.460 ;
        RECT 38.715 46.440 39.295 46.610 ;
        RECT 43.505 46.410 43.895 47.180 ;
        RECT 44.435 47.170 44.665 47.320 ;
        RECT 44.425 46.430 44.795 47.170 ;
        RECT 47.725 46.990 48.155 51.960 ;
        RECT 48.665 51.950 48.895 52.015 ;
        RECT 49.805 51.950 50.035 52.015 ;
        RECT 48.605 46.950 49.005 51.950 ;
        RECT 49.685 46.950 50.085 51.950 ;
        RECT 50.595 51.920 50.825 52.015 ;
        RECT 55.045 51.970 55.275 52.075 ;
        RECT 50.535 46.950 50.965 51.920 ;
        RECT 54.915 50.250 55.285 51.970 ;
        RECT 55.835 51.850 56.065 52.075 ;
        RECT 59.125 51.940 59.355 51.995 ;
        RECT 55.045 50.075 55.275 50.250 ;
        RECT 55.825 50.170 56.195 51.850 ;
        RECT 55.835 50.075 56.065 50.170 ;
        RECT 55.195 49.630 55.915 49.890 ;
        RECT 48.155 46.580 48.615 46.810 ;
        RECT 50.085 46.690 50.545 46.810 ;
        RECT 49.935 46.580 50.545 46.690 ;
        RECT 52.965 46.610 53.735 47.680 ;
        RECT 55.055 47.450 55.775 47.710 ;
        RECT 54.895 47.160 55.125 47.300 ;
        RECT 43.645 46.320 43.875 46.410 ;
        RECT 44.435 46.320 44.665 46.430 ;
        RECT 49.935 46.410 50.515 46.580 ;
        RECT 54.755 46.390 55.145 47.160 ;
        RECT 55.685 47.150 55.915 47.300 ;
        RECT 55.675 46.410 56.045 47.150 ;
        RECT 58.975 46.970 59.405 51.940 ;
        RECT 59.915 51.930 60.145 51.995 ;
        RECT 61.055 51.930 61.285 51.995 ;
        RECT 59.855 46.930 60.255 51.930 ;
        RECT 60.935 46.930 61.335 51.930 ;
        RECT 61.845 51.900 62.075 51.995 ;
        RECT 66.265 51.960 66.495 52.065 ;
        RECT 61.785 46.930 62.215 51.900 ;
        RECT 66.135 50.240 66.505 51.960 ;
        RECT 67.055 51.840 67.285 52.065 ;
        RECT 70.345 51.930 70.575 51.985 ;
        RECT 66.265 50.065 66.495 50.240 ;
        RECT 67.045 50.160 67.415 51.840 ;
        RECT 67.055 50.065 67.285 50.160 ;
        RECT 66.415 49.620 67.135 49.880 ;
        RECT 59.405 46.560 59.865 46.790 ;
        RECT 61.335 46.670 61.795 46.790 ;
        RECT 61.185 46.560 61.795 46.670 ;
        RECT 64.185 46.600 64.955 47.670 ;
        RECT 66.275 47.440 66.995 47.700 ;
        RECT 66.115 47.150 66.345 47.290 ;
        RECT 54.895 46.300 55.125 46.390 ;
        RECT 55.685 46.300 55.915 46.410 ;
        RECT 61.185 46.390 61.765 46.560 ;
        RECT 65.975 46.380 66.365 47.150 ;
        RECT 66.905 47.140 67.135 47.290 ;
        RECT 66.895 46.400 67.265 47.140 ;
        RECT 70.195 46.960 70.625 51.930 ;
        RECT 71.135 51.920 71.365 51.985 ;
        RECT 72.275 51.920 72.505 51.985 ;
        RECT 71.075 46.920 71.475 51.920 ;
        RECT 72.155 46.920 72.555 51.920 ;
        RECT 73.065 51.890 73.295 51.985 ;
        RECT 77.505 51.950 77.735 52.055 ;
        RECT 73.005 46.920 73.435 51.890 ;
        RECT 77.375 50.230 77.745 51.950 ;
        RECT 78.295 51.830 78.525 52.055 ;
        RECT 81.585 51.920 81.815 51.975 ;
        RECT 77.505 50.055 77.735 50.230 ;
        RECT 78.285 50.150 78.655 51.830 ;
        RECT 78.295 50.055 78.525 50.150 ;
        RECT 77.655 49.610 78.375 49.870 ;
        RECT 70.625 46.550 71.085 46.780 ;
        RECT 72.555 46.660 73.015 46.780 ;
        RECT 72.405 46.550 73.015 46.660 ;
        RECT 75.425 46.590 76.195 47.660 ;
        RECT 77.515 47.430 78.235 47.690 ;
        RECT 77.355 47.140 77.585 47.280 ;
        RECT 66.115 46.290 66.345 46.380 ;
        RECT 66.905 46.290 67.135 46.400 ;
        RECT 72.405 46.380 72.985 46.550 ;
        RECT 77.215 46.370 77.605 47.140 ;
        RECT 78.145 47.130 78.375 47.280 ;
        RECT 78.135 46.390 78.505 47.130 ;
        RECT 81.435 46.950 81.865 51.920 ;
        RECT 82.375 51.910 82.605 51.975 ;
        RECT 83.515 51.910 83.745 51.975 ;
        RECT 82.315 46.910 82.715 51.910 ;
        RECT 83.395 46.910 83.795 51.910 ;
        RECT 84.305 51.880 84.535 51.975 ;
        RECT 88.755 51.960 88.985 52.065 ;
        RECT 84.245 46.910 84.675 51.880 ;
        RECT 88.625 50.240 88.995 51.960 ;
        RECT 89.545 51.840 89.775 52.065 ;
        RECT 92.835 51.930 93.065 51.985 ;
        RECT 88.755 50.065 88.985 50.240 ;
        RECT 89.535 50.160 89.905 51.840 ;
        RECT 89.545 50.065 89.775 50.160 ;
        RECT 88.905 49.620 89.625 49.880 ;
        RECT 81.865 46.540 82.325 46.770 ;
        RECT 83.795 46.650 84.255 46.770 ;
        RECT 83.645 46.540 84.255 46.650 ;
        RECT 86.675 46.600 87.445 47.670 ;
        RECT 88.765 47.440 89.485 47.700 ;
        RECT 88.605 47.150 88.835 47.290 ;
        RECT 77.355 46.280 77.585 46.370 ;
        RECT 78.145 46.280 78.375 46.390 ;
        RECT 83.645 46.370 84.225 46.540 ;
        RECT 88.465 46.380 88.855 47.150 ;
        RECT 89.395 47.140 89.625 47.290 ;
        RECT 89.385 46.400 89.755 47.140 ;
        RECT 92.685 46.960 93.115 51.930 ;
        RECT 93.625 51.920 93.855 51.985 ;
        RECT 94.765 51.920 94.995 51.985 ;
        RECT 93.565 46.920 93.965 51.920 ;
        RECT 94.645 46.920 95.045 51.920 ;
        RECT 95.555 51.890 95.785 51.985 ;
        RECT 100.035 51.950 100.265 52.055 ;
        RECT 95.495 46.920 95.925 51.890 ;
        RECT 99.905 50.230 100.275 51.950 ;
        RECT 100.825 51.830 101.055 52.055 ;
        RECT 104.115 51.920 104.345 51.975 ;
        RECT 100.035 50.055 100.265 50.230 ;
        RECT 100.815 50.150 101.185 51.830 ;
        RECT 100.825 50.055 101.055 50.150 ;
        RECT 100.185 49.610 100.905 49.870 ;
        RECT 93.115 46.550 93.575 46.780 ;
        RECT 95.045 46.660 95.505 46.780 ;
        RECT 94.895 46.550 95.505 46.660 ;
        RECT 97.955 46.590 98.725 47.660 ;
        RECT 100.045 47.430 100.765 47.690 ;
        RECT 99.885 47.140 100.115 47.280 ;
        RECT 88.605 46.290 88.835 46.380 ;
        RECT 89.395 46.290 89.625 46.400 ;
        RECT 94.895 46.380 95.475 46.550 ;
        RECT 99.745 46.370 100.135 47.140 ;
        RECT 100.675 47.130 100.905 47.280 ;
        RECT 100.665 46.390 101.035 47.130 ;
        RECT 103.965 46.950 104.395 51.920 ;
        RECT 104.905 51.910 105.135 51.975 ;
        RECT 106.045 51.910 106.275 51.975 ;
        RECT 104.845 46.910 105.245 51.910 ;
        RECT 105.925 46.910 106.325 51.910 ;
        RECT 106.835 51.880 107.065 51.975 ;
        RECT 111.305 51.950 111.535 52.055 ;
        RECT 106.775 46.910 107.205 51.880 ;
        RECT 111.175 50.230 111.545 51.950 ;
        RECT 112.095 51.830 112.325 52.055 ;
        RECT 115.385 51.920 115.615 51.975 ;
        RECT 111.305 50.055 111.535 50.230 ;
        RECT 112.085 50.150 112.455 51.830 ;
        RECT 112.095 50.055 112.325 50.150 ;
        RECT 111.455 49.610 112.175 49.870 ;
        RECT 104.395 46.540 104.855 46.770 ;
        RECT 106.325 46.650 106.785 46.770 ;
        RECT 106.175 46.540 106.785 46.650 ;
        RECT 109.225 46.590 109.995 47.660 ;
        RECT 111.315 47.430 112.035 47.690 ;
        RECT 111.155 47.140 111.385 47.280 ;
        RECT 99.885 46.280 100.115 46.370 ;
        RECT 100.675 46.280 100.905 46.390 ;
        RECT 106.175 46.370 106.755 46.540 ;
        RECT 111.015 46.370 111.405 47.140 ;
        RECT 111.945 47.130 112.175 47.280 ;
        RECT 111.935 46.390 112.305 47.130 ;
        RECT 115.235 46.950 115.665 51.920 ;
        RECT 116.175 51.910 116.405 51.975 ;
        RECT 117.315 51.910 117.545 51.975 ;
        RECT 116.115 46.910 116.515 51.910 ;
        RECT 117.195 46.910 117.595 51.910 ;
        RECT 118.105 51.880 118.335 51.975 ;
        RECT 122.555 51.950 122.785 52.055 ;
        RECT 118.045 46.910 118.475 51.880 ;
        RECT 122.425 50.230 122.795 51.950 ;
        RECT 123.345 51.830 123.575 52.055 ;
        RECT 126.635 51.920 126.865 51.975 ;
        RECT 122.555 50.055 122.785 50.230 ;
        RECT 123.335 50.150 123.705 51.830 ;
        RECT 123.345 50.055 123.575 50.150 ;
        RECT 122.705 49.610 123.425 49.870 ;
        RECT 115.665 46.540 116.125 46.770 ;
        RECT 117.595 46.650 118.055 46.770 ;
        RECT 117.445 46.540 118.055 46.650 ;
        RECT 120.475 46.590 121.245 47.660 ;
        RECT 122.565 47.430 123.285 47.690 ;
        RECT 122.405 47.140 122.635 47.280 ;
        RECT 111.155 46.280 111.385 46.370 ;
        RECT 111.945 46.280 112.175 46.390 ;
        RECT 117.445 46.370 118.025 46.540 ;
        RECT 122.265 46.370 122.655 47.140 ;
        RECT 123.195 47.130 123.425 47.280 ;
        RECT 123.185 46.390 123.555 47.130 ;
        RECT 126.485 46.950 126.915 51.920 ;
        RECT 127.425 51.910 127.655 51.975 ;
        RECT 128.565 51.910 128.795 51.975 ;
        RECT 127.365 46.910 127.765 51.910 ;
        RECT 128.445 46.910 128.845 51.910 ;
        RECT 129.355 51.880 129.585 51.975 ;
        RECT 129.295 46.910 129.725 51.880 ;
        RECT 126.915 46.540 127.375 46.770 ;
        RECT 128.845 46.650 129.305 46.770 ;
        RECT 128.695 46.540 129.305 46.650 ;
        RECT 122.405 46.280 122.635 46.370 ;
        RECT 123.195 46.280 123.425 46.390 ;
        RECT 128.695 46.370 129.275 46.540 ;
        RECT 21.505 45.950 21.965 46.180 ;
        RECT 32.705 45.960 33.165 46.190 ;
        RECT 43.925 45.930 44.385 46.160 ;
        RECT 55.175 45.910 55.635 46.140 ;
        RECT 66.395 45.900 66.855 46.130 ;
        RECT 77.635 45.890 78.095 46.120 ;
        RECT 88.885 45.900 89.345 46.130 ;
        RECT 100.165 45.890 100.625 46.120 ;
        RECT 111.435 45.890 111.895 46.120 ;
        RECT 122.685 45.890 123.145 46.120 ;
        RECT 29.055 45.020 41.225 45.030 ;
        RECT 17.855 45.005 41.225 45.020 ;
        RECT 15.900 45.000 41.225 45.005 ;
        RECT 15.900 44.980 52.445 45.000 ;
        RECT 15.900 44.970 63.695 44.980 ;
        RECT 15.900 44.960 74.915 44.970 ;
        RECT 85.235 44.960 97.405 44.970 ;
        RECT 15.900 43.880 131.205 44.960 ;
        RECT 15.900 43.870 30.025 43.880 ;
        RECT 15.900 43.855 18.690 43.870 ;
        RECT 15.900 41.620 17.050 43.855 ;
        RECT 40.275 43.850 131.205 43.880 ;
        RECT 51.525 43.830 131.205 43.850 ;
        RECT 62.745 43.820 131.205 43.830 ;
        RECT 73.985 43.810 86.155 43.820 ;
        RECT 96.515 43.810 131.205 43.820 ;
        RECT 29.015 43.330 41.185 43.340 ;
        RECT 17.815 43.310 41.185 43.330 ;
        RECT 142.830 43.320 144.150 43.340 ;
        RECT 17.815 43.290 52.405 43.310 ;
        RECT 140.750 43.300 144.150 43.320 ;
        RECT 17.815 43.280 63.655 43.290 ;
        RECT 119.895 43.280 144.150 43.300 ;
        RECT 17.815 43.270 74.875 43.280 ;
        RECT 85.195 43.270 97.365 43.280 ;
        RECT 108.685 43.270 144.150 43.280 ;
        RECT 17.815 42.180 144.150 43.270 ;
        RECT 18.755 42.150 144.150 42.180 ;
        RECT 18.755 42.120 131.165 42.150 ;
        RECT 18.755 42.090 109.655 42.120 ;
        RECT 18.755 42.080 98.445 42.090 ;
        RECT 41.325 42.070 98.445 42.080 ;
        RECT 142.830 42.070 144.150 42.150 ;
        RECT 41.325 42.060 87.205 42.070 ;
        RECT 75.035 42.050 87.205 42.060 ;
        RECT 15.900 41.540 19.685 41.620 ;
        RECT 142.070 41.610 146.210 41.640 ;
        RECT 119.855 41.590 146.210 41.610 ;
        RECT 108.645 41.550 146.210 41.590 ;
        RECT 15.900 41.520 42.165 41.540 ;
        RECT 97.445 41.530 146.210 41.550 ;
        RECT 15.900 41.510 75.875 41.520 ;
        RECT 86.235 41.510 146.210 41.530 ;
        RECT 15.900 40.500 146.210 41.510 ;
        RECT 15.900 40.480 142.320 40.500 ;
        RECT 15.900 40.470 140.920 40.480 ;
        RECT 18.715 40.460 140.920 40.470 ;
        RECT 142.070 40.460 142.250 40.480 ;
        RECT 18.715 40.440 120.815 40.460 ;
        RECT 18.715 40.400 109.615 40.440 ;
        RECT 18.715 40.390 98.405 40.400 ;
        RECT 41.285 40.380 98.405 40.390 ;
        RECT 41.285 40.370 87.165 40.380 ;
        RECT 74.995 40.360 87.165 40.370 ;
        RECT 26.775 39.230 27.235 39.460 ;
        RECT 38.055 39.230 38.515 39.460 ;
        RECT 49.345 39.210 49.805 39.440 ;
        RECT 60.565 39.210 61.025 39.440 ;
        RECT 71.765 39.210 72.225 39.440 ;
        RECT 83.055 39.200 83.515 39.430 ;
        RECT 94.295 39.220 94.755 39.450 ;
        RECT 105.505 39.240 105.965 39.470 ;
        RECT 116.705 39.280 117.165 39.510 ;
        RECT 127.915 39.300 128.375 39.530 ;
        RECT 20.645 38.810 21.225 38.980 ;
        RECT 26.495 38.960 26.725 39.070 ;
        RECT 27.285 38.980 27.515 39.070 ;
        RECT 20.615 38.700 21.225 38.810 ;
        RECT 20.615 38.580 21.075 38.700 ;
        RECT 22.545 38.580 23.005 38.810 ;
        RECT 20.195 33.470 20.625 38.440 ;
        RECT 20.335 33.375 20.565 33.470 ;
        RECT 21.075 33.440 21.475 38.440 ;
        RECT 22.155 33.440 22.555 38.440 ;
        RECT 21.125 33.375 21.355 33.440 ;
        RECT 22.265 33.375 22.495 33.440 ;
        RECT 23.005 33.430 23.435 38.400 ;
        RECT 26.365 38.220 26.735 38.960 ;
        RECT 26.495 38.070 26.725 38.220 ;
        RECT 27.265 38.210 27.655 38.980 ;
        RECT 31.925 38.810 32.505 38.980 ;
        RECT 37.775 38.960 38.005 39.070 ;
        RECT 38.565 38.980 38.795 39.070 ;
        RECT 27.285 38.070 27.515 38.210 ;
        RECT 26.635 37.660 27.355 37.920 ;
        RECT 28.675 37.690 29.445 38.760 ;
        RECT 31.895 38.700 32.505 38.810 ;
        RECT 31.895 38.580 32.355 38.700 ;
        RECT 33.825 38.580 34.285 38.810 ;
        RECT 26.495 35.480 27.215 35.740 ;
        RECT 26.345 35.200 26.575 35.295 ;
        RECT 26.215 33.520 26.585 35.200 ;
        RECT 27.135 35.120 27.365 35.295 ;
        RECT 23.055 33.375 23.285 33.430 ;
        RECT 26.345 33.295 26.575 33.520 ;
        RECT 27.125 33.400 27.495 35.120 ;
        RECT 31.475 33.470 31.905 38.440 ;
        RECT 27.135 33.295 27.365 33.400 ;
        RECT 31.615 33.375 31.845 33.470 ;
        RECT 32.355 33.440 32.755 38.440 ;
        RECT 33.435 33.440 33.835 38.440 ;
        RECT 32.405 33.375 32.635 33.440 ;
        RECT 33.545 33.375 33.775 33.440 ;
        RECT 34.285 33.430 34.715 38.400 ;
        RECT 37.645 38.220 38.015 38.960 ;
        RECT 37.775 38.070 38.005 38.220 ;
        RECT 38.545 38.210 38.935 38.980 ;
        RECT 43.215 38.790 43.795 38.960 ;
        RECT 49.065 38.940 49.295 39.050 ;
        RECT 49.855 38.960 50.085 39.050 ;
        RECT 38.565 38.070 38.795 38.210 ;
        RECT 37.915 37.660 38.635 37.920 ;
        RECT 39.955 37.690 40.725 38.760 ;
        RECT 43.185 38.680 43.795 38.790 ;
        RECT 43.185 38.560 43.645 38.680 ;
        RECT 45.115 38.560 45.575 38.790 ;
        RECT 37.775 35.480 38.495 35.740 ;
        RECT 37.625 35.200 37.855 35.295 ;
        RECT 37.495 33.520 37.865 35.200 ;
        RECT 38.415 35.120 38.645 35.295 ;
        RECT 34.335 33.375 34.565 33.430 ;
        RECT 37.625 33.295 37.855 33.520 ;
        RECT 38.405 33.400 38.775 35.120 ;
        RECT 42.765 33.450 43.195 38.420 ;
        RECT 38.415 33.295 38.645 33.400 ;
        RECT 42.905 33.355 43.135 33.450 ;
        RECT 43.645 33.420 44.045 38.420 ;
        RECT 44.725 33.420 45.125 38.420 ;
        RECT 43.695 33.355 43.925 33.420 ;
        RECT 44.835 33.355 45.065 33.420 ;
        RECT 45.575 33.410 46.005 38.380 ;
        RECT 48.935 38.200 49.305 38.940 ;
        RECT 49.065 38.050 49.295 38.200 ;
        RECT 49.835 38.190 50.225 38.960 ;
        RECT 54.435 38.790 55.015 38.960 ;
        RECT 60.285 38.940 60.515 39.050 ;
        RECT 61.075 38.960 61.305 39.050 ;
        RECT 49.855 38.050 50.085 38.190 ;
        RECT 49.205 37.640 49.925 37.900 ;
        RECT 51.245 37.670 52.015 38.740 ;
        RECT 54.405 38.680 55.015 38.790 ;
        RECT 54.405 38.560 54.865 38.680 ;
        RECT 56.335 38.560 56.795 38.790 ;
        RECT 49.065 35.460 49.785 35.720 ;
        RECT 48.915 35.180 49.145 35.275 ;
        RECT 48.785 33.500 49.155 35.180 ;
        RECT 49.705 35.100 49.935 35.275 ;
        RECT 45.625 33.355 45.855 33.410 ;
        RECT 48.915 33.275 49.145 33.500 ;
        RECT 49.695 33.380 50.065 35.100 ;
        RECT 53.985 33.450 54.415 38.420 ;
        RECT 49.705 33.275 49.935 33.380 ;
        RECT 54.125 33.355 54.355 33.450 ;
        RECT 54.865 33.420 55.265 38.420 ;
        RECT 55.945 33.420 56.345 38.420 ;
        RECT 54.915 33.355 55.145 33.420 ;
        RECT 56.055 33.355 56.285 33.420 ;
        RECT 56.795 33.410 57.225 38.380 ;
        RECT 60.155 38.200 60.525 38.940 ;
        RECT 60.285 38.050 60.515 38.200 ;
        RECT 61.055 38.190 61.445 38.960 ;
        RECT 65.635 38.790 66.215 38.960 ;
        RECT 71.485 38.940 71.715 39.050 ;
        RECT 72.275 38.960 72.505 39.050 ;
        RECT 61.075 38.050 61.305 38.190 ;
        RECT 60.425 37.640 61.145 37.900 ;
        RECT 62.465 37.670 63.235 38.740 ;
        RECT 65.605 38.680 66.215 38.790 ;
        RECT 65.605 38.560 66.065 38.680 ;
        RECT 67.535 38.560 67.995 38.790 ;
        RECT 60.285 35.460 61.005 35.720 ;
        RECT 60.135 35.180 60.365 35.275 ;
        RECT 60.005 33.500 60.375 35.180 ;
        RECT 60.925 35.100 61.155 35.275 ;
        RECT 56.845 33.355 57.075 33.410 ;
        RECT 60.135 33.275 60.365 33.500 ;
        RECT 60.915 33.380 61.285 35.100 ;
        RECT 65.185 33.450 65.615 38.420 ;
        RECT 60.925 33.275 61.155 33.380 ;
        RECT 65.325 33.355 65.555 33.450 ;
        RECT 66.065 33.420 66.465 38.420 ;
        RECT 67.145 33.420 67.545 38.420 ;
        RECT 66.115 33.355 66.345 33.420 ;
        RECT 67.255 33.355 67.485 33.420 ;
        RECT 67.995 33.410 68.425 38.380 ;
        RECT 71.355 38.200 71.725 38.940 ;
        RECT 71.485 38.050 71.715 38.200 ;
        RECT 72.255 38.190 72.645 38.960 ;
        RECT 76.925 38.780 77.505 38.950 ;
        RECT 82.775 38.930 83.005 39.040 ;
        RECT 83.565 38.950 83.795 39.040 ;
        RECT 72.275 38.050 72.505 38.190 ;
        RECT 71.625 37.640 72.345 37.900 ;
        RECT 73.665 37.670 74.435 38.740 ;
        RECT 76.895 38.670 77.505 38.780 ;
        RECT 76.895 38.550 77.355 38.670 ;
        RECT 78.825 38.550 79.285 38.780 ;
        RECT 71.485 35.460 72.205 35.720 ;
        RECT 71.335 35.180 71.565 35.275 ;
        RECT 71.205 33.500 71.575 35.180 ;
        RECT 72.125 35.100 72.355 35.275 ;
        RECT 68.045 33.355 68.275 33.410 ;
        RECT 71.335 33.275 71.565 33.500 ;
        RECT 72.115 33.380 72.485 35.100 ;
        RECT 76.475 33.440 76.905 38.410 ;
        RECT 72.125 33.275 72.355 33.380 ;
        RECT 76.615 33.345 76.845 33.440 ;
        RECT 77.355 33.410 77.755 38.410 ;
        RECT 78.435 33.410 78.835 38.410 ;
        RECT 77.405 33.345 77.635 33.410 ;
        RECT 78.545 33.345 78.775 33.410 ;
        RECT 79.285 33.400 79.715 38.370 ;
        RECT 82.645 38.190 83.015 38.930 ;
        RECT 82.775 38.040 83.005 38.190 ;
        RECT 83.545 38.180 83.935 38.950 ;
        RECT 88.165 38.800 88.745 38.970 ;
        RECT 94.015 38.950 94.245 39.060 ;
        RECT 94.805 38.970 95.035 39.060 ;
        RECT 83.565 38.040 83.795 38.180 ;
        RECT 82.915 37.630 83.635 37.890 ;
        RECT 84.955 37.660 85.725 38.730 ;
        RECT 88.135 38.690 88.745 38.800 ;
        RECT 88.135 38.570 88.595 38.690 ;
        RECT 90.065 38.570 90.525 38.800 ;
        RECT 82.775 35.450 83.495 35.710 ;
        RECT 82.625 35.170 82.855 35.265 ;
        RECT 82.495 33.490 82.865 35.170 ;
        RECT 83.415 35.090 83.645 35.265 ;
        RECT 79.335 33.345 79.565 33.400 ;
        RECT 82.625 33.265 82.855 33.490 ;
        RECT 83.405 33.370 83.775 35.090 ;
        RECT 87.715 33.460 88.145 38.430 ;
        RECT 83.415 33.265 83.645 33.370 ;
        RECT 87.855 33.365 88.085 33.460 ;
        RECT 88.595 33.430 88.995 38.430 ;
        RECT 89.675 33.430 90.075 38.430 ;
        RECT 88.645 33.365 88.875 33.430 ;
        RECT 89.785 33.365 90.015 33.430 ;
        RECT 90.525 33.420 90.955 38.390 ;
        RECT 93.885 38.210 94.255 38.950 ;
        RECT 94.015 38.060 94.245 38.210 ;
        RECT 94.785 38.200 95.175 38.970 ;
        RECT 99.375 38.820 99.955 38.990 ;
        RECT 105.225 38.970 105.455 39.080 ;
        RECT 106.015 38.990 106.245 39.080 ;
        RECT 94.805 38.060 95.035 38.200 ;
        RECT 94.155 37.650 94.875 37.910 ;
        RECT 96.195 37.680 96.965 38.750 ;
        RECT 99.345 38.710 99.955 38.820 ;
        RECT 99.345 38.590 99.805 38.710 ;
        RECT 101.275 38.590 101.735 38.820 ;
        RECT 94.015 35.470 94.735 35.730 ;
        RECT 93.865 35.190 94.095 35.285 ;
        RECT 93.735 33.510 94.105 35.190 ;
        RECT 94.655 35.110 94.885 35.285 ;
        RECT 90.575 33.365 90.805 33.420 ;
        RECT 93.865 33.285 94.095 33.510 ;
        RECT 94.645 33.390 95.015 35.110 ;
        RECT 98.925 33.480 99.355 38.450 ;
        RECT 94.655 33.285 94.885 33.390 ;
        RECT 99.065 33.385 99.295 33.480 ;
        RECT 99.805 33.450 100.205 38.450 ;
        RECT 100.885 33.450 101.285 38.450 ;
        RECT 99.855 33.385 100.085 33.450 ;
        RECT 100.995 33.385 101.225 33.450 ;
        RECT 101.735 33.440 102.165 38.410 ;
        RECT 105.095 38.230 105.465 38.970 ;
        RECT 105.225 38.080 105.455 38.230 ;
        RECT 105.995 38.220 106.385 38.990 ;
        RECT 110.575 38.860 111.155 39.030 ;
        RECT 116.425 39.010 116.655 39.120 ;
        RECT 117.215 39.030 117.445 39.120 ;
        RECT 106.015 38.080 106.245 38.220 ;
        RECT 105.365 37.670 106.085 37.930 ;
        RECT 107.405 37.700 108.175 38.770 ;
        RECT 110.545 38.750 111.155 38.860 ;
        RECT 110.545 38.630 111.005 38.750 ;
        RECT 112.475 38.630 112.935 38.860 ;
        RECT 105.225 35.490 105.945 35.750 ;
        RECT 105.075 35.210 105.305 35.305 ;
        RECT 104.945 33.530 105.315 35.210 ;
        RECT 105.865 35.130 106.095 35.305 ;
        RECT 101.785 33.385 102.015 33.440 ;
        RECT 105.075 33.305 105.305 33.530 ;
        RECT 105.855 33.410 106.225 35.130 ;
        RECT 110.125 33.520 110.555 38.490 ;
        RECT 110.265 33.425 110.495 33.520 ;
        RECT 111.005 33.490 111.405 38.490 ;
        RECT 112.085 33.490 112.485 38.490 ;
        RECT 111.055 33.425 111.285 33.490 ;
        RECT 112.195 33.425 112.425 33.490 ;
        RECT 112.935 33.480 113.365 38.450 ;
        RECT 116.295 38.270 116.665 39.010 ;
        RECT 116.425 38.120 116.655 38.270 ;
        RECT 117.195 38.260 117.585 39.030 ;
        RECT 121.785 38.880 122.365 39.050 ;
        RECT 127.635 39.030 127.865 39.140 ;
        RECT 128.425 39.050 128.655 39.140 ;
        RECT 117.215 38.120 117.445 38.260 ;
        RECT 116.565 37.710 117.285 37.970 ;
        RECT 118.605 37.740 119.375 38.810 ;
        RECT 121.755 38.770 122.365 38.880 ;
        RECT 121.755 38.650 122.215 38.770 ;
        RECT 123.685 38.650 124.145 38.880 ;
        RECT 116.425 35.530 117.145 35.790 ;
        RECT 116.275 35.250 116.505 35.345 ;
        RECT 116.145 33.570 116.515 35.250 ;
        RECT 117.065 35.170 117.295 35.345 ;
        RECT 112.985 33.425 113.215 33.480 ;
        RECT 105.865 33.305 106.095 33.410 ;
        RECT 116.275 33.345 116.505 33.570 ;
        RECT 117.055 33.450 117.425 35.170 ;
        RECT 121.335 33.540 121.765 38.510 ;
        RECT 117.065 33.345 117.295 33.450 ;
        RECT 121.475 33.445 121.705 33.540 ;
        RECT 122.215 33.510 122.615 38.510 ;
        RECT 123.295 33.510 123.695 38.510 ;
        RECT 122.265 33.445 122.495 33.510 ;
        RECT 123.405 33.445 123.635 33.510 ;
        RECT 124.145 33.500 124.575 38.470 ;
        RECT 127.505 38.290 127.875 39.030 ;
        RECT 127.635 38.140 127.865 38.290 ;
        RECT 128.405 38.280 128.795 39.050 ;
        RECT 128.425 38.140 128.655 38.280 ;
        RECT 127.775 37.730 128.495 37.990 ;
        RECT 129.815 37.760 130.585 38.830 ;
        RECT 142.850 37.630 144.170 38.900 ;
        RECT 127.635 35.550 128.355 35.810 ;
        RECT 127.485 35.270 127.715 35.365 ;
        RECT 127.355 33.590 127.725 35.270 ;
        RECT 128.275 35.190 128.505 35.365 ;
        RECT 124.195 33.445 124.425 33.500 ;
        RECT 127.485 33.365 127.715 33.590 ;
        RECT 128.265 33.470 128.635 35.190 ;
        RECT 128.275 33.365 128.505 33.470 ;
        RECT 20.615 32.940 21.075 33.170 ;
        RECT 22.545 33.130 23.005 33.170 ;
        RECT 22.485 32.850 23.115 33.130 ;
        RECT 26.625 32.860 27.085 33.090 ;
        RECT 31.895 32.940 32.355 33.170 ;
        RECT 33.825 33.130 34.285 33.170 ;
        RECT 33.765 32.850 34.395 33.130 ;
        RECT 37.905 32.860 38.365 33.090 ;
        RECT 43.185 32.920 43.645 33.150 ;
        RECT 45.115 33.110 45.575 33.150 ;
        RECT 45.055 32.830 45.685 33.110 ;
        RECT 49.195 32.840 49.655 33.070 ;
        RECT 54.405 32.920 54.865 33.150 ;
        RECT 56.335 33.110 56.795 33.150 ;
        RECT 56.275 32.830 56.905 33.110 ;
        RECT 60.415 32.840 60.875 33.070 ;
        RECT 65.605 32.920 66.065 33.150 ;
        RECT 67.535 33.110 67.995 33.150 ;
        RECT 67.475 32.830 68.105 33.110 ;
        RECT 71.615 32.840 72.075 33.070 ;
        RECT 76.895 32.910 77.355 33.140 ;
        RECT 78.825 33.100 79.285 33.140 ;
        RECT 78.765 32.820 79.395 33.100 ;
        RECT 82.905 32.830 83.365 33.060 ;
        RECT 88.135 32.930 88.595 33.160 ;
        RECT 90.065 33.120 90.525 33.160 ;
        RECT 90.005 32.840 90.635 33.120 ;
        RECT 94.145 32.850 94.605 33.080 ;
        RECT 99.345 32.950 99.805 33.180 ;
        RECT 101.275 33.140 101.735 33.180 ;
        RECT 101.215 32.860 101.845 33.140 ;
        RECT 105.355 32.870 105.815 33.100 ;
        RECT 110.545 32.990 111.005 33.220 ;
        RECT 112.475 33.180 112.935 33.220 ;
        RECT 112.415 32.900 113.045 33.180 ;
        RECT 116.555 32.910 117.015 33.140 ;
        RECT 121.755 33.010 122.215 33.240 ;
        RECT 123.685 33.200 124.145 33.240 ;
        RECT 123.625 32.920 124.255 33.200 ;
        RECT 127.765 32.930 128.225 33.160 ;
        RECT 23.185 30.880 27.925 31.180 ;
        RECT 34.465 30.880 39.205 31.180 ;
        RECT 45.755 30.860 50.495 31.160 ;
        RECT 56.975 30.860 61.715 31.160 ;
        RECT 68.175 30.860 72.915 31.160 ;
        RECT 79.465 30.850 84.205 31.150 ;
        RECT 90.705 30.870 95.445 31.170 ;
        RECT 101.915 30.890 106.655 31.190 ;
        RECT 113.115 30.930 117.855 31.230 ;
        RECT 124.325 30.950 129.065 31.250 ;
        RECT 19.485 20.270 19.905 30.160 ;
        RECT 19.585 20.090 19.815 20.270 ;
        RECT 20.805 20.260 21.175 30.210 ;
        RECT 20.875 20.090 21.105 20.260 ;
        RECT 21.935 20.220 22.305 30.170 ;
        RECT 27.255 20.270 27.615 30.190 ;
        RECT 30.765 20.270 31.185 30.160 ;
        RECT 22.015 20.090 22.245 20.220 ;
        RECT 27.305 20.090 27.535 20.270 ;
        RECT 30.865 20.090 31.095 20.270 ;
        RECT 32.085 20.260 32.455 30.210 ;
        RECT 32.155 20.090 32.385 20.260 ;
        RECT 33.215 20.220 33.585 30.170 ;
        RECT 38.535 20.270 38.895 30.190 ;
        RECT 33.295 20.090 33.525 20.220 ;
        RECT 38.585 20.090 38.815 20.270 ;
        RECT 42.055 20.250 42.475 30.140 ;
        RECT 42.155 20.070 42.385 20.250 ;
        RECT 43.375 20.240 43.745 30.190 ;
        RECT 43.445 20.070 43.675 20.240 ;
        RECT 44.505 20.200 44.875 30.150 ;
        RECT 49.825 20.250 50.185 30.170 ;
        RECT 53.275 20.250 53.695 30.140 ;
        RECT 44.585 20.070 44.815 20.200 ;
        RECT 49.875 20.070 50.105 20.250 ;
        RECT 53.375 20.070 53.605 20.250 ;
        RECT 54.595 20.240 54.965 30.190 ;
        RECT 54.665 20.070 54.895 20.240 ;
        RECT 55.725 20.200 56.095 30.150 ;
        RECT 61.045 20.250 61.405 30.170 ;
        RECT 64.475 20.250 64.895 30.140 ;
        RECT 55.805 20.070 56.035 20.200 ;
        RECT 61.095 20.070 61.325 20.250 ;
        RECT 64.575 20.070 64.805 20.250 ;
        RECT 65.795 20.240 66.165 30.190 ;
        RECT 65.865 20.070 66.095 20.240 ;
        RECT 66.925 20.200 67.295 30.150 ;
        RECT 72.245 20.250 72.605 30.170 ;
        RECT 67.005 20.070 67.235 20.200 ;
        RECT 72.295 20.070 72.525 20.250 ;
        RECT 75.765 20.240 76.185 30.130 ;
        RECT 75.865 20.060 76.095 20.240 ;
        RECT 77.085 20.230 77.455 30.180 ;
        RECT 77.155 20.060 77.385 20.230 ;
        RECT 78.215 20.190 78.585 30.140 ;
        RECT 83.535 20.240 83.895 30.160 ;
        RECT 87.005 20.260 87.425 30.150 ;
        RECT 78.295 20.060 78.525 20.190 ;
        RECT 83.585 20.060 83.815 20.240 ;
        RECT 87.105 20.080 87.335 20.260 ;
        RECT 88.325 20.250 88.695 30.200 ;
        RECT 88.395 20.080 88.625 20.250 ;
        RECT 89.455 20.210 89.825 30.160 ;
        RECT 94.775 20.260 95.135 30.180 ;
        RECT 98.215 20.280 98.635 30.170 ;
        RECT 89.535 20.080 89.765 20.210 ;
        RECT 94.825 20.080 95.055 20.260 ;
        RECT 98.315 20.100 98.545 20.280 ;
        RECT 99.535 20.270 99.905 30.220 ;
        RECT 99.605 20.100 99.835 20.270 ;
        RECT 100.665 20.230 101.035 30.180 ;
        RECT 105.985 20.280 106.345 30.200 ;
        RECT 109.415 20.320 109.835 30.210 ;
        RECT 100.745 20.100 100.975 20.230 ;
        RECT 106.035 20.100 106.265 20.280 ;
        RECT 109.515 20.140 109.745 20.320 ;
        RECT 110.735 20.310 111.105 30.260 ;
        RECT 110.805 20.140 111.035 20.310 ;
        RECT 111.865 20.270 112.235 30.220 ;
        RECT 117.185 20.320 117.545 30.240 ;
        RECT 120.625 20.340 121.045 30.230 ;
        RECT 111.945 20.140 112.175 20.270 ;
        RECT 117.235 20.140 117.465 20.320 ;
        RECT 120.725 20.160 120.955 20.340 ;
        RECT 121.945 20.330 122.315 30.280 ;
        RECT 122.015 20.160 122.245 20.330 ;
        RECT 123.075 20.290 123.445 30.240 ;
        RECT 128.395 20.340 128.755 30.260 ;
        RECT 123.155 20.160 123.385 20.290 ;
        RECT 128.445 20.160 128.675 20.340 ;
        RECT 132.345 20.170 132.755 30.180 ;
        RECT 137.735 30.120 137.965 30.130 ;
        RECT 132.445 20.130 132.675 20.170 ;
        RECT 137.665 20.080 138.055 30.120 ;
        RECT 19.775 19.610 20.925 19.920 ;
        RECT 22.185 19.620 27.335 19.900 ;
        RECT 31.055 19.610 32.205 19.920 ;
        RECT 33.465 19.620 38.615 19.900 ;
        RECT 42.345 19.590 43.495 19.900 ;
        RECT 44.755 19.600 49.905 19.880 ;
        RECT 53.565 19.590 54.715 19.900 ;
        RECT 55.975 19.600 61.125 19.880 ;
        RECT 64.765 19.590 65.915 19.900 ;
        RECT 67.175 19.600 72.325 19.880 ;
        RECT 76.055 19.580 77.205 19.890 ;
        RECT 78.465 19.590 83.615 19.870 ;
        RECT 87.295 19.600 88.445 19.910 ;
        RECT 89.705 19.610 94.855 19.890 ;
        RECT 98.505 19.620 99.655 19.930 ;
        RECT 100.915 19.630 106.065 19.910 ;
        RECT 109.705 19.660 110.855 19.970 ;
        RECT 112.115 19.670 117.265 19.950 ;
        RECT 120.915 19.680 122.065 19.990 ;
        RECT 123.325 19.690 128.475 19.970 ;
        RECT 132.635 19.640 138.025 19.930 ;
        RECT 142.940 19.110 144.080 37.630 ;
        RECT 13.940 18.460 17.635 18.530 ;
        RECT 117.755 18.510 131.425 18.530 ;
        RECT 106.545 18.470 131.425 18.510 ;
        RECT 13.940 18.440 41.565 18.460 ;
        RECT 95.345 18.450 131.425 18.470 ;
        RECT 13.940 18.430 75.275 18.440 ;
        RECT 84.135 18.430 131.425 18.450 ;
        RECT 13.940 17.380 131.425 18.430 ;
        RECT 142.890 17.990 144.140 19.110 ;
        RECT 145.070 18.880 146.210 40.500 ;
        RECT 145.030 17.960 146.250 18.880 ;
        RECT 13.950 17.370 15.100 17.380 ;
        RECT 16.615 17.360 120.215 17.380 ;
        RECT 16.615 17.320 109.015 17.360 ;
        RECT 16.615 17.310 97.805 17.320 ;
        RECT 39.185 17.300 97.805 17.310 ;
        RECT 39.185 17.290 86.565 17.300 ;
        RECT 72.895 17.280 86.565 17.290 ;
        RECT 117.765 16.950 140.620 16.960 ;
        RECT 142.040 16.950 148.010 16.980 ;
        RECT 117.765 16.940 148.010 16.950 ;
        RECT 106.555 16.900 148.010 16.940 ;
        RECT 16.625 16.870 41.575 16.890 ;
        RECT 95.355 16.880 148.010 16.900 ;
        RECT 16.625 16.860 75.285 16.870 ;
        RECT 84.145 16.860 148.010 16.880 ;
        RECT 16.625 15.840 148.010 16.860 ;
        RECT 16.625 15.820 142.660 15.840 ;
        RECT 16.625 15.810 140.620 15.820 ;
        RECT 142.040 15.810 142.660 15.820 ;
        RECT 16.625 15.790 120.225 15.810 ;
        RECT 16.625 15.750 109.025 15.790 ;
        RECT 16.625 15.740 97.815 15.750 ;
        RECT 39.195 15.730 97.815 15.740 ;
        RECT 39.195 15.720 86.575 15.730 ;
        RECT 72.905 15.710 86.575 15.720 ;
        RECT 131.215 15.460 132.585 15.470 ;
        RECT 12.290 15.390 17.625 15.450 ;
        RECT 117.795 15.440 132.785 15.460 ;
        RECT 106.585 15.400 132.785 15.440 ;
        RECT 12.290 15.370 41.585 15.390 ;
        RECT 95.385 15.380 132.785 15.400 ;
        RECT 12.290 15.360 75.295 15.370 ;
        RECT 84.175 15.360 132.785 15.380 ;
        RECT 12.290 14.320 132.785 15.360 ;
        RECT 142.905 15.040 144.045 15.050 ;
        RECT 12.290 14.310 131.445 14.320 ;
        RECT 12.290 14.300 120.235 14.310 ;
        RECT 12.320 14.280 13.470 14.300 ;
        RECT 16.655 14.290 120.235 14.300 ;
        RECT 16.655 14.250 109.035 14.290 ;
        RECT 16.655 14.240 97.825 14.250 ;
        RECT 39.225 14.230 97.825 14.240 ;
        RECT 39.225 14.220 86.585 14.230 ;
        RECT 72.935 14.210 86.585 14.220 ;
        RECT 142.850 13.920 144.100 15.040 ;
        RECT 145.020 14.870 146.160 14.980 ;
        RECT 144.980 13.950 146.200 14.870 ;
        RECT 16.965 13.800 17.435 13.810 ;
        RECT 10.800 13.780 17.435 13.800 ;
        RECT 10.800 13.720 17.555 13.780 ;
        RECT 117.845 13.770 131.445 13.790 ;
        RECT 106.635 13.730 131.445 13.770 ;
        RECT 10.800 13.700 41.585 13.720 ;
        RECT 95.435 13.710 131.445 13.730 ;
        RECT 10.800 13.690 75.295 13.700 ;
        RECT 84.225 13.690 131.445 13.710 ;
        RECT 10.800 12.650 131.445 13.690 ;
        RECT 16.705 12.640 131.445 12.650 ;
        RECT 16.705 12.620 120.235 12.640 ;
        RECT 16.705 12.580 109.035 12.620 ;
        RECT 16.705 12.570 97.825 12.580 ;
        RECT 39.275 12.560 97.825 12.570 ;
        RECT 39.275 12.550 86.585 12.560 ;
        RECT 72.985 12.540 86.585 12.550 ;
        RECT 128.755 12.240 130.465 12.250 ;
        RECT 117.545 12.220 119.255 12.230 ;
        RECT 106.345 12.180 108.055 12.190 ;
        RECT 27.615 12.170 29.325 12.180 ;
        RECT 38.895 12.170 40.605 12.180 ;
        RECT 25.675 11.030 29.325 12.170 ;
        RECT 36.955 11.030 40.605 12.170 ;
        RECT 95.135 12.160 96.845 12.170 ;
        RECT 50.185 12.150 51.895 12.160 ;
        RECT 61.405 12.150 63.115 12.160 ;
        RECT 72.605 12.150 74.315 12.160 ;
        RECT 25.675 11.020 27.625 11.030 ;
        RECT 36.955 11.020 38.905 11.030 ;
        RECT 48.245 11.010 51.895 12.150 ;
        RECT 59.465 11.010 63.115 12.150 ;
        RECT 70.665 11.010 74.315 12.150 ;
        RECT 83.895 12.140 85.605 12.150 ;
        RECT 48.245 11.000 50.195 11.010 ;
        RECT 59.465 11.000 61.415 11.010 ;
        RECT 70.665 11.000 72.615 11.010 ;
        RECT 81.955 11.000 85.605 12.140 ;
        RECT 93.195 11.020 96.845 12.160 ;
        RECT 104.405 11.040 108.055 12.180 ;
        RECT 115.605 11.080 119.255 12.220 ;
        RECT 126.815 11.100 130.465 12.240 ;
        RECT 126.815 11.090 128.765 11.100 ;
        RECT 115.605 11.070 117.555 11.080 ;
        RECT 104.405 11.030 106.355 11.040 ;
        RECT 93.195 11.010 95.145 11.020 ;
        RECT 81.955 10.990 83.905 11.000 ;
        RECT 142.905 8.580 144.045 13.920 ;
        RECT 74.420 7.440 144.045 8.580 ;
        RECT 74.420 1.410 75.560 7.440 ;
        RECT 145.020 6.630 146.160 13.950 ;
        RECT 93.650 5.490 146.160 6.630 ;
        RECT 93.650 1.480 94.790 5.490 ;
        RECT 146.870 4.560 148.010 15.840 ;
        RECT 113.130 3.420 148.010 4.560 ;
        RECT 113.130 1.610 114.270 3.420 ;
        RECT 149.460 2.770 150.600 64.660 ;
        RECT 131.940 1.880 150.600 2.770 ;
        RECT 131.800 1.630 150.600 1.880 ;
        RECT 74.290 0.160 75.680 1.410 ;
        RECT 93.500 0.230 94.890 1.480 ;
        RECT 112.900 0.360 114.290 1.610 ;
        RECT 131.800 1.380 133.490 1.630 ;
        RECT 151.730 1.420 152.870 66.900 ;
        RECT 131.800 0.430 133.540 1.380 ;
        RECT 113.130 0.330 114.270 0.360 ;
        RECT 151.600 0.300 152.970 1.420 ;
        RECT 93.650 0.150 94.790 0.230 ;
      LAYER met2 ;
        RECT 135.390 223.830 136.740 225.230 ;
        RECT 138.180 223.760 139.530 225.160 ;
        RECT 143.230 223.790 144.580 225.190 ;
        RECT 46.880 211.105 48.760 211.475 ;
        RECT 76.880 211.105 78.760 211.475 ;
        RECT 106.880 211.105 108.760 211.475 ;
        RECT 31.880 208.385 33.760 208.755 ;
        RECT 61.880 208.385 63.760 208.755 ;
        RECT 91.880 208.385 93.760 208.755 ;
        RECT 121.880 208.385 123.760 208.755 ;
        RECT 46.880 205.665 48.760 206.035 ;
        RECT 76.880 205.665 78.760 206.035 ;
        RECT 106.880 205.665 108.760 206.035 ;
        RECT 31.880 202.945 33.760 203.315 ;
        RECT 61.880 202.945 63.760 203.315 ;
        RECT 91.880 202.945 93.760 203.315 ;
        RECT 121.880 202.945 123.760 203.315 ;
        RECT 72.720 201.780 72.980 202.100 ;
        RECT 72.260 201.440 72.520 201.760 ;
        RECT 64.900 200.760 65.160 201.080 ;
        RECT 46.880 200.225 48.760 200.595 ;
        RECT 64.960 199.720 65.100 200.760 ;
        RECT 52.480 199.400 52.740 199.720 ;
        RECT 64.900 199.400 65.160 199.720 ;
        RECT 71.340 199.400 71.600 199.720 ;
        RECT 46.040 198.720 46.300 199.040 ;
        RECT 49.260 198.720 49.520 199.040 ;
        RECT 31.880 197.505 33.760 197.875 ;
        RECT 31.320 196.000 31.580 196.320 ;
        RECT 29.480 193.960 29.740 194.280 ;
        RECT 28.100 193.280 28.360 193.600 ;
        RECT 28.160 188.500 28.300 193.280 ;
        RECT 29.540 191.560 29.680 193.960 ;
        RECT 29.480 191.240 29.740 191.560 ;
        RECT 31.380 190.880 31.520 196.000 ;
        RECT 34.540 195.320 34.800 195.640 ;
        RECT 42.820 195.320 43.080 195.640 ;
        RECT 43.740 195.320 44.000 195.640 ;
        RECT 34.600 194.280 34.740 195.320 ;
        RECT 42.880 194.280 43.020 195.320 ;
        RECT 34.540 193.960 34.800 194.280 ;
        RECT 42.820 193.960 43.080 194.280 ;
        RECT 37.760 192.600 38.020 192.920 ;
        RECT 40.060 192.600 40.320 192.920 ;
        RECT 31.880 192.065 33.760 192.435 ;
        RECT 31.320 190.560 31.580 190.880 ;
        RECT 28.100 188.180 28.360 188.500 ;
        RECT 28.160 183.060 28.300 188.180 ;
        RECT 29.480 187.160 29.740 187.480 ;
        RECT 29.540 186.120 29.680 187.160 ;
        RECT 29.480 185.800 29.740 186.120 ;
        RECT 31.380 185.440 31.520 190.560 ;
        RECT 37.820 190.540 37.960 192.600 ;
        RECT 37.760 190.220 38.020 190.540 ;
        RECT 40.120 190.200 40.260 192.600 ;
        RECT 43.280 190.900 43.540 191.220 ;
        RECT 32.240 189.880 32.500 190.200 ;
        RECT 36.840 189.880 37.100 190.200 ;
        RECT 40.060 189.880 40.320 190.200 ;
        RECT 32.300 188.840 32.440 189.880 ;
        RECT 32.240 188.520 32.500 188.840 ;
        RECT 36.900 188.160 37.040 189.880 ;
        RECT 36.840 187.840 37.100 188.160 ;
        RECT 31.880 186.625 33.760 186.995 ;
        RECT 31.320 185.120 31.580 185.440 ;
        RECT 35.920 185.120 36.180 185.440 ;
        RECT 31.780 184.440 32.040 184.760 ;
        RECT 31.840 183.400 31.980 184.440 ;
        RECT 31.780 183.080 32.040 183.400 ;
        RECT 28.100 182.740 28.360 183.060 ;
        RECT 29.480 182.400 29.740 182.720 ;
        RECT 29.540 180.680 29.680 182.400 ;
        RECT 31.880 181.185 33.760 181.555 ;
        RECT 29.480 180.360 29.740 180.680 ;
        RECT 31.880 175.745 33.760 176.115 ;
        RECT 26.260 174.580 26.520 174.900 ;
        RECT 24.880 174.240 25.140 174.560 ;
        RECT 24.420 173.900 24.680 174.220 ;
        RECT 24.480 172.860 24.620 173.900 ;
        RECT 24.420 172.540 24.680 172.860 ;
        RECT 24.940 169.800 25.080 174.240 ;
        RECT 26.320 170.140 26.460 174.580 ;
        RECT 29.940 173.560 30.200 173.880 ;
        RECT 26.720 170.840 26.980 171.160 ;
        RECT 26.260 169.820 26.520 170.140 ;
        RECT 24.880 169.480 25.140 169.800 ;
        RECT 23.040 168.800 23.300 169.120 ;
        RECT 23.100 167.420 23.240 168.800 ;
        RECT 23.040 167.100 23.300 167.420 ;
        RECT 26.780 167.080 26.920 170.840 ;
        RECT 26.720 166.760 26.980 167.080 ;
        RECT 30.000 166.400 30.140 173.560 ;
        RECT 34.540 172.200 34.800 172.520 ;
        RECT 30.860 170.840 31.120 171.160 ;
        RECT 29.940 166.080 30.200 166.400 ;
        RECT 30.400 166.080 30.660 166.400 ;
        RECT 29.480 163.360 29.740 163.680 ;
        RECT 25.800 162.680 26.060 163.000 ;
        RECT 28.100 162.680 28.360 163.000 ;
        RECT 25.860 161.640 26.000 162.680 ;
        RECT 28.160 161.980 28.300 162.680 ;
        RECT 28.100 161.660 28.360 161.980 ;
        RECT 25.800 161.320 26.060 161.640 ;
        RECT 28.160 160.140 28.300 161.660 ;
        RECT 29.540 160.280 29.680 163.360 ;
        RECT 30.000 163.340 30.140 166.080 ;
        RECT 30.460 164.020 30.600 166.080 ;
        RECT 30.920 164.020 31.060 170.840 ;
        RECT 31.880 170.305 33.760 170.675 ;
        RECT 33.610 169.285 33.890 169.655 ;
        RECT 33.680 169.120 33.820 169.285 ;
        RECT 33.620 168.800 33.880 169.120 ;
        RECT 34.080 168.460 34.340 168.780 ;
        RECT 31.320 165.400 31.580 165.720 ;
        RECT 30.400 163.700 30.660 164.020 ;
        RECT 30.860 163.700 31.120 164.020 ;
        RECT 29.940 163.020 30.200 163.340 ;
        RECT 28.160 160.000 28.760 160.140 ;
        RECT 26.720 157.920 26.980 158.240 ;
        RECT 26.260 157.240 26.520 157.560 ;
        RECT 26.320 156.200 26.460 157.240 ;
        RECT 26.260 155.880 26.520 156.200 ;
        RECT 26.780 152.540 26.920 157.920 ;
        RECT 28.100 157.240 28.360 157.560 ;
        RECT 28.160 156.540 28.300 157.240 ;
        RECT 28.100 156.220 28.360 156.540 ;
        RECT 28.620 152.800 28.760 160.000 ;
        RECT 29.480 159.960 29.740 160.280 ;
        RECT 29.540 158.920 29.680 159.960 ;
        RECT 29.480 158.600 29.740 158.920 ;
        RECT 30.460 157.900 30.600 163.700 ;
        RECT 31.380 163.680 31.520 165.400 ;
        RECT 31.880 164.865 33.760 165.235 ;
        RECT 34.140 164.700 34.280 168.460 ;
        RECT 34.080 164.380 34.340 164.700 ;
        RECT 34.600 164.360 34.740 172.200 ;
        RECT 35.460 171.520 35.720 171.840 ;
        RECT 35.520 169.800 35.660 171.520 ;
        RECT 35.980 171.500 36.120 185.120 ;
        RECT 36.900 184.760 37.040 187.840 ;
        RECT 37.300 184.780 37.560 185.100 ;
        RECT 36.840 184.440 37.100 184.760 ;
        RECT 37.360 182.040 37.500 184.780 ;
        RECT 38.680 184.440 38.940 184.760 ;
        RECT 37.300 181.720 37.560 182.040 ;
        RECT 37.760 174.920 38.020 175.240 ;
        RECT 36.380 173.900 36.640 174.220 ;
        RECT 35.920 171.180 36.180 171.500 ;
        RECT 35.460 169.480 35.720 169.800 ;
        RECT 35.000 169.140 35.260 169.460 ;
        RECT 35.060 166.740 35.200 169.140 ;
        RECT 35.000 166.420 35.260 166.740 ;
        RECT 35.000 165.740 35.260 166.060 ;
        RECT 34.540 164.040 34.800 164.360 ;
        RECT 35.060 164.020 35.200 165.740 ;
        RECT 35.000 163.700 35.260 164.020 ;
        RECT 31.320 163.360 31.580 163.680 ;
        RECT 33.620 162.680 33.880 163.000 ;
        RECT 33.680 161.300 33.820 162.680 ;
        RECT 33.620 160.980 33.880 161.300 ;
        RECT 35.520 160.960 35.660 169.480 ;
        RECT 35.920 166.760 36.180 167.080 ;
        RECT 35.980 164.360 36.120 166.760 ;
        RECT 35.920 164.040 36.180 164.360 ;
        RECT 35.920 163.360 36.180 163.680 ;
        RECT 31.320 160.640 31.580 160.960 ;
        RECT 35.460 160.640 35.720 160.960 ;
        RECT 30.400 157.580 30.660 157.900 ;
        RECT 29.480 157.240 29.740 157.560 ;
        RECT 26.320 152.400 26.920 152.540 ;
        RECT 28.560 152.480 28.820 152.800 ;
        RECT 25.800 150.440 26.060 150.760 ;
        RECT 25.860 148.380 26.000 150.440 ;
        RECT 25.800 148.060 26.060 148.380 ;
        RECT 26.320 147.360 26.460 152.400 ;
        RECT 26.720 151.800 26.980 152.120 ;
        RECT 26.780 150.080 26.920 151.800 ;
        RECT 28.620 150.330 28.760 152.480 ;
        RECT 29.540 152.460 29.680 157.240 ;
        RECT 30.460 153.140 30.600 157.580 ;
        RECT 31.380 155.520 31.520 160.640 ;
        RECT 35.460 159.960 35.720 160.280 ;
        RECT 31.880 159.425 33.760 159.795 ;
        RECT 35.520 157.900 35.660 159.960 ;
        RECT 35.460 157.580 35.720 157.900 ;
        RECT 33.620 157.240 33.880 157.560 ;
        RECT 33.680 155.860 33.820 157.240 ;
        RECT 33.620 155.540 33.880 155.860 ;
        RECT 35.980 155.520 36.120 163.360 ;
        RECT 31.320 155.200 31.580 155.520 ;
        RECT 35.920 155.200 36.180 155.520 ;
        RECT 31.880 153.985 33.760 154.355 ;
        RECT 30.400 152.820 30.660 153.140 ;
        RECT 32.240 152.820 32.500 153.140 ;
        RECT 29.480 152.140 29.740 152.460 ;
        RECT 29.540 151.100 29.680 152.140 ;
        RECT 29.480 150.780 29.740 151.100 ;
        RECT 29.020 150.330 29.280 150.420 ;
        RECT 28.620 150.190 29.280 150.330 ;
        RECT 29.020 150.100 29.280 150.190 ;
        RECT 32.300 150.080 32.440 152.820 ;
        RECT 33.160 151.800 33.420 152.120 ;
        RECT 33.220 150.080 33.360 151.800 ;
        RECT 35.920 150.100 36.180 150.420 ;
        RECT 26.720 149.760 26.980 150.080 ;
        RECT 32.240 149.760 32.500 150.080 ;
        RECT 33.160 149.760 33.420 150.080 ;
        RECT 31.320 149.420 31.580 149.740 ;
        RECT 31.380 148.380 31.520 149.420 ;
        RECT 34.080 149.080 34.340 149.400 ;
        RECT 31.880 148.545 33.760 148.915 ;
        RECT 31.320 148.060 31.580 148.380 ;
        RECT 34.140 147.700 34.280 149.080 ;
        RECT 35.980 147.700 36.120 150.100 ;
        RECT 34.080 147.380 34.340 147.700 ;
        RECT 35.920 147.380 36.180 147.700 ;
        RECT 26.260 147.040 26.520 147.360 ;
        RECT 26.320 144.980 26.460 147.040 ;
        RECT 30.400 146.700 30.660 147.020 ;
        RECT 30.460 145.660 30.600 146.700 ;
        RECT 30.400 145.340 30.660 145.660 ;
        RECT 26.260 144.660 26.520 144.980 ;
        RECT 30.860 143.980 31.120 144.300 ;
        RECT 27.640 139.560 27.900 139.880 ;
        RECT 27.700 137.500 27.840 139.560 ;
        RECT 29.480 138.200 29.740 138.520 ;
        RECT 27.640 137.180 27.900 137.500 ;
        RECT 29.020 137.180 29.280 137.500 ;
        RECT 27.640 136.160 27.900 136.480 ;
        RECT 26.720 134.120 26.980 134.440 ;
        RECT 26.780 132.060 26.920 134.120 ;
        RECT 26.720 131.740 26.980 132.060 ;
        RECT 26.720 130.950 26.980 131.040 ;
        RECT 27.700 130.950 27.840 136.160 ;
        RECT 29.080 134.780 29.220 137.180 ;
        RECT 29.540 136.480 29.680 138.200 ;
        RECT 29.940 136.840 30.200 137.160 ;
        RECT 29.480 136.160 29.740 136.480 ;
        RECT 29.020 134.460 29.280 134.780 ;
        RECT 29.080 131.040 29.220 134.460 ;
        RECT 29.540 131.380 29.680 136.160 ;
        RECT 29.480 131.060 29.740 131.380 ;
        RECT 26.720 130.810 27.840 130.950 ;
        RECT 26.720 130.720 26.980 130.810 ;
        RECT 29.020 130.720 29.280 131.040 ;
        RECT 26.780 125.940 26.920 130.720 ;
        RECT 29.080 125.940 29.220 130.720 ;
        RECT 30.000 130.700 30.140 136.840 ;
        RECT 29.940 130.380 30.200 130.700 ;
        RECT 29.480 128.000 29.740 128.320 ;
        RECT 26.720 125.620 26.980 125.940 ;
        RECT 29.020 125.620 29.280 125.940 ;
        RECT 29.540 124.920 29.680 128.000 ;
        RECT 30.000 127.980 30.140 130.380 ;
        RECT 30.400 128.340 30.660 128.660 ;
        RECT 30.460 127.980 30.600 128.340 ;
        RECT 29.940 127.660 30.200 127.980 ;
        RECT 30.400 127.660 30.660 127.980 ;
        RECT 30.000 126.620 30.140 127.660 ;
        RECT 29.940 126.300 30.200 126.620 ;
        RECT 23.500 124.600 23.760 124.920 ;
        RECT 25.340 124.600 25.600 124.920 ;
        RECT 27.180 124.600 27.440 124.920 ;
        RECT 29.480 124.600 29.740 124.920 ;
        RECT 23.560 123.560 23.700 124.600 ;
        RECT 23.500 123.240 23.760 123.560 ;
        RECT 25.400 119.820 25.540 124.600 ;
        RECT 27.240 122.880 27.380 124.600 ;
        RECT 29.540 123.900 29.680 124.600 ;
        RECT 30.460 123.900 30.600 127.660 ;
        RECT 29.480 123.580 29.740 123.900 ;
        RECT 30.400 123.580 30.660 123.900 ;
        RECT 27.180 122.560 27.440 122.880 ;
        RECT 30.460 121.180 30.600 123.580 ;
        RECT 30.400 120.860 30.660 121.180 ;
        RECT 25.340 119.500 25.600 119.820 ;
        RECT 25.800 114.060 26.060 114.380 ;
        RECT 25.860 113.020 26.000 114.060 ;
        RECT 27.180 113.720 27.440 114.040 ;
        RECT 27.640 113.720 27.900 114.040 ;
        RECT 25.800 112.700 26.060 113.020 ;
        RECT 24.420 111.680 24.680 112.000 ;
        RECT 24.480 107.240 24.620 111.680 ;
        RECT 24.420 106.920 24.680 107.240 ;
        RECT 21.660 105.560 21.920 105.880 ;
        RECT 21.720 94.980 21.860 105.560 ;
        RECT 27.240 94.980 27.380 113.720 ;
        RECT 27.700 112.340 27.840 113.720 ;
        RECT 27.640 112.020 27.900 112.340 ;
        RECT 30.920 109.280 31.060 143.980 ;
        RECT 31.880 143.105 33.760 143.475 ;
        RECT 34.080 139.220 34.340 139.540 ;
        RECT 35.000 139.220 35.260 139.540 ;
        RECT 31.320 138.880 31.580 139.200 ;
        RECT 31.380 134.100 31.520 138.880 ;
        RECT 31.880 137.665 33.760 138.035 ;
        RECT 34.140 137.160 34.280 139.220 ;
        RECT 34.080 136.840 34.340 137.160 ;
        RECT 35.060 136.480 35.200 139.220 ;
        RECT 35.980 139.200 36.120 147.380 ;
        RECT 35.920 138.880 36.180 139.200 ;
        RECT 35.460 138.200 35.720 138.520 ;
        RECT 35.000 136.160 35.260 136.480 ;
        RECT 35.520 136.140 35.660 138.200 ;
        RECT 35.980 136.820 36.120 138.880 ;
        RECT 35.920 136.500 36.180 136.820 ;
        RECT 35.460 135.820 35.720 136.140 ;
        RECT 35.000 134.460 35.260 134.780 ;
        RECT 31.320 133.780 31.580 134.100 ;
        RECT 34.080 133.780 34.340 134.100 ;
        RECT 31.380 131.380 31.520 133.780 ;
        RECT 31.880 132.225 33.760 132.595 ;
        RECT 34.140 132.060 34.280 133.780 ;
        RECT 34.540 133.100 34.800 133.420 ;
        RECT 34.080 131.740 34.340 132.060 ;
        RECT 31.320 131.060 31.580 131.380 ;
        RECT 34.600 129.340 34.740 133.100 ;
        RECT 34.540 129.020 34.800 129.340 ;
        RECT 34.080 128.000 34.340 128.320 ;
        RECT 31.320 127.320 31.580 127.640 ;
        RECT 31.380 117.780 31.520 127.320 ;
        RECT 31.880 126.785 33.760 127.155 ;
        RECT 33.620 125.620 33.880 125.940 ;
        RECT 33.680 122.880 33.820 125.620 ;
        RECT 33.620 122.560 33.880 122.880 ;
        RECT 34.140 122.200 34.280 128.000 ;
        RECT 34.540 122.900 34.800 123.220 ;
        RECT 34.080 121.880 34.340 122.200 ;
        RECT 31.880 121.345 33.760 121.715 ;
        RECT 34.600 120.500 34.740 122.900 ;
        RECT 35.060 122.620 35.200 134.460 ;
        RECT 36.440 133.760 36.580 173.900 ;
        RECT 37.300 163.360 37.560 163.680 ;
        RECT 37.360 161.300 37.500 163.360 ;
        RECT 37.300 160.980 37.560 161.300 ;
        RECT 36.840 143.640 37.100 143.960 ;
        RECT 35.920 133.440 36.180 133.760 ;
        RECT 36.380 133.440 36.640 133.760 ;
        RECT 35.980 124.920 36.120 133.440 ;
        RECT 36.380 132.760 36.640 133.080 ;
        RECT 36.440 129.000 36.580 132.760 ;
        RECT 36.900 129.340 37.040 143.640 ;
        RECT 37.300 138.880 37.560 139.200 ;
        RECT 37.360 137.500 37.500 138.880 ;
        RECT 37.300 137.180 37.560 137.500 ;
        RECT 37.820 133.760 37.960 174.920 ;
        RECT 38.740 174.560 38.880 184.440 ;
        RECT 40.120 177.620 40.260 189.880 ;
        RECT 43.340 185.780 43.480 190.900 ;
        RECT 43.800 190.200 43.940 195.320 ;
        RECT 46.100 193.940 46.240 198.720 ;
        RECT 46.500 196.340 46.760 196.660 ;
        RECT 46.040 193.620 46.300 193.940 ;
        RECT 46.560 191.220 46.700 196.340 ;
        RECT 46.880 194.785 48.760 195.155 ;
        RECT 49.320 194.620 49.460 198.720 ;
        RECT 51.100 195.660 51.360 195.980 ;
        RECT 50.180 195.320 50.440 195.640 ;
        RECT 49.260 194.300 49.520 194.620 ;
        RECT 50.240 193.940 50.380 195.320 ;
        RECT 49.720 193.620 49.980 193.940 ;
        RECT 50.180 193.620 50.440 193.940 ;
        RECT 49.260 193.280 49.520 193.600 ;
        RECT 46.500 190.900 46.760 191.220 ;
        RECT 43.740 189.880 44.000 190.200 ;
        RECT 46.040 189.880 46.300 190.200 ;
        RECT 43.280 185.460 43.540 185.780 ;
        RECT 40.520 184.780 40.780 185.100 ;
        RECT 40.580 183.740 40.720 184.780 ;
        RECT 44.200 184.440 44.460 184.760 ;
        RECT 40.520 183.420 40.780 183.740 ;
        RECT 40.580 180.000 40.720 183.420 ;
        RECT 44.260 183.400 44.400 184.440 ;
        RECT 44.200 183.080 44.460 183.400 ;
        RECT 40.980 181.720 41.240 182.040 ;
        RECT 40.520 179.680 40.780 180.000 ;
        RECT 40.580 178.300 40.720 179.680 ;
        RECT 41.040 179.320 41.180 181.720 ;
        RECT 45.120 179.680 45.380 180.000 ;
        RECT 44.660 179.340 44.920 179.660 ;
        RECT 40.980 179.000 41.240 179.320 ;
        RECT 40.520 177.980 40.780 178.300 ;
        RECT 39.600 177.300 39.860 177.620 ;
        RECT 40.060 177.300 40.320 177.620 ;
        RECT 39.660 174.560 39.800 177.300 ;
        RECT 41.040 174.560 41.180 179.000 ;
        RECT 44.720 177.620 44.860 179.340 ;
        RECT 41.900 177.300 42.160 177.620 ;
        RECT 44.660 177.530 44.920 177.620 ;
        RECT 44.260 177.390 44.920 177.530 ;
        RECT 41.440 176.960 41.700 177.280 ;
        RECT 38.680 174.240 38.940 174.560 ;
        RECT 39.600 174.240 39.860 174.560 ;
        RECT 40.980 174.240 41.240 174.560 ;
        RECT 39.660 166.820 39.800 174.240 ;
        RECT 41.500 173.940 41.640 176.960 ;
        RECT 41.960 174.560 42.100 177.300 ;
        RECT 44.260 176.940 44.400 177.390 ;
        RECT 44.660 177.300 44.920 177.390 ;
        RECT 44.200 176.620 44.460 176.940 ;
        RECT 44.660 176.620 44.920 176.940 ;
        RECT 42.360 176.280 42.620 176.600 ;
        RECT 41.900 174.240 42.160 174.560 ;
        RECT 41.500 173.800 42.100 173.940 ;
        RECT 40.060 168.460 40.320 168.780 ;
        RECT 40.120 167.420 40.260 168.460 ;
        RECT 40.060 167.100 40.320 167.420 ;
        RECT 39.140 166.420 39.400 166.740 ;
        RECT 39.660 166.680 40.260 166.820 ;
        RECT 39.200 164.700 39.340 166.420 ;
        RECT 40.120 164.700 40.260 166.680 ;
        RECT 39.140 164.380 39.400 164.700 ;
        RECT 40.060 164.380 40.320 164.700 ;
        RECT 40.120 161.890 40.260 164.380 ;
        RECT 40.520 163.020 40.780 163.340 ;
        RECT 38.280 161.750 40.260 161.890 ;
        RECT 38.280 161.300 38.420 161.750 ;
        RECT 40.580 161.640 40.720 163.020 ;
        RECT 38.220 160.980 38.480 161.300 ;
        RECT 38.680 160.980 38.940 161.300 ;
        RECT 39.140 160.980 39.400 161.300 ;
        RECT 39.590 161.125 39.870 161.495 ;
        RECT 40.520 161.320 40.780 161.640 ;
        RECT 41.960 161.210 42.100 173.800 ;
        RECT 39.600 160.980 39.860 161.125 ;
        RECT 41.500 161.070 42.100 161.210 ;
        RECT 38.740 156.200 38.880 160.980 ;
        RECT 39.200 160.815 39.340 160.980 ;
        RECT 39.130 160.445 39.410 160.815 ;
        RECT 40.060 160.640 40.320 160.960 ;
        RECT 39.140 158.940 39.400 159.260 ;
        RECT 38.680 155.880 38.940 156.200 ;
        RECT 39.200 155.520 39.340 158.940 ;
        RECT 39.140 155.200 39.400 155.520 ;
        RECT 39.200 151.100 39.340 155.200 ;
        RECT 39.140 150.780 39.400 151.100 ;
        RECT 39.140 149.080 39.400 149.400 ;
        RECT 38.220 140.920 38.480 141.240 ;
        RECT 37.760 133.440 38.020 133.760 ;
        RECT 37.760 132.760 38.020 133.080 ;
        RECT 36.840 129.020 37.100 129.340 ;
        RECT 36.380 128.680 36.640 129.000 ;
        RECT 36.380 124.940 36.640 125.260 ;
        RECT 35.920 124.600 36.180 124.920 ;
        RECT 35.980 123.220 36.120 124.600 ;
        RECT 35.920 122.900 36.180 123.220 ;
        RECT 35.060 122.480 36.120 122.620 ;
        RECT 34.540 120.410 34.800 120.500 ;
        RECT 34.540 120.270 35.660 120.410 ;
        RECT 34.540 120.180 34.800 120.270 ;
        RECT 32.240 119.840 32.500 120.160 ;
        RECT 32.300 118.460 32.440 119.840 ;
        RECT 32.240 118.140 32.500 118.460 ;
        RECT 31.320 117.460 31.580 117.780 ;
        RECT 31.880 115.905 33.760 116.275 ;
        RECT 35.520 114.720 35.660 120.270 ;
        RECT 35.980 114.720 36.120 122.480 ;
        RECT 36.440 121.180 36.580 124.940 ;
        RECT 36.380 120.860 36.640 121.180 ;
        RECT 35.460 114.400 35.720 114.720 ;
        RECT 35.920 114.400 36.180 114.720 ;
        RECT 31.320 112.700 31.580 113.020 ;
        RECT 30.860 108.960 31.120 109.280 ;
        RECT 21.650 92.980 21.930 94.980 ;
        RECT 27.170 92.980 27.450 94.980 ;
        RECT 31.380 94.740 31.520 112.700 ;
        RECT 35.520 112.000 35.660 114.400 ;
        RECT 35.920 113.720 36.180 114.040 ;
        RECT 35.980 113.020 36.120 113.720 ;
        RECT 35.920 112.700 36.180 113.020 ;
        RECT 36.840 112.700 37.100 113.020 ;
        RECT 35.460 111.680 35.720 112.000 ;
        RECT 36.900 111.910 37.040 112.700 ;
        RECT 37.820 112.340 37.960 132.760 ;
        RECT 38.280 114.720 38.420 140.920 ;
        RECT 38.680 139.220 38.940 139.540 ;
        RECT 38.740 137.500 38.880 139.220 ;
        RECT 38.680 137.180 38.940 137.500 ;
        RECT 39.200 134.780 39.340 149.080 ;
        RECT 40.120 142.260 40.260 160.640 ;
        RECT 40.980 150.100 41.240 150.420 ;
        RECT 41.040 147.360 41.180 150.100 ;
        RECT 40.980 147.040 41.240 147.360 ;
        RECT 40.520 146.360 40.780 146.680 ;
        RECT 40.060 141.940 40.320 142.260 ;
        RECT 39.600 138.200 39.860 138.520 ;
        RECT 39.660 136.820 39.800 138.200 ;
        RECT 39.600 136.500 39.860 136.820 ;
        RECT 39.140 134.460 39.400 134.780 ;
        RECT 40.580 134.100 40.720 146.360 ;
        RECT 41.500 144.640 41.640 161.070 ;
        RECT 41.900 157.920 42.160 158.240 ;
        RECT 41.960 156.540 42.100 157.920 ;
        RECT 41.900 156.220 42.160 156.540 ;
        RECT 41.900 152.140 42.160 152.460 ;
        RECT 41.960 150.420 42.100 152.140 ;
        RECT 41.900 150.100 42.160 150.420 ;
        RECT 41.900 149.080 42.160 149.400 ;
        RECT 41.960 147.360 42.100 149.080 ;
        RECT 41.900 147.040 42.160 147.360 ;
        RECT 41.900 145.000 42.160 145.320 ;
        RECT 41.440 144.320 41.700 144.640 ;
        RECT 41.960 140.220 42.100 145.000 ;
        RECT 42.420 144.640 42.560 176.280 ;
        RECT 44.260 174.220 44.400 176.620 ;
        RECT 44.200 173.900 44.460 174.220 ;
        RECT 44.720 172.520 44.860 176.620 ;
        RECT 45.180 175.580 45.320 179.680 ;
        RECT 45.580 179.000 45.840 179.320 ;
        RECT 45.120 175.260 45.380 175.580 ;
        RECT 44.660 172.200 44.920 172.520 ;
        RECT 45.180 172.180 45.320 175.260 ;
        RECT 45.120 171.860 45.380 172.180 ;
        RECT 43.740 171.520 44.000 171.840 ;
        RECT 42.820 170.840 43.080 171.160 ;
        RECT 42.880 167.080 43.020 170.840 ;
        RECT 43.800 169.120 43.940 171.520 ;
        RECT 44.660 170.840 44.920 171.160 ;
        RECT 43.740 168.800 44.000 169.120 ;
        RECT 42.820 166.760 43.080 167.080 ;
        RECT 42.820 166.080 43.080 166.400 ;
        RECT 42.880 163.000 43.020 166.080 ;
        RECT 42.820 162.680 43.080 163.000 ;
        RECT 42.880 156.540 43.020 162.680 ;
        RECT 43.800 160.140 43.940 168.800 ;
        RECT 43.340 160.000 43.940 160.140 ;
        RECT 43.340 158.580 43.480 160.000 ;
        RECT 43.280 158.260 43.540 158.580 ;
        RECT 44.200 157.920 44.460 158.240 ;
        RECT 42.820 156.220 43.080 156.540 ;
        RECT 44.260 155.860 44.400 157.920 ;
        RECT 44.200 155.540 44.460 155.860 ;
        RECT 44.260 153.480 44.400 155.540 ;
        RECT 44.200 153.160 44.460 153.480 ;
        RECT 43.730 152.540 44.010 152.655 ;
        RECT 44.200 152.540 44.460 152.800 ;
        RECT 43.730 152.480 44.460 152.540 ;
        RECT 43.730 152.400 44.400 152.480 ;
        RECT 43.730 152.285 44.010 152.400 ;
        RECT 43.280 151.800 43.540 152.120 ;
        RECT 42.810 150.245 43.090 150.615 ;
        RECT 42.820 150.100 43.080 150.245 ;
        RECT 42.820 149.080 43.080 149.400 ;
        RECT 42.880 144.980 43.020 149.080 ;
        RECT 43.340 144.980 43.480 151.800 ;
        RECT 43.800 150.420 43.940 152.285 ;
        RECT 44.200 151.800 44.460 152.120 ;
        RECT 43.740 150.100 44.000 150.420 ;
        RECT 44.260 150.080 44.400 151.800 ;
        RECT 44.200 149.935 44.460 150.080 ;
        RECT 44.190 149.565 44.470 149.935 ;
        RECT 44.260 147.700 44.400 149.565 ;
        RECT 44.200 147.380 44.460 147.700 ;
        RECT 42.820 144.660 43.080 144.980 ;
        RECT 43.280 144.660 43.540 144.980 ;
        RECT 42.360 144.320 42.620 144.640 ;
        RECT 42.820 143.640 43.080 143.960 ;
        RECT 44.200 143.640 44.460 143.960 ;
        RECT 41.900 139.900 42.160 140.220 ;
        RECT 41.900 139.220 42.160 139.540 ;
        RECT 41.960 137.500 42.100 139.220 ;
        RECT 41.900 137.180 42.160 137.500 ;
        RECT 40.520 133.780 40.780 134.100 ;
        RECT 42.360 133.100 42.620 133.420 ;
        RECT 42.420 128.660 42.560 133.100 ;
        RECT 42.880 130.270 43.020 143.640 ;
        RECT 43.740 142.620 44.000 142.940 ;
        RECT 43.270 135.965 43.550 136.335 ;
        RECT 43.340 134.440 43.480 135.965 ;
        RECT 43.280 134.120 43.540 134.440 ;
        RECT 43.340 131.040 43.480 134.120 ;
        RECT 43.280 130.720 43.540 131.040 ;
        RECT 42.880 130.130 43.480 130.270 ;
        RECT 42.360 128.340 42.620 128.660 ;
        RECT 42.820 128.000 43.080 128.320 ;
        RECT 42.880 126.620 43.020 128.000 ;
        RECT 42.820 126.300 43.080 126.620 ;
        RECT 42.880 125.600 43.020 126.300 ;
        RECT 40.060 125.280 40.320 125.600 ;
        RECT 42.820 125.510 43.080 125.600 ;
        RECT 42.420 125.370 43.080 125.510 ;
        RECT 40.120 123.560 40.260 125.280 ;
        RECT 40.060 123.240 40.320 123.560 ;
        RECT 42.420 122.880 42.560 125.370 ;
        RECT 42.820 125.280 43.080 125.370 ;
        RECT 42.820 123.240 43.080 123.560 ;
        RECT 42.360 122.560 42.620 122.880 ;
        RECT 42.880 121.180 43.020 123.240 ;
        RECT 42.820 120.860 43.080 121.180 ;
        RECT 43.340 114.720 43.480 130.130 ;
        RECT 43.800 128.660 43.940 142.620 ;
        RECT 44.260 140.220 44.400 143.640 ;
        RECT 44.720 141.580 44.860 170.840 ;
        RECT 45.120 168.800 45.380 169.120 ;
        RECT 45.180 165.720 45.320 168.800 ;
        RECT 45.120 165.400 45.380 165.720 ;
        RECT 45.180 163.340 45.320 165.400 ;
        RECT 45.120 163.020 45.380 163.340 ;
        RECT 45.120 159.960 45.380 160.280 ;
        RECT 45.180 144.980 45.320 159.960 ;
        RECT 45.120 144.660 45.380 144.980 ;
        RECT 45.640 144.640 45.780 179.000 ;
        RECT 46.100 172.180 46.240 189.880 ;
        RECT 46.880 189.345 48.760 189.715 ;
        RECT 46.500 187.160 46.760 187.480 ;
        RECT 46.560 184.760 46.700 187.160 ;
        RECT 46.500 184.440 46.760 184.760 ;
        RECT 46.560 180.340 46.700 184.440 ;
        RECT 46.880 183.905 48.760 184.275 ;
        RECT 49.320 183.060 49.460 193.280 ;
        RECT 49.780 191.900 49.920 193.620 ;
        RECT 49.720 191.580 49.980 191.900 ;
        RECT 49.720 184.440 49.980 184.760 ;
        RECT 49.780 183.060 49.920 184.440 ;
        RECT 49.260 182.740 49.520 183.060 ;
        RECT 49.720 182.740 49.980 183.060 ;
        RECT 46.500 180.020 46.760 180.340 ;
        RECT 48.340 179.680 48.600 180.000 ;
        RECT 48.400 179.320 48.540 179.680 ;
        RECT 48.340 179.000 48.600 179.320 ;
        RECT 46.880 178.465 48.760 178.835 ;
        RECT 47.880 177.300 48.140 177.620 ;
        RECT 48.330 177.445 48.610 177.815 ;
        RECT 48.340 177.300 48.600 177.445 ;
        RECT 47.940 176.940 48.080 177.300 ;
        RECT 47.880 176.620 48.140 176.940 ;
        RECT 46.500 176.280 46.760 176.600 ;
        RECT 46.040 171.860 46.300 172.180 ;
        RECT 46.040 164.040 46.300 164.360 ;
        RECT 46.100 161.300 46.240 164.040 ;
        RECT 46.040 160.980 46.300 161.300 ;
        RECT 46.040 159.960 46.300 160.280 ;
        RECT 46.100 158.580 46.240 159.960 ;
        RECT 46.040 158.260 46.300 158.580 ;
        RECT 46.560 157.980 46.700 176.280 ;
        RECT 48.400 175.580 48.540 177.300 ;
        RECT 48.340 175.260 48.600 175.580 ;
        RECT 46.880 173.025 48.760 173.395 ;
        RECT 47.410 172.005 47.690 172.375 ;
        RECT 47.420 171.860 47.680 172.005 ;
        RECT 47.480 169.655 47.620 171.860 ;
        RECT 47.410 169.285 47.690 169.655 ;
        RECT 49.320 168.780 49.460 182.740 ;
        RECT 50.180 179.680 50.440 180.000 ;
        RECT 50.240 178.300 50.380 179.680 ;
        RECT 50.180 177.980 50.440 178.300 ;
        RECT 50.240 177.620 50.380 177.980 ;
        RECT 51.160 177.620 51.300 195.660 ;
        RECT 52.540 194.620 52.680 199.400 ;
        RECT 63.520 198.950 63.780 199.040 ;
        RECT 63.520 198.810 64.180 198.950 ;
        RECT 63.520 198.720 63.780 198.810 ;
        RECT 54.780 198.040 55.040 198.360 ;
        RECT 54.840 195.980 54.980 198.040 ;
        RECT 61.880 197.505 63.760 197.875 ;
        RECT 54.780 195.660 55.040 195.980 ;
        RECT 56.160 195.320 56.420 195.640 ;
        RECT 61.220 195.320 61.480 195.640 ;
        RECT 52.480 194.300 52.740 194.620 ;
        RECT 56.220 192.920 56.360 195.320 ;
        RECT 61.280 194.280 61.420 195.320 ;
        RECT 57.540 193.960 57.800 194.280 ;
        RECT 61.220 193.960 61.480 194.280 ;
        RECT 56.160 192.600 56.420 192.920 ;
        RECT 54.780 190.560 55.040 190.880 ;
        RECT 53.400 189.880 53.660 190.200 ;
        RECT 53.460 188.840 53.600 189.880 ;
        RECT 53.400 188.520 53.660 188.840 ;
        RECT 54.840 186.460 54.980 190.560 ;
        RECT 54.780 186.140 55.040 186.460 ;
        RECT 52.020 185.460 52.280 185.780 ;
        RECT 52.080 181.020 52.220 185.460 ;
        RECT 54.320 184.440 54.580 184.760 ;
        RECT 52.020 180.700 52.280 181.020 ;
        RECT 51.560 180.360 51.820 180.680 ;
        RECT 51.620 179.320 51.760 180.360 ;
        RECT 52.080 180.340 52.220 180.700 ;
        RECT 52.020 180.020 52.280 180.340 ;
        RECT 54.380 179.660 54.520 184.440 ;
        RECT 56.220 179.660 56.360 192.600 ;
        RECT 57.600 191.900 57.740 193.960 ;
        RECT 64.040 193.600 64.180 198.810 ;
        RECT 71.400 198.360 71.540 199.400 ;
        RECT 72.320 199.040 72.460 201.440 ;
        RECT 72.260 198.720 72.520 199.040 ;
        RECT 71.340 198.040 71.600 198.360 ;
        RECT 72.260 198.040 72.520 198.360 ;
        RECT 71.400 196.660 71.540 198.040 ;
        RECT 72.320 196.660 72.460 198.040 ;
        RECT 72.780 197.340 72.920 201.780 ;
        RECT 76.880 200.225 78.760 200.595 ;
        RECT 106.880 200.225 108.760 200.595 ;
        RECT 77.780 199.400 78.040 199.720 ;
        RECT 100.780 199.400 101.040 199.720 ;
        RECT 111.360 199.400 111.620 199.720 ;
        RECT 121.020 199.400 121.280 199.720 ;
        RECT 74.100 199.060 74.360 199.380 ;
        RECT 75.020 199.060 75.280 199.380 ;
        RECT 72.720 197.020 72.980 197.340 ;
        RECT 71.340 196.340 71.600 196.660 ;
        RECT 72.260 196.570 72.520 196.660 ;
        RECT 71.860 196.430 72.520 196.570 ;
        RECT 67.200 195.320 67.460 195.640 ;
        RECT 70.880 195.320 71.140 195.640 ;
        RECT 67.260 194.280 67.400 195.320 ;
        RECT 67.200 193.960 67.460 194.280 ;
        RECT 58.000 193.280 58.260 193.600 ;
        RECT 63.980 193.280 64.240 193.600 ;
        RECT 57.540 191.580 57.800 191.900 ;
        RECT 58.060 190.880 58.200 193.280 ;
        RECT 61.880 192.065 63.760 192.435 ;
        RECT 58.000 190.560 58.260 190.880 ;
        RECT 61.220 190.560 61.480 190.880 ;
        RECT 56.620 189.880 56.880 190.200 ;
        RECT 56.680 188.840 56.820 189.880 ;
        RECT 56.620 188.520 56.880 188.840 ;
        RECT 57.080 188.520 57.340 188.840 ;
        RECT 57.140 185.440 57.280 188.520 ;
        RECT 61.280 188.500 61.420 190.560 ;
        RECT 61.220 188.180 61.480 188.500 ;
        RECT 57.080 185.120 57.340 185.440 ;
        RECT 56.620 182.740 56.880 183.060 ;
        RECT 56.680 181.020 56.820 182.740 ;
        RECT 56.620 180.700 56.880 181.020 ;
        RECT 54.320 179.340 54.580 179.660 ;
        RECT 56.160 179.340 56.420 179.660 ;
        RECT 59.840 179.340 60.100 179.660 ;
        RECT 51.560 179.000 51.820 179.320 ;
        RECT 53.860 179.000 54.120 179.320 ;
        RECT 51.620 177.620 51.760 179.000 ;
        RECT 53.920 178.300 54.060 179.000 ;
        RECT 53.860 177.980 54.120 178.300 ;
        RECT 50.180 177.300 50.440 177.620 ;
        RECT 51.100 177.300 51.360 177.620 ;
        RECT 51.560 177.300 51.820 177.620 ;
        RECT 52.010 177.530 52.290 177.815 ;
        RECT 52.010 177.445 52.680 177.530 ;
        RECT 52.020 177.390 52.680 177.445 ;
        RECT 52.020 177.300 52.280 177.390 ;
        RECT 50.240 175.580 50.380 177.300 ;
        RECT 51.620 176.940 51.760 177.300 ;
        RECT 51.560 176.620 51.820 176.940 ;
        RECT 50.180 175.260 50.440 175.580 ;
        RECT 51.620 175.095 51.760 176.620 ;
        RECT 51.550 174.725 51.830 175.095 ;
        RECT 52.020 174.920 52.280 175.240 ;
        RECT 51.100 173.900 51.360 174.220 ;
        RECT 50.640 169.480 50.900 169.800 ;
        RECT 50.180 168.800 50.440 169.120 ;
        RECT 49.260 168.460 49.520 168.780 ;
        RECT 46.880 167.585 48.760 167.955 ;
        RECT 49.320 166.740 49.460 168.460 ;
        RECT 49.720 168.120 49.980 168.440 ;
        RECT 49.260 166.420 49.520 166.740 ;
        RECT 47.880 166.080 48.140 166.400 ;
        RECT 47.940 164.700 48.080 166.080 ;
        RECT 49.260 165.400 49.520 165.720 ;
        RECT 47.880 164.380 48.140 164.700 ;
        RECT 46.880 162.145 48.760 162.515 ;
        RECT 48.340 161.660 48.600 161.980 ;
        RECT 46.950 161.125 47.230 161.495 ;
        RECT 46.960 160.980 47.220 161.125 ;
        RECT 47.420 160.815 47.680 160.960 ;
        RECT 47.410 160.445 47.690 160.815 ;
        RECT 46.100 157.840 46.700 157.980 ;
        RECT 47.480 158.150 47.620 160.445 ;
        RECT 48.400 158.240 48.540 161.660 ;
        RECT 49.320 161.640 49.460 165.400 ;
        RECT 49.780 163.680 49.920 168.120 ;
        RECT 50.240 165.720 50.380 168.800 ;
        RECT 50.180 165.400 50.440 165.720 ;
        RECT 50.700 164.020 50.840 169.480 ;
        RECT 50.640 163.700 50.900 164.020 ;
        RECT 49.720 163.360 49.980 163.680 ;
        RECT 49.260 161.380 49.520 161.640 ;
        RECT 48.860 161.320 49.520 161.380 ;
        RECT 48.860 161.240 49.460 161.320 ;
        RECT 48.860 158.580 49.000 161.240 ;
        RECT 50.700 160.620 50.840 163.700 ;
        RECT 50.640 160.300 50.900 160.620 ;
        RECT 49.260 159.960 49.520 160.280 ;
        RECT 48.800 158.260 49.060 158.580 ;
        RECT 47.880 158.150 48.140 158.240 ;
        RECT 47.480 158.010 48.140 158.150 ;
        RECT 46.100 145.060 46.240 157.840 ;
        RECT 47.480 157.470 47.620 158.010 ;
        RECT 47.880 157.920 48.140 158.010 ;
        RECT 48.340 157.920 48.600 158.240 ;
        RECT 46.560 157.330 47.620 157.470 ;
        RECT 46.560 155.860 46.700 157.330 ;
        RECT 46.880 156.705 48.760 157.075 ;
        RECT 46.500 155.540 46.760 155.860 ;
        RECT 48.340 154.520 48.600 154.840 ;
        RECT 48.400 152.800 48.540 154.520 ;
        RECT 48.340 152.480 48.600 152.800 ;
        RECT 46.880 151.265 48.760 151.635 ;
        RECT 46.490 150.245 46.770 150.615 ;
        RECT 46.500 150.100 46.760 150.245 ;
        RECT 46.560 147.360 46.700 150.100 ;
        RECT 46.500 147.040 46.760 147.360 ;
        RECT 46.880 145.825 48.760 146.195 ;
        RECT 46.100 144.920 48.080 145.060 ;
        RECT 49.320 144.980 49.460 159.960 ;
        RECT 49.720 157.920 49.980 158.240 ;
        RECT 49.780 155.860 49.920 157.920 ;
        RECT 50.180 157.240 50.440 157.560 ;
        RECT 49.720 155.540 49.980 155.860 ;
        RECT 49.720 153.500 49.980 153.820 ;
        RECT 47.940 144.640 48.080 144.920 ;
        RECT 49.260 144.660 49.520 144.980 ;
        RECT 45.580 144.320 45.840 144.640 ;
        RECT 47.880 144.320 48.140 144.640 ;
        RECT 45.580 143.640 45.840 143.960 ;
        RECT 46.500 143.640 46.760 143.960 ;
        RECT 48.340 143.640 48.600 143.960 ;
        RECT 48.800 143.640 49.060 143.960 ;
        RECT 45.120 141.600 45.380 141.920 ;
        RECT 44.660 141.260 44.920 141.580 ;
        RECT 44.200 139.900 44.460 140.220 ;
        RECT 45.180 136.140 45.320 141.600 ;
        RECT 45.120 135.820 45.380 136.140 ;
        RECT 44.200 135.480 44.460 135.800 ;
        RECT 44.260 133.760 44.400 135.480 ;
        RECT 44.200 133.440 44.460 133.760 ;
        RECT 44.260 132.060 44.400 133.440 ;
        RECT 44.200 131.740 44.460 132.060 ;
        RECT 43.740 128.340 44.000 128.660 ;
        RECT 44.660 124.600 44.920 124.920 ;
        RECT 44.720 122.200 44.860 124.600 ;
        RECT 44.660 121.880 44.920 122.200 ;
        RECT 45.640 119.220 45.780 143.640 ;
        RECT 46.040 141.600 46.300 141.920 ;
        RECT 46.100 139.540 46.240 141.600 ;
        RECT 46.560 140.220 46.700 143.640 ;
        RECT 48.400 142.340 48.540 143.640 ;
        RECT 48.860 142.940 49.000 143.640 ;
        RECT 48.800 142.620 49.060 142.940 ;
        RECT 48.400 142.200 49.460 142.340 ;
        RECT 46.880 140.385 48.760 140.755 ;
        RECT 46.500 139.900 46.760 140.220 ;
        RECT 46.040 139.220 46.300 139.540 ;
        RECT 46.040 135.480 46.300 135.800 ;
        RECT 46.100 130.700 46.240 135.480 ;
        RECT 46.880 134.945 48.760 135.315 ;
        RECT 49.320 130.780 49.460 142.200 ;
        RECT 49.780 139.200 49.920 153.500 ;
        RECT 50.240 147.360 50.380 157.240 ;
        RECT 50.640 153.160 50.900 153.480 ;
        RECT 50.700 152.540 50.840 153.160 ;
        RECT 51.160 153.140 51.300 173.900 ;
        RECT 51.560 169.140 51.820 169.460 ;
        RECT 51.620 158.580 51.760 169.140 ;
        RECT 51.560 158.260 51.820 158.580 ;
        RECT 51.560 157.240 51.820 157.560 ;
        RECT 51.100 152.820 51.360 153.140 ;
        RECT 51.620 152.800 51.760 157.240 ;
        RECT 52.080 153.140 52.220 174.920 ;
        RECT 52.540 174.560 52.680 177.390 ;
        RECT 52.940 176.280 53.200 176.600 ;
        RECT 52.480 174.240 52.740 174.560 ;
        RECT 52.480 160.300 52.740 160.620 ;
        RECT 52.540 158.240 52.680 160.300 ;
        RECT 52.480 157.920 52.740 158.240 ;
        RECT 52.480 153.500 52.740 153.820 ;
        RECT 52.020 152.820 52.280 153.140 ;
        RECT 50.700 152.400 51.300 152.540 ;
        RECT 51.560 152.480 51.820 152.800 ;
        RECT 50.640 151.800 50.900 152.120 ;
        RECT 50.700 150.420 50.840 151.800 ;
        RECT 50.640 150.100 50.900 150.420 ;
        RECT 51.160 149.820 51.300 152.400 ;
        RECT 50.700 149.680 51.300 149.820 ;
        RECT 50.180 147.040 50.440 147.360 ;
        RECT 50.180 146.360 50.440 146.680 ;
        RECT 50.240 145.320 50.380 146.360 ;
        RECT 50.180 145.000 50.440 145.320 ;
        RECT 49.720 138.880 49.980 139.200 ;
        RECT 50.180 138.880 50.440 139.200 ;
        RECT 50.240 138.260 50.380 138.880 ;
        RECT 49.780 138.120 50.380 138.260 ;
        RECT 49.780 133.760 49.920 138.120 ;
        RECT 50.180 135.480 50.440 135.800 ;
        RECT 49.720 133.440 49.980 133.760 ;
        RECT 49.720 132.760 49.980 133.080 ;
        RECT 49.780 131.720 49.920 132.760 ;
        RECT 49.720 131.400 49.980 131.720 ;
        RECT 50.240 131.380 50.380 135.480 ;
        RECT 50.180 131.060 50.440 131.380 ;
        RECT 46.040 130.380 46.300 130.700 ;
        RECT 49.320 130.640 50.380 130.780 ;
        RECT 49.260 130.040 49.520 130.360 ;
        RECT 46.880 129.505 48.760 129.875 ;
        RECT 49.320 129.000 49.460 130.040 ;
        RECT 49.260 128.680 49.520 129.000 ;
        RECT 49.260 128.000 49.520 128.320 ;
        RECT 46.040 124.600 46.300 124.920 ;
        RECT 46.100 120.160 46.240 124.600 ;
        RECT 46.880 124.065 48.760 124.435 ;
        RECT 49.320 123.220 49.460 128.000 ;
        RECT 49.260 122.900 49.520 123.220 ;
        RECT 46.500 122.560 46.760 122.880 ;
        RECT 46.560 121.180 46.700 122.560 ;
        RECT 46.500 120.860 46.760 121.180 ;
        RECT 46.040 119.840 46.300 120.160 ;
        RECT 45.640 119.080 46.240 119.220 ;
        RECT 38.220 114.400 38.480 114.720 ;
        RECT 43.280 114.400 43.540 114.720 ;
        RECT 40.060 114.060 40.320 114.380 ;
        RECT 38.680 113.720 38.940 114.040 ;
        RECT 37.760 112.020 38.020 112.340 ;
        RECT 36.670 111.770 37.040 111.910 ;
        RECT 31.880 110.465 33.760 110.835 ;
        RECT 35.520 110.300 35.660 111.680 ;
        RECT 36.670 111.060 36.810 111.770 ;
        RECT 35.980 110.920 36.810 111.060 ;
        RECT 33.620 109.980 33.880 110.300 ;
        RECT 35.460 109.980 35.720 110.300 ;
        RECT 32.240 108.280 32.500 108.600 ;
        RECT 32.300 107.240 32.440 108.280 ;
        RECT 32.240 106.920 32.500 107.240 ;
        RECT 33.680 106.900 33.820 109.980 ;
        RECT 35.980 109.620 36.120 110.920 ;
        RECT 35.920 109.300 36.180 109.620 ;
        RECT 38.740 109.280 38.880 113.720 ;
        RECT 40.120 112.340 40.260 114.060 ;
        RECT 46.100 113.020 46.240 119.080 ;
        RECT 46.880 118.625 48.760 118.995 ;
        RECT 49.320 114.460 49.460 122.900 ;
        RECT 50.240 114.720 50.380 130.640 ;
        RECT 50.700 115.060 50.840 149.680 ;
        RECT 52.020 148.060 52.280 148.380 ;
        RECT 52.080 139.200 52.220 148.060 ;
        RECT 52.020 138.880 52.280 139.200 ;
        RECT 52.540 137.500 52.680 153.500 ;
        RECT 53.000 147.700 53.140 176.280 ;
        RECT 53.920 174.900 54.060 177.980 ;
        RECT 54.380 177.960 54.520 179.340 ;
        RECT 54.320 177.640 54.580 177.960 ;
        RECT 58.920 177.640 59.180 177.960 ;
        RECT 58.460 176.960 58.720 177.280 ;
        RECT 56.620 175.260 56.880 175.580 ;
        RECT 56.680 175.095 56.820 175.260 ;
        RECT 53.860 174.580 54.120 174.900 ;
        RECT 55.230 174.725 55.510 175.095 ;
        RECT 56.610 174.725 56.890 175.095 ;
        RECT 55.300 174.560 55.440 174.725 ;
        RECT 56.680 174.560 56.820 174.725 ;
        RECT 55.240 174.240 55.500 174.560 ;
        RECT 56.620 174.240 56.880 174.560 ;
        RECT 55.300 173.880 55.440 174.240 ;
        RECT 55.240 173.560 55.500 173.880 ;
        RECT 58.520 171.840 58.660 176.960 ;
        RECT 58.980 175.580 59.120 177.640 ;
        RECT 58.920 175.260 59.180 175.580 ;
        RECT 59.900 174.560 60.040 179.340 ;
        RECT 60.290 174.725 60.570 175.095 ;
        RECT 60.360 174.560 60.500 174.725 ;
        RECT 61.280 174.560 61.420 188.180 ;
        RECT 64.040 188.160 64.180 193.280 ;
        RECT 69.500 190.900 69.760 191.220 ;
        RECT 63.980 187.840 64.240 188.160 ;
        RECT 61.880 186.625 63.760 186.995 ;
        RECT 64.040 185.440 64.180 187.840 ;
        RECT 63.980 185.120 64.240 185.440 ;
        RECT 62.600 184.780 62.860 185.100 ;
        RECT 62.660 183.740 62.800 184.780 ;
        RECT 62.600 183.420 62.860 183.740 ;
        RECT 61.880 181.185 63.760 181.555 ;
        RECT 64.040 177.280 64.180 185.120 ;
        RECT 69.560 184.760 69.700 190.900 ;
        RECT 70.940 190.880 71.080 195.320 ;
        RECT 70.880 190.560 71.140 190.880 ;
        RECT 70.420 189.880 70.680 190.200 ;
        RECT 70.480 184.760 70.620 189.880 ;
        RECT 71.400 188.500 71.540 196.340 ;
        RECT 71.860 190.880 72.000 196.430 ;
        RECT 72.260 196.340 72.520 196.430 ;
        RECT 72.260 193.960 72.520 194.280 ;
        RECT 72.320 191.900 72.460 193.960 ;
        RECT 72.780 191.900 72.920 197.020 ;
        RECT 73.640 196.340 73.900 196.660 ;
        RECT 73.700 194.620 73.840 196.340 ;
        RECT 74.160 194.620 74.300 199.060 ;
        RECT 75.080 196.660 75.220 199.060 ;
        RECT 75.480 198.720 75.740 199.040 ;
        RECT 75.020 196.340 75.280 196.660 ;
        RECT 74.560 196.000 74.820 196.320 ;
        RECT 73.640 194.530 73.900 194.620 ;
        RECT 73.240 194.390 73.900 194.530 ;
        RECT 72.260 191.580 72.520 191.900 ;
        RECT 72.720 191.580 72.980 191.900 ;
        RECT 73.240 191.560 73.380 194.390 ;
        RECT 73.640 194.300 73.900 194.390 ;
        RECT 74.100 194.300 74.360 194.620 ;
        RECT 74.620 193.940 74.760 196.000 ;
        RECT 75.020 195.320 75.280 195.640 ;
        RECT 74.560 193.620 74.820 193.940 ;
        RECT 73.180 191.470 73.440 191.560 ;
        RECT 73.180 191.330 73.840 191.470 ;
        RECT 73.180 191.240 73.440 191.330 ;
        RECT 71.800 190.560 72.060 190.880 ;
        RECT 71.340 188.180 71.600 188.500 ;
        RECT 69.500 184.440 69.760 184.760 ;
        RECT 70.420 184.440 70.680 184.760 ;
        RECT 64.440 179.000 64.700 179.320 ;
        RECT 69.040 179.000 69.300 179.320 ;
        RECT 64.500 177.620 64.640 179.000 ;
        RECT 64.440 177.300 64.700 177.620 ;
        RECT 63.980 176.960 64.240 177.280 ;
        RECT 68.580 177.190 68.840 177.280 ;
        RECT 69.100 177.190 69.240 179.000 ;
        RECT 69.560 177.280 69.700 184.440 ;
        RECT 70.480 177.620 70.620 184.440 ;
        RECT 71.400 183.060 71.540 188.180 ;
        RECT 73.180 187.160 73.440 187.480 ;
        RECT 73.240 185.780 73.380 187.160 ;
        RECT 73.180 185.460 73.440 185.780 ;
        RECT 72.720 184.780 72.980 185.100 ;
        RECT 72.780 183.740 72.920 184.780 ;
        RECT 73.240 183.740 73.380 185.460 ;
        RECT 73.700 185.100 73.840 191.330 ;
        RECT 74.620 191.220 74.760 193.620 ;
        RECT 75.080 193.600 75.220 195.320 ;
        RECT 75.020 193.280 75.280 193.600 ;
        RECT 74.560 190.900 74.820 191.220 ;
        RECT 74.100 190.560 74.360 190.880 ;
        RECT 74.160 185.180 74.300 190.560 ;
        RECT 75.080 185.780 75.220 193.280 ;
        RECT 75.540 192.920 75.680 198.720 ;
        RECT 75.940 198.380 76.200 198.700 ;
        RECT 76.000 195.980 76.140 198.380 ;
        RECT 77.840 197.340 77.980 199.400 ;
        RECT 81.000 199.060 81.260 199.380 ;
        RECT 81.060 198.700 81.200 199.060 ;
        RECT 81.920 198.720 82.180 199.040 ;
        RECT 81.000 198.380 81.260 198.700 ;
        RECT 79.160 198.040 79.420 198.360 ;
        RECT 77.780 197.020 78.040 197.340 ;
        RECT 76.400 196.680 76.660 197.000 ;
        RECT 75.940 195.660 76.200 195.980 ;
        RECT 75.480 192.600 75.740 192.920 ;
        RECT 75.020 185.460 75.280 185.780 ;
        RECT 73.640 184.780 73.900 185.100 ;
        RECT 74.160 185.040 74.760 185.180 ;
        RECT 72.720 183.420 72.980 183.740 ;
        RECT 73.180 183.420 73.440 183.740 ;
        RECT 73.700 183.400 73.840 184.780 ;
        RECT 74.100 184.440 74.360 184.760 ;
        RECT 73.640 183.080 73.900 183.400 ;
        RECT 71.340 182.740 71.600 183.060 ;
        RECT 72.720 181.720 72.980 182.040 ;
        RECT 71.340 179.680 71.600 180.000 ;
        RECT 70.420 177.300 70.680 177.620 ;
        RECT 66.270 176.765 66.550 177.135 ;
        RECT 68.580 177.050 69.240 177.190 ;
        RECT 68.580 176.960 68.840 177.050 ;
        RECT 69.500 176.960 69.760 177.280 ;
        RECT 66.340 176.600 66.480 176.765 ;
        RECT 63.980 176.280 64.240 176.600 ;
        RECT 66.280 176.280 66.540 176.600 ;
        RECT 67.660 176.280 67.920 176.600 ;
        RECT 61.880 175.745 63.760 176.115 ;
        RECT 64.040 175.580 64.180 176.280 ;
        RECT 63.980 175.260 64.240 175.580 ;
        RECT 66.340 174.900 66.480 176.280 ;
        RECT 66.280 174.580 66.540 174.900 ;
        RECT 67.720 174.560 67.860 176.280 ;
        RECT 68.570 175.405 68.850 175.775 ;
        RECT 68.580 175.260 68.840 175.405 ;
        RECT 58.920 174.240 59.180 174.560 ;
        RECT 59.840 174.240 60.100 174.560 ;
        RECT 60.300 174.240 60.560 174.560 ;
        RECT 61.220 174.240 61.480 174.560 ;
        RECT 67.660 174.240 67.920 174.560 ;
        RECT 58.980 174.030 59.120 174.240 ;
        RECT 58.920 173.710 59.180 174.030 ;
        RECT 55.700 171.520 55.960 171.840 ;
        RECT 58.460 171.520 58.720 171.840 ;
        RECT 53.860 171.180 54.120 171.500 ;
        RECT 53.920 169.460 54.060 171.180 ;
        RECT 55.760 170.140 55.900 171.520 ;
        RECT 55.700 169.820 55.960 170.140 ;
        RECT 53.860 169.140 54.120 169.460 ;
        RECT 53.400 166.760 53.660 167.080 ;
        RECT 53.460 164.700 53.600 166.760 ;
        RECT 53.400 164.380 53.660 164.700 ;
        RECT 53.920 163.680 54.060 169.140 ;
        RECT 58.520 169.120 58.660 171.520 ;
        RECT 61.280 169.460 61.420 174.240 ;
        RECT 69.560 171.840 69.700 176.960 ;
        RECT 70.480 175.580 70.620 177.300 ;
        RECT 71.400 176.600 71.540 179.680 ;
        RECT 71.800 179.000 72.060 179.320 ;
        RECT 71.340 176.280 71.600 176.600 ;
        RECT 70.420 175.260 70.680 175.580 ;
        RECT 69.500 171.520 69.760 171.840 ;
        RECT 70.480 171.500 70.620 175.260 ;
        RECT 71.400 174.560 71.540 176.280 ;
        RECT 71.860 175.240 72.000 179.000 ;
        RECT 72.260 176.960 72.520 177.280 ;
        RECT 72.320 175.580 72.460 176.960 ;
        RECT 72.260 175.260 72.520 175.580 ;
        RECT 71.800 174.920 72.060 175.240 ;
        RECT 71.340 174.240 71.600 174.560 ;
        RECT 71.860 172.520 72.000 174.920 ;
        RECT 72.320 174.900 72.460 175.260 ;
        RECT 72.260 174.580 72.520 174.900 ;
        RECT 71.800 172.200 72.060 172.520 ;
        RECT 70.420 171.180 70.680 171.500 ;
        RECT 72.260 171.015 72.520 171.160 ;
        RECT 61.880 170.305 63.760 170.675 ;
        RECT 72.250 170.645 72.530 171.015 ;
        RECT 69.500 169.820 69.760 170.140 ;
        RECT 61.220 169.140 61.480 169.460 ;
        RECT 58.460 168.800 58.720 169.120 ;
        RECT 60.300 168.800 60.560 169.120 ;
        RECT 58.520 166.400 58.660 168.800 ;
        RECT 60.360 166.740 60.500 168.800 ;
        RECT 60.300 166.420 60.560 166.740 ;
        RECT 64.440 166.420 64.700 166.740 ;
        RECT 57.080 166.080 57.340 166.400 ;
        RECT 58.460 166.080 58.720 166.400 ;
        RECT 57.140 164.700 57.280 166.080 ;
        RECT 58.000 165.400 58.260 165.720 ;
        RECT 57.080 164.380 57.340 164.700 ;
        RECT 53.860 163.360 54.120 163.680 ;
        RECT 54.320 163.360 54.580 163.680 ;
        RECT 54.380 161.980 54.520 163.360 ;
        RECT 58.060 163.000 58.200 165.400 ;
        RECT 58.520 164.020 58.660 166.080 ;
        RECT 61.880 164.865 63.760 165.235 ;
        RECT 58.460 163.700 58.720 164.020 ;
        RECT 58.000 162.680 58.260 163.000 ;
        RECT 59.840 162.910 60.100 163.000 ;
        RECT 59.840 162.770 60.500 162.910 ;
        RECT 59.840 162.680 60.100 162.770 ;
        RECT 54.320 161.660 54.580 161.980 ;
        RECT 58.060 161.640 58.200 162.680 ;
        RECT 58.000 161.320 58.260 161.640 ;
        RECT 53.400 160.980 53.660 161.300 ;
        RECT 53.460 149.740 53.600 160.980 ;
        RECT 57.080 158.600 57.340 158.920 ;
        RECT 57.140 156.200 57.280 158.600 ;
        RECT 58.060 158.240 58.200 161.320 ;
        RECT 60.360 160.960 60.500 162.770 ;
        RECT 62.140 162.680 62.400 163.000 ;
        RECT 62.200 161.980 62.340 162.680 ;
        RECT 64.500 161.980 64.640 166.420 ;
        RECT 65.820 165.400 66.080 165.720 ;
        RECT 65.880 164.020 66.020 165.400 ;
        RECT 65.820 163.700 66.080 164.020 ;
        RECT 62.140 161.660 62.400 161.980 ;
        RECT 64.440 161.660 64.700 161.980 ;
        RECT 61.220 160.980 61.480 161.300 ;
        RECT 59.840 160.640 60.100 160.960 ;
        RECT 60.300 160.640 60.560 160.960 ;
        RECT 58.460 158.600 58.720 158.920 ;
        RECT 58.000 157.920 58.260 158.240 ;
        RECT 57.540 157.580 57.800 157.900 ;
        RECT 57.080 155.880 57.340 156.200 ;
        RECT 54.780 152.480 55.040 152.800 ;
        RECT 56.620 152.480 56.880 152.800 ;
        RECT 53.400 149.420 53.660 149.740 ;
        RECT 53.400 148.060 53.660 148.380 ;
        RECT 52.940 147.380 53.200 147.700 ;
        RECT 53.460 145.320 53.600 148.060 ;
        RECT 54.840 148.040 54.980 152.480 ;
        RECT 55.700 151.800 55.960 152.120 ;
        RECT 55.760 148.380 55.900 151.800 ;
        RECT 55.700 148.060 55.960 148.380 ;
        RECT 54.320 147.720 54.580 148.040 ;
        RECT 54.780 147.720 55.040 148.040 ;
        RECT 53.400 145.000 53.660 145.320 ;
        RECT 54.380 145.060 54.520 147.720 ;
        RECT 54.840 145.660 54.980 147.720 ;
        RECT 55.760 147.360 55.900 148.060 ;
        RECT 56.680 147.360 56.820 152.480 ;
        RECT 57.600 152.460 57.740 157.580 ;
        RECT 58.520 155.260 58.660 158.600 ;
        RECT 59.900 158.580 60.040 160.640 ;
        RECT 59.840 158.260 60.100 158.580 ;
        RECT 59.380 157.920 59.640 158.240 ;
        RECT 58.060 155.120 58.660 155.260 ;
        RECT 58.060 154.840 58.200 155.120 ;
        RECT 58.000 154.520 58.260 154.840 ;
        RECT 57.540 152.140 57.800 152.460 ;
        RECT 57.540 147.610 57.800 147.700 ;
        RECT 58.060 147.610 58.200 154.520 ;
        RECT 58.460 152.480 58.720 152.800 ;
        RECT 58.520 150.760 58.660 152.480 ;
        RECT 58.460 150.440 58.720 150.760 ;
        RECT 58.520 148.040 58.660 150.440 ;
        RECT 58.920 150.100 59.180 150.420 ;
        RECT 58.460 147.720 58.720 148.040 ;
        RECT 57.540 147.470 58.200 147.610 ;
        RECT 57.540 147.380 57.800 147.470 ;
        RECT 55.700 147.040 55.960 147.360 ;
        RECT 56.620 147.040 56.880 147.360 ;
        RECT 55.760 146.680 55.900 147.040 ;
        RECT 55.700 146.360 55.960 146.680 ;
        RECT 54.780 145.340 55.040 145.660 ;
        RECT 54.380 144.920 54.980 145.060 ;
        RECT 53.400 139.220 53.660 139.540 ;
        RECT 53.460 137.500 53.600 139.220 ;
        RECT 53.860 138.880 54.120 139.200 ;
        RECT 52.480 137.180 52.740 137.500 ;
        RECT 53.400 137.180 53.660 137.500 ;
        RECT 51.560 136.500 51.820 136.820 ;
        RECT 51.100 136.160 51.360 136.480 ;
        RECT 51.160 133.500 51.300 136.160 ;
        RECT 51.620 134.780 51.760 136.500 ;
        RECT 53.460 136.480 53.600 137.180 ;
        RECT 52.020 136.160 52.280 136.480 ;
        RECT 53.400 136.160 53.660 136.480 ;
        RECT 52.080 134.780 52.220 136.160 ;
        RECT 52.940 135.820 53.200 136.140 ;
        RECT 51.560 134.460 51.820 134.780 ;
        RECT 52.020 134.460 52.280 134.780 ;
        RECT 53.000 133.760 53.140 135.820 ;
        RECT 51.160 133.360 51.760 133.500 ;
        RECT 52.940 133.440 53.200 133.760 ;
        RECT 51.100 132.760 51.360 133.080 ;
        RECT 51.160 128.660 51.300 132.760 ;
        RECT 51.620 132.140 51.760 133.360 ;
        RECT 51.620 132.000 52.220 132.140 ;
        RECT 51.560 131.060 51.820 131.380 ;
        RECT 51.100 128.340 51.360 128.660 ;
        RECT 51.620 125.940 51.760 131.060 ;
        RECT 52.080 131.040 52.220 132.000 ;
        RECT 52.020 130.720 52.280 131.040 ;
        RECT 51.560 125.620 51.820 125.940 ;
        RECT 52.080 120.500 52.220 130.720 ;
        RECT 52.480 130.380 52.740 130.700 ;
        RECT 52.540 124.920 52.680 130.380 ;
        RECT 53.000 130.360 53.140 133.440 ;
        RECT 53.920 130.700 54.060 138.880 ;
        RECT 53.860 130.380 54.120 130.700 ;
        RECT 52.940 130.040 53.200 130.360 ;
        RECT 53.000 129.340 53.140 130.040 ;
        RECT 52.940 129.020 53.200 129.340 ;
        RECT 52.480 124.600 52.740 124.920 ;
        RECT 54.320 124.600 54.580 124.920 ;
        RECT 52.540 123.900 52.680 124.600 ;
        RECT 52.480 123.580 52.740 123.900 ;
        RECT 53.400 123.240 53.660 123.560 ;
        RECT 53.460 121.180 53.600 123.240 ;
        RECT 53.400 120.860 53.660 121.180 ;
        RECT 52.020 120.180 52.280 120.500 ;
        RECT 54.380 120.160 54.520 124.600 ;
        RECT 54.320 119.840 54.580 120.160 ;
        RECT 54.840 115.400 54.980 144.920 ;
        RECT 55.240 144.660 55.500 144.980 ;
        RECT 55.760 144.890 55.900 146.360 ;
        RECT 56.160 144.890 56.420 144.980 ;
        RECT 55.760 144.750 56.420 144.890 ;
        RECT 56.160 144.660 56.420 144.750 ;
        RECT 56.680 144.890 56.820 147.040 ;
        RECT 57.600 145.660 57.740 147.380 ;
        RECT 58.520 147.360 58.660 147.720 ;
        RECT 58.460 147.040 58.720 147.360 ;
        RECT 58.980 147.100 59.120 150.100 ;
        RECT 59.440 149.400 59.580 157.920 ;
        RECT 59.900 154.840 60.040 158.260 ;
        RECT 60.360 157.900 60.500 160.640 ;
        RECT 61.280 157.900 61.420 160.980 ;
        RECT 66.280 159.960 66.540 160.280 ;
        RECT 61.880 159.425 63.760 159.795 ;
        RECT 62.600 158.260 62.860 158.580 ;
        RECT 60.300 157.580 60.560 157.900 ;
        RECT 61.220 157.580 61.480 157.900 ;
        RECT 62.660 155.860 62.800 158.260 ;
        RECT 66.340 157.900 66.480 159.960 ;
        RECT 63.980 157.580 64.240 157.900 ;
        RECT 66.280 157.580 66.540 157.900 ;
        RECT 62.600 155.540 62.860 155.860 ;
        RECT 59.840 154.520 60.100 154.840 ;
        RECT 59.900 153.480 60.040 154.520 ;
        RECT 61.880 153.985 63.760 154.355 ;
        RECT 59.840 153.160 60.100 153.480 ;
        RECT 59.380 149.080 59.640 149.400 ;
        RECT 58.980 146.960 59.580 147.100 ;
        RECT 57.540 145.340 57.800 145.660 ;
        RECT 57.080 144.890 57.340 144.980 ;
        RECT 56.680 144.750 57.340 144.890 ;
        RECT 55.300 144.380 55.440 144.660 ;
        RECT 56.680 144.380 56.820 144.750 ;
        RECT 57.080 144.660 57.340 144.750 ;
        RECT 55.300 144.240 56.820 144.380 ;
        RECT 57.540 143.980 57.800 144.300 ;
        RECT 55.700 135.480 55.960 135.800 ;
        RECT 55.760 133.760 55.900 135.480 ;
        RECT 57.600 134.780 57.740 143.980 ;
        RECT 57.540 134.460 57.800 134.780 ;
        RECT 56.160 133.780 56.420 134.100 ;
        RECT 55.700 133.440 55.960 133.760 ;
        RECT 55.760 131.380 55.900 133.440 ;
        RECT 56.220 132.060 56.360 133.780 ;
        RECT 56.160 131.740 56.420 132.060 ;
        RECT 55.700 131.060 55.960 131.380 ;
        RECT 57.600 129.340 57.740 134.460 ;
        RECT 57.540 129.020 57.800 129.340 ;
        RECT 57.600 125.600 57.740 129.020 ;
        RECT 58.000 128.000 58.260 128.320 ;
        RECT 57.540 125.280 57.800 125.600 ;
        RECT 58.060 123.220 58.200 128.000 ;
        RECT 58.000 122.900 58.260 123.220 ;
        RECT 56.160 122.560 56.420 122.880 ;
        RECT 56.220 121.180 56.360 122.560 ;
        RECT 56.160 120.860 56.420 121.180 ;
        RECT 58.060 120.500 58.200 122.900 ;
        RECT 58.920 122.560 59.180 122.880 ;
        RECT 58.000 120.180 58.260 120.500 ;
        RECT 58.980 120.160 59.120 122.560 ;
        RECT 58.920 119.840 59.180 120.160 ;
        RECT 54.780 115.080 55.040 115.400 ;
        RECT 50.640 114.740 50.900 115.060 ;
        RECT 49.320 114.320 49.920 114.460 ;
        RECT 50.180 114.400 50.440 114.720 ;
        RECT 46.500 113.720 46.760 114.040 ;
        RECT 49.260 113.720 49.520 114.040 ;
        RECT 43.740 112.700 44.000 113.020 ;
        RECT 46.040 112.700 46.300 113.020 ;
        RECT 40.060 112.020 40.320 112.340 ;
        RECT 42.820 111.680 43.080 112.000 ;
        RECT 42.880 109.620 43.020 111.680 ;
        RECT 42.820 109.300 43.080 109.620 ;
        RECT 38.680 108.960 38.940 109.280 ;
        RECT 38.220 108.280 38.480 108.600 ;
        RECT 33.620 106.580 33.880 106.900 ;
        RECT 31.880 105.025 33.760 105.395 ;
        RECT 32.300 95.280 32.900 95.420 ;
        RECT 32.300 94.740 32.440 95.280 ;
        RECT 32.760 94.980 32.900 95.280 ;
        RECT 38.280 94.980 38.420 108.280 ;
        RECT 43.800 94.980 43.940 112.700 ;
        RECT 46.560 112.680 46.700 113.720 ;
        RECT 46.880 113.185 48.760 113.555 ;
        RECT 46.500 112.360 46.760 112.680 ;
        RECT 49.320 108.940 49.460 113.720 ;
        RECT 49.780 112.340 49.920 114.320 ;
        RECT 57.540 114.060 57.800 114.380 ;
        RECT 57.080 113.720 57.340 114.040 ;
        RECT 57.140 113.020 57.280 113.720 ;
        RECT 54.780 112.700 55.040 113.020 ;
        RECT 57.080 112.700 57.340 113.020 ;
        RECT 53.860 112.360 54.120 112.680 ;
        RECT 49.720 112.020 49.980 112.340 ;
        RECT 53.920 110.300 54.060 112.360 ;
        RECT 53.860 109.980 54.120 110.300 ;
        RECT 49.260 108.620 49.520 108.940 ;
        RECT 49.720 108.280 49.980 108.600 ;
        RECT 46.880 107.745 48.760 108.115 ;
        RECT 49.780 102.220 49.920 108.280 ;
        RECT 49.320 102.080 49.920 102.220 ;
        RECT 49.320 94.980 49.460 102.080 ;
        RECT 54.840 94.980 54.980 112.700 ;
        RECT 57.600 109.280 57.740 114.060 ;
        RECT 59.440 112.680 59.580 146.960 ;
        RECT 59.900 144.640 60.040 153.160 ;
        RECT 64.040 153.140 64.180 157.580 ;
        RECT 64.440 157.240 64.700 157.560 ;
        RECT 64.500 155.860 64.640 157.240 ;
        RECT 68.120 155.880 68.380 156.200 ;
        RECT 64.440 155.540 64.700 155.860 ;
        RECT 66.740 155.540 67.000 155.860 ;
        RECT 66.800 153.820 66.940 155.540 ;
        RECT 68.180 155.180 68.320 155.880 ;
        RECT 68.120 154.860 68.380 155.180 ;
        RECT 68.580 154.520 68.840 154.840 ;
        RECT 66.740 153.500 67.000 153.820 ;
        RECT 62.140 152.820 62.400 153.140 ;
        RECT 63.980 152.820 64.240 153.140 ;
        RECT 65.350 152.965 65.630 153.335 ;
        RECT 68.640 153.140 68.780 154.520 ;
        RECT 65.360 152.820 65.620 152.965 ;
        RECT 68.580 152.820 68.840 153.140 ;
        RECT 62.200 152.460 62.340 152.820 ;
        RECT 62.140 152.140 62.400 152.460 ;
        RECT 65.360 151.800 65.620 152.120 ;
        RECT 61.220 150.100 61.480 150.420 ;
        RECT 61.280 149.400 61.420 150.100 ;
        RECT 61.220 149.080 61.480 149.400 ;
        RECT 61.280 147.360 61.420 149.080 ;
        RECT 61.880 148.545 63.760 148.915 ;
        RECT 61.220 147.040 61.480 147.360 ;
        RECT 65.420 146.680 65.560 151.800 ;
        RECT 67.660 150.780 67.920 151.100 ;
        RECT 67.200 149.080 67.460 149.400 ;
        RECT 67.260 147.360 67.400 149.080 ;
        RECT 67.200 147.040 67.460 147.360 ;
        RECT 60.760 146.360 61.020 146.680 ;
        RECT 65.360 146.360 65.620 146.680 ;
        RECT 59.840 144.320 60.100 144.640 ;
        RECT 60.300 144.320 60.560 144.640 ;
        RECT 59.900 133.760 60.040 144.320 ;
        RECT 60.360 141.240 60.500 144.320 ;
        RECT 60.820 141.580 60.960 146.360 ;
        RECT 65.420 145.660 65.560 146.360 ;
        RECT 65.360 145.340 65.620 145.660 ;
        RECT 67.200 145.000 67.460 145.320 ;
        RECT 66.740 144.660 67.000 144.980 ;
        RECT 61.220 143.640 61.480 143.960 ;
        RECT 64.440 143.640 64.700 143.960 ;
        RECT 60.760 141.260 61.020 141.580 ;
        RECT 60.300 140.920 60.560 141.240 ;
        RECT 60.360 134.100 60.500 140.920 ;
        RECT 61.280 139.540 61.420 143.640 ;
        RECT 61.880 143.105 63.760 143.475 ;
        RECT 64.500 142.260 64.640 143.640 ;
        RECT 64.440 141.940 64.700 142.260 ;
        RECT 63.520 141.600 63.780 141.920 ;
        RECT 63.980 141.600 64.240 141.920 ;
        RECT 63.580 140.220 63.720 141.600 ;
        RECT 63.520 139.900 63.780 140.220 ;
        RECT 61.220 139.220 61.480 139.540 ;
        RECT 61.880 137.665 63.760 138.035 ;
        RECT 60.300 133.780 60.560 134.100 ;
        RECT 59.840 133.440 60.100 133.760 ;
        RECT 59.900 131.720 60.040 133.440 ;
        RECT 61.220 132.760 61.480 133.080 ;
        RECT 59.840 131.400 60.100 131.720 ;
        RECT 61.280 131.380 61.420 132.760 ;
        RECT 61.880 132.225 63.760 132.595 ;
        RECT 63.520 131.400 63.780 131.720 ;
        RECT 61.220 131.060 61.480 131.380 ;
        RECT 60.760 130.040 61.020 130.360 ;
        RECT 60.820 128.660 60.960 130.040 ;
        RECT 60.760 128.340 61.020 128.660 ;
        RECT 63.580 128.060 63.720 131.400 ;
        RECT 64.040 131.040 64.180 141.600 ;
        RECT 64.500 140.220 64.640 141.940 ;
        RECT 64.440 139.900 64.700 140.220 ;
        RECT 65.820 136.160 66.080 136.480 ;
        RECT 65.880 134.100 66.020 136.160 ;
        RECT 65.820 133.780 66.080 134.100 ;
        RECT 66.800 131.040 66.940 144.660 ;
        RECT 67.260 139.540 67.400 145.000 ;
        RECT 67.720 144.980 67.860 150.780 ;
        RECT 67.660 144.660 67.920 144.980 ;
        RECT 69.560 144.640 69.700 169.820 ;
        RECT 72.260 169.140 72.520 169.460 ;
        RECT 71.800 168.800 72.060 169.120 ;
        RECT 70.880 163.360 71.140 163.680 ;
        RECT 70.410 161.125 70.690 161.495 ;
        RECT 70.420 160.980 70.680 161.125 ;
        RECT 70.940 158.580 71.080 163.360 ;
        RECT 71.860 161.980 72.000 168.800 ;
        RECT 71.800 161.660 72.060 161.980 ;
        RECT 71.340 159.960 71.600 160.280 ;
        RECT 71.800 159.960 72.060 160.280 ;
        RECT 70.420 158.260 70.680 158.580 ;
        RECT 70.880 158.260 71.140 158.580 ;
        RECT 70.480 156.200 70.620 158.260 ;
        RECT 70.420 155.880 70.680 156.200 ;
        RECT 70.880 154.860 71.140 155.180 ;
        RECT 70.940 150.760 71.080 154.860 ;
        RECT 71.400 153.820 71.540 159.960 ;
        RECT 71.340 153.500 71.600 153.820 ;
        RECT 71.400 152.655 71.540 153.500 ;
        RECT 71.330 152.285 71.610 152.655 ;
        RECT 70.880 150.440 71.140 150.760 ;
        RECT 70.420 150.100 70.680 150.420 ;
        RECT 70.480 145.660 70.620 150.100 ;
        RECT 71.860 149.935 72.000 159.960 ;
        RECT 71.790 149.565 72.070 149.935 ;
        RECT 71.860 148.380 72.000 149.565 ;
        RECT 71.800 148.060 72.060 148.380 ;
        RECT 70.420 145.340 70.680 145.660 ;
        RECT 72.320 145.570 72.460 169.140 ;
        RECT 72.780 165.460 72.920 181.720 ;
        RECT 73.640 179.340 73.900 179.660 ;
        RECT 73.180 177.980 73.440 178.300 ;
        RECT 73.240 174.980 73.380 177.980 ;
        RECT 73.700 175.580 73.840 179.340 ;
        RECT 73.640 175.260 73.900 175.580 ;
        RECT 73.240 174.840 73.840 174.980 ;
        RECT 73.180 174.240 73.440 174.560 ;
        RECT 73.240 166.400 73.380 174.240 ;
        RECT 73.700 172.860 73.840 174.840 ;
        RECT 73.640 172.540 73.900 172.860 ;
        RECT 73.640 170.840 73.900 171.160 ;
        RECT 73.180 166.080 73.440 166.400 ;
        RECT 72.780 165.320 73.380 165.460 ;
        RECT 73.240 158.660 73.380 165.320 ;
        RECT 73.700 159.340 73.840 170.840 ;
        RECT 74.160 167.080 74.300 184.440 ;
        RECT 74.620 182.380 74.760 185.040 ;
        RECT 75.020 183.080 75.280 183.400 ;
        RECT 74.560 182.060 74.820 182.380 ;
        RECT 74.620 178.300 74.760 182.060 ;
        RECT 75.080 179.320 75.220 183.080 ;
        RECT 75.020 179.000 75.280 179.320 ;
        RECT 75.080 178.300 75.220 179.000 ;
        RECT 74.560 177.980 74.820 178.300 ;
        RECT 75.020 177.980 75.280 178.300 ;
        RECT 74.620 175.580 74.760 177.980 ;
        RECT 75.020 177.300 75.280 177.620 ;
        RECT 74.560 175.260 74.820 175.580 ;
        RECT 74.560 173.900 74.820 174.220 ;
        RECT 74.100 166.760 74.360 167.080 ;
        RECT 74.160 161.495 74.300 166.760 ;
        RECT 74.620 166.740 74.760 173.900 ;
        RECT 75.080 173.880 75.220 177.300 ;
        RECT 75.540 174.560 75.680 192.600 ;
        RECT 76.000 190.200 76.140 195.660 ;
        RECT 76.460 193.940 76.600 196.680 ;
        RECT 79.220 196.320 79.360 198.040 ;
        RECT 79.160 196.000 79.420 196.320 ;
        RECT 76.880 194.785 78.760 195.155 ;
        RECT 81.060 194.620 81.200 198.380 ;
        RECT 80.080 194.300 80.340 194.620 ;
        RECT 81.000 194.300 81.260 194.620 ;
        RECT 80.140 193.940 80.280 194.300 ;
        RECT 76.400 193.620 76.660 193.940 ;
        RECT 80.080 193.620 80.340 193.940 ;
        RECT 76.460 190.540 76.600 193.620 ;
        RECT 81.980 192.920 82.120 198.720 ;
        RECT 82.380 198.040 82.640 198.360 ;
        RECT 98.480 198.040 98.740 198.360 ;
        RECT 82.440 196.660 82.580 198.040 ;
        RECT 91.880 197.505 93.760 197.875 ;
        RECT 86.120 196.660 86.720 196.740 ;
        RECT 82.380 196.340 82.640 196.660 ;
        RECT 86.120 196.600 86.780 196.660 ;
        RECT 86.120 194.620 86.260 196.600 ;
        RECT 86.520 196.340 86.780 196.600 ;
        RECT 88.360 196.230 88.620 196.320 ;
        RECT 88.360 196.090 89.020 196.230 ;
        RECT 88.360 196.000 88.620 196.090 ;
        RECT 86.520 195.320 86.780 195.640 ;
        RECT 86.580 194.620 86.720 195.320 ;
        RECT 86.060 194.300 86.320 194.620 ;
        RECT 86.520 194.300 86.780 194.620 ;
        RECT 84.680 193.620 84.940 193.940 ;
        RECT 77.320 192.600 77.580 192.920 ;
        RECT 81.920 192.600 82.180 192.920 ;
        RECT 77.380 191.900 77.520 192.600 ;
        RECT 77.320 191.580 77.580 191.900 ;
        RECT 81.980 191.220 82.120 192.600 ;
        RECT 84.740 191.900 84.880 193.620 ;
        RECT 88.880 193.600 89.020 196.090 ;
        RECT 98.020 195.320 98.280 195.640 ;
        RECT 98.080 193.940 98.220 195.320 ;
        RECT 98.540 194.280 98.680 198.040 ;
        RECT 100.840 197.340 100.980 199.400 ;
        RECT 110.440 199.060 110.700 199.380 ;
        RECT 105.840 198.720 106.100 199.040 ;
        RECT 109.060 198.720 109.320 199.040 ;
        RECT 105.900 197.340 106.040 198.720 ;
        RECT 100.780 197.020 101.040 197.340 ;
        RECT 105.840 197.020 106.100 197.340 ;
        RECT 103.080 196.000 103.340 196.320 ;
        RECT 103.140 194.620 103.280 196.000 ;
        RECT 106.880 194.785 108.760 195.155 ;
        RECT 103.080 194.300 103.340 194.620 ;
        RECT 98.480 193.960 98.740 194.280 ;
        RECT 90.660 193.620 90.920 193.940 ;
        RECT 96.640 193.620 96.900 193.940 ;
        RECT 98.020 193.620 98.280 193.940 ;
        RECT 88.820 193.280 89.080 193.600 ;
        RECT 84.680 191.580 84.940 191.900 ;
        RECT 81.920 190.900 82.180 191.220 ;
        RECT 76.400 190.220 76.660 190.540 ;
        RECT 75.940 189.880 76.200 190.200 ;
        RECT 81.000 189.880 81.260 190.200 ;
        RECT 86.060 189.880 86.320 190.200 ;
        RECT 76.880 189.345 78.760 189.715 ;
        RECT 81.060 188.840 81.200 189.880 ;
        RECT 81.000 188.520 81.260 188.840 ;
        RECT 85.600 188.520 85.860 188.840 ;
        RECT 85.140 187.840 85.400 188.160 ;
        RECT 85.200 185.780 85.340 187.840 ;
        RECT 85.140 185.460 85.400 185.780 ;
        RECT 76.400 184.780 76.660 185.100 ;
        RECT 83.760 184.780 84.020 185.100 ;
        RECT 76.460 183.740 76.600 184.780 ;
        RECT 76.880 183.905 78.760 184.275 ;
        RECT 83.820 183.740 83.960 184.780 ;
        RECT 85.660 184.760 85.800 188.520 ;
        RECT 86.120 188.160 86.260 189.880 ;
        RECT 86.060 187.840 86.320 188.160 ;
        RECT 85.600 184.440 85.860 184.760 ;
        RECT 76.400 183.420 76.660 183.740 ;
        RECT 83.760 183.420 84.020 183.740 ;
        RECT 84.220 183.420 84.480 183.740 ;
        RECT 79.160 182.740 79.420 183.060 ;
        RECT 76.400 182.060 76.660 182.380 ;
        RECT 75.940 176.620 76.200 176.940 ;
        RECT 76.000 175.095 76.140 176.620 ;
        RECT 75.930 174.725 76.210 175.095 ;
        RECT 75.480 174.240 75.740 174.560 ;
        RECT 75.020 173.560 75.280 173.880 ;
        RECT 75.080 169.120 75.220 173.560 ;
        RECT 75.540 172.180 75.680 174.240 ;
        RECT 75.480 171.860 75.740 172.180 ;
        RECT 75.020 168.800 75.280 169.120 ;
        RECT 74.560 166.420 74.820 166.740 ;
        RECT 74.620 163.680 74.760 166.420 ;
        RECT 75.080 165.720 75.220 168.800 ;
        RECT 75.480 168.460 75.740 168.780 ;
        RECT 75.540 166.060 75.680 168.460 ;
        RECT 76.460 168.440 76.600 182.060 ;
        RECT 76.880 178.465 78.760 178.835 ;
        RECT 78.700 176.280 78.960 176.600 ;
        RECT 78.760 174.900 78.900 176.280 ;
        RECT 78.700 174.580 78.960 174.900 ;
        RECT 79.220 174.560 79.360 182.740 ;
        RECT 81.460 180.700 81.720 181.020 ;
        RECT 81.520 180.340 81.660 180.700 ;
        RECT 81.460 180.020 81.720 180.340 ;
        RECT 80.540 179.680 80.800 180.000 ;
        RECT 80.600 177.530 80.740 179.680 ;
        RECT 81.520 178.300 81.660 180.020 ;
        RECT 82.380 179.000 82.640 179.320 ;
        RECT 81.460 177.980 81.720 178.300 ;
        RECT 81.520 177.620 81.660 177.980 ;
        RECT 81.000 177.530 81.260 177.620 ;
        RECT 80.600 177.390 81.260 177.530 ;
        RECT 81.000 177.300 81.260 177.390 ;
        RECT 81.460 177.300 81.720 177.620 ;
        RECT 81.920 177.300 82.180 177.620 ;
        RECT 81.060 177.135 81.200 177.300 ;
        RECT 80.990 176.765 81.270 177.135 ;
        RECT 79.620 176.280 79.880 176.600 ;
        RECT 79.160 174.240 79.420 174.560 ;
        RECT 76.880 173.025 78.760 173.395 ;
        RECT 76.400 168.120 76.660 168.440 ;
        RECT 75.940 166.080 76.200 166.400 ;
        RECT 75.480 165.740 75.740 166.060 ;
        RECT 75.020 165.400 75.280 165.720 ;
        RECT 74.560 163.360 74.820 163.680 ;
        RECT 74.620 161.640 74.760 163.360 ;
        RECT 75.080 163.340 75.220 165.400 ;
        RECT 75.020 163.020 75.280 163.340 ;
        RECT 74.090 161.125 74.370 161.495 ;
        RECT 74.560 161.320 74.820 161.640 ;
        RECT 75.080 161.300 75.220 163.020 ;
        RECT 74.100 160.980 74.360 161.125 ;
        RECT 75.020 160.980 75.280 161.300 ;
        RECT 73.700 159.260 74.300 159.340 ;
        RECT 73.640 159.200 74.300 159.260 ;
        RECT 73.640 158.940 73.900 159.200 ;
        RECT 73.240 158.520 73.840 158.660 ;
        RECT 73.700 158.240 73.840 158.520 ;
        RECT 73.640 157.920 73.900 158.240 ;
        RECT 73.700 155.860 73.840 157.920 ;
        RECT 73.640 155.540 73.900 155.860 ;
        RECT 72.720 154.860 72.980 155.180 ;
        RECT 72.780 151.100 72.920 154.860 ;
        RECT 73.180 152.480 73.440 152.800 ;
        RECT 72.720 150.780 72.980 151.100 ;
        RECT 73.240 150.420 73.380 152.480 ;
        RECT 73.700 150.420 73.840 155.540 ;
        RECT 74.160 153.140 74.300 159.200 ;
        RECT 75.080 158.240 75.220 160.980 ;
        RECT 76.000 160.140 76.140 166.080 ;
        RECT 75.540 160.000 76.140 160.140 ;
        RECT 75.540 158.580 75.680 160.000 ;
        RECT 75.480 158.260 75.740 158.580 ;
        RECT 75.020 157.920 75.280 158.240 ;
        RECT 74.560 157.240 74.820 157.560 ;
        RECT 74.620 156.200 74.760 157.240 ;
        RECT 74.560 155.880 74.820 156.200 ;
        RECT 75.080 155.860 75.220 157.920 ;
        RECT 75.020 155.540 75.280 155.860 ;
        RECT 75.540 155.260 75.680 158.260 ;
        RECT 76.460 157.980 76.600 168.120 ;
        RECT 76.880 167.585 78.760 167.955 ;
        RECT 79.160 162.680 79.420 163.000 ;
        RECT 76.880 162.145 78.760 162.515 ;
        RECT 79.220 161.300 79.360 162.680 ;
        RECT 79.160 161.210 79.420 161.300 ;
        RECT 78.760 161.070 79.420 161.210 ;
        RECT 76.860 159.960 77.120 160.280 ;
        RECT 76.920 158.920 77.060 159.960 ;
        RECT 76.860 158.600 77.120 158.920 ;
        RECT 78.760 158.240 78.900 161.070 ;
        RECT 79.160 160.980 79.420 161.070 ;
        RECT 79.160 160.300 79.420 160.620 ;
        RECT 79.220 159.260 79.360 160.300 ;
        RECT 79.160 158.940 79.420 159.260 ;
        RECT 79.220 158.240 79.360 158.940 ;
        RECT 75.080 155.120 75.680 155.260 ;
        RECT 76.000 157.840 76.600 157.980 ;
        RECT 78.700 157.920 78.960 158.240 ;
        RECT 79.160 157.920 79.420 158.240 ;
        RECT 74.100 152.820 74.360 153.140 ;
        RECT 74.100 152.140 74.360 152.460 ;
        RECT 73.180 150.100 73.440 150.420 ;
        RECT 73.640 150.100 73.900 150.420 ;
        RECT 73.640 149.420 73.900 149.740 ;
        RECT 72.720 149.080 72.980 149.400 ;
        RECT 72.780 147.700 72.920 149.080 ;
        RECT 72.720 147.380 72.980 147.700 ;
        RECT 72.320 145.430 72.920 145.570 ;
        RECT 69.960 144.660 70.220 144.980 ;
        RECT 72.260 144.660 72.520 144.980 ;
        RECT 68.120 144.320 68.380 144.640 ;
        RECT 69.500 144.320 69.760 144.640 ;
        RECT 68.180 142.940 68.320 144.320 ;
        RECT 68.120 142.620 68.380 142.940 ;
        RECT 68.180 139.540 68.320 142.620 ;
        RECT 69.560 139.540 69.700 144.320 ;
        RECT 70.020 142.260 70.160 144.660 ;
        RECT 70.880 143.980 71.140 144.300 ;
        RECT 69.960 141.940 70.220 142.260 ;
        RECT 70.020 139.540 70.160 141.940 ;
        RECT 70.940 139.880 71.080 143.980 ;
        RECT 71.800 143.640 72.060 143.960 ;
        RECT 71.860 141.580 72.000 143.640 ;
        RECT 71.800 141.260 72.060 141.580 ;
        RECT 70.880 139.560 71.140 139.880 ;
        RECT 67.200 139.220 67.460 139.540 ;
        RECT 68.120 139.220 68.380 139.540 ;
        RECT 69.500 139.220 69.760 139.540 ;
        RECT 69.960 139.220 70.220 139.540 ;
        RECT 67.260 137.160 67.400 139.220 ;
        RECT 67.200 136.840 67.460 137.160 ;
        RECT 68.180 136.820 68.320 139.220 ;
        RECT 68.120 136.500 68.380 136.820 ;
        RECT 68.180 134.780 68.320 136.500 ;
        RECT 69.560 136.480 69.700 139.220 ;
        RECT 69.500 136.160 69.760 136.480 ;
        RECT 68.580 135.820 68.840 136.140 ;
        RECT 68.120 134.460 68.380 134.780 ;
        RECT 67.200 133.780 67.460 134.100 ;
        RECT 63.980 130.720 64.240 131.040 ;
        RECT 66.740 130.720 67.000 131.040 ;
        RECT 64.040 128.660 64.180 130.720 ;
        RECT 66.800 129.340 66.940 130.720 ;
        RECT 67.260 130.360 67.400 133.780 ;
        RECT 67.200 130.040 67.460 130.360 ;
        RECT 66.740 129.020 67.000 129.340 ;
        RECT 63.980 128.340 64.240 128.660 ;
        RECT 63.580 127.920 64.180 128.060 ;
        RECT 61.880 126.785 63.760 127.155 ;
        RECT 64.040 125.940 64.180 127.920 ;
        RECT 63.980 125.620 64.240 125.940 ;
        RECT 67.260 124.920 67.400 130.040 ;
        RECT 68.640 124.920 68.780 135.820 ;
        RECT 69.560 134.100 69.700 136.160 ;
        RECT 69.500 133.780 69.760 134.100 ;
        RECT 70.880 128.680 71.140 129.000 ;
        RECT 70.420 128.340 70.680 128.660 ;
        RECT 70.480 125.940 70.620 128.340 ;
        RECT 70.420 125.620 70.680 125.940 ;
        RECT 64.900 124.600 65.160 124.920 ;
        RECT 67.200 124.600 67.460 124.920 ;
        RECT 68.580 124.600 68.840 124.920 ;
        RECT 64.960 123.220 65.100 124.600 ;
        RECT 67.260 123.900 67.400 124.600 ;
        RECT 67.200 123.580 67.460 123.900 ;
        RECT 64.900 122.900 65.160 123.220 ;
        RECT 63.980 121.880 64.240 122.200 ;
        RECT 64.440 121.880 64.700 122.200 ;
        RECT 61.880 121.345 63.760 121.715 ;
        RECT 64.040 121.090 64.180 121.880 ;
        RECT 63.580 120.950 64.180 121.090 ;
        RECT 60.300 119.840 60.560 120.160 ;
        RECT 59.380 112.360 59.640 112.680 ;
        RECT 60.360 112.000 60.500 119.840 ;
        RECT 63.580 119.820 63.720 120.950 ;
        RECT 64.500 120.500 64.640 121.880 ;
        RECT 68.640 121.180 68.780 124.600 ;
        RECT 69.500 123.240 69.760 123.560 ;
        RECT 69.560 121.180 69.700 123.240 ;
        RECT 70.480 122.880 70.620 125.620 ;
        RECT 70.940 125.600 71.080 128.680 ;
        RECT 72.320 125.600 72.460 144.660 ;
        RECT 72.780 131.380 72.920 145.430 ;
        RECT 73.700 142.940 73.840 149.420 ;
        RECT 74.160 147.215 74.300 152.140 ;
        RECT 74.560 149.080 74.820 149.400 ;
        RECT 74.090 146.845 74.370 147.215 ;
        RECT 74.620 145.320 74.760 149.080 ;
        RECT 74.560 145.000 74.820 145.320 ;
        RECT 73.640 142.620 73.900 142.940 ;
        RECT 74.620 142.260 74.760 145.000 ;
        RECT 74.560 141.940 74.820 142.260 ;
        RECT 73.640 141.600 73.900 141.920 ;
        RECT 73.700 140.220 73.840 141.600 ;
        RECT 73.640 139.900 73.900 140.220 ;
        RECT 75.080 139.200 75.220 155.120 ;
        RECT 75.480 147.040 75.740 147.360 ;
        RECT 75.540 142.260 75.680 147.040 ;
        RECT 76.000 144.980 76.140 157.840 ;
        RECT 76.400 157.240 76.660 157.560 ;
        RECT 76.460 150.420 76.600 157.240 ;
        RECT 76.880 156.705 78.760 157.075 ;
        RECT 79.160 153.500 79.420 153.820 ;
        RECT 76.880 151.265 78.760 151.635 ;
        RECT 76.400 150.100 76.660 150.420 ;
        RECT 76.880 145.825 78.760 146.195 ;
        RECT 75.940 144.660 76.200 144.980 ;
        RECT 76.400 144.320 76.660 144.640 ;
        RECT 75.480 141.940 75.740 142.260 ;
        RECT 75.020 138.880 75.280 139.200 ;
        RECT 73.630 136.645 73.910 137.015 ;
        RECT 73.700 136.480 73.840 136.645 ;
        RECT 73.640 136.390 73.900 136.480 ;
        RECT 73.240 136.250 73.900 136.390 ;
        RECT 73.240 134.440 73.380 136.250 ;
        RECT 73.640 136.160 73.900 136.250 ;
        RECT 73.640 135.480 73.900 135.800 ;
        RECT 73.180 134.120 73.440 134.440 ;
        RECT 73.700 133.080 73.840 135.480 ;
        RECT 75.080 133.760 75.220 138.880 ;
        RECT 75.020 133.440 75.280 133.760 ;
        RECT 73.640 132.760 73.900 133.080 ;
        RECT 72.720 131.060 72.980 131.380 ;
        RECT 73.700 131.040 73.840 132.760 ;
        RECT 73.640 130.720 73.900 131.040 ;
        RECT 72.720 130.040 72.980 130.360 ;
        RECT 74.560 130.040 74.820 130.360 ;
        RECT 72.780 125.600 72.920 130.040 ;
        RECT 73.640 128.000 73.900 128.320 ;
        RECT 73.700 126.620 73.840 128.000 ;
        RECT 73.640 126.300 73.900 126.620 ;
        RECT 74.620 125.600 74.760 130.040 ;
        RECT 70.880 125.280 71.140 125.600 ;
        RECT 72.260 125.280 72.520 125.600 ;
        RECT 72.720 125.280 72.980 125.600 ;
        RECT 74.560 125.280 74.820 125.600 ;
        RECT 71.340 124.600 71.600 124.920 ;
        RECT 70.420 122.560 70.680 122.880 ;
        RECT 68.580 120.860 68.840 121.180 ;
        RECT 69.500 120.860 69.760 121.180 ;
        RECT 64.440 120.180 64.700 120.500 ;
        RECT 70.480 120.160 70.620 122.560 ;
        RECT 71.400 120.160 71.540 124.600 ;
        RECT 73.180 122.560 73.440 122.880 ;
        RECT 73.240 121.180 73.380 122.560 ;
        RECT 73.180 120.860 73.440 121.180 ;
        RECT 70.420 119.840 70.680 120.160 ;
        RECT 71.340 119.840 71.600 120.160 ;
        RECT 63.520 119.500 63.780 119.820 ;
        RECT 61.880 115.905 63.760 116.275 ;
        RECT 70.480 115.740 70.620 119.840 ;
        RECT 70.420 115.420 70.680 115.740 ;
        RECT 64.900 114.740 65.160 115.060 ;
        RECT 64.960 112.340 65.100 114.740 ;
        RECT 70.480 114.720 70.620 115.420 ;
        RECT 75.080 115.060 75.220 133.440 ;
        RECT 75.540 128.320 75.680 141.940 ;
        RECT 76.460 139.880 76.600 144.320 ;
        RECT 76.880 140.385 78.760 140.755 ;
        RECT 76.400 139.560 76.660 139.880 ;
        RECT 79.220 137.500 79.360 153.500 ;
        RECT 79.680 150.420 79.820 176.280 ;
        RECT 81.060 174.560 81.200 176.765 ;
        RECT 81.520 174.900 81.660 177.300 ;
        RECT 81.980 175.580 82.120 177.300 ;
        RECT 81.920 175.260 82.180 175.580 ;
        RECT 81.460 174.580 81.720 174.900 ;
        RECT 81.000 174.240 81.260 174.560 ;
        RECT 81.910 174.045 82.190 174.415 ;
        RECT 81.920 173.900 82.180 174.045 ;
        RECT 80.080 168.800 80.340 169.120 ;
        RECT 80.140 165.720 80.280 168.800 ;
        RECT 80.080 165.400 80.340 165.720 ;
        RECT 80.140 158.240 80.280 165.400 ;
        RECT 81.920 159.960 82.180 160.280 ;
        RECT 80.080 157.920 80.340 158.240 ;
        RECT 81.000 157.240 81.260 157.560 ;
        RECT 81.060 152.800 81.200 157.240 ;
        RECT 81.460 155.880 81.720 156.200 ;
        RECT 81.000 152.480 81.260 152.800 ;
        RECT 80.540 152.140 80.800 152.460 ;
        RECT 80.080 151.800 80.340 152.120 ;
        RECT 79.620 150.100 79.880 150.420 ;
        RECT 79.160 137.180 79.420 137.500 ;
        RECT 78.700 136.390 78.960 136.480 ;
        RECT 78.700 136.250 79.360 136.390 ;
        RECT 78.700 136.160 78.960 136.250 ;
        RECT 76.880 134.945 78.760 135.315 ;
        RECT 76.860 134.120 77.120 134.440 ;
        RECT 76.920 132.060 77.060 134.120 ;
        RECT 79.220 133.080 79.360 136.250 ;
        RECT 79.160 132.760 79.420 133.080 ;
        RECT 76.860 131.740 77.120 132.060 ;
        RECT 76.400 130.720 76.660 131.040 ;
        RECT 75.480 128.000 75.740 128.320 ;
        RECT 75.540 123.220 75.680 128.000 ;
        RECT 76.460 125.600 76.600 130.720 ;
        RECT 76.880 129.505 78.760 129.875 ;
        RECT 79.620 128.855 79.880 129.000 ;
        RECT 79.610 128.485 79.890 128.855 ;
        RECT 76.400 125.510 76.660 125.600 ;
        RECT 76.000 125.370 76.660 125.510 ;
        RECT 76.000 123.900 76.140 125.370 ;
        RECT 76.400 125.280 76.660 125.370 ;
        RECT 76.400 124.600 76.660 124.920 ;
        RECT 79.620 124.600 79.880 124.920 ;
        RECT 75.940 123.580 76.200 123.900 ;
        RECT 76.460 123.220 76.600 124.600 ;
        RECT 76.880 124.065 78.760 124.435 ;
        RECT 79.680 123.560 79.820 124.600 ;
        RECT 79.620 123.240 79.880 123.560 ;
        RECT 75.480 122.900 75.740 123.220 ;
        RECT 76.400 122.900 76.660 123.220 ;
        RECT 75.020 114.740 75.280 115.060 ;
        RECT 70.420 114.400 70.680 114.720 ;
        RECT 73.640 113.720 73.900 114.040 ;
        RECT 73.700 112.680 73.840 113.720 ;
        RECT 73.640 112.360 73.900 112.680 ;
        RECT 75.540 112.340 75.680 122.900 ;
        RECT 76.880 118.625 78.760 118.995 ;
        RECT 79.620 114.400 79.880 114.720 ;
        RECT 80.140 114.630 80.280 151.800 ;
        RECT 80.600 150.080 80.740 152.140 ;
        RECT 80.540 149.760 80.800 150.080 ;
        RECT 80.540 149.080 80.800 149.400 ;
        RECT 81.520 149.140 81.660 155.880 ;
        RECT 80.600 137.500 80.740 149.080 ;
        RECT 81.060 149.000 81.660 149.140 ;
        RECT 81.060 141.920 81.200 149.000 ;
        RECT 81.980 147.360 82.120 159.960 ;
        RECT 82.440 147.700 82.580 179.000 ;
        RECT 82.840 176.620 83.100 176.940 ;
        RECT 83.300 176.620 83.560 176.940 ;
        RECT 83.760 176.620 84.020 176.940 ;
        RECT 82.900 174.220 83.040 176.620 ;
        RECT 82.840 173.900 83.100 174.220 ;
        RECT 82.840 170.840 83.100 171.160 ;
        RECT 82.900 169.800 83.040 170.840 ;
        RECT 82.840 169.480 83.100 169.800 ;
        RECT 82.900 164.020 83.040 169.480 ;
        RECT 82.840 163.700 83.100 164.020 ;
        RECT 82.840 160.980 83.100 161.300 ;
        RECT 82.900 159.260 83.040 160.980 ;
        RECT 82.840 158.940 83.100 159.260 ;
        RECT 82.900 158.240 83.040 158.940 ;
        RECT 82.840 157.920 83.100 158.240 ;
        RECT 82.840 157.240 83.100 157.560 ;
        RECT 82.900 155.860 83.040 157.240 ;
        RECT 82.840 155.540 83.100 155.860 ;
        RECT 83.360 153.140 83.500 176.620 ;
        RECT 83.820 175.775 83.960 176.620 ;
        RECT 83.750 175.405 84.030 175.775 ;
        RECT 84.280 174.560 84.420 183.420 ;
        RECT 85.660 182.720 85.800 184.440 ;
        RECT 85.600 182.400 85.860 182.720 ;
        RECT 85.660 180.000 85.800 182.400 ;
        RECT 85.600 179.680 85.860 180.000 ;
        RECT 85.600 175.490 85.860 175.580 ;
        RECT 86.120 175.490 86.260 187.840 ;
        RECT 88.880 185.780 89.020 193.280 ;
        RECT 89.280 192.600 89.540 192.920 ;
        RECT 89.340 190.200 89.480 192.600 ;
        RECT 90.200 190.220 90.460 190.540 ;
        RECT 89.280 189.880 89.540 190.200 ;
        RECT 89.740 187.500 90.000 187.820 ;
        RECT 89.800 185.780 89.940 187.500 ;
        RECT 88.820 185.460 89.080 185.780 ;
        RECT 89.740 185.460 90.000 185.780 ;
        RECT 88.880 184.670 89.020 185.460 ;
        RECT 88.880 184.530 89.480 184.670 ;
        RECT 89.340 182.380 89.480 184.530 ;
        RECT 89.800 182.720 89.940 185.460 ;
        RECT 89.740 182.400 90.000 182.720 ;
        RECT 86.980 182.060 87.240 182.380 ;
        RECT 89.280 182.060 89.540 182.380 ;
        RECT 86.520 179.680 86.780 180.000 ;
        RECT 86.580 177.620 86.720 179.680 ;
        RECT 87.040 177.620 87.180 182.060 ;
        RECT 86.520 177.300 86.780 177.620 ;
        RECT 86.980 177.300 87.240 177.620 ;
        RECT 85.600 175.350 86.260 175.490 ;
        RECT 85.600 175.260 85.860 175.350 ;
        RECT 86.980 175.260 87.240 175.580 ;
        RECT 84.680 174.580 84.940 174.900 ;
        RECT 84.220 174.240 84.480 174.560 ;
        RECT 84.740 172.860 84.880 174.580 ;
        RECT 84.680 172.540 84.940 172.860 ;
        RECT 83.760 172.200 84.020 172.520 ;
        RECT 83.820 169.120 83.960 172.200 ;
        RECT 87.040 171.840 87.180 175.260 ;
        RECT 89.340 174.900 89.480 182.060 ;
        RECT 89.800 181.020 89.940 182.400 ;
        RECT 89.740 180.700 90.000 181.020 ;
        RECT 90.260 177.960 90.400 190.220 ;
        RECT 90.720 188.500 90.860 193.620 ;
        RECT 91.880 192.065 93.760 192.435 ;
        RECT 96.700 191.900 96.840 193.620 ;
        RECT 96.640 191.580 96.900 191.900 ;
        RECT 91.580 190.900 91.840 191.220 ;
        RECT 90.660 188.180 90.920 188.500 ;
        RECT 90.720 179.660 90.860 188.180 ;
        RECT 91.120 187.840 91.380 188.160 ;
        RECT 91.180 185.100 91.320 187.840 ;
        RECT 91.640 187.820 91.780 190.900 ;
        RECT 93.420 190.560 93.680 190.880 ;
        RECT 93.480 189.180 93.620 190.560 ;
        RECT 98.080 190.540 98.220 193.620 ;
        RECT 106.300 192.940 106.560 193.260 ;
        RECT 98.020 190.220 98.280 190.540 ;
        RECT 105.840 189.880 106.100 190.200 ;
        RECT 93.420 188.860 93.680 189.180 ;
        RECT 91.580 187.500 91.840 187.820 ;
        RECT 98.940 187.160 99.200 187.480 ;
        RECT 91.880 186.625 93.760 186.995 ;
        RECT 96.180 185.120 96.440 185.440 ;
        RECT 91.120 184.780 91.380 185.100 ;
        RECT 94.340 184.780 94.600 185.100 ;
        RECT 93.880 184.440 94.140 184.760 ;
        RECT 93.940 183.740 94.080 184.440 ;
        RECT 93.880 183.420 94.140 183.740 ;
        RECT 93.880 181.720 94.140 182.040 ;
        RECT 91.880 181.185 93.760 181.555 ;
        RECT 93.940 180.000 94.080 181.720 ;
        RECT 94.400 181.020 94.540 184.780 ;
        RECT 96.240 182.720 96.380 185.120 ;
        RECT 99.000 184.760 99.140 187.160 ;
        RECT 105.900 185.440 106.040 189.880 ;
        RECT 106.360 185.780 106.500 192.940 ;
        RECT 109.120 191.220 109.260 198.720 ;
        RECT 110.500 196.660 110.640 199.060 ;
        RECT 110.900 198.720 111.160 199.040 ;
        RECT 110.440 196.340 110.700 196.660 ;
        RECT 109.980 196.000 110.240 196.320 ;
        RECT 110.040 194.280 110.180 196.000 ;
        RECT 109.980 193.960 110.240 194.280 ;
        RECT 109.060 190.900 109.320 191.220 ;
        RECT 106.880 189.345 108.760 189.715 ;
        RECT 109.120 188.160 109.260 190.900 ;
        RECT 110.040 189.180 110.180 193.960 ;
        RECT 110.500 193.940 110.640 196.340 ;
        RECT 110.440 193.620 110.700 193.940 ;
        RECT 109.980 188.860 110.240 189.180 ;
        RECT 109.980 188.180 110.240 188.500 ;
        RECT 109.060 187.840 109.320 188.160 ;
        RECT 106.300 185.460 106.560 185.780 ;
        RECT 105.840 185.120 106.100 185.440 ;
        RECT 98.940 184.440 99.200 184.760 ;
        RECT 100.320 184.440 100.580 184.760 ;
        RECT 97.560 183.080 97.820 183.400 ;
        RECT 96.180 182.400 96.440 182.720 ;
        RECT 94.340 180.700 94.600 181.020 ;
        RECT 97.620 180.680 97.760 183.080 ;
        RECT 96.640 180.590 96.900 180.680 ;
        RECT 96.640 180.450 97.300 180.590 ;
        RECT 96.640 180.360 96.900 180.450 ;
        RECT 93.880 179.680 94.140 180.000 ;
        RECT 90.660 179.340 90.920 179.660 ;
        RECT 90.720 177.960 90.860 179.340 ;
        RECT 90.200 177.640 90.460 177.960 ;
        RECT 90.660 177.640 90.920 177.960 ;
        RECT 97.160 177.620 97.300 180.450 ;
        RECT 97.560 180.360 97.820 180.680 ;
        RECT 99.000 177.960 99.140 184.440 ;
        RECT 100.380 180.000 100.520 184.440 ;
        RECT 106.880 183.905 108.760 184.275 ;
        RECT 101.240 183.080 101.500 183.400 ;
        RECT 101.300 181.020 101.440 183.080 ;
        RECT 106.300 182.740 106.560 183.060 ;
        RECT 101.240 180.700 101.500 181.020 ;
        RECT 103.540 180.020 103.800 180.340 ;
        RECT 100.320 179.680 100.580 180.000 ;
        RECT 103.600 179.660 103.740 180.020 ;
        RECT 106.360 180.000 106.500 182.740 ;
        RECT 106.300 179.680 106.560 180.000 ;
        RECT 103.540 179.340 103.800 179.660 ;
        RECT 103.080 179.000 103.340 179.320 ;
        RECT 103.140 177.960 103.280 179.000 ;
        RECT 98.940 177.640 99.200 177.960 ;
        RECT 103.080 177.640 103.340 177.960 ;
        RECT 94.800 177.300 95.060 177.620 ;
        RECT 97.100 177.300 97.360 177.620 ;
        RECT 91.880 175.745 93.760 176.115 ;
        RECT 94.860 174.900 95.000 177.300 ;
        RECT 106.360 177.280 106.500 179.680 ;
        RECT 106.880 178.465 108.760 178.835 ;
        RECT 108.590 177.445 108.870 177.815 ;
        RECT 109.120 177.620 109.260 187.840 ;
        RECT 110.040 186.460 110.180 188.180 ;
        RECT 109.980 186.140 110.240 186.460 ;
        RECT 109.520 185.120 109.780 185.440 ;
        RECT 109.580 180.000 109.720 185.120 ;
        RECT 109.980 182.740 110.240 183.060 ;
        RECT 109.520 179.680 109.780 180.000 ;
        RECT 109.520 179.175 109.780 179.320 ;
        RECT 109.510 178.805 109.790 179.175 ;
        RECT 110.040 177.620 110.180 182.740 ;
        RECT 110.500 177.815 110.640 193.620 ;
        RECT 110.960 193.600 111.100 198.720 ;
        RECT 111.420 194.620 111.560 199.400 ;
        RECT 116.880 199.060 117.140 199.380 ;
        RECT 111.820 198.380 112.080 198.700 ;
        RECT 111.880 194.620 112.020 198.380 ;
        RECT 116.940 194.620 117.080 199.060 ;
        RECT 118.720 198.950 118.980 199.040 ;
        RECT 118.320 198.810 118.980 198.950 ;
        RECT 118.320 196.320 118.460 198.810 ;
        RECT 118.720 198.720 118.980 198.810 ;
        RECT 119.640 198.040 119.900 198.360 ;
        RECT 119.700 196.320 119.840 198.040 ;
        RECT 118.260 196.000 118.520 196.320 ;
        RECT 119.640 196.000 119.900 196.320 ;
        RECT 111.360 194.300 111.620 194.620 ;
        RECT 111.820 194.300 112.080 194.620 ;
        RECT 116.880 194.300 117.140 194.620 ;
        RECT 110.900 193.280 111.160 193.600 ;
        RECT 110.900 182.400 111.160 182.720 ;
        RECT 110.960 180.000 111.100 182.400 ;
        RECT 110.900 179.680 111.160 180.000 ;
        RECT 106.300 176.960 106.560 177.280 ;
        RECT 106.760 176.960 107.020 177.280 ;
        RECT 99.400 176.620 99.660 176.940 ;
        RECT 89.280 174.580 89.540 174.900 ;
        RECT 94.800 174.580 95.060 174.900 ;
        RECT 86.980 171.520 87.240 171.840 ;
        RECT 83.760 168.800 84.020 169.120 ;
        RECT 85.140 168.120 85.400 168.440 ;
        RECT 84.220 165.400 84.480 165.720 ;
        RECT 84.280 163.340 84.420 165.400 ;
        RECT 84.220 163.020 84.480 163.340 ;
        RECT 83.760 157.580 84.020 157.900 ;
        RECT 83.820 156.540 83.960 157.580 ;
        RECT 83.760 156.220 84.020 156.540 ;
        RECT 84.280 155.860 84.420 163.020 ;
        RECT 85.200 163.000 85.340 168.120 ;
        RECT 85.140 162.680 85.400 163.000 ;
        RECT 85.200 161.640 85.340 162.680 ;
        RECT 85.140 161.320 85.400 161.640 ;
        RECT 84.680 160.980 84.940 161.300 ;
        RECT 84.740 158.920 84.880 160.980 ;
        RECT 84.680 158.600 84.940 158.920 ;
        RECT 84.740 158.240 84.880 158.600 ;
        RECT 87.040 158.580 87.180 171.520 ;
        RECT 88.820 170.840 89.080 171.160 ;
        RECT 88.880 167.420 89.020 170.840 ;
        RECT 89.340 168.440 89.480 174.580 ;
        RECT 91.120 173.900 91.380 174.220 ;
        RECT 91.180 172.860 91.320 173.900 ;
        RECT 91.120 172.540 91.380 172.860 ;
        RECT 94.340 171.860 94.600 172.180 ;
        RECT 91.880 170.305 93.760 170.675 ;
        RECT 90.200 169.480 90.460 169.800 ;
        RECT 89.280 168.120 89.540 168.440 ;
        RECT 88.820 167.100 89.080 167.420 ;
        RECT 89.340 166.400 89.480 168.120 ;
        RECT 89.740 166.760 90.000 167.080 ;
        RECT 89.280 166.080 89.540 166.400 ;
        RECT 89.800 164.360 89.940 166.760 ;
        RECT 90.260 166.740 90.400 169.480 ;
        RECT 94.400 169.460 94.540 171.860 ;
        RECT 91.580 169.140 91.840 169.460 ;
        RECT 94.340 169.140 94.600 169.460 ;
        RECT 91.640 166.740 91.780 169.140 ;
        RECT 90.200 166.420 90.460 166.740 ;
        RECT 91.580 166.420 91.840 166.740 ;
        RECT 91.120 165.400 91.380 165.720 ;
        RECT 93.880 165.400 94.140 165.720 ;
        RECT 89.740 164.040 90.000 164.360 ;
        RECT 91.180 163.340 91.320 165.400 ;
        RECT 91.880 164.865 93.760 165.235 ;
        RECT 93.940 164.020 94.080 165.400 ;
        RECT 94.860 164.700 95.000 174.580 ;
        RECT 98.940 174.130 99.200 174.220 ;
        RECT 99.460 174.130 99.600 176.620 ;
        RECT 99.860 176.280 100.120 176.600 ;
        RECT 104.000 176.280 104.260 176.600 ;
        RECT 98.940 173.990 99.600 174.130 ;
        RECT 98.940 173.900 99.200 173.990 ;
        RECT 96.630 172.005 96.910 172.375 ;
        RECT 98.930 172.005 99.210 172.375 ;
        RECT 96.700 169.120 96.840 172.005 ;
        RECT 98.940 171.860 99.200 172.005 ;
        RECT 96.640 168.800 96.900 169.120 ;
        RECT 95.720 166.080 95.980 166.400 ;
        RECT 94.800 164.380 95.060 164.700 ;
        RECT 95.780 164.020 95.920 166.080 ;
        RECT 98.020 165.400 98.280 165.720 ;
        RECT 98.080 164.360 98.220 165.400 ;
        RECT 98.020 164.040 98.280 164.360 ;
        RECT 93.880 163.700 94.140 164.020 ;
        RECT 95.720 163.700 95.980 164.020 ;
        RECT 91.120 163.020 91.380 163.340 ;
        RECT 91.880 159.425 93.760 159.795 ;
        RECT 86.980 158.260 87.240 158.580 ;
        RECT 84.680 157.920 84.940 158.240 ;
        RECT 94.340 157.920 94.600 158.240 ;
        RECT 84.740 155.860 84.880 157.920 ;
        RECT 93.880 157.240 94.140 157.560 ;
        RECT 86.980 156.220 87.240 156.540 ;
        RECT 84.220 155.540 84.480 155.860 ;
        RECT 84.680 155.540 84.940 155.860 ;
        RECT 87.040 154.840 87.180 156.220 ;
        RECT 93.940 156.200 94.080 157.240 ;
        RECT 93.880 155.880 94.140 156.200 ;
        RECT 86.980 154.520 87.240 154.840 ;
        RECT 90.660 154.520 90.920 154.840 ;
        RECT 85.600 153.160 85.860 153.480 ;
        RECT 83.300 152.820 83.560 153.140 ;
        RECT 85.660 152.800 85.800 153.160 ;
        RECT 84.220 152.480 84.480 152.800 ;
        RECT 85.600 152.480 85.860 152.800 ;
        RECT 84.280 151.100 84.420 152.480 ;
        RECT 85.660 151.180 85.800 152.480 ;
        RECT 84.220 150.780 84.480 151.100 ;
        RECT 84.740 151.040 86.260 151.180 ;
        RECT 83.760 149.760 84.020 150.080 ;
        RECT 82.840 148.060 83.100 148.380 ;
        RECT 82.380 147.380 82.640 147.700 ;
        RECT 81.920 147.040 82.180 147.360 ;
        RECT 82.380 146.700 82.640 147.020 ;
        RECT 81.450 145.485 81.730 145.855 ;
        RECT 82.440 145.660 82.580 146.700 ;
        RECT 81.520 142.260 81.660 145.485 ;
        RECT 82.380 145.340 82.640 145.660 ;
        RECT 81.920 143.640 82.180 143.960 ;
        RECT 81.460 141.940 81.720 142.260 ;
        RECT 81.980 141.920 82.120 143.640 ;
        RECT 82.380 142.620 82.640 142.940 ;
        RECT 81.000 141.600 81.260 141.920 ;
        RECT 81.920 141.600 82.180 141.920 ;
        RECT 81.460 140.920 81.720 141.240 ;
        RECT 81.000 138.880 81.260 139.200 ;
        RECT 80.540 137.180 80.800 137.500 ;
        RECT 81.060 130.780 81.200 138.880 ;
        RECT 80.600 130.700 81.200 130.780 ;
        RECT 80.540 130.640 81.200 130.700 ;
        RECT 80.540 130.380 80.800 130.640 ;
        RECT 80.600 126.620 80.740 130.380 ;
        RECT 80.540 126.300 80.800 126.620 ;
        RECT 80.600 120.160 80.740 126.300 ;
        RECT 80.540 119.840 80.800 120.160 ;
        RECT 81.520 115.740 81.660 140.920 ;
        RECT 81.920 139.220 82.180 139.540 ;
        RECT 81.980 136.480 82.120 139.220 ;
        RECT 82.440 137.500 82.580 142.620 ;
        RECT 82.900 139.200 83.040 148.060 ;
        RECT 83.820 145.660 83.960 149.760 ;
        RECT 83.760 145.340 84.020 145.660 ;
        RECT 83.760 144.890 84.020 144.980 ;
        RECT 84.280 144.890 84.420 150.780 ;
        RECT 84.740 150.420 84.880 151.040 ;
        RECT 84.680 150.100 84.940 150.420 ;
        RECT 85.140 150.100 85.400 150.420 ;
        RECT 85.200 144.980 85.340 150.100 ;
        RECT 85.600 146.360 85.860 146.680 ;
        RECT 83.760 144.750 84.420 144.890 ;
        RECT 83.760 144.660 84.020 144.750 ;
        RECT 85.140 144.660 85.400 144.980 ;
        RECT 84.680 143.980 84.940 144.300 ;
        RECT 84.740 142.340 84.880 143.980 ;
        RECT 85.200 142.940 85.340 144.660 ;
        RECT 85.140 142.620 85.400 142.940 ;
        RECT 84.740 142.200 85.340 142.340 ;
        RECT 85.200 141.240 85.340 142.200 ;
        RECT 85.140 140.920 85.400 141.240 ;
        RECT 82.840 138.880 83.100 139.200 ;
        RECT 82.380 137.180 82.640 137.500 ;
        RECT 85.200 137.160 85.340 140.920 ;
        RECT 85.140 136.840 85.400 137.160 ;
        RECT 82.380 136.500 82.640 136.820 ;
        RECT 81.920 136.160 82.180 136.480 ;
        RECT 82.440 130.360 82.580 136.500 ;
        RECT 84.680 136.160 84.940 136.480 ;
        RECT 85.140 136.160 85.400 136.480 ;
        RECT 84.220 132.760 84.480 133.080 ;
        RECT 84.280 131.720 84.420 132.760 ;
        RECT 84.220 131.400 84.480 131.720 ;
        RECT 82.840 130.380 83.100 130.700 ;
        RECT 82.380 130.040 82.640 130.360 ;
        RECT 82.900 120.500 83.040 130.380 ;
        RECT 83.760 130.040 84.020 130.360 ;
        RECT 83.820 123.900 83.960 130.040 ;
        RECT 84.740 125.940 84.880 136.160 ;
        RECT 85.200 132.060 85.340 136.160 ;
        RECT 85.140 131.740 85.400 132.060 ;
        RECT 84.680 125.620 84.940 125.940 ;
        RECT 83.760 123.580 84.020 123.900 ;
        RECT 84.740 120.500 84.880 125.620 ;
        RECT 85.660 123.300 85.800 146.360 ;
        RECT 86.120 144.980 86.260 151.040 ;
        RECT 87.040 150.080 87.180 154.520 ;
        RECT 90.720 153.140 90.860 154.520 ;
        RECT 91.880 153.985 93.760 154.355 ;
        RECT 94.400 153.140 94.540 157.920 ;
        RECT 95.780 155.520 95.920 163.700 ;
        RECT 98.020 156.220 98.280 156.540 ;
        RECT 96.640 155.540 96.900 155.860 ;
        RECT 95.720 155.200 95.980 155.520 ;
        RECT 95.780 153.140 95.920 155.200 ;
        RECT 90.660 152.820 90.920 153.140 ;
        RECT 94.340 152.820 94.600 153.140 ;
        RECT 95.720 152.820 95.980 153.140 ;
        RECT 87.440 152.480 87.700 152.800 ;
        RECT 86.980 149.760 87.240 150.080 ;
        RECT 87.040 149.400 87.180 149.760 ;
        RECT 86.980 149.080 87.240 149.400 ;
        RECT 86.060 144.660 86.320 144.980 ;
        RECT 86.060 142.620 86.320 142.940 ;
        RECT 86.120 142.260 86.260 142.620 ;
        RECT 87.040 142.260 87.180 149.080 ;
        RECT 86.060 141.940 86.320 142.260 ;
        RECT 86.980 141.940 87.240 142.260 ;
        RECT 86.510 141.405 86.790 141.775 ;
        RECT 86.520 141.260 86.780 141.405 ;
        RECT 86.060 140.920 86.320 141.240 ;
        RECT 86.120 136.820 86.260 140.920 ;
        RECT 86.060 136.500 86.320 136.820 ;
        RECT 87.040 136.140 87.180 141.940 ;
        RECT 87.500 139.540 87.640 152.480 ;
        RECT 90.720 152.120 90.860 152.820 ;
        RECT 87.900 151.800 88.160 152.120 ;
        RECT 90.660 151.800 90.920 152.120 ;
        RECT 87.960 150.760 88.100 151.800 ;
        RECT 90.720 151.100 90.860 151.800 ;
        RECT 90.660 150.780 90.920 151.100 ;
        RECT 87.900 150.440 88.160 150.760 ;
        RECT 87.900 149.420 88.160 149.740 ;
        RECT 87.960 149.140 88.100 149.420 ;
        RECT 87.960 149.000 88.560 149.140 ;
        RECT 87.900 141.940 88.160 142.260 ;
        RECT 87.440 139.220 87.700 139.540 ;
        RECT 87.500 136.480 87.640 139.220 ;
        RECT 87.440 136.160 87.700 136.480 ;
        RECT 86.980 135.820 87.240 136.140 ;
        RECT 86.060 135.480 86.320 135.800 ;
        RECT 86.120 134.100 86.260 135.480 ;
        RECT 86.060 133.780 86.320 134.100 ;
        RECT 87.960 133.760 88.100 141.940 ;
        RECT 87.900 133.440 88.160 133.760 ;
        RECT 87.960 127.980 88.100 133.440 ;
        RECT 87.900 127.660 88.160 127.980 ;
        RECT 87.960 125.940 88.100 127.660 ;
        RECT 87.900 125.620 88.160 125.940 ;
        RECT 86.520 125.280 86.780 125.600 ;
        RECT 86.060 124.600 86.320 124.920 ;
        RECT 86.120 123.900 86.260 124.600 ;
        RECT 86.580 123.900 86.720 125.280 ;
        RECT 86.060 123.580 86.320 123.900 ;
        RECT 86.520 123.580 86.780 123.900 ;
        RECT 85.660 123.160 86.260 123.300 ;
        RECT 85.600 122.560 85.860 122.880 ;
        RECT 85.660 121.180 85.800 122.560 ;
        RECT 85.600 120.860 85.860 121.180 ;
        RECT 82.840 120.180 83.100 120.500 ;
        RECT 84.680 120.180 84.940 120.500 ;
        RECT 81.460 115.420 81.720 115.740 ;
        RECT 86.120 114.720 86.260 123.160 ;
        RECT 87.960 120.500 88.100 125.620 ;
        RECT 87.900 120.180 88.160 120.500 ;
        RECT 80.540 114.630 80.800 114.720 ;
        RECT 80.140 114.490 80.800 114.630 ;
        RECT 80.540 114.400 80.800 114.490 ;
        RECT 86.060 114.400 86.320 114.720 ;
        RECT 79.160 114.060 79.420 114.380 ;
        RECT 76.880 113.185 78.760 113.555 ;
        RECT 79.220 112.340 79.360 114.060 ;
        RECT 64.900 112.020 65.160 112.340 ;
        RECT 68.120 112.020 68.380 112.340 ;
        RECT 75.480 112.020 75.740 112.340 ;
        RECT 79.160 112.020 79.420 112.340 ;
        RECT 60.300 111.680 60.560 112.000 ;
        RECT 60.360 110.300 60.500 111.680 ;
        RECT 63.980 111.000 64.240 111.320 ;
        RECT 65.820 111.000 66.080 111.320 ;
        RECT 61.880 110.465 63.760 110.835 ;
        RECT 60.300 109.980 60.560 110.300 ;
        RECT 64.040 109.620 64.180 111.000 ;
        RECT 65.880 109.620 66.020 111.000 ;
        RECT 63.980 109.300 64.240 109.620 ;
        RECT 65.820 109.300 66.080 109.620 ;
        RECT 57.540 108.960 57.800 109.280 ;
        RECT 57.600 106.900 57.740 108.960 ;
        RECT 66.280 108.620 66.540 108.940 ;
        RECT 60.300 108.280 60.560 108.600 ;
        RECT 65.820 108.280 66.080 108.600 ;
        RECT 57.540 106.580 57.800 106.900 ;
        RECT 60.360 94.980 60.500 108.280 ;
        RECT 61.880 105.025 63.760 105.395 ;
        RECT 65.880 94.980 66.020 108.280 ;
        RECT 66.340 107.580 66.480 108.620 ;
        RECT 68.180 107.580 68.320 112.020 ;
        RECT 71.340 111.680 71.600 112.000 ;
        RECT 75.540 111.840 75.680 112.020 ;
        RECT 75.540 111.700 76.600 111.840 ;
        RECT 66.280 107.260 66.540 107.580 ;
        RECT 68.120 107.260 68.380 107.580 ;
        RECT 71.400 94.980 71.540 111.680 ;
        RECT 76.460 109.620 76.600 111.700 ;
        RECT 78.240 111.680 78.500 112.000 ;
        RECT 76.400 109.300 76.660 109.620 ;
        RECT 78.300 109.280 78.440 111.680 ;
        RECT 79.680 111.320 79.820 114.400 ;
        RECT 80.540 113.720 80.800 114.040 ;
        RECT 83.760 113.720 84.020 114.040 ;
        RECT 86.980 113.720 87.240 114.040 ;
        RECT 80.600 112.680 80.740 113.720 ;
        RECT 82.380 112.700 82.640 113.020 ;
        RECT 80.540 112.360 80.800 112.680 ;
        RECT 79.620 111.000 79.880 111.320 ;
        RECT 78.240 108.960 78.500 109.280 ;
        RECT 76.400 108.280 76.660 108.600 ;
        RECT 76.460 102.220 76.600 108.280 ;
        RECT 76.880 107.745 78.760 108.115 ;
        RECT 76.460 102.080 77.060 102.220 ;
        RECT 76.920 94.980 77.060 102.080 ;
        RECT 82.440 94.980 82.580 112.700 ;
        RECT 83.820 109.620 83.960 113.720 ;
        RECT 87.040 109.620 87.180 113.720 ;
        RECT 87.960 112.340 88.100 120.180 ;
        RECT 88.420 112.340 88.560 149.000 ;
        RECT 91.880 148.545 93.760 148.915 ;
        RECT 94.400 143.960 94.540 152.820 ;
        RECT 95.260 152.480 95.520 152.800 ;
        RECT 95.320 151.100 95.460 152.480 ;
        RECT 96.700 151.100 96.840 155.540 ;
        RECT 98.080 153.480 98.220 156.220 ;
        RECT 98.020 153.160 98.280 153.480 ;
        RECT 98.480 151.800 98.740 152.120 ;
        RECT 98.540 151.100 98.680 151.800 ;
        RECT 95.260 150.780 95.520 151.100 ;
        RECT 96.640 150.780 96.900 151.100 ;
        RECT 98.480 150.780 98.740 151.100 ;
        RECT 94.340 143.640 94.600 143.960 ;
        RECT 91.880 143.105 93.760 143.475 ;
        RECT 93.880 141.940 94.140 142.260 ;
        RECT 96.180 141.940 96.440 142.260 ;
        RECT 88.820 141.260 89.080 141.580 ;
        RECT 88.880 140.220 89.020 141.260 ;
        RECT 88.820 139.900 89.080 140.220 ;
        RECT 91.120 139.560 91.380 139.880 ;
        RECT 90.200 138.200 90.460 138.520 ;
        RECT 90.260 137.160 90.400 138.200 ;
        RECT 91.180 137.500 91.320 139.560 ;
        RECT 91.880 137.665 93.760 138.035 ;
        RECT 93.940 137.500 94.080 141.940 ;
        RECT 96.240 138.520 96.380 141.940 ;
        RECT 97.560 141.600 97.820 141.920 ;
        RECT 98.480 141.600 98.740 141.920 ;
        RECT 97.100 140.920 97.360 141.240 ;
        RECT 97.160 139.540 97.300 140.920 ;
        RECT 97.100 139.220 97.360 139.540 ;
        RECT 96.180 138.200 96.440 138.520 ;
        RECT 91.120 137.180 91.380 137.500 ;
        RECT 93.880 137.180 94.140 137.500 ;
        RECT 90.200 136.840 90.460 137.160 ;
        RECT 90.660 136.160 90.920 136.480 ;
        RECT 90.720 131.040 90.860 136.160 ;
        RECT 96.240 136.140 96.380 138.200 ;
        RECT 97.620 137.500 97.760 141.600 ;
        RECT 98.540 140.220 98.680 141.600 ;
        RECT 98.480 139.900 98.740 140.220 ;
        RECT 97.560 137.180 97.820 137.500 ;
        RECT 96.180 135.820 96.440 136.140 ;
        RECT 98.480 135.480 98.740 135.800 ;
        RECT 91.880 132.225 93.760 132.595 ;
        RECT 95.720 131.060 95.980 131.380 ;
        RECT 90.660 130.720 90.920 131.040 ;
        RECT 94.340 130.040 94.600 130.360 ;
        RECT 94.400 128.660 94.540 130.040 ;
        RECT 94.340 128.340 94.600 128.660 ;
        RECT 91.880 126.785 93.760 127.155 ;
        RECT 95.780 125.940 95.920 131.060 ;
        RECT 96.180 130.380 96.440 130.700 ;
        RECT 96.640 130.380 96.900 130.700 ;
        RECT 96.240 129.000 96.380 130.380 ;
        RECT 96.700 129.340 96.840 130.380 ;
        RECT 96.640 129.020 96.900 129.340 ;
        RECT 96.180 128.680 96.440 129.000 ;
        RECT 95.720 125.620 95.980 125.940 ;
        RECT 89.280 125.280 89.540 125.600 ;
        RECT 89.340 123.220 89.480 125.280 ;
        RECT 89.740 124.600 90.000 124.920 ;
        RECT 90.660 124.600 90.920 124.920 ;
        RECT 92.960 124.600 93.220 124.920 ;
        RECT 89.800 123.560 89.940 124.600 ;
        RECT 89.740 123.240 90.000 123.560 ;
        RECT 90.720 123.220 90.860 124.600 ;
        RECT 93.020 123.900 93.160 124.600 ;
        RECT 92.960 123.580 93.220 123.900 ;
        RECT 89.280 122.900 89.540 123.220 ;
        RECT 90.660 122.900 90.920 123.220 ;
        RECT 89.740 121.880 90.000 122.200 ;
        RECT 93.880 121.880 94.140 122.200 ;
        RECT 89.800 119.820 89.940 121.880 ;
        RECT 91.880 121.345 93.760 121.715 ;
        RECT 93.940 120.500 94.080 121.880 ;
        RECT 93.880 120.180 94.140 120.500 ;
        RECT 89.740 119.500 90.000 119.820 ;
        RECT 91.880 115.905 93.760 116.275 ;
        RECT 90.200 114.060 90.460 114.380 ;
        RECT 90.260 112.340 90.400 114.060 ;
        RECT 94.340 113.720 94.600 114.040 ;
        RECT 96.640 113.720 96.900 114.040 ;
        RECT 93.880 112.700 94.140 113.020 ;
        RECT 87.900 112.020 88.160 112.340 ;
        RECT 88.360 112.020 88.620 112.340 ;
        RECT 90.200 112.020 90.460 112.340 ;
        RECT 87.960 110.300 88.100 112.020 ;
        RECT 89.740 111.680 90.000 112.000 ;
        RECT 87.900 109.980 88.160 110.300 ;
        RECT 83.760 109.300 84.020 109.620 ;
        RECT 86.980 109.300 87.240 109.620 ;
        RECT 87.960 106.900 88.100 109.980 ;
        RECT 89.800 108.940 89.940 111.680 ;
        RECT 91.880 110.465 93.760 110.835 ;
        RECT 89.740 108.620 90.000 108.940 ;
        RECT 88.360 108.280 88.620 108.600 ;
        RECT 87.900 106.580 88.160 106.900 ;
        RECT 88.420 106.300 88.560 108.280 ;
        RECT 87.960 106.160 88.560 106.300 ;
        RECT 87.960 94.980 88.100 106.160 ;
        RECT 91.880 105.025 93.760 105.395 ;
        RECT 93.940 104.260 94.080 112.700 ;
        RECT 94.400 112.680 94.540 113.720 ;
        RECT 96.180 112.700 96.440 113.020 ;
        RECT 94.340 112.360 94.600 112.680 ;
        RECT 96.240 106.560 96.380 112.700 ;
        RECT 96.700 112.680 96.840 113.720 ;
        RECT 98.540 112.680 98.680 135.480 ;
        RECT 99.000 128.855 99.140 171.860 ;
        RECT 99.400 168.120 99.660 168.440 ;
        RECT 99.460 167.080 99.600 168.120 ;
        RECT 99.400 166.760 99.660 167.080 ;
        RECT 99.400 154.520 99.660 154.840 ;
        RECT 99.460 136.480 99.600 154.520 ;
        RECT 99.920 136.820 100.060 176.280 ;
        RECT 100.780 174.580 101.040 174.900 ;
        RECT 100.840 163.680 100.980 174.580 ;
        RECT 101.240 168.800 101.500 169.120 ;
        RECT 101.300 164.700 101.440 168.800 ;
        RECT 103.080 168.120 103.340 168.440 ;
        RECT 103.140 166.740 103.280 168.120 ;
        RECT 103.080 166.420 103.340 166.740 ;
        RECT 101.240 164.380 101.500 164.700 ;
        RECT 103.540 163.700 103.800 164.020 ;
        RECT 100.780 163.360 101.040 163.680 ;
        RECT 100.840 160.960 100.980 163.360 ;
        RECT 101.700 162.680 101.960 163.000 ;
        RECT 100.780 160.640 101.040 160.960 ;
        RECT 101.760 155.860 101.900 162.680 ;
        RECT 103.600 161.980 103.740 163.700 ;
        RECT 103.540 161.660 103.800 161.980 ;
        RECT 100.780 155.540 101.040 155.860 ;
        RECT 101.240 155.540 101.500 155.860 ;
        RECT 101.700 155.540 101.960 155.860 ;
        RECT 100.840 153.820 100.980 155.540 ;
        RECT 100.780 153.500 101.040 153.820 ;
        RECT 101.300 152.655 101.440 155.540 ;
        RECT 103.070 152.965 103.350 153.335 ;
        RECT 103.140 152.800 103.280 152.965 ;
        RECT 101.230 152.285 101.510 152.655 ;
        RECT 103.080 152.480 103.340 152.800 ;
        RECT 101.300 148.040 101.440 152.285 ;
        RECT 102.620 151.800 102.880 152.120 ;
        RECT 102.680 150.760 102.820 151.800 ;
        RECT 102.620 150.440 102.880 150.760 ;
        RECT 101.240 147.720 101.500 148.040 ;
        RECT 104.060 147.700 104.200 176.280 ;
        RECT 106.820 175.580 106.960 176.960 ;
        RECT 108.140 176.620 108.400 176.940 ;
        RECT 106.760 175.260 107.020 175.580 ;
        RECT 108.200 174.560 108.340 176.620 ;
        RECT 108.660 175.240 108.800 177.445 ;
        RECT 109.060 177.300 109.320 177.620 ;
        RECT 109.980 177.300 110.240 177.620 ;
        RECT 110.430 177.445 110.710 177.815 ;
        RECT 108.600 174.920 108.860 175.240 ;
        RECT 108.140 174.240 108.400 174.560 ;
        RECT 106.880 173.025 108.760 173.395 ;
        RECT 109.120 172.520 109.260 177.300 ;
        RECT 110.040 174.810 110.180 177.300 ;
        RECT 110.960 176.940 111.100 179.680 ;
        RECT 111.420 177.620 111.560 194.300 ;
        RECT 111.880 186.120 112.020 194.300 ;
        RECT 118.320 191.220 118.460 196.000 ;
        RECT 121.080 194.620 121.220 199.400 ;
        RECT 121.880 197.505 123.760 197.875 ;
        RECT 121.020 194.300 121.280 194.620 ;
        RECT 121.880 192.065 123.760 192.435 ;
        RECT 118.260 190.900 118.520 191.220 ;
        RECT 112.280 190.220 112.540 190.540 ;
        RECT 115.960 190.220 116.220 190.540 ;
        RECT 112.340 189.180 112.480 190.220 ;
        RECT 112.280 188.860 112.540 189.180 ;
        RECT 115.500 187.160 115.760 187.480 ;
        RECT 111.820 186.030 112.080 186.120 ;
        RECT 111.820 185.890 112.480 186.030 ;
        RECT 111.820 185.800 112.080 185.890 ;
        RECT 112.340 183.060 112.480 185.890 ;
        RECT 115.560 185.100 115.700 187.160 ;
        RECT 115.500 184.780 115.760 185.100 ;
        RECT 113.200 184.440 113.460 184.760 ;
        RECT 115.040 184.440 115.300 184.760 ;
        RECT 112.740 183.080 113.000 183.400 ;
        RECT 111.820 182.740 112.080 183.060 ;
        RECT 112.280 182.740 112.540 183.060 ;
        RECT 111.880 180.000 112.020 182.740 ;
        RECT 112.280 181.720 112.540 182.040 ;
        RECT 111.820 179.680 112.080 180.000 ;
        RECT 111.880 178.300 112.020 179.680 ;
        RECT 111.820 177.980 112.080 178.300 ;
        RECT 111.360 177.300 111.620 177.620 ;
        RECT 110.900 176.620 111.160 176.940 ;
        RECT 111.880 175.580 112.020 177.980 ;
        RECT 111.820 175.260 112.080 175.580 ;
        RECT 110.440 174.810 110.700 174.900 ;
        RECT 111.360 174.810 111.620 174.900 ;
        RECT 110.040 174.670 110.700 174.810 ;
        RECT 110.440 174.580 110.700 174.670 ;
        RECT 110.960 174.670 111.620 174.810 ;
        RECT 110.960 174.220 111.100 174.670 ;
        RECT 111.360 174.580 111.620 174.670 ;
        RECT 110.900 173.900 111.160 174.220 ;
        RECT 111.360 173.900 111.620 174.220 ;
        RECT 109.060 172.200 109.320 172.520 ;
        RECT 109.120 169.120 109.260 172.200 ;
        RECT 109.060 168.800 109.320 169.120 ;
        RECT 106.300 168.460 106.560 168.780 ;
        RECT 105.840 168.120 106.100 168.440 ;
        RECT 105.900 163.340 106.040 168.120 ;
        RECT 106.360 166.400 106.500 168.460 ;
        RECT 106.880 167.585 108.760 167.955 ;
        RECT 109.120 166.400 109.260 168.800 ;
        RECT 110.440 168.120 110.700 168.440 ;
        RECT 110.500 167.080 110.640 168.120 ;
        RECT 110.440 166.760 110.700 167.080 ;
        RECT 106.300 166.080 106.560 166.400 ;
        RECT 109.060 166.080 109.320 166.400 ;
        RECT 105.840 163.020 106.100 163.340 ;
        RECT 104.920 162.680 105.180 163.000 ;
        RECT 106.360 162.740 106.500 166.080 ;
        RECT 109.120 163.680 109.260 166.080 ;
        RECT 109.060 163.360 109.320 163.680 ;
        RECT 104.980 161.640 105.120 162.680 ;
        RECT 105.900 162.600 106.500 162.740 ;
        RECT 105.900 161.980 106.040 162.600 ;
        RECT 105.840 161.660 106.100 161.980 ;
        RECT 104.920 161.320 105.180 161.640 ;
        RECT 105.380 157.920 105.640 158.240 ;
        RECT 105.440 155.520 105.580 157.920 ;
        RECT 106.360 156.200 106.500 162.600 ;
        RECT 106.880 162.145 108.760 162.515 ;
        RECT 109.520 157.920 109.780 158.240 ;
        RECT 106.880 156.705 108.760 157.075 ;
        RECT 109.580 156.540 109.720 157.920 ;
        RECT 109.980 157.240 110.240 157.560 ;
        RECT 110.440 157.240 110.700 157.560 ;
        RECT 110.040 156.540 110.180 157.240 ;
        RECT 107.220 156.220 107.480 156.540 ;
        RECT 109.520 156.220 109.780 156.540 ;
        RECT 109.980 156.220 110.240 156.540 ;
        RECT 106.300 155.880 106.560 156.200 ;
        RECT 107.280 155.860 107.420 156.220 ;
        RECT 107.220 155.540 107.480 155.860 ;
        RECT 107.670 155.685 107.950 156.055 ;
        RECT 109.520 155.770 109.780 155.860 ;
        RECT 110.040 155.770 110.180 156.220 ;
        RECT 105.380 155.200 105.640 155.520 ;
        RECT 105.440 152.800 105.580 155.200 ;
        RECT 106.300 154.520 106.560 154.840 ;
        RECT 106.760 154.520 107.020 154.840 ;
        RECT 105.380 152.480 105.640 152.800 ;
        RECT 105.840 152.140 106.100 152.460 ;
        RECT 104.460 151.800 104.720 152.120 ;
        RECT 104.520 150.760 104.660 151.800 ;
        RECT 104.460 150.440 104.720 150.760 ;
        RECT 104.000 147.380 104.260 147.700 ;
        RECT 105.900 147.360 106.040 152.140 ;
        RECT 105.840 147.040 106.100 147.360 ;
        RECT 102.160 143.640 102.420 143.960 ;
        RECT 102.220 141.920 102.360 143.640 ;
        RECT 105.840 141.940 106.100 142.260 ;
        RECT 100.320 141.775 100.580 141.920 ;
        RECT 100.310 141.405 100.590 141.775 ;
        RECT 102.160 141.600 102.420 141.920 ;
        RECT 104.460 141.600 104.720 141.920 ;
        RECT 100.780 140.920 101.040 141.240 ;
        RECT 102.620 140.920 102.880 141.240 ;
        RECT 99.860 136.500 100.120 136.820 ;
        RECT 100.840 136.480 100.980 140.920 ;
        RECT 102.680 139.880 102.820 140.920 ;
        RECT 104.520 140.220 104.660 141.600 ;
        RECT 104.920 141.260 105.180 141.580 ;
        RECT 104.460 139.900 104.720 140.220 ;
        RECT 102.620 139.560 102.880 139.880 ;
        RECT 104.980 138.520 105.120 141.260 ;
        RECT 105.900 139.620 106.040 141.940 ;
        RECT 106.360 139.790 106.500 154.520 ;
        RECT 106.820 152.800 106.960 154.520 ;
        RECT 107.280 153.820 107.420 155.540 ;
        RECT 107.220 153.500 107.480 153.820 ;
        RECT 107.280 152.800 107.420 153.500 ;
        RECT 107.740 153.140 107.880 155.685 ;
        RECT 109.520 155.630 110.180 155.770 ;
        RECT 109.520 155.540 109.780 155.630 ;
        RECT 108.600 155.090 108.860 155.180 ;
        RECT 108.200 154.950 108.860 155.090 ;
        RECT 107.680 152.820 107.940 153.140 ;
        RECT 106.760 152.655 107.020 152.800 ;
        RECT 106.750 152.285 107.030 152.655 ;
        RECT 107.220 152.480 107.480 152.800 ;
        RECT 108.200 152.460 108.340 154.950 ;
        RECT 108.600 154.860 108.860 154.950 ;
        RECT 109.980 153.160 110.240 153.480 ;
        RECT 110.500 153.220 110.640 157.240 ;
        RECT 110.960 156.200 111.100 173.900 ;
        RECT 110.900 155.880 111.160 156.200 ;
        RECT 108.600 152.655 108.860 152.800 ;
        RECT 110.040 152.710 110.180 153.160 ;
        RECT 110.500 153.080 111.100 153.220 ;
        RECT 108.140 152.140 108.400 152.460 ;
        RECT 108.590 152.285 108.870 152.655 ;
        RECT 110.040 152.570 110.640 152.710 ;
        RECT 108.600 152.030 108.860 152.120 ;
        RECT 108.600 151.890 109.720 152.030 ;
        RECT 108.600 151.800 108.860 151.890 ;
        RECT 106.880 151.265 108.760 151.635 ;
        RECT 108.140 150.100 108.400 150.420 ;
        RECT 108.200 146.930 108.340 150.100 ;
        RECT 109.060 149.080 109.320 149.400 ;
        RECT 109.120 147.700 109.260 149.080 ;
        RECT 109.060 147.380 109.320 147.700 ;
        RECT 109.580 147.360 109.720 151.890 ;
        RECT 109.980 151.800 110.240 152.120 ;
        RECT 110.040 150.760 110.180 151.800 ;
        RECT 109.980 150.440 110.240 150.760 ;
        RECT 110.040 149.255 110.180 150.440 ;
        RECT 110.500 150.420 110.640 152.570 ;
        RECT 110.440 150.100 110.700 150.420 ;
        RECT 110.440 149.420 110.700 149.740 ;
        RECT 109.970 148.885 110.250 149.255 ;
        RECT 109.980 147.720 110.240 148.040 ;
        RECT 109.520 147.040 109.780 147.360 ;
        RECT 109.060 146.930 109.320 147.020 ;
        RECT 108.200 146.790 109.320 146.930 ;
        RECT 109.060 146.700 109.320 146.790 ;
        RECT 106.880 145.825 108.760 146.195 ;
        RECT 108.140 144.320 108.400 144.640 ;
        RECT 108.200 141.920 108.340 144.320 ;
        RECT 109.120 144.300 109.260 146.700 ;
        RECT 110.040 146.420 110.180 147.720 ;
        RECT 109.580 146.280 110.180 146.420 ;
        RECT 109.060 143.980 109.320 144.300 ;
        RECT 108.140 141.600 108.400 141.920 ;
        RECT 108.600 141.490 108.860 141.580 ;
        RECT 108.600 141.350 109.260 141.490 ;
        RECT 108.600 141.260 108.860 141.350 ;
        RECT 106.880 140.385 108.760 140.755 ;
        RECT 109.120 140.220 109.260 141.350 ;
        RECT 108.140 139.900 108.400 140.220 ;
        RECT 109.060 139.900 109.320 140.220 ;
        RECT 106.360 139.650 106.960 139.790 ;
        RECT 105.440 139.480 106.040 139.620 ;
        RECT 105.440 138.520 105.580 139.480 ;
        RECT 105.840 138.880 106.100 139.200 ;
        RECT 104.920 138.200 105.180 138.520 ;
        RECT 105.380 138.200 105.640 138.520 ;
        RECT 102.160 137.180 102.420 137.500 ;
        RECT 99.400 136.160 99.660 136.480 ;
        RECT 100.780 136.160 101.040 136.480 ;
        RECT 98.930 128.485 99.210 128.855 ;
        RECT 98.940 128.340 99.200 128.485 ;
        RECT 102.220 125.600 102.360 137.180 ;
        RECT 105.440 137.160 105.580 138.200 ;
        RECT 105.380 136.840 105.640 137.160 ;
        RECT 105.380 135.480 105.640 135.800 ;
        RECT 103.080 131.060 103.340 131.380 ;
        RECT 103.140 125.600 103.280 131.060 ;
        RECT 102.160 125.280 102.420 125.600 ;
        RECT 103.080 125.280 103.340 125.600 ;
        RECT 101.240 124.600 101.500 124.920 ;
        RECT 104.920 124.600 105.180 124.920 ;
        RECT 99.400 122.560 99.660 122.880 ;
        RECT 99.460 121.180 99.600 122.560 ;
        RECT 99.400 120.860 99.660 121.180 ;
        RECT 101.300 120.160 101.440 124.600 ;
        RECT 104.980 123.560 105.120 124.600 ;
        RECT 104.920 123.240 105.180 123.560 ;
        RECT 101.240 119.840 101.500 120.160 ;
        RECT 105.440 115.400 105.580 135.480 ;
        RECT 105.900 131.040 106.040 138.880 ;
        RECT 106.300 137.180 106.560 137.500 ;
        RECT 106.360 132.060 106.500 137.180 ;
        RECT 106.820 136.140 106.960 139.650 ;
        RECT 106.760 135.820 107.020 136.140 ;
        RECT 108.200 135.800 108.340 139.900 ;
        RECT 108.590 138.685 108.870 139.055 ;
        RECT 108.660 136.820 108.800 138.685 ;
        RECT 109.120 137.500 109.260 139.900 ;
        RECT 109.060 137.180 109.320 137.500 ;
        RECT 108.600 136.500 108.860 136.820 ;
        RECT 108.140 135.480 108.400 135.800 ;
        RECT 106.880 134.945 108.760 135.315 ;
        RECT 109.580 134.780 109.720 146.280 ;
        RECT 110.500 145.320 110.640 149.420 ;
        RECT 110.960 149.400 111.100 153.080 ;
        RECT 110.900 149.080 111.160 149.400 ;
        RECT 110.900 148.060 111.160 148.380 ;
        RECT 110.440 145.000 110.700 145.320 ;
        RECT 110.440 143.980 110.700 144.300 ;
        RECT 110.500 142.600 110.640 143.980 ;
        RECT 110.440 142.280 110.700 142.600 ;
        RECT 110.500 141.775 110.640 142.280 ;
        RECT 110.430 141.405 110.710 141.775 ;
        RECT 109.980 140.920 110.240 141.240 ;
        RECT 110.040 139.540 110.180 140.920 ;
        RECT 109.980 139.220 110.240 139.540 ;
        RECT 109.980 137.180 110.240 137.500 ;
        RECT 110.040 136.480 110.180 137.180 ;
        RECT 109.980 136.160 110.240 136.480 ;
        RECT 110.500 136.140 110.640 141.405 ;
        RECT 110.440 135.820 110.700 136.140 ;
        RECT 109.520 134.460 109.780 134.780 ;
        RECT 110.960 134.440 111.100 148.060 ;
        RECT 111.420 144.980 111.560 173.900 ;
        RECT 111.820 157.240 112.080 157.560 ;
        RECT 111.880 144.980 112.020 157.240 ;
        RECT 112.340 147.700 112.480 181.720 ;
        RECT 112.800 180.000 112.940 183.080 ;
        RECT 113.260 180.340 113.400 184.440 ;
        RECT 115.100 183.060 115.240 184.440 ;
        RECT 116.020 183.740 116.160 190.220 ;
        RECT 118.320 188.160 118.460 190.900 ;
        RECT 119.180 190.560 119.440 190.880 ;
        RECT 118.260 187.840 118.520 188.160 ;
        RECT 119.240 186.460 119.380 190.560 ;
        RECT 123.320 189.880 123.580 190.200 ;
        RECT 123.380 188.840 123.520 189.880 ;
        RECT 123.320 188.520 123.580 188.840 ;
        RECT 124.700 187.840 124.960 188.160 ;
        RECT 121.880 186.625 123.760 186.995 ;
        RECT 119.180 186.140 119.440 186.460 ;
        RECT 115.960 183.420 116.220 183.740 ;
        RECT 115.040 182.740 115.300 183.060 ;
        RECT 121.880 181.185 123.760 181.555 ;
        RECT 113.200 180.020 113.460 180.340 ;
        RECT 124.240 180.020 124.500 180.340 ;
        RECT 112.740 179.680 113.000 180.000 ;
        RECT 116.880 179.680 117.140 180.000 ;
        RECT 114.580 179.000 114.840 179.320 ;
        RECT 112.740 174.580 113.000 174.900 ;
        RECT 112.800 171.840 112.940 174.580 ;
        RECT 113.200 173.560 113.460 173.880 ;
        RECT 113.260 172.520 113.400 173.560 ;
        RECT 113.200 172.200 113.460 172.520 ;
        RECT 112.740 171.520 113.000 171.840 ;
        RECT 112.800 169.460 112.940 171.520 ;
        RECT 112.740 169.140 113.000 169.460 ;
        RECT 112.800 164.020 112.940 169.140 ;
        RECT 112.740 163.700 113.000 164.020 ;
        RECT 112.800 160.960 112.940 163.700 ;
        RECT 112.740 160.640 113.000 160.960 ;
        RECT 113.260 158.240 113.400 172.200 ;
        RECT 114.120 165.400 114.380 165.720 ;
        RECT 114.180 164.700 114.320 165.400 ;
        RECT 114.120 164.380 114.380 164.700 ;
        RECT 112.740 157.920 113.000 158.240 ;
        RECT 113.200 157.920 113.460 158.240 ;
        RECT 114.120 157.920 114.380 158.240 ;
        RECT 112.800 155.520 112.940 157.920 ;
        RECT 114.180 156.540 114.320 157.920 ;
        RECT 114.120 156.220 114.380 156.540 ;
        RECT 112.740 155.200 113.000 155.520 ;
        RECT 114.120 152.820 114.380 153.140 ;
        RECT 112.730 152.285 113.010 152.655 ;
        RECT 112.800 150.420 112.940 152.285 ;
        RECT 113.200 151.800 113.460 152.120 ;
        RECT 113.660 151.800 113.920 152.120 ;
        RECT 112.740 150.100 113.000 150.420 ;
        RECT 113.260 149.740 113.400 151.800 ;
        RECT 113.720 151.100 113.860 151.800 ;
        RECT 113.660 150.780 113.920 151.100 ;
        RECT 114.180 150.500 114.320 152.820 ;
        RECT 113.720 150.360 114.320 150.500 ;
        RECT 113.200 149.420 113.460 149.740 ;
        RECT 112.740 149.080 113.000 149.400 ;
        RECT 112.280 147.380 112.540 147.700 ;
        RECT 112.800 147.100 112.940 149.080 ;
        RECT 113.190 148.885 113.470 149.255 ;
        RECT 113.260 147.360 113.400 148.885 ;
        RECT 112.340 146.960 112.940 147.100 ;
        RECT 113.200 147.040 113.460 147.360 ;
        RECT 111.360 144.660 111.620 144.980 ;
        RECT 111.820 144.660 112.080 144.980 ;
        RECT 111.820 143.640 112.080 143.960 ;
        RECT 111.360 142.620 111.620 142.940 ;
        RECT 111.420 136.820 111.560 142.620 ;
        RECT 111.360 136.500 111.620 136.820 ;
        RECT 111.360 135.480 111.620 135.800 ;
        RECT 110.900 134.120 111.160 134.440 ;
        RECT 107.220 133.780 107.480 134.100 ;
        RECT 106.300 131.740 106.560 132.060 ;
        RECT 107.280 131.040 107.420 133.780 ;
        RECT 110.440 133.440 110.700 133.760 ;
        RECT 110.900 133.440 111.160 133.760 ;
        RECT 105.840 130.720 106.100 131.040 ;
        RECT 107.220 130.720 107.480 131.040 ;
        RECT 109.520 130.720 109.780 131.040 ;
        RECT 105.900 129.340 106.040 130.720 ;
        RECT 106.880 129.505 108.760 129.875 ;
        RECT 105.840 129.020 106.100 129.340 ;
        RECT 105.900 123.900 106.040 129.020 ;
        RECT 109.060 128.000 109.320 128.320 ;
        RECT 106.300 125.280 106.560 125.600 ;
        RECT 105.840 123.580 106.100 123.900 ;
        RECT 106.360 122.880 106.500 125.280 ;
        RECT 109.120 124.920 109.260 128.000 ;
        RECT 109.580 125.600 109.720 130.720 ;
        RECT 110.500 125.600 110.640 133.440 ;
        RECT 110.960 130.700 111.100 133.440 ;
        RECT 110.900 130.380 111.160 130.700 ;
        RECT 109.520 125.280 109.780 125.600 ;
        RECT 110.440 125.280 110.700 125.600 ;
        RECT 109.060 124.600 109.320 124.920 ;
        RECT 106.880 124.065 108.760 124.435 ;
        RECT 106.300 122.560 106.560 122.880 ;
        RECT 109.120 122.200 109.260 124.600 ;
        RECT 110.900 122.900 111.160 123.220 ;
        RECT 109.060 121.880 109.320 122.200 ;
        RECT 109.120 121.180 109.260 121.880 ;
        RECT 109.060 120.860 109.320 121.180 ;
        RECT 110.960 120.500 111.100 122.900 ;
        RECT 110.900 120.180 111.160 120.500 ;
        RECT 106.880 118.625 108.760 118.995 ;
        RECT 105.380 115.080 105.640 115.400 ;
        RECT 109.520 115.080 109.780 115.400 ;
        RECT 98.940 113.720 99.200 114.040 ;
        RECT 105.380 113.720 105.640 114.040 ;
        RECT 109.060 113.720 109.320 114.040 ;
        RECT 96.640 112.360 96.900 112.680 ;
        RECT 98.480 112.360 98.740 112.680 ;
        RECT 99.000 107.240 99.140 113.720 ;
        RECT 104.460 112.700 104.720 113.020 ;
        RECT 98.940 106.920 99.200 107.240 ;
        RECT 96.180 106.240 96.440 106.560 ;
        RECT 98.940 105.560 99.200 105.880 ;
        RECT 93.480 104.120 94.080 104.260 ;
        RECT 93.480 94.980 93.620 104.120 ;
        RECT 99.000 94.980 99.140 105.560 ;
        RECT 104.520 94.980 104.660 112.700 ;
        RECT 105.440 112.680 105.580 113.720 ;
        RECT 106.880 113.185 108.760 113.555 ;
        RECT 105.380 112.360 105.640 112.680 ;
        RECT 109.120 108.940 109.260 113.720 ;
        RECT 109.580 112.680 109.720 115.080 ;
        RECT 110.960 115.060 111.100 120.180 ;
        RECT 110.900 114.970 111.160 115.060 ;
        RECT 110.500 114.830 111.160 114.970 ;
        RECT 109.520 112.360 109.780 112.680 ;
        RECT 110.500 112.340 110.640 114.830 ;
        RECT 110.900 114.740 111.160 114.830 ;
        RECT 111.420 112.340 111.560 135.480 ;
        RECT 111.880 134.780 112.020 143.640 ;
        RECT 112.340 136.480 112.480 146.960 ;
        RECT 113.260 145.570 113.400 147.040 ;
        RECT 112.800 145.430 113.400 145.570 ;
        RECT 112.800 142.940 112.940 145.430 ;
        RECT 113.720 145.060 113.860 150.360 ;
        RECT 114.120 149.080 114.380 149.400 ;
        RECT 114.180 147.360 114.320 149.080 ;
        RECT 114.120 147.040 114.380 147.360 ;
        RECT 113.260 144.920 113.860 145.060 ;
        RECT 112.740 142.620 113.000 142.940 ;
        RECT 113.260 142.260 113.400 144.920 ;
        RECT 114.180 142.260 114.320 147.040 ;
        RECT 113.200 141.940 113.460 142.260 ;
        RECT 114.120 141.940 114.380 142.260 ;
        RECT 112.740 141.260 113.000 141.580 ;
        RECT 112.800 140.220 112.940 141.260 ;
        RECT 112.740 139.900 113.000 140.220 ;
        RECT 113.260 138.860 113.400 141.940 ;
        RECT 113.660 140.920 113.920 141.240 ;
        RECT 113.200 138.540 113.460 138.860 ;
        RECT 113.200 137.180 113.460 137.500 ;
        RECT 112.280 136.160 112.540 136.480 ;
        RECT 111.820 134.460 112.080 134.780 ;
        RECT 112.280 133.780 112.540 134.100 ;
        RECT 112.340 128.660 112.480 133.780 ;
        RECT 112.740 133.100 113.000 133.420 ;
        RECT 112.800 130.360 112.940 133.100 ;
        RECT 112.740 130.040 113.000 130.360 ;
        RECT 112.800 129.000 112.940 130.040 ;
        RECT 113.260 129.340 113.400 137.180 ;
        RECT 113.720 136.480 113.860 140.920 ;
        RECT 114.120 138.200 114.380 138.520 ;
        RECT 114.180 136.480 114.320 138.200 ;
        RECT 114.640 136.820 114.780 179.000 ;
        RECT 116.940 177.620 117.080 179.680 ;
        RECT 117.340 179.000 117.600 179.320 ;
        RECT 116.880 177.300 117.140 177.620 ;
        RECT 115.500 176.960 115.760 177.280 ;
        RECT 115.560 175.580 115.700 176.960 ;
        RECT 115.500 175.260 115.760 175.580 ;
        RECT 116.420 170.840 116.680 171.160 ;
        RECT 115.960 169.480 116.220 169.800 ;
        RECT 116.020 168.780 116.160 169.480 ;
        RECT 115.500 168.460 115.760 168.780 ;
        RECT 115.960 168.460 116.220 168.780 ;
        RECT 115.040 168.120 115.300 168.440 ;
        RECT 115.100 163.680 115.240 168.120 ;
        RECT 115.560 165.720 115.700 168.460 ;
        RECT 115.500 165.400 115.760 165.720 ;
        RECT 115.040 163.360 115.300 163.680 ;
        RECT 116.020 155.860 116.160 168.460 ;
        RECT 116.480 163.340 116.620 170.840 ;
        RECT 116.940 169.120 117.080 177.300 ;
        RECT 117.400 172.520 117.540 179.000 ;
        RECT 124.300 178.300 124.440 180.020 ;
        RECT 124.760 179.660 124.900 187.840 ;
        RECT 124.700 179.340 124.960 179.660 ;
        RECT 124.240 177.980 124.500 178.300 ;
        RECT 118.260 176.280 118.520 176.600 ;
        RECT 117.800 174.920 118.060 175.240 ;
        RECT 117.340 172.200 117.600 172.520 ;
        RECT 117.860 171.840 118.000 174.920 ;
        RECT 118.320 174.220 118.460 176.280 ;
        RECT 121.880 175.745 123.760 176.115 ;
        RECT 124.760 174.900 124.900 179.340 ;
        RECT 124.700 174.580 124.960 174.900 ;
        RECT 118.260 173.900 118.520 174.220 ;
        RECT 121.940 173.900 122.200 174.220 ;
        RECT 122.850 174.045 123.130 174.415 ;
        RECT 122.000 172.860 122.140 173.900 ;
        RECT 121.940 172.540 122.200 172.860 ;
        RECT 122.920 172.520 123.060 174.045 ;
        RECT 135.630 173.380 136.780 174.600 ;
        RECT 122.860 172.200 123.120 172.520 ;
        RECT 117.800 171.520 118.060 171.840 ;
        RECT 118.720 171.180 118.980 171.500 ;
        RECT 118.780 169.120 118.920 171.180 ;
        RECT 121.880 170.305 123.760 170.675 ;
        RECT 129.290 170.560 133.760 172.150 ;
        RECT 116.880 168.800 117.140 169.120 ;
        RECT 118.720 168.800 118.980 169.120 ;
        RECT 117.340 168.120 117.600 168.440 ;
        RECT 117.400 166.740 117.540 168.120 ;
        RECT 117.340 166.420 117.600 166.740 ;
        RECT 116.880 165.400 117.140 165.720 ;
        RECT 116.420 163.020 116.680 163.340 ;
        RECT 116.480 156.055 116.620 163.020 ;
        RECT 116.940 163.000 117.080 165.400 ;
        RECT 116.880 162.680 117.140 163.000 ;
        RECT 116.940 158.580 117.080 162.680 ;
        RECT 118.780 161.300 118.920 168.800 ;
        RECT 121.480 166.760 121.740 167.080 ;
        RECT 121.540 164.700 121.680 166.760 ;
        RECT 135.630 166.640 136.740 173.380 ;
        RECT 126.080 166.080 126.340 166.400 ;
        RECT 121.880 164.865 123.760 165.235 ;
        RECT 121.480 164.380 121.740 164.700 ;
        RECT 118.720 160.980 118.980 161.300 ;
        RECT 117.340 160.640 117.600 160.960 ;
        RECT 117.400 159.260 117.540 160.640 ;
        RECT 121.880 159.425 123.760 159.795 ;
        RECT 117.340 158.940 117.600 159.260 ;
        RECT 116.880 158.260 117.140 158.580 ;
        RECT 115.960 155.540 116.220 155.860 ;
        RECT 116.410 155.685 116.690 156.055 ;
        RECT 116.020 153.335 116.160 155.540 ;
        RECT 117.400 155.260 117.540 158.940 ;
        RECT 124.240 155.880 124.500 156.200 ;
        RECT 116.940 155.120 117.540 155.260 ;
        RECT 115.950 152.965 116.230 153.335 ;
        RECT 115.500 150.100 115.760 150.420 ;
        RECT 115.040 147.720 115.300 148.040 ;
        RECT 114.580 136.500 114.840 136.820 ;
        RECT 113.660 136.160 113.920 136.480 ;
        RECT 114.120 136.160 114.380 136.480 ;
        RECT 115.100 136.220 115.240 147.720 ;
        RECT 115.560 147.360 115.700 150.100 ;
        RECT 116.020 147.360 116.160 152.965 ;
        RECT 115.500 147.040 115.760 147.360 ;
        RECT 115.960 147.040 116.220 147.360 ;
        RECT 115.560 144.640 115.700 147.040 ;
        RECT 115.500 144.320 115.760 144.640 ;
        RECT 115.960 143.640 116.220 143.960 ;
        RECT 114.640 136.080 115.240 136.220 ;
        RECT 113.660 131.060 113.920 131.380 ;
        RECT 113.200 129.020 113.460 129.340 ;
        RECT 112.740 128.680 113.000 129.000 ;
        RECT 112.280 128.340 112.540 128.660 ;
        RECT 112.800 126.280 112.940 128.680 ;
        RECT 113.720 126.620 113.860 131.060 ;
        RECT 113.660 126.300 113.920 126.620 ;
        RECT 112.740 125.960 113.000 126.280 ;
        RECT 113.660 124.940 113.920 125.260 ;
        RECT 112.280 124.600 112.540 124.920 ;
        RECT 112.340 123.220 112.480 124.600 ;
        RECT 113.720 123.220 113.860 124.940 ;
        RECT 112.280 122.900 112.540 123.220 ;
        RECT 113.660 122.900 113.920 123.220 ;
        RECT 113.660 121.880 113.920 122.200 ;
        RECT 113.720 119.820 113.860 121.880 ;
        RECT 113.660 119.500 113.920 119.820 ;
        RECT 114.640 112.340 114.780 136.080 ;
        RECT 115.040 121.880 115.300 122.200 ;
        RECT 115.100 117.780 115.240 121.880 ;
        RECT 115.500 120.180 115.760 120.500 ;
        RECT 115.560 118.460 115.700 120.180 ;
        RECT 115.500 118.140 115.760 118.460 ;
        RECT 115.040 117.460 115.300 117.780 ;
        RECT 116.020 117.440 116.160 143.640 ;
        RECT 116.420 140.920 116.680 141.240 ;
        RECT 116.480 136.820 116.620 140.920 ;
        RECT 116.420 136.500 116.680 136.820 ;
        RECT 116.940 131.040 117.080 155.120 ;
        RECT 117.340 154.520 117.600 154.840 ;
        RECT 117.400 153.820 117.540 154.520 ;
        RECT 121.880 153.985 123.760 154.355 ;
        RECT 124.300 153.820 124.440 155.880 ;
        RECT 126.140 155.520 126.280 166.080 ;
        RECT 135.630 165.420 136.780 166.640 ;
        RECT 126.080 155.200 126.340 155.520 ;
        RECT 117.340 153.500 117.600 153.820 ;
        RECT 124.240 153.500 124.500 153.820 ;
        RECT 117.400 152.800 117.540 153.500 ;
        RECT 117.340 152.480 117.600 152.800 ;
        RECT 118.260 152.140 118.520 152.460 ;
        RECT 118.320 149.400 118.460 152.140 ;
        RECT 124.240 151.800 124.500 152.120 ;
        RECT 120.560 150.440 120.820 150.760 ;
        RECT 118.260 149.080 118.520 149.400 ;
        RECT 120.620 148.380 120.760 150.440 ;
        RECT 124.300 150.420 124.440 151.800 ;
        RECT 126.140 150.420 126.280 155.200 ;
        RECT 124.240 150.100 124.500 150.420 ;
        RECT 126.080 150.100 126.340 150.420 ;
        RECT 121.880 148.545 123.760 148.915 ;
        RECT 120.560 148.060 120.820 148.380 ;
        RECT 120.100 147.040 120.360 147.360 ;
        RECT 119.640 146.700 119.900 147.020 ;
        RECT 118.260 143.640 118.520 143.960 ;
        RECT 118.320 139.880 118.460 143.640 ;
        RECT 118.260 139.560 118.520 139.880 ;
        RECT 119.700 139.440 119.840 146.700 ;
        RECT 120.160 144.980 120.300 147.040 ;
        RECT 120.100 144.660 120.360 144.980 ;
        RECT 120.100 143.640 120.360 143.960 ;
        RECT 120.160 141.580 120.300 143.640 ;
        RECT 121.880 143.105 123.760 143.475 ;
        RECT 123.320 141.940 123.580 142.260 ;
        RECT 120.100 141.260 120.360 141.580 ;
        RECT 121.940 139.440 122.200 139.540 ;
        RECT 119.700 139.300 120.300 139.440 ;
        RECT 116.880 130.720 117.140 131.040 ;
        RECT 116.420 125.280 116.680 125.600 ;
        RECT 116.480 123.900 116.620 125.280 ;
        RECT 116.420 123.580 116.680 123.900 ;
        RECT 116.940 123.300 117.080 130.720 ;
        RECT 118.720 130.040 118.980 130.360 ;
        RECT 118.780 129.000 118.920 130.040 ;
        RECT 118.720 128.680 118.980 129.000 ;
        RECT 117.800 126.300 118.060 126.620 ;
        RECT 116.480 123.220 117.080 123.300 ;
        RECT 116.420 123.160 117.080 123.220 ;
        RECT 116.420 122.900 116.680 123.160 ;
        RECT 117.860 122.880 118.000 126.300 ;
        RECT 119.640 124.940 119.900 125.260 ;
        RECT 119.700 123.900 119.840 124.940 ;
        RECT 119.640 123.580 119.900 123.900 ;
        RECT 117.800 122.560 118.060 122.880 ;
        RECT 120.160 118.120 120.300 139.300 ;
        RECT 121.540 139.300 122.200 139.440 ;
        RECT 121.540 137.500 121.680 139.300 ;
        RECT 121.940 139.220 122.200 139.300 ;
        RECT 123.380 138.520 123.520 141.940 ;
        RECT 124.700 141.600 124.960 141.920 ;
        RECT 124.760 139.200 124.900 141.600 ;
        RECT 135.630 141.200 136.780 141.270 ;
        RECT 135.630 140.180 136.800 141.200 ;
        RECT 124.700 138.940 124.960 139.200 ;
        RECT 124.300 138.880 124.960 138.940 ;
        RECT 124.300 138.800 124.900 138.880 ;
        RECT 123.320 138.200 123.580 138.520 ;
        RECT 121.880 137.665 123.760 138.035 ;
        RECT 121.480 137.180 121.740 137.500 ;
        RECT 121.880 132.225 123.760 132.595 ;
        RECT 122.860 130.040 123.120 130.360 ;
        RECT 122.920 128.660 123.060 130.040 ;
        RECT 124.300 128.660 124.440 138.800 ;
        RECT 124.700 138.200 124.960 138.520 ;
        RECT 124.760 137.500 124.900 138.200 ;
        RECT 129.140 138.175 134.100 139.455 ;
        RECT 124.700 137.180 124.960 137.500 ;
        RECT 135.640 133.320 136.800 140.180 ;
        RECT 122.860 128.340 123.120 128.660 ;
        RECT 124.240 128.340 124.500 128.660 ;
        RECT 121.880 126.785 123.760 127.155 ;
        RECT 124.300 125.600 124.440 128.340 ;
        RECT 124.240 125.280 124.500 125.600 ;
        RECT 121.880 121.345 123.760 121.715 ;
        RECT 124.300 120.160 124.440 125.280 ;
        RECT 124.240 119.840 124.500 120.160 ;
        RECT 120.100 117.800 120.360 118.120 ;
        RECT 116.880 117.460 117.140 117.780 ;
        RECT 115.960 117.120 116.220 117.440 ;
        RECT 116.940 114.720 117.080 117.460 ;
        RECT 124.700 116.780 124.960 117.100 ;
        RECT 119.640 116.440 119.900 116.760 ;
        RECT 121.480 116.440 121.740 116.760 ;
        RECT 116.880 114.400 117.140 114.720 ;
        RECT 116.940 112.340 117.080 114.400 ;
        RECT 118.260 112.700 118.520 113.020 ;
        RECT 110.440 112.020 110.700 112.340 ;
        RECT 111.360 112.020 111.620 112.340 ;
        RECT 114.580 112.020 114.840 112.340 ;
        RECT 116.880 112.020 117.140 112.340 ;
        RECT 114.120 111.680 114.380 112.000 ;
        RECT 116.420 111.680 116.680 112.000 ;
        RECT 112.280 111.000 112.540 111.320 ;
        RECT 112.340 109.620 112.480 111.000 ;
        RECT 114.180 109.620 114.320 111.680 ;
        RECT 112.280 109.300 112.540 109.620 ;
        RECT 114.120 109.300 114.380 109.620 ;
        RECT 116.480 109.280 116.620 111.680 ;
        RECT 118.320 109.620 118.460 112.700 ;
        RECT 119.700 112.680 119.840 116.440 ;
        RECT 121.540 115.060 121.680 116.440 ;
        RECT 121.880 115.905 123.760 116.275 ;
        RECT 121.480 114.740 121.740 115.060 ;
        RECT 124.760 112.680 124.900 116.780 ;
        RECT 126.540 113.720 126.800 114.040 ;
        RECT 119.640 112.360 119.900 112.680 ;
        RECT 124.700 112.360 124.960 112.680 ;
        RECT 121.020 111.680 121.280 112.000 ;
        RECT 124.700 111.680 124.960 112.000 ;
        RECT 118.260 109.300 118.520 109.620 ;
        RECT 116.420 108.960 116.680 109.280 ;
        RECT 109.060 108.620 109.320 108.940 ;
        RECT 109.520 108.280 109.780 108.600 ;
        RECT 115.500 108.280 115.760 108.600 ;
        RECT 106.880 107.745 108.760 108.115 ;
        RECT 109.580 107.660 109.720 108.280 ;
        RECT 109.580 107.520 110.180 107.660 ;
        RECT 110.040 94.980 110.180 107.520 ;
        RECT 115.560 94.980 115.700 108.280 ;
        RECT 121.080 94.980 121.220 111.680 ;
        RECT 124.240 111.000 124.500 111.320 ;
        RECT 121.880 110.465 123.760 110.835 ;
        RECT 124.300 109.960 124.440 111.000 ;
        RECT 124.760 110.300 124.900 111.680 ;
        RECT 124.700 109.980 124.960 110.300 ;
        RECT 124.240 109.640 124.500 109.960 ;
        RECT 121.880 105.025 123.760 105.395 ;
        RECT 126.600 94.980 126.740 113.720 ;
        RECT 131.130 111.485 131.410 111.855 ;
        RECT 131.200 109.280 131.340 111.485 ;
        RECT 131.140 108.960 131.400 109.280 ;
        RECT 129.750 105.580 133.160 106.650 ;
        RECT 31.380 94.600 32.440 94.740 ;
        RECT 32.690 92.980 32.970 94.980 ;
        RECT 38.210 92.980 38.490 94.980 ;
        RECT 43.730 92.980 44.010 94.980 ;
        RECT 49.250 92.980 49.530 94.980 ;
        RECT 54.770 92.980 55.050 94.980 ;
        RECT 60.290 92.980 60.570 94.980 ;
        RECT 65.810 92.980 66.090 94.980 ;
        RECT 71.330 92.980 71.610 94.980 ;
        RECT 76.850 92.980 77.130 94.980 ;
        RECT 82.370 92.980 82.650 94.980 ;
        RECT 87.890 92.980 88.170 94.980 ;
        RECT 93.410 92.980 93.690 94.980 ;
        RECT 98.930 92.980 99.210 94.980 ;
        RECT 104.450 92.980 104.730 94.980 ;
        RECT 109.970 92.980 110.250 94.980 ;
        RECT 115.490 92.980 115.770 94.980 ;
        RECT 121.010 92.980 121.290 94.980 ;
        RECT 126.530 92.980 126.810 94.980 ;
        RECT 13.920 85.550 15.140 89.420 ;
        RECT 19.910 85.980 21.130 89.850 ;
        RECT 67.730 89.640 68.670 89.840 ;
        RECT 25.730 85.120 26.950 88.990 ;
        RECT 31.780 85.510 33.000 89.380 ;
        RECT 37.750 88.780 38.970 89.290 ;
        RECT 37.680 88.620 38.970 88.780 ;
        RECT 43.810 88.630 45.030 89.530 ;
        RECT 49.740 88.640 50.960 89.040 ;
        RECT 37.680 86.810 39.070 88.620 ;
        RECT 37.750 85.420 38.970 86.810 ;
        RECT 43.810 86.720 45.140 88.630 ;
        RECT 49.740 86.920 51.010 88.640 ;
        RECT 43.810 85.660 45.030 86.720 ;
        RECT 49.740 85.170 50.960 86.920 ;
        RECT 55.530 85.320 56.750 89.190 ;
        RECT 61.720 88.640 62.940 88.870 ;
        RECT 61.720 86.600 63.130 88.640 ;
        RECT 61.720 85.000 62.940 86.600 ;
        RECT 67.580 85.770 68.800 89.640 ;
        RECT 73.850 84.290 75.070 88.160 ;
        RECT 79.730 84.310 80.950 88.180 ;
        RECT 74.090 80.440 74.370 84.290 ;
        RECT 20.140 80.160 74.370 80.440 ;
        RECT 20.140 75.650 20.420 80.160 ;
        RECT 80.070 79.800 80.350 84.310 ;
        RECT 85.470 84.100 86.690 87.970 ;
        RECT 91.460 84.500 92.680 88.320 ;
        RECT 97.600 84.630 98.820 88.500 ;
        RECT 103.650 84.740 104.870 88.610 ;
        RECT 109.620 85.420 110.840 89.290 ;
        RECT 115.740 85.700 116.960 89.570 ;
        RECT 121.520 85.700 122.740 89.570 ;
        RECT 31.380 79.520 80.350 79.800 ;
        RECT 31.380 75.850 31.660 79.520 ;
        RECT 86.050 79.170 86.330 84.100 ;
        RECT 42.510 78.890 86.330 79.170 ;
        RECT 3.960 71.320 6.050 73.240 ;
        RECT 19.330 73.120 21.890 75.650 ;
        RECT 28.185 73.180 30.255 74.460 ;
        RECT 30.670 73.320 33.230 75.850 ;
        RECT 42.510 75.750 42.790 78.890 ;
        RECT 92.030 78.570 92.310 84.500 ;
        RECT 53.830 78.290 92.310 78.570 ;
        RECT 53.830 75.820 54.110 78.290 ;
        RECT 98.010 77.990 98.290 84.630 ;
        RECT 64.900 77.710 98.290 77.990 ;
        RECT 19.005 71.800 19.865 72.640 ;
        RECT 15.560 68.610 16.990 71.210 ;
        RECT 19.305 68.570 19.845 71.800 ;
        RECT 20.145 70.600 20.555 73.120 ;
        RECT 30.205 71.810 31.065 72.650 ;
        RECT 19.325 47.770 19.825 68.570 ;
        RECT 20.165 49.090 20.555 70.600 ;
        RECT 20.955 70.010 21.845 70.740 ;
        RECT 21.055 65.190 21.315 70.010 ;
        RECT 22.695 68.620 25.405 69.470 ;
        RECT 22.895 65.840 24.825 68.620 ;
        RECT 30.505 68.580 31.045 71.810 ;
        RECT 31.345 70.610 31.755 73.320 ;
        RECT 39.475 73.150 41.545 74.430 ;
        RECT 41.910 73.220 44.470 75.750 ;
        RECT 41.425 71.780 42.285 72.620 ;
        RECT 27.795 67.130 28.915 67.810 ;
        RECT 28.075 65.850 28.745 67.130 ;
        RECT 21.455 65.460 26.505 65.840 ;
        RECT 27.865 65.440 28.915 65.850 ;
        RECT 21.055 63.640 21.435 65.190 ;
        RECT 21.175 55.800 21.435 63.640 ;
        RECT 26.485 63.200 26.755 65.240 ;
        RECT 27.615 63.200 27.885 65.200 ;
        RECT 26.485 56.510 27.885 63.200 ;
        RECT 21.085 55.290 21.445 55.800 ;
        RECT 21.065 54.860 21.445 55.290 ;
        RECT 26.485 55.190 26.755 56.510 ;
        RECT 27.615 55.150 27.885 56.510 ;
        RECT 28.885 55.260 29.205 65.190 ;
        RECT 28.885 55.200 29.215 55.260 ;
        RECT 21.065 54.580 21.315 54.860 ;
        RECT 20.865 54.180 25.505 54.580 ;
        RECT 26.405 54.290 27.535 54.300 ;
        RECT 28.895 54.290 29.215 55.200 ;
        RECT 21.065 52.060 21.315 54.180 ;
        RECT 25.765 53.490 26.125 54.110 ;
        RECT 25.845 52.610 26.105 53.490 ;
        RECT 26.385 53.240 29.215 54.290 ;
        RECT 25.675 52.230 26.205 52.610 ;
        RECT 21.065 51.970 21.565 52.060 ;
        RECT 21.055 51.240 21.565 51.970 ;
        RECT 21.295 50.240 21.565 51.240 ;
        RECT 22.205 50.990 22.475 51.940 ;
        RECT 22.205 50.840 22.675 50.990 ;
        RECT 22.205 50.160 22.765 50.840 ;
        RECT 22.285 50.150 22.765 50.160 ;
        RECT 21.575 49.620 22.195 49.980 ;
        RECT 21.615 49.090 22.045 49.620 ;
        RECT 20.165 48.670 22.045 49.090 ;
        RECT 22.535 48.960 22.765 50.150 ;
        RECT 21.615 47.800 22.045 48.670 ;
        RECT 22.455 48.360 22.835 48.960 ;
        RECT 19.325 47.060 20.015 47.770 ;
        RECT 21.435 47.440 22.055 47.800 ;
        RECT 21.135 47.060 21.425 47.250 ;
        RECT 19.325 46.620 21.425 47.060 ;
        RECT 19.325 46.600 20.015 46.620 ;
        RECT 21.135 46.380 21.425 46.620 ;
        RECT 22.055 46.990 22.325 47.240 ;
        RECT 22.535 46.990 22.765 48.360 ;
        RECT 25.355 47.010 25.685 52.030 ;
        RECT 26.405 52.020 27.535 53.240 ;
        RECT 28.895 53.220 29.215 53.240 ;
        RECT 22.055 46.880 22.765 46.990 ;
        RECT 25.345 46.960 25.685 47.010 ;
        RECT 26.235 47.780 27.615 52.020 ;
        RECT 22.055 46.570 22.715 46.880 ;
        RECT 22.055 46.400 22.325 46.570 ;
        RECT 25.345 45.000 25.625 46.960 ;
        RECT 26.235 46.920 26.535 47.780 ;
        RECT 27.315 46.920 27.615 47.780 ;
        RECT 28.165 46.920 28.495 51.990 ;
        RECT 27.565 46.380 28.045 46.760 ;
        RECT 27.665 45.760 27.915 46.380 ;
        RECT 27.565 45.160 27.945 45.760 ;
        RECT 24.825 44.230 25.925 45.000 ;
        RECT 28.215 44.930 28.495 46.920 ;
        RECT 30.525 47.780 31.025 68.580 ;
        RECT 31.365 49.100 31.755 70.610 ;
        RECT 32.155 70.020 33.045 70.750 ;
        RECT 32.255 65.200 32.515 70.020 ;
        RECT 33.895 68.630 36.605 69.480 ;
        RECT 34.095 65.850 36.025 68.630 ;
        RECT 41.725 68.550 42.265 71.780 ;
        RECT 42.565 70.580 42.975 73.220 ;
        RECT 50.055 73.090 52.125 74.370 ;
        RECT 53.150 73.290 55.710 75.820 ;
        RECT 64.900 75.810 65.180 77.710 ;
        RECT 103.990 77.230 104.270 84.740 ;
        RECT 76.140 76.950 104.270 77.230 ;
        RECT 52.675 71.760 53.535 72.600 ;
        RECT 38.995 67.140 40.115 67.820 ;
        RECT 39.275 65.860 39.945 67.140 ;
        RECT 32.655 65.470 37.705 65.850 ;
        RECT 39.065 65.450 40.115 65.860 ;
        RECT 32.255 63.650 32.635 65.200 ;
        RECT 32.375 55.810 32.635 63.650 ;
        RECT 37.685 63.210 37.955 65.250 ;
        RECT 38.815 63.210 39.085 65.210 ;
        RECT 37.685 56.520 39.085 63.210 ;
        RECT 32.285 55.300 32.645 55.810 ;
        RECT 32.265 54.870 32.645 55.300 ;
        RECT 37.685 55.200 37.955 56.520 ;
        RECT 38.815 55.160 39.085 56.520 ;
        RECT 40.085 55.270 40.405 65.200 ;
        RECT 40.085 55.210 40.415 55.270 ;
        RECT 32.265 54.590 32.515 54.870 ;
        RECT 32.065 54.190 36.705 54.590 ;
        RECT 37.605 54.300 38.735 54.310 ;
        RECT 40.095 54.300 40.415 55.210 ;
        RECT 32.265 52.070 32.515 54.190 ;
        RECT 36.965 53.500 37.325 54.120 ;
        RECT 37.045 52.620 37.305 53.500 ;
        RECT 37.585 53.250 40.415 54.300 ;
        RECT 36.875 52.240 37.405 52.620 ;
        RECT 32.265 51.980 32.765 52.070 ;
        RECT 32.255 51.250 32.765 51.980 ;
        RECT 32.495 50.250 32.765 51.250 ;
        RECT 33.405 51.000 33.675 51.950 ;
        RECT 33.405 50.850 33.875 51.000 ;
        RECT 33.405 50.170 33.965 50.850 ;
        RECT 33.485 50.160 33.965 50.170 ;
        RECT 32.775 49.630 33.395 49.990 ;
        RECT 32.815 49.100 33.245 49.630 ;
        RECT 31.365 48.680 33.245 49.100 ;
        RECT 33.735 48.970 33.965 50.160 ;
        RECT 32.815 47.810 33.245 48.680 ;
        RECT 33.655 48.370 34.035 48.970 ;
        RECT 30.525 47.070 31.215 47.780 ;
        RECT 32.635 47.450 33.255 47.810 ;
        RECT 32.335 47.070 32.625 47.260 ;
        RECT 30.525 46.630 32.625 47.070 ;
        RECT 30.525 46.610 31.215 46.630 ;
        RECT 32.335 46.390 32.625 46.630 ;
        RECT 33.255 47.000 33.525 47.250 ;
        RECT 33.735 47.000 33.965 48.370 ;
        RECT 36.555 47.020 36.885 52.040 ;
        RECT 37.605 52.030 38.735 53.250 ;
        RECT 40.095 53.230 40.415 53.250 ;
        RECT 33.255 46.890 33.965 47.000 ;
        RECT 36.545 46.970 36.885 47.020 ;
        RECT 37.435 47.790 38.815 52.030 ;
        RECT 33.255 46.580 33.915 46.890 ;
        RECT 33.255 46.410 33.525 46.580 ;
        RECT 36.545 45.010 36.825 46.970 ;
        RECT 37.435 46.930 37.735 47.790 ;
        RECT 38.515 46.930 38.815 47.790 ;
        RECT 39.365 46.930 39.695 52.000 ;
        RECT 38.765 46.390 39.245 46.770 ;
        RECT 38.865 45.770 39.115 46.390 ;
        RECT 38.765 45.170 39.145 45.770 ;
        RECT 28.215 43.200 28.515 44.930 ;
        RECT 36.025 44.240 37.125 45.010 ;
        RECT 39.415 44.940 39.695 46.930 ;
        RECT 41.745 47.750 42.245 68.550 ;
        RECT 42.585 49.070 42.975 70.580 ;
        RECT 43.375 69.990 44.265 70.720 ;
        RECT 43.475 65.170 43.735 69.990 ;
        RECT 45.115 68.600 47.825 69.450 ;
        RECT 45.315 65.820 47.245 68.600 ;
        RECT 52.975 68.530 53.515 71.760 ;
        RECT 53.815 70.560 54.225 73.290 ;
        RECT 61.475 73.120 63.545 74.400 ;
        RECT 64.400 73.280 66.960 75.810 ;
        RECT 76.140 75.740 76.420 76.950 ;
        RECT 109.970 76.610 110.250 85.420 ;
        RECT 87.580 76.330 110.250 76.610 ;
        RECT 87.580 75.760 87.860 76.330 ;
        RECT 115.950 76.030 116.230 85.700 ;
        RECT 98.850 75.840 116.230 76.030 ;
        RECT 63.895 71.750 64.755 72.590 ;
        RECT 50.215 67.110 51.335 67.790 ;
        RECT 50.495 65.830 51.165 67.110 ;
        RECT 43.875 65.440 48.925 65.820 ;
        RECT 50.285 65.420 51.335 65.830 ;
        RECT 43.475 63.620 43.855 65.170 ;
        RECT 43.595 55.780 43.855 63.620 ;
        RECT 48.905 63.180 49.175 65.220 ;
        RECT 50.035 63.180 50.305 65.180 ;
        RECT 48.905 56.490 50.305 63.180 ;
        RECT 43.505 55.270 43.865 55.780 ;
        RECT 43.485 54.840 43.865 55.270 ;
        RECT 48.905 55.170 49.175 56.490 ;
        RECT 50.035 55.130 50.305 56.490 ;
        RECT 51.305 55.240 51.625 65.170 ;
        RECT 51.305 55.180 51.635 55.240 ;
        RECT 43.485 54.560 43.735 54.840 ;
        RECT 43.285 54.160 47.925 54.560 ;
        RECT 48.825 54.270 49.955 54.280 ;
        RECT 51.315 54.270 51.635 55.180 ;
        RECT 43.485 52.040 43.735 54.160 ;
        RECT 48.185 53.470 48.545 54.090 ;
        RECT 48.265 52.590 48.525 53.470 ;
        RECT 48.805 53.220 51.635 54.270 ;
        RECT 48.095 52.210 48.625 52.590 ;
        RECT 43.485 51.950 43.985 52.040 ;
        RECT 43.475 51.220 43.985 51.950 ;
        RECT 43.715 50.220 43.985 51.220 ;
        RECT 44.625 50.970 44.895 51.920 ;
        RECT 44.625 50.820 45.095 50.970 ;
        RECT 44.625 50.140 45.185 50.820 ;
        RECT 44.705 50.130 45.185 50.140 ;
        RECT 43.995 49.600 44.615 49.960 ;
        RECT 44.035 49.070 44.465 49.600 ;
        RECT 42.585 48.650 44.465 49.070 ;
        RECT 44.955 48.940 45.185 50.130 ;
        RECT 44.035 47.780 44.465 48.650 ;
        RECT 44.875 48.340 45.255 48.940 ;
        RECT 41.745 47.040 42.435 47.750 ;
        RECT 43.855 47.420 44.475 47.780 ;
        RECT 43.555 47.040 43.845 47.230 ;
        RECT 41.745 46.600 43.845 47.040 ;
        RECT 41.745 46.580 42.435 46.600 ;
        RECT 43.555 46.360 43.845 46.600 ;
        RECT 44.475 46.970 44.745 47.220 ;
        RECT 44.955 46.970 45.185 48.340 ;
        RECT 47.775 46.990 48.105 52.010 ;
        RECT 48.825 52.000 49.955 53.220 ;
        RECT 51.315 53.200 51.635 53.220 ;
        RECT 44.475 46.860 45.185 46.970 ;
        RECT 47.765 46.940 48.105 46.990 ;
        RECT 48.655 47.760 50.035 52.000 ;
        RECT 44.475 46.550 45.135 46.860 ;
        RECT 44.475 46.380 44.745 46.550 ;
        RECT 47.765 44.980 48.045 46.940 ;
        RECT 48.655 46.900 48.955 47.760 ;
        RECT 49.735 46.900 50.035 47.760 ;
        RECT 50.585 46.900 50.915 51.970 ;
        RECT 49.985 46.360 50.465 46.740 ;
        RECT 50.085 45.740 50.335 46.360 ;
        RECT 49.985 45.140 50.365 45.740 ;
        RECT 39.415 43.210 39.715 44.940 ;
        RECT 47.245 44.210 48.345 44.980 ;
        RECT 50.635 44.910 50.915 46.900 ;
        RECT 52.995 47.730 53.495 68.530 ;
        RECT 53.835 49.050 54.225 70.560 ;
        RECT 54.625 69.970 55.515 70.700 ;
        RECT 54.725 65.150 54.985 69.970 ;
        RECT 56.365 68.580 59.075 69.430 ;
        RECT 56.565 65.800 58.495 68.580 ;
        RECT 64.195 68.520 64.735 71.750 ;
        RECT 65.035 70.550 65.445 73.280 ;
        RECT 72.585 73.130 74.655 74.410 ;
        RECT 75.550 73.210 78.110 75.740 ;
        RECT 75.135 71.740 75.995 72.580 ;
        RECT 61.465 67.090 62.585 67.770 ;
        RECT 61.745 65.810 62.415 67.090 ;
        RECT 55.125 65.420 60.175 65.800 ;
        RECT 61.535 65.400 62.585 65.810 ;
        RECT 54.725 63.600 55.105 65.150 ;
        RECT 54.845 55.760 55.105 63.600 ;
        RECT 60.155 63.160 60.425 65.200 ;
        RECT 61.285 63.160 61.555 65.160 ;
        RECT 60.155 56.470 61.555 63.160 ;
        RECT 54.755 55.250 55.115 55.760 ;
        RECT 54.735 54.820 55.115 55.250 ;
        RECT 60.155 55.150 60.425 56.470 ;
        RECT 61.285 55.110 61.555 56.470 ;
        RECT 62.555 55.220 62.875 65.150 ;
        RECT 62.555 55.160 62.885 55.220 ;
        RECT 54.735 54.540 54.985 54.820 ;
        RECT 54.535 54.140 59.175 54.540 ;
        RECT 60.075 54.250 61.205 54.260 ;
        RECT 62.565 54.250 62.885 55.160 ;
        RECT 54.735 52.020 54.985 54.140 ;
        RECT 59.435 53.450 59.795 54.070 ;
        RECT 59.515 52.570 59.775 53.450 ;
        RECT 60.055 53.200 62.885 54.250 ;
        RECT 59.345 52.190 59.875 52.570 ;
        RECT 54.735 51.930 55.235 52.020 ;
        RECT 54.725 51.200 55.235 51.930 ;
        RECT 54.965 50.200 55.235 51.200 ;
        RECT 55.875 50.950 56.145 51.900 ;
        RECT 55.875 50.800 56.345 50.950 ;
        RECT 55.875 50.120 56.435 50.800 ;
        RECT 55.955 50.110 56.435 50.120 ;
        RECT 55.245 49.580 55.865 49.940 ;
        RECT 55.285 49.050 55.715 49.580 ;
        RECT 53.835 48.630 55.715 49.050 ;
        RECT 56.205 48.920 56.435 50.110 ;
        RECT 55.285 47.760 55.715 48.630 ;
        RECT 56.125 48.320 56.505 48.920 ;
        RECT 52.995 47.020 53.685 47.730 ;
        RECT 55.105 47.400 55.725 47.760 ;
        RECT 54.805 47.020 55.095 47.210 ;
        RECT 52.995 46.580 55.095 47.020 ;
        RECT 52.995 46.560 53.685 46.580 ;
        RECT 54.805 46.340 55.095 46.580 ;
        RECT 55.725 46.950 55.995 47.200 ;
        RECT 56.205 46.950 56.435 48.320 ;
        RECT 59.025 46.970 59.355 51.990 ;
        RECT 60.075 51.980 61.205 53.200 ;
        RECT 62.565 53.180 62.885 53.200 ;
        RECT 55.725 46.840 56.435 46.950 ;
        RECT 59.015 46.920 59.355 46.970 ;
        RECT 59.905 47.740 61.285 51.980 ;
        RECT 55.725 46.530 56.385 46.840 ;
        RECT 55.725 46.360 55.995 46.530 ;
        RECT 59.015 44.960 59.295 46.920 ;
        RECT 59.905 46.880 60.205 47.740 ;
        RECT 60.985 46.880 61.285 47.740 ;
        RECT 61.835 46.880 62.165 51.950 ;
        RECT 61.235 46.340 61.715 46.720 ;
        RECT 61.335 45.720 61.585 46.340 ;
        RECT 61.235 45.120 61.615 45.720 ;
        RECT 19.865 42.210 21.245 42.780 ;
        RECT 27.495 42.630 28.875 43.200 ;
        RECT 31.145 42.210 32.525 42.780 ;
        RECT 38.695 42.640 40.075 43.210 ;
        RECT 50.635 43.180 50.935 44.910 ;
        RECT 58.495 44.190 59.595 44.960 ;
        RECT 61.885 44.890 62.165 46.880 ;
        RECT 64.215 47.720 64.715 68.520 ;
        RECT 65.055 49.040 65.445 70.550 ;
        RECT 65.845 69.960 66.735 70.690 ;
        RECT 65.945 65.140 66.205 69.960 ;
        RECT 67.585 68.570 70.295 69.420 ;
        RECT 67.785 65.790 69.715 68.570 ;
        RECT 75.435 68.510 75.975 71.740 ;
        RECT 76.275 70.540 76.685 73.210 ;
        RECT 83.855 73.120 85.925 74.400 ;
        RECT 86.850 73.230 89.410 75.760 ;
        RECT 98.150 75.750 116.230 75.840 ;
        RECT 86.385 71.750 87.245 72.590 ;
        RECT 72.685 67.080 73.805 67.760 ;
        RECT 72.965 65.800 73.635 67.080 ;
        RECT 66.345 65.410 71.395 65.790 ;
        RECT 72.755 65.390 73.805 65.800 ;
        RECT 65.945 63.590 66.325 65.140 ;
        RECT 66.065 55.750 66.325 63.590 ;
        RECT 71.375 63.150 71.645 65.190 ;
        RECT 72.505 63.150 72.775 65.150 ;
        RECT 71.375 56.460 72.775 63.150 ;
        RECT 65.975 55.240 66.335 55.750 ;
        RECT 65.955 54.810 66.335 55.240 ;
        RECT 71.375 55.140 71.645 56.460 ;
        RECT 72.505 55.100 72.775 56.460 ;
        RECT 73.775 55.210 74.095 65.140 ;
        RECT 73.775 55.150 74.105 55.210 ;
        RECT 65.955 54.530 66.205 54.810 ;
        RECT 65.755 54.130 70.395 54.530 ;
        RECT 71.295 54.240 72.425 54.250 ;
        RECT 73.785 54.240 74.105 55.150 ;
        RECT 65.955 52.010 66.205 54.130 ;
        RECT 70.655 53.440 71.015 54.060 ;
        RECT 70.735 52.560 70.995 53.440 ;
        RECT 71.275 53.190 74.105 54.240 ;
        RECT 70.565 52.180 71.095 52.560 ;
        RECT 65.955 51.920 66.455 52.010 ;
        RECT 65.945 51.190 66.455 51.920 ;
        RECT 66.185 50.190 66.455 51.190 ;
        RECT 67.095 50.940 67.365 51.890 ;
        RECT 67.095 50.790 67.565 50.940 ;
        RECT 67.095 50.110 67.655 50.790 ;
        RECT 67.175 50.100 67.655 50.110 ;
        RECT 66.465 49.570 67.085 49.930 ;
        RECT 66.505 49.040 66.935 49.570 ;
        RECT 65.055 48.620 66.935 49.040 ;
        RECT 67.425 48.910 67.655 50.100 ;
        RECT 66.505 47.750 66.935 48.620 ;
        RECT 67.345 48.310 67.725 48.910 ;
        RECT 64.215 47.010 64.905 47.720 ;
        RECT 66.325 47.390 66.945 47.750 ;
        RECT 66.025 47.010 66.315 47.200 ;
        RECT 64.215 46.570 66.315 47.010 ;
        RECT 64.215 46.550 64.905 46.570 ;
        RECT 66.025 46.330 66.315 46.570 ;
        RECT 66.945 46.940 67.215 47.190 ;
        RECT 67.425 46.940 67.655 48.310 ;
        RECT 70.245 46.960 70.575 51.980 ;
        RECT 71.295 51.970 72.425 53.190 ;
        RECT 73.785 53.170 74.105 53.190 ;
        RECT 66.945 46.830 67.655 46.940 ;
        RECT 70.235 46.910 70.575 46.960 ;
        RECT 71.125 47.730 72.505 51.970 ;
        RECT 66.945 46.520 67.605 46.830 ;
        RECT 66.945 46.350 67.215 46.520 ;
        RECT 70.235 44.950 70.515 46.910 ;
        RECT 71.125 46.870 71.425 47.730 ;
        RECT 72.205 46.870 72.505 47.730 ;
        RECT 73.055 46.870 73.385 51.940 ;
        RECT 72.455 46.330 72.935 46.710 ;
        RECT 72.555 45.710 72.805 46.330 ;
        RECT 72.455 45.110 72.835 45.710 ;
        RECT 20.225 40.480 20.525 42.210 ;
        RECT 20.245 38.490 20.525 40.480 ;
        RECT 22.815 40.410 23.915 41.180 ;
        RECT 31.505 40.480 31.805 42.210 ;
        RECT 42.435 42.190 43.815 42.760 ;
        RECT 49.915 42.610 51.295 43.180 ;
        RECT 61.885 43.160 62.185 44.890 ;
        RECT 69.715 44.180 70.815 44.950 ;
        RECT 73.105 44.880 73.385 46.870 ;
        RECT 75.455 47.710 75.955 68.510 ;
        RECT 76.295 49.030 76.685 70.540 ;
        RECT 77.085 69.950 77.975 70.680 ;
        RECT 77.185 65.130 77.445 69.950 ;
        RECT 78.825 68.560 81.535 69.410 ;
        RECT 79.025 65.780 80.955 68.560 ;
        RECT 86.685 68.520 87.225 71.750 ;
        RECT 87.525 70.550 87.935 73.230 ;
        RECT 95.045 73.060 97.115 74.340 ;
        RECT 98.150 73.310 100.710 75.750 ;
        RECT 109.390 75.480 111.950 75.560 ;
        RECT 121.930 75.480 122.210 85.700 ;
        RECT 127.550 85.510 128.770 89.380 ;
        RECT 127.910 76.040 128.190 85.510 ;
        RECT 133.380 76.580 136.010 77.880 ;
        RECT 137.240 76.560 139.870 77.860 ;
        RECT 109.390 75.200 122.210 75.480 ;
        RECT 97.665 71.740 98.525 72.580 ;
        RECT 83.925 67.070 85.045 67.750 ;
        RECT 84.205 65.790 84.875 67.070 ;
        RECT 77.585 65.400 82.635 65.780 ;
        RECT 83.995 65.380 85.045 65.790 ;
        RECT 77.185 63.580 77.565 65.130 ;
        RECT 77.305 55.740 77.565 63.580 ;
        RECT 82.615 63.140 82.885 65.180 ;
        RECT 83.745 63.140 84.015 65.140 ;
        RECT 82.615 56.450 84.015 63.140 ;
        RECT 77.215 55.230 77.575 55.740 ;
        RECT 77.195 54.800 77.575 55.230 ;
        RECT 82.615 55.130 82.885 56.450 ;
        RECT 83.745 55.090 84.015 56.450 ;
        RECT 85.015 55.200 85.335 65.130 ;
        RECT 85.015 55.140 85.345 55.200 ;
        RECT 77.195 54.520 77.445 54.800 ;
        RECT 76.995 54.120 81.635 54.520 ;
        RECT 82.535 54.230 83.665 54.240 ;
        RECT 85.025 54.230 85.345 55.140 ;
        RECT 77.195 52.000 77.445 54.120 ;
        RECT 81.895 53.430 82.255 54.050 ;
        RECT 81.975 52.550 82.235 53.430 ;
        RECT 82.515 53.180 85.345 54.230 ;
        RECT 81.805 52.170 82.335 52.550 ;
        RECT 77.195 51.910 77.695 52.000 ;
        RECT 77.185 51.180 77.695 51.910 ;
        RECT 77.425 50.180 77.695 51.180 ;
        RECT 78.335 50.930 78.605 51.880 ;
        RECT 78.335 50.780 78.805 50.930 ;
        RECT 78.335 50.100 78.895 50.780 ;
        RECT 78.415 50.090 78.895 50.100 ;
        RECT 77.705 49.560 78.325 49.920 ;
        RECT 77.745 49.030 78.175 49.560 ;
        RECT 76.295 48.610 78.175 49.030 ;
        RECT 78.665 48.900 78.895 50.090 ;
        RECT 77.745 47.740 78.175 48.610 ;
        RECT 78.585 48.300 78.965 48.900 ;
        RECT 75.455 47.000 76.145 47.710 ;
        RECT 77.565 47.380 78.185 47.740 ;
        RECT 77.265 47.000 77.555 47.190 ;
        RECT 75.455 46.560 77.555 47.000 ;
        RECT 75.455 46.540 76.145 46.560 ;
        RECT 77.265 46.320 77.555 46.560 ;
        RECT 78.185 46.930 78.455 47.180 ;
        RECT 78.665 46.930 78.895 48.300 ;
        RECT 81.485 46.950 81.815 51.970 ;
        RECT 82.535 51.960 83.665 53.180 ;
        RECT 85.025 53.160 85.345 53.180 ;
        RECT 78.185 46.820 78.895 46.930 ;
        RECT 81.475 46.900 81.815 46.950 ;
        RECT 82.365 47.720 83.745 51.960 ;
        RECT 78.185 46.510 78.845 46.820 ;
        RECT 78.185 46.340 78.455 46.510 ;
        RECT 81.475 44.940 81.755 46.900 ;
        RECT 82.365 46.860 82.665 47.720 ;
        RECT 83.445 46.860 83.745 47.720 ;
        RECT 84.295 46.860 84.625 51.930 ;
        RECT 83.695 46.320 84.175 46.700 ;
        RECT 83.795 45.700 84.045 46.320 ;
        RECT 83.695 45.100 84.075 45.700 ;
        RECT 53.655 42.190 55.035 42.760 ;
        RECT 61.165 42.590 62.545 43.160 ;
        RECT 73.105 43.150 73.405 44.880 ;
        RECT 80.955 44.170 82.055 44.940 ;
        RECT 84.345 44.870 84.625 46.860 ;
        RECT 86.705 47.720 87.205 68.520 ;
        RECT 87.545 49.040 87.935 70.550 ;
        RECT 88.335 69.960 89.225 70.690 ;
        RECT 88.435 65.140 88.695 69.960 ;
        RECT 90.075 68.570 92.785 69.420 ;
        RECT 90.275 65.790 92.205 68.570 ;
        RECT 97.965 68.510 98.505 71.740 ;
        RECT 98.805 70.540 99.215 73.310 ;
        RECT 106.455 73.110 108.525 74.390 ;
        RECT 109.390 73.030 111.950 75.200 ;
        RECT 125.760 74.810 128.190 76.040 ;
        RECT 121.290 74.790 128.190 74.810 ;
        RECT 120.600 74.530 128.190 74.790 ;
        RECT 117.655 73.110 119.725 74.390 ;
        RECT 120.600 73.180 128.160 74.530 ;
        RECT 129.505 73.190 131.575 74.470 ;
        RECT 120.600 73.110 126.160 73.180 ;
        RECT 108.935 71.740 109.795 72.580 ;
        RECT 95.175 67.080 96.295 67.760 ;
        RECT 95.455 65.800 96.125 67.080 ;
        RECT 88.835 65.410 93.885 65.790 ;
        RECT 95.245 65.390 96.295 65.800 ;
        RECT 88.435 63.590 88.815 65.140 ;
        RECT 88.555 55.750 88.815 63.590 ;
        RECT 93.865 63.150 94.135 65.190 ;
        RECT 94.995 63.150 95.265 65.150 ;
        RECT 93.865 56.460 95.265 63.150 ;
        RECT 88.465 55.240 88.825 55.750 ;
        RECT 88.445 54.810 88.825 55.240 ;
        RECT 93.865 55.140 94.135 56.460 ;
        RECT 94.995 55.100 95.265 56.460 ;
        RECT 96.265 55.210 96.585 65.140 ;
        RECT 96.265 55.150 96.595 55.210 ;
        RECT 88.445 54.530 88.695 54.810 ;
        RECT 88.245 54.130 92.885 54.530 ;
        RECT 93.785 54.240 94.915 54.250 ;
        RECT 96.275 54.240 96.595 55.150 ;
        RECT 88.445 52.010 88.695 54.130 ;
        RECT 93.145 53.440 93.505 54.060 ;
        RECT 93.225 52.560 93.485 53.440 ;
        RECT 93.765 53.190 96.595 54.240 ;
        RECT 93.055 52.180 93.585 52.560 ;
        RECT 88.445 51.920 88.945 52.010 ;
        RECT 88.435 51.190 88.945 51.920 ;
        RECT 88.675 50.190 88.945 51.190 ;
        RECT 89.585 50.940 89.855 51.890 ;
        RECT 89.585 50.790 90.055 50.940 ;
        RECT 89.585 50.110 90.145 50.790 ;
        RECT 89.665 50.100 90.145 50.110 ;
        RECT 88.955 49.570 89.575 49.930 ;
        RECT 88.995 49.040 89.425 49.570 ;
        RECT 87.545 48.620 89.425 49.040 ;
        RECT 89.915 48.910 90.145 50.100 ;
        RECT 88.995 47.750 89.425 48.620 ;
        RECT 89.835 48.310 90.215 48.910 ;
        RECT 86.705 47.010 87.395 47.720 ;
        RECT 88.815 47.390 89.435 47.750 ;
        RECT 88.515 47.010 88.805 47.200 ;
        RECT 86.705 46.570 88.805 47.010 ;
        RECT 86.705 46.550 87.395 46.570 ;
        RECT 88.515 46.330 88.805 46.570 ;
        RECT 89.435 46.940 89.705 47.190 ;
        RECT 89.915 46.940 90.145 48.310 ;
        RECT 92.735 46.960 93.065 51.980 ;
        RECT 93.785 51.970 94.915 53.190 ;
        RECT 96.275 53.170 96.595 53.190 ;
        RECT 89.435 46.830 90.145 46.940 ;
        RECT 92.725 46.910 93.065 46.960 ;
        RECT 93.615 47.730 94.995 51.970 ;
        RECT 89.435 46.520 90.095 46.830 ;
        RECT 89.435 46.350 89.705 46.520 ;
        RECT 92.725 44.950 93.005 46.910 ;
        RECT 93.615 46.870 93.915 47.730 ;
        RECT 94.695 46.870 94.995 47.730 ;
        RECT 95.545 46.870 95.875 51.940 ;
        RECT 94.945 46.330 95.425 46.710 ;
        RECT 95.045 45.710 95.295 46.330 ;
        RECT 94.945 45.110 95.325 45.710 ;
        RECT 64.855 42.190 66.235 42.760 ;
        RECT 72.385 42.580 73.765 43.150 ;
        RECT 84.345 43.140 84.645 44.870 ;
        RECT 92.205 44.180 93.305 44.950 ;
        RECT 95.595 44.880 95.875 46.870 ;
        RECT 97.985 47.710 98.485 68.510 ;
        RECT 98.825 49.030 99.215 70.540 ;
        RECT 99.615 69.950 100.505 70.680 ;
        RECT 99.715 65.130 99.975 69.950 ;
        RECT 101.355 68.560 104.065 69.410 ;
        RECT 101.555 65.780 103.485 68.560 ;
        RECT 109.235 68.510 109.775 71.740 ;
        RECT 110.075 70.540 110.485 73.030 ;
        RECT 120.185 71.740 121.045 72.580 ;
        RECT 106.455 67.070 107.575 67.750 ;
        RECT 106.735 65.790 107.405 67.070 ;
        RECT 100.115 65.400 105.165 65.780 ;
        RECT 106.525 65.380 107.575 65.790 ;
        RECT 99.715 63.580 100.095 65.130 ;
        RECT 99.835 55.740 100.095 63.580 ;
        RECT 105.145 63.140 105.415 65.180 ;
        RECT 106.275 63.140 106.545 65.140 ;
        RECT 105.145 56.450 106.545 63.140 ;
        RECT 99.745 55.230 100.105 55.740 ;
        RECT 99.725 54.800 100.105 55.230 ;
        RECT 105.145 55.130 105.415 56.450 ;
        RECT 106.275 55.090 106.545 56.450 ;
        RECT 107.545 55.200 107.865 65.130 ;
        RECT 107.545 55.140 107.875 55.200 ;
        RECT 99.725 54.520 99.975 54.800 ;
        RECT 99.525 54.120 104.165 54.520 ;
        RECT 105.065 54.230 106.195 54.240 ;
        RECT 107.555 54.230 107.875 55.140 ;
        RECT 99.725 52.000 99.975 54.120 ;
        RECT 104.425 53.430 104.785 54.050 ;
        RECT 104.505 52.550 104.765 53.430 ;
        RECT 105.045 53.180 107.875 54.230 ;
        RECT 104.335 52.170 104.865 52.550 ;
        RECT 99.725 51.910 100.225 52.000 ;
        RECT 99.715 51.180 100.225 51.910 ;
        RECT 99.955 50.180 100.225 51.180 ;
        RECT 100.865 50.930 101.135 51.880 ;
        RECT 100.865 50.780 101.335 50.930 ;
        RECT 100.865 50.100 101.425 50.780 ;
        RECT 100.945 50.090 101.425 50.100 ;
        RECT 100.235 49.560 100.855 49.920 ;
        RECT 100.275 49.030 100.705 49.560 ;
        RECT 98.825 48.610 100.705 49.030 ;
        RECT 101.195 48.900 101.425 50.090 ;
        RECT 100.275 47.740 100.705 48.610 ;
        RECT 101.115 48.300 101.495 48.900 ;
        RECT 97.985 47.000 98.675 47.710 ;
        RECT 100.095 47.380 100.715 47.740 ;
        RECT 99.795 47.000 100.085 47.190 ;
        RECT 97.985 46.560 100.085 47.000 ;
        RECT 97.985 46.540 98.675 46.560 ;
        RECT 99.795 46.320 100.085 46.560 ;
        RECT 100.715 46.930 100.985 47.180 ;
        RECT 101.195 46.930 101.425 48.300 ;
        RECT 104.015 46.950 104.345 51.970 ;
        RECT 105.065 51.960 106.195 53.180 ;
        RECT 107.555 53.160 107.875 53.180 ;
        RECT 100.715 46.820 101.425 46.930 ;
        RECT 104.005 46.900 104.345 46.950 ;
        RECT 104.895 47.720 106.275 51.960 ;
        RECT 100.715 46.510 101.375 46.820 ;
        RECT 100.715 46.340 100.985 46.510 ;
        RECT 104.005 44.940 104.285 46.900 ;
        RECT 104.895 46.860 105.195 47.720 ;
        RECT 105.975 46.860 106.275 47.720 ;
        RECT 106.825 46.860 107.155 51.930 ;
        RECT 106.225 46.320 106.705 46.700 ;
        RECT 106.325 45.700 106.575 46.320 ;
        RECT 106.225 45.100 106.605 45.700 ;
        RECT 95.595 43.150 95.895 44.880 ;
        RECT 103.485 44.170 104.585 44.940 ;
        RECT 106.875 44.870 107.155 46.860 ;
        RECT 109.255 47.710 109.755 68.510 ;
        RECT 110.095 49.030 110.485 70.540 ;
        RECT 110.885 69.950 111.775 70.680 ;
        RECT 110.985 65.130 111.245 69.950 ;
        RECT 112.625 68.560 115.335 69.410 ;
        RECT 112.825 65.780 114.755 68.560 ;
        RECT 120.485 68.510 121.025 71.740 ;
        RECT 121.325 70.540 121.735 73.110 ;
        RECT 132.925 70.810 133.225 70.900 ;
        RECT 117.725 67.070 118.845 67.750 ;
        RECT 118.005 65.790 118.675 67.070 ;
        RECT 111.385 65.400 116.435 65.780 ;
        RECT 117.795 65.380 118.845 65.790 ;
        RECT 110.985 63.580 111.365 65.130 ;
        RECT 111.105 55.740 111.365 63.580 ;
        RECT 116.415 63.140 116.685 65.180 ;
        RECT 117.545 63.140 117.815 65.140 ;
        RECT 116.415 56.450 117.815 63.140 ;
        RECT 111.015 55.230 111.375 55.740 ;
        RECT 110.995 54.800 111.375 55.230 ;
        RECT 116.415 55.130 116.685 56.450 ;
        RECT 117.545 55.090 117.815 56.450 ;
        RECT 118.815 55.200 119.135 65.130 ;
        RECT 118.815 55.140 119.145 55.200 ;
        RECT 110.995 54.520 111.245 54.800 ;
        RECT 110.795 54.120 115.435 54.520 ;
        RECT 116.335 54.230 117.465 54.240 ;
        RECT 118.825 54.230 119.145 55.140 ;
        RECT 110.995 52.000 111.245 54.120 ;
        RECT 115.695 53.430 116.055 54.050 ;
        RECT 115.775 52.550 116.035 53.430 ;
        RECT 116.315 53.180 119.145 54.230 ;
        RECT 115.605 52.170 116.135 52.550 ;
        RECT 110.995 51.910 111.495 52.000 ;
        RECT 110.985 51.180 111.495 51.910 ;
        RECT 111.225 50.180 111.495 51.180 ;
        RECT 112.135 50.930 112.405 51.880 ;
        RECT 112.135 50.780 112.605 50.930 ;
        RECT 112.135 50.100 112.695 50.780 ;
        RECT 112.215 50.090 112.695 50.100 ;
        RECT 111.505 49.560 112.125 49.920 ;
        RECT 111.545 49.030 111.975 49.560 ;
        RECT 110.095 48.610 111.975 49.030 ;
        RECT 112.465 48.900 112.695 50.090 ;
        RECT 111.545 47.740 111.975 48.610 ;
        RECT 112.385 48.300 112.765 48.900 ;
        RECT 109.255 47.000 109.945 47.710 ;
        RECT 111.365 47.380 111.985 47.740 ;
        RECT 111.065 47.000 111.355 47.190 ;
        RECT 109.255 46.560 111.355 47.000 ;
        RECT 109.255 46.540 109.945 46.560 ;
        RECT 111.065 46.320 111.355 46.560 ;
        RECT 111.985 46.930 112.255 47.180 ;
        RECT 112.465 46.930 112.695 48.300 ;
        RECT 115.285 46.950 115.615 51.970 ;
        RECT 116.335 51.960 117.465 53.180 ;
        RECT 118.825 53.160 119.145 53.180 ;
        RECT 111.985 46.820 112.695 46.930 ;
        RECT 115.275 46.900 115.615 46.950 ;
        RECT 116.165 47.720 117.545 51.960 ;
        RECT 111.985 46.510 112.645 46.820 ;
        RECT 111.985 46.340 112.255 46.510 ;
        RECT 115.275 44.940 115.555 46.900 ;
        RECT 116.165 46.860 116.465 47.720 ;
        RECT 117.245 46.860 117.545 47.720 ;
        RECT 118.095 46.860 118.425 51.930 ;
        RECT 117.495 46.320 117.975 46.700 ;
        RECT 117.595 45.700 117.845 46.320 ;
        RECT 117.495 45.100 117.875 45.700 ;
        RECT 20.795 39.650 21.175 40.250 ;
        RECT 20.825 39.030 21.075 39.650 ;
        RECT 20.695 38.650 21.175 39.030 ;
        RECT 20.245 33.420 20.575 38.490 ;
        RECT 21.125 37.630 21.425 38.490 ;
        RECT 22.205 37.630 22.505 38.490 ;
        RECT 23.115 38.450 23.395 40.410 ;
        RECT 26.415 38.840 26.685 39.010 ;
        RECT 26.025 38.530 26.685 38.840 ;
        RECT 21.125 33.390 22.505 37.630 ;
        RECT 23.055 38.400 23.395 38.450 ;
        RECT 25.975 38.420 26.685 38.530 ;
        RECT 19.525 32.170 19.845 32.190 ;
        RECT 21.205 32.170 22.335 33.390 ;
        RECT 23.055 33.380 23.385 38.400 ;
        RECT 25.975 37.050 26.205 38.420 ;
        RECT 26.415 38.170 26.685 38.420 ;
        RECT 27.315 38.790 27.605 39.030 ;
        RECT 28.725 38.790 29.415 38.810 ;
        RECT 27.315 38.350 29.415 38.790 ;
        RECT 27.315 38.160 27.605 38.350 ;
        RECT 26.685 37.610 27.305 37.970 ;
        RECT 28.725 37.640 29.415 38.350 ;
        RECT 25.905 36.450 26.285 37.050 ;
        RECT 26.695 36.740 27.125 37.610 ;
        RECT 25.975 35.260 26.205 36.450 ;
        RECT 26.695 36.320 28.575 36.740 ;
        RECT 26.695 35.790 27.125 36.320 ;
        RECT 26.545 35.430 27.165 35.790 ;
        RECT 25.975 35.250 26.455 35.260 ;
        RECT 25.975 34.570 26.535 35.250 ;
        RECT 26.065 34.420 26.535 34.570 ;
        RECT 26.265 33.470 26.535 34.420 ;
        RECT 27.175 34.170 27.445 35.170 ;
        RECT 27.175 33.440 27.685 34.170 ;
        RECT 27.175 33.350 27.675 33.440 ;
        RECT 22.535 32.800 23.065 33.180 ;
        RECT 19.525 31.120 22.355 32.170 ;
        RECT 22.635 31.920 22.895 32.800 ;
        RECT 22.615 31.300 22.975 31.920 ;
        RECT 27.425 31.230 27.675 33.350 ;
        RECT 19.525 30.210 19.845 31.120 ;
        RECT 21.205 31.110 22.335 31.120 ;
        RECT 23.235 30.830 27.875 31.230 ;
        RECT 27.425 30.550 27.675 30.830 ;
        RECT 19.525 30.150 19.855 30.210 ;
        RECT 19.535 20.220 19.855 30.150 ;
        RECT 20.855 28.900 21.125 30.260 ;
        RECT 21.985 28.900 22.255 30.220 ;
        RECT 27.295 30.120 27.675 30.550 ;
        RECT 27.295 29.610 27.655 30.120 ;
        RECT 20.855 22.210 22.255 28.900 ;
        RECT 20.855 20.210 21.125 22.210 ;
        RECT 21.985 20.170 22.255 22.210 ;
        RECT 27.305 21.770 27.565 29.610 ;
        RECT 27.305 20.220 27.685 21.770 ;
        RECT 19.825 19.560 20.875 19.970 ;
        RECT 22.235 19.570 27.285 19.950 ;
        RECT 19.995 18.280 20.665 19.560 ;
        RECT 19.825 17.600 20.945 18.280 ;
        RECT 23.915 16.790 25.845 19.570 ;
        RECT 23.335 15.940 26.045 16.790 ;
        RECT 27.425 15.400 27.685 20.220 ;
        RECT 26.895 14.670 27.785 15.400 ;
        RECT 28.185 14.810 28.575 36.320 ;
        RECT 28.915 16.840 29.415 37.640 ;
        RECT 31.525 38.490 31.805 40.480 ;
        RECT 34.095 40.410 35.195 41.180 ;
        RECT 42.795 40.460 43.095 42.190 ;
        RECT 32.075 39.650 32.455 40.250 ;
        RECT 32.105 39.030 32.355 39.650 ;
        RECT 31.975 38.650 32.455 39.030 ;
        RECT 31.525 33.420 31.855 38.490 ;
        RECT 32.405 37.630 32.705 38.490 ;
        RECT 33.485 37.630 33.785 38.490 ;
        RECT 34.395 38.450 34.675 40.410 ;
        RECT 37.695 38.840 37.965 39.010 ;
        RECT 37.305 38.530 37.965 38.840 ;
        RECT 32.405 33.390 33.785 37.630 ;
        RECT 34.335 38.400 34.675 38.450 ;
        RECT 37.255 38.420 37.965 38.530 ;
        RECT 30.805 32.170 31.125 32.190 ;
        RECT 32.485 32.170 33.615 33.390 ;
        RECT 34.335 33.380 34.665 38.400 ;
        RECT 37.255 37.050 37.485 38.420 ;
        RECT 37.695 38.170 37.965 38.420 ;
        RECT 38.595 38.790 38.885 39.030 ;
        RECT 40.005 38.790 40.695 38.810 ;
        RECT 38.595 38.350 40.695 38.790 ;
        RECT 38.595 38.160 38.885 38.350 ;
        RECT 37.965 37.610 38.585 37.970 ;
        RECT 40.005 37.640 40.695 38.350 ;
        RECT 37.185 36.450 37.565 37.050 ;
        RECT 37.975 36.740 38.405 37.610 ;
        RECT 37.255 35.260 37.485 36.450 ;
        RECT 37.975 36.320 39.855 36.740 ;
        RECT 37.975 35.790 38.405 36.320 ;
        RECT 37.825 35.430 38.445 35.790 ;
        RECT 37.255 35.250 37.735 35.260 ;
        RECT 37.255 34.570 37.815 35.250 ;
        RECT 37.345 34.420 37.815 34.570 ;
        RECT 37.545 33.470 37.815 34.420 ;
        RECT 38.455 34.170 38.725 35.170 ;
        RECT 38.455 33.440 38.965 34.170 ;
        RECT 38.455 33.350 38.955 33.440 ;
        RECT 33.815 32.800 34.345 33.180 ;
        RECT 30.805 31.120 33.635 32.170 ;
        RECT 33.915 31.920 34.175 32.800 ;
        RECT 33.895 31.300 34.255 31.920 ;
        RECT 38.705 31.230 38.955 33.350 ;
        RECT 30.805 30.210 31.125 31.120 ;
        RECT 32.485 31.110 33.615 31.120 ;
        RECT 34.515 30.830 39.155 31.230 ;
        RECT 38.705 30.550 38.955 30.830 ;
        RECT 30.805 30.150 31.135 30.210 ;
        RECT 30.815 20.220 31.135 30.150 ;
        RECT 32.135 28.900 32.405 30.260 ;
        RECT 33.265 28.900 33.535 30.220 ;
        RECT 38.575 30.120 38.955 30.550 ;
        RECT 38.575 29.610 38.935 30.120 ;
        RECT 32.135 22.210 33.535 28.900 ;
        RECT 32.135 20.210 32.405 22.210 ;
        RECT 33.265 20.170 33.535 22.210 ;
        RECT 38.585 21.770 38.845 29.610 ;
        RECT 38.585 20.220 38.965 21.770 ;
        RECT 31.105 19.560 32.155 19.970 ;
        RECT 33.515 19.570 38.565 19.950 ;
        RECT 31.275 18.280 31.945 19.560 ;
        RECT 31.105 17.600 32.225 18.280 ;
        RECT 28.185 12.290 28.595 14.810 ;
        RECT 28.895 13.610 29.435 16.840 ;
        RECT 35.195 16.790 37.125 19.570 ;
        RECT 34.615 15.940 37.325 16.790 ;
        RECT 38.705 15.400 38.965 20.220 ;
        RECT 38.175 14.670 39.065 15.400 ;
        RECT 39.465 14.810 39.855 36.320 ;
        RECT 40.195 16.840 40.695 37.640 ;
        RECT 42.815 38.470 43.095 40.460 ;
        RECT 45.385 40.390 46.485 41.160 ;
        RECT 54.015 40.460 54.315 42.190 ;
        RECT 43.365 39.630 43.745 40.230 ;
        RECT 43.395 39.010 43.645 39.630 ;
        RECT 43.265 38.630 43.745 39.010 ;
        RECT 42.815 33.400 43.145 38.470 ;
        RECT 43.695 37.610 43.995 38.470 ;
        RECT 44.775 37.610 45.075 38.470 ;
        RECT 45.685 38.430 45.965 40.390 ;
        RECT 48.985 38.820 49.255 38.990 ;
        RECT 48.595 38.510 49.255 38.820 ;
        RECT 43.695 33.370 45.075 37.610 ;
        RECT 45.625 38.380 45.965 38.430 ;
        RECT 48.545 38.400 49.255 38.510 ;
        RECT 42.095 32.150 42.415 32.170 ;
        RECT 43.775 32.150 44.905 33.370 ;
        RECT 45.625 33.360 45.955 38.380 ;
        RECT 48.545 37.030 48.775 38.400 ;
        RECT 48.985 38.150 49.255 38.400 ;
        RECT 49.885 38.770 50.175 39.010 ;
        RECT 51.295 38.770 51.985 38.790 ;
        RECT 49.885 38.330 51.985 38.770 ;
        RECT 49.885 38.140 50.175 38.330 ;
        RECT 49.255 37.590 49.875 37.950 ;
        RECT 51.295 37.620 51.985 38.330 ;
        RECT 48.475 36.430 48.855 37.030 ;
        RECT 49.265 36.720 49.695 37.590 ;
        RECT 48.545 35.240 48.775 36.430 ;
        RECT 49.265 36.300 51.145 36.720 ;
        RECT 49.265 35.770 49.695 36.300 ;
        RECT 49.115 35.410 49.735 35.770 ;
        RECT 48.545 35.230 49.025 35.240 ;
        RECT 48.545 34.550 49.105 35.230 ;
        RECT 48.635 34.400 49.105 34.550 ;
        RECT 48.835 33.450 49.105 34.400 ;
        RECT 49.745 34.150 50.015 35.150 ;
        RECT 49.745 33.420 50.255 34.150 ;
        RECT 49.745 33.330 50.245 33.420 ;
        RECT 45.105 32.780 45.635 33.160 ;
        RECT 42.095 31.100 44.925 32.150 ;
        RECT 45.205 31.900 45.465 32.780 ;
        RECT 45.185 31.280 45.545 31.900 ;
        RECT 49.995 31.210 50.245 33.330 ;
        RECT 42.095 30.190 42.415 31.100 ;
        RECT 43.775 31.090 44.905 31.100 ;
        RECT 45.805 30.810 50.445 31.210 ;
        RECT 49.995 30.530 50.245 30.810 ;
        RECT 42.095 30.130 42.425 30.190 ;
        RECT 42.105 20.200 42.425 30.130 ;
        RECT 43.425 28.880 43.695 30.240 ;
        RECT 44.555 28.880 44.825 30.200 ;
        RECT 49.865 30.100 50.245 30.530 ;
        RECT 49.865 29.590 50.225 30.100 ;
        RECT 43.425 22.190 44.825 28.880 ;
        RECT 43.425 20.190 43.695 22.190 ;
        RECT 44.555 20.150 44.825 22.190 ;
        RECT 49.875 21.750 50.135 29.590 ;
        RECT 49.875 20.200 50.255 21.750 ;
        RECT 42.395 19.540 43.445 19.950 ;
        RECT 44.805 19.550 49.855 19.930 ;
        RECT 42.565 18.260 43.235 19.540 ;
        RECT 42.395 17.580 43.515 18.260 ;
        RECT 28.875 12.770 29.735 13.610 ;
        RECT 28.185 11.950 30.415 12.290 ;
        RECT 39.465 11.990 39.875 14.810 ;
        RECT 40.175 13.610 40.715 16.840 ;
        RECT 46.485 16.770 48.415 19.550 ;
        RECT 45.905 15.920 48.615 16.770 ;
        RECT 49.995 15.380 50.255 20.200 ;
        RECT 49.465 14.650 50.355 15.380 ;
        RECT 50.755 14.790 51.145 36.300 ;
        RECT 51.485 16.820 51.985 37.620 ;
        RECT 54.035 38.470 54.315 40.460 ;
        RECT 56.605 40.390 57.705 41.160 ;
        RECT 65.215 40.460 65.515 42.190 ;
        RECT 76.145 42.180 77.525 42.750 ;
        RECT 83.625 42.570 85.005 43.140 ;
        RECT 87.385 42.200 88.765 42.770 ;
        RECT 94.875 42.580 96.255 43.150 ;
        RECT 106.875 43.140 107.175 44.870 ;
        RECT 114.755 44.170 115.855 44.940 ;
        RECT 118.145 44.870 118.425 46.860 ;
        RECT 120.505 47.710 121.005 68.510 ;
        RECT 121.345 49.030 121.735 70.540 ;
        RECT 122.135 69.950 123.025 70.680 ;
        RECT 132.615 70.040 134.265 70.810 ;
        RECT 122.235 65.130 122.495 69.950 ;
        RECT 123.875 68.560 126.585 69.410 ;
        RECT 124.075 65.780 126.005 68.560 ;
        RECT 128.975 67.070 130.095 67.750 ;
        RECT 129.255 65.790 129.925 67.070 ;
        RECT 122.635 65.400 127.685 65.780 ;
        RECT 129.045 65.380 130.095 65.790 ;
        RECT 132.925 65.180 133.225 70.040 ;
        RECT 137.675 68.690 139.075 69.460 ;
        RECT 138.385 65.740 138.645 68.690 ;
        RECT 149.410 68.420 150.690 69.620 ;
        RECT 149.480 65.810 150.640 68.420 ;
        RECT 133.365 65.380 138.645 65.740 ;
        RECT 122.235 63.580 122.615 65.130 ;
        RECT 122.355 55.740 122.615 63.580 ;
        RECT 127.665 63.140 127.935 65.180 ;
        RECT 128.795 63.140 129.065 65.140 ;
        RECT 127.665 56.450 129.065 63.140 ;
        RECT 122.265 55.230 122.625 55.740 ;
        RECT 122.245 54.800 122.625 55.230 ;
        RECT 127.665 55.130 127.935 56.450 ;
        RECT 128.795 55.090 129.065 56.450 ;
        RECT 130.065 55.200 130.385 65.130 ;
        RECT 132.925 61.010 133.355 65.180 ;
        RECT 138.385 65.150 138.645 65.380 ;
        RECT 138.385 64.770 138.675 65.150 ;
        RECT 130.065 55.140 130.395 55.200 ;
        RECT 133.055 55.190 133.355 61.010 ;
        RECT 122.245 54.520 122.495 54.800 ;
        RECT 122.045 54.120 126.685 54.520 ;
        RECT 127.585 54.230 128.715 54.240 ;
        RECT 130.075 54.230 130.395 55.140 ;
        RECT 138.395 55.080 138.675 64.770 ;
        RECT 149.390 64.610 150.670 65.810 ;
        RECT 122.245 52.000 122.495 54.120 ;
        RECT 126.945 53.430 127.305 54.050 ;
        RECT 127.025 52.550 127.285 53.430 ;
        RECT 127.565 53.180 130.395 54.230 ;
        RECT 126.855 52.170 127.385 52.550 ;
        RECT 122.245 51.910 122.745 52.000 ;
        RECT 122.235 51.180 122.745 51.910 ;
        RECT 122.475 50.180 122.745 51.180 ;
        RECT 123.385 50.930 123.655 51.880 ;
        RECT 123.385 50.780 123.855 50.930 ;
        RECT 123.385 50.100 123.945 50.780 ;
        RECT 123.465 50.090 123.945 50.100 ;
        RECT 122.755 49.560 123.375 49.920 ;
        RECT 122.795 49.030 123.225 49.560 ;
        RECT 121.345 48.610 123.225 49.030 ;
        RECT 123.715 48.900 123.945 50.090 ;
        RECT 122.795 47.740 123.225 48.610 ;
        RECT 123.635 48.300 124.015 48.900 ;
        RECT 120.505 47.000 121.195 47.710 ;
        RECT 122.615 47.380 123.235 47.740 ;
        RECT 122.315 47.000 122.605 47.190 ;
        RECT 120.505 46.560 122.605 47.000 ;
        RECT 120.505 46.540 121.195 46.560 ;
        RECT 122.315 46.320 122.605 46.560 ;
        RECT 123.235 46.930 123.505 47.180 ;
        RECT 123.715 46.930 123.945 48.300 ;
        RECT 126.535 46.950 126.865 51.970 ;
        RECT 127.585 51.960 128.715 53.180 ;
        RECT 130.075 53.160 130.395 53.180 ;
        RECT 123.235 46.820 123.945 46.930 ;
        RECT 126.525 46.900 126.865 46.950 ;
        RECT 127.415 47.720 128.795 51.960 ;
        RECT 123.235 46.510 123.895 46.820 ;
        RECT 123.235 46.340 123.505 46.510 ;
        RECT 126.525 44.940 126.805 46.900 ;
        RECT 127.415 46.860 127.715 47.720 ;
        RECT 128.495 46.860 128.795 47.720 ;
        RECT 129.345 46.860 129.675 51.930 ;
        RECT 128.745 46.320 129.225 46.700 ;
        RECT 128.845 45.700 129.095 46.320 ;
        RECT 128.745 45.100 129.125 45.700 ;
        RECT 118.145 43.140 118.445 44.870 ;
        RECT 126.005 44.170 127.105 44.940 ;
        RECT 129.395 44.870 129.675 46.860 ;
        RECT 129.395 43.140 129.695 44.870 ;
        RECT 98.595 42.220 99.975 42.790 ;
        RECT 106.155 42.570 107.535 43.140 ;
        RECT 109.795 42.260 111.175 42.830 ;
        RECT 117.425 42.570 118.805 43.140 ;
        RECT 121.005 42.280 122.385 42.850 ;
        RECT 128.675 42.570 130.055 43.140 ;
        RECT 54.585 39.630 54.965 40.230 ;
        RECT 54.615 39.010 54.865 39.630 ;
        RECT 54.485 38.630 54.965 39.010 ;
        RECT 54.035 33.400 54.365 38.470 ;
        RECT 54.915 37.610 55.215 38.470 ;
        RECT 55.995 37.610 56.295 38.470 ;
        RECT 56.905 38.430 57.185 40.390 ;
        RECT 60.205 38.820 60.475 38.990 ;
        RECT 59.815 38.510 60.475 38.820 ;
        RECT 54.915 33.370 56.295 37.610 ;
        RECT 56.845 38.380 57.185 38.430 ;
        RECT 59.765 38.400 60.475 38.510 ;
        RECT 53.315 32.150 53.635 32.170 ;
        RECT 54.995 32.150 56.125 33.370 ;
        RECT 56.845 33.360 57.175 38.380 ;
        RECT 59.765 37.030 59.995 38.400 ;
        RECT 60.205 38.150 60.475 38.400 ;
        RECT 61.105 38.770 61.395 39.010 ;
        RECT 62.515 38.770 63.205 38.790 ;
        RECT 61.105 38.330 63.205 38.770 ;
        RECT 61.105 38.140 61.395 38.330 ;
        RECT 60.475 37.590 61.095 37.950 ;
        RECT 62.515 37.620 63.205 38.330 ;
        RECT 59.695 36.430 60.075 37.030 ;
        RECT 60.485 36.720 60.915 37.590 ;
        RECT 59.765 35.240 59.995 36.430 ;
        RECT 60.485 36.300 62.365 36.720 ;
        RECT 60.485 35.770 60.915 36.300 ;
        RECT 60.335 35.410 60.955 35.770 ;
        RECT 59.765 35.230 60.245 35.240 ;
        RECT 59.765 34.550 60.325 35.230 ;
        RECT 59.855 34.400 60.325 34.550 ;
        RECT 60.055 33.450 60.325 34.400 ;
        RECT 60.965 34.150 61.235 35.150 ;
        RECT 60.965 33.420 61.475 34.150 ;
        RECT 60.965 33.330 61.465 33.420 ;
        RECT 56.325 32.780 56.855 33.160 ;
        RECT 53.315 31.100 56.145 32.150 ;
        RECT 56.425 31.900 56.685 32.780 ;
        RECT 56.405 31.280 56.765 31.900 ;
        RECT 61.215 31.210 61.465 33.330 ;
        RECT 53.315 30.190 53.635 31.100 ;
        RECT 54.995 31.090 56.125 31.100 ;
        RECT 57.025 30.810 61.665 31.210 ;
        RECT 61.215 30.530 61.465 30.810 ;
        RECT 53.315 30.130 53.645 30.190 ;
        RECT 53.325 20.200 53.645 30.130 ;
        RECT 54.645 28.880 54.915 30.240 ;
        RECT 55.775 28.880 56.045 30.200 ;
        RECT 61.085 30.100 61.465 30.530 ;
        RECT 61.085 29.590 61.445 30.100 ;
        RECT 54.645 22.190 56.045 28.880 ;
        RECT 54.645 20.190 54.915 22.190 ;
        RECT 55.775 20.150 56.045 22.190 ;
        RECT 61.095 21.750 61.355 29.590 ;
        RECT 61.095 20.200 61.475 21.750 ;
        RECT 53.615 19.540 54.665 19.950 ;
        RECT 56.025 19.550 61.075 19.930 ;
        RECT 53.785 18.260 54.455 19.540 ;
        RECT 53.615 17.580 54.735 18.260 ;
        RECT 40.155 12.770 41.015 13.610 ;
        RECT 50.755 12.170 51.165 14.790 ;
        RECT 51.465 13.590 52.005 16.820 ;
        RECT 57.705 16.770 59.635 19.550 ;
        RECT 57.125 15.920 59.835 16.770 ;
        RECT 61.215 15.380 61.475 20.200 ;
        RECT 60.685 14.650 61.575 15.380 ;
        RECT 61.975 14.790 62.365 36.300 ;
        RECT 62.705 16.820 63.205 37.620 ;
        RECT 65.235 38.470 65.515 40.460 ;
        RECT 67.805 40.390 68.905 41.160 ;
        RECT 76.505 40.450 76.805 42.180 ;
        RECT 65.785 39.630 66.165 40.230 ;
        RECT 65.815 39.010 66.065 39.630 ;
        RECT 65.685 38.630 66.165 39.010 ;
        RECT 65.235 33.400 65.565 38.470 ;
        RECT 66.115 37.610 66.415 38.470 ;
        RECT 67.195 37.610 67.495 38.470 ;
        RECT 68.105 38.430 68.385 40.390 ;
        RECT 71.405 38.820 71.675 38.990 ;
        RECT 71.015 38.510 71.675 38.820 ;
        RECT 66.115 33.370 67.495 37.610 ;
        RECT 68.045 38.380 68.385 38.430 ;
        RECT 70.965 38.400 71.675 38.510 ;
        RECT 64.515 32.150 64.835 32.170 ;
        RECT 66.195 32.150 67.325 33.370 ;
        RECT 68.045 33.360 68.375 38.380 ;
        RECT 70.965 37.030 71.195 38.400 ;
        RECT 71.405 38.150 71.675 38.400 ;
        RECT 72.305 38.770 72.595 39.010 ;
        RECT 73.715 38.770 74.405 38.790 ;
        RECT 72.305 38.330 74.405 38.770 ;
        RECT 72.305 38.140 72.595 38.330 ;
        RECT 71.675 37.590 72.295 37.950 ;
        RECT 73.715 37.620 74.405 38.330 ;
        RECT 70.895 36.430 71.275 37.030 ;
        RECT 71.685 36.720 72.115 37.590 ;
        RECT 70.965 35.240 71.195 36.430 ;
        RECT 71.685 36.300 73.565 36.720 ;
        RECT 71.685 35.770 72.115 36.300 ;
        RECT 71.535 35.410 72.155 35.770 ;
        RECT 70.965 35.230 71.445 35.240 ;
        RECT 70.965 34.550 71.525 35.230 ;
        RECT 71.055 34.400 71.525 34.550 ;
        RECT 71.255 33.450 71.525 34.400 ;
        RECT 72.165 34.150 72.435 35.150 ;
        RECT 72.165 33.420 72.675 34.150 ;
        RECT 72.165 33.330 72.665 33.420 ;
        RECT 67.525 32.780 68.055 33.160 ;
        RECT 64.515 31.100 67.345 32.150 ;
        RECT 67.625 31.900 67.885 32.780 ;
        RECT 67.605 31.280 67.965 31.900 ;
        RECT 72.415 31.210 72.665 33.330 ;
        RECT 64.515 30.190 64.835 31.100 ;
        RECT 66.195 31.090 67.325 31.100 ;
        RECT 68.225 30.810 72.865 31.210 ;
        RECT 72.415 30.530 72.665 30.810 ;
        RECT 64.515 30.130 64.845 30.190 ;
        RECT 64.525 20.200 64.845 30.130 ;
        RECT 65.845 28.880 66.115 30.240 ;
        RECT 66.975 28.880 67.245 30.200 ;
        RECT 72.285 30.100 72.665 30.530 ;
        RECT 72.285 29.590 72.645 30.100 ;
        RECT 65.845 22.190 67.245 28.880 ;
        RECT 65.845 20.190 66.115 22.190 ;
        RECT 66.975 20.150 67.245 22.190 ;
        RECT 72.295 21.750 72.555 29.590 ;
        RECT 72.295 20.200 72.675 21.750 ;
        RECT 64.815 19.540 65.865 19.950 ;
        RECT 67.225 19.550 72.275 19.930 ;
        RECT 64.985 18.260 65.655 19.540 ;
        RECT 64.815 17.580 65.935 18.260 ;
        RECT 51.445 12.750 52.305 13.590 ;
        RECT 27.865 11.130 30.415 11.950 ;
        RECT 28.395 11.090 30.415 11.130 ;
        RECT 39.115 10.980 41.565 11.990 ;
        RECT 50.335 10.970 52.355 12.170 ;
        RECT 61.975 12.160 62.385 14.790 ;
        RECT 62.685 13.590 63.225 16.820 ;
        RECT 68.905 16.770 70.835 19.550 ;
        RECT 68.325 15.920 71.035 16.770 ;
        RECT 72.415 15.380 72.675 20.200 ;
        RECT 71.885 14.650 72.775 15.380 ;
        RECT 73.175 14.790 73.565 36.300 ;
        RECT 73.905 16.820 74.405 37.620 ;
        RECT 76.525 38.460 76.805 40.450 ;
        RECT 79.095 40.380 80.195 41.150 ;
        RECT 87.745 40.470 88.045 42.200 ;
        RECT 77.075 39.620 77.455 40.220 ;
        RECT 77.105 39.000 77.355 39.620 ;
        RECT 76.975 38.620 77.455 39.000 ;
        RECT 76.525 33.390 76.855 38.460 ;
        RECT 77.405 37.600 77.705 38.460 ;
        RECT 78.485 37.600 78.785 38.460 ;
        RECT 79.395 38.420 79.675 40.380 ;
        RECT 82.695 38.810 82.965 38.980 ;
        RECT 82.305 38.500 82.965 38.810 ;
        RECT 77.405 33.360 78.785 37.600 ;
        RECT 79.335 38.370 79.675 38.420 ;
        RECT 82.255 38.390 82.965 38.500 ;
        RECT 75.805 32.140 76.125 32.160 ;
        RECT 77.485 32.140 78.615 33.360 ;
        RECT 79.335 33.350 79.665 38.370 ;
        RECT 82.255 37.020 82.485 38.390 ;
        RECT 82.695 38.140 82.965 38.390 ;
        RECT 83.595 38.760 83.885 39.000 ;
        RECT 85.005 38.760 85.695 38.780 ;
        RECT 83.595 38.320 85.695 38.760 ;
        RECT 83.595 38.130 83.885 38.320 ;
        RECT 82.965 37.580 83.585 37.940 ;
        RECT 85.005 37.610 85.695 38.320 ;
        RECT 82.185 36.420 82.565 37.020 ;
        RECT 82.975 36.710 83.405 37.580 ;
        RECT 82.255 35.230 82.485 36.420 ;
        RECT 82.975 36.290 84.855 36.710 ;
        RECT 82.975 35.760 83.405 36.290 ;
        RECT 82.825 35.400 83.445 35.760 ;
        RECT 82.255 35.220 82.735 35.230 ;
        RECT 82.255 34.540 82.815 35.220 ;
        RECT 82.345 34.390 82.815 34.540 ;
        RECT 82.545 33.440 82.815 34.390 ;
        RECT 83.455 34.140 83.725 35.140 ;
        RECT 83.455 33.410 83.965 34.140 ;
        RECT 83.455 33.320 83.955 33.410 ;
        RECT 78.815 32.770 79.345 33.150 ;
        RECT 75.805 31.090 78.635 32.140 ;
        RECT 78.915 31.890 79.175 32.770 ;
        RECT 78.895 31.270 79.255 31.890 ;
        RECT 83.705 31.200 83.955 33.320 ;
        RECT 75.805 30.180 76.125 31.090 ;
        RECT 77.485 31.080 78.615 31.090 ;
        RECT 79.515 30.800 84.155 31.200 ;
        RECT 83.705 30.520 83.955 30.800 ;
        RECT 75.805 30.120 76.135 30.180 ;
        RECT 75.815 20.190 76.135 30.120 ;
        RECT 77.135 28.870 77.405 30.230 ;
        RECT 78.265 28.870 78.535 30.190 ;
        RECT 83.575 30.090 83.955 30.520 ;
        RECT 83.575 29.580 83.935 30.090 ;
        RECT 77.135 22.180 78.535 28.870 ;
        RECT 77.135 20.180 77.405 22.180 ;
        RECT 78.265 20.140 78.535 22.180 ;
        RECT 83.585 21.740 83.845 29.580 ;
        RECT 83.585 20.190 83.965 21.740 ;
        RECT 76.105 19.530 77.155 19.940 ;
        RECT 78.515 19.540 83.565 19.920 ;
        RECT 76.275 18.250 76.945 19.530 ;
        RECT 76.105 17.570 77.225 18.250 ;
        RECT 62.665 12.750 63.525 13.590 ;
        RECT 73.175 12.190 73.585 14.790 ;
        RECT 73.885 13.590 74.425 16.820 ;
        RECT 80.195 16.760 82.125 19.540 ;
        RECT 79.615 15.910 82.325 16.760 ;
        RECT 83.705 15.370 83.965 20.190 ;
        RECT 83.175 14.640 84.065 15.370 ;
        RECT 84.465 14.780 84.855 36.290 ;
        RECT 85.195 16.810 85.695 37.610 ;
        RECT 87.765 38.480 88.045 40.470 ;
        RECT 90.335 40.400 91.435 41.170 ;
        RECT 98.955 40.490 99.255 42.220 ;
        RECT 88.315 39.640 88.695 40.240 ;
        RECT 88.345 39.020 88.595 39.640 ;
        RECT 88.215 38.640 88.695 39.020 ;
        RECT 87.765 33.410 88.095 38.480 ;
        RECT 88.645 37.620 88.945 38.480 ;
        RECT 89.725 37.620 90.025 38.480 ;
        RECT 90.635 38.440 90.915 40.400 ;
        RECT 93.935 38.830 94.205 39.000 ;
        RECT 93.545 38.520 94.205 38.830 ;
        RECT 88.645 33.380 90.025 37.620 ;
        RECT 90.575 38.390 90.915 38.440 ;
        RECT 93.495 38.410 94.205 38.520 ;
        RECT 87.045 32.160 87.365 32.180 ;
        RECT 88.725 32.160 89.855 33.380 ;
        RECT 90.575 33.370 90.905 38.390 ;
        RECT 93.495 37.040 93.725 38.410 ;
        RECT 93.935 38.160 94.205 38.410 ;
        RECT 94.835 38.780 95.125 39.020 ;
        RECT 96.245 38.780 96.935 38.800 ;
        RECT 94.835 38.340 96.935 38.780 ;
        RECT 94.835 38.150 95.125 38.340 ;
        RECT 94.205 37.600 94.825 37.960 ;
        RECT 96.245 37.630 96.935 38.340 ;
        RECT 93.425 36.440 93.805 37.040 ;
        RECT 94.215 36.730 94.645 37.600 ;
        RECT 93.495 35.250 93.725 36.440 ;
        RECT 94.215 36.310 96.095 36.730 ;
        RECT 94.215 35.780 94.645 36.310 ;
        RECT 94.065 35.420 94.685 35.780 ;
        RECT 93.495 35.240 93.975 35.250 ;
        RECT 93.495 34.560 94.055 35.240 ;
        RECT 93.585 34.410 94.055 34.560 ;
        RECT 93.785 33.460 94.055 34.410 ;
        RECT 94.695 34.160 94.965 35.160 ;
        RECT 94.695 33.430 95.205 34.160 ;
        RECT 94.695 33.340 95.195 33.430 ;
        RECT 90.055 32.790 90.585 33.170 ;
        RECT 87.045 31.110 89.875 32.160 ;
        RECT 90.155 31.910 90.415 32.790 ;
        RECT 90.135 31.290 90.495 31.910 ;
        RECT 94.945 31.220 95.195 33.340 ;
        RECT 87.045 30.200 87.365 31.110 ;
        RECT 88.725 31.100 89.855 31.110 ;
        RECT 90.755 30.820 95.395 31.220 ;
        RECT 94.945 30.540 95.195 30.820 ;
        RECT 87.045 30.140 87.375 30.200 ;
        RECT 87.055 20.210 87.375 30.140 ;
        RECT 88.375 28.890 88.645 30.250 ;
        RECT 89.505 28.890 89.775 30.210 ;
        RECT 94.815 30.110 95.195 30.540 ;
        RECT 94.815 29.600 95.175 30.110 ;
        RECT 88.375 22.200 89.775 28.890 ;
        RECT 88.375 20.200 88.645 22.200 ;
        RECT 89.505 20.160 89.775 22.200 ;
        RECT 94.825 21.760 95.085 29.600 ;
        RECT 94.825 20.210 95.205 21.760 ;
        RECT 87.345 19.550 88.395 19.960 ;
        RECT 89.755 19.560 94.805 19.940 ;
        RECT 87.515 18.270 88.185 19.550 ;
        RECT 87.345 17.590 88.465 18.270 ;
        RECT 73.865 12.750 74.725 13.590 ;
        RECT 61.415 10.960 63.435 12.160 ;
        RECT 72.725 10.990 74.745 12.190 ;
        RECT 84.465 12.180 84.875 14.780 ;
        RECT 85.175 13.580 85.715 16.810 ;
        RECT 91.435 16.780 93.365 19.560 ;
        RECT 90.855 15.930 93.565 16.780 ;
        RECT 94.945 15.390 95.205 20.210 ;
        RECT 94.415 14.660 95.305 15.390 ;
        RECT 95.705 14.800 96.095 36.310 ;
        RECT 96.435 16.830 96.935 37.630 ;
        RECT 98.975 38.500 99.255 40.490 ;
        RECT 101.545 40.420 102.645 41.190 ;
        RECT 110.155 40.530 110.455 42.260 ;
        RECT 99.525 39.660 99.905 40.260 ;
        RECT 99.555 39.040 99.805 39.660 ;
        RECT 99.425 38.660 99.905 39.040 ;
        RECT 98.975 33.430 99.305 38.500 ;
        RECT 99.855 37.640 100.155 38.500 ;
        RECT 100.935 37.640 101.235 38.500 ;
        RECT 101.845 38.460 102.125 40.420 ;
        RECT 105.145 38.850 105.415 39.020 ;
        RECT 104.755 38.540 105.415 38.850 ;
        RECT 99.855 33.400 101.235 37.640 ;
        RECT 101.785 38.410 102.125 38.460 ;
        RECT 104.705 38.430 105.415 38.540 ;
        RECT 98.255 32.180 98.575 32.200 ;
        RECT 99.935 32.180 101.065 33.400 ;
        RECT 101.785 33.390 102.115 38.410 ;
        RECT 104.705 37.060 104.935 38.430 ;
        RECT 105.145 38.180 105.415 38.430 ;
        RECT 106.045 38.800 106.335 39.040 ;
        RECT 107.455 38.800 108.145 38.820 ;
        RECT 106.045 38.360 108.145 38.800 ;
        RECT 106.045 38.170 106.335 38.360 ;
        RECT 105.415 37.620 106.035 37.980 ;
        RECT 107.455 37.650 108.145 38.360 ;
        RECT 104.635 36.460 105.015 37.060 ;
        RECT 105.425 36.750 105.855 37.620 ;
        RECT 104.705 35.270 104.935 36.460 ;
        RECT 105.425 36.330 107.305 36.750 ;
        RECT 105.425 35.800 105.855 36.330 ;
        RECT 105.275 35.440 105.895 35.800 ;
        RECT 104.705 35.260 105.185 35.270 ;
        RECT 104.705 34.580 105.265 35.260 ;
        RECT 104.795 34.430 105.265 34.580 ;
        RECT 104.995 33.480 105.265 34.430 ;
        RECT 105.905 34.180 106.175 35.180 ;
        RECT 105.905 33.450 106.415 34.180 ;
        RECT 105.905 33.360 106.405 33.450 ;
        RECT 101.265 32.810 101.795 33.190 ;
        RECT 98.255 31.130 101.085 32.180 ;
        RECT 101.365 31.930 101.625 32.810 ;
        RECT 101.345 31.310 101.705 31.930 ;
        RECT 106.155 31.240 106.405 33.360 ;
        RECT 98.255 30.220 98.575 31.130 ;
        RECT 99.935 31.120 101.065 31.130 ;
        RECT 101.965 30.840 106.605 31.240 ;
        RECT 106.155 30.560 106.405 30.840 ;
        RECT 98.255 30.160 98.585 30.220 ;
        RECT 98.265 20.230 98.585 30.160 ;
        RECT 99.585 28.910 99.855 30.270 ;
        RECT 100.715 28.910 100.985 30.230 ;
        RECT 106.025 30.130 106.405 30.560 ;
        RECT 106.025 29.620 106.385 30.130 ;
        RECT 99.585 22.220 100.985 28.910 ;
        RECT 99.585 20.220 99.855 22.220 ;
        RECT 100.715 20.180 100.985 22.220 ;
        RECT 106.035 21.780 106.295 29.620 ;
        RECT 106.035 20.230 106.415 21.780 ;
        RECT 98.555 19.570 99.605 19.980 ;
        RECT 100.965 19.580 106.015 19.960 ;
        RECT 98.725 18.290 99.395 19.570 ;
        RECT 98.555 17.610 99.675 18.290 ;
        RECT 85.155 12.740 86.015 13.580 ;
        RECT 95.705 12.180 96.115 14.800 ;
        RECT 96.415 13.600 96.955 16.830 ;
        RECT 102.645 16.800 104.575 19.580 ;
        RECT 102.065 15.950 104.775 16.800 ;
        RECT 106.155 15.410 106.415 20.230 ;
        RECT 105.625 14.680 106.515 15.410 ;
        RECT 106.915 14.820 107.305 36.330 ;
        RECT 107.645 16.850 108.145 37.650 ;
        RECT 110.175 38.540 110.455 40.530 ;
        RECT 112.745 40.460 113.845 41.230 ;
        RECT 121.365 40.550 121.665 42.280 ;
        RECT 142.880 42.020 144.100 43.390 ;
        RECT 110.725 39.700 111.105 40.300 ;
        RECT 110.755 39.080 111.005 39.700 ;
        RECT 110.625 38.700 111.105 39.080 ;
        RECT 110.175 33.470 110.505 38.540 ;
        RECT 111.055 37.680 111.355 38.540 ;
        RECT 112.135 37.680 112.435 38.540 ;
        RECT 113.045 38.500 113.325 40.460 ;
        RECT 116.345 38.890 116.615 39.060 ;
        RECT 115.955 38.580 116.615 38.890 ;
        RECT 111.055 33.440 112.435 37.680 ;
        RECT 112.985 38.450 113.325 38.500 ;
        RECT 115.905 38.470 116.615 38.580 ;
        RECT 109.455 32.220 109.775 32.240 ;
        RECT 111.135 32.220 112.265 33.440 ;
        RECT 112.985 33.430 113.315 38.450 ;
        RECT 115.905 37.100 116.135 38.470 ;
        RECT 116.345 38.220 116.615 38.470 ;
        RECT 117.245 38.840 117.535 39.080 ;
        RECT 118.655 38.840 119.345 38.860 ;
        RECT 117.245 38.400 119.345 38.840 ;
        RECT 117.245 38.210 117.535 38.400 ;
        RECT 116.615 37.660 117.235 38.020 ;
        RECT 118.655 37.690 119.345 38.400 ;
        RECT 115.835 36.500 116.215 37.100 ;
        RECT 116.625 36.790 117.055 37.660 ;
        RECT 115.905 35.310 116.135 36.500 ;
        RECT 116.625 36.370 118.505 36.790 ;
        RECT 116.625 35.840 117.055 36.370 ;
        RECT 116.475 35.480 117.095 35.840 ;
        RECT 115.905 35.300 116.385 35.310 ;
        RECT 115.905 34.620 116.465 35.300 ;
        RECT 115.995 34.470 116.465 34.620 ;
        RECT 116.195 33.520 116.465 34.470 ;
        RECT 117.105 34.220 117.375 35.220 ;
        RECT 117.105 33.490 117.615 34.220 ;
        RECT 117.105 33.400 117.605 33.490 ;
        RECT 112.465 32.850 112.995 33.230 ;
        RECT 109.455 31.170 112.285 32.220 ;
        RECT 112.565 31.970 112.825 32.850 ;
        RECT 112.545 31.350 112.905 31.970 ;
        RECT 117.355 31.280 117.605 33.400 ;
        RECT 109.455 30.260 109.775 31.170 ;
        RECT 111.135 31.160 112.265 31.170 ;
        RECT 113.165 30.880 117.805 31.280 ;
        RECT 117.355 30.600 117.605 30.880 ;
        RECT 109.455 30.200 109.785 30.260 ;
        RECT 109.465 20.270 109.785 30.200 ;
        RECT 110.785 28.950 111.055 30.310 ;
        RECT 111.915 28.950 112.185 30.270 ;
        RECT 117.225 30.170 117.605 30.600 ;
        RECT 117.225 29.660 117.585 30.170 ;
        RECT 110.785 22.260 112.185 28.950 ;
        RECT 110.785 20.260 111.055 22.260 ;
        RECT 111.915 20.220 112.185 22.260 ;
        RECT 117.235 21.820 117.495 29.660 ;
        RECT 117.235 20.270 117.615 21.820 ;
        RECT 109.755 19.610 110.805 20.020 ;
        RECT 112.165 19.620 117.215 20.000 ;
        RECT 109.925 18.330 110.595 19.610 ;
        RECT 109.755 17.650 110.875 18.330 ;
        RECT 96.395 12.760 97.255 13.600 ;
        RECT 106.915 12.230 107.325 14.820 ;
        RECT 107.625 13.620 108.165 16.850 ;
        RECT 113.845 16.840 115.775 19.620 ;
        RECT 113.265 15.990 115.975 16.840 ;
        RECT 117.355 15.450 117.615 20.270 ;
        RECT 116.825 14.720 117.715 15.450 ;
        RECT 118.115 14.860 118.505 36.370 ;
        RECT 118.845 16.890 119.345 37.690 ;
        RECT 121.385 38.560 121.665 40.550 ;
        RECT 123.955 40.480 125.055 41.250 ;
        RECT 121.935 39.720 122.315 40.320 ;
        RECT 121.965 39.100 122.215 39.720 ;
        RECT 121.835 38.720 122.315 39.100 ;
        RECT 121.385 33.490 121.715 38.560 ;
        RECT 122.265 37.700 122.565 38.560 ;
        RECT 123.345 37.700 123.645 38.560 ;
        RECT 124.255 38.520 124.535 40.480 ;
        RECT 127.555 38.910 127.825 39.080 ;
        RECT 127.165 38.600 127.825 38.910 ;
        RECT 122.265 33.460 123.645 37.700 ;
        RECT 124.195 38.470 124.535 38.520 ;
        RECT 127.115 38.490 127.825 38.600 ;
        RECT 120.665 32.240 120.985 32.260 ;
        RECT 122.345 32.240 123.475 33.460 ;
        RECT 124.195 33.450 124.525 38.470 ;
        RECT 127.115 37.120 127.345 38.490 ;
        RECT 127.555 38.240 127.825 38.490 ;
        RECT 128.455 38.860 128.745 39.100 ;
        RECT 142.940 38.950 144.100 42.020 ;
        RECT 129.865 38.860 130.555 38.880 ;
        RECT 128.455 38.420 130.555 38.860 ;
        RECT 128.455 38.230 128.745 38.420 ;
        RECT 127.825 37.680 128.445 38.040 ;
        RECT 129.865 37.710 130.555 38.420 ;
        RECT 127.045 36.520 127.425 37.120 ;
        RECT 127.835 36.810 128.265 37.680 ;
        RECT 127.115 35.330 127.345 36.520 ;
        RECT 127.835 36.390 129.715 36.810 ;
        RECT 127.835 35.860 128.265 36.390 ;
        RECT 127.685 35.500 128.305 35.860 ;
        RECT 127.115 35.320 127.595 35.330 ;
        RECT 127.115 34.640 127.675 35.320 ;
        RECT 127.205 34.490 127.675 34.640 ;
        RECT 127.405 33.540 127.675 34.490 ;
        RECT 128.315 34.240 128.585 35.240 ;
        RECT 128.315 33.510 128.825 34.240 ;
        RECT 128.315 33.420 128.815 33.510 ;
        RECT 123.675 32.870 124.205 33.250 ;
        RECT 120.665 31.190 123.495 32.240 ;
        RECT 123.775 31.990 124.035 32.870 ;
        RECT 123.755 31.370 124.115 31.990 ;
        RECT 128.565 31.300 128.815 33.420 ;
        RECT 120.665 30.280 120.985 31.190 ;
        RECT 122.345 31.180 123.475 31.190 ;
        RECT 124.375 30.900 129.015 31.300 ;
        RECT 128.565 30.620 128.815 30.900 ;
        RECT 120.665 30.220 120.995 30.280 ;
        RECT 120.675 20.290 120.995 30.220 ;
        RECT 121.995 28.970 122.265 30.330 ;
        RECT 123.125 28.970 123.395 30.290 ;
        RECT 128.435 30.190 128.815 30.620 ;
        RECT 128.435 29.680 128.795 30.190 ;
        RECT 121.995 22.280 123.395 28.970 ;
        RECT 121.995 20.280 122.265 22.280 ;
        RECT 123.125 20.240 123.395 22.280 ;
        RECT 128.445 21.840 128.705 29.680 ;
        RECT 128.445 20.290 128.825 21.840 ;
        RECT 120.965 19.630 122.015 20.040 ;
        RECT 123.375 19.640 128.425 20.020 ;
        RECT 121.135 18.350 121.805 19.630 ;
        RECT 120.965 17.670 122.085 18.350 ;
        RECT 107.605 12.780 108.465 13.620 ;
        RECT 118.115 12.230 118.525 14.860 ;
        RECT 118.825 13.660 119.365 16.890 ;
        RECT 125.055 16.860 126.985 19.640 ;
        RECT 124.475 16.010 127.185 16.860 ;
        RECT 128.565 15.470 128.825 20.290 ;
        RECT 128.035 14.740 128.925 15.470 ;
        RECT 129.325 14.880 129.715 36.390 ;
        RECT 130.055 16.910 130.555 37.710 ;
        RECT 142.900 37.580 144.120 38.950 ;
        RECT 132.395 24.340 132.705 30.230 ;
        RECT 132.195 20.120 132.705 24.340 ;
        RECT 118.805 12.820 119.665 13.660 ;
        RECT 129.325 12.260 129.735 14.880 ;
        RECT 130.035 13.680 130.575 16.910 ;
        RECT 132.195 15.510 132.505 20.120 ;
        RECT 137.715 19.980 138.005 30.170 ;
        RECT 132.685 19.590 138.005 19.980 ;
        RECT 137.715 16.940 138.005 19.590 ;
        RECT 142.940 17.940 144.090 19.160 ;
        RECT 145.080 18.760 146.200 18.930 ;
        RECT 137.395 15.890 138.295 16.940 ;
        RECT 137.715 15.720 138.005 15.890 ;
        RECT 131.975 14.270 132.735 15.510 ;
        RECT 142.940 15.090 144.050 17.940 ;
        RECT 142.900 13.870 144.050 15.090 ;
        RECT 145.070 14.920 146.200 18.760 ;
        RECT 145.030 13.970 146.200 14.920 ;
        RECT 145.030 13.900 146.150 13.970 ;
        RECT 130.015 12.840 130.875 13.680 ;
        RECT 83.845 10.980 85.865 12.180 ;
        RECT 95.145 10.980 97.165 12.180 ;
        RECT 106.335 11.030 108.355 12.230 ;
        RECT 117.565 11.030 119.585 12.230 ;
        RECT 128.865 11.060 130.885 12.260 ;
        RECT 74.340 0.110 75.630 1.460 ;
        RECT 93.550 0.180 94.840 1.530 ;
        RECT 112.950 0.310 114.240 1.660 ;
        RECT 131.850 0.380 133.490 1.930 ;
        RECT 151.650 0.250 152.920 1.470 ;
      LAYER met3 ;
        RECT 135.340 223.855 136.790 225.205 ;
        RECT 138.130 223.785 139.580 225.135 ;
        RECT 143.180 223.815 144.630 225.165 ;
        RECT 46.830 211.125 48.810 211.455 ;
        RECT 76.830 211.125 78.810 211.455 ;
        RECT 106.830 211.125 108.810 211.455 ;
        RECT 31.830 208.405 33.810 208.735 ;
        RECT 61.830 208.405 63.810 208.735 ;
        RECT 91.830 208.405 93.810 208.735 ;
        RECT 121.830 208.405 123.810 208.735 ;
        RECT 46.830 205.685 48.810 206.015 ;
        RECT 76.830 205.685 78.810 206.015 ;
        RECT 106.830 205.685 108.810 206.015 ;
        RECT 31.830 202.965 33.810 203.295 ;
        RECT 61.830 202.965 63.810 203.295 ;
        RECT 91.830 202.965 93.810 203.295 ;
        RECT 121.830 202.965 123.810 203.295 ;
        RECT 46.830 200.245 48.810 200.575 ;
        RECT 76.830 200.245 78.810 200.575 ;
        RECT 106.830 200.245 108.810 200.575 ;
        RECT 31.830 197.525 33.810 197.855 ;
        RECT 61.830 197.525 63.810 197.855 ;
        RECT 91.830 197.525 93.810 197.855 ;
        RECT 121.830 197.525 123.810 197.855 ;
        RECT 46.830 194.805 48.810 195.135 ;
        RECT 76.830 194.805 78.810 195.135 ;
        RECT 106.830 194.805 108.810 195.135 ;
        RECT 31.830 192.085 33.810 192.415 ;
        RECT 61.830 192.085 63.810 192.415 ;
        RECT 91.830 192.085 93.810 192.415 ;
        RECT 121.830 192.085 123.810 192.415 ;
        RECT 46.830 189.365 48.810 189.695 ;
        RECT 76.830 189.365 78.810 189.695 ;
        RECT 106.830 189.365 108.810 189.695 ;
        RECT 31.830 186.645 33.810 186.975 ;
        RECT 61.830 186.645 63.810 186.975 ;
        RECT 91.830 186.645 93.810 186.975 ;
        RECT 121.830 186.645 123.810 186.975 ;
        RECT 46.830 183.925 48.810 184.255 ;
        RECT 76.830 183.925 78.810 184.255 ;
        RECT 106.830 183.925 108.810 184.255 ;
        RECT 31.830 181.205 33.810 181.535 ;
        RECT 61.830 181.205 63.810 181.535 ;
        RECT 91.830 181.205 93.810 181.535 ;
        RECT 121.830 181.205 123.810 181.535 ;
        RECT 109.485 179.150 109.815 179.155 ;
        RECT 109.485 179.140 110.070 179.150 ;
        RECT 109.260 178.840 110.070 179.140 ;
        RECT 109.485 178.830 110.070 178.840 ;
        RECT 109.485 178.825 109.815 178.830 ;
        RECT 46.830 178.485 48.810 178.815 ;
        RECT 76.830 178.485 78.810 178.815 ;
        RECT 106.830 178.485 108.810 178.815 ;
        RECT 48.305 177.780 48.635 177.795 ;
        RECT 51.985 177.780 52.315 177.795 ;
        RECT 48.305 177.480 52.315 177.780 ;
        RECT 48.305 177.465 48.635 177.480 ;
        RECT 51.985 177.465 52.315 177.480 ;
        RECT 108.565 177.780 108.895 177.795 ;
        RECT 110.405 177.780 110.735 177.795 ;
        RECT 108.565 177.480 110.735 177.780 ;
        RECT 108.565 177.465 108.895 177.480 ;
        RECT 110.405 177.465 110.735 177.480 ;
        RECT 66.245 177.100 66.575 177.115 ;
        RECT 80.965 177.100 81.295 177.115 ;
        RECT 66.245 176.800 81.295 177.100 ;
        RECT 66.245 176.785 66.575 176.800 ;
        RECT 80.965 176.785 81.295 176.800 ;
        RECT 31.830 175.765 33.810 176.095 ;
        RECT 61.830 175.765 63.810 176.095 ;
        RECT 91.830 175.765 93.810 176.095 ;
        RECT 121.830 175.765 123.810 176.095 ;
        RECT 68.545 175.740 68.875 175.755 ;
        RECT 83.725 175.740 84.055 175.755 ;
        RECT 68.545 175.440 84.055 175.740 ;
        RECT 68.545 175.425 68.875 175.440 ;
        RECT 83.725 175.425 84.055 175.440 ;
        RECT 51.525 175.060 51.855 175.075 ;
        RECT 55.205 175.060 55.535 175.075 ;
        RECT 51.525 174.760 55.535 175.060 ;
        RECT 51.525 174.745 51.855 174.760 ;
        RECT 55.205 174.745 55.535 174.760 ;
        RECT 56.585 175.060 56.915 175.075 ;
        RECT 60.265 175.060 60.595 175.075 ;
        RECT 75.905 175.060 76.235 175.075 ;
        RECT 56.585 174.760 76.235 175.060 ;
        RECT 56.585 174.745 56.915 174.760 ;
        RECT 60.265 174.745 60.595 174.760 ;
        RECT 75.905 174.745 76.235 174.760 ;
        RECT 81.170 174.380 81.550 174.390 ;
        RECT 81.885 174.380 82.215 174.395 ;
        RECT 81.170 174.080 82.215 174.380 ;
        RECT 81.170 174.070 81.550 174.080 ;
        RECT 81.885 174.065 82.215 174.080 ;
        RECT 122.825 174.380 123.155 174.395 ;
        RECT 131.340 174.380 133.340 174.530 ;
        RECT 122.825 174.080 133.340 174.380 ;
        RECT 122.825 174.065 123.155 174.080 ;
        RECT 131.340 173.930 133.340 174.080 ;
        RECT 46.830 173.045 48.810 173.375 ;
        RECT 76.830 173.045 78.810 173.375 ;
        RECT 106.830 173.045 108.810 173.375 ;
        RECT 47.385 172.340 47.715 172.355 ;
        RECT 64.610 172.340 64.990 172.350 ;
        RECT 96.605 172.340 96.935 172.355 ;
        RECT 98.905 172.340 99.235 172.355 ;
        RECT 47.385 172.040 99.235 172.340 ;
        RECT 47.385 172.025 47.715 172.040 ;
        RECT 64.610 172.030 64.990 172.040 ;
        RECT 96.605 172.025 96.935 172.040 ;
        RECT 98.905 172.025 99.235 172.040 ;
        RECT 72.225 170.980 72.555 170.995 ;
        RECT 72.890 170.980 73.270 170.990 ;
        RECT 72.225 170.680 73.270 170.980 ;
        RECT 72.225 170.665 72.555 170.680 ;
        RECT 72.890 170.670 73.270 170.680 ;
        RECT 31.830 170.325 33.810 170.655 ;
        RECT 61.830 170.325 63.810 170.655 ;
        RECT 91.830 170.325 93.810 170.655 ;
        RECT 121.830 170.325 123.810 170.655 ;
        RECT 129.240 170.585 133.810 172.125 ;
        RECT 33.585 169.620 33.915 169.635 ;
        RECT 47.385 169.620 47.715 169.635 ;
        RECT 33.585 169.320 47.715 169.620 ;
        RECT 33.585 169.305 33.915 169.320 ;
        RECT 47.385 169.305 47.715 169.320 ;
        RECT 46.830 167.605 48.810 167.935 ;
        RECT 76.830 167.605 78.810 167.935 ;
        RECT 106.830 167.605 108.810 167.935 ;
        RECT 31.830 164.885 33.810 165.215 ;
        RECT 61.830 164.885 63.810 165.215 ;
        RECT 91.830 164.885 93.810 165.215 ;
        RECT 121.830 164.885 123.810 165.215 ;
        RECT 46.830 162.165 48.810 162.495 ;
        RECT 76.830 162.165 78.810 162.495 ;
        RECT 106.830 162.165 108.810 162.495 ;
        RECT 39.565 161.460 39.895 161.475 ;
        RECT 46.925 161.460 47.255 161.475 ;
        RECT 39.565 161.160 47.255 161.460 ;
        RECT 39.565 161.145 39.895 161.160 ;
        RECT 46.925 161.145 47.255 161.160 ;
        RECT 70.385 161.460 70.715 161.475 ;
        RECT 74.065 161.460 74.395 161.475 ;
        RECT 70.385 161.160 74.395 161.460 ;
        RECT 70.385 161.145 70.715 161.160 ;
        RECT 74.065 161.145 74.395 161.160 ;
        RECT 39.105 160.780 39.435 160.795 ;
        RECT 47.385 160.780 47.715 160.795 ;
        RECT 39.105 160.480 47.715 160.780 ;
        RECT 39.105 160.465 39.435 160.480 ;
        RECT 47.385 160.465 47.715 160.480 ;
        RECT 31.830 159.445 33.810 159.775 ;
        RECT 61.830 159.445 63.810 159.775 ;
        RECT 91.830 159.445 93.810 159.775 ;
        RECT 121.830 159.445 123.810 159.775 ;
        RECT 46.830 156.725 48.810 157.055 ;
        RECT 76.830 156.725 78.810 157.055 ;
        RECT 106.830 156.725 108.810 157.055 ;
        RECT 107.645 156.020 107.975 156.035 ;
        RECT 116.385 156.020 116.715 156.035 ;
        RECT 107.645 155.720 116.715 156.020 ;
        RECT 107.645 155.705 107.975 155.720 ;
        RECT 116.385 155.705 116.715 155.720 ;
        RECT 31.830 154.005 33.810 154.335 ;
        RECT 61.830 154.005 63.810 154.335 ;
        RECT 91.830 154.005 93.810 154.335 ;
        RECT 121.830 154.005 123.810 154.335 ;
        RECT 64.610 153.300 64.990 153.310 ;
        RECT 65.325 153.300 65.655 153.315 ;
        RECT 64.610 153.000 65.655 153.300 ;
        RECT 64.610 152.990 64.990 153.000 ;
        RECT 65.325 152.985 65.655 153.000 ;
        RECT 103.045 153.300 103.375 153.315 ;
        RECT 115.925 153.300 116.255 153.315 ;
        RECT 103.045 153.000 116.255 153.300 ;
        RECT 103.045 152.985 103.375 153.000 ;
        RECT 115.925 152.985 116.255 153.000 ;
        RECT 43.705 152.620 44.035 152.635 ;
        RECT 71.305 152.620 71.635 152.635 ;
        RECT 43.705 152.320 71.635 152.620 ;
        RECT 43.705 152.305 44.035 152.320 ;
        RECT 71.305 152.305 71.635 152.320 ;
        RECT 101.205 152.620 101.535 152.635 ;
        RECT 106.725 152.620 107.055 152.635 ;
        RECT 101.205 152.320 107.055 152.620 ;
        RECT 101.205 152.305 101.535 152.320 ;
        RECT 106.725 152.305 107.055 152.320 ;
        RECT 108.565 152.620 108.895 152.635 ;
        RECT 112.705 152.620 113.035 152.635 ;
        RECT 108.565 152.320 113.035 152.620 ;
        RECT 108.565 152.305 108.895 152.320 ;
        RECT 112.705 152.305 113.035 152.320 ;
        RECT 46.830 151.285 48.810 151.615 ;
        RECT 76.830 151.285 78.810 151.615 ;
        RECT 106.830 151.285 108.810 151.615 ;
        RECT 42.785 150.580 43.115 150.595 ;
        RECT 46.465 150.580 46.795 150.595 ;
        RECT 42.785 150.280 46.795 150.580 ;
        RECT 42.785 150.265 43.115 150.280 ;
        RECT 46.465 150.265 46.795 150.280 ;
        RECT 44.165 149.900 44.495 149.915 ;
        RECT 71.765 149.900 72.095 149.915 ;
        RECT 44.165 149.600 72.095 149.900 ;
        RECT 44.165 149.585 44.495 149.600 ;
        RECT 71.765 149.585 72.095 149.600 ;
        RECT 109.945 149.220 110.275 149.235 ;
        RECT 113.165 149.220 113.495 149.235 ;
        RECT 109.945 148.920 113.495 149.220 ;
        RECT 109.945 148.905 110.275 148.920 ;
        RECT 113.165 148.905 113.495 148.920 ;
        RECT 31.830 148.565 33.810 148.895 ;
        RECT 61.830 148.565 63.810 148.895 ;
        RECT 91.830 148.565 93.810 148.895 ;
        RECT 121.830 148.565 123.810 148.895 ;
        RECT 74.065 147.180 74.395 147.195 ;
        RECT 74.065 146.880 119.690 147.180 ;
        RECT 74.065 146.865 74.395 146.880 ;
        RECT 46.830 145.845 48.810 146.175 ;
        RECT 76.830 145.845 78.810 146.175 ;
        RECT 106.830 145.845 108.810 146.175 ;
        RECT 81.425 145.830 81.755 145.835 ;
        RECT 81.170 145.820 81.755 145.830 ;
        RECT 80.970 145.520 81.755 145.820 ;
        RECT 81.170 145.510 81.755 145.520 ;
        RECT 81.425 145.505 81.755 145.510 ;
        RECT 119.390 144.460 119.690 146.880 ;
        RECT 119.390 144.160 124.750 144.460 ;
        RECT 31.830 143.125 33.810 143.455 ;
        RECT 61.830 143.125 63.810 143.455 ;
        RECT 91.830 143.125 93.810 143.455 ;
        RECT 121.830 143.125 123.810 143.455 ;
        RECT 124.450 143.100 124.750 144.160 ;
        RECT 131.340 143.100 133.340 143.250 ;
        RECT 124.450 142.800 133.340 143.100 ;
        RECT 131.340 142.650 133.340 142.800 ;
        RECT 86.485 141.740 86.815 141.755 ;
        RECT 100.285 141.740 100.615 141.755 ;
        RECT 110.405 141.740 110.735 141.755 ;
        RECT 86.485 141.440 110.735 141.740 ;
        RECT 86.485 141.425 86.815 141.440 ;
        RECT 100.285 141.425 100.615 141.440 ;
        RECT 110.405 141.425 110.735 141.440 ;
        RECT 46.830 140.405 48.810 140.735 ;
        RECT 76.830 140.405 78.810 140.735 ;
        RECT 106.830 140.405 108.810 140.735 ;
        RECT 108.565 139.020 108.895 139.035 ;
        RECT 109.690 139.020 110.070 139.030 ;
        RECT 108.565 138.720 110.070 139.020 ;
        RECT 108.565 138.705 108.895 138.720 ;
        RECT 109.690 138.710 110.070 138.720 ;
        RECT 129.090 138.200 134.150 139.430 ;
        RECT 31.830 137.685 33.810 138.015 ;
        RECT 61.830 137.685 63.810 138.015 ;
        RECT 91.830 137.685 93.810 138.015 ;
        RECT 121.830 137.685 123.810 138.015 ;
        RECT 72.890 136.980 73.270 136.990 ;
        RECT 73.605 136.980 73.935 136.995 ;
        RECT 72.890 136.680 73.935 136.980 ;
        RECT 72.890 136.670 73.270 136.680 ;
        RECT 73.605 136.665 73.935 136.680 ;
        RECT 43.245 136.300 43.575 136.315 ;
        RECT 64.610 136.300 64.990 136.310 ;
        RECT 43.245 136.000 64.990 136.300 ;
        RECT 43.245 135.985 43.575 136.000 ;
        RECT 64.610 135.990 64.990 136.000 ;
        RECT 46.830 134.965 48.810 135.295 ;
        RECT 76.830 134.965 78.810 135.295 ;
        RECT 106.830 134.965 108.810 135.295 ;
        RECT 31.830 132.245 33.810 132.575 ;
        RECT 61.830 132.245 63.810 132.575 ;
        RECT 91.830 132.245 93.810 132.575 ;
        RECT 121.830 132.245 123.810 132.575 ;
        RECT 46.830 129.525 48.810 129.855 ;
        RECT 76.830 129.525 78.810 129.855 ;
        RECT 106.830 129.525 108.810 129.855 ;
        RECT 79.585 128.820 79.915 128.835 ;
        RECT 98.905 128.820 99.235 128.835 ;
        RECT 79.585 128.520 99.235 128.820 ;
        RECT 79.585 128.505 79.915 128.520 ;
        RECT 98.905 128.505 99.235 128.520 ;
        RECT 31.830 126.805 33.810 127.135 ;
        RECT 61.830 126.805 63.810 127.135 ;
        RECT 91.830 126.805 93.810 127.135 ;
        RECT 121.830 126.805 123.810 127.135 ;
        RECT 46.830 124.085 48.810 124.415 ;
        RECT 76.830 124.085 78.810 124.415 ;
        RECT 106.830 124.085 108.810 124.415 ;
        RECT 31.830 121.365 33.810 121.695 ;
        RECT 61.830 121.365 63.810 121.695 ;
        RECT 91.830 121.365 93.810 121.695 ;
        RECT 121.830 121.365 123.810 121.695 ;
        RECT 46.830 118.645 48.810 118.975 ;
        RECT 76.830 118.645 78.810 118.975 ;
        RECT 106.830 118.645 108.810 118.975 ;
        RECT 31.830 115.925 33.810 116.255 ;
        RECT 61.830 115.925 63.810 116.255 ;
        RECT 91.830 115.925 93.810 116.255 ;
        RECT 121.830 115.925 123.810 116.255 ;
        RECT 46.830 113.205 48.810 113.535 ;
        RECT 76.830 113.205 78.810 113.535 ;
        RECT 106.830 113.205 108.810 113.535 ;
        RECT 131.340 111.835 133.340 111.970 ;
        RECT 131.105 111.505 133.340 111.835 ;
        RECT 131.340 111.370 133.340 111.505 ;
        RECT 31.830 110.485 33.810 110.815 ;
        RECT 61.830 110.485 63.810 110.815 ;
        RECT 91.830 110.485 93.810 110.815 ;
        RECT 121.830 110.485 123.810 110.815 ;
        RECT 46.830 107.765 48.810 108.095 ;
        RECT 76.830 107.765 78.810 108.095 ;
        RECT 106.830 107.765 108.810 108.095 ;
        RECT 129.700 105.605 133.210 106.625 ;
        RECT 31.830 105.045 33.810 105.375 ;
        RECT 61.830 105.045 63.810 105.375 ;
        RECT 91.830 105.045 93.810 105.375 ;
        RECT 121.830 105.045 123.810 105.375 ;
        RECT 37.630 88.620 38.970 88.755 ;
        RECT 13.950 87.980 14.980 88.515 ;
        RECT 13.950 87.500 14.990 87.980 ;
        RECT 13.950 87.175 14.980 87.500 ;
        RECT 14.070 86.570 14.810 87.175 ;
        RECT 20.050 87.105 20.920 88.515 ;
        RECT 14.070 75.715 14.700 86.570 ;
        RECT 20.170 77.115 20.800 87.105 ;
        RECT 25.910 87.055 26.860 88.515 ;
        RECT 26.070 78.385 26.700 87.055 ;
        RECT 31.730 86.965 32.910 88.585 ;
        RECT 32.005 79.615 32.635 86.965 ;
        RECT 37.630 86.835 39.120 88.620 ;
        RECT 38.060 81.125 38.690 86.835 ;
        RECT 43.790 86.745 45.190 88.605 ;
        RECT 49.710 86.945 51.060 88.615 ;
        RECT 44.175 82.625 44.805 86.745 ;
        RECT 50.070 83.875 50.700 86.945 ;
        RECT 55.530 86.785 56.750 88.545 ;
        RECT 55.825 85.115 56.455 86.785 ;
        RECT 61.670 86.625 63.180 88.615 ;
        RECT 67.680 88.305 68.720 89.815 ;
        RECT 67.885 87.225 68.515 88.305 ;
        RECT 62.110 86.175 62.740 86.625 ;
        RECT 67.885 86.595 130.605 87.225 ;
        RECT 62.110 85.545 118.855 86.175 ;
        RECT 55.825 84.485 107.605 85.115 ;
        RECT 50.070 83.245 96.285 83.875 ;
        RECT 44.175 81.995 85.055 82.625 ;
        RECT 38.060 80.495 73.765 81.125 ;
        RECT 32.005 78.985 62.635 79.615 ;
        RECT 26.070 77.755 51.245 78.385 ;
        RECT 20.170 76.485 40.645 77.115 ;
        RECT 14.070 75.660 29.295 75.715 ;
        RECT 40.015 75.710 40.645 76.485 ;
        RECT 14.070 75.085 30.410 75.660 ;
        RECT 27.850 74.670 30.410 75.085 ;
        RECT 3.910 71.345 6.100 73.215 ;
        RECT 27.850 73.120 30.450 74.670 ;
        RECT 39.060 74.510 41.620 75.710 ;
        RECT 50.615 75.580 51.245 77.755 ;
        RECT 62.005 75.690 62.635 78.985 ;
        RECT 49.930 74.650 52.490 75.580 ;
        RECT 0.970 70.330 3.070 70.430 ;
        RECT 15.510 70.330 17.040 71.185 ;
        RECT 0.960 68.750 17.040 70.330 ;
        RECT 0.970 68.710 3.070 68.750 ;
        RECT 15.510 68.635 17.040 68.750 ;
        RECT 20.145 54.060 20.605 54.135 ;
        RECT 25.715 54.060 26.175 54.085 ;
        RECT 20.145 53.620 26.175 54.060 ;
        RECT 20.145 53.565 20.605 53.620 ;
        RECT 25.715 53.515 26.175 53.620 ;
        RECT 22.405 48.870 22.885 48.935 ;
        RECT 22.405 48.550 24.205 48.870 ;
        RECT 22.405 48.385 22.885 48.550 ;
        RECT 23.635 45.710 24.195 48.550 ;
        RECT 27.515 45.710 27.995 45.735 ;
        RECT 23.635 45.290 27.995 45.710 ;
        RECT 23.635 45.280 24.195 45.290 ;
        RECT 27.515 45.185 27.995 45.290 ;
        RECT 20.745 40.120 21.225 40.225 ;
        RECT 24.545 40.120 25.105 40.130 ;
        RECT 20.745 39.700 25.105 40.120 ;
        RECT 20.745 39.675 21.225 39.700 ;
        RECT 24.545 36.860 25.105 39.700 ;
        RECT 25.855 36.860 26.335 37.025 ;
        RECT 24.535 36.540 26.335 36.860 ;
        RECT 25.855 36.475 26.335 36.540 ;
        RECT 22.565 31.790 23.025 31.895 ;
        RECT 28.135 31.790 28.595 31.845 ;
        RECT 22.565 31.350 28.595 31.790 ;
        RECT 22.565 31.325 23.025 31.350 ;
        RECT 28.135 31.275 28.595 31.350 ;
        RECT 29.765 12.265 30.255 73.120 ;
        RECT 38.960 73.080 41.730 74.510 ;
        RECT 31.345 54.070 31.805 54.145 ;
        RECT 36.915 54.070 37.375 54.095 ;
        RECT 31.345 53.630 37.375 54.070 ;
        RECT 31.345 53.575 31.805 53.630 ;
        RECT 36.915 53.525 37.375 53.630 ;
        RECT 33.605 48.880 34.085 48.945 ;
        RECT 33.605 48.560 35.405 48.880 ;
        RECT 33.605 48.395 34.085 48.560 ;
        RECT 34.835 45.720 35.395 48.560 ;
        RECT 38.715 45.720 39.195 45.745 ;
        RECT 34.835 45.300 39.195 45.720 ;
        RECT 34.835 45.290 35.395 45.300 ;
        RECT 38.715 45.195 39.195 45.300 ;
        RECT 32.025 40.120 32.505 40.225 ;
        RECT 35.825 40.120 36.385 40.130 ;
        RECT 32.025 39.700 36.385 40.120 ;
        RECT 32.025 39.675 32.505 39.700 ;
        RECT 35.825 36.860 36.385 39.700 ;
        RECT 37.135 36.860 37.615 37.025 ;
        RECT 35.815 36.540 37.615 36.860 ;
        RECT 37.135 36.475 37.615 36.540 ;
        RECT 33.845 31.790 34.305 31.895 ;
        RECT 39.415 31.790 39.875 31.845 ;
        RECT 33.845 31.350 39.875 31.790 ;
        RECT 33.845 31.325 34.305 31.350 ;
        RECT 39.415 31.275 39.875 31.350 ;
        RECT 41.055 12.360 41.545 73.080 ;
        RECT 49.930 73.030 52.530 74.650 ;
        RECT 61.330 74.530 63.890 75.690 ;
        RECT 73.135 75.580 73.765 80.495 ;
        RECT 84.425 75.690 85.055 81.995 ;
        RECT 72.340 74.980 74.900 75.580 ;
        RECT 42.565 54.040 43.025 54.115 ;
        RECT 48.135 54.040 48.595 54.065 ;
        RECT 42.565 53.600 48.595 54.040 ;
        RECT 42.565 53.545 43.025 53.600 ;
        RECT 48.135 53.495 48.595 53.600 ;
        RECT 44.825 48.850 45.305 48.915 ;
        RECT 44.825 48.530 46.625 48.850 ;
        RECT 44.825 48.365 45.305 48.530 ;
        RECT 46.055 45.690 46.615 48.530 ;
        RECT 49.935 45.690 50.415 45.715 ;
        RECT 46.055 45.270 50.415 45.690 ;
        RECT 46.055 45.260 46.615 45.270 ;
        RECT 49.935 45.165 50.415 45.270 ;
        RECT 43.315 40.100 43.795 40.205 ;
        RECT 47.115 40.100 47.675 40.110 ;
        RECT 43.315 39.680 47.675 40.100 ;
        RECT 43.315 39.655 43.795 39.680 ;
        RECT 47.115 36.840 47.675 39.680 ;
        RECT 48.425 36.840 48.905 37.005 ;
        RECT 47.105 36.520 48.905 36.840 ;
        RECT 48.425 36.455 48.905 36.520 ;
        RECT 45.135 31.770 45.595 31.875 ;
        RECT 50.705 31.770 51.165 31.825 ;
        RECT 45.135 31.330 51.165 31.770 ;
        RECT 45.135 31.305 45.595 31.330 ;
        RECT 50.705 31.255 51.165 31.330 ;
        RECT 41.055 12.350 41.555 12.360 ;
        RECT 28.345 11.115 30.465 12.265 ;
        RECT 41.065 11.965 41.555 12.350 ;
        RECT 51.635 12.145 52.125 73.030 ;
        RECT 61.260 73.010 64.060 74.530 ;
        RECT 72.340 73.050 75.020 74.980 ;
        RECT 83.730 74.540 86.290 75.690 ;
        RECT 95.655 75.580 96.285 83.245 ;
        RECT 106.975 75.640 107.605 84.485 ;
        RECT 118.225 75.650 118.855 85.545 ;
        RECT 129.975 75.650 130.605 86.595 ;
        RECT 133.330 76.605 136.060 77.855 ;
        RECT 137.190 76.585 139.920 77.835 ;
        RECT 53.815 54.020 54.275 54.095 ;
        RECT 59.385 54.020 59.845 54.045 ;
        RECT 53.815 53.580 59.845 54.020 ;
        RECT 53.815 53.525 54.275 53.580 ;
        RECT 59.385 53.475 59.845 53.580 ;
        RECT 56.075 48.830 56.555 48.895 ;
        RECT 56.075 48.510 57.875 48.830 ;
        RECT 56.075 48.345 56.555 48.510 ;
        RECT 57.305 45.670 57.865 48.510 ;
        RECT 61.185 45.670 61.665 45.695 ;
        RECT 57.305 45.250 61.665 45.670 ;
        RECT 57.305 45.240 57.865 45.250 ;
        RECT 61.185 45.145 61.665 45.250 ;
        RECT 54.535 40.100 55.015 40.205 ;
        RECT 58.335 40.100 58.895 40.110 ;
        RECT 54.535 39.680 58.895 40.100 ;
        RECT 54.535 39.655 55.015 39.680 ;
        RECT 58.335 36.840 58.895 39.680 ;
        RECT 59.645 36.840 60.125 37.005 ;
        RECT 58.325 36.520 60.125 36.840 ;
        RECT 59.645 36.455 60.125 36.520 ;
        RECT 56.355 31.770 56.815 31.875 ;
        RECT 61.925 31.770 62.385 31.825 ;
        RECT 56.355 31.330 62.385 31.770 ;
        RECT 56.355 31.305 56.815 31.330 ;
        RECT 61.925 31.255 62.385 31.330 ;
        RECT 29.765 11.100 30.255 11.115 ;
        RECT 39.065 11.005 41.615 11.965 ;
        RECT 50.285 10.995 52.405 12.145 ;
        RECT 62.915 12.135 63.405 73.010 ;
        RECT 65.035 54.010 65.495 54.085 ;
        RECT 70.605 54.010 71.065 54.035 ;
        RECT 65.035 53.570 71.065 54.010 ;
        RECT 65.035 53.515 65.495 53.570 ;
        RECT 70.605 53.465 71.065 53.570 ;
        RECT 67.295 48.820 67.775 48.885 ;
        RECT 67.295 48.500 69.095 48.820 ;
        RECT 67.295 48.335 67.775 48.500 ;
        RECT 68.525 45.660 69.085 48.500 ;
        RECT 72.405 45.660 72.885 45.685 ;
        RECT 68.525 45.240 72.885 45.660 ;
        RECT 68.525 45.230 69.085 45.240 ;
        RECT 72.405 45.135 72.885 45.240 ;
        RECT 65.735 40.100 66.215 40.205 ;
        RECT 69.535 40.100 70.095 40.110 ;
        RECT 65.735 39.680 70.095 40.100 ;
        RECT 65.735 39.655 66.215 39.680 ;
        RECT 69.535 36.840 70.095 39.680 ;
        RECT 70.845 36.840 71.325 37.005 ;
        RECT 69.525 36.520 71.325 36.840 ;
        RECT 70.845 36.455 71.325 36.520 ;
        RECT 67.555 31.770 68.015 31.875 ;
        RECT 73.125 31.770 73.585 31.825 ;
        RECT 67.555 31.330 73.585 31.770 ;
        RECT 67.555 31.305 68.015 31.330 ;
        RECT 73.125 31.255 73.585 31.330 ;
        RECT 74.055 12.165 74.545 73.050 ;
        RECT 83.690 73.000 86.290 74.540 ;
        RECT 94.960 74.710 97.520 75.580 ;
        RECT 94.960 73.020 97.570 74.710 ;
        RECT 106.340 74.460 108.900 75.640 ;
        RECT 117.470 74.720 120.030 75.650 ;
        RECT 76.275 54.000 76.735 54.075 ;
        RECT 81.845 54.000 82.305 54.025 ;
        RECT 76.275 53.560 82.305 54.000 ;
        RECT 76.275 53.505 76.735 53.560 ;
        RECT 81.845 53.455 82.305 53.560 ;
        RECT 78.535 48.810 79.015 48.875 ;
        RECT 78.535 48.490 80.335 48.810 ;
        RECT 78.535 48.325 79.015 48.490 ;
        RECT 79.765 45.650 80.325 48.490 ;
        RECT 83.645 45.650 84.125 45.675 ;
        RECT 79.765 45.230 84.125 45.650 ;
        RECT 79.765 45.220 80.325 45.230 ;
        RECT 83.645 45.125 84.125 45.230 ;
        RECT 77.025 40.090 77.505 40.195 ;
        RECT 80.825 40.090 81.385 40.100 ;
        RECT 77.025 39.670 81.385 40.090 ;
        RECT 77.025 39.645 77.505 39.670 ;
        RECT 80.825 36.830 81.385 39.670 ;
        RECT 82.135 36.830 82.615 36.995 ;
        RECT 80.815 36.510 82.615 36.830 ;
        RECT 82.135 36.445 82.615 36.510 ;
        RECT 78.845 31.760 79.305 31.865 ;
        RECT 84.415 31.760 84.875 31.815 ;
        RECT 78.845 31.320 84.875 31.760 ;
        RECT 78.845 31.295 79.305 31.320 ;
        RECT 84.415 31.245 84.875 31.320 ;
        RECT 61.365 10.985 63.485 12.135 ;
        RECT 72.675 11.015 74.795 12.165 ;
        RECT 85.375 12.155 85.865 73.000 ;
        RECT 87.525 54.010 87.985 54.085 ;
        RECT 93.095 54.010 93.555 54.035 ;
        RECT 87.525 53.570 93.555 54.010 ;
        RECT 87.525 53.515 87.985 53.570 ;
        RECT 93.095 53.465 93.555 53.570 ;
        RECT 89.785 48.820 90.265 48.885 ;
        RECT 89.785 48.500 91.585 48.820 ;
        RECT 89.785 48.335 90.265 48.500 ;
        RECT 91.015 45.660 91.575 48.500 ;
        RECT 94.895 45.660 95.375 45.685 ;
        RECT 91.015 45.240 95.375 45.660 ;
        RECT 91.015 45.230 91.575 45.240 ;
        RECT 94.895 45.135 95.375 45.240 ;
        RECT 88.265 40.110 88.745 40.215 ;
        RECT 92.065 40.110 92.625 40.120 ;
        RECT 88.265 39.690 92.625 40.110 ;
        RECT 88.265 39.665 88.745 39.690 ;
        RECT 92.065 36.850 92.625 39.690 ;
        RECT 93.375 36.850 93.855 37.015 ;
        RECT 92.055 36.530 93.855 36.850 ;
        RECT 93.375 36.465 93.855 36.530 ;
        RECT 90.085 31.780 90.545 31.885 ;
        RECT 95.655 31.780 96.115 31.835 ;
        RECT 90.085 31.340 96.115 31.780 ;
        RECT 90.085 31.315 90.545 31.340 ;
        RECT 95.655 31.265 96.115 31.340 ;
        RECT 96.605 12.155 97.095 73.020 ;
        RECT 106.150 73.000 109.060 74.460 ;
        RECT 117.470 73.070 120.000 74.720 ;
        RECT 129.290 74.650 131.850 75.650 ;
        RECT 129.300 73.140 131.820 74.650 ;
        RECT 98.805 54.000 99.265 54.075 ;
        RECT 104.375 54.000 104.835 54.025 ;
        RECT 98.805 53.560 104.835 54.000 ;
        RECT 98.805 53.505 99.265 53.560 ;
        RECT 104.375 53.455 104.835 53.560 ;
        RECT 101.065 48.810 101.545 48.875 ;
        RECT 101.065 48.490 102.865 48.810 ;
        RECT 101.065 48.325 101.545 48.490 ;
        RECT 102.295 45.650 102.855 48.490 ;
        RECT 106.175 45.650 106.655 45.675 ;
        RECT 102.295 45.230 106.655 45.650 ;
        RECT 102.295 45.220 102.855 45.230 ;
        RECT 106.175 45.125 106.655 45.230 ;
        RECT 99.475 40.130 99.955 40.235 ;
        RECT 103.275 40.130 103.835 40.140 ;
        RECT 99.475 39.710 103.835 40.130 ;
        RECT 99.475 39.685 99.955 39.710 ;
        RECT 103.275 36.870 103.835 39.710 ;
        RECT 104.585 36.870 105.065 37.035 ;
        RECT 103.265 36.550 105.065 36.870 ;
        RECT 104.585 36.485 105.065 36.550 ;
        RECT 101.295 31.800 101.755 31.905 ;
        RECT 106.865 31.800 107.325 31.855 ;
        RECT 101.295 31.360 107.325 31.800 ;
        RECT 101.295 31.335 101.755 31.360 ;
        RECT 106.865 31.285 107.325 31.360 ;
        RECT 107.865 12.205 108.355 73.000 ;
        RECT 110.075 54.000 110.535 54.075 ;
        RECT 115.645 54.000 116.105 54.025 ;
        RECT 110.075 53.560 116.105 54.000 ;
        RECT 110.075 53.505 110.535 53.560 ;
        RECT 115.645 53.455 116.105 53.560 ;
        RECT 112.335 48.810 112.815 48.875 ;
        RECT 112.335 48.490 114.135 48.810 ;
        RECT 112.335 48.325 112.815 48.490 ;
        RECT 113.565 45.650 114.125 48.490 ;
        RECT 117.445 45.650 117.925 45.675 ;
        RECT 113.565 45.230 117.925 45.650 ;
        RECT 113.565 45.220 114.125 45.230 ;
        RECT 117.445 45.125 117.925 45.230 ;
        RECT 110.675 40.170 111.155 40.275 ;
        RECT 114.475 40.170 115.035 40.180 ;
        RECT 110.675 39.750 115.035 40.170 ;
        RECT 110.675 39.725 111.155 39.750 ;
        RECT 114.475 36.910 115.035 39.750 ;
        RECT 115.785 36.910 116.265 37.075 ;
        RECT 114.465 36.590 116.265 36.910 ;
        RECT 115.785 36.525 116.265 36.590 ;
        RECT 112.495 31.840 112.955 31.945 ;
        RECT 118.065 31.840 118.525 31.895 ;
        RECT 112.495 31.400 118.525 31.840 ;
        RECT 112.495 31.375 112.955 31.400 ;
        RECT 118.065 31.325 118.525 31.400 ;
        RECT 119.085 12.205 119.575 73.070 ;
        RECT 121.325 54.000 121.785 54.075 ;
        RECT 126.895 54.000 127.355 54.025 ;
        RECT 121.325 53.560 127.355 54.000 ;
        RECT 121.325 53.505 121.785 53.560 ;
        RECT 126.895 53.455 127.355 53.560 ;
        RECT 123.585 48.810 124.065 48.875 ;
        RECT 123.585 48.490 125.385 48.810 ;
        RECT 123.585 48.325 124.065 48.490 ;
        RECT 124.815 45.650 125.375 48.490 ;
        RECT 128.695 45.650 129.175 45.675 ;
        RECT 124.815 45.230 129.175 45.650 ;
        RECT 124.815 45.220 125.375 45.230 ;
        RECT 128.695 45.125 129.175 45.230 ;
        RECT 121.885 40.190 122.365 40.295 ;
        RECT 125.685 40.190 126.245 40.200 ;
        RECT 121.885 39.770 126.245 40.190 ;
        RECT 121.885 39.745 122.365 39.770 ;
        RECT 125.685 36.930 126.245 39.770 ;
        RECT 126.995 36.930 127.475 37.095 ;
        RECT 125.675 36.610 127.475 36.930 ;
        RECT 126.995 36.545 127.475 36.610 ;
        RECT 123.705 31.860 124.165 31.965 ;
        RECT 129.275 31.860 129.735 31.915 ;
        RECT 123.705 31.420 129.735 31.860 ;
        RECT 123.705 31.395 124.165 31.420 ;
        RECT 129.275 31.345 129.735 31.420 ;
        RECT 130.335 12.235 130.825 73.140 ;
        RECT 74.055 11.010 74.545 11.015 ;
        RECT 83.795 11.005 85.915 12.155 ;
        RECT 95.095 11.005 97.215 12.155 ;
        RECT 106.285 11.055 108.405 12.205 ;
        RECT 117.515 11.055 119.635 12.205 ;
        RECT 128.815 11.085 130.935 12.235 ;
        RECT 107.865 11.010 108.355 11.055 ;
        RECT 119.085 11.050 119.575 11.055 ;
        RECT 85.375 11.000 85.865 11.005 ;
        RECT 96.605 10.980 97.095 11.005 ;
        RECT 74.290 0.135 75.680 1.435 ;
        RECT 93.500 0.205 94.890 1.505 ;
        RECT 112.900 0.335 114.290 1.635 ;
        RECT 131.800 0.405 133.540 1.905 ;
        RECT 151.600 0.275 152.970 1.445 ;
      LAYER met4 ;
        RECT 30.420 225.130 30.670 225.140 ;
        RECT 30.300 224.760 30.670 225.130 ;
        RECT 30.970 224.760 33.430 225.140 ;
        RECT 33.730 224.760 36.190 225.140 ;
        RECT 36.490 224.760 38.950 225.140 ;
        RECT 39.250 224.760 41.710 225.140 ;
        RECT 42.010 224.760 44.470 225.140 ;
        RECT 44.770 224.760 47.230 225.140 ;
        RECT 47.530 224.760 49.990 225.140 ;
        RECT 50.290 224.760 52.750 225.140 ;
        RECT 53.050 224.760 55.510 225.140 ;
        RECT 55.810 224.760 58.270 225.140 ;
        RECT 58.570 224.760 61.030 225.140 ;
        RECT 61.330 224.760 63.790 225.140 ;
        RECT 64.090 224.760 66.550 225.140 ;
        RECT 66.850 224.760 69.310 225.140 ;
        RECT 69.610 224.760 72.070 225.140 ;
        RECT 72.370 224.760 74.830 225.140 ;
        RECT 75.130 224.760 77.590 225.140 ;
        RECT 77.890 224.760 80.350 225.140 ;
        RECT 80.650 224.760 83.110 225.140 ;
        RECT 83.410 224.760 85.870 225.140 ;
        RECT 86.170 224.760 88.630 225.140 ;
        RECT 88.930 224.760 91.390 225.140 ;
        RECT 91.690 224.760 94.150 225.140 ;
        RECT 94.450 224.760 96.910 225.140 ;
        RECT 97.210 224.760 99.670 225.140 ;
        RECT 99.970 224.760 102.430 225.140 ;
        RECT 102.730 224.760 105.190 225.140 ;
        RECT 105.490 224.760 107.950 225.140 ;
        RECT 108.250 224.760 110.710 225.140 ;
        RECT 111.010 224.760 113.470 225.140 ;
        RECT 113.770 224.760 116.230 225.140 ;
        RECT 116.530 224.760 118.990 225.140 ;
        RECT 119.290 224.760 121.750 225.140 ;
        RECT 122.050 224.760 124.510 225.140 ;
        RECT 124.810 224.760 127.270 225.140 ;
        RECT 127.570 224.760 130.030 225.140 ;
        RECT 130.330 224.760 132.790 225.140 ;
        RECT 133.090 224.760 133.520 225.140 ;
        RECT 30.300 224.240 133.520 224.760 ;
        RECT 135.385 224.760 135.550 225.185 ;
        RECT 135.850 224.760 136.745 225.185 ;
        RECT 30.300 219.100 31.660 224.240 ;
        RECT 135.385 223.875 136.745 224.760 ;
        RECT 138.175 224.760 138.310 225.115 ;
        RECT 138.610 224.760 139.535 225.115 ;
        RECT 138.175 223.805 139.535 224.760 ;
        RECT 143.225 224.760 143.830 225.145 ;
        RECT 144.130 224.760 144.585 225.145 ;
        RECT 143.225 223.835 144.585 224.760 ;
        RECT 6.000 218.040 31.660 219.100 ;
        RECT 30.300 217.960 31.660 218.040 ;
        RECT 31.820 104.970 33.820 211.530 ;
        RECT 46.820 104.970 48.820 211.530 ;
        RECT 61.820 104.970 63.820 211.530 ;
        RECT 64.635 172.025 64.965 172.355 ;
        RECT 64.650 153.315 64.950 172.025 ;
        RECT 72.915 170.665 73.245 170.995 ;
        RECT 64.635 152.985 64.965 153.315 ;
        RECT 64.650 136.315 64.950 152.985 ;
        RECT 72.930 136.995 73.230 170.665 ;
        RECT 72.915 136.665 73.245 136.995 ;
        RECT 64.635 135.985 64.965 136.315 ;
        RECT 76.820 104.970 78.820 211.530 ;
        RECT 81.195 174.065 81.525 174.395 ;
        RECT 81.210 145.835 81.510 174.065 ;
        RECT 81.195 145.505 81.525 145.835 ;
        RECT 91.820 104.970 93.820 211.530 ;
        RECT 106.820 104.970 108.820 211.530 ;
        RECT 109.715 178.825 110.045 179.155 ;
        RECT 109.730 139.035 110.030 178.825 ;
        RECT 109.715 138.705 110.045 139.035 ;
        RECT 121.820 104.970 123.820 211.530 ;
        RECT 118.110 97.700 120.130 99.670 ;
        RECT 121.810 97.750 123.830 99.720 ;
        RECT 118.130 93.980 120.130 97.700 ;
        RECT 121.820 96.830 123.820 97.750 ;
        RECT 121.820 94.830 139.410 96.830 ;
        RECT 118.130 91.980 135.580 93.980 ;
        RECT 133.580 77.835 135.580 91.980 ;
        RECT 133.375 76.625 136.015 77.835 ;
        RECT 137.410 77.815 139.410 94.830 ;
        RECT 137.235 76.605 139.875 77.815 ;
        RECT 3.955 71.365 4.000 73.195 ;
        RECT 6.000 71.365 6.055 73.195 ;
        RECT 3.000 68.705 3.025 70.435 ;
        RECT 15.555 68.655 16.995 71.165 ;
        RECT 74.335 1.000 75.635 1.415 ;
        RECT 74.335 0.155 74.530 1.000 ;
        RECT 75.430 0.155 75.635 1.000 ;
        RECT 93.545 1.000 94.845 1.485 ;
        RECT 93.545 0.225 93.850 1.000 ;
        RECT 94.750 0.225 94.845 1.000 ;
        RECT 112.945 1.000 114.245 1.615 ;
        RECT 112.945 0.355 113.170 1.000 ;
        RECT 114.070 0.355 114.245 1.000 ;
        RECT 131.845 1.000 133.495 1.885 ;
        RECT 131.845 0.425 132.490 1.000 ;
        RECT 133.390 0.425 133.495 1.000 ;
        RECT 151.645 1.000 152.925 1.425 ;
        RECT 151.645 0.295 151.810 1.000 ;
        RECT 152.710 0.295 152.925 1.000 ;
  END
END tt_um_08_sws
END LIBRARY

