VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_08_sws
  CLASS BLOCK ;
  FOREIGN tt_um_08_sws ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    ANTENNAGATEAREA 200.000000 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    ANTENNAGATEAREA 550.000000 ;
    ANTENNADIFFAREA 2.900000 ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    ANTENNAGATEAREA 550.000000 ;
    ANTENNADIFFAREA 2.900000 ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    ANTENNADIFFAREA 29.000000 ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    ANTENNADIFFAREA 29.000000 ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    ANTENNADIFFAREA 394.109192 ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 29.985 211.185 30.155 211.375 ;
        RECT 31.420 211.235 31.540 211.345 ;
        RECT 36.885 211.185 37.055 211.375 ;
        RECT 38.725 211.185 38.895 211.375 ;
        RECT 44.245 211.185 44.415 211.375 ;
        RECT 49.765 211.185 49.935 211.375 ;
        RECT 51.605 211.185 51.775 211.375 ;
        RECT 57.125 211.185 57.295 211.375 ;
        RECT 62.645 211.185 62.815 211.375 ;
        RECT 64.485 211.185 64.655 211.375 ;
        RECT 70.005 211.185 70.175 211.375 ;
        RECT 75.525 211.185 75.695 211.375 ;
        RECT 77.365 211.185 77.535 211.375 ;
        RECT 82.885 211.185 83.055 211.375 ;
        RECT 88.405 211.185 88.575 211.375 ;
        RECT 90.245 211.185 90.415 211.375 ;
        RECT 95.765 211.185 95.935 211.375 ;
        RECT 101.285 211.185 101.455 211.375 ;
        RECT 103.125 211.185 103.295 211.375 ;
        RECT 108.645 211.185 108.815 211.375 ;
        RECT 114.165 211.185 114.335 211.375 ;
        RECT 115.140 211.235 115.260 211.345 ;
        RECT 120.605 211.185 120.775 211.375 ;
        RECT 126.125 211.185 126.295 211.375 ;
        RECT 127.505 211.185 127.675 211.375 ;
        RECT 29.845 210.375 31.215 211.185 ;
        RECT 31.685 210.375 37.195 211.185 ;
        RECT 37.215 210.315 37.645 211.100 ;
        RECT 37.665 210.375 39.035 211.185 ;
        RECT 39.045 210.375 44.555 211.185 ;
        RECT 44.565 210.375 50.075 211.185 ;
        RECT 50.095 210.315 50.525 211.100 ;
        RECT 50.545 210.375 51.915 211.185 ;
        RECT 51.925 210.375 57.435 211.185 ;
        RECT 57.445 210.375 62.955 211.185 ;
        RECT 62.975 210.315 63.405 211.100 ;
        RECT 63.425 210.375 64.795 211.185 ;
        RECT 64.805 210.375 70.315 211.185 ;
        RECT 70.325 210.375 75.835 211.185 ;
        RECT 75.855 210.315 76.285 211.100 ;
        RECT 76.305 210.375 77.675 211.185 ;
        RECT 77.685 210.375 83.195 211.185 ;
        RECT 83.205 210.375 88.715 211.185 ;
        RECT 88.735 210.315 89.165 211.100 ;
        RECT 89.185 210.375 90.555 211.185 ;
        RECT 90.565 210.375 96.075 211.185 ;
        RECT 96.085 210.375 101.595 211.185 ;
        RECT 101.615 210.315 102.045 211.100 ;
        RECT 102.065 210.375 103.435 211.185 ;
        RECT 103.445 210.375 108.955 211.185 ;
        RECT 108.965 210.375 114.475 211.185 ;
        RECT 114.495 210.315 114.925 211.100 ;
        RECT 115.405 210.375 120.915 211.185 ;
        RECT 120.925 210.375 126.435 211.185 ;
        RECT 126.445 210.375 127.815 211.185 ;
      LAYER nwell ;
        RECT 29.650 207.155 128.010 209.985 ;
      LAYER pwell ;
        RECT 29.845 205.955 31.215 206.765 ;
        RECT 31.685 205.955 33.515 206.765 ;
        RECT 33.525 205.955 39.035 206.765 ;
        RECT 39.045 205.955 44.555 206.765 ;
        RECT 44.565 205.955 50.075 206.765 ;
        RECT 50.095 206.040 50.525 206.825 ;
        RECT 51.465 205.955 55.135 206.765 ;
        RECT 55.145 205.955 60.655 206.765 ;
        RECT 60.665 205.955 66.175 206.765 ;
        RECT 66.185 206.635 67.105 206.865 ;
        RECT 69.935 206.635 70.865 206.855 ;
        RECT 66.185 205.955 75.375 206.635 ;
        RECT 75.855 206.040 76.285 206.825 ;
        RECT 76.305 205.955 77.675 206.735 ;
        RECT 78.145 206.665 79.075 206.865 ;
        RECT 80.410 206.665 81.355 206.865 ;
        RECT 78.145 206.185 81.355 206.665 ;
        RECT 78.285 205.985 81.355 206.185 ;
        RECT 29.985 205.745 30.155 205.955 ;
        RECT 31.420 205.795 31.540 205.905 ;
        RECT 33.205 205.765 33.375 205.955 ;
        RECT 36.885 205.745 37.055 205.935 ;
        RECT 37.860 205.795 37.980 205.905 ;
        RECT 38.725 205.765 38.895 205.955 ;
        RECT 40.565 205.745 40.735 205.935 ;
        RECT 44.245 205.765 44.415 205.955 ;
        RECT 46.085 205.745 46.255 205.935 ;
        RECT 49.765 205.765 49.935 205.955 ;
        RECT 51.145 205.800 51.305 205.910 ;
        RECT 51.605 205.745 51.775 205.935 ;
        RECT 54.825 205.765 54.995 205.955 ;
        RECT 57.125 205.745 57.295 205.935 ;
        RECT 60.345 205.765 60.515 205.955 ;
        RECT 62.645 205.745 62.815 205.935 ;
        RECT 65.865 205.765 66.035 205.955 ;
        RECT 66.785 205.745 66.955 205.935 ;
        RECT 68.165 205.745 68.335 205.935 ;
        RECT 75.065 205.765 75.235 205.955 ;
        RECT 75.580 205.795 75.700 205.905 ;
        RECT 76.445 205.765 76.615 205.955 ;
        RECT 77.880 205.795 78.000 205.905 ;
        RECT 78.285 205.765 78.455 205.985 ;
        RECT 80.410 205.955 81.355 205.985 ;
        RECT 81.365 206.635 82.285 206.865 ;
        RECT 85.115 206.635 86.045 206.855 ;
        RECT 81.365 205.955 90.555 206.635 ;
        RECT 91.495 205.955 92.845 206.865 ;
        RECT 93.325 205.955 96.075 206.765 ;
        RECT 96.085 205.955 101.595 206.765 ;
        RECT 101.615 206.040 102.045 206.825 ;
        RECT 102.525 205.955 104.355 206.765 ;
        RECT 104.365 205.955 109.875 206.765 ;
        RECT 109.885 205.955 115.395 206.765 ;
        RECT 115.405 205.955 120.915 206.765 ;
        RECT 120.925 205.955 126.435 206.765 ;
        RECT 126.445 205.955 127.815 206.765 ;
        RECT 78.745 205.745 78.915 205.935 ;
        RECT 81.965 205.745 82.135 205.935 ;
        RECT 84.265 205.745 84.435 205.935 ;
        RECT 85.185 205.790 85.345 205.900 ;
        RECT 85.645 205.745 85.815 205.935 ;
        RECT 90.245 205.745 90.415 205.955 ;
        RECT 91.165 205.800 91.325 205.910 ;
        RECT 91.630 205.745 91.800 205.935 ;
        RECT 92.545 205.765 92.715 205.955 ;
        RECT 93.005 205.905 93.175 205.935 ;
        RECT 93.005 205.795 93.180 205.905 ;
        RECT 93.005 205.745 93.175 205.795 ;
        RECT 95.305 205.745 95.475 205.935 ;
        RECT 95.765 205.905 95.935 205.955 ;
        RECT 95.765 205.795 95.940 205.905 ;
        RECT 95.765 205.765 95.935 205.795 ;
        RECT 97.605 205.745 97.775 205.935 ;
        RECT 101.285 205.765 101.455 205.955 ;
        RECT 102.260 205.795 102.380 205.905 ;
        RECT 103.125 205.745 103.295 205.935 ;
        RECT 104.045 205.765 104.215 205.955 ;
        RECT 108.645 205.745 108.815 205.935 ;
        RECT 109.565 205.765 109.735 205.955 ;
        RECT 114.165 205.745 114.335 205.935 ;
        RECT 115.085 205.905 115.255 205.955 ;
        RECT 115.085 205.795 115.260 205.905 ;
        RECT 115.085 205.765 115.255 205.795 ;
        RECT 120.605 205.745 120.775 205.955 ;
        RECT 126.125 205.745 126.295 205.955 ;
        RECT 127.505 205.745 127.675 205.955 ;
        RECT 29.845 204.935 31.215 205.745 ;
        RECT 31.685 204.935 37.195 205.745 ;
        RECT 37.215 204.875 37.645 205.660 ;
        RECT 38.125 204.935 40.875 205.745 ;
        RECT 40.885 204.935 46.395 205.745 ;
        RECT 46.405 204.935 51.915 205.745 ;
        RECT 51.925 204.935 57.435 205.745 ;
        RECT 57.445 204.935 62.955 205.745 ;
        RECT 62.975 204.875 63.405 205.660 ;
        RECT 63.425 204.935 67.095 205.745 ;
        RECT 67.115 204.835 68.465 205.745 ;
        RECT 68.685 205.065 79.055 205.745 ;
        RECT 68.685 204.835 70.895 205.065 ;
        RECT 73.615 204.845 74.545 205.065 ;
        RECT 79.065 204.835 82.175 205.745 ;
        RECT 82.285 205.065 84.575 205.745 ;
        RECT 82.285 204.835 83.205 205.065 ;
        RECT 85.605 204.835 88.715 205.745 ;
        RECT 88.735 204.875 89.165 205.660 ;
        RECT 89.195 204.835 90.545 205.745 ;
        RECT 90.565 204.835 91.915 205.745 ;
        RECT 92.875 204.835 94.225 205.745 ;
        RECT 94.245 204.965 95.615 205.745 ;
        RECT 96.085 204.935 97.915 205.745 ;
        RECT 97.925 204.935 103.435 205.745 ;
        RECT 103.445 204.935 108.955 205.745 ;
        RECT 108.965 204.935 114.475 205.745 ;
        RECT 114.495 204.875 114.925 205.660 ;
        RECT 115.405 204.935 120.915 205.745 ;
        RECT 120.925 204.935 126.435 205.745 ;
        RECT 126.445 204.935 127.815 205.745 ;
      LAYER nwell ;
        RECT 29.650 201.715 128.010 204.545 ;
      LAYER pwell ;
        RECT 29.845 200.515 31.215 201.325 ;
        RECT 31.685 200.515 33.515 201.325 ;
        RECT 33.525 200.515 39.035 201.325 ;
        RECT 39.045 200.515 44.555 201.325 ;
        RECT 44.565 200.515 50.075 201.325 ;
        RECT 50.095 200.600 50.525 201.385 ;
        RECT 50.545 200.515 51.915 201.325 ;
        RECT 51.925 200.515 57.435 201.325 ;
        RECT 57.445 200.515 62.955 201.325 ;
        RECT 62.965 200.515 68.475 201.325 ;
        RECT 68.495 200.515 69.845 201.425 ;
        RECT 72.520 201.195 73.440 201.425 ;
        RECT 69.975 200.515 73.440 201.195 ;
        RECT 74.005 200.515 75.835 201.325 ;
        RECT 75.855 200.600 76.285 201.385 ;
        RECT 76.305 201.225 77.235 201.425 ;
        RECT 78.570 201.225 79.515 201.425 ;
        RECT 76.305 200.745 79.515 201.225 ;
        RECT 76.445 200.545 79.515 200.745 ;
        RECT 29.985 200.305 30.155 200.515 ;
        RECT 31.420 200.355 31.540 200.465 ;
        RECT 33.205 200.325 33.375 200.515 ;
        RECT 36.885 200.305 37.055 200.495 ;
        RECT 38.725 200.325 38.895 200.515 ;
        RECT 41.025 200.305 41.195 200.495 ;
        RECT 44.245 200.325 44.415 200.515 ;
        RECT 46.545 200.305 46.715 200.495 ;
        RECT 49.765 200.325 49.935 200.515 ;
        RECT 51.605 200.325 51.775 200.515 ;
        RECT 52.065 200.305 52.235 200.495 ;
        RECT 52.525 200.305 52.695 200.495 ;
        RECT 56.205 200.305 56.375 200.495 ;
        RECT 57.125 200.325 57.295 200.515 ;
        RECT 59.940 200.355 60.060 200.465 ;
        RECT 62.645 200.305 62.815 200.515 ;
        RECT 63.620 200.355 63.740 200.465 ;
        RECT 65.405 200.305 65.575 200.495 ;
        RECT 65.865 200.305 66.035 200.495 ;
        RECT 68.165 200.325 68.335 200.515 ;
        RECT 68.625 200.325 68.795 200.515 ;
        RECT 70.005 200.325 70.175 200.515 ;
        RECT 75.525 200.495 75.695 200.515 ;
        RECT 72.305 200.305 72.475 200.495 ;
        RECT 73.740 200.355 73.860 200.465 ;
        RECT 75.520 200.325 75.695 200.495 ;
        RECT 76.040 200.355 76.160 200.465 ;
        RECT 76.445 200.325 76.615 200.545 ;
        RECT 78.570 200.515 79.515 200.545 ;
        RECT 79.525 201.195 80.445 201.425 ;
        RECT 83.275 201.195 84.205 201.415 ;
        RECT 88.725 201.195 89.645 201.425 ;
        RECT 92.475 201.195 93.405 201.415 ;
        RECT 79.525 200.515 88.715 201.195 ;
        RECT 88.725 200.515 97.915 201.195 ;
        RECT 97.925 200.515 101.595 201.325 ;
        RECT 101.615 200.600 102.045 201.385 ;
        RECT 102.985 200.515 106.655 201.325 ;
        RECT 109.320 201.195 110.240 201.425 ;
        RECT 106.775 200.515 110.240 201.195 ;
        RECT 110.345 201.195 111.265 201.425 ;
        RECT 114.095 201.195 115.025 201.415 ;
        RECT 110.345 200.515 119.535 201.195 ;
        RECT 119.545 200.515 120.915 201.325 ;
        RECT 120.925 200.515 126.435 201.325 ;
        RECT 126.445 200.515 127.815 201.325 ;
        RECT 75.520 200.305 75.690 200.325 ;
        RECT 77.825 200.305 77.995 200.495 ;
        RECT 78.290 200.305 78.460 200.495 ;
        RECT 83.805 200.305 83.975 200.495 ;
        RECT 84.725 200.350 84.885 200.460 ;
        RECT 85.185 200.305 85.355 200.495 ;
        RECT 88.405 200.325 88.575 200.515 ;
        RECT 91.165 200.325 91.335 200.495 ;
        RECT 91.165 200.305 91.330 200.325 ;
        RECT 91.625 200.305 91.795 200.495 ;
        RECT 94.385 200.305 94.555 200.495 ;
        RECT 95.765 200.305 95.935 200.495 ;
        RECT 96.225 200.305 96.395 200.495 ;
        RECT 97.605 200.325 97.775 200.515 ;
        RECT 98.985 200.305 99.155 200.495 ;
        RECT 99.445 200.305 99.615 200.495 ;
        RECT 101.285 200.325 101.455 200.515 ;
        RECT 102.665 200.360 102.825 200.470 ;
        RECT 106.345 200.325 106.515 200.515 ;
        RECT 106.805 200.325 106.975 200.515 ;
        RECT 109.565 200.305 109.735 200.495 ;
        RECT 110.080 200.355 110.200 200.465 ;
        RECT 113.890 200.305 114.060 200.495 ;
        RECT 116.005 200.305 116.175 200.495 ;
        RECT 116.520 200.355 116.640 200.465 ;
        RECT 116.925 200.305 117.095 200.495 ;
        RECT 118.765 200.350 118.925 200.460 ;
        RECT 119.225 200.305 119.395 200.515 ;
        RECT 120.605 200.465 120.775 200.515 ;
        RECT 120.605 200.355 120.780 200.465 ;
        RECT 120.605 200.325 120.775 200.355 ;
        RECT 126.125 200.305 126.295 200.515 ;
        RECT 127.505 200.305 127.675 200.515 ;
        RECT 29.845 199.495 31.215 200.305 ;
        RECT 31.685 199.495 37.195 200.305 ;
        RECT 37.215 199.435 37.645 200.220 ;
        RECT 37.665 199.495 41.335 200.305 ;
        RECT 41.345 199.495 46.855 200.305 ;
        RECT 46.865 199.495 52.375 200.305 ;
        RECT 52.495 199.625 55.960 200.305 ;
        RECT 56.175 199.625 59.640 200.305 ;
        RECT 55.040 199.395 55.960 199.625 ;
        RECT 58.720 199.395 59.640 199.625 ;
        RECT 60.205 199.495 62.955 200.305 ;
        RECT 62.975 199.435 63.405 200.220 ;
        RECT 63.885 199.495 65.715 200.305 ;
        RECT 65.735 199.395 67.085 200.305 ;
        RECT 67.105 199.495 72.615 200.305 ;
        RECT 72.915 199.395 75.835 200.305 ;
        RECT 76.305 199.625 78.135 200.305 ;
        RECT 76.305 199.395 77.650 199.625 ;
        RECT 78.145 199.395 80.435 200.305 ;
        RECT 80.445 199.625 84.115 200.305 ;
        RECT 85.155 199.625 88.620 200.305 ;
        RECT 80.445 199.395 81.375 199.625 ;
        RECT 87.700 199.395 88.620 199.625 ;
        RECT 88.735 199.435 89.165 200.220 ;
        RECT 89.495 199.625 91.330 200.305 ;
        RECT 91.485 199.625 93.315 200.305 ;
        RECT 89.495 199.395 90.425 199.625 ;
        RECT 93.335 199.395 94.685 200.305 ;
        RECT 94.705 199.495 96.075 200.305 ;
        RECT 96.085 199.525 97.455 200.305 ;
        RECT 97.465 199.495 99.295 200.305 ;
        RECT 99.315 199.395 100.665 200.305 ;
        RECT 100.685 199.625 109.875 200.305 ;
        RECT 110.575 199.625 114.475 200.305 ;
        RECT 100.685 199.395 101.605 199.625 ;
        RECT 104.435 199.405 105.365 199.625 ;
        RECT 113.545 199.395 114.475 199.625 ;
        RECT 114.495 199.435 114.925 200.220 ;
        RECT 114.955 199.395 116.305 200.305 ;
        RECT 116.795 199.395 118.145 200.305 ;
        RECT 119.085 199.525 120.455 200.305 ;
        RECT 120.925 199.495 126.435 200.305 ;
        RECT 126.445 199.495 127.815 200.305 ;
      LAYER nwell ;
        RECT 29.650 196.275 128.010 199.105 ;
      LAYER pwell ;
        RECT 29.845 195.075 31.215 195.885 ;
        RECT 32.145 195.075 37.655 195.885 ;
        RECT 37.665 195.075 43.175 195.885 ;
        RECT 43.185 195.075 48.695 195.885 ;
        RECT 48.705 195.075 50.075 195.855 ;
        RECT 50.095 195.160 50.525 195.945 ;
        RECT 51.005 195.075 52.375 195.855 ;
        RECT 52.395 195.075 53.745 195.985 ;
        RECT 56.420 195.755 57.340 195.985 ;
        RECT 53.875 195.075 57.340 195.755 ;
        RECT 57.455 195.075 58.805 195.985 ;
        RECT 58.825 195.075 60.195 195.855 ;
        RECT 60.300 195.755 61.220 195.985 ;
        RECT 67.085 195.755 68.015 195.985 ;
        RECT 60.300 195.075 63.765 195.755 ;
        RECT 64.115 195.075 68.015 195.755 ;
        RECT 68.025 195.075 69.395 195.855 ;
        RECT 70.325 195.075 75.835 195.885 ;
        RECT 75.855 195.160 76.285 195.945 ;
        RECT 77.225 195.075 80.895 195.885 ;
        RECT 80.915 195.755 83.915 195.985 ;
        RECT 86.875 195.755 87.795 195.985 ;
        RECT 80.915 195.665 85.495 195.755 ;
        RECT 80.905 195.305 85.495 195.665 ;
        RECT 80.905 195.115 81.835 195.305 ;
        RECT 80.915 195.075 81.835 195.115 ;
        RECT 83.925 195.075 85.495 195.305 ;
        RECT 85.505 195.075 87.795 195.755 ;
        RECT 87.805 195.075 89.635 195.755 ;
        RECT 89.645 195.075 92.395 195.885 ;
        RECT 92.415 195.075 93.765 195.985 ;
        RECT 96.440 195.755 97.360 195.985 ;
        RECT 100.665 195.755 101.595 195.985 ;
        RECT 93.895 195.075 97.360 195.755 ;
        RECT 97.695 195.075 101.595 195.755 ;
        RECT 101.615 195.160 102.045 195.945 ;
        RECT 102.065 195.075 105.735 195.885 ;
        RECT 105.745 195.075 107.115 195.855 ;
        RECT 107.125 195.075 108.495 195.885 ;
        RECT 108.505 195.075 109.875 195.855 ;
        RECT 113.085 195.755 114.015 195.985 ;
        RECT 110.115 195.075 114.015 195.755 ;
        RECT 114.025 195.755 114.945 195.985 ;
        RECT 117.775 195.755 118.705 195.975 ;
        RECT 114.025 195.075 123.215 195.755 ;
        RECT 123.685 195.075 126.435 195.885 ;
        RECT 126.445 195.075 127.815 195.885 ;
        RECT 29.985 194.865 30.155 195.075 ;
        RECT 31.420 194.915 31.540 195.025 ;
        RECT 31.825 194.920 31.985 195.030 ;
        RECT 36.885 194.865 37.055 195.055 ;
        RECT 37.345 194.885 37.515 195.075 ;
        RECT 42.865 194.865 43.035 195.075 ;
        RECT 43.325 194.865 43.495 195.055 ;
        RECT 44.705 194.865 44.875 195.055 ;
        RECT 48.385 194.885 48.555 195.075 ;
        RECT 49.765 194.885 49.935 195.075 ;
        RECT 50.740 194.915 50.860 195.025 ;
        RECT 52.065 194.885 52.235 195.075 ;
        RECT 53.445 194.885 53.615 195.075 ;
        RECT 53.905 194.885 54.075 195.075 ;
        RECT 58.505 194.885 58.675 195.075 ;
        RECT 58.965 194.885 59.135 195.075 ;
        RECT 62.645 194.865 62.815 195.055 ;
        RECT 63.565 194.885 63.735 195.075 ;
        RECT 67.430 194.885 67.600 195.075 ;
        RECT 68.165 194.885 68.335 195.075 ;
        RECT 70.005 194.920 70.165 195.030 ;
        RECT 72.305 194.865 72.475 195.055 ;
        RECT 73.225 194.910 73.385 195.020 ;
        RECT 73.685 194.865 73.855 195.055 ;
        RECT 75.525 194.885 75.695 195.075 ;
        RECT 76.905 194.920 77.065 195.030 ;
        RECT 78.745 194.885 78.915 195.055 ;
        RECT 80.585 194.885 80.755 195.075 ;
        RECT 81.965 194.885 82.135 195.055 ;
        RECT 85.185 194.885 85.355 195.075 ;
        RECT 85.645 194.885 85.815 195.075 ;
        RECT 87.945 194.885 88.115 195.075 ;
        RECT 75.625 194.865 75.695 194.885 ;
        RECT 78.845 194.865 78.915 194.885 ;
        RECT 82.065 194.865 82.135 194.885 ;
        RECT 88.405 194.865 88.575 195.055 ;
        RECT 89.325 194.865 89.495 195.055 ;
        RECT 92.085 194.885 92.255 195.075 ;
        RECT 92.545 194.885 92.715 195.075 ;
        RECT 93.925 194.885 94.095 195.075 ;
        RECT 99.905 194.865 100.075 195.055 ;
        RECT 100.420 194.915 100.540 195.025 ;
        RECT 101.010 194.885 101.180 195.075 ;
        RECT 104.045 194.865 104.215 195.055 ;
        RECT 104.505 194.865 104.675 195.055 ;
        RECT 105.425 194.885 105.595 195.075 ;
        RECT 105.885 194.865 106.055 195.075 ;
        RECT 108.185 194.885 108.355 195.075 ;
        RECT 108.645 194.885 108.815 195.075 ;
        RECT 112.785 194.865 112.955 195.055 ;
        RECT 113.245 194.865 113.415 195.055 ;
        RECT 113.430 194.885 113.600 195.075 ;
        RECT 118.305 194.865 118.475 195.055 ;
        RECT 118.820 194.915 118.940 195.025 ;
        RECT 120.605 194.865 120.775 195.055 ;
        RECT 122.905 194.885 123.075 195.075 ;
        RECT 123.420 194.915 123.540 195.025 ;
        RECT 126.125 194.865 126.295 195.075 ;
        RECT 127.505 194.865 127.675 195.075 ;
        RECT 29.845 194.055 31.215 194.865 ;
        RECT 31.685 194.055 37.195 194.865 ;
        RECT 37.215 193.995 37.645 194.780 ;
        RECT 37.665 194.055 43.175 194.865 ;
        RECT 43.195 193.955 44.545 194.865 ;
        RECT 44.565 194.185 53.755 194.865 ;
        RECT 49.075 193.965 50.005 194.185 ;
        RECT 52.835 193.955 53.755 194.185 ;
        RECT 53.765 194.185 62.955 194.865 ;
        RECT 53.765 193.955 54.685 194.185 ;
        RECT 57.515 193.965 58.445 194.185 ;
        RECT 62.975 193.995 63.405 194.780 ;
        RECT 63.425 194.185 72.615 194.865 ;
        RECT 73.545 194.185 75.375 194.865 ;
        RECT 63.425 193.955 64.345 194.185 ;
        RECT 67.175 193.965 68.105 194.185 ;
        RECT 74.030 193.955 75.375 194.185 ;
        RECT 75.625 194.635 77.895 194.865 ;
        RECT 78.845 194.635 81.115 194.865 ;
        RECT 82.065 194.635 84.335 194.865 ;
        RECT 75.625 193.955 78.380 194.635 ;
        RECT 78.845 193.955 81.600 194.635 ;
        RECT 82.065 193.955 84.820 194.635 ;
        RECT 85.045 194.055 88.715 194.865 ;
        RECT 88.735 193.995 89.165 194.780 ;
        RECT 89.195 193.955 90.545 194.865 ;
        RECT 90.935 194.185 100.215 194.865 ;
        RECT 90.935 194.065 93.270 194.185 ;
        RECT 90.935 193.955 91.855 194.065 ;
        RECT 97.935 193.965 98.855 194.185 ;
        RECT 100.685 194.055 104.355 194.865 ;
        RECT 104.375 193.955 105.725 194.865 ;
        RECT 105.855 194.185 109.320 194.865 ;
        RECT 108.400 193.955 109.320 194.185 ;
        RECT 109.520 194.185 112.985 194.865 ;
        RECT 109.520 193.955 110.440 194.185 ;
        RECT 113.105 194.085 114.475 194.865 ;
        RECT 114.495 193.995 114.925 194.780 ;
        RECT 115.040 194.185 118.505 194.865 ;
        RECT 115.040 193.955 115.960 194.185 ;
        RECT 119.085 194.055 120.915 194.865 ;
        RECT 120.925 194.055 126.435 194.865 ;
        RECT 126.445 194.055 127.815 194.865 ;
      LAYER nwell ;
        RECT 29.650 190.835 128.010 193.665 ;
      LAYER pwell ;
        RECT 29.845 189.635 31.215 190.445 ;
        RECT 31.225 189.635 36.735 190.445 ;
        RECT 39.400 190.315 40.320 190.545 ;
        RECT 36.855 189.635 40.320 190.315 ;
        RECT 40.795 190.435 41.715 190.545 ;
        RECT 40.795 190.315 43.130 190.435 ;
        RECT 47.795 190.315 48.715 190.535 ;
        RECT 40.795 189.635 50.075 190.315 ;
        RECT 50.095 189.720 50.525 190.505 ;
        RECT 50.545 190.315 51.475 190.545 ;
        RECT 50.545 189.635 54.445 190.315 ;
        RECT 55.155 189.635 56.505 190.545 ;
        RECT 56.525 190.315 57.455 190.545 ;
        RECT 63.865 190.315 64.795 190.545 ;
        RECT 56.525 189.635 60.425 190.315 ;
        RECT 60.895 189.635 64.795 190.315 ;
        RECT 64.805 190.315 65.725 190.545 ;
        RECT 68.555 190.315 69.485 190.535 ;
        RECT 74.490 190.315 75.835 190.545 ;
        RECT 64.805 189.635 73.995 190.315 ;
        RECT 74.005 189.635 75.835 190.315 ;
        RECT 75.855 189.720 76.285 190.505 ;
        RECT 78.805 190.315 81.805 190.545 ;
        RECT 77.225 190.225 81.805 190.315 ;
        RECT 77.225 189.865 81.815 190.225 ;
        RECT 77.225 189.635 78.795 189.865 ;
        RECT 80.885 189.675 81.815 189.865 ;
        RECT 80.885 189.635 81.805 189.675 ;
        RECT 81.825 189.635 83.195 190.445 ;
        RECT 86.405 190.315 87.335 190.545 ;
        RECT 83.435 189.635 87.335 190.315 ;
        RECT 87.715 190.435 88.635 190.545 ;
        RECT 87.715 190.315 90.050 190.435 ;
        RECT 94.715 190.315 95.635 190.535 ;
        RECT 87.715 189.635 96.995 190.315 ;
        RECT 97.005 189.635 98.375 190.415 ;
        RECT 98.395 189.635 99.745 190.545 ;
        RECT 99.765 189.635 101.595 190.445 ;
        RECT 101.615 189.720 102.045 190.505 ;
        RECT 102.525 190.315 103.445 190.545 ;
        RECT 106.275 190.315 107.205 190.535 ;
        RECT 115.845 190.315 116.775 190.545 ;
        RECT 102.525 189.635 111.715 190.315 ;
        RECT 112.875 189.635 116.775 190.315 ;
        RECT 116.785 190.315 117.705 190.545 ;
        RECT 120.535 190.315 121.465 190.535 ;
        RECT 116.785 189.635 125.975 190.315 ;
        RECT 126.445 189.635 127.815 190.445 ;
        RECT 29.985 189.425 30.155 189.635 ;
        RECT 31.420 189.475 31.540 189.585 ;
        RECT 34.125 189.425 34.295 189.615 ;
        RECT 34.585 189.425 34.755 189.615 ;
        RECT 35.965 189.425 36.135 189.615 ;
        RECT 36.425 189.445 36.595 189.635 ;
        RECT 36.885 189.445 37.055 189.635 ;
        RECT 46.545 189.425 46.715 189.615 ;
        RECT 49.765 189.445 49.935 189.635 ;
        RECT 50.410 189.425 50.580 189.615 ;
        RECT 50.960 189.445 51.130 189.635 ;
        RECT 51.145 189.425 51.315 189.615 ;
        RECT 54.880 189.475 55.000 189.585 ;
        RECT 55.285 189.445 55.455 189.635 ;
        RECT 56.940 189.445 57.110 189.635 ;
        RECT 61.265 189.425 61.435 189.615 ;
        RECT 62.645 189.425 62.815 189.615 ;
        RECT 63.620 189.475 63.740 189.585 ;
        RECT 64.025 189.425 64.195 189.615 ;
        RECT 64.210 189.445 64.380 189.635 ;
        RECT 68.625 189.425 68.795 189.615 ;
        RECT 72.305 189.425 72.475 189.615 ;
        RECT 73.685 189.445 73.855 189.635 ;
        RECT 74.145 189.445 74.315 189.635 ;
        RECT 75.525 189.445 75.695 189.615 ;
        RECT 76.905 189.480 77.065 189.590 ;
        RECT 77.365 189.445 77.535 189.635 ;
        RECT 78.285 189.425 78.455 189.615 ;
        RECT 78.745 189.445 78.915 189.615 ;
        RECT 78.845 189.425 78.915 189.445 ;
        RECT 81.970 189.425 82.140 189.615 ;
        RECT 82.885 189.445 83.055 189.635 ;
        RECT 86.750 189.445 86.920 189.635 ;
        RECT 88.130 189.425 88.300 189.615 ;
        RECT 89.785 189.470 89.945 189.580 ;
        RECT 90.245 189.425 90.415 189.615 ;
        RECT 96.685 189.445 96.855 189.635 ;
        RECT 98.065 189.445 98.235 189.635 ;
        RECT 98.525 189.445 98.695 189.635 ;
        RECT 101.285 189.445 101.455 189.635 ;
        RECT 102.260 189.475 102.380 189.585 ;
        RECT 108.185 189.425 108.355 189.615 ;
        RECT 108.920 189.425 109.090 189.615 ;
        RECT 111.405 189.445 111.575 189.635 ;
        RECT 112.325 189.480 112.485 189.590 ;
        RECT 112.785 189.425 112.955 189.615 ;
        RECT 114.220 189.475 114.340 189.585 ;
        RECT 116.190 189.445 116.360 189.635 ;
        RECT 123.825 189.425 123.995 189.615 ;
        RECT 124.340 189.475 124.460 189.585 ;
        RECT 125.665 189.445 125.835 189.635 ;
        RECT 126.125 189.585 126.295 189.615 ;
        RECT 126.125 189.475 126.300 189.585 ;
        RECT 126.125 189.425 126.295 189.475 ;
        RECT 127.505 189.425 127.675 189.635 ;
        RECT 29.845 188.615 31.215 189.425 ;
        RECT 31.685 188.615 34.435 189.425 ;
        RECT 34.455 188.515 35.805 189.425 ;
        RECT 35.835 188.515 37.185 189.425 ;
        RECT 37.215 188.555 37.645 189.340 ;
        RECT 37.665 188.745 46.855 189.425 ;
        RECT 47.095 188.745 50.995 189.425 ;
        RECT 37.665 188.515 38.585 188.745 ;
        RECT 41.415 188.525 42.345 188.745 ;
        RECT 50.065 188.515 50.995 188.745 ;
        RECT 51.005 188.645 52.375 189.425 ;
        RECT 52.385 188.745 61.575 189.425 ;
        RECT 52.385 188.515 53.305 188.745 ;
        RECT 56.135 188.525 57.065 188.745 ;
        RECT 61.595 188.515 62.945 189.425 ;
        RECT 62.975 188.555 63.405 189.340 ;
        RECT 63.885 188.645 65.255 189.425 ;
        RECT 65.360 188.745 68.825 189.425 ;
        RECT 69.040 188.745 72.505 189.425 ;
        RECT 73.005 188.745 75.430 189.425 ;
        RECT 75.855 188.745 78.595 189.425 ;
        RECT 78.845 189.195 81.115 189.425 ;
        RECT 65.360 188.515 66.280 188.745 ;
        RECT 69.040 188.515 69.960 188.745 ;
        RECT 78.845 188.515 81.600 189.195 ;
        RECT 81.825 188.515 84.435 189.425 ;
        RECT 84.815 188.745 88.715 189.425 ;
        RECT 87.785 188.515 88.715 188.745 ;
        RECT 88.735 188.555 89.165 189.340 ;
        RECT 90.105 188.745 99.210 189.425 ;
        RECT 99.305 188.745 108.495 189.425 ;
        RECT 108.505 188.745 112.405 189.425 ;
        RECT 99.305 188.515 100.225 188.745 ;
        RECT 103.055 188.525 103.985 188.745 ;
        RECT 108.505 188.515 109.435 188.745 ;
        RECT 112.655 188.515 114.005 189.425 ;
        RECT 114.495 188.555 114.925 189.340 ;
        RECT 114.945 188.745 124.135 189.425 ;
        RECT 114.945 188.515 115.865 188.745 ;
        RECT 118.695 188.525 119.625 188.745 ;
        RECT 124.605 188.615 126.435 189.425 ;
        RECT 126.445 188.615 127.815 189.425 ;
      LAYER nwell ;
        RECT 29.650 185.395 128.010 188.225 ;
      LAYER pwell ;
        RECT 29.845 184.195 31.215 185.005 ;
        RECT 33.880 184.875 34.800 185.105 ;
        RECT 31.335 184.195 34.800 184.875 ;
        RECT 34.905 184.875 35.825 185.105 ;
        RECT 38.655 184.875 39.585 185.095 ;
        RECT 47.305 184.875 48.235 185.105 ;
        RECT 34.905 184.195 44.095 184.875 ;
        RECT 44.335 184.195 48.235 184.875 ;
        RECT 48.715 184.195 50.065 185.105 ;
        RECT 50.095 184.280 50.525 185.065 ;
        RECT 54.120 184.875 55.040 185.105 ;
        RECT 51.575 184.195 55.040 184.875 ;
        RECT 55.340 184.195 58.815 185.105 ;
        RECT 71.225 184.875 72.155 185.105 ;
        RECT 58.910 184.195 68.015 184.875 ;
        RECT 68.255 184.195 72.155 184.875 ;
        RECT 72.260 184.875 73.180 185.105 ;
        RECT 72.260 184.195 75.725 184.875 ;
        RECT 75.855 184.280 76.285 185.065 ;
        RECT 79.550 184.875 80.895 185.105 ;
        RECT 76.315 184.195 79.055 184.875 ;
        RECT 79.065 184.195 80.895 184.875 ;
        RECT 81.365 184.195 84.840 185.105 ;
        RECT 88.245 184.875 89.175 185.105 ;
        RECT 85.275 184.195 89.175 184.875 ;
        RECT 89.185 184.875 90.105 185.105 ;
        RECT 92.935 184.875 93.865 185.095 ;
        RECT 89.185 184.195 98.375 184.875 ;
        RECT 98.385 184.195 99.755 184.975 ;
        RECT 100.225 184.195 101.595 184.975 ;
        RECT 101.615 184.280 102.045 185.065 ;
        RECT 102.065 184.875 102.995 185.105 ;
        RECT 106.300 184.875 107.220 185.105 ;
        RECT 102.065 184.195 105.965 184.875 ;
        RECT 106.300 184.195 109.765 184.875 ;
        RECT 109.885 184.195 113.360 185.105 ;
        RECT 117.225 184.875 118.155 185.105 ;
        RECT 114.255 184.195 118.155 184.875 ;
        RECT 118.260 184.875 119.180 185.105 ;
        RECT 118.260 184.195 121.725 184.875 ;
        RECT 121.845 184.195 123.215 184.975 ;
        RECT 123.225 184.195 124.595 184.975 ;
        RECT 124.605 184.195 126.435 185.005 ;
        RECT 126.445 184.195 127.815 185.005 ;
        RECT 29.985 183.985 30.155 184.195 ;
        RECT 31.365 184.005 31.535 184.195 ;
        RECT 31.825 184.030 31.985 184.140 ;
        RECT 33.205 183.985 33.375 184.175 ;
        RECT 33.665 183.985 33.835 184.175 ;
        RECT 38.265 184.030 38.425 184.140 ;
        RECT 38.725 183.985 38.895 184.175 ;
        RECT 40.380 183.985 40.550 184.175 ;
        RECT 43.785 184.005 43.955 184.195 ;
        RECT 47.650 184.005 47.820 184.195 ;
        RECT 48.440 184.035 48.560 184.145 ;
        RECT 48.845 184.005 49.015 184.195 ;
        RECT 51.145 184.040 51.305 184.150 ;
        RECT 51.605 184.005 51.775 184.195 ;
        RECT 52.985 183.985 53.155 184.175 ;
        RECT 53.720 183.985 53.890 184.175 ;
        RECT 57.585 183.985 57.755 184.175 ;
        RECT 58.500 184.005 58.670 184.195 ;
        RECT 59.020 184.035 59.140 184.145 ;
        RECT 62.640 183.985 62.810 184.175 ;
        RECT 63.620 184.035 63.740 184.145 ;
        RECT 67.430 183.985 67.600 184.175 ;
        RECT 67.705 184.005 67.875 184.195 ;
        RECT 71.570 184.005 71.740 184.195 ;
        RECT 75.525 184.005 75.695 184.195 ;
        RECT 76.905 183.985 77.075 184.175 ;
        RECT 77.365 183.985 77.535 184.175 ;
        RECT 78.745 184.005 78.915 184.195 ;
        RECT 79.205 184.005 79.375 184.195 ;
        RECT 80.130 183.985 80.300 184.175 ;
        RECT 81.100 184.035 81.220 184.145 ;
        RECT 81.510 184.005 81.680 184.195 ;
        RECT 83.810 183.985 83.980 184.175 ;
        RECT 87.485 183.985 87.655 184.175 ;
        RECT 88.590 184.005 88.760 184.195 ;
        RECT 98.065 184.005 98.235 184.195 ;
        RECT 99.445 184.005 99.615 184.195 ;
        RECT 99.900 184.145 100.070 184.175 ;
        RECT 99.900 184.035 100.080 184.145 ;
        RECT 99.900 183.985 100.070 184.035 ;
        RECT 100.365 184.005 100.535 184.195 ;
        RECT 102.480 184.005 102.650 184.195 ;
        RECT 103.585 183.985 103.755 184.175 ;
        RECT 104.050 183.985 104.220 184.175 ;
        RECT 107.730 183.985 107.900 184.175 ;
        RECT 109.565 184.005 109.735 184.195 ;
        RECT 110.030 184.005 110.200 184.195 ;
        RECT 111.460 184.035 111.580 184.145 ;
        RECT 111.865 183.985 112.035 184.175 ;
        RECT 113.245 183.985 113.415 184.175 ;
        RECT 113.760 184.035 113.880 184.145 ;
        RECT 115.090 183.985 115.260 184.175 ;
        RECT 117.570 184.005 117.740 184.195 ;
        RECT 118.765 183.985 118.935 184.175 ;
        RECT 121.525 184.005 121.695 184.195 ;
        RECT 121.985 184.005 122.155 184.195 ;
        RECT 122.445 183.985 122.615 184.175 ;
        RECT 123.365 184.005 123.535 184.195 ;
        RECT 126.125 183.985 126.295 184.195 ;
        RECT 127.505 183.985 127.675 184.195 ;
        RECT 29.845 183.175 31.215 183.985 ;
        RECT 32.155 183.075 33.505 183.985 ;
        RECT 33.635 183.305 37.100 183.985 ;
        RECT 36.180 183.075 37.100 183.305 ;
        RECT 37.215 183.115 37.645 183.900 ;
        RECT 38.585 183.205 39.955 183.985 ;
        RECT 39.965 183.305 43.865 183.985 ;
        RECT 44.105 183.305 53.295 183.985 ;
        RECT 53.305 183.305 57.205 183.985 ;
        RECT 39.965 183.075 40.895 183.305 ;
        RECT 44.105 183.075 45.025 183.305 ;
        RECT 47.855 183.085 48.785 183.305 ;
        RECT 53.305 183.075 54.235 183.305 ;
        RECT 57.445 183.205 58.815 183.985 ;
        RECT 59.480 183.075 62.955 183.985 ;
        RECT 62.975 183.115 63.405 183.900 ;
        RECT 64.115 183.305 68.015 183.985 ;
        RECT 67.085 183.075 68.015 183.305 ;
        RECT 68.025 183.305 77.215 183.985 ;
        RECT 68.025 183.075 68.945 183.305 ;
        RECT 71.775 183.085 72.705 183.305 ;
        RECT 77.225 183.075 79.945 183.985 ;
        RECT 79.985 183.075 83.460 183.985 ;
        RECT 83.665 183.075 87.140 183.985 ;
        RECT 87.355 183.075 88.705 183.985 ;
        RECT 88.735 183.115 89.165 183.900 ;
        RECT 89.205 183.075 100.215 183.985 ;
        RECT 100.320 183.305 103.785 183.985 ;
        RECT 100.320 183.075 101.240 183.305 ;
        RECT 103.905 183.075 107.380 183.985 ;
        RECT 107.585 183.075 111.060 183.985 ;
        RECT 111.735 183.075 113.085 183.985 ;
        RECT 113.115 183.075 114.465 183.985 ;
        RECT 114.495 183.115 114.925 183.900 ;
        RECT 114.945 183.075 118.420 183.985 ;
        RECT 118.735 183.305 122.200 183.985 ;
        RECT 121.280 183.075 122.200 183.305 ;
        RECT 122.305 183.205 123.675 183.985 ;
        RECT 123.685 183.175 126.435 183.985 ;
        RECT 126.445 183.175 127.815 183.985 ;
      LAYER nwell ;
        RECT 29.650 179.955 128.010 182.785 ;
      LAYER pwell ;
        RECT 29.845 178.755 31.215 179.565 ;
        RECT 31.685 178.755 35.160 179.665 ;
        RECT 35.560 178.755 39.035 179.665 ;
        RECT 39.045 178.755 42.520 179.665 ;
        RECT 45.380 179.435 46.300 179.665 ;
        RECT 42.835 178.755 46.300 179.435 ;
        RECT 46.600 178.755 50.075 179.665 ;
        RECT 50.095 178.840 50.525 179.625 ;
        RECT 50.740 178.755 54.215 179.665 ;
        RECT 54.225 178.755 57.700 179.665 ;
        RECT 58.000 179.435 58.920 179.665 ;
        RECT 64.240 179.435 65.160 179.665 ;
        RECT 58.000 178.755 61.465 179.435 ;
        RECT 61.695 178.755 65.160 179.435 ;
        RECT 65.265 178.755 67.095 179.565 ;
        RECT 67.105 178.755 70.580 179.665 ;
        RECT 70.785 178.755 72.155 179.535 ;
        RECT 72.165 179.435 73.510 179.665 ;
        RECT 74.005 179.435 75.350 179.665 ;
        RECT 72.165 178.755 73.995 179.435 ;
        RECT 74.005 178.755 75.835 179.435 ;
        RECT 75.855 178.840 76.285 179.625 ;
        RECT 76.305 179.435 77.650 179.665 ;
        RECT 76.305 178.755 78.135 179.435 ;
        RECT 78.145 178.755 79.515 179.565 ;
        RECT 79.525 178.755 82.135 179.665 ;
        RECT 82.480 178.755 85.955 179.665 ;
        RECT 86.335 179.555 87.255 179.665 ;
        RECT 86.335 179.435 88.670 179.555 ;
        RECT 93.335 179.435 94.255 179.655 ;
        RECT 86.335 178.755 95.615 179.435 ;
        RECT 95.635 178.755 96.985 179.665 ;
        RECT 100.580 179.435 101.500 179.665 ;
        RECT 98.035 178.755 101.500 179.435 ;
        RECT 101.615 178.840 102.045 179.625 ;
        RECT 102.065 178.755 103.435 179.535 ;
        RECT 103.905 178.755 105.735 179.565 ;
        RECT 105.940 178.755 109.415 179.665 ;
        RECT 109.425 178.755 112.900 179.665 ;
        RECT 115.760 179.435 116.680 179.665 ;
        RECT 113.215 178.755 116.680 179.435 ;
        RECT 116.785 179.435 117.705 179.665 ;
        RECT 120.535 179.435 121.465 179.655 ;
        RECT 116.785 178.755 125.975 179.435 ;
        RECT 126.445 178.755 127.815 179.565 ;
        RECT 29.985 178.545 30.155 178.755 ;
        RECT 31.420 178.595 31.540 178.705 ;
        RECT 31.830 178.565 32.000 178.755 ;
        RECT 34.125 178.545 34.295 178.735 ;
        RECT 34.585 178.545 34.755 178.735 ;
        RECT 35.965 178.545 36.135 178.735 ;
        RECT 37.805 178.545 37.975 178.735 ;
        RECT 38.720 178.565 38.890 178.755 ;
        RECT 39.190 178.565 39.360 178.755 ;
        RECT 42.865 178.565 43.035 178.755 ;
        RECT 47.010 178.545 47.180 178.735 ;
        RECT 49.760 178.565 49.930 178.755 ;
        RECT 50.685 178.545 50.855 178.735 ;
        RECT 53.900 178.565 54.070 178.755 ;
        RECT 54.370 178.565 54.540 178.755 ;
        RECT 59.940 178.595 60.060 178.705 ;
        RECT 60.345 178.545 60.515 178.735 ;
        RECT 61.265 178.565 61.435 178.755 ;
        RECT 61.725 178.565 61.895 178.755 ;
        RECT 62.645 178.545 62.815 178.735 ;
        RECT 63.565 178.545 63.735 178.735 ;
        RECT 66.785 178.565 66.955 178.755 ;
        RECT 67.250 178.565 67.420 178.755 ;
        RECT 70.465 178.545 70.635 178.735 ;
        RECT 70.925 178.565 71.095 178.755 ;
        RECT 71.845 178.545 72.015 178.735 ;
        RECT 73.685 178.565 73.855 178.755 ;
        RECT 74.605 178.545 74.775 178.735 ;
        RECT 75.525 178.565 75.695 178.755 ;
        RECT 76.445 178.545 76.615 178.735 ;
        RECT 76.905 178.545 77.075 178.735 ;
        RECT 77.825 178.565 77.995 178.755 ;
        RECT 79.205 178.565 79.375 178.755 ;
        RECT 79.670 178.735 79.840 178.755 ;
        RECT 79.665 178.565 79.840 178.735 ;
        RECT 82.480 178.595 82.600 178.705 ;
        RECT 79.665 178.545 79.835 178.565 ;
        RECT 84.265 178.545 84.435 178.735 ;
        RECT 85.640 178.565 85.810 178.755 ;
        RECT 87.945 178.545 88.115 178.735 ;
        RECT 88.460 178.595 88.580 178.705 ;
        RECT 89.325 178.545 89.495 178.735 ;
        RECT 90.705 178.545 90.875 178.735 ;
        RECT 95.305 178.545 95.475 178.755 ;
        RECT 95.765 178.565 95.935 178.755 ;
        RECT 96.225 178.590 96.385 178.700 ;
        RECT 97.605 178.600 97.765 178.710 ;
        RECT 98.065 178.565 98.235 178.755 ;
        RECT 102.205 178.565 102.375 178.755 ;
        RECT 103.640 178.595 103.760 178.705 ;
        RECT 105.425 178.545 105.595 178.755 ;
        RECT 105.885 178.545 106.055 178.735 ;
        RECT 107.320 178.595 107.440 178.705 ;
        RECT 109.100 178.565 109.270 178.755 ;
        RECT 109.570 178.565 109.740 178.755 ;
        RECT 110.025 178.545 110.195 178.735 ;
        RECT 113.245 178.565 113.415 178.755 ;
        RECT 113.890 178.545 114.060 178.735 ;
        RECT 115.085 178.545 115.255 178.735 ;
        RECT 125.205 178.545 125.375 178.735 ;
        RECT 125.665 178.565 125.835 178.755 ;
        RECT 126.180 178.700 126.300 178.705 ;
        RECT 126.125 178.595 126.300 178.700 ;
        RECT 126.125 178.590 126.285 178.595 ;
        RECT 127.505 178.545 127.675 178.755 ;
        RECT 29.845 177.735 31.215 178.545 ;
        RECT 31.685 177.735 34.435 178.545 ;
        RECT 34.445 177.765 35.815 178.545 ;
        RECT 35.835 177.635 37.185 178.545 ;
        RECT 37.215 177.675 37.645 178.460 ;
        RECT 37.665 177.865 46.855 178.545 ;
        RECT 42.175 177.645 43.105 177.865 ;
        RECT 45.935 177.635 46.855 177.865 ;
        RECT 46.865 177.635 50.340 178.545 ;
        RECT 50.545 177.865 59.735 178.545 ;
        RECT 55.055 177.645 55.985 177.865 ;
        RECT 58.815 177.635 59.735 177.865 ;
        RECT 60.205 177.765 61.575 178.545 ;
        RECT 61.585 177.735 62.955 178.545 ;
        RECT 62.975 177.675 63.405 178.460 ;
        RECT 63.535 177.865 67.000 178.545 ;
        RECT 66.080 177.635 67.000 177.865 ;
        RECT 67.105 177.735 70.775 178.545 ;
        RECT 70.795 177.635 72.145 178.545 ;
        RECT 72.165 177.735 74.915 178.545 ;
        RECT 74.925 177.865 76.755 178.545 ;
        RECT 76.765 177.865 79.505 178.545 ;
        RECT 74.925 177.635 76.270 177.865 ;
        RECT 79.525 177.635 82.245 178.545 ;
        RECT 82.745 177.735 84.575 178.545 ;
        RECT 84.680 177.865 88.145 178.545 ;
        RECT 84.680 177.635 85.600 177.865 ;
        RECT 88.735 177.675 89.165 178.460 ;
        RECT 89.195 177.635 90.545 178.545 ;
        RECT 90.675 177.865 94.140 178.545 ;
        RECT 93.220 177.635 94.140 177.865 ;
        RECT 94.245 177.765 95.615 178.545 ;
        RECT 96.545 177.865 105.735 178.545 ;
        RECT 96.545 177.635 97.465 177.865 ;
        RECT 100.295 177.645 101.225 177.865 ;
        RECT 105.755 177.635 107.105 178.545 ;
        RECT 107.585 177.735 110.335 178.545 ;
        RECT 110.575 177.865 114.475 178.545 ;
        RECT 113.545 177.635 114.475 177.865 ;
        RECT 114.495 177.675 114.925 178.460 ;
        RECT 114.955 177.635 116.305 178.545 ;
        RECT 116.325 177.865 125.515 178.545 ;
        RECT 116.325 177.635 117.245 177.865 ;
        RECT 120.075 177.645 121.005 177.865 ;
        RECT 126.445 177.735 127.815 178.545 ;
      LAYER nwell ;
        RECT 29.650 174.515 128.010 177.345 ;
      LAYER pwell ;
        RECT 29.845 173.315 31.215 174.125 ;
        RECT 31.595 174.115 32.515 174.225 ;
        RECT 31.595 173.995 33.930 174.115 ;
        RECT 38.595 173.995 39.515 174.215 ;
        RECT 41.440 173.995 42.360 174.225 ;
        RECT 45.120 173.995 46.040 174.225 ;
        RECT 31.595 173.315 40.875 173.995 ;
        RECT 41.440 173.315 44.905 173.995 ;
        RECT 45.120 173.315 48.585 173.995 ;
        RECT 48.715 173.315 50.065 174.225 ;
        RECT 50.095 173.400 50.525 174.185 ;
        RECT 50.545 173.315 52.375 174.125 ;
        RECT 52.395 173.315 53.745 174.225 ;
        RECT 53.765 173.995 54.685 174.225 ;
        RECT 57.515 173.995 58.445 174.215 ;
        RECT 62.965 173.995 63.895 174.225 ;
        RECT 53.765 173.315 62.955 173.995 ;
        RECT 62.965 173.315 66.865 173.995 ;
        RECT 67.105 173.315 69.855 174.125 ;
        RECT 69.875 173.315 71.225 174.225 ;
        RECT 71.245 173.315 72.615 174.095 ;
        RECT 73.225 173.315 75.835 174.225 ;
        RECT 75.855 173.400 76.285 174.185 ;
        RECT 76.905 173.315 79.515 174.225 ;
        RECT 80.445 173.315 83.185 173.995 ;
        RECT 83.205 173.315 85.035 174.125 ;
        RECT 85.415 174.115 86.335 174.225 ;
        RECT 85.415 173.995 87.750 174.115 ;
        RECT 92.415 173.995 93.335 174.215 ;
        RECT 85.415 173.315 94.695 173.995 ;
        RECT 95.635 173.315 96.985 174.225 ;
        RECT 100.205 173.995 101.135 174.225 ;
        RECT 97.235 173.315 101.135 173.995 ;
        RECT 101.615 173.400 102.045 174.185 ;
        RECT 102.065 173.315 105.225 174.225 ;
        RECT 106.205 173.995 107.125 174.225 ;
        RECT 109.955 173.995 110.885 174.215 ;
        RECT 119.065 173.995 119.995 174.225 ;
        RECT 106.205 173.315 115.395 173.995 ;
        RECT 116.095 173.315 119.995 173.995 ;
        RECT 120.100 173.995 121.020 174.225 ;
        RECT 120.100 173.315 123.565 173.995 ;
        RECT 123.685 173.315 125.515 173.995 ;
        RECT 126.445 173.315 127.815 174.125 ;
        RECT 29.985 173.105 30.155 173.315 ;
        RECT 34.585 173.105 34.755 173.295 ;
        RECT 35.965 173.105 36.135 173.295 ;
        RECT 36.885 173.150 37.045 173.260 ;
        RECT 38.265 173.150 38.425 173.260 ;
        RECT 39.645 173.105 39.815 173.295 ;
        RECT 40.565 173.125 40.735 173.315 ;
        RECT 41.025 173.265 41.195 173.295 ;
        RECT 41.025 173.155 41.200 173.265 ;
        RECT 41.025 173.105 41.195 173.155 ;
        RECT 41.760 173.105 41.930 173.295 ;
        RECT 44.705 173.125 44.875 173.315 ;
        RECT 45.680 173.155 45.800 173.265 ;
        RECT 46.085 173.105 46.255 173.295 ;
        RECT 48.385 173.125 48.555 173.315 ;
        RECT 48.845 173.125 49.015 173.315 ;
        RECT 50.040 173.105 50.210 173.295 ;
        RECT 52.065 173.125 52.235 173.315 ;
        RECT 52.525 173.125 52.695 173.315 ;
        RECT 62.645 173.105 62.815 173.315 ;
        RECT 63.380 173.125 63.550 173.315 ;
        RECT 63.565 173.105 63.735 173.295 ;
        RECT 69.545 173.125 69.715 173.315 ;
        RECT 70.925 173.125 71.095 173.315 ;
        RECT 71.385 173.125 71.555 173.315 ;
        RECT 72.820 173.155 72.940 173.265 ;
        RECT 73.685 173.105 73.855 173.295 ;
        RECT 74.605 173.150 74.765 173.260 ;
        RECT 75.520 173.125 75.690 173.315 ;
        RECT 76.500 173.155 76.620 173.265 ;
        RECT 77.365 173.105 77.535 173.295 ;
        RECT 77.880 173.155 78.000 173.265 ;
        RECT 79.200 173.125 79.370 173.315 ;
        RECT 79.665 173.105 79.835 173.295 ;
        RECT 80.125 173.265 80.285 173.270 ;
        RECT 80.125 173.160 80.300 173.265 ;
        RECT 80.180 173.155 80.300 173.160 ;
        RECT 80.585 173.125 80.755 173.315 ;
        RECT 82.885 173.105 83.055 173.295 ;
        RECT 84.265 173.105 84.435 173.295 ;
        RECT 84.725 173.125 84.895 173.315 ;
        RECT 88.130 173.105 88.300 173.295 ;
        RECT 89.785 173.150 89.945 173.260 ;
        RECT 90.245 173.105 90.415 173.295 ;
        RECT 94.385 173.125 94.555 173.315 ;
        RECT 95.305 173.160 95.465 173.270 ;
        RECT 95.765 173.125 95.935 173.315 ;
        RECT 100.550 173.125 100.720 173.315 ;
        RECT 101.340 173.155 101.460 173.265 ;
        RECT 104.965 173.125 105.135 173.315 ;
        RECT 105.885 173.160 106.045 173.270 ;
        RECT 108.645 173.105 108.815 173.295 ;
        RECT 110.025 173.105 110.195 173.295 ;
        RECT 113.705 173.105 113.875 173.295 ;
        RECT 114.220 173.155 114.340 173.265 ;
        RECT 115.085 173.125 115.255 173.315 ;
        RECT 115.600 173.260 115.720 173.265 ;
        RECT 115.545 173.155 115.720 173.260 ;
        RECT 115.545 173.150 115.705 173.155 ;
        RECT 119.410 173.105 119.580 173.315 ;
        RECT 120.145 173.105 120.315 173.295 ;
        RECT 121.525 173.105 121.695 173.295 ;
        RECT 122.905 173.105 123.075 173.295 ;
        RECT 123.365 173.125 123.535 173.315 ;
        RECT 124.340 173.155 124.460 173.265 ;
        RECT 125.205 173.125 125.375 173.315 ;
        RECT 126.125 173.105 126.295 173.295 ;
        RECT 127.505 173.105 127.675 173.315 ;
        RECT 29.845 172.295 31.215 173.105 ;
        RECT 31.225 172.295 34.895 173.105 ;
        RECT 34.915 172.195 36.265 173.105 ;
        RECT 37.215 172.235 37.645 173.020 ;
        RECT 38.585 172.325 39.955 173.105 ;
        RECT 39.965 172.325 41.335 173.105 ;
        RECT 41.345 172.425 45.245 173.105 ;
        RECT 46.055 172.425 49.520 173.105 ;
        RECT 41.345 172.195 42.275 172.425 ;
        RECT 48.600 172.195 49.520 172.425 ;
        RECT 49.625 172.425 53.525 173.105 ;
        RECT 53.850 172.425 62.955 173.105 ;
        RECT 49.625 172.195 50.555 172.425 ;
        RECT 62.975 172.235 63.405 173.020 ;
        RECT 63.435 172.195 64.785 173.105 ;
        RECT 64.805 172.425 73.995 173.105 ;
        RECT 74.935 172.425 77.675 173.105 ;
        RECT 78.145 172.425 79.975 173.105 ;
        RECT 64.805 172.195 65.725 172.425 ;
        RECT 68.555 172.205 69.485 172.425 ;
        RECT 78.145 172.195 79.490 172.425 ;
        RECT 80.445 172.295 83.195 173.105 ;
        RECT 83.215 172.195 84.565 173.105 ;
        RECT 84.815 172.425 88.715 173.105 ;
        RECT 87.785 172.195 88.715 172.425 ;
        RECT 88.735 172.235 89.165 173.020 ;
        RECT 90.105 172.425 99.210 173.105 ;
        RECT 99.675 172.425 108.955 173.105 ;
        RECT 99.675 172.305 102.010 172.425 ;
        RECT 99.675 172.195 100.595 172.305 ;
        RECT 106.675 172.205 107.595 172.425 ;
        RECT 108.965 172.325 110.335 173.105 ;
        RECT 110.440 172.425 113.905 173.105 ;
        RECT 110.440 172.195 111.360 172.425 ;
        RECT 114.495 172.235 114.925 173.020 ;
        RECT 116.095 172.425 119.995 173.105 ;
        RECT 119.065 172.195 119.995 172.425 ;
        RECT 120.015 172.195 121.365 173.105 ;
        RECT 121.385 172.325 122.755 173.105 ;
        RECT 122.765 172.325 124.135 173.105 ;
        RECT 124.605 172.295 126.435 173.105 ;
        RECT 126.445 172.295 127.815 173.105 ;
      LAYER nwell ;
        RECT 29.650 169.075 128.010 171.905 ;
      LAYER pwell ;
        RECT 29.845 167.875 31.215 168.685 ;
        RECT 31.595 168.675 32.515 168.785 ;
        RECT 31.595 168.555 33.930 168.675 ;
        RECT 38.595 168.555 39.515 168.775 ;
        RECT 40.885 168.555 41.815 168.785 ;
        RECT 31.595 167.875 40.875 168.555 ;
        RECT 40.885 167.875 44.785 168.555 ;
        RECT 45.025 167.875 46.395 168.685 ;
        RECT 46.600 167.875 50.075 168.785 ;
        RECT 50.095 167.960 50.525 168.745 ;
        RECT 51.005 167.875 52.375 168.655 ;
        RECT 52.580 167.875 56.055 168.785 ;
        RECT 58.720 168.555 59.640 168.785 ;
        RECT 56.175 167.875 59.640 168.555 ;
        RECT 59.840 167.875 63.710 168.785 ;
        RECT 63.885 167.875 66.635 168.685 ;
        RECT 66.645 168.555 67.565 168.785 ;
        RECT 70.395 168.555 71.325 168.775 ;
        RECT 66.645 167.875 75.835 168.555 ;
        RECT 75.855 167.960 76.285 168.745 ;
        RECT 77.225 168.555 78.570 168.785 ;
        RECT 79.065 168.555 80.410 168.785 ;
        RECT 77.225 167.875 79.055 168.555 ;
        RECT 79.065 167.875 80.895 168.555 ;
        RECT 80.905 167.875 82.275 168.685 ;
        RECT 82.285 167.875 85.760 168.785 ;
        RECT 89.165 168.555 90.095 168.785 ;
        RECT 86.195 167.875 90.095 168.555 ;
        RECT 90.565 167.875 91.935 168.655 ;
        RECT 91.945 167.875 93.315 168.685 ;
        RECT 95.980 168.555 96.900 168.785 ;
        RECT 100.205 168.555 101.135 168.785 ;
        RECT 93.435 167.875 96.900 168.555 ;
        RECT 97.235 167.875 101.135 168.555 ;
        RECT 101.615 167.960 102.045 168.745 ;
        RECT 102.065 167.875 103.435 168.685 ;
        RECT 106.645 168.555 107.575 168.785 ;
        RECT 103.675 167.875 107.575 168.555 ;
        RECT 107.585 167.875 108.955 168.685 ;
        RECT 108.965 167.875 110.335 168.655 ;
        RECT 113.545 168.555 114.475 168.785 ;
        RECT 110.575 167.875 114.475 168.555 ;
        RECT 114.945 167.875 116.775 168.685 ;
        RECT 116.785 168.555 117.705 168.785 ;
        RECT 120.535 168.555 121.465 168.775 ;
        RECT 116.785 167.875 125.975 168.555 ;
        RECT 126.445 167.875 127.815 168.685 ;
        RECT 29.985 167.665 30.155 167.875 ;
        RECT 31.420 167.715 31.540 167.825 ;
        RECT 34.125 167.665 34.295 167.855 ;
        RECT 35.505 167.665 35.675 167.855 ;
        RECT 36.885 167.665 37.055 167.855 ;
        RECT 37.805 167.665 37.975 167.855 ;
        RECT 40.565 167.685 40.735 167.875 ;
        RECT 41.300 167.685 41.470 167.875 ;
        RECT 46.085 167.855 46.255 167.875 ;
        RECT 42.405 167.665 42.575 167.855 ;
        RECT 46.080 167.685 46.255 167.855 ;
        RECT 49.760 167.685 49.930 167.875 ;
        RECT 46.080 167.665 46.250 167.685 ;
        RECT 49.950 167.665 50.120 167.855 ;
        RECT 50.685 167.825 50.855 167.855 ;
        RECT 50.685 167.715 50.860 167.825 ;
        RECT 50.685 167.665 50.855 167.715 ;
        RECT 51.145 167.685 51.315 167.875 ;
        RECT 55.280 167.665 55.450 167.855 ;
        RECT 55.740 167.685 55.910 167.875 ;
        RECT 56.020 167.665 56.190 167.855 ;
        RECT 56.205 167.685 56.375 167.875 ;
        RECT 63.565 167.855 63.710 167.875 ;
        RECT 59.940 167.715 60.060 167.825 ;
        RECT 62.645 167.665 62.815 167.855 ;
        RECT 63.565 167.685 63.735 167.855 ;
        RECT 64.945 167.665 65.115 167.855 ;
        RECT 65.680 167.665 65.850 167.855 ;
        RECT 66.325 167.685 66.495 167.875 ;
        RECT 72.950 167.665 73.120 167.855 ;
        RECT 73.740 167.715 73.860 167.825 ;
        RECT 75.525 167.685 75.695 167.875 ;
        RECT 76.440 167.665 76.610 167.855 ;
        RECT 76.905 167.825 77.065 167.830 ;
        RECT 76.905 167.720 77.080 167.825 ;
        RECT 76.960 167.715 77.080 167.720 ;
        RECT 78.745 167.665 78.915 167.875 ;
        RECT 80.585 167.665 80.755 167.875 ;
        RECT 81.050 167.665 81.220 167.855 ;
        RECT 81.965 167.685 82.135 167.875 ;
        RECT 82.430 167.685 82.600 167.875 ;
        RECT 88.130 167.665 88.300 167.855 ;
        RECT 89.510 167.685 89.680 167.875 ;
        RECT 89.785 167.710 89.945 167.820 ;
        RECT 90.300 167.715 90.420 167.825 ;
        RECT 90.705 167.685 90.875 167.875 ;
        RECT 91.165 167.665 91.335 167.855 ;
        RECT 91.625 167.665 91.795 167.855 ;
        RECT 93.005 167.825 93.175 167.875 ;
        RECT 93.005 167.715 93.180 167.825 ;
        RECT 93.005 167.685 93.175 167.715 ;
        RECT 93.465 167.685 93.635 167.875 ;
        RECT 100.550 167.685 100.720 167.875 ;
        RECT 101.340 167.715 101.460 167.825 ;
        RECT 102.665 167.665 102.835 167.855 ;
        RECT 103.125 167.685 103.295 167.875 ;
        RECT 104.045 167.665 104.215 167.855 ;
        RECT 104.560 167.715 104.680 167.825 ;
        RECT 106.345 167.665 106.515 167.855 ;
        RECT 106.990 167.685 107.160 167.875 ;
        RECT 108.645 167.685 108.815 167.875 ;
        RECT 109.105 167.855 109.275 167.875 ;
        RECT 109.100 167.685 109.275 167.855 ;
        RECT 29.845 166.855 31.215 167.665 ;
        RECT 31.685 166.855 34.435 167.665 ;
        RECT 34.455 166.755 35.805 167.665 ;
        RECT 35.825 166.855 37.195 167.665 ;
        RECT 37.215 166.795 37.645 167.580 ;
        RECT 37.665 166.885 39.035 167.665 ;
        RECT 39.045 166.855 42.715 167.665 ;
        RECT 42.920 166.755 46.395 167.665 ;
        RECT 46.635 166.985 50.535 167.665 ;
        RECT 49.605 166.755 50.535 166.985 ;
        RECT 50.555 166.755 51.905 167.665 ;
        RECT 52.120 166.755 55.595 167.665 ;
        RECT 55.605 166.985 59.505 167.665 ;
        RECT 55.605 166.755 56.535 166.985 ;
        RECT 60.205 166.855 62.955 167.665 ;
        RECT 62.975 166.795 63.405 167.580 ;
        RECT 63.425 166.855 65.255 167.665 ;
        RECT 65.265 166.985 69.165 167.665 ;
        RECT 69.635 166.985 73.535 167.665 ;
        RECT 65.265 166.755 66.195 166.985 ;
        RECT 72.605 166.755 73.535 166.985 ;
        RECT 74.145 166.755 76.755 167.665 ;
        RECT 77.225 166.985 79.055 167.665 ;
        RECT 77.225 166.755 78.570 166.985 ;
        RECT 79.065 166.855 80.895 167.665 ;
        RECT 80.905 166.755 84.380 167.665 ;
        RECT 84.815 166.985 88.715 167.665 ;
        RECT 87.785 166.755 88.715 166.985 ;
        RECT 88.735 166.795 89.165 167.580 ;
        RECT 90.115 166.755 91.465 167.665 ;
        RECT 91.485 166.885 92.855 167.665 ;
        RECT 93.695 166.985 102.975 167.665 ;
        RECT 93.695 166.865 96.030 166.985 ;
        RECT 93.695 166.755 94.615 166.865 ;
        RECT 100.695 166.765 101.615 166.985 ;
        RECT 102.985 166.885 104.355 167.665 ;
        RECT 104.825 166.855 106.655 167.665 ;
        RECT 106.665 167.635 107.610 167.665 ;
        RECT 109.100 167.635 109.270 167.685 ;
        RECT 109.570 167.665 109.740 167.855 ;
        RECT 113.890 167.685 114.060 167.875 ;
        RECT 114.165 167.665 114.335 167.855 ;
        RECT 114.680 167.715 114.800 167.825 ;
        RECT 115.085 167.665 115.255 167.855 ;
        RECT 116.465 167.685 116.635 167.875 ;
        RECT 121.060 167.665 121.230 167.855 ;
        RECT 123.820 167.665 123.990 167.855 ;
        RECT 124.340 167.715 124.460 167.825 ;
        RECT 125.665 167.685 125.835 167.875 ;
        RECT 126.125 167.825 126.295 167.855 ;
        RECT 126.125 167.715 126.300 167.825 ;
        RECT 126.125 167.665 126.295 167.715 ;
        RECT 127.505 167.665 127.675 167.875 ;
        RECT 106.665 166.955 109.415 167.635 ;
        RECT 106.665 166.755 107.610 166.955 ;
        RECT 109.425 166.755 112.900 167.665 ;
        RECT 113.105 166.855 114.475 167.665 ;
        RECT 114.495 166.795 114.925 167.580 ;
        RECT 115.055 166.985 118.520 167.665 ;
        RECT 117.600 166.755 118.520 166.985 ;
        RECT 118.765 166.755 121.375 167.665 ;
        RECT 121.525 166.755 124.135 167.665 ;
        RECT 124.605 166.855 126.435 167.665 ;
        RECT 126.445 166.855 127.815 167.665 ;
      LAYER nwell ;
        RECT 29.650 163.635 128.010 166.465 ;
      LAYER pwell ;
        RECT 29.845 162.435 31.215 163.245 ;
        RECT 35.345 163.115 36.275 163.345 ;
        RECT 39.485 163.115 40.415 163.345 ;
        RECT 32.375 162.435 36.275 163.115 ;
        RECT 36.515 162.435 40.415 163.115 ;
        RECT 40.795 163.235 41.715 163.345 ;
        RECT 40.795 163.115 43.130 163.235 ;
        RECT 47.795 163.115 48.715 163.335 ;
        RECT 40.795 162.435 50.075 163.115 ;
        RECT 50.095 162.520 50.525 163.305 ;
        RECT 50.915 163.235 51.835 163.345 ;
        RECT 50.915 163.115 53.250 163.235 ;
        RECT 57.915 163.115 58.835 163.335 ;
        RECT 62.860 163.115 63.780 163.345 ;
        RECT 50.915 162.435 60.195 163.115 ;
        RECT 60.315 162.435 63.780 163.115 ;
        RECT 63.885 162.435 67.360 163.345 ;
        RECT 67.565 162.435 71.040 163.345 ;
        RECT 71.245 162.435 72.615 163.245 ;
        RECT 72.625 162.435 73.995 163.215 ;
        RECT 74.005 163.115 75.350 163.345 ;
        RECT 74.005 162.435 75.835 163.115 ;
        RECT 75.855 162.520 76.285 163.305 ;
        RECT 76.765 163.115 78.110 163.345 ;
        RECT 79.090 163.115 80.435 163.345 ;
        RECT 76.765 162.435 78.595 163.115 ;
        RECT 78.605 162.435 80.435 163.115 ;
        RECT 80.445 162.435 81.815 163.245 ;
        RECT 81.825 162.435 85.300 163.345 ;
        RECT 85.875 163.235 86.795 163.345 ;
        RECT 85.875 163.115 88.210 163.235 ;
        RECT 92.875 163.115 93.795 163.335 ;
        RECT 85.875 162.435 95.155 163.115 ;
        RECT 95.165 162.435 96.535 163.245 ;
        RECT 96.555 162.435 97.905 163.345 ;
        RECT 98.120 162.435 101.595 163.345 ;
        RECT 101.615 162.520 102.045 163.305 ;
        RECT 102.065 162.435 103.895 163.245 ;
        RECT 104.100 162.435 107.575 163.345 ;
        RECT 107.585 162.435 111.060 163.345 ;
        RECT 111.265 162.435 114.740 163.345 ;
        RECT 115.140 162.435 118.615 163.345 ;
        RECT 119.085 162.435 120.915 163.245 ;
        RECT 120.925 162.435 126.435 163.245 ;
        RECT 126.445 162.435 127.815 163.245 ;
        RECT 29.985 162.225 30.155 162.435 ;
        RECT 31.825 162.270 31.985 162.390 ;
        RECT 35.505 162.225 35.675 162.415 ;
        RECT 35.690 162.245 35.860 162.435 ;
        RECT 36.885 162.225 37.055 162.415 ;
        RECT 39.830 162.245 40.000 162.435 ;
        RECT 40.105 162.225 40.275 162.415 ;
        RECT 41.485 162.225 41.655 162.415 ;
        RECT 41.945 162.225 42.115 162.415 ;
        RECT 46.540 162.225 46.710 162.415 ;
        RECT 49.765 162.245 49.935 162.435 ;
        RECT 50.220 162.225 50.390 162.415 ;
        RECT 51.605 162.225 51.775 162.415 ;
        RECT 52.120 162.275 52.240 162.385 ;
        RECT 53.905 162.225 54.075 162.415 ;
        RECT 54.365 162.225 54.535 162.415 ;
        RECT 55.750 162.225 55.920 162.415 ;
        RECT 59.430 162.225 59.600 162.415 ;
        RECT 59.885 162.245 60.055 162.435 ;
        RECT 60.345 162.245 60.515 162.435 ;
        RECT 63.620 162.275 63.740 162.385 ;
        RECT 64.030 162.245 64.200 162.435 ;
        RECT 67.710 162.415 67.880 162.435 ;
        RECT 66.325 162.225 66.495 162.415 ;
        RECT 67.705 162.245 67.880 162.415 ;
        RECT 67.705 162.225 67.875 162.245 ;
        RECT 68.165 162.225 68.335 162.415 ;
        RECT 70.925 162.225 71.095 162.415 ;
        RECT 72.305 162.245 72.475 162.435 ;
        RECT 72.765 162.225 72.935 162.435 ;
        RECT 75.525 162.245 75.695 162.435 ;
        RECT 76.500 162.275 76.620 162.385 ;
        RECT 78.285 162.245 78.455 162.435 ;
        RECT 78.745 162.245 78.915 162.435 ;
        RECT 81.505 162.245 81.675 162.435 ;
        RECT 81.970 162.415 82.140 162.435 ;
        RECT 81.965 162.245 82.140 162.415 ;
        RECT 82.480 162.275 82.600 162.385 ;
        RECT 81.965 162.225 82.135 162.245 ;
        RECT 82.890 162.225 83.060 162.415 ;
        RECT 86.620 162.275 86.740 162.385 ;
        RECT 88.405 162.225 88.575 162.415 ;
        RECT 91.625 162.225 91.795 162.415 ;
        RECT 93.005 162.225 93.175 162.415 ;
        RECT 93.520 162.275 93.640 162.385 ;
        RECT 94.845 162.245 95.015 162.435 ;
        RECT 96.225 162.225 96.395 162.435 ;
        RECT 96.685 162.245 96.855 162.435 ;
        RECT 101.280 162.245 101.450 162.435 ;
        RECT 103.585 162.245 103.755 162.435 ;
        RECT 107.260 162.415 107.430 162.435 ;
        RECT 105.425 162.225 105.595 162.415 ;
        RECT 106.805 162.225 106.975 162.415 ;
        RECT 107.260 162.245 107.440 162.415 ;
        RECT 107.730 162.245 107.900 162.435 ;
        RECT 107.270 162.225 107.440 162.245 ;
        RECT 110.945 162.225 111.115 162.415 ;
        RECT 111.410 162.245 111.580 162.435 ;
        RECT 115.545 162.270 115.705 162.380 ;
        RECT 116.005 162.225 116.175 162.415 ;
        RECT 118.300 162.245 118.470 162.435 ;
        RECT 118.820 162.275 118.940 162.385 ;
        RECT 120.605 162.245 120.775 162.435 ;
        RECT 126.125 162.225 126.295 162.435 ;
        RECT 127.505 162.225 127.675 162.435 ;
        RECT 29.845 161.415 31.215 162.225 ;
        RECT 32.145 161.415 35.815 162.225 ;
        RECT 35.835 161.315 37.185 162.225 ;
        RECT 37.215 161.355 37.645 162.140 ;
        RECT 37.665 161.415 40.415 162.225 ;
        RECT 40.425 161.445 41.795 162.225 ;
        RECT 41.815 161.315 43.165 162.225 ;
        RECT 43.380 161.315 46.855 162.225 ;
        RECT 47.060 161.315 50.535 162.225 ;
        RECT 50.545 161.445 51.915 162.225 ;
        RECT 52.385 161.415 54.215 162.225 ;
        RECT 54.225 161.445 55.595 162.225 ;
        RECT 55.605 161.315 59.080 162.225 ;
        RECT 59.285 161.315 62.760 162.225 ;
        RECT 62.975 161.355 63.405 162.140 ;
        RECT 63.885 161.415 66.635 162.225 ;
        RECT 66.655 161.315 68.005 162.225 ;
        RECT 68.025 161.445 69.395 162.225 ;
        RECT 69.405 161.415 71.235 162.225 ;
        RECT 71.245 161.545 73.075 162.225 ;
        RECT 73.170 161.545 82.275 162.225 ;
        RECT 71.245 161.315 72.590 161.545 ;
        RECT 82.745 161.315 86.220 162.225 ;
        RECT 86.885 161.415 88.715 162.225 ;
        RECT 88.735 161.355 89.165 162.140 ;
        RECT 89.185 161.415 91.935 162.225 ;
        RECT 91.955 161.315 93.305 162.225 ;
        RECT 93.785 161.415 96.535 162.225 ;
        RECT 96.545 161.545 105.735 162.225 ;
        RECT 96.545 161.315 97.465 161.545 ;
        RECT 100.295 161.325 101.225 161.545 ;
        RECT 105.745 161.415 107.115 162.225 ;
        RECT 107.125 161.315 110.600 162.225 ;
        RECT 110.915 161.545 114.380 162.225 ;
        RECT 113.460 161.315 114.380 161.545 ;
        RECT 114.495 161.355 114.925 162.140 ;
        RECT 115.875 161.315 117.225 162.225 ;
        RECT 117.245 161.545 126.435 162.225 ;
        RECT 117.245 161.315 118.165 161.545 ;
        RECT 120.995 161.325 121.925 161.545 ;
        RECT 126.445 161.415 127.815 162.225 ;
      LAYER nwell ;
        RECT 29.650 158.195 128.010 161.025 ;
      LAYER pwell ;
        RECT 29.845 156.995 31.215 157.805 ;
        RECT 32.515 157.795 33.435 157.905 ;
        RECT 32.515 157.675 34.850 157.795 ;
        RECT 39.515 157.675 40.435 157.895 ;
        RECT 32.515 156.995 41.795 157.675 ;
        RECT 41.805 156.995 44.555 157.805 ;
        RECT 44.565 156.995 50.075 157.805 ;
        RECT 50.095 157.080 50.525 157.865 ;
        RECT 51.005 156.995 52.835 157.805 ;
        RECT 52.845 157.705 53.790 157.905 ;
        RECT 52.845 157.025 55.595 157.705 ;
        RECT 52.845 156.995 53.790 157.025 ;
        RECT 29.985 156.785 30.155 156.995 ;
        RECT 31.825 156.840 31.985 156.950 ;
        RECT 33.665 156.785 33.835 156.975 ;
        RECT 34.125 156.785 34.295 156.975 ;
        RECT 36.885 156.785 37.055 156.975 ;
        RECT 37.805 156.785 37.975 156.975 ;
        RECT 39.645 156.830 39.805 156.940 ;
        RECT 41.485 156.805 41.655 156.995 ;
        RECT 44.245 156.805 44.415 156.995 ;
        RECT 45.165 156.785 45.335 156.975 ;
        RECT 29.845 155.975 31.215 156.785 ;
        RECT 31.225 155.975 33.975 156.785 ;
        RECT 33.995 155.875 35.345 156.785 ;
        RECT 35.365 155.975 37.195 156.785 ;
        RECT 37.215 155.915 37.645 156.700 ;
        RECT 37.665 156.005 39.035 156.785 ;
        RECT 39.965 155.975 45.475 156.785 ;
        RECT 45.485 156.755 46.430 156.785 ;
        RECT 47.920 156.755 48.090 156.975 ;
        RECT 48.390 156.785 48.560 156.975 ;
        RECT 49.765 156.805 49.935 156.995 ;
        RECT 50.740 156.835 50.860 156.945 ;
        RECT 52.525 156.805 52.695 156.995 ;
        RECT 55.280 156.805 55.450 157.025 ;
        RECT 55.605 156.995 59.275 157.805 ;
        RECT 59.285 156.995 62.760 157.905 ;
        RECT 63.335 157.795 64.255 157.905 ;
        RECT 63.335 157.675 65.670 157.795 ;
        RECT 70.335 157.675 71.255 157.895 ;
        RECT 63.335 156.995 72.615 157.675 ;
        RECT 73.085 156.995 75.835 157.805 ;
        RECT 75.855 157.080 76.285 157.865 ;
        RECT 76.305 157.675 77.650 157.905 ;
        RECT 78.630 157.675 79.975 157.905 ;
        RECT 76.305 156.995 78.135 157.675 ;
        RECT 78.145 156.995 79.975 157.675 ;
        RECT 79.985 156.995 82.705 157.905 ;
        RECT 82.745 157.705 83.690 157.905 ;
        RECT 82.745 157.025 85.495 157.705 ;
        RECT 82.745 156.995 83.690 157.025 ;
        RECT 58.965 156.805 59.135 156.995 ;
        RECT 59.430 156.805 59.600 156.995 ;
        RECT 61.265 156.785 61.435 156.975 ;
        RECT 62.645 156.785 62.815 156.975 ;
        RECT 66.970 156.785 67.140 156.975 ;
        RECT 68.165 156.830 68.325 156.940 ;
        RECT 72.030 156.785 72.200 156.975 ;
        RECT 72.305 156.805 72.475 156.995 ;
        RECT 72.820 156.835 72.940 156.945 ;
        RECT 73.685 156.785 73.855 156.975 ;
        RECT 74.605 156.830 74.765 156.940 ;
        RECT 75.525 156.805 75.695 156.995 ;
        RECT 77.365 156.785 77.535 156.975 ;
        RECT 77.825 156.945 77.995 156.995 ;
        RECT 77.825 156.835 78.000 156.945 ;
        RECT 77.825 156.805 77.995 156.835 ;
        RECT 78.285 156.785 78.455 156.995 ;
        RECT 80.125 156.805 80.295 156.995 ;
        RECT 84.260 156.785 84.430 156.975 ;
        RECT 85.180 156.805 85.350 157.025 ;
        RECT 85.965 156.995 87.795 157.805 ;
        RECT 88.175 157.795 89.095 157.905 ;
        RECT 88.175 157.675 90.510 157.795 ;
        RECT 95.175 157.675 96.095 157.895 ;
        RECT 88.175 156.995 97.455 157.675 ;
        RECT 97.465 156.995 99.295 157.805 ;
        RECT 99.315 156.995 100.665 157.905 ;
        RECT 101.615 157.080 102.045 157.865 ;
        RECT 102.065 156.995 105.735 157.805 ;
        RECT 105.745 157.705 106.690 157.905 ;
        RECT 105.745 157.025 108.495 157.705 ;
        RECT 105.745 156.995 106.690 157.025 ;
        RECT 85.700 156.835 85.820 156.945 ;
        RECT 87.485 156.805 87.655 156.995 ;
        RECT 88.130 156.785 88.300 156.975 ;
        RECT 90.245 156.785 90.415 156.975 ;
        RECT 91.625 156.785 91.795 156.975 ;
        RECT 92.140 156.835 92.260 156.945 ;
        RECT 92.545 156.785 92.715 156.975 ;
        RECT 93.925 156.785 94.095 156.975 ;
        RECT 97.145 156.805 97.315 156.995 ;
        RECT 98.985 156.805 99.155 156.995 ;
        RECT 100.365 156.805 100.535 156.995 ;
        RECT 101.010 156.785 101.180 156.975 ;
        RECT 101.285 156.840 101.445 156.950 ;
        RECT 101.745 156.785 101.915 156.975 ;
        RECT 104.045 156.785 104.215 156.975 ;
        RECT 105.425 156.805 105.595 156.995 ;
        RECT 108.180 156.975 108.350 157.025 ;
        RECT 108.505 156.995 111.980 157.905 ;
        RECT 113.105 157.675 114.035 157.905 ;
        RECT 120.445 157.675 121.375 157.905 ;
        RECT 113.105 156.995 117.005 157.675 ;
        RECT 117.475 156.995 121.375 157.675 ;
        RECT 122.305 156.995 123.675 157.775 ;
        RECT 123.685 156.995 125.055 157.775 ;
        RECT 125.065 156.995 126.435 157.805 ;
        RECT 126.445 156.995 127.815 157.805 ;
        RECT 107.725 156.785 107.895 156.975 ;
        RECT 108.180 156.805 108.360 156.975 ;
        RECT 108.650 156.805 108.820 156.995 ;
        RECT 45.485 156.075 48.235 156.755 ;
        RECT 45.485 155.875 46.430 156.075 ;
        RECT 48.245 155.875 51.720 156.785 ;
        RECT 52.295 156.105 61.575 156.785 ;
        RECT 52.295 155.985 54.630 156.105 ;
        RECT 52.295 155.875 53.215 155.985 ;
        RECT 59.295 155.885 60.215 156.105 ;
        RECT 61.595 155.875 62.945 156.785 ;
        RECT 62.975 155.915 63.405 156.700 ;
        RECT 63.655 156.105 67.555 156.785 ;
        RECT 68.715 156.105 72.615 156.785 ;
        RECT 66.625 155.875 67.555 156.105 ;
        RECT 71.685 155.875 72.615 156.105 ;
        RECT 72.635 155.875 73.985 156.785 ;
        RECT 74.935 156.105 77.675 156.785 ;
        RECT 78.145 156.105 80.885 156.785 ;
        RECT 81.100 155.875 84.575 156.785 ;
        RECT 84.815 156.105 88.715 156.785 ;
        RECT 87.785 155.875 88.715 156.105 ;
        RECT 88.735 155.915 89.165 156.700 ;
        RECT 89.185 155.975 90.555 156.785 ;
        RECT 90.575 155.875 91.925 156.785 ;
        RECT 92.405 156.005 93.775 156.785 ;
        RECT 93.895 156.105 97.360 156.785 ;
        RECT 97.695 156.105 101.595 156.785 ;
        RECT 96.440 155.875 97.360 156.105 ;
        RECT 100.665 155.875 101.595 156.105 ;
        RECT 101.605 156.005 102.975 156.785 ;
        RECT 102.985 155.975 104.355 156.785 ;
        RECT 104.365 155.975 108.035 156.785 ;
        RECT 108.190 156.755 108.360 156.805 ;
        RECT 110.945 156.785 111.115 156.975 ;
        RECT 112.785 156.840 112.945 156.950 ;
        RECT 113.520 156.805 113.690 156.995 ;
        RECT 115.140 156.835 115.260 156.945 ;
        RECT 115.545 156.785 115.715 156.975 ;
        RECT 120.790 156.805 120.960 156.995 ;
        RECT 121.985 156.840 122.145 156.950 ;
        RECT 122.445 156.805 122.615 156.995 ;
        RECT 123.825 156.805 123.995 156.995 ;
        RECT 126.125 156.785 126.295 156.995 ;
        RECT 127.505 156.785 127.675 156.995 ;
        RECT 109.850 156.755 110.795 156.785 ;
        RECT 108.045 156.075 110.795 156.755 ;
        RECT 110.915 156.105 114.380 156.785 ;
        RECT 109.850 155.875 110.795 156.075 ;
        RECT 113.460 155.875 114.380 156.105 ;
        RECT 114.495 155.915 114.925 156.700 ;
        RECT 115.415 155.875 116.765 156.785 ;
        RECT 117.155 156.105 126.435 156.785 ;
        RECT 117.155 155.985 119.490 156.105 ;
        RECT 117.155 155.875 118.075 155.985 ;
        RECT 124.155 155.885 125.075 156.105 ;
        RECT 126.445 155.975 127.815 156.785 ;
      LAYER nwell ;
        RECT 29.650 152.755 128.010 155.585 ;
      LAYER pwell ;
        RECT 29.845 151.555 31.215 152.365 ;
        RECT 31.595 152.355 32.515 152.465 ;
        RECT 31.595 152.235 33.930 152.355 ;
        RECT 38.595 152.235 39.515 152.455 ;
        RECT 31.595 151.555 40.875 152.235 ;
        RECT 41.345 151.555 43.175 152.365 ;
        RECT 43.185 151.555 44.555 152.335 ;
        RECT 44.565 152.265 45.510 152.465 ;
        RECT 49.130 152.265 50.075 152.465 ;
        RECT 44.565 151.585 47.315 152.265 ;
        RECT 47.325 151.585 50.075 152.265 ;
        RECT 50.095 151.640 50.525 152.425 ;
        RECT 51.685 152.375 52.635 152.465 ;
        RECT 44.565 151.555 45.510 151.585 ;
        RECT 29.985 151.345 30.155 151.555 ;
        RECT 31.420 151.395 31.540 151.505 ;
        RECT 32.745 151.345 32.915 151.535 ;
        RECT 36.610 151.345 36.780 151.535 ;
        RECT 40.565 151.365 40.735 151.555 ;
        RECT 41.080 151.395 41.200 151.505 ;
        RECT 42.865 151.365 43.035 151.555 ;
        RECT 43.325 151.365 43.495 151.555 ;
        RECT 47.000 151.535 47.170 151.585 ;
        RECT 47.000 151.365 47.175 151.535 ;
        RECT 47.470 151.365 47.640 151.585 ;
        RECT 49.130 151.555 50.075 151.585 ;
        RECT 50.705 151.555 52.635 152.375 ;
        RECT 52.845 151.555 56.320 152.465 ;
        RECT 56.895 152.355 57.815 152.465 ;
        RECT 56.895 152.235 59.230 152.355 ;
        RECT 63.895 152.235 64.815 152.455 ;
        RECT 66.645 152.235 67.565 152.465 ;
        RECT 70.395 152.235 71.325 152.455 ;
        RECT 56.895 151.555 66.175 152.235 ;
        RECT 66.645 151.555 75.835 152.235 ;
        RECT 75.855 151.640 76.285 152.425 ;
        RECT 76.305 151.555 77.675 152.335 ;
        RECT 78.170 152.235 79.515 152.465 ;
        RECT 81.330 152.265 82.275 152.465 ;
        RECT 77.685 151.555 79.515 152.235 ;
        RECT 79.525 151.585 82.275 152.265 ;
        RECT 50.705 151.535 50.855 151.555 ;
        RECT 49.305 151.365 49.475 151.535 ;
        RECT 50.685 151.365 50.855 151.535 ;
        RECT 51.605 151.365 51.775 151.535 ;
        RECT 52.525 151.390 52.685 151.500 ;
        RECT 47.005 151.345 47.175 151.365 ;
        RECT 49.305 151.345 49.455 151.365 ;
        RECT 51.605 151.345 51.755 151.365 ;
        RECT 52.990 151.345 53.160 151.555 ;
        RECT 57.125 151.390 57.285 151.500 ;
        RECT 60.990 151.345 61.160 151.535 ;
        RECT 62.645 151.345 62.815 151.535 ;
        RECT 64.485 151.345 64.655 151.535 ;
        RECT 64.950 151.345 65.120 151.535 ;
        RECT 65.865 151.365 66.035 151.555 ;
        RECT 66.380 151.395 66.500 151.505 ;
        RECT 68.625 151.345 68.795 151.535 ;
        RECT 75.525 151.365 75.695 151.555 ;
        RECT 77.365 151.365 77.535 151.555 ;
        RECT 77.825 151.365 77.995 151.555 ;
        RECT 79.205 151.345 79.375 151.535 ;
        RECT 79.670 151.365 79.840 151.585 ;
        RECT 81.330 151.555 82.275 151.585 ;
        RECT 82.285 151.555 85.760 152.465 ;
        RECT 86.335 152.355 87.255 152.465 ;
        RECT 86.335 152.235 88.670 152.355 ;
        RECT 93.335 152.235 94.255 152.455 ;
        RECT 86.335 151.555 95.615 152.235 ;
        RECT 96.085 151.555 97.915 152.365 ;
        RECT 97.925 151.555 101.400 152.465 ;
        RECT 101.615 151.640 102.045 152.425 ;
        RECT 102.065 151.555 107.575 152.365 ;
        RECT 107.585 151.555 111.060 152.465 ;
        RECT 111.460 151.555 114.935 152.465 ;
        RECT 115.405 151.555 117.235 152.365 ;
        RECT 120.445 152.235 121.375 152.465 ;
        RECT 117.475 151.555 121.375 152.235 ;
        RECT 121.385 151.555 122.755 152.365 ;
        RECT 122.765 151.555 126.435 152.365 ;
        RECT 126.445 151.555 127.815 152.365 ;
        RECT 80.585 151.345 80.755 151.535 ;
        RECT 82.430 151.365 82.600 151.555 ;
        RECT 84.265 151.345 84.435 151.535 ;
        RECT 88.130 151.345 88.300 151.535 ;
        RECT 89.380 151.395 89.500 151.505 ;
        RECT 91.165 151.345 91.335 151.535 ;
        RECT 91.625 151.345 91.795 151.535 ;
        RECT 93.060 151.395 93.180 151.505 ;
        RECT 95.305 151.365 95.475 151.555 ;
        RECT 95.820 151.395 95.940 151.505 ;
        RECT 96.685 151.345 96.855 151.535 ;
        RECT 97.605 151.365 97.775 151.555 ;
        RECT 98.070 151.365 98.240 151.555 ;
        RECT 106.345 151.345 106.515 151.535 ;
        RECT 107.265 151.365 107.435 151.555 ;
        RECT 107.730 151.535 107.900 151.555 ;
        RECT 107.725 151.365 107.900 151.535 ;
        RECT 107.725 151.345 107.895 151.365 ;
        RECT 108.190 151.345 108.360 151.535 ;
        RECT 112.785 151.345 112.955 151.535 ;
        RECT 113.245 151.345 113.415 151.535 ;
        RECT 114.620 151.365 114.790 151.555 ;
        RECT 115.140 151.395 115.260 151.505 ;
        RECT 115.545 151.345 115.715 151.535 ;
        RECT 116.925 151.365 117.095 151.555 ;
        RECT 120.790 151.365 120.960 151.555 ;
        RECT 122.445 151.365 122.615 151.555 ;
        RECT 126.125 151.345 126.295 151.555 ;
        RECT 127.505 151.345 127.675 151.555 ;
        RECT 29.845 150.535 31.215 151.345 ;
        RECT 31.695 150.435 33.045 151.345 ;
        RECT 33.295 150.665 37.195 151.345 ;
        RECT 36.265 150.435 37.195 150.665 ;
        RECT 37.215 150.475 37.645 151.260 ;
        RECT 38.035 150.665 47.315 151.345 ;
        RECT 38.035 150.545 40.370 150.665 ;
        RECT 38.035 150.435 38.955 150.545 ;
        RECT 45.035 150.445 45.955 150.665 ;
        RECT 47.525 150.525 49.455 151.345 ;
        RECT 49.825 150.525 51.755 151.345 ;
        RECT 47.525 150.435 48.475 150.525 ;
        RECT 49.825 150.435 50.775 150.525 ;
        RECT 52.845 150.435 56.320 151.345 ;
        RECT 57.675 150.665 61.575 151.345 ;
        RECT 60.645 150.435 61.575 150.665 ;
        RECT 61.585 150.565 62.955 151.345 ;
        RECT 62.975 150.475 63.405 151.260 ;
        RECT 63.425 150.535 64.795 151.345 ;
        RECT 64.805 150.435 68.280 151.345 ;
        RECT 68.495 150.435 69.845 151.345 ;
        RECT 70.235 150.665 79.515 151.345 ;
        RECT 70.235 150.545 72.570 150.665 ;
        RECT 70.235 150.435 71.155 150.545 ;
        RECT 77.235 150.445 78.155 150.665 ;
        RECT 79.525 150.565 80.895 151.345 ;
        RECT 80.905 150.535 84.575 151.345 ;
        RECT 84.815 150.665 88.715 151.345 ;
        RECT 87.785 150.435 88.715 150.665 ;
        RECT 88.735 150.475 89.165 151.260 ;
        RECT 89.645 150.535 91.475 151.345 ;
        RECT 91.485 150.565 92.855 151.345 ;
        RECT 93.325 150.535 96.995 151.345 ;
        RECT 97.375 150.665 106.655 151.345 ;
        RECT 97.375 150.545 99.710 150.665 ;
        RECT 97.375 150.435 98.295 150.545 ;
        RECT 104.375 150.445 105.295 150.665 ;
        RECT 106.665 150.535 108.035 151.345 ;
        RECT 108.045 150.435 111.520 151.345 ;
        RECT 111.725 150.535 113.095 151.345 ;
        RECT 113.115 150.435 114.465 151.345 ;
        RECT 114.495 150.475 114.925 151.260 ;
        RECT 115.415 150.435 116.765 151.345 ;
        RECT 117.155 150.665 126.435 151.345 ;
        RECT 117.155 150.545 119.490 150.665 ;
        RECT 117.155 150.435 118.075 150.545 ;
        RECT 124.155 150.445 125.075 150.665 ;
        RECT 126.445 150.535 127.815 151.345 ;
      LAYER nwell ;
        RECT 29.650 147.315 128.010 150.145 ;
      LAYER pwell ;
        RECT 29.845 146.115 31.215 146.925 ;
        RECT 31.595 146.915 32.515 147.025 ;
        RECT 31.595 146.795 33.930 146.915 ;
        RECT 38.595 146.795 39.515 147.015 ;
        RECT 31.595 146.115 40.875 146.795 ;
        RECT 40.885 146.115 42.715 146.925 ;
        RECT 42.725 146.795 43.655 147.025 ;
        RECT 47.065 146.935 48.015 147.025 ;
        RECT 42.725 146.115 46.625 146.795 ;
        RECT 47.065 146.115 48.995 146.935 ;
        RECT 50.095 146.200 50.525 146.985 ;
        RECT 51.015 146.115 52.365 147.025 ;
        RECT 52.385 146.825 53.330 147.025 ;
        RECT 52.385 146.145 55.135 146.825 ;
        RECT 61.020 146.795 61.940 147.025 ;
        RECT 52.385 146.115 53.330 146.145 ;
        RECT 29.985 145.905 30.155 146.115 ;
        RECT 31.420 145.955 31.540 146.065 ;
        RECT 32.745 145.905 32.915 146.095 ;
        RECT 36.610 145.905 36.780 146.095 ;
        RECT 37.805 145.905 37.975 146.095 ;
        RECT 40.565 145.925 40.735 146.115 ;
        RECT 42.405 145.905 42.575 146.115 ;
        RECT 43.140 145.925 43.310 146.115 ;
        RECT 48.845 146.095 48.995 146.115 ;
        RECT 47.925 145.905 48.095 146.095 ;
        RECT 48.845 145.925 49.015 146.095 ;
        RECT 49.765 145.960 49.925 146.070 ;
        RECT 50.740 145.955 50.860 146.065 ;
        RECT 52.065 145.925 52.235 146.115 ;
        RECT 53.445 145.905 53.615 146.095 ;
        RECT 54.820 145.925 54.990 146.145 ;
        RECT 55.525 146.115 57.950 146.795 ;
        RECT 58.475 146.115 61.940 146.795 ;
        RECT 62.045 146.115 64.795 146.925 ;
        RECT 67.460 146.795 68.380 147.025 ;
        RECT 64.915 146.115 68.380 146.795 ;
        RECT 68.945 146.115 70.775 146.925 ;
        RECT 73.985 146.795 74.915 147.025 ;
        RECT 71.015 146.115 74.915 146.795 ;
        RECT 75.855 146.200 76.285 146.985 ;
        RECT 77.225 146.115 80.895 146.925 ;
        RECT 80.905 146.115 86.415 146.925 ;
        RECT 86.795 146.915 87.715 147.025 ;
        RECT 86.795 146.795 89.130 146.915 ;
        RECT 93.795 146.795 94.715 147.015 ;
        RECT 86.795 146.115 96.075 146.795 ;
        RECT 96.085 146.115 97.455 146.925 ;
        RECT 97.475 146.115 98.825 147.025 ;
        RECT 100.650 146.825 101.595 147.025 ;
        RECT 98.845 146.145 101.595 146.825 ;
        RECT 101.615 146.200 102.045 146.985 ;
        RECT 106.185 146.795 107.115 147.025 ;
        RECT 108.930 146.825 109.875 147.025 ;
        RECT 58.045 145.925 58.215 146.095 ;
        RECT 58.505 145.925 58.675 146.115 ;
        RECT 62.645 145.905 62.815 146.095 ;
        RECT 63.620 145.955 63.740 146.065 ;
        RECT 64.485 145.925 64.655 146.115 ;
        RECT 64.945 145.925 65.115 146.115 ;
        RECT 66.785 145.905 66.955 146.095 ;
        RECT 67.250 145.905 67.420 146.095 ;
        RECT 68.680 145.955 68.800 146.065 ;
        RECT 70.465 145.925 70.635 146.115 ;
        RECT 70.980 145.955 71.100 146.065 ;
        RECT 74.330 145.925 74.500 146.115 ;
        RECT 80.585 146.095 80.755 146.115 ;
        RECT 74.605 145.905 74.775 146.095 ;
        RECT 75.065 145.905 75.235 146.095 ;
        RECT 75.525 145.960 75.685 146.070 ;
        RECT 76.905 145.960 77.065 146.070 ;
        RECT 77.825 145.905 77.995 146.095 ;
        RECT 80.580 145.925 80.755 146.095 ;
        RECT 29.845 145.095 31.215 145.905 ;
        RECT 31.695 144.995 33.045 145.905 ;
        RECT 33.295 145.225 37.195 145.905 ;
        RECT 36.265 144.995 37.195 145.225 ;
        RECT 37.215 145.035 37.645 145.820 ;
        RECT 37.665 145.125 39.035 145.905 ;
        RECT 39.045 145.095 42.715 145.905 ;
        RECT 42.725 145.095 48.235 145.905 ;
        RECT 48.245 145.095 53.755 145.905 ;
        RECT 53.850 145.225 62.955 145.905 ;
        RECT 62.975 145.035 63.405 145.820 ;
        RECT 63.885 144.995 67.095 145.905 ;
        RECT 67.105 144.995 70.580 145.905 ;
        RECT 71.245 145.095 74.915 145.905 ;
        RECT 74.925 145.125 76.295 145.905 ;
        RECT 76.305 145.225 78.135 145.905 ;
        RECT 78.145 145.875 79.090 145.905 ;
        RECT 80.580 145.875 80.750 145.925 ;
        RECT 81.050 145.905 81.220 146.095 ;
        RECT 86.105 145.925 86.275 146.115 ;
        RECT 88.130 145.905 88.300 146.095 ;
        RECT 92.730 145.905 92.900 146.095 ;
        RECT 93.465 145.905 93.635 146.095 ;
        RECT 95.765 145.925 95.935 146.115 ;
        RECT 97.145 145.925 97.315 146.115 ;
        RECT 97.605 145.925 97.775 146.115 ;
        RECT 98.990 145.925 99.160 146.145 ;
        RECT 100.650 146.115 101.595 146.145 ;
        RECT 103.215 146.115 107.115 146.795 ;
        RECT 107.125 146.145 109.875 146.825 ;
        RECT 102.665 146.065 102.825 146.070 ;
        RECT 102.665 145.960 102.840 146.065 ;
        RECT 102.720 145.955 102.840 145.960 ;
        RECT 104.505 145.905 104.675 146.095 ;
        RECT 105.885 145.905 106.055 146.095 ;
        RECT 106.530 145.925 106.700 146.115 ;
        RECT 107.270 145.925 107.440 146.145 ;
        RECT 108.930 146.115 109.875 146.145 ;
        RECT 109.885 146.825 110.830 147.025 ;
        RECT 113.935 146.915 114.855 147.025 ;
        RECT 109.885 146.145 112.635 146.825 ;
        RECT 113.935 146.795 116.270 146.915 ;
        RECT 120.935 146.795 121.855 147.015 ;
        RECT 109.885 146.115 110.830 146.145 ;
        RECT 108.645 145.905 108.815 146.095 ;
        RECT 112.320 145.925 112.490 146.145 ;
        RECT 113.935 146.115 123.215 146.795 ;
        RECT 123.225 146.115 124.595 146.895 ;
        RECT 124.605 146.115 126.435 146.925 ;
        RECT 126.445 146.115 127.815 146.925 ;
        RECT 113.245 145.960 113.405 146.070 ;
        RECT 114.165 145.905 114.335 146.095 ;
        RECT 118.490 145.905 118.660 146.095 ;
        RECT 119.280 145.955 119.400 146.065 ;
        RECT 119.685 145.905 119.855 146.095 ;
        RECT 122.905 145.925 123.075 146.115 ;
        RECT 123.365 145.925 123.535 146.115 ;
        RECT 126.125 145.905 126.295 146.115 ;
        RECT 127.505 145.905 127.675 146.115 ;
        RECT 78.145 145.195 80.895 145.875 ;
        RECT 78.145 144.995 79.090 145.195 ;
        RECT 80.905 144.995 84.380 145.905 ;
        RECT 84.815 145.225 88.715 145.905 ;
        RECT 87.785 144.995 88.715 145.225 ;
        RECT 88.735 145.035 89.165 145.820 ;
        RECT 89.415 145.225 93.315 145.905 ;
        RECT 93.325 145.225 102.430 145.905 ;
        RECT 92.385 144.995 93.315 145.225 ;
        RECT 102.985 145.095 104.815 145.905 ;
        RECT 104.825 145.125 106.195 145.905 ;
        RECT 106.205 145.095 108.955 145.905 ;
        RECT 108.965 145.095 114.475 145.905 ;
        RECT 114.495 145.035 114.925 145.820 ;
        RECT 115.175 145.225 119.075 145.905 ;
        RECT 118.145 144.995 119.075 145.225 ;
        RECT 119.545 145.125 120.915 145.905 ;
        RECT 120.925 145.095 126.435 145.905 ;
        RECT 126.445 145.095 127.815 145.905 ;
      LAYER nwell ;
        RECT 29.650 141.875 128.010 144.705 ;
      LAYER pwell ;
        RECT 29.845 140.675 31.215 141.485 ;
        RECT 32.515 141.475 33.435 141.585 ;
        RECT 32.515 141.355 34.850 141.475 ;
        RECT 39.515 141.355 40.435 141.575 ;
        RECT 32.515 140.675 41.795 141.355 ;
        RECT 41.805 140.675 44.555 141.485 ;
        RECT 44.575 140.675 45.925 141.585 ;
        RECT 45.945 141.355 46.875 141.585 ;
        RECT 45.945 140.675 49.845 141.355 ;
        RECT 50.095 140.760 50.525 141.545 ;
        RECT 54.905 141.495 55.855 141.585 ;
        RECT 51.005 140.675 53.755 141.485 ;
        RECT 53.925 140.675 55.855 141.495 ;
        RECT 56.065 141.385 57.010 141.585 ;
        RECT 56.065 140.705 58.815 141.385 ;
        RECT 56.065 140.675 57.010 140.705 ;
        RECT 29.985 140.465 30.155 140.675 ;
        RECT 31.420 140.515 31.540 140.625 ;
        RECT 31.825 140.520 31.985 140.630 ;
        RECT 32.745 140.465 32.915 140.655 ;
        RECT 36.610 140.465 36.780 140.655 ;
        RECT 38.725 140.465 38.895 140.655 ;
        RECT 39.185 140.465 39.355 140.655 ;
        RECT 41.025 140.510 41.185 140.620 ;
        RECT 41.485 140.465 41.655 140.675 ;
        RECT 42.865 140.465 43.035 140.655 ;
        RECT 44.245 140.485 44.415 140.675 ;
        RECT 44.705 140.485 44.875 140.675 ;
        RECT 46.360 140.485 46.530 140.675 ;
        RECT 50.740 140.515 50.860 140.625 ;
        RECT 53.445 140.485 53.615 140.675 ;
        RECT 53.925 140.655 54.075 140.675 ;
        RECT 53.905 140.485 54.075 140.655 ;
        RECT 54.825 140.465 54.995 140.655 ;
        RECT 56.205 140.465 56.375 140.655 ;
        RECT 58.500 140.485 58.670 140.705 ;
        RECT 59.285 140.675 62.955 141.485 ;
        RECT 64.770 141.385 65.715 141.585 ;
        RECT 62.965 140.705 65.715 141.385 ;
        RECT 58.960 140.625 59.130 140.655 ;
        RECT 58.960 140.515 59.140 140.625 ;
        RECT 29.845 139.655 31.215 140.465 ;
        RECT 31.695 139.555 33.045 140.465 ;
        RECT 33.295 139.785 37.195 140.465 ;
        RECT 36.265 139.555 37.195 139.785 ;
        RECT 37.215 139.595 37.645 140.380 ;
        RECT 37.665 139.655 39.035 140.465 ;
        RECT 39.045 139.685 40.415 140.465 ;
        RECT 41.345 139.685 42.715 140.465 ;
        RECT 42.725 139.785 52.005 140.465 ;
        RECT 52.395 139.785 55.135 140.465 ;
        RECT 44.085 139.565 45.005 139.785 ;
        RECT 49.670 139.665 52.005 139.785 ;
        RECT 55.145 139.685 56.515 140.465 ;
        RECT 56.525 140.435 57.470 140.465 ;
        RECT 58.960 140.435 59.130 140.515 ;
        RECT 59.430 140.465 59.600 140.655 ;
        RECT 62.645 140.485 62.815 140.675 ;
        RECT 63.110 140.485 63.280 140.705 ;
        RECT 64.770 140.675 65.715 140.705 ;
        RECT 65.725 140.675 69.200 141.585 ;
        RECT 70.335 140.675 71.685 141.585 ;
        RECT 74.905 141.355 75.835 141.585 ;
        RECT 71.935 140.675 75.835 141.355 ;
        RECT 75.855 140.760 76.285 141.545 ;
        RECT 78.805 141.495 79.755 141.585 ;
        RECT 76.765 140.675 78.595 141.355 ;
        RECT 78.805 140.675 80.735 141.495 ;
        RECT 81.365 141.385 82.310 141.585 ;
        RECT 81.365 140.705 84.115 141.385 ;
        RECT 81.365 140.675 82.310 140.705 ;
        RECT 63.620 140.515 63.740 140.625 ;
        RECT 56.525 139.755 59.275 140.435 ;
        RECT 51.085 139.555 52.005 139.665 ;
        RECT 56.525 139.555 57.470 139.755 ;
        RECT 59.285 139.555 62.760 140.465 ;
        RECT 64.030 140.435 64.200 140.655 ;
        RECT 65.870 140.485 66.040 140.675 ;
        RECT 66.790 140.465 66.960 140.655 ;
        RECT 70.005 140.520 70.165 140.630 ;
        RECT 70.465 140.485 70.635 140.675 ;
        RECT 75.250 140.485 75.420 140.675 ;
        RECT 76.500 140.515 76.620 140.625 ;
        RECT 78.285 140.485 78.455 140.675 ;
        RECT 80.585 140.655 80.735 140.675 ;
        RECT 79.665 140.465 79.835 140.655 ;
        RECT 80.125 140.465 80.295 140.655 ;
        RECT 80.585 140.485 80.755 140.655 ;
        RECT 81.100 140.515 81.220 140.625 ;
        RECT 83.800 140.485 83.970 140.705 ;
        RECT 84.125 140.675 87.600 141.585 ;
        RECT 88.725 140.675 90.095 141.455 ;
        RECT 90.115 140.675 91.465 141.585 ;
        RECT 91.855 141.475 92.775 141.585 ;
        RECT 91.855 141.355 94.190 141.475 ;
        RECT 98.855 141.355 99.775 141.575 ;
        RECT 91.855 140.675 101.135 141.355 ;
        RECT 101.615 140.760 102.045 141.545 ;
        RECT 107.805 141.495 108.755 141.585 ;
        RECT 111.485 141.495 112.435 141.585 ;
        RECT 102.985 140.675 106.655 141.485 ;
        RECT 106.825 140.675 108.755 141.495 ;
        RECT 108.965 140.675 110.335 141.485 ;
        RECT 110.505 140.675 112.435 141.495 ;
        RECT 112.845 141.495 113.795 141.585 ;
        RECT 112.845 140.675 114.775 141.495 ;
        RECT 118.145 141.355 119.075 141.585 ;
        RECT 115.175 140.675 119.075 141.355 ;
        RECT 119.085 140.675 120.915 141.485 ;
        RECT 120.925 140.675 126.435 141.485 ;
        RECT 126.445 140.675 127.815 141.485 ;
        RECT 84.270 140.485 84.440 140.675 ;
        RECT 86.105 140.465 86.275 140.655 ;
        RECT 88.405 140.485 88.575 140.655 ;
        RECT 88.865 140.485 89.035 140.675 ;
        RECT 89.380 140.515 89.500 140.625 ;
        RECT 91.165 140.485 91.335 140.675 ;
        RECT 88.405 140.465 88.555 140.485 ;
        RECT 92.085 140.465 92.255 140.655 ;
        RECT 92.545 140.465 92.715 140.655 ;
        RECT 93.925 140.465 94.095 140.655 ;
        RECT 96.225 140.465 96.395 140.655 ;
        RECT 96.740 140.515 96.860 140.625 ;
        RECT 97.145 140.485 97.315 140.655 ;
        RECT 100.825 140.485 100.995 140.675 ;
        RECT 101.340 140.515 101.460 140.625 ;
        RECT 102.205 140.485 102.375 140.655 ;
        RECT 102.665 140.520 102.825 140.630 ;
        RECT 97.165 140.465 97.315 140.485 ;
        RECT 103.585 140.465 103.755 140.655 ;
        RECT 104.045 140.485 104.215 140.655 ;
        RECT 106.345 140.485 106.515 140.675 ;
        RECT 106.825 140.655 106.975 140.675 ;
        RECT 106.805 140.485 106.975 140.655 ;
        RECT 110.025 140.485 110.195 140.675 ;
        RECT 110.505 140.655 110.655 140.675 ;
        RECT 114.625 140.655 114.775 140.675 ;
        RECT 110.485 140.485 110.655 140.655 ;
        RECT 104.065 140.465 104.215 140.485 ;
        RECT 106.365 140.465 106.515 140.485 ;
        RECT 112.050 140.465 112.220 140.655 ;
        RECT 114.165 140.465 114.335 140.655 ;
        RECT 114.625 140.485 114.795 140.655 ;
        RECT 116.465 140.465 116.635 140.655 ;
        RECT 118.490 140.485 118.660 140.675 ;
        RECT 120.605 140.485 120.775 140.675 ;
        RECT 126.125 140.465 126.295 140.675 ;
        RECT 127.505 140.465 127.675 140.675 ;
        RECT 65.690 140.435 66.635 140.465 ;
        RECT 62.975 139.595 63.405 140.380 ;
        RECT 63.885 139.755 66.635 140.435 ;
        RECT 65.690 139.555 66.635 139.755 ;
        RECT 66.645 139.555 70.120 140.465 ;
        RECT 70.695 139.785 79.975 140.465 ;
        RECT 79.985 139.785 82.725 140.465 ;
        RECT 70.695 139.665 73.030 139.785 ;
        RECT 70.695 139.555 71.615 139.665 ;
        RECT 77.695 139.565 78.615 139.785 ;
        RECT 82.745 139.655 86.415 140.465 ;
        RECT 86.625 139.645 88.555 140.465 ;
        RECT 86.625 139.555 87.575 139.645 ;
        RECT 88.735 139.595 89.165 140.380 ;
        RECT 89.645 139.655 92.395 140.465 ;
        RECT 92.405 139.685 93.775 140.465 ;
        RECT 93.785 139.685 95.155 140.465 ;
        RECT 95.175 139.555 96.525 140.465 ;
        RECT 97.165 139.645 99.095 140.465 ;
        RECT 99.685 139.785 102.110 140.465 ;
        RECT 102.525 139.655 103.895 140.465 ;
        RECT 104.065 139.645 105.995 140.465 ;
        RECT 106.365 139.645 108.295 140.465 ;
        RECT 108.735 139.785 112.635 140.465 ;
        RECT 98.145 139.555 99.095 139.645 ;
        RECT 105.045 139.555 105.995 139.645 ;
        RECT 107.345 139.555 108.295 139.645 ;
        RECT 111.705 139.555 112.635 139.785 ;
        RECT 112.645 139.655 114.475 140.465 ;
        RECT 114.495 139.595 114.925 140.380 ;
        RECT 114.945 139.655 116.775 140.465 ;
        RECT 117.155 139.785 126.435 140.465 ;
        RECT 117.155 139.665 119.490 139.785 ;
        RECT 117.155 139.555 118.075 139.665 ;
        RECT 124.155 139.565 125.075 139.785 ;
        RECT 126.445 139.655 127.815 140.465 ;
      LAYER nwell ;
        RECT 29.650 136.435 128.010 139.265 ;
      LAYER pwell ;
        RECT 29.845 135.235 31.215 136.045 ;
        RECT 31.685 135.235 33.515 136.045 ;
        RECT 33.525 135.235 39.035 136.045 ;
        RECT 39.055 135.235 40.405 136.145 ;
        RECT 40.795 136.035 41.715 136.145 ;
        RECT 40.795 135.915 43.130 136.035 ;
        RECT 47.795 135.915 48.715 136.135 ;
        RECT 40.795 135.235 50.075 135.915 ;
        RECT 50.095 135.320 50.525 136.105 ;
        RECT 53.745 135.915 54.675 136.145 ;
        RECT 56.285 136.055 57.235 136.145 ;
        RECT 50.775 135.235 54.675 135.915 ;
        RECT 55.305 135.235 57.235 136.055 ;
        RECT 57.530 135.235 66.635 135.915 ;
        RECT 66.645 135.235 70.315 136.045 ;
        RECT 73.525 135.915 74.455 136.145 ;
        RECT 70.555 135.235 74.455 135.915 ;
        RECT 74.465 135.235 75.835 136.045 ;
        RECT 75.855 135.320 76.285 136.105 ;
        RECT 80.645 136.055 81.595 136.145 ;
        RECT 82.945 136.055 83.895 136.145 ;
        RECT 85.245 136.055 86.195 136.145 ;
        RECT 76.765 135.235 80.435 136.045 ;
        RECT 80.645 135.235 82.575 136.055 ;
        RECT 82.945 135.235 84.875 136.055 ;
        RECT 85.245 135.235 87.175 136.055 ;
        RECT 100.205 135.915 101.135 136.145 ;
        RECT 87.805 135.235 96.910 135.915 ;
        RECT 97.235 135.235 101.135 135.915 ;
        RECT 101.615 135.320 102.045 136.105 ;
        RECT 102.075 135.235 103.425 136.145 ;
        RECT 103.815 136.035 104.735 136.145 ;
        RECT 103.815 135.915 106.150 136.035 ;
        RECT 110.815 135.915 111.735 136.135 ;
        RECT 103.815 135.235 113.095 135.915 ;
        RECT 113.105 135.235 114.475 136.015 ;
        RECT 114.495 135.235 115.845 136.145 ;
        RECT 116.235 136.035 117.155 136.145 ;
        RECT 116.235 135.915 118.570 136.035 ;
        RECT 123.235 135.915 124.155 136.135 ;
        RECT 116.235 135.235 125.515 135.915 ;
        RECT 126.445 135.235 127.815 136.045 ;
        RECT 29.985 135.025 30.155 135.235 ;
        RECT 31.420 135.075 31.540 135.185 ;
        RECT 32.745 135.025 32.915 135.215 ;
        RECT 33.205 135.045 33.375 135.235 ;
        RECT 33.480 135.025 33.650 135.215 ;
        RECT 37.805 135.025 37.975 135.215 ;
        RECT 38.725 135.045 38.895 135.235 ;
        RECT 39.185 135.045 39.355 135.235 ;
        RECT 47.465 135.025 47.635 135.215 ;
        RECT 49.765 135.045 49.935 135.235 ;
        RECT 54.090 135.045 54.260 135.235 ;
        RECT 55.305 135.215 55.455 135.235 ;
        RECT 54.880 135.075 55.000 135.185 ;
        RECT 55.285 135.045 55.455 135.215 ;
        RECT 57.585 135.070 57.745 135.180 ;
        RECT 58.045 135.045 58.215 135.215 ;
        RECT 58.065 135.025 58.215 135.045 ;
        RECT 29.845 134.215 31.215 135.025 ;
        RECT 31.225 134.215 33.055 135.025 ;
        RECT 33.065 134.345 36.965 135.025 ;
        RECT 33.065 134.115 33.995 134.345 ;
        RECT 37.215 134.155 37.645 134.940 ;
        RECT 37.665 134.345 46.945 135.025 ;
        RECT 47.325 134.345 56.605 135.025 ;
        RECT 39.025 134.125 39.945 134.345 ;
        RECT 44.610 134.225 46.945 134.345 ;
        RECT 46.025 134.115 46.945 134.225 ;
        RECT 48.685 134.125 49.605 134.345 ;
        RECT 54.270 134.225 56.605 134.345 ;
        RECT 55.685 134.115 56.605 134.225 ;
        RECT 58.065 134.205 59.995 135.025 ;
        RECT 60.350 134.995 60.520 135.215 ;
        RECT 63.620 135.075 63.740 135.185 ;
        RECT 64.030 135.025 64.200 135.215 ;
        RECT 66.325 135.045 66.495 135.235 ;
        RECT 67.705 135.025 67.875 135.215 ;
        RECT 70.005 135.045 70.175 135.235 ;
        RECT 72.490 135.025 72.660 135.215 ;
        RECT 73.870 135.045 74.040 135.235 ;
        RECT 74.145 135.025 74.315 135.215 ;
        RECT 75.525 135.025 75.695 135.235 ;
        RECT 76.500 135.180 76.620 135.185 ;
        RECT 76.445 135.075 76.620 135.180 ;
        RECT 76.445 135.070 76.605 135.075 ;
        RECT 80.125 135.025 80.295 135.235 ;
        RECT 82.425 135.215 82.575 135.235 ;
        RECT 84.725 135.215 84.875 135.235 ;
        RECT 87.025 135.215 87.175 135.235 ;
        RECT 80.585 135.025 80.755 135.215 ;
        RECT 81.965 135.025 82.135 135.215 ;
        RECT 82.425 135.045 82.595 135.215 ;
        RECT 84.725 135.045 84.895 135.215 ;
        RECT 86.750 135.025 86.920 135.215 ;
        RECT 87.025 135.045 87.195 135.215 ;
        RECT 87.485 135.185 87.655 135.215 ;
        RECT 87.485 135.075 87.660 135.185 ;
        RECT 87.485 135.025 87.655 135.075 ;
        RECT 87.945 135.045 88.115 135.235 ;
        RECT 92.730 135.025 92.900 135.215 ;
        RECT 95.765 135.025 95.935 135.215 ;
        RECT 100.550 135.045 100.720 135.235 ;
        RECT 101.340 135.075 101.460 135.185 ;
        RECT 102.205 135.045 102.375 135.235 ;
        RECT 105.425 135.025 105.595 135.215 ;
        RECT 106.160 135.025 106.330 135.215 ;
        RECT 110.485 135.070 110.645 135.180 ;
        RECT 112.785 135.045 112.955 135.235 ;
        RECT 114.165 135.025 114.335 135.235 ;
        RECT 114.625 135.045 114.795 135.235 ;
        RECT 118.490 135.025 118.660 135.215 ;
        RECT 119.225 135.025 119.395 135.215 ;
        RECT 120.660 135.075 120.780 135.185 ;
        RECT 121.065 135.025 121.235 135.215 ;
        RECT 122.445 135.025 122.615 135.215 ;
        RECT 125.205 135.045 125.375 135.235 ;
        RECT 126.125 135.025 126.295 135.215 ;
        RECT 127.505 135.025 127.675 135.235 ;
        RECT 62.010 134.995 62.955 135.025 ;
        RECT 60.205 134.315 62.955 134.995 ;
        RECT 59.045 134.115 59.995 134.205 ;
        RECT 62.010 134.115 62.955 134.315 ;
        RECT 62.975 134.155 63.405 134.940 ;
        RECT 63.885 134.115 67.360 135.025 ;
        RECT 67.575 134.115 68.925 135.025 ;
        RECT 69.175 134.345 73.075 135.025 ;
        RECT 72.145 134.115 73.075 134.345 ;
        RECT 73.095 134.115 74.445 135.025 ;
        RECT 74.465 134.245 75.835 135.025 ;
        RECT 76.765 134.215 80.435 135.025 ;
        RECT 80.455 134.115 81.805 135.025 ;
        RECT 81.835 134.115 83.185 135.025 ;
        RECT 83.435 134.345 87.335 135.025 ;
        RECT 86.405 134.115 87.335 134.345 ;
        RECT 87.355 134.115 88.705 135.025 ;
        RECT 88.735 134.155 89.165 134.940 ;
        RECT 89.415 134.345 93.315 135.025 ;
        RECT 93.335 134.345 96.075 135.025 ;
        RECT 96.455 134.345 105.735 135.025 ;
        RECT 105.745 134.345 109.645 135.025 ;
        RECT 92.385 134.115 93.315 134.345 ;
        RECT 96.455 134.225 98.790 134.345 ;
        RECT 96.455 134.115 97.375 134.225 ;
        RECT 103.455 134.125 104.375 134.345 ;
        RECT 105.745 134.115 106.675 134.345 ;
        RECT 110.805 134.215 114.475 135.025 ;
        RECT 114.495 134.155 114.925 134.940 ;
        RECT 115.175 134.345 119.075 135.025 ;
        RECT 118.145 134.115 119.075 134.345 ;
        RECT 119.095 134.115 120.445 135.025 ;
        RECT 120.925 134.245 122.295 135.025 ;
        RECT 122.305 134.245 123.675 135.025 ;
        RECT 123.685 134.215 126.435 135.025 ;
        RECT 126.445 134.215 127.815 135.025 ;
      LAYER nwell ;
        RECT 29.650 130.995 128.010 133.825 ;
      LAYER pwell ;
        RECT 29.845 129.795 31.215 130.605 ;
        RECT 32.155 129.795 33.505 130.705 ;
        RECT 33.525 129.795 34.895 130.575 ;
        RECT 38.105 130.475 39.035 130.705 ;
        RECT 40.405 130.475 41.325 130.695 ;
        RECT 47.405 130.595 48.325 130.705 ;
        RECT 45.990 130.475 48.325 130.595 ;
        RECT 35.135 129.795 39.035 130.475 ;
        RECT 39.045 129.795 48.325 130.475 ;
        RECT 48.705 129.795 50.075 130.575 ;
        RECT 50.095 129.880 50.525 130.665 ;
        RECT 50.545 130.475 51.475 130.705 ;
        RECT 56.745 130.615 57.695 130.705 ;
        RECT 50.545 129.795 54.445 130.475 ;
        RECT 55.765 129.795 57.695 130.615 ;
        RECT 61.105 130.475 62.035 130.705 ;
        RECT 65.245 130.475 66.175 130.705 ;
        RECT 58.135 129.795 62.035 130.475 ;
        RECT 62.275 129.795 66.175 130.475 ;
        RECT 66.555 130.595 67.475 130.705 ;
        RECT 66.555 130.475 68.890 130.595 ;
        RECT 73.555 130.475 74.475 130.695 ;
        RECT 66.555 129.795 75.835 130.475 ;
        RECT 75.855 129.880 76.285 130.665 ;
        RECT 79.505 130.475 80.435 130.705 ;
        RECT 76.535 129.795 80.435 130.475 ;
        RECT 80.815 130.595 81.735 130.705 ;
        RECT 80.815 130.475 83.150 130.595 ;
        RECT 87.815 130.475 88.735 130.695 ;
        RECT 92.315 130.595 93.235 130.705 ;
        RECT 80.815 129.795 90.095 130.475 ;
        RECT 90.105 129.795 91.475 130.575 ;
        RECT 92.315 130.475 94.650 130.595 ;
        RECT 99.315 130.475 100.235 130.695 ;
        RECT 92.315 129.795 101.595 130.475 ;
        RECT 101.615 129.880 102.045 130.665 ;
        RECT 102.075 129.795 103.425 130.705 ;
        RECT 103.445 129.795 104.815 130.575 ;
        RECT 104.825 129.795 106.195 130.605 ;
        RECT 109.405 130.475 110.335 130.705 ;
        RECT 106.435 129.795 110.335 130.475 ;
        RECT 110.345 129.795 111.715 130.575 ;
        RECT 115.845 130.475 116.775 130.705 ;
        RECT 112.875 129.795 116.775 130.475 ;
        RECT 117.255 129.795 118.605 130.705 ;
        RECT 118.625 129.795 119.995 130.575 ;
        RECT 120.925 129.795 126.435 130.605 ;
        RECT 126.445 129.795 127.815 130.605 ;
        RECT 29.985 129.585 30.155 129.795 ;
        RECT 31.420 129.635 31.540 129.745 ;
        RECT 31.825 129.640 31.985 129.750 ;
        RECT 33.205 129.605 33.375 129.795 ;
        RECT 33.665 129.605 33.835 129.795 ;
        RECT 35.045 129.585 35.215 129.775 ;
        RECT 35.505 129.585 35.675 129.775 ;
        RECT 36.940 129.635 37.060 129.745 ;
        RECT 37.860 129.635 37.980 129.745 ;
        RECT 38.265 129.585 38.435 129.775 ;
        RECT 38.450 129.605 38.620 129.795 ;
        RECT 39.185 129.605 39.355 129.795 ;
        RECT 39.645 129.585 39.815 129.775 ;
        RECT 41.025 129.585 41.195 129.775 ;
        RECT 42.405 129.585 42.575 129.775 ;
        RECT 48.845 129.605 49.015 129.795 ;
        RECT 50.960 129.605 51.130 129.795 ;
        RECT 55.765 129.775 55.915 129.795 ;
        RECT 52.985 129.585 53.155 129.775 ;
        RECT 55.285 129.640 55.445 129.750 ;
        RECT 55.745 129.605 55.915 129.775 ;
        RECT 61.450 129.605 61.620 129.795 ;
        RECT 62.645 129.585 62.815 129.775 ;
        RECT 64.485 129.585 64.655 129.775 ;
        RECT 65.590 129.605 65.760 129.795 ;
        RECT 65.865 129.585 66.035 129.775 ;
        RECT 66.325 129.585 66.495 129.775 ;
        RECT 67.760 129.635 67.880 129.745 ;
        RECT 75.525 129.605 75.695 129.795 ;
        RECT 77.365 129.585 77.535 129.775 ;
        RECT 78.745 129.585 78.915 129.775 ;
        RECT 79.850 129.605 80.020 129.795 ;
        RECT 88.405 129.585 88.575 129.775 ;
        RECT 89.785 129.605 89.955 129.795 ;
        RECT 91.165 129.605 91.335 129.795 ;
        RECT 91.680 129.635 91.800 129.745 ;
        RECT 98.525 129.585 98.695 129.775 ;
        RECT 99.040 129.635 99.160 129.745 ;
        RECT 100.365 129.585 100.535 129.775 ;
        RECT 100.880 129.635 101.000 129.745 ;
        RECT 101.285 129.605 101.455 129.795 ;
        RECT 102.205 129.605 102.375 129.795 ;
        RECT 104.505 129.585 104.675 129.795 ;
        RECT 105.885 129.605 106.055 129.795 ;
        RECT 109.750 129.605 109.920 129.795 ;
        RECT 110.485 129.605 110.655 129.795 ;
        RECT 112.325 129.640 112.485 129.750 ;
        RECT 114.165 129.585 114.335 129.775 ;
        RECT 116.190 129.605 116.360 129.795 ;
        RECT 116.980 129.635 117.100 129.745 ;
        RECT 117.385 129.605 117.555 129.795 ;
        RECT 118.765 129.605 118.935 129.795 ;
        RECT 120.605 129.640 120.765 129.750 ;
        RECT 124.285 129.585 124.455 129.775 ;
        RECT 126.125 129.585 126.295 129.795 ;
        RECT 127.505 129.585 127.675 129.795 ;
        RECT 29.845 128.775 31.215 129.585 ;
        RECT 31.685 128.775 35.355 129.585 ;
        RECT 35.375 128.675 36.725 129.585 ;
        RECT 37.215 128.715 37.645 129.500 ;
        RECT 38.125 128.805 39.495 129.585 ;
        RECT 39.515 128.675 40.865 129.585 ;
        RECT 40.885 128.805 42.255 129.585 ;
        RECT 42.275 128.675 43.625 129.585 ;
        RECT 44.015 128.905 53.295 129.585 ;
        RECT 53.675 128.905 62.955 129.585 ;
        RECT 44.015 128.785 46.350 128.905 ;
        RECT 44.015 128.675 44.935 128.785 ;
        RECT 51.015 128.685 51.935 128.905 ;
        RECT 53.675 128.785 56.010 128.905 ;
        RECT 53.675 128.675 54.595 128.785 ;
        RECT 60.675 128.685 61.595 128.905 ;
        RECT 62.975 128.715 63.405 129.500 ;
        RECT 63.425 128.805 64.795 129.585 ;
        RECT 64.815 128.675 66.165 129.585 ;
        RECT 66.185 128.805 67.555 129.585 ;
        RECT 68.395 128.905 77.675 129.585 ;
        RECT 68.395 128.785 70.730 128.905 ;
        RECT 68.395 128.675 69.315 128.785 ;
        RECT 75.395 128.685 76.315 128.905 ;
        RECT 77.685 128.775 79.055 129.585 ;
        RECT 79.435 128.905 88.715 129.585 ;
        RECT 79.435 128.785 81.770 128.905 ;
        RECT 79.435 128.675 80.355 128.785 ;
        RECT 86.435 128.685 87.355 128.905 ;
        RECT 88.735 128.715 89.165 129.500 ;
        RECT 89.555 128.905 98.835 129.585 ;
        RECT 89.555 128.785 91.890 128.905 ;
        RECT 89.555 128.675 90.475 128.785 ;
        RECT 96.555 128.685 97.475 128.905 ;
        RECT 99.305 128.805 100.675 129.585 ;
        RECT 101.145 128.775 104.815 129.585 ;
        RECT 105.195 128.905 114.475 129.585 ;
        RECT 105.195 128.785 107.530 128.905 ;
        RECT 105.195 128.675 106.115 128.785 ;
        RECT 112.195 128.685 113.115 128.905 ;
        RECT 114.495 128.715 114.925 129.500 ;
        RECT 115.315 128.905 124.595 129.585 ;
        RECT 115.315 128.785 117.650 128.905 ;
        RECT 115.315 128.675 116.235 128.785 ;
        RECT 122.315 128.685 123.235 128.905 ;
        RECT 124.605 128.775 126.435 129.585 ;
        RECT 126.445 128.775 127.815 129.585 ;
      LAYER nwell ;
        RECT 29.650 125.555 128.010 128.385 ;
      LAYER pwell ;
        RECT 29.845 124.355 31.215 125.165 ;
        RECT 31.225 124.355 33.975 125.165 ;
        RECT 34.185 125.035 36.395 125.265 ;
        RECT 39.115 125.035 40.045 125.255 ;
        RECT 45.025 125.035 45.955 125.265 ;
        RECT 34.185 124.355 44.555 125.035 ;
        RECT 45.025 124.355 48.925 125.035 ;
        RECT 50.095 124.440 50.525 125.225 ;
        RECT 51.145 124.355 53.755 125.265 ;
        RECT 55.365 125.175 56.315 125.265 ;
        RECT 57.665 125.175 58.615 125.265 ;
        RECT 54.385 124.355 56.315 125.175 ;
        RECT 56.685 124.355 58.615 125.175 ;
        RECT 59.195 125.155 60.115 125.265 ;
        RECT 59.195 125.035 61.530 125.155 ;
        RECT 66.195 125.035 67.115 125.255 ;
        RECT 59.195 124.355 68.475 125.035 ;
        RECT 68.485 124.355 69.855 125.165 ;
        RECT 69.865 124.355 73.535 125.165 ;
        RECT 73.545 124.355 74.915 125.135 ;
        RECT 75.855 124.440 76.285 125.225 ;
        RECT 76.305 124.355 81.815 125.165 ;
        RECT 81.825 124.355 87.335 125.165 ;
        RECT 87.345 124.355 88.715 125.135 ;
        RECT 88.725 124.355 90.095 125.165 ;
        RECT 90.105 124.355 95.615 125.165 ;
        RECT 95.635 124.355 96.985 125.265 ;
        RECT 97.925 124.355 101.595 125.165 ;
        RECT 101.615 124.440 102.045 125.225 ;
        RECT 102.985 124.355 108.495 125.165 ;
        RECT 108.515 124.355 109.865 125.265 ;
        RECT 110.805 124.355 114.475 125.165 ;
        RECT 114.485 124.355 119.995 125.165 ;
        RECT 120.015 124.355 121.365 125.265 ;
        RECT 121.385 124.355 122.755 125.135 ;
        RECT 122.765 124.355 124.135 125.135 ;
        RECT 124.605 124.355 126.435 125.165 ;
        RECT 126.445 124.355 127.815 125.165 ;
        RECT 29.985 124.145 30.155 124.355 ;
        RECT 31.420 124.195 31.540 124.305 ;
        RECT 33.665 124.165 33.835 124.355 ;
        RECT 36.885 124.145 37.055 124.335 ;
        RECT 44.245 124.165 44.415 124.355 ;
        RECT 44.760 124.195 44.880 124.305 ;
        RECT 45.440 124.165 45.610 124.355 ;
        RECT 47.925 124.145 48.095 124.335 ;
        RECT 49.305 124.145 49.475 124.335 ;
        RECT 49.765 124.305 49.925 124.310 ;
        RECT 49.765 124.200 49.940 124.305 ;
        RECT 49.820 124.195 49.940 124.200 ;
        RECT 50.740 124.195 50.860 124.305 ;
        RECT 51.605 124.145 51.775 124.335 ;
        RECT 53.440 124.165 53.610 124.355 ;
        RECT 54.385 124.335 54.535 124.355 ;
        RECT 56.685 124.335 56.835 124.355 ;
        RECT 53.960 124.195 54.080 124.305 ;
        RECT 54.365 124.165 54.535 124.335 ;
        RECT 56.665 124.165 56.835 124.335 ;
        RECT 57.125 124.145 57.295 124.335 ;
        RECT 58.505 124.145 58.675 124.335 ;
        RECT 59.020 124.195 59.140 124.305 ;
        RECT 62.645 124.145 62.815 124.335 ;
        RECT 64.025 124.190 64.185 124.300 ;
        RECT 64.485 124.145 64.655 124.335 ;
        RECT 66.785 124.145 66.955 124.335 ;
        RECT 68.165 124.165 68.335 124.355 ;
        RECT 69.545 124.165 69.715 124.355 ;
        RECT 70.465 124.145 70.635 124.335 ;
        RECT 70.930 124.145 71.100 124.335 ;
        RECT 73.225 124.165 73.395 124.355 ;
        RECT 73.685 124.165 73.855 124.355 ;
        RECT 74.605 124.145 74.775 124.335 ;
        RECT 75.525 124.200 75.685 124.310 ;
        RECT 78.285 124.145 78.455 124.335 ;
        RECT 81.505 124.165 81.675 124.355 ;
        RECT 83.805 124.145 83.975 124.335 ;
        RECT 85.185 124.145 85.355 124.335 ;
        RECT 85.700 124.195 85.820 124.305 ;
        RECT 86.110 124.145 86.280 124.335 ;
        RECT 87.025 124.165 87.195 124.355 ;
        RECT 87.485 124.165 87.655 124.355 ;
        RECT 89.380 124.195 89.500 124.305 ;
        RECT 89.785 124.165 89.955 124.355 ;
        RECT 93.005 124.145 93.175 124.335 ;
        RECT 94.385 124.145 94.555 124.335 ;
        RECT 94.845 124.145 95.015 124.335 ;
        RECT 95.305 124.165 95.475 124.355 ;
        RECT 96.685 124.165 96.855 124.355 ;
        RECT 97.605 124.200 97.765 124.310 ;
        RECT 98.525 124.145 98.695 124.335 ;
        RECT 98.985 124.145 99.155 124.335 ;
        RECT 101.285 124.165 101.455 124.355 ;
        RECT 102.665 124.145 102.835 124.335 ;
        RECT 103.125 124.145 103.295 124.335 ;
        RECT 104.560 124.195 104.680 124.305 ;
        RECT 108.185 124.145 108.355 124.355 ;
        RECT 108.645 124.145 108.815 124.335 ;
        RECT 109.565 124.165 109.735 124.355 ;
        RECT 110.080 124.195 110.200 124.305 ;
        RECT 110.485 124.200 110.645 124.310 ;
        RECT 111.865 124.145 112.035 124.335 ;
        RECT 112.325 124.145 112.495 124.335 ;
        RECT 114.165 124.165 114.335 124.355 ;
        RECT 115.545 124.190 115.705 124.300 ;
        RECT 116.005 124.145 116.175 124.335 ;
        RECT 119.685 124.165 119.855 124.355 ;
        RECT 120.145 124.165 120.315 124.355 ;
        RECT 121.525 124.165 121.695 124.355 ;
        RECT 123.825 124.165 123.995 124.355 ;
        RECT 124.340 124.195 124.460 124.305 ;
        RECT 126.125 124.165 126.295 124.355 ;
        RECT 127.505 124.145 127.675 124.355 ;
        RECT 29.845 123.335 31.215 124.145 ;
        RECT 31.685 123.335 37.195 124.145 ;
        RECT 37.215 123.275 37.645 124.060 ;
        RECT 37.865 123.465 48.235 124.145 ;
        RECT 37.865 123.235 40.075 123.465 ;
        RECT 42.795 123.245 43.725 123.465 ;
        RECT 48.245 123.365 49.615 124.145 ;
        RECT 50.085 123.335 51.915 124.145 ;
        RECT 51.925 123.335 57.435 124.145 ;
        RECT 57.455 123.235 58.805 124.145 ;
        RECT 59.285 123.335 62.955 124.145 ;
        RECT 62.975 123.275 63.405 124.060 ;
        RECT 64.345 123.365 65.715 124.145 ;
        RECT 65.725 123.335 67.095 124.145 ;
        RECT 67.105 123.335 70.775 124.145 ;
        RECT 70.785 123.235 73.395 124.145 ;
        RECT 73.545 123.335 74.915 124.145 ;
        RECT 74.925 123.335 78.595 124.145 ;
        RECT 78.605 123.335 84.115 124.145 ;
        RECT 84.135 123.235 85.485 124.145 ;
        RECT 85.965 123.235 88.575 124.145 ;
        RECT 88.735 123.275 89.165 124.060 ;
        RECT 89.645 123.335 93.315 124.145 ;
        RECT 93.335 123.235 94.685 124.145 ;
        RECT 94.705 123.365 96.075 124.145 ;
        RECT 96.085 123.335 98.835 124.145 ;
        RECT 98.845 123.365 100.215 124.145 ;
        RECT 100.225 123.335 102.975 124.145 ;
        RECT 102.985 123.365 104.355 124.145 ;
        RECT 104.825 123.335 108.495 124.145 ;
        RECT 108.505 123.365 109.875 124.145 ;
        RECT 110.345 123.335 112.175 124.145 ;
        RECT 112.185 123.365 113.555 124.145 ;
        RECT 114.495 123.275 114.925 124.060 ;
        RECT 115.865 123.465 126.235 124.145 ;
        RECT 120.375 123.245 121.305 123.465 ;
        RECT 124.025 123.235 126.235 123.465 ;
        RECT 126.445 123.335 127.815 124.145 ;
      LAYER nwell ;
        RECT 29.650 120.115 128.010 122.945 ;
      LAYER pwell ;
        RECT 29.845 118.915 31.215 119.725 ;
        RECT 31.225 118.915 36.735 119.725 ;
        RECT 36.745 118.915 38.115 119.695 ;
        RECT 38.125 118.915 39.495 119.695 ;
        RECT 39.705 119.595 41.915 119.825 ;
        RECT 44.635 119.595 45.565 119.815 ;
        RECT 39.705 118.915 50.075 119.595 ;
        RECT 50.095 119.000 50.525 119.785 ;
        RECT 50.545 118.915 51.915 119.695 ;
        RECT 52.855 118.915 54.205 119.825 ;
        RECT 54.225 118.915 55.595 119.725 ;
        RECT 55.605 118.915 56.975 119.695 ;
        RECT 56.985 118.915 58.355 119.695 ;
        RECT 58.565 119.595 60.775 119.825 ;
        RECT 63.495 119.595 64.425 119.815 ;
        RECT 58.565 118.915 68.935 119.595 ;
        RECT 68.945 118.915 70.315 119.695 ;
        RECT 70.795 118.915 72.145 119.825 ;
        RECT 72.175 118.915 73.525 119.825 ;
        RECT 73.545 118.915 74.915 119.695 ;
        RECT 75.855 119.000 76.285 119.785 ;
        RECT 76.305 118.915 77.675 119.725 ;
        RECT 77.685 118.915 79.055 119.695 ;
        RECT 79.265 119.595 81.475 119.825 ;
        RECT 84.195 119.595 85.125 119.815 ;
        RECT 79.265 118.915 89.635 119.595 ;
        RECT 89.645 118.915 91.015 119.695 ;
        RECT 91.225 119.595 93.435 119.825 ;
        RECT 96.155 119.595 97.085 119.815 ;
        RECT 91.225 118.915 101.595 119.595 ;
        RECT 101.615 119.000 102.045 119.785 ;
        RECT 103.185 119.595 105.395 119.825 ;
        RECT 108.115 119.595 109.045 119.815 ;
        RECT 103.185 118.915 113.555 119.595 ;
        RECT 113.565 118.915 114.935 119.695 ;
        RECT 116.065 119.595 118.275 119.825 ;
        RECT 120.995 119.595 121.925 119.815 ;
        RECT 116.065 118.915 126.435 119.595 ;
        RECT 126.445 118.915 127.815 119.725 ;
        RECT 29.985 118.705 30.155 118.915 ;
        RECT 31.420 118.755 31.540 118.865 ;
        RECT 35.045 118.705 35.215 118.895 ;
        RECT 36.425 118.705 36.595 118.915 ;
        RECT 36.885 118.865 37.055 118.915 ;
        RECT 36.885 118.755 37.060 118.865 ;
        RECT 36.885 118.725 37.055 118.755 ;
        RECT 37.805 118.705 37.975 118.895 ;
        RECT 38.265 118.725 38.435 118.915 ;
        RECT 39.185 118.705 39.355 118.895 ;
        RECT 40.565 118.705 40.735 118.895 ;
        RECT 41.945 118.705 42.115 118.895 ;
        RECT 49.765 118.725 49.935 118.915 ;
        RECT 51.605 118.725 51.775 118.915 ;
        RECT 52.525 118.760 52.685 118.870 ;
        RECT 53.905 118.725 54.075 118.915 ;
        RECT 55.285 118.725 55.455 118.915 ;
        RECT 56.665 118.725 56.835 118.915 ;
        RECT 57.125 118.725 57.295 118.915 ;
        RECT 62.645 118.705 62.815 118.895 ;
        RECT 68.625 118.725 68.795 118.915 ;
        RECT 69.085 118.725 69.255 118.915 ;
        RECT 70.520 118.755 70.640 118.865 ;
        RECT 70.925 118.725 71.095 118.915 ;
        RECT 72.305 118.725 72.475 118.915 ;
        RECT 73.685 118.705 73.855 118.915 ;
        RECT 75.525 118.760 75.685 118.870 ;
        RECT 77.365 118.725 77.535 118.915 ;
        RECT 77.825 118.725 77.995 118.915 ;
        RECT 84.265 118.705 84.435 118.895 ;
        RECT 84.780 118.755 84.900 118.865 ;
        RECT 85.185 118.705 85.355 118.895 ;
        RECT 87.485 118.705 87.655 118.895 ;
        RECT 88.405 118.750 88.565 118.860 ;
        RECT 89.325 118.725 89.495 118.915 ;
        RECT 89.785 118.725 89.955 118.915 ;
        RECT 99.445 118.705 99.615 118.895 ;
        RECT 101.285 118.725 101.455 118.915 ;
        RECT 102.665 118.760 102.825 118.870 ;
        RECT 110.025 118.705 110.195 118.895 ;
        RECT 111.405 118.705 111.575 118.895 ;
        RECT 112.785 118.705 112.955 118.895 ;
        RECT 113.245 118.725 113.415 118.915 ;
        RECT 114.165 118.705 114.335 118.895 ;
        RECT 114.625 118.725 114.795 118.915 ;
        RECT 115.545 118.760 115.705 118.870 ;
        RECT 125.205 118.705 125.375 118.895 ;
        RECT 126.125 118.725 126.295 118.915 ;
        RECT 127.505 118.705 127.675 118.915 ;
        RECT 29.845 117.895 31.215 118.705 ;
        RECT 31.685 117.895 35.355 118.705 ;
        RECT 35.375 117.795 36.725 118.705 ;
        RECT 37.215 117.835 37.645 118.620 ;
        RECT 37.675 117.795 39.025 118.705 ;
        RECT 39.055 117.795 40.405 118.705 ;
        RECT 40.435 117.795 41.785 118.705 ;
        RECT 41.805 118.025 52.175 118.705 ;
        RECT 46.315 117.805 47.245 118.025 ;
        RECT 49.965 117.795 52.175 118.025 ;
        RECT 52.585 118.025 62.955 118.705 ;
        RECT 52.585 117.795 54.795 118.025 ;
        RECT 57.515 117.805 58.445 118.025 ;
        RECT 62.975 117.835 63.405 118.620 ;
        RECT 63.625 118.025 73.995 118.705 ;
        RECT 74.205 118.025 84.575 118.705 ;
        RECT 63.625 117.795 65.835 118.025 ;
        RECT 68.555 117.805 69.485 118.025 ;
        RECT 74.205 117.795 76.415 118.025 ;
        RECT 79.135 117.805 80.065 118.025 ;
        RECT 85.045 117.925 86.415 118.705 ;
        RECT 86.435 117.795 87.785 118.705 ;
        RECT 88.735 117.835 89.165 118.620 ;
        RECT 89.385 118.025 99.755 118.705 ;
        RECT 99.965 118.025 110.335 118.705 ;
        RECT 89.385 117.795 91.595 118.025 ;
        RECT 94.315 117.805 95.245 118.025 ;
        RECT 99.965 117.795 102.175 118.025 ;
        RECT 104.895 117.805 105.825 118.025 ;
        RECT 110.355 117.795 111.705 118.705 ;
        RECT 111.735 117.795 113.085 118.705 ;
        RECT 113.105 117.895 114.475 118.705 ;
        RECT 114.495 117.835 114.925 118.620 ;
        RECT 115.145 118.025 125.515 118.705 ;
        RECT 115.145 117.795 117.355 118.025 ;
        RECT 120.075 117.805 121.005 118.025 ;
        RECT 126.445 117.895 127.815 118.705 ;
      LAYER nwell ;
        RECT 29.650 114.675 128.010 117.505 ;
      LAYER pwell ;
        RECT 29.845 113.475 31.215 114.285 ;
        RECT 31.685 113.475 37.195 114.285 ;
        RECT 37.215 113.560 37.645 114.345 ;
        RECT 38.325 114.155 40.535 114.385 ;
        RECT 43.255 114.155 44.185 114.375 ;
        RECT 38.325 113.475 48.695 114.155 ;
        RECT 48.705 113.475 50.075 114.285 ;
        RECT 50.095 113.560 50.525 114.345 ;
        RECT 50.545 113.475 51.915 114.285 ;
        RECT 51.925 113.475 57.435 114.285 ;
        RECT 57.455 113.475 58.805 114.385 ;
        RECT 58.825 113.475 61.575 114.285 ;
        RECT 61.595 113.475 62.945 114.385 ;
        RECT 62.975 113.560 63.405 114.345 ;
        RECT 63.895 113.475 65.245 114.385 ;
        RECT 65.465 114.155 67.675 114.385 ;
        RECT 70.395 114.155 71.325 114.375 ;
        RECT 65.465 113.475 75.835 114.155 ;
        RECT 75.855 113.560 76.285 114.345 ;
        RECT 76.305 113.475 81.815 114.285 ;
        RECT 81.825 113.475 87.335 114.285 ;
        RECT 87.355 113.475 88.705 114.385 ;
        RECT 88.735 113.560 89.165 114.345 ;
        RECT 89.385 114.155 91.595 114.385 ;
        RECT 94.315 114.155 95.245 114.375 ;
        RECT 89.385 113.475 99.755 114.155 ;
        RECT 99.775 113.475 101.125 114.385 ;
        RECT 101.615 113.560 102.045 114.345 ;
        RECT 102.535 113.475 103.885 114.385 ;
        RECT 104.105 114.155 106.315 114.385 ;
        RECT 109.035 114.155 109.965 114.375 ;
        RECT 104.105 113.475 114.475 114.155 ;
        RECT 114.495 113.560 114.925 114.345 ;
        RECT 114.945 113.475 117.695 114.285 ;
        RECT 117.715 113.475 119.065 114.385 ;
        RECT 120.015 113.475 121.365 114.385 ;
        RECT 121.385 113.475 125.055 114.285 ;
        RECT 125.065 113.475 126.435 114.255 ;
        RECT 126.445 113.475 127.815 114.285 ;
        RECT 29.985 113.285 30.155 113.475 ;
        RECT 31.420 113.315 31.540 113.425 ;
        RECT 36.885 113.285 37.055 113.475 ;
        RECT 37.860 113.315 37.980 113.425 ;
        RECT 48.385 113.285 48.555 113.475 ;
        RECT 49.765 113.285 49.935 113.475 ;
        RECT 51.605 113.285 51.775 113.475 ;
        RECT 57.125 113.285 57.295 113.475 ;
        RECT 58.505 113.285 58.675 113.475 ;
        RECT 61.265 113.285 61.435 113.475 ;
        RECT 61.725 113.285 61.895 113.475 ;
        RECT 63.620 113.315 63.740 113.425 ;
        RECT 64.025 113.285 64.195 113.475 ;
        RECT 75.525 113.285 75.695 113.475 ;
        RECT 81.505 113.285 81.675 113.475 ;
        RECT 87.025 113.285 87.195 113.475 ;
        RECT 87.485 113.285 87.655 113.475 ;
        RECT 99.445 113.285 99.615 113.475 ;
        RECT 100.825 113.285 100.995 113.475 ;
        RECT 101.340 113.315 101.460 113.425 ;
        RECT 102.260 113.315 102.380 113.425 ;
        RECT 102.665 113.285 102.835 113.475 ;
        RECT 114.165 113.285 114.335 113.475 ;
        RECT 117.385 113.285 117.555 113.475 ;
        RECT 117.845 113.285 118.015 113.475 ;
        RECT 119.685 113.320 119.845 113.430 ;
        RECT 121.065 113.285 121.235 113.475 ;
        RECT 124.745 113.285 124.915 113.475 ;
        RECT 126.115 113.285 126.285 113.475 ;
        RECT 127.505 113.285 127.675 113.475 ;
      LAYER nwell ;
        RECT 20.485 54.580 29.875 66.420 ;
        RECT 31.685 54.590 41.075 66.430 ;
        RECT 42.905 54.560 52.295 66.400 ;
        RECT 54.155 54.540 63.545 66.380 ;
        RECT 65.375 54.530 74.765 66.370 ;
        RECT 76.615 54.520 86.005 66.360 ;
        RECT 87.865 54.530 97.255 66.370 ;
        RECT 99.145 54.520 108.535 66.360 ;
        RECT 110.415 54.520 119.805 66.360 ;
        RECT 121.665 54.520 131.055 66.360 ;
        RECT 132.415 54.490 139.375 66.330 ;
        RECT 20.655 49.020 23.115 53.210 ;
      LAYER pwell ;
        RECT 20.555 45.340 22.915 48.340 ;
      LAYER nwell ;
        RECT 24.735 45.940 29.125 53.130 ;
        RECT 31.855 49.030 34.315 53.220 ;
      LAYER pwell ;
        RECT 31.755 45.350 34.115 48.350 ;
      LAYER nwell ;
        RECT 35.935 45.950 40.325 53.140 ;
        RECT 43.075 49.000 45.535 53.190 ;
      LAYER pwell ;
        RECT 42.975 45.320 45.335 48.320 ;
      LAYER nwell ;
        RECT 47.155 45.920 51.545 53.110 ;
        RECT 54.325 48.980 56.785 53.170 ;
      LAYER pwell ;
        RECT 54.225 45.300 56.585 48.300 ;
      LAYER nwell ;
        RECT 58.405 45.900 62.795 53.090 ;
        RECT 65.545 48.970 68.005 53.160 ;
      LAYER pwell ;
        RECT 65.445 45.290 67.805 48.290 ;
      LAYER nwell ;
        RECT 69.625 45.890 74.015 53.080 ;
        RECT 76.785 48.960 79.245 53.150 ;
      LAYER pwell ;
        RECT 76.685 45.280 79.045 48.280 ;
      LAYER nwell ;
        RECT 80.865 45.880 85.255 53.070 ;
        RECT 88.035 48.970 90.495 53.160 ;
      LAYER pwell ;
        RECT 87.935 45.290 90.295 48.290 ;
      LAYER nwell ;
        RECT 92.115 45.890 96.505 53.080 ;
        RECT 99.315 48.960 101.775 53.150 ;
      LAYER pwell ;
        RECT 99.215 45.280 101.575 48.280 ;
      LAYER nwell ;
        RECT 103.395 45.880 107.785 53.070 ;
        RECT 110.585 48.960 113.045 53.150 ;
      LAYER pwell ;
        RECT 110.485 45.280 112.845 48.280 ;
      LAYER nwell ;
        RECT 114.665 45.880 119.055 53.070 ;
        RECT 121.835 48.960 124.295 53.150 ;
      LAYER pwell ;
        RECT 121.735 45.280 124.095 48.280 ;
      LAYER nwell ;
        RECT 125.915 45.880 130.305 53.070 ;
        RECT 19.615 32.280 24.005 39.470 ;
      LAYER pwell ;
        RECT 25.825 37.070 28.185 40.070 ;
      LAYER nwell ;
        RECT 25.625 32.200 28.085 36.390 ;
        RECT 30.895 32.280 35.285 39.470 ;
      LAYER pwell ;
        RECT 37.105 37.070 39.465 40.070 ;
      LAYER nwell ;
        RECT 36.905 32.200 39.365 36.390 ;
        RECT 42.185 32.260 46.575 39.450 ;
      LAYER pwell ;
        RECT 48.395 37.050 50.755 40.050 ;
      LAYER nwell ;
        RECT 48.195 32.180 50.655 36.370 ;
        RECT 53.405 32.260 57.795 39.450 ;
      LAYER pwell ;
        RECT 59.615 37.050 61.975 40.050 ;
      LAYER nwell ;
        RECT 59.415 32.180 61.875 36.370 ;
        RECT 64.605 32.260 68.995 39.450 ;
      LAYER pwell ;
        RECT 70.815 37.050 73.175 40.050 ;
      LAYER nwell ;
        RECT 70.615 32.180 73.075 36.370 ;
        RECT 75.895 32.250 80.285 39.440 ;
      LAYER pwell ;
        RECT 82.105 37.040 84.465 40.040 ;
      LAYER nwell ;
        RECT 81.905 32.170 84.365 36.360 ;
        RECT 87.135 32.270 91.525 39.460 ;
      LAYER pwell ;
        RECT 93.345 37.060 95.705 40.060 ;
      LAYER nwell ;
        RECT 93.145 32.190 95.605 36.380 ;
        RECT 98.345 32.290 102.735 39.480 ;
      LAYER pwell ;
        RECT 104.555 37.080 106.915 40.080 ;
      LAYER nwell ;
        RECT 104.355 32.210 106.815 36.400 ;
        RECT 109.545 32.330 113.935 39.520 ;
      LAYER pwell ;
        RECT 115.755 37.120 118.115 40.120 ;
      LAYER nwell ;
        RECT 115.555 32.250 118.015 36.440 ;
        RECT 120.755 32.350 125.145 39.540 ;
      LAYER pwell ;
        RECT 126.965 37.140 129.325 40.140 ;
      LAYER nwell ;
        RECT 126.765 32.270 129.225 36.460 ;
        RECT 18.865 18.990 28.255 30.830 ;
        RECT 30.145 18.990 39.535 30.830 ;
        RECT 41.435 18.970 50.825 30.810 ;
        RECT 52.655 18.970 62.045 30.810 ;
        RECT 63.855 18.970 73.245 30.810 ;
        RECT 75.145 18.960 84.535 30.800 ;
        RECT 86.385 18.980 95.775 30.820 ;
        RECT 97.595 19.000 106.985 30.840 ;
        RECT 108.795 19.040 118.185 30.880 ;
        RECT 120.005 19.060 129.395 30.900 ;
        RECT 131.725 19.030 138.685 30.870 ;
      LAYER li1 ;
        RECT 29.840 211.205 127.820 211.375 ;
        RECT 29.925 210.455 31.135 211.205 ;
        RECT 31.770 210.660 37.115 211.205 ;
        RECT 29.925 209.915 30.445 210.455 ;
        RECT 30.615 209.745 31.135 210.285 ;
        RECT 29.925 208.655 31.135 209.745 ;
        RECT 33.360 209.090 33.710 210.340 ;
        RECT 35.190 209.830 35.530 210.660 ;
        RECT 37.285 210.480 37.575 211.205 ;
        RECT 37.745 210.455 38.955 211.205 ;
        RECT 39.130 210.660 44.475 211.205 ;
        RECT 44.650 210.660 49.995 211.205 ;
        RECT 31.770 208.655 37.115 209.090 ;
        RECT 37.285 208.655 37.575 209.820 ;
        RECT 37.745 209.745 38.265 210.285 ;
        RECT 38.435 209.915 38.955 210.455 ;
        RECT 37.745 208.655 38.955 209.745 ;
        RECT 40.720 209.090 41.070 210.340 ;
        RECT 42.550 209.830 42.890 210.660 ;
        RECT 46.240 209.090 46.590 210.340 ;
        RECT 48.070 209.830 48.410 210.660 ;
        RECT 50.165 210.480 50.455 211.205 ;
        RECT 50.625 210.455 51.835 211.205 ;
        RECT 52.010 210.660 57.355 211.205 ;
        RECT 57.530 210.660 62.875 211.205 ;
        RECT 39.130 208.655 44.475 209.090 ;
        RECT 44.650 208.655 49.995 209.090 ;
        RECT 50.165 208.655 50.455 209.820 ;
        RECT 50.625 209.745 51.145 210.285 ;
        RECT 51.315 209.915 51.835 210.455 ;
        RECT 50.625 208.655 51.835 209.745 ;
        RECT 53.600 209.090 53.950 210.340 ;
        RECT 55.430 209.830 55.770 210.660 ;
        RECT 59.120 209.090 59.470 210.340 ;
        RECT 60.950 209.830 61.290 210.660 ;
        RECT 63.045 210.480 63.335 211.205 ;
        RECT 63.505 210.455 64.715 211.205 ;
        RECT 64.890 210.660 70.235 211.205 ;
        RECT 70.410 210.660 75.755 211.205 ;
        RECT 52.010 208.655 57.355 209.090 ;
        RECT 57.530 208.655 62.875 209.090 ;
        RECT 63.045 208.655 63.335 209.820 ;
        RECT 63.505 209.745 64.025 210.285 ;
        RECT 64.195 209.915 64.715 210.455 ;
        RECT 63.505 208.655 64.715 209.745 ;
        RECT 66.480 209.090 66.830 210.340 ;
        RECT 68.310 209.830 68.650 210.660 ;
        RECT 72.000 209.090 72.350 210.340 ;
        RECT 73.830 209.830 74.170 210.660 ;
        RECT 75.925 210.480 76.215 211.205 ;
        RECT 76.385 210.455 77.595 211.205 ;
        RECT 77.770 210.660 83.115 211.205 ;
        RECT 83.290 210.660 88.635 211.205 ;
        RECT 64.890 208.655 70.235 209.090 ;
        RECT 70.410 208.655 75.755 209.090 ;
        RECT 75.925 208.655 76.215 209.820 ;
        RECT 76.385 209.745 76.905 210.285 ;
        RECT 77.075 209.915 77.595 210.455 ;
        RECT 76.385 208.655 77.595 209.745 ;
        RECT 79.360 209.090 79.710 210.340 ;
        RECT 81.190 209.830 81.530 210.660 ;
        RECT 84.880 209.090 85.230 210.340 ;
        RECT 86.710 209.830 87.050 210.660 ;
        RECT 88.805 210.480 89.095 211.205 ;
        RECT 89.265 210.455 90.475 211.205 ;
        RECT 90.650 210.660 95.995 211.205 ;
        RECT 96.170 210.660 101.515 211.205 ;
        RECT 77.770 208.655 83.115 209.090 ;
        RECT 83.290 208.655 88.635 209.090 ;
        RECT 88.805 208.655 89.095 209.820 ;
        RECT 89.265 209.745 89.785 210.285 ;
        RECT 89.955 209.915 90.475 210.455 ;
        RECT 89.265 208.655 90.475 209.745 ;
        RECT 92.240 209.090 92.590 210.340 ;
        RECT 94.070 209.830 94.410 210.660 ;
        RECT 97.760 209.090 98.110 210.340 ;
        RECT 99.590 209.830 99.930 210.660 ;
        RECT 101.685 210.480 101.975 211.205 ;
        RECT 102.145 210.455 103.355 211.205 ;
        RECT 103.530 210.660 108.875 211.205 ;
        RECT 109.050 210.660 114.395 211.205 ;
        RECT 90.650 208.655 95.995 209.090 ;
        RECT 96.170 208.655 101.515 209.090 ;
        RECT 101.685 208.655 101.975 209.820 ;
        RECT 102.145 209.745 102.665 210.285 ;
        RECT 102.835 209.915 103.355 210.455 ;
        RECT 102.145 208.655 103.355 209.745 ;
        RECT 105.120 209.090 105.470 210.340 ;
        RECT 106.950 209.830 107.290 210.660 ;
        RECT 110.640 209.090 110.990 210.340 ;
        RECT 112.470 209.830 112.810 210.660 ;
        RECT 114.565 210.480 114.855 211.205 ;
        RECT 115.490 210.660 120.835 211.205 ;
        RECT 121.010 210.660 126.355 211.205 ;
        RECT 103.530 208.655 108.875 209.090 ;
        RECT 109.050 208.655 114.395 209.090 ;
        RECT 114.565 208.655 114.855 209.820 ;
        RECT 117.080 209.090 117.430 210.340 ;
        RECT 118.910 209.830 119.250 210.660 ;
        RECT 122.600 209.090 122.950 210.340 ;
        RECT 124.430 209.830 124.770 210.660 ;
        RECT 126.525 210.455 127.735 211.205 ;
        RECT 126.525 209.745 127.045 210.285 ;
        RECT 127.215 209.915 127.735 210.455 ;
        RECT 115.490 208.655 120.835 209.090 ;
        RECT 121.010 208.655 126.355 209.090 ;
        RECT 126.525 208.655 127.735 209.745 ;
        RECT 29.840 208.485 127.820 208.655 ;
        RECT 29.925 207.395 31.135 208.485 ;
        RECT 29.925 206.685 30.445 207.225 ;
        RECT 30.615 206.855 31.135 207.395 ;
        RECT 31.765 207.395 33.435 208.485 ;
        RECT 33.610 208.050 38.955 208.485 ;
        RECT 39.130 208.050 44.475 208.485 ;
        RECT 44.650 208.050 49.995 208.485 ;
        RECT 31.765 206.875 32.515 207.395 ;
        RECT 32.685 206.705 33.435 207.225 ;
        RECT 35.200 206.800 35.550 208.050 ;
        RECT 29.925 205.935 31.135 206.685 ;
        RECT 31.765 205.935 33.435 206.705 ;
        RECT 37.030 206.480 37.370 207.310 ;
        RECT 40.720 206.800 41.070 208.050 ;
        RECT 42.550 206.480 42.890 207.310 ;
        RECT 46.240 206.800 46.590 208.050 ;
        RECT 50.165 207.320 50.455 208.485 ;
        RECT 51.545 207.395 55.055 208.485 ;
        RECT 55.230 208.050 60.575 208.485 ;
        RECT 60.750 208.050 66.095 208.485 ;
        RECT 48.070 206.480 48.410 207.310 ;
        RECT 51.545 206.875 53.235 207.395 ;
        RECT 53.405 206.705 55.055 207.225 ;
        RECT 56.820 206.800 57.170 208.050 ;
        RECT 33.610 205.935 38.955 206.480 ;
        RECT 39.130 205.935 44.475 206.480 ;
        RECT 44.650 205.935 49.995 206.480 ;
        RECT 50.165 205.935 50.455 206.660 ;
        RECT 51.545 205.935 55.055 206.705 ;
        RECT 58.650 206.480 58.990 207.310 ;
        RECT 62.340 206.800 62.690 208.050 ;
        RECT 64.170 206.480 64.510 207.310 ;
        RECT 66.270 207.295 66.525 208.175 ;
        RECT 66.695 207.345 67.000 208.485 ;
        RECT 67.340 208.105 67.670 208.485 ;
        RECT 67.850 207.935 68.020 208.225 ;
        RECT 68.190 208.025 68.440 208.485 ;
        RECT 67.220 207.765 68.020 207.935 ;
        RECT 68.610 207.975 69.480 208.315 ;
        RECT 66.270 206.645 66.480 207.295 ;
        RECT 67.220 207.175 67.390 207.765 ;
        RECT 68.610 207.595 68.780 207.975 ;
        RECT 69.715 207.855 69.885 208.315 ;
        RECT 70.055 208.025 70.425 208.485 ;
        RECT 70.720 207.885 70.890 208.225 ;
        RECT 71.060 208.055 71.390 208.485 ;
        RECT 71.625 207.885 71.795 208.225 ;
        RECT 67.560 207.425 68.780 207.595 ;
        RECT 68.950 207.515 69.410 207.805 ;
        RECT 69.715 207.685 70.275 207.855 ;
        RECT 70.720 207.715 71.795 207.885 ;
        RECT 71.965 207.985 72.645 208.315 ;
        RECT 72.860 207.985 73.110 208.315 ;
        RECT 73.280 208.025 73.530 208.485 ;
        RECT 70.105 207.545 70.275 207.685 ;
        RECT 68.950 207.505 69.915 207.515 ;
        RECT 68.610 207.335 68.780 207.425 ;
        RECT 69.240 207.345 69.915 207.505 ;
        RECT 66.650 207.145 67.390 207.175 ;
        RECT 66.650 206.845 67.565 207.145 ;
        RECT 67.240 206.670 67.565 206.845 ;
        RECT 55.230 205.935 60.575 206.480 ;
        RECT 60.750 205.935 66.095 206.480 ;
        RECT 66.270 206.115 66.525 206.645 ;
        RECT 66.695 205.935 67.000 206.395 ;
        RECT 67.245 206.315 67.565 206.670 ;
        RECT 67.735 206.885 68.275 207.255 ;
        RECT 68.610 207.165 69.015 207.335 ;
        RECT 67.735 206.485 67.975 206.885 ;
        RECT 68.455 206.715 68.675 206.995 ;
        RECT 68.145 206.545 68.675 206.715 ;
        RECT 68.145 206.315 68.315 206.545 ;
        RECT 68.845 206.385 69.015 207.165 ;
        RECT 69.185 206.555 69.535 207.175 ;
        RECT 69.705 206.555 69.915 207.345 ;
        RECT 70.105 207.375 71.605 207.545 ;
        RECT 70.105 206.685 70.275 207.375 ;
        RECT 71.965 207.205 72.135 207.985 ;
        RECT 72.940 207.855 73.110 207.985 ;
        RECT 70.445 207.035 72.135 207.205 ;
        RECT 72.305 207.425 72.770 207.815 ;
        RECT 72.940 207.685 73.335 207.855 ;
        RECT 70.445 206.855 70.615 207.035 ;
        RECT 67.245 206.145 68.315 206.315 ;
        RECT 68.485 205.935 68.675 206.375 ;
        RECT 68.845 206.105 69.795 206.385 ;
        RECT 70.105 206.295 70.365 206.685 ;
        RECT 70.785 206.615 71.575 206.865 ;
        RECT 70.015 206.125 70.365 206.295 ;
        RECT 70.575 205.935 70.905 206.395 ;
        RECT 71.780 206.325 71.950 207.035 ;
        RECT 72.305 206.835 72.475 207.425 ;
        RECT 72.120 206.615 72.475 206.835 ;
        RECT 72.645 206.615 72.995 207.235 ;
        RECT 73.165 206.325 73.335 207.685 ;
        RECT 73.700 207.515 74.025 208.300 ;
        RECT 73.505 206.465 73.965 207.515 ;
        RECT 71.780 206.155 72.635 206.325 ;
        RECT 72.840 206.155 73.335 206.325 ;
        RECT 73.505 205.935 73.835 206.295 ;
        RECT 74.195 206.195 74.365 208.315 ;
        RECT 74.535 207.985 74.865 208.485 ;
        RECT 75.035 207.815 75.290 208.315 ;
        RECT 74.540 207.645 75.290 207.815 ;
        RECT 74.540 206.655 74.770 207.645 ;
        RECT 74.940 206.825 75.290 207.475 ;
        RECT 75.925 207.320 76.215 208.485 ;
        RECT 76.475 207.555 76.645 208.315 ;
        RECT 76.825 207.725 77.155 208.485 ;
        RECT 76.475 207.385 77.140 207.555 ;
        RECT 77.325 207.410 77.595 208.315 ;
        RECT 76.970 207.240 77.140 207.385 ;
        RECT 76.405 206.835 76.735 207.205 ;
        RECT 76.970 206.910 77.255 207.240 ;
        RECT 74.540 206.485 75.290 206.655 ;
        RECT 74.535 205.935 74.865 206.315 ;
        RECT 75.035 206.195 75.290 206.485 ;
        RECT 75.925 205.935 76.215 206.660 ;
        RECT 76.970 206.655 77.140 206.910 ;
        RECT 76.475 206.485 77.140 206.655 ;
        RECT 77.425 206.610 77.595 207.410 ;
        RECT 78.225 207.345 78.485 208.485 ;
        RECT 78.725 207.975 80.340 208.305 ;
        RECT 78.735 207.175 78.905 207.735 ;
        RECT 79.165 207.635 80.340 207.805 ;
        RECT 80.510 207.685 80.790 208.485 ;
        RECT 79.165 207.345 79.495 207.635 ;
        RECT 80.170 207.515 80.340 207.635 ;
        RECT 79.665 207.175 79.910 207.465 ;
        RECT 80.170 207.345 80.830 207.515 ;
        RECT 81.000 207.345 81.275 208.315 ;
        RECT 80.660 207.175 80.830 207.345 ;
        RECT 78.230 206.925 78.565 207.175 ;
        RECT 78.735 206.845 79.450 207.175 ;
        RECT 79.665 206.845 80.490 207.175 ;
        RECT 80.660 206.845 80.935 207.175 ;
        RECT 78.735 206.755 78.985 206.845 ;
        RECT 76.475 206.105 76.645 206.485 ;
        RECT 76.825 205.935 77.155 206.315 ;
        RECT 77.335 206.105 77.595 206.610 ;
        RECT 78.225 205.935 78.485 206.755 ;
        RECT 78.655 206.335 78.985 206.755 ;
        RECT 80.660 206.675 80.830 206.845 ;
        RECT 79.165 206.505 80.830 206.675 ;
        RECT 81.105 206.610 81.275 207.345 ;
        RECT 79.165 206.105 79.425 206.505 ;
        RECT 79.595 205.935 79.925 206.335 ;
        RECT 80.095 206.155 80.265 206.505 ;
        RECT 80.435 205.935 80.810 206.335 ;
        RECT 81.000 206.265 81.275 206.610 ;
        RECT 81.450 207.295 81.705 208.175 ;
        RECT 81.875 207.345 82.180 208.485 ;
        RECT 82.520 208.105 82.850 208.485 ;
        RECT 83.030 207.935 83.200 208.225 ;
        RECT 83.370 208.025 83.620 208.485 ;
        RECT 82.400 207.765 83.200 207.935 ;
        RECT 83.790 207.975 84.660 208.315 ;
        RECT 81.450 206.645 81.660 207.295 ;
        RECT 82.400 207.175 82.570 207.765 ;
        RECT 83.790 207.595 83.960 207.975 ;
        RECT 84.895 207.855 85.065 208.315 ;
        RECT 85.235 208.025 85.605 208.485 ;
        RECT 85.900 207.885 86.070 208.225 ;
        RECT 86.240 208.055 86.570 208.485 ;
        RECT 86.805 207.885 86.975 208.225 ;
        RECT 82.740 207.425 83.960 207.595 ;
        RECT 84.130 207.515 84.590 207.805 ;
        RECT 84.895 207.685 85.455 207.855 ;
        RECT 85.900 207.715 86.975 207.885 ;
        RECT 87.145 207.985 87.825 208.315 ;
        RECT 88.040 207.985 88.290 208.315 ;
        RECT 88.460 208.025 88.710 208.485 ;
        RECT 85.285 207.545 85.455 207.685 ;
        RECT 84.130 207.505 85.095 207.515 ;
        RECT 83.790 207.335 83.960 207.425 ;
        RECT 84.420 207.345 85.095 207.505 ;
        RECT 81.830 207.145 82.570 207.175 ;
        RECT 81.830 206.845 82.745 207.145 ;
        RECT 82.420 206.670 82.745 206.845 ;
        RECT 81.450 206.115 81.705 206.645 ;
        RECT 81.875 205.935 82.180 206.395 ;
        RECT 82.425 206.315 82.745 206.670 ;
        RECT 82.915 206.885 83.455 207.255 ;
        RECT 83.790 207.165 84.195 207.335 ;
        RECT 82.915 206.485 83.155 206.885 ;
        RECT 83.635 206.715 83.855 206.995 ;
        RECT 83.325 206.545 83.855 206.715 ;
        RECT 83.325 206.315 83.495 206.545 ;
        RECT 84.025 206.385 84.195 207.165 ;
        RECT 84.365 206.555 84.715 207.175 ;
        RECT 84.885 206.555 85.095 207.345 ;
        RECT 85.285 207.375 86.785 207.545 ;
        RECT 85.285 206.685 85.455 207.375 ;
        RECT 87.145 207.205 87.315 207.985 ;
        RECT 88.120 207.855 88.290 207.985 ;
        RECT 85.625 207.035 87.315 207.205 ;
        RECT 87.485 207.425 87.950 207.815 ;
        RECT 88.120 207.685 88.515 207.855 ;
        RECT 85.625 206.855 85.795 207.035 ;
        RECT 82.425 206.145 83.495 206.315 ;
        RECT 83.665 205.935 83.855 206.375 ;
        RECT 84.025 206.105 84.975 206.385 ;
        RECT 85.285 206.295 85.545 206.685 ;
        RECT 85.965 206.615 86.755 206.865 ;
        RECT 85.195 206.125 85.545 206.295 ;
        RECT 85.755 205.935 86.085 206.395 ;
        RECT 86.960 206.325 87.130 207.035 ;
        RECT 87.485 206.835 87.655 207.425 ;
        RECT 87.300 206.615 87.655 206.835 ;
        RECT 87.825 206.615 88.175 207.235 ;
        RECT 88.345 206.325 88.515 207.685 ;
        RECT 88.880 207.515 89.205 208.300 ;
        RECT 88.685 206.465 89.145 207.515 ;
        RECT 86.960 206.155 87.815 206.325 ;
        RECT 88.020 206.155 88.515 206.325 ;
        RECT 88.685 205.935 89.015 206.295 ;
        RECT 89.375 206.195 89.545 208.315 ;
        RECT 89.715 207.985 90.045 208.485 ;
        RECT 90.215 207.815 90.470 208.315 ;
        RECT 89.720 207.645 90.470 207.815 ;
        RECT 89.720 206.655 89.950 207.645 ;
        RECT 90.120 206.825 90.470 207.475 ;
        RECT 91.625 207.345 91.835 208.485 ;
        RECT 92.005 207.335 92.335 208.315 ;
        RECT 92.505 207.345 92.735 208.485 ;
        RECT 93.405 207.395 95.995 208.485 ;
        RECT 96.170 208.050 101.515 208.485 ;
        RECT 89.720 206.485 90.470 206.655 ;
        RECT 89.715 205.935 90.045 206.315 ;
        RECT 90.215 206.195 90.470 206.485 ;
        RECT 91.625 205.935 91.835 206.755 ;
        RECT 92.005 206.735 92.255 207.335 ;
        RECT 92.425 206.925 92.755 207.175 ;
        RECT 93.405 206.875 94.615 207.395 ;
        RECT 92.005 206.105 92.335 206.735 ;
        RECT 92.505 205.935 92.735 206.755 ;
        RECT 94.785 206.705 95.995 207.225 ;
        RECT 97.760 206.800 98.110 208.050 ;
        RECT 101.685 207.320 101.975 208.485 ;
        RECT 102.605 207.395 104.275 208.485 ;
        RECT 104.450 208.050 109.795 208.485 ;
        RECT 109.970 208.050 115.315 208.485 ;
        RECT 115.490 208.050 120.835 208.485 ;
        RECT 121.010 208.050 126.355 208.485 ;
        RECT 93.405 205.935 95.995 206.705 ;
        RECT 99.590 206.480 99.930 207.310 ;
        RECT 102.605 206.875 103.355 207.395 ;
        RECT 103.525 206.705 104.275 207.225 ;
        RECT 106.040 206.800 106.390 208.050 ;
        RECT 96.170 205.935 101.515 206.480 ;
        RECT 101.685 205.935 101.975 206.660 ;
        RECT 102.605 205.935 104.275 206.705 ;
        RECT 107.870 206.480 108.210 207.310 ;
        RECT 111.560 206.800 111.910 208.050 ;
        RECT 113.390 206.480 113.730 207.310 ;
        RECT 117.080 206.800 117.430 208.050 ;
        RECT 118.910 206.480 119.250 207.310 ;
        RECT 122.600 206.800 122.950 208.050 ;
        RECT 126.525 207.395 127.735 208.485 ;
        RECT 124.430 206.480 124.770 207.310 ;
        RECT 126.525 206.855 127.045 207.395 ;
        RECT 127.215 206.685 127.735 207.225 ;
        RECT 104.450 205.935 109.795 206.480 ;
        RECT 109.970 205.935 115.315 206.480 ;
        RECT 115.490 205.935 120.835 206.480 ;
        RECT 121.010 205.935 126.355 206.480 ;
        RECT 126.525 205.935 127.735 206.685 ;
        RECT 29.840 205.765 127.820 205.935 ;
        RECT 29.925 205.015 31.135 205.765 ;
        RECT 31.770 205.220 37.115 205.765 ;
        RECT 29.925 204.475 30.445 205.015 ;
        RECT 30.615 204.305 31.135 204.845 ;
        RECT 29.925 203.215 31.135 204.305 ;
        RECT 33.360 203.650 33.710 204.900 ;
        RECT 35.190 204.390 35.530 205.220 ;
        RECT 37.285 205.040 37.575 205.765 ;
        RECT 38.205 204.995 40.795 205.765 ;
        RECT 40.970 205.220 46.315 205.765 ;
        RECT 46.490 205.220 51.835 205.765 ;
        RECT 52.010 205.220 57.355 205.765 ;
        RECT 57.530 205.220 62.875 205.765 ;
        RECT 31.770 203.215 37.115 203.650 ;
        RECT 37.285 203.215 37.575 204.380 ;
        RECT 38.205 204.305 39.415 204.825 ;
        RECT 39.585 204.475 40.795 204.995 ;
        RECT 38.205 203.215 40.795 204.305 ;
        RECT 42.560 203.650 42.910 204.900 ;
        RECT 44.390 204.390 44.730 205.220 ;
        RECT 48.080 203.650 48.430 204.900 ;
        RECT 49.910 204.390 50.250 205.220 ;
        RECT 53.600 203.650 53.950 204.900 ;
        RECT 55.430 204.390 55.770 205.220 ;
        RECT 59.120 203.650 59.470 204.900 ;
        RECT 60.950 204.390 61.290 205.220 ;
        RECT 63.045 205.040 63.335 205.765 ;
        RECT 63.505 204.995 67.015 205.765 ;
        RECT 40.970 203.215 46.315 203.650 ;
        RECT 46.490 203.215 51.835 203.650 ;
        RECT 52.010 203.215 57.355 203.650 ;
        RECT 57.530 203.215 62.875 203.650 ;
        RECT 63.045 203.215 63.335 204.380 ;
        RECT 63.505 204.305 65.195 204.825 ;
        RECT 65.365 204.475 67.015 204.995 ;
        RECT 67.245 204.945 67.455 205.765 ;
        RECT 67.625 204.965 67.955 205.595 ;
        RECT 67.625 204.365 67.875 204.965 ;
        RECT 68.125 204.945 68.355 205.765 ;
        RECT 68.875 205.295 69.045 205.765 ;
        RECT 69.215 205.115 69.545 205.595 ;
        RECT 69.715 205.295 69.885 205.765 ;
        RECT 70.055 205.115 70.385 205.595 ;
        RECT 68.620 204.945 70.385 205.115 ;
        RECT 70.555 204.955 70.725 205.765 ;
        RECT 70.925 205.385 71.995 205.555 ;
        RECT 70.925 205.030 71.245 205.385 ;
        RECT 68.045 204.525 68.375 204.775 ;
        RECT 68.620 204.395 69.030 204.945 ;
        RECT 70.920 204.775 71.245 205.030 ;
        RECT 69.215 204.565 71.245 204.775 ;
        RECT 70.900 204.555 71.245 204.565 ;
        RECT 71.415 204.815 71.655 205.215 ;
        RECT 71.825 205.155 71.995 205.385 ;
        RECT 72.165 205.325 72.355 205.765 ;
        RECT 72.525 205.315 73.475 205.595 ;
        RECT 73.695 205.405 74.045 205.575 ;
        RECT 71.825 204.985 72.355 205.155 ;
        RECT 63.505 203.215 67.015 204.305 ;
        RECT 67.245 203.215 67.455 204.355 ;
        RECT 67.625 203.385 67.955 204.365 ;
        RECT 68.125 203.215 68.355 204.355 ;
        RECT 68.620 204.225 70.345 204.395 ;
        RECT 68.875 203.215 69.045 204.055 ;
        RECT 69.255 203.385 69.505 204.225 ;
        RECT 69.715 203.215 69.885 204.055 ;
        RECT 70.055 203.385 70.345 204.225 ;
        RECT 70.555 203.215 70.725 204.275 ;
        RECT 70.900 203.935 71.070 204.555 ;
        RECT 71.415 204.445 71.955 204.815 ;
        RECT 72.135 204.705 72.355 204.985 ;
        RECT 72.525 204.535 72.695 205.315 ;
        RECT 72.290 204.365 72.695 204.535 ;
        RECT 72.865 204.525 73.215 205.145 ;
        RECT 72.290 204.275 72.460 204.365 ;
        RECT 73.385 204.355 73.595 205.145 ;
        RECT 71.240 204.105 72.460 204.275 ;
        RECT 72.920 204.195 73.595 204.355 ;
        RECT 70.900 203.765 71.700 203.935 ;
        RECT 71.020 203.215 71.350 203.595 ;
        RECT 71.530 203.475 71.700 203.765 ;
        RECT 72.290 203.725 72.460 204.105 ;
        RECT 72.630 204.185 73.595 204.195 ;
        RECT 73.785 205.015 74.045 205.405 ;
        RECT 74.255 205.305 74.585 205.765 ;
        RECT 75.460 205.375 76.315 205.545 ;
        RECT 76.520 205.375 77.015 205.545 ;
        RECT 77.185 205.405 77.515 205.765 ;
        RECT 73.785 204.325 73.955 205.015 ;
        RECT 74.125 204.665 74.295 204.845 ;
        RECT 74.465 204.835 75.255 205.085 ;
        RECT 75.460 204.665 75.630 205.375 ;
        RECT 75.800 204.865 76.155 205.085 ;
        RECT 74.125 204.495 75.815 204.665 ;
        RECT 72.630 203.895 73.090 204.185 ;
        RECT 73.785 204.155 75.285 204.325 ;
        RECT 73.785 204.015 73.955 204.155 ;
        RECT 73.395 203.845 73.955 204.015 ;
        RECT 71.870 203.215 72.120 203.675 ;
        RECT 72.290 203.385 73.160 203.725 ;
        RECT 73.395 203.385 73.565 203.845 ;
        RECT 74.400 203.815 75.475 203.985 ;
        RECT 73.735 203.215 74.105 203.675 ;
        RECT 74.400 203.475 74.570 203.815 ;
        RECT 74.740 203.215 75.070 203.645 ;
        RECT 75.305 203.475 75.475 203.815 ;
        RECT 75.645 203.715 75.815 204.495 ;
        RECT 75.985 204.275 76.155 204.865 ;
        RECT 76.325 204.465 76.675 205.085 ;
        RECT 75.985 203.885 76.450 204.275 ;
        RECT 76.845 204.015 77.015 205.375 ;
        RECT 77.185 204.185 77.645 205.235 ;
        RECT 76.620 203.845 77.015 204.015 ;
        RECT 76.620 203.715 76.790 203.845 ;
        RECT 75.645 203.385 76.325 203.715 ;
        RECT 76.540 203.385 76.790 203.715 ;
        RECT 76.960 203.215 77.210 203.675 ;
        RECT 77.380 203.400 77.705 204.185 ;
        RECT 77.875 203.385 78.045 205.505 ;
        RECT 78.215 205.385 78.545 205.765 ;
        RECT 78.715 205.215 78.970 205.505 ;
        RECT 78.220 205.045 78.970 205.215 ;
        RECT 78.220 204.055 78.450 205.045 ;
        RECT 79.145 205.025 79.465 205.505 ;
        RECT 79.635 205.195 79.865 205.595 ;
        RECT 80.035 205.375 80.385 205.765 ;
        RECT 79.635 205.115 80.145 205.195 ;
        RECT 80.555 205.115 80.885 205.595 ;
        RECT 79.635 205.025 80.885 205.115 ;
        RECT 78.620 204.225 78.970 204.875 ;
        RECT 79.145 204.095 79.315 205.025 ;
        RECT 79.975 204.945 80.885 205.025 ;
        RECT 81.055 204.945 81.225 205.765 ;
        RECT 81.730 205.025 82.195 205.570 ;
        RECT 79.485 204.435 79.655 204.855 ;
        RECT 79.885 204.605 80.485 204.775 ;
        RECT 79.485 204.265 80.145 204.435 ;
        RECT 78.220 203.885 78.970 204.055 ;
        RECT 79.145 203.895 79.805 204.095 ;
        RECT 79.975 204.065 80.145 204.265 ;
        RECT 80.315 204.405 80.485 204.605 ;
        RECT 80.655 204.575 81.350 204.775 ;
        RECT 81.610 204.405 81.855 204.855 ;
        RECT 80.315 204.235 81.855 204.405 ;
        RECT 82.025 204.065 82.195 205.025 ;
        RECT 79.975 203.895 82.195 204.065 ;
        RECT 82.365 205.115 82.625 205.595 ;
        RECT 82.795 205.225 83.045 205.765 ;
        RECT 82.365 204.085 82.535 205.115 ;
        RECT 83.215 205.085 83.435 205.545 ;
        RECT 83.185 205.060 83.435 205.085 ;
        RECT 82.705 204.465 82.935 204.860 ;
        RECT 83.105 204.635 83.435 205.060 ;
        RECT 83.605 205.385 84.495 205.555 ;
        RECT 83.605 204.660 83.775 205.385 ;
        RECT 83.945 204.830 84.495 205.215 ;
        RECT 85.585 205.025 86.050 205.570 ;
        RECT 83.605 204.590 84.495 204.660 ;
        RECT 83.600 204.565 84.495 204.590 ;
        RECT 83.590 204.550 84.495 204.565 ;
        RECT 83.585 204.535 84.495 204.550 ;
        RECT 83.575 204.530 84.495 204.535 ;
        RECT 83.570 204.520 84.495 204.530 ;
        RECT 83.565 204.510 84.495 204.520 ;
        RECT 83.555 204.505 84.495 204.510 ;
        RECT 83.545 204.495 84.495 204.505 ;
        RECT 83.535 204.490 84.495 204.495 ;
        RECT 83.535 204.485 83.870 204.490 ;
        RECT 83.520 204.480 83.870 204.485 ;
        RECT 83.505 204.470 83.870 204.480 ;
        RECT 83.480 204.465 83.870 204.470 ;
        RECT 82.705 204.460 83.870 204.465 ;
        RECT 82.705 204.425 83.840 204.460 ;
        RECT 82.705 204.400 83.805 204.425 ;
        RECT 82.705 204.370 83.775 204.400 ;
        RECT 82.705 204.340 83.755 204.370 ;
        RECT 82.705 204.310 83.735 204.340 ;
        RECT 82.705 204.300 83.665 204.310 ;
        RECT 82.705 204.290 83.640 204.300 ;
        RECT 82.705 204.275 83.620 204.290 ;
        RECT 82.705 204.260 83.600 204.275 ;
        RECT 82.810 204.250 83.595 204.260 ;
        RECT 82.810 204.215 83.580 204.250 ;
        RECT 78.215 203.215 78.545 203.715 ;
        RECT 78.715 203.385 78.970 203.885 ;
        RECT 79.635 203.725 79.805 203.895 ;
        RECT 79.165 203.215 79.465 203.725 ;
        RECT 79.635 203.555 80.015 203.725 ;
        RECT 80.595 203.215 81.225 203.725 ;
        RECT 81.395 203.385 81.725 203.895 ;
        RECT 81.895 203.215 82.195 203.725 ;
        RECT 82.365 203.385 82.640 204.085 ;
        RECT 82.810 203.965 83.565 204.215 ;
        RECT 83.735 203.895 84.065 204.140 ;
        RECT 84.235 204.040 84.495 204.490 ;
        RECT 85.585 204.065 85.755 205.025 ;
        RECT 86.555 204.945 86.725 205.765 ;
        RECT 86.895 205.115 87.225 205.595 ;
        RECT 87.395 205.375 87.745 205.765 ;
        RECT 87.915 205.195 88.145 205.595 ;
        RECT 87.635 205.115 88.145 205.195 ;
        RECT 86.895 205.025 88.145 205.115 ;
        RECT 88.315 205.025 88.635 205.505 ;
        RECT 88.805 205.040 89.095 205.765 ;
        RECT 86.895 204.945 87.805 205.025 ;
        RECT 85.925 204.405 86.170 204.855 ;
        RECT 86.430 204.575 87.125 204.775 ;
        RECT 87.295 204.605 87.895 204.775 ;
        RECT 87.295 204.405 87.465 204.605 ;
        RECT 88.125 204.435 88.295 204.855 ;
        RECT 85.925 204.235 87.465 204.405 ;
        RECT 87.635 204.265 88.295 204.435 ;
        RECT 87.635 204.065 87.805 204.265 ;
        RECT 88.465 204.095 88.635 205.025 ;
        RECT 89.325 204.945 89.535 205.765 ;
        RECT 89.705 204.965 90.035 205.595 ;
        RECT 85.585 203.895 87.805 204.065 ;
        RECT 87.975 203.895 88.635 204.095 ;
        RECT 83.880 203.870 84.065 203.895 ;
        RECT 83.880 203.770 84.495 203.870 ;
        RECT 82.810 203.215 83.065 203.760 ;
        RECT 83.235 203.385 83.715 203.725 ;
        RECT 83.890 203.215 84.495 203.770 ;
        RECT 85.585 203.215 85.885 203.725 ;
        RECT 86.055 203.385 86.385 203.895 ;
        RECT 87.975 203.725 88.145 203.895 ;
        RECT 86.555 203.215 87.185 203.725 ;
        RECT 87.765 203.555 88.145 203.725 ;
        RECT 88.315 203.215 88.615 203.725 ;
        RECT 88.805 203.215 89.095 204.380 ;
        RECT 89.705 204.365 89.955 204.965 ;
        RECT 90.205 204.945 90.435 205.765 ;
        RECT 90.645 204.965 91.340 205.595 ;
        RECT 91.545 204.965 91.855 205.765 ;
        RECT 91.165 204.915 91.340 204.965 ;
        RECT 92.985 204.945 93.215 205.765 ;
        RECT 93.385 204.965 93.715 205.595 ;
        RECT 90.125 204.525 90.455 204.775 ;
        RECT 90.665 204.525 91.000 204.775 ;
        RECT 91.170 204.365 91.340 204.915 ;
        RECT 91.510 204.525 91.845 204.795 ;
        RECT 92.965 204.525 93.295 204.775 ;
        RECT 93.465 204.365 93.715 204.965 ;
        RECT 93.885 204.945 94.095 205.765 ;
        RECT 94.325 205.090 94.585 205.595 ;
        RECT 94.765 205.385 95.095 205.765 ;
        RECT 95.275 205.215 95.445 205.595 ;
        RECT 89.325 203.215 89.535 204.355 ;
        RECT 89.705 203.385 90.035 204.365 ;
        RECT 90.205 203.215 90.435 204.355 ;
        RECT 90.645 203.215 90.905 204.355 ;
        RECT 91.075 203.385 91.405 204.365 ;
        RECT 91.575 203.215 91.855 204.355 ;
        RECT 92.985 203.215 93.215 204.355 ;
        RECT 93.385 203.385 93.715 204.365 ;
        RECT 93.885 203.215 94.095 204.355 ;
        RECT 94.325 204.290 94.495 205.090 ;
        RECT 94.780 205.045 95.445 205.215 ;
        RECT 94.780 204.790 94.950 205.045 ;
        RECT 96.165 204.995 97.835 205.765 ;
        RECT 98.010 205.220 103.355 205.765 ;
        RECT 103.530 205.220 108.875 205.765 ;
        RECT 109.050 205.220 114.395 205.765 ;
        RECT 94.665 204.460 94.950 204.790 ;
        RECT 95.185 204.495 95.515 204.865 ;
        RECT 94.780 204.315 94.950 204.460 ;
        RECT 94.325 203.385 94.595 204.290 ;
        RECT 94.780 204.145 95.445 204.315 ;
        RECT 94.765 203.215 95.095 203.975 ;
        RECT 95.275 203.385 95.445 204.145 ;
        RECT 96.165 204.305 96.915 204.825 ;
        RECT 97.085 204.475 97.835 204.995 ;
        RECT 96.165 203.215 97.835 204.305 ;
        RECT 99.600 203.650 99.950 204.900 ;
        RECT 101.430 204.390 101.770 205.220 ;
        RECT 105.120 203.650 105.470 204.900 ;
        RECT 106.950 204.390 107.290 205.220 ;
        RECT 110.640 203.650 110.990 204.900 ;
        RECT 112.470 204.390 112.810 205.220 ;
        RECT 114.565 205.040 114.855 205.765 ;
        RECT 115.490 205.220 120.835 205.765 ;
        RECT 121.010 205.220 126.355 205.765 ;
        RECT 98.010 203.215 103.355 203.650 ;
        RECT 103.530 203.215 108.875 203.650 ;
        RECT 109.050 203.215 114.395 203.650 ;
        RECT 114.565 203.215 114.855 204.380 ;
        RECT 117.080 203.650 117.430 204.900 ;
        RECT 118.910 204.390 119.250 205.220 ;
        RECT 122.600 203.650 122.950 204.900 ;
        RECT 124.430 204.390 124.770 205.220 ;
        RECT 126.525 205.015 127.735 205.765 ;
        RECT 126.525 204.305 127.045 204.845 ;
        RECT 127.215 204.475 127.735 205.015 ;
        RECT 115.490 203.215 120.835 203.650 ;
        RECT 121.010 203.215 126.355 203.650 ;
        RECT 126.525 203.215 127.735 204.305 ;
        RECT 29.840 203.045 127.820 203.215 ;
        RECT 29.925 201.955 31.135 203.045 ;
        RECT 29.925 201.245 30.445 201.785 ;
        RECT 30.615 201.415 31.135 201.955 ;
        RECT 31.765 201.955 33.435 203.045 ;
        RECT 33.610 202.610 38.955 203.045 ;
        RECT 39.130 202.610 44.475 203.045 ;
        RECT 44.650 202.610 49.995 203.045 ;
        RECT 31.765 201.435 32.515 201.955 ;
        RECT 32.685 201.265 33.435 201.785 ;
        RECT 35.200 201.360 35.550 202.610 ;
        RECT 29.925 200.495 31.135 201.245 ;
        RECT 31.765 200.495 33.435 201.265 ;
        RECT 37.030 201.040 37.370 201.870 ;
        RECT 40.720 201.360 41.070 202.610 ;
        RECT 42.550 201.040 42.890 201.870 ;
        RECT 46.240 201.360 46.590 202.610 ;
        RECT 50.165 201.880 50.455 203.045 ;
        RECT 50.625 201.955 51.835 203.045 ;
        RECT 52.010 202.610 57.355 203.045 ;
        RECT 57.530 202.610 62.875 203.045 ;
        RECT 63.050 202.610 68.395 203.045 ;
        RECT 48.070 201.040 48.410 201.870 ;
        RECT 50.625 201.415 51.145 201.955 ;
        RECT 51.315 201.245 51.835 201.785 ;
        RECT 53.600 201.360 53.950 202.610 ;
        RECT 33.610 200.495 38.955 201.040 ;
        RECT 39.130 200.495 44.475 201.040 ;
        RECT 44.650 200.495 49.995 201.040 ;
        RECT 50.165 200.495 50.455 201.220 ;
        RECT 50.625 200.495 51.835 201.245 ;
        RECT 55.430 201.040 55.770 201.870 ;
        RECT 59.120 201.360 59.470 202.610 ;
        RECT 60.950 201.040 61.290 201.870 ;
        RECT 64.640 201.360 64.990 202.610 ;
        RECT 68.605 201.905 68.835 203.045 ;
        RECT 69.005 201.895 69.335 202.875 ;
        RECT 69.505 201.905 69.715 203.045 ;
        RECT 70.060 202.415 70.345 202.875 ;
        RECT 70.515 202.585 70.785 203.045 ;
        RECT 70.060 202.195 71.015 202.415 ;
        RECT 66.470 201.040 66.810 201.870 ;
        RECT 68.585 201.485 68.915 201.735 ;
        RECT 52.010 200.495 57.355 201.040 ;
        RECT 57.530 200.495 62.875 201.040 ;
        RECT 63.050 200.495 68.395 201.040 ;
        RECT 68.605 200.495 68.835 201.315 ;
        RECT 69.085 201.295 69.335 201.895 ;
        RECT 69.945 201.465 70.635 202.025 ;
        RECT 69.005 200.665 69.335 201.295 ;
        RECT 69.505 200.495 69.715 201.315 ;
        RECT 70.805 201.295 71.015 202.195 ;
        RECT 70.060 201.125 71.015 201.295 ;
        RECT 71.185 202.025 71.585 202.875 ;
        RECT 71.775 202.415 72.055 202.875 ;
        RECT 72.575 202.585 72.900 203.045 ;
        RECT 71.775 202.195 72.900 202.415 ;
        RECT 71.185 201.465 72.280 202.025 ;
        RECT 72.450 201.735 72.900 202.195 ;
        RECT 73.070 201.905 73.455 202.875 ;
        RECT 70.060 200.665 70.345 201.125 ;
        RECT 70.515 200.495 70.785 200.955 ;
        RECT 71.185 200.665 71.585 201.465 ;
        RECT 72.450 201.405 73.005 201.735 ;
        RECT 72.450 201.295 72.900 201.405 ;
        RECT 71.775 201.125 72.900 201.295 ;
        RECT 73.175 201.235 73.455 201.905 ;
        RECT 74.085 201.955 75.755 203.045 ;
        RECT 74.085 201.435 74.835 201.955 ;
        RECT 75.925 201.880 76.215 203.045 ;
        RECT 76.385 201.905 76.645 203.045 ;
        RECT 76.885 202.535 78.500 202.865 ;
        RECT 75.005 201.265 75.755 201.785 ;
        RECT 76.895 201.735 77.065 202.295 ;
        RECT 77.325 202.195 78.500 202.365 ;
        RECT 78.670 202.245 78.950 203.045 ;
        RECT 77.325 201.905 77.655 202.195 ;
        RECT 78.330 202.075 78.500 202.195 ;
        RECT 77.825 201.735 78.070 202.025 ;
        RECT 78.330 201.905 78.990 202.075 ;
        RECT 79.160 201.905 79.435 202.875 ;
        RECT 78.820 201.735 78.990 201.905 ;
        RECT 76.390 201.485 76.725 201.735 ;
        RECT 76.895 201.405 77.610 201.735 ;
        RECT 77.825 201.405 78.650 201.735 ;
        RECT 78.820 201.405 79.095 201.735 ;
        RECT 76.895 201.315 77.145 201.405 ;
        RECT 71.775 200.665 72.055 201.125 ;
        RECT 72.575 200.495 72.900 200.955 ;
        RECT 73.070 200.665 73.455 201.235 ;
        RECT 74.085 200.495 75.755 201.265 ;
        RECT 75.925 200.495 76.215 201.220 ;
        RECT 76.385 200.495 76.645 201.315 ;
        RECT 76.815 200.895 77.145 201.315 ;
        RECT 78.820 201.235 78.990 201.405 ;
        RECT 77.325 201.065 78.990 201.235 ;
        RECT 79.265 201.170 79.435 201.905 ;
        RECT 77.325 200.665 77.585 201.065 ;
        RECT 77.755 200.495 78.085 200.895 ;
        RECT 78.255 200.715 78.425 201.065 ;
        RECT 78.595 200.495 78.970 200.895 ;
        RECT 79.160 200.825 79.435 201.170 ;
        RECT 79.610 201.855 79.865 202.735 ;
        RECT 80.035 201.905 80.340 203.045 ;
        RECT 80.680 202.665 81.010 203.045 ;
        RECT 81.190 202.495 81.360 202.785 ;
        RECT 81.530 202.585 81.780 203.045 ;
        RECT 80.560 202.325 81.360 202.495 ;
        RECT 81.950 202.535 82.820 202.875 ;
        RECT 79.610 201.205 79.820 201.855 ;
        RECT 80.560 201.735 80.730 202.325 ;
        RECT 81.950 202.155 82.120 202.535 ;
        RECT 83.055 202.415 83.225 202.875 ;
        RECT 83.395 202.585 83.765 203.045 ;
        RECT 84.060 202.445 84.230 202.785 ;
        RECT 84.400 202.615 84.730 203.045 ;
        RECT 84.965 202.445 85.135 202.785 ;
        RECT 80.900 201.985 82.120 202.155 ;
        RECT 82.290 202.075 82.750 202.365 ;
        RECT 83.055 202.245 83.615 202.415 ;
        RECT 84.060 202.275 85.135 202.445 ;
        RECT 85.305 202.545 85.985 202.875 ;
        RECT 86.200 202.545 86.450 202.875 ;
        RECT 86.620 202.585 86.870 203.045 ;
        RECT 83.445 202.105 83.615 202.245 ;
        RECT 82.290 202.065 83.255 202.075 ;
        RECT 81.950 201.895 82.120 201.985 ;
        RECT 82.580 201.905 83.255 202.065 ;
        RECT 79.990 201.705 80.730 201.735 ;
        RECT 79.990 201.405 80.905 201.705 ;
        RECT 80.580 201.230 80.905 201.405 ;
        RECT 79.610 200.675 79.865 201.205 ;
        RECT 80.035 200.495 80.340 200.955 ;
        RECT 80.585 200.875 80.905 201.230 ;
        RECT 81.075 201.445 81.615 201.815 ;
        RECT 81.950 201.725 82.355 201.895 ;
        RECT 81.075 201.045 81.315 201.445 ;
        RECT 81.795 201.275 82.015 201.555 ;
        RECT 81.485 201.105 82.015 201.275 ;
        RECT 81.485 200.875 81.655 201.105 ;
        RECT 82.185 200.945 82.355 201.725 ;
        RECT 82.525 201.115 82.875 201.735 ;
        RECT 83.045 201.115 83.255 201.905 ;
        RECT 83.445 201.935 84.945 202.105 ;
        RECT 83.445 201.245 83.615 201.935 ;
        RECT 85.305 201.765 85.475 202.545 ;
        RECT 86.280 202.415 86.450 202.545 ;
        RECT 83.785 201.595 85.475 201.765 ;
        RECT 85.645 201.985 86.110 202.375 ;
        RECT 86.280 202.245 86.675 202.415 ;
        RECT 83.785 201.415 83.955 201.595 ;
        RECT 80.585 200.705 81.655 200.875 ;
        RECT 81.825 200.495 82.015 200.935 ;
        RECT 82.185 200.665 83.135 200.945 ;
        RECT 83.445 200.855 83.705 201.245 ;
        RECT 84.125 201.175 84.915 201.425 ;
        RECT 83.355 200.685 83.705 200.855 ;
        RECT 83.915 200.495 84.245 200.955 ;
        RECT 85.120 200.885 85.290 201.595 ;
        RECT 85.645 201.395 85.815 201.985 ;
        RECT 85.460 201.175 85.815 201.395 ;
        RECT 85.985 201.175 86.335 201.795 ;
        RECT 86.505 200.885 86.675 202.245 ;
        RECT 87.040 202.075 87.365 202.860 ;
        RECT 86.845 201.025 87.305 202.075 ;
        RECT 85.120 200.715 85.975 200.885 ;
        RECT 86.180 200.715 86.675 200.885 ;
        RECT 86.845 200.495 87.175 200.855 ;
        RECT 87.535 200.755 87.705 202.875 ;
        RECT 87.875 202.545 88.205 203.045 ;
        RECT 88.375 202.375 88.630 202.875 ;
        RECT 87.880 202.205 88.630 202.375 ;
        RECT 87.880 201.215 88.110 202.205 ;
        RECT 88.280 201.385 88.630 202.035 ;
        RECT 88.810 201.855 89.065 202.735 ;
        RECT 89.235 201.905 89.540 203.045 ;
        RECT 89.880 202.665 90.210 203.045 ;
        RECT 90.390 202.495 90.560 202.785 ;
        RECT 90.730 202.585 90.980 203.045 ;
        RECT 89.760 202.325 90.560 202.495 ;
        RECT 91.150 202.535 92.020 202.875 ;
        RECT 87.880 201.045 88.630 201.215 ;
        RECT 87.875 200.495 88.205 200.875 ;
        RECT 88.375 200.755 88.630 201.045 ;
        RECT 88.810 201.205 89.020 201.855 ;
        RECT 89.760 201.735 89.930 202.325 ;
        RECT 91.150 202.155 91.320 202.535 ;
        RECT 92.255 202.415 92.425 202.875 ;
        RECT 92.595 202.585 92.965 203.045 ;
        RECT 93.260 202.445 93.430 202.785 ;
        RECT 93.600 202.615 93.930 203.045 ;
        RECT 94.165 202.445 94.335 202.785 ;
        RECT 90.100 201.985 91.320 202.155 ;
        RECT 91.490 202.075 91.950 202.365 ;
        RECT 92.255 202.245 92.815 202.415 ;
        RECT 93.260 202.275 94.335 202.445 ;
        RECT 94.505 202.545 95.185 202.875 ;
        RECT 95.400 202.545 95.650 202.875 ;
        RECT 95.820 202.585 96.070 203.045 ;
        RECT 92.645 202.105 92.815 202.245 ;
        RECT 91.490 202.065 92.455 202.075 ;
        RECT 91.150 201.895 91.320 201.985 ;
        RECT 91.780 201.905 92.455 202.065 ;
        RECT 89.190 201.705 89.930 201.735 ;
        RECT 89.190 201.405 90.105 201.705 ;
        RECT 89.780 201.230 90.105 201.405 ;
        RECT 88.810 200.675 89.065 201.205 ;
        RECT 89.235 200.495 89.540 200.955 ;
        RECT 89.785 200.875 90.105 201.230 ;
        RECT 90.275 201.445 90.815 201.815 ;
        RECT 91.150 201.725 91.555 201.895 ;
        RECT 90.275 201.045 90.515 201.445 ;
        RECT 90.995 201.275 91.215 201.555 ;
        RECT 90.685 201.105 91.215 201.275 ;
        RECT 90.685 200.875 90.855 201.105 ;
        RECT 91.385 200.945 91.555 201.725 ;
        RECT 91.725 201.115 92.075 201.735 ;
        RECT 92.245 201.115 92.455 201.905 ;
        RECT 92.645 201.935 94.145 202.105 ;
        RECT 92.645 201.245 92.815 201.935 ;
        RECT 94.505 201.765 94.675 202.545 ;
        RECT 95.480 202.415 95.650 202.545 ;
        RECT 92.985 201.595 94.675 201.765 ;
        RECT 94.845 201.985 95.310 202.375 ;
        RECT 95.480 202.245 95.875 202.415 ;
        RECT 92.985 201.415 93.155 201.595 ;
        RECT 89.785 200.705 90.855 200.875 ;
        RECT 91.025 200.495 91.215 200.935 ;
        RECT 91.385 200.665 92.335 200.945 ;
        RECT 92.645 200.855 92.905 201.245 ;
        RECT 93.325 201.175 94.115 201.425 ;
        RECT 92.555 200.685 92.905 200.855 ;
        RECT 93.115 200.495 93.445 200.955 ;
        RECT 94.320 200.885 94.490 201.595 ;
        RECT 94.845 201.395 95.015 201.985 ;
        RECT 94.660 201.175 95.015 201.395 ;
        RECT 95.185 201.175 95.535 201.795 ;
        RECT 95.705 200.885 95.875 202.245 ;
        RECT 96.240 202.075 96.565 202.860 ;
        RECT 96.045 201.025 96.505 202.075 ;
        RECT 94.320 200.715 95.175 200.885 ;
        RECT 95.380 200.715 95.875 200.885 ;
        RECT 96.045 200.495 96.375 200.855 ;
        RECT 96.735 200.755 96.905 202.875 ;
        RECT 97.075 202.545 97.405 203.045 ;
        RECT 97.575 202.375 97.830 202.875 ;
        RECT 97.080 202.205 97.830 202.375 ;
        RECT 97.080 201.215 97.310 202.205 ;
        RECT 97.480 201.385 97.830 202.035 ;
        RECT 98.005 201.955 101.515 203.045 ;
        RECT 98.005 201.435 99.695 201.955 ;
        RECT 101.685 201.880 101.975 203.045 ;
        RECT 103.065 201.955 106.575 203.045 ;
        RECT 106.860 202.415 107.145 202.875 ;
        RECT 107.315 202.585 107.585 203.045 ;
        RECT 106.860 202.195 107.815 202.415 ;
        RECT 99.865 201.265 101.515 201.785 ;
        RECT 103.065 201.435 104.755 201.955 ;
        RECT 104.925 201.265 106.575 201.785 ;
        RECT 106.745 201.465 107.435 202.025 ;
        RECT 107.605 201.295 107.815 202.195 ;
        RECT 97.080 201.045 97.830 201.215 ;
        RECT 97.075 200.495 97.405 200.875 ;
        RECT 97.575 200.755 97.830 201.045 ;
        RECT 98.005 200.495 101.515 201.265 ;
        RECT 101.685 200.495 101.975 201.220 ;
        RECT 103.065 200.495 106.575 201.265 ;
        RECT 106.860 201.125 107.815 201.295 ;
        RECT 107.985 202.025 108.385 202.875 ;
        RECT 108.575 202.415 108.855 202.875 ;
        RECT 109.375 202.585 109.700 203.045 ;
        RECT 108.575 202.195 109.700 202.415 ;
        RECT 107.985 201.465 109.080 202.025 ;
        RECT 109.250 201.735 109.700 202.195 ;
        RECT 109.870 201.905 110.255 202.875 ;
        RECT 106.860 200.665 107.145 201.125 ;
        RECT 107.315 200.495 107.585 200.955 ;
        RECT 107.985 200.665 108.385 201.465 ;
        RECT 109.250 201.405 109.805 201.735 ;
        RECT 109.250 201.295 109.700 201.405 ;
        RECT 108.575 201.125 109.700 201.295 ;
        RECT 109.975 201.235 110.255 201.905 ;
        RECT 108.575 200.665 108.855 201.125 ;
        RECT 109.375 200.495 109.700 200.955 ;
        RECT 109.870 200.665 110.255 201.235 ;
        RECT 110.430 201.855 110.685 202.735 ;
        RECT 110.855 201.905 111.160 203.045 ;
        RECT 111.500 202.665 111.830 203.045 ;
        RECT 112.010 202.495 112.180 202.785 ;
        RECT 112.350 202.585 112.600 203.045 ;
        RECT 111.380 202.325 112.180 202.495 ;
        RECT 112.770 202.535 113.640 202.875 ;
        RECT 110.430 201.205 110.640 201.855 ;
        RECT 111.380 201.735 111.550 202.325 ;
        RECT 112.770 202.155 112.940 202.535 ;
        RECT 113.875 202.415 114.045 202.875 ;
        RECT 114.215 202.585 114.585 203.045 ;
        RECT 114.880 202.445 115.050 202.785 ;
        RECT 115.220 202.615 115.550 203.045 ;
        RECT 115.785 202.445 115.955 202.785 ;
        RECT 111.720 201.985 112.940 202.155 ;
        RECT 113.110 202.075 113.570 202.365 ;
        RECT 113.875 202.245 114.435 202.415 ;
        RECT 114.880 202.275 115.955 202.445 ;
        RECT 116.125 202.545 116.805 202.875 ;
        RECT 117.020 202.545 117.270 202.875 ;
        RECT 117.440 202.585 117.690 203.045 ;
        RECT 114.265 202.105 114.435 202.245 ;
        RECT 113.110 202.065 114.075 202.075 ;
        RECT 112.770 201.895 112.940 201.985 ;
        RECT 113.400 201.905 114.075 202.065 ;
        RECT 110.810 201.705 111.550 201.735 ;
        RECT 110.810 201.405 111.725 201.705 ;
        RECT 111.400 201.230 111.725 201.405 ;
        RECT 110.430 200.675 110.685 201.205 ;
        RECT 110.855 200.495 111.160 200.955 ;
        RECT 111.405 200.875 111.725 201.230 ;
        RECT 111.895 201.445 112.435 201.815 ;
        RECT 112.770 201.725 113.175 201.895 ;
        RECT 111.895 201.045 112.135 201.445 ;
        RECT 112.615 201.275 112.835 201.555 ;
        RECT 112.305 201.105 112.835 201.275 ;
        RECT 112.305 200.875 112.475 201.105 ;
        RECT 113.005 200.945 113.175 201.725 ;
        RECT 113.345 201.115 113.695 201.735 ;
        RECT 113.865 201.115 114.075 201.905 ;
        RECT 114.265 201.935 115.765 202.105 ;
        RECT 114.265 201.245 114.435 201.935 ;
        RECT 116.125 201.765 116.295 202.545 ;
        RECT 117.100 202.415 117.270 202.545 ;
        RECT 114.605 201.595 116.295 201.765 ;
        RECT 116.465 201.985 116.930 202.375 ;
        RECT 117.100 202.245 117.495 202.415 ;
        RECT 114.605 201.415 114.775 201.595 ;
        RECT 111.405 200.705 112.475 200.875 ;
        RECT 112.645 200.495 112.835 200.935 ;
        RECT 113.005 200.665 113.955 200.945 ;
        RECT 114.265 200.855 114.525 201.245 ;
        RECT 114.945 201.175 115.735 201.425 ;
        RECT 114.175 200.685 114.525 200.855 ;
        RECT 114.735 200.495 115.065 200.955 ;
        RECT 115.940 200.885 116.110 201.595 ;
        RECT 116.465 201.395 116.635 201.985 ;
        RECT 116.280 201.175 116.635 201.395 ;
        RECT 116.805 201.175 117.155 201.795 ;
        RECT 117.325 200.885 117.495 202.245 ;
        RECT 117.860 202.075 118.185 202.860 ;
        RECT 117.665 201.025 118.125 202.075 ;
        RECT 115.940 200.715 116.795 200.885 ;
        RECT 117.000 200.715 117.495 200.885 ;
        RECT 117.665 200.495 117.995 200.855 ;
        RECT 118.355 200.755 118.525 202.875 ;
        RECT 118.695 202.545 119.025 203.045 ;
        RECT 119.195 202.375 119.450 202.875 ;
        RECT 118.700 202.205 119.450 202.375 ;
        RECT 118.700 201.215 118.930 202.205 ;
        RECT 119.100 201.385 119.450 202.035 ;
        RECT 119.625 201.955 120.835 203.045 ;
        RECT 121.010 202.610 126.355 203.045 ;
        RECT 119.625 201.415 120.145 201.955 ;
        RECT 120.315 201.245 120.835 201.785 ;
        RECT 122.600 201.360 122.950 202.610 ;
        RECT 126.525 201.955 127.735 203.045 ;
        RECT 118.700 201.045 119.450 201.215 ;
        RECT 118.695 200.495 119.025 200.875 ;
        RECT 119.195 200.755 119.450 201.045 ;
        RECT 119.625 200.495 120.835 201.245 ;
        RECT 124.430 201.040 124.770 201.870 ;
        RECT 126.525 201.415 127.045 201.955 ;
        RECT 127.215 201.245 127.735 201.785 ;
        RECT 121.010 200.495 126.355 201.040 ;
        RECT 126.525 200.495 127.735 201.245 ;
        RECT 29.840 200.325 127.820 200.495 ;
        RECT 29.925 199.575 31.135 200.325 ;
        RECT 31.770 199.780 37.115 200.325 ;
        RECT 29.925 199.035 30.445 199.575 ;
        RECT 30.615 198.865 31.135 199.405 ;
        RECT 29.925 197.775 31.135 198.865 ;
        RECT 33.360 198.210 33.710 199.460 ;
        RECT 35.190 198.950 35.530 199.780 ;
        RECT 37.285 199.600 37.575 200.325 ;
        RECT 37.745 199.555 41.255 200.325 ;
        RECT 41.430 199.780 46.775 200.325 ;
        RECT 46.950 199.780 52.295 200.325 ;
        RECT 31.770 197.775 37.115 198.210 ;
        RECT 37.285 197.775 37.575 198.940 ;
        RECT 37.745 198.865 39.435 199.385 ;
        RECT 39.605 199.035 41.255 199.555 ;
        RECT 37.745 197.775 41.255 198.865 ;
        RECT 43.020 198.210 43.370 199.460 ;
        RECT 44.850 198.950 45.190 199.780 ;
        RECT 48.540 198.210 48.890 199.460 ;
        RECT 50.370 198.950 50.710 199.780 ;
        RECT 52.580 199.695 52.865 200.155 ;
        RECT 53.035 199.865 53.305 200.325 ;
        RECT 52.580 199.525 53.535 199.695 ;
        RECT 52.465 198.795 53.155 199.355 ;
        RECT 53.325 198.625 53.535 199.525 ;
        RECT 52.580 198.405 53.535 198.625 ;
        RECT 53.705 199.355 54.105 200.155 ;
        RECT 54.295 199.695 54.575 200.155 ;
        RECT 55.095 199.865 55.420 200.325 ;
        RECT 54.295 199.525 55.420 199.695 ;
        RECT 55.590 199.585 55.975 200.155 ;
        RECT 54.970 199.415 55.420 199.525 ;
        RECT 53.705 198.795 54.800 199.355 ;
        RECT 54.970 199.085 55.525 199.415 ;
        RECT 41.430 197.775 46.775 198.210 ;
        RECT 46.950 197.775 52.295 198.210 ;
        RECT 52.580 197.945 52.865 198.405 ;
        RECT 53.035 197.775 53.305 198.235 ;
        RECT 53.705 197.945 54.105 198.795 ;
        RECT 54.970 198.625 55.420 199.085 ;
        RECT 55.695 198.915 55.975 199.585 ;
        RECT 56.260 199.695 56.545 200.155 ;
        RECT 56.715 199.865 56.985 200.325 ;
        RECT 56.260 199.525 57.215 199.695 ;
        RECT 54.295 198.405 55.420 198.625 ;
        RECT 54.295 197.945 54.575 198.405 ;
        RECT 55.095 197.775 55.420 198.235 ;
        RECT 55.590 197.945 55.975 198.915 ;
        RECT 56.145 198.795 56.835 199.355 ;
        RECT 57.005 198.625 57.215 199.525 ;
        RECT 56.260 198.405 57.215 198.625 ;
        RECT 57.385 199.355 57.785 200.155 ;
        RECT 57.975 199.695 58.255 200.155 ;
        RECT 58.775 199.865 59.100 200.325 ;
        RECT 57.975 199.525 59.100 199.695 ;
        RECT 59.270 199.585 59.655 200.155 ;
        RECT 58.650 199.415 59.100 199.525 ;
        RECT 57.385 198.795 58.480 199.355 ;
        RECT 58.650 199.085 59.205 199.415 ;
        RECT 56.260 197.945 56.545 198.405 ;
        RECT 56.715 197.775 56.985 198.235 ;
        RECT 57.385 197.945 57.785 198.795 ;
        RECT 58.650 198.625 59.100 199.085 ;
        RECT 59.375 198.915 59.655 199.585 ;
        RECT 60.285 199.555 62.875 200.325 ;
        RECT 63.045 199.600 63.335 200.325 ;
        RECT 63.965 199.555 65.635 200.325 ;
        RECT 57.975 198.405 59.100 198.625 ;
        RECT 57.975 197.945 58.255 198.405 ;
        RECT 58.775 197.775 59.100 198.235 ;
        RECT 59.270 197.945 59.655 198.915 ;
        RECT 60.285 198.865 61.495 199.385 ;
        RECT 61.665 199.035 62.875 199.555 ;
        RECT 60.285 197.775 62.875 198.865 ;
        RECT 63.045 197.775 63.335 198.940 ;
        RECT 63.965 198.865 64.715 199.385 ;
        RECT 64.885 199.035 65.635 199.555 ;
        RECT 65.845 199.505 66.075 200.325 ;
        RECT 66.245 199.525 66.575 200.155 ;
        RECT 65.825 199.085 66.155 199.335 ;
        RECT 66.325 198.925 66.575 199.525 ;
        RECT 66.745 199.505 66.955 200.325 ;
        RECT 67.190 199.780 72.535 200.325 ;
        RECT 73.035 199.925 73.365 200.325 ;
        RECT 63.965 197.775 65.635 198.865 ;
        RECT 65.845 197.775 66.075 198.915 ;
        RECT 66.245 197.945 66.575 198.925 ;
        RECT 66.745 197.775 66.955 198.915 ;
        RECT 68.780 198.210 69.130 199.460 ;
        RECT 70.610 198.950 70.950 199.780 ;
        RECT 73.535 199.755 73.865 200.095 ;
        RECT 74.915 199.925 75.245 200.325 ;
        RECT 72.880 199.585 75.245 199.755 ;
        RECT 75.415 199.600 75.745 200.110 ;
        RECT 72.880 198.585 73.050 199.585 ;
        RECT 75.075 199.415 75.245 199.585 ;
        RECT 73.220 198.755 73.465 199.415 ;
        RECT 73.680 198.755 73.945 199.415 ;
        RECT 74.140 198.755 74.425 199.415 ;
        RECT 74.600 199.085 74.905 199.415 ;
        RECT 75.075 199.085 75.385 199.415 ;
        RECT 74.600 198.755 74.815 199.085 ;
        RECT 72.880 198.415 73.335 198.585 ;
        RECT 67.190 197.775 72.535 198.210 ;
        RECT 73.005 197.985 73.335 198.415 ;
        RECT 73.515 198.415 74.805 198.585 ;
        RECT 73.515 197.995 73.765 198.415 ;
        RECT 73.995 197.775 74.325 198.245 ;
        RECT 74.555 197.995 74.805 198.415 ;
        RECT 74.995 197.775 75.245 198.915 ;
        RECT 75.555 198.835 75.745 199.600 ;
        RECT 76.390 199.485 76.650 200.325 ;
        RECT 76.825 199.580 77.080 200.155 ;
        RECT 77.250 199.945 77.580 200.325 ;
        RECT 77.795 199.775 77.965 200.155 ;
        RECT 77.250 199.605 77.965 199.775 ;
        RECT 75.415 197.985 75.745 198.835 ;
        RECT 76.390 197.775 76.650 198.925 ;
        RECT 76.825 198.850 76.995 199.580 ;
        RECT 77.250 199.415 77.420 199.605 ;
        RECT 78.230 199.585 78.565 200.325 ;
        RECT 77.165 199.085 77.420 199.415 ;
        RECT 77.250 198.875 77.420 199.085 ;
        RECT 77.700 199.055 78.055 199.425 ;
        RECT 78.735 199.415 78.950 200.110 ;
        RECT 79.140 199.585 79.490 200.110 ;
        RECT 79.660 199.585 80.355 200.155 ;
        RECT 80.530 200.070 80.865 200.115 ;
        RECT 80.525 199.605 80.865 200.070 ;
        RECT 81.035 199.945 81.365 200.325 ;
        RECT 79.285 199.415 79.490 199.585 ;
        RECT 78.250 199.085 78.535 199.415 ;
        RECT 78.735 199.085 79.115 199.415 ;
        RECT 79.285 199.085 79.595 199.415 ;
        RECT 79.765 198.915 79.935 199.585 ;
        RECT 76.825 197.945 77.080 198.850 ;
        RECT 77.250 198.705 77.965 198.875 ;
        RECT 77.250 197.775 77.580 198.535 ;
        RECT 77.795 197.945 77.965 198.705 ;
        RECT 78.225 197.775 78.485 198.915 ;
        RECT 78.655 198.745 79.935 198.915 ;
        RECT 80.115 198.745 80.355 199.415 ;
        RECT 80.525 198.915 80.695 199.605 ;
        RECT 80.865 199.085 81.125 199.415 ;
        RECT 78.655 197.945 78.985 198.745 ;
        RECT 79.155 197.775 79.325 198.575 ;
        RECT 79.525 197.945 79.855 198.745 ;
        RECT 80.055 197.775 80.335 198.575 ;
        RECT 80.525 197.945 80.785 198.915 ;
        RECT 80.955 198.535 81.125 199.085 ;
        RECT 81.295 198.715 81.635 199.745 ;
        RECT 81.825 199.645 82.095 199.990 ;
        RECT 81.825 199.475 82.135 199.645 ;
        RECT 81.825 198.715 82.095 199.475 ;
        RECT 82.320 198.715 82.600 199.990 ;
        RECT 82.800 199.825 83.030 200.155 ;
        RECT 83.275 199.945 83.605 200.325 ;
        RECT 82.800 198.535 82.970 199.825 ;
        RECT 83.775 199.755 83.950 200.155 ;
        RECT 83.320 199.585 83.950 199.755 ;
        RECT 85.240 199.695 85.525 200.155 ;
        RECT 85.695 199.865 85.965 200.325 ;
        RECT 83.320 199.415 83.490 199.585 ;
        RECT 85.240 199.525 86.195 199.695 ;
        RECT 83.140 199.085 83.490 199.415 ;
        RECT 80.955 198.365 82.970 198.535 ;
        RECT 83.320 198.565 83.490 199.085 ;
        RECT 83.670 198.735 84.035 199.415 ;
        RECT 85.125 198.795 85.815 199.355 ;
        RECT 85.985 198.625 86.195 199.525 ;
        RECT 83.320 198.395 83.950 198.565 ;
        RECT 80.980 197.775 81.310 198.185 ;
        RECT 81.510 197.945 81.680 198.365 ;
        RECT 81.895 197.775 82.565 198.185 ;
        RECT 82.800 197.945 82.970 198.365 ;
        RECT 83.275 197.775 83.605 198.215 ;
        RECT 83.775 197.945 83.950 198.395 ;
        RECT 85.240 198.405 86.195 198.625 ;
        RECT 86.365 199.355 86.765 200.155 ;
        RECT 86.955 199.695 87.235 200.155 ;
        RECT 87.755 199.865 88.080 200.325 ;
        RECT 86.955 199.525 88.080 199.695 ;
        RECT 88.250 199.585 88.635 200.155 ;
        RECT 88.805 199.600 89.095 200.325 ;
        RECT 87.630 199.415 88.080 199.525 ;
        RECT 86.365 198.795 87.460 199.355 ;
        RECT 87.630 199.085 88.185 199.415 ;
        RECT 85.240 197.945 85.525 198.405 ;
        RECT 85.695 197.775 85.965 198.235 ;
        RECT 86.365 197.945 86.765 198.795 ;
        RECT 87.630 198.625 88.080 199.085 ;
        RECT 88.355 198.915 88.635 199.585 ;
        RECT 89.300 199.585 89.915 200.155 ;
        RECT 90.085 199.815 90.300 200.325 ;
        RECT 90.530 199.815 90.810 200.145 ;
        RECT 90.990 199.815 91.230 200.325 ;
        RECT 91.565 199.825 91.825 200.155 ;
        RECT 92.035 199.845 92.310 200.325 ;
        RECT 86.955 198.405 88.080 198.625 ;
        RECT 86.955 197.945 87.235 198.405 ;
        RECT 87.755 197.775 88.080 198.235 ;
        RECT 88.250 197.945 88.635 198.915 ;
        RECT 88.805 197.775 89.095 198.940 ;
        RECT 89.300 198.565 89.615 199.585 ;
        RECT 89.785 198.915 89.955 199.415 ;
        RECT 90.205 199.085 90.470 199.645 ;
        RECT 90.640 198.915 90.810 199.815 ;
        RECT 90.980 199.085 91.335 199.645 ;
        RECT 91.565 198.915 91.735 199.825 ;
        RECT 92.520 199.755 92.725 200.155 ;
        RECT 92.895 199.925 93.230 200.325 ;
        RECT 91.905 199.085 92.265 199.665 ;
        RECT 92.520 199.585 93.205 199.755 ;
        RECT 92.445 198.915 92.695 199.415 ;
        RECT 89.785 198.745 91.210 198.915 ;
        RECT 89.300 197.945 89.835 198.565 ;
        RECT 90.005 197.775 90.335 198.575 ;
        RECT 90.820 198.570 91.210 198.745 ;
        RECT 91.565 198.745 92.695 198.915 ;
        RECT 91.565 197.975 91.835 198.745 ;
        RECT 92.865 198.555 93.205 199.585 ;
        RECT 93.465 199.505 93.675 200.325 ;
        RECT 93.845 199.525 94.175 200.155 ;
        RECT 93.845 198.925 94.095 199.525 ;
        RECT 94.345 199.505 94.575 200.325 ;
        RECT 94.785 199.575 95.995 200.325 ;
        RECT 96.255 199.775 96.425 200.155 ;
        RECT 96.605 199.945 96.935 200.325 ;
        RECT 96.255 199.605 96.920 199.775 ;
        RECT 97.115 199.650 97.375 200.155 ;
        RECT 94.265 199.085 94.595 199.335 ;
        RECT 92.005 197.775 92.335 198.555 ;
        RECT 92.540 198.380 93.205 198.555 ;
        RECT 92.540 197.975 92.725 198.380 ;
        RECT 92.895 197.775 93.230 198.200 ;
        RECT 93.465 197.775 93.675 198.915 ;
        RECT 93.845 197.945 94.175 198.925 ;
        RECT 94.345 197.775 94.575 198.915 ;
        RECT 94.785 198.865 95.305 199.405 ;
        RECT 95.475 199.035 95.995 199.575 ;
        RECT 96.185 199.055 96.515 199.425 ;
        RECT 96.750 199.350 96.920 199.605 ;
        RECT 96.750 199.020 97.035 199.350 ;
        RECT 96.750 198.875 96.920 199.020 ;
        RECT 94.785 197.775 95.995 198.865 ;
        RECT 96.255 198.705 96.920 198.875 ;
        RECT 97.205 198.850 97.375 199.650 ;
        RECT 97.545 199.555 99.215 200.325 ;
        RECT 96.255 197.945 96.425 198.705 ;
        RECT 96.605 197.775 96.935 198.535 ;
        RECT 97.105 197.945 97.375 198.850 ;
        RECT 97.545 198.865 98.295 199.385 ;
        RECT 98.465 199.035 99.215 199.555 ;
        RECT 99.425 199.505 99.655 200.325 ;
        RECT 99.825 199.525 100.155 200.155 ;
        RECT 99.405 199.085 99.735 199.335 ;
        RECT 99.905 198.925 100.155 199.525 ;
        RECT 100.325 199.505 100.535 200.325 ;
        RECT 100.770 199.615 101.025 200.145 ;
        RECT 101.195 199.865 101.500 200.325 ;
        RECT 101.745 199.945 102.815 200.115 ;
        RECT 97.545 197.775 99.215 198.865 ;
        RECT 99.425 197.775 99.655 198.915 ;
        RECT 99.825 197.945 100.155 198.925 ;
        RECT 100.770 198.965 100.980 199.615 ;
        RECT 101.745 199.590 102.065 199.945 ;
        RECT 101.740 199.415 102.065 199.590 ;
        RECT 101.150 199.115 102.065 199.415 ;
        RECT 102.235 199.375 102.475 199.775 ;
        RECT 102.645 199.715 102.815 199.945 ;
        RECT 102.985 199.885 103.175 200.325 ;
        RECT 103.345 199.875 104.295 200.155 ;
        RECT 104.515 199.965 104.865 200.135 ;
        RECT 102.645 199.545 103.175 199.715 ;
        RECT 101.150 199.085 101.890 199.115 ;
        RECT 100.325 197.775 100.535 198.915 ;
        RECT 100.770 198.085 101.025 198.965 ;
        RECT 101.195 197.775 101.500 198.915 ;
        RECT 101.720 198.495 101.890 199.085 ;
        RECT 102.235 199.005 102.775 199.375 ;
        RECT 102.955 199.265 103.175 199.545 ;
        RECT 103.345 199.095 103.515 199.875 ;
        RECT 103.110 198.925 103.515 199.095 ;
        RECT 103.685 199.085 104.035 199.705 ;
        RECT 103.110 198.835 103.280 198.925 ;
        RECT 104.205 198.915 104.415 199.705 ;
        RECT 102.060 198.665 103.280 198.835 ;
        RECT 103.740 198.755 104.415 198.915 ;
        RECT 101.720 198.325 102.520 198.495 ;
        RECT 101.840 197.775 102.170 198.155 ;
        RECT 102.350 198.035 102.520 198.325 ;
        RECT 103.110 198.285 103.280 198.665 ;
        RECT 103.450 198.745 104.415 198.755 ;
        RECT 104.605 199.575 104.865 199.965 ;
        RECT 105.075 199.865 105.405 200.325 ;
        RECT 106.280 199.935 107.135 200.105 ;
        RECT 107.340 199.935 107.835 200.105 ;
        RECT 108.005 199.965 108.335 200.325 ;
        RECT 104.605 198.885 104.775 199.575 ;
        RECT 104.945 199.225 105.115 199.405 ;
        RECT 105.285 199.395 106.075 199.645 ;
        RECT 106.280 199.225 106.450 199.935 ;
        RECT 106.620 199.425 106.975 199.645 ;
        RECT 104.945 199.055 106.635 199.225 ;
        RECT 103.450 198.455 103.910 198.745 ;
        RECT 104.605 198.715 106.105 198.885 ;
        RECT 104.605 198.575 104.775 198.715 ;
        RECT 104.215 198.405 104.775 198.575 ;
        RECT 102.690 197.775 102.940 198.235 ;
        RECT 103.110 197.945 103.980 198.285 ;
        RECT 104.215 197.945 104.385 198.405 ;
        RECT 105.220 198.375 106.295 198.545 ;
        RECT 104.555 197.775 104.925 198.235 ;
        RECT 105.220 198.035 105.390 198.375 ;
        RECT 105.560 197.775 105.890 198.205 ;
        RECT 106.125 198.035 106.295 198.375 ;
        RECT 106.465 198.275 106.635 199.055 ;
        RECT 106.805 198.835 106.975 199.425 ;
        RECT 107.145 199.025 107.495 199.645 ;
        RECT 106.805 198.445 107.270 198.835 ;
        RECT 107.665 198.575 107.835 199.935 ;
        RECT 108.005 198.745 108.465 199.795 ;
        RECT 107.440 198.405 107.835 198.575 ;
        RECT 107.440 198.275 107.610 198.405 ;
        RECT 106.465 197.945 107.145 198.275 ;
        RECT 107.360 197.945 107.610 198.275 ;
        RECT 107.780 197.775 108.030 198.235 ;
        RECT 108.200 197.960 108.525 198.745 ;
        RECT 108.695 197.945 108.865 200.065 ;
        RECT 109.035 199.945 109.365 200.325 ;
        RECT 109.535 199.775 109.790 200.065 ;
        RECT 109.040 199.605 109.790 199.775 ;
        RECT 109.040 198.615 109.270 199.605 ;
        RECT 110.700 199.515 110.945 200.120 ;
        RECT 111.165 199.790 111.675 200.325 ;
        RECT 109.440 198.785 109.790 199.435 ;
        RECT 110.425 199.345 111.655 199.515 ;
        RECT 109.040 198.445 109.790 198.615 ;
        RECT 109.035 197.775 109.365 198.275 ;
        RECT 109.535 197.945 109.790 198.445 ;
        RECT 110.425 198.535 110.765 199.345 ;
        RECT 110.935 198.780 111.685 198.970 ;
        RECT 110.425 198.125 110.940 198.535 ;
        RECT 111.175 197.775 111.345 198.535 ;
        RECT 111.515 198.115 111.685 198.780 ;
        RECT 111.855 198.795 112.045 200.155 ;
        RECT 112.215 199.305 112.490 200.155 ;
        RECT 112.680 199.790 113.210 200.155 ;
        RECT 113.635 199.925 113.965 200.325 ;
        RECT 113.035 199.755 113.210 199.790 ;
        RECT 112.215 199.135 112.495 199.305 ;
        RECT 112.215 198.995 112.490 199.135 ;
        RECT 112.695 198.795 112.865 199.595 ;
        RECT 111.855 198.625 112.865 198.795 ;
        RECT 113.035 199.585 113.965 199.755 ;
        RECT 114.135 199.585 114.390 200.155 ;
        RECT 114.565 199.600 114.855 200.325 ;
        RECT 113.035 198.455 113.205 199.585 ;
        RECT 113.795 199.415 113.965 199.585 ;
        RECT 112.080 198.285 113.205 198.455 ;
        RECT 113.375 199.085 113.570 199.415 ;
        RECT 113.795 199.085 114.050 199.415 ;
        RECT 113.375 198.115 113.545 199.085 ;
        RECT 114.220 198.915 114.390 199.585 ;
        RECT 115.085 199.505 115.295 200.325 ;
        RECT 115.465 199.525 115.795 200.155 ;
        RECT 111.515 197.945 113.545 198.115 ;
        RECT 113.715 197.775 113.885 198.915 ;
        RECT 114.055 197.945 114.390 198.915 ;
        RECT 114.565 197.775 114.855 198.940 ;
        RECT 115.465 198.925 115.715 199.525 ;
        RECT 115.965 199.505 116.195 200.325 ;
        RECT 116.905 199.505 117.135 200.325 ;
        RECT 117.305 199.525 117.635 200.155 ;
        RECT 115.885 199.085 116.215 199.335 ;
        RECT 116.885 199.085 117.215 199.335 ;
        RECT 117.385 198.925 117.635 199.525 ;
        RECT 117.805 199.505 118.015 200.325 ;
        RECT 119.255 199.775 119.425 200.155 ;
        RECT 119.605 199.945 119.935 200.325 ;
        RECT 119.255 199.605 119.920 199.775 ;
        RECT 120.115 199.650 120.375 200.155 ;
        RECT 121.010 199.780 126.355 200.325 ;
        RECT 119.185 199.055 119.515 199.425 ;
        RECT 119.750 199.350 119.920 199.605 ;
        RECT 115.085 197.775 115.295 198.915 ;
        RECT 115.465 197.945 115.795 198.925 ;
        RECT 115.965 197.775 116.195 198.915 ;
        RECT 116.905 197.775 117.135 198.915 ;
        RECT 117.305 197.945 117.635 198.925 ;
        RECT 119.750 199.020 120.035 199.350 ;
        RECT 117.805 197.775 118.015 198.915 ;
        RECT 119.750 198.875 119.920 199.020 ;
        RECT 119.255 198.705 119.920 198.875 ;
        RECT 120.205 198.850 120.375 199.650 ;
        RECT 119.255 197.945 119.425 198.705 ;
        RECT 119.605 197.775 119.935 198.535 ;
        RECT 120.105 197.945 120.375 198.850 ;
        RECT 122.600 198.210 122.950 199.460 ;
        RECT 124.430 198.950 124.770 199.780 ;
        RECT 126.525 199.575 127.735 200.325 ;
        RECT 126.525 198.865 127.045 199.405 ;
        RECT 127.215 199.035 127.735 199.575 ;
        RECT 121.010 197.775 126.355 198.210 ;
        RECT 126.525 197.775 127.735 198.865 ;
        RECT 29.840 197.605 127.820 197.775 ;
        RECT 29.925 196.515 31.135 197.605 ;
        RECT 32.230 197.170 37.575 197.605 ;
        RECT 37.750 197.170 43.095 197.605 ;
        RECT 43.270 197.170 48.615 197.605 ;
        RECT 29.925 195.805 30.445 196.345 ;
        RECT 30.615 195.975 31.135 196.515 ;
        RECT 33.820 195.920 34.170 197.170 ;
        RECT 29.925 195.055 31.135 195.805 ;
        RECT 35.650 195.600 35.990 196.430 ;
        RECT 39.340 195.920 39.690 197.170 ;
        RECT 41.170 195.600 41.510 196.430 ;
        RECT 44.860 195.920 45.210 197.170 ;
        RECT 48.785 196.530 49.055 197.435 ;
        RECT 49.225 196.845 49.555 197.605 ;
        RECT 49.735 196.675 49.905 197.435 ;
        RECT 46.690 195.600 47.030 196.430 ;
        RECT 48.785 195.730 48.955 196.530 ;
        RECT 49.240 196.505 49.905 196.675 ;
        RECT 49.240 196.360 49.410 196.505 ;
        RECT 50.165 196.440 50.455 197.605 ;
        RECT 51.085 196.530 51.355 197.435 ;
        RECT 51.525 196.845 51.855 197.605 ;
        RECT 52.035 196.675 52.205 197.435 ;
        RECT 49.125 196.030 49.410 196.360 ;
        RECT 49.240 195.775 49.410 196.030 ;
        RECT 49.645 195.955 49.975 196.325 ;
        RECT 32.230 195.055 37.575 195.600 ;
        RECT 37.750 195.055 43.095 195.600 ;
        RECT 43.270 195.055 48.615 195.600 ;
        RECT 48.785 195.225 49.045 195.730 ;
        RECT 49.240 195.605 49.905 195.775 ;
        RECT 49.225 195.055 49.555 195.435 ;
        RECT 49.735 195.225 49.905 195.605 ;
        RECT 50.165 195.055 50.455 195.780 ;
        RECT 51.085 195.730 51.255 196.530 ;
        RECT 51.540 196.505 52.205 196.675 ;
        RECT 51.540 196.360 51.710 196.505 ;
        RECT 52.525 196.465 52.735 197.605 ;
        RECT 51.425 196.030 51.710 196.360 ;
        RECT 52.905 196.455 53.235 197.435 ;
        RECT 53.405 196.465 53.635 197.605 ;
        RECT 53.960 196.975 54.245 197.435 ;
        RECT 54.415 197.145 54.685 197.605 ;
        RECT 53.960 196.755 54.915 196.975 ;
        RECT 51.540 195.775 51.710 196.030 ;
        RECT 51.945 195.955 52.275 196.325 ;
        RECT 51.085 195.225 51.345 195.730 ;
        RECT 51.540 195.605 52.205 195.775 ;
        RECT 51.525 195.055 51.855 195.435 ;
        RECT 52.035 195.225 52.205 195.605 ;
        RECT 52.525 195.055 52.735 195.875 ;
        RECT 52.905 195.855 53.155 196.455 ;
        RECT 53.325 196.045 53.655 196.295 ;
        RECT 53.845 196.025 54.535 196.585 ;
        RECT 52.905 195.225 53.235 195.855 ;
        RECT 53.405 195.055 53.635 195.875 ;
        RECT 54.705 195.855 54.915 196.755 ;
        RECT 53.960 195.685 54.915 195.855 ;
        RECT 55.085 196.585 55.485 197.435 ;
        RECT 55.675 196.975 55.955 197.435 ;
        RECT 56.475 197.145 56.800 197.605 ;
        RECT 55.675 196.755 56.800 196.975 ;
        RECT 55.085 196.025 56.180 196.585 ;
        RECT 56.350 196.295 56.800 196.755 ;
        RECT 56.970 196.465 57.355 197.435 ;
        RECT 57.585 196.465 57.795 197.605 ;
        RECT 53.960 195.225 54.245 195.685 ;
        RECT 54.415 195.055 54.685 195.515 ;
        RECT 55.085 195.225 55.485 196.025 ;
        RECT 56.350 195.965 56.905 196.295 ;
        RECT 56.350 195.855 56.800 195.965 ;
        RECT 55.675 195.685 56.800 195.855 ;
        RECT 57.075 195.795 57.355 196.465 ;
        RECT 57.965 196.455 58.295 197.435 ;
        RECT 58.465 196.465 58.695 197.605 ;
        RECT 58.995 196.675 59.165 197.435 ;
        RECT 59.345 196.845 59.675 197.605 ;
        RECT 58.995 196.505 59.660 196.675 ;
        RECT 59.845 196.530 60.115 197.435 ;
        RECT 55.675 195.225 55.955 195.685 ;
        RECT 56.475 195.055 56.800 195.515 ;
        RECT 56.970 195.225 57.355 195.795 ;
        RECT 57.585 195.055 57.795 195.875 ;
        RECT 57.965 195.855 58.215 196.455 ;
        RECT 59.490 196.360 59.660 196.505 ;
        RECT 58.385 196.045 58.715 196.295 ;
        RECT 58.925 195.955 59.255 196.325 ;
        RECT 59.490 196.030 59.775 196.360 ;
        RECT 57.965 195.225 58.295 195.855 ;
        RECT 58.465 195.055 58.695 195.875 ;
        RECT 59.490 195.775 59.660 196.030 ;
        RECT 58.995 195.605 59.660 195.775 ;
        RECT 59.945 195.730 60.115 196.530 ;
        RECT 58.995 195.225 59.165 195.605 ;
        RECT 59.345 195.055 59.675 195.435 ;
        RECT 59.855 195.225 60.115 195.730 ;
        RECT 60.285 196.465 60.670 197.435 ;
        RECT 60.840 197.145 61.165 197.605 ;
        RECT 61.685 196.975 61.965 197.435 ;
        RECT 60.840 196.755 61.965 196.975 ;
        RECT 60.285 195.795 60.565 196.465 ;
        RECT 60.840 196.295 61.290 196.755 ;
        RECT 62.155 196.585 62.555 197.435 ;
        RECT 62.955 197.145 63.225 197.605 ;
        RECT 63.395 196.975 63.680 197.435 ;
        RECT 60.735 195.965 61.290 196.295 ;
        RECT 61.460 196.025 62.555 196.585 ;
        RECT 60.840 195.855 61.290 195.965 ;
        RECT 60.285 195.225 60.670 195.795 ;
        RECT 60.840 195.685 61.965 195.855 ;
        RECT 60.840 195.055 61.165 195.515 ;
        RECT 61.685 195.225 61.965 195.685 ;
        RECT 62.155 195.225 62.555 196.025 ;
        RECT 62.725 196.755 63.680 196.975 ;
        RECT 63.965 196.845 64.480 197.255 ;
        RECT 64.715 196.845 64.885 197.605 ;
        RECT 65.055 197.265 67.085 197.435 ;
        RECT 62.725 195.855 62.935 196.755 ;
        RECT 63.105 196.025 63.795 196.585 ;
        RECT 63.965 196.035 64.305 196.845 ;
        RECT 65.055 196.600 65.225 197.265 ;
        RECT 65.620 196.925 66.745 197.095 ;
        RECT 64.475 196.410 65.225 196.600 ;
        RECT 65.395 196.585 66.405 196.755 ;
        RECT 63.965 195.865 65.195 196.035 ;
        RECT 62.725 195.685 63.680 195.855 ;
        RECT 62.955 195.055 63.225 195.515 ;
        RECT 63.395 195.225 63.680 195.685 ;
        RECT 64.240 195.260 64.485 195.865 ;
        RECT 64.705 195.055 65.215 195.590 ;
        RECT 65.395 195.225 65.585 196.585 ;
        RECT 65.755 195.905 66.030 196.385 ;
        RECT 65.755 195.735 66.035 195.905 ;
        RECT 66.235 195.785 66.405 196.585 ;
        RECT 66.575 195.795 66.745 196.925 ;
        RECT 66.915 196.295 67.085 197.265 ;
        RECT 67.255 196.465 67.425 197.605 ;
        RECT 67.595 196.465 67.930 197.435 ;
        RECT 68.195 196.675 68.365 197.435 ;
        RECT 68.545 196.845 68.875 197.605 ;
        RECT 68.195 196.505 68.860 196.675 ;
        RECT 69.045 196.530 69.315 197.435 ;
        RECT 70.410 197.170 75.755 197.605 ;
        RECT 66.915 195.965 67.110 196.295 ;
        RECT 67.335 195.965 67.590 196.295 ;
        RECT 67.335 195.795 67.505 195.965 ;
        RECT 67.760 195.795 67.930 196.465 ;
        RECT 68.690 196.360 68.860 196.505 ;
        RECT 68.125 195.955 68.455 196.325 ;
        RECT 68.690 196.030 68.975 196.360 ;
        RECT 65.755 195.225 66.030 195.735 ;
        RECT 66.575 195.625 67.505 195.795 ;
        RECT 66.575 195.590 66.750 195.625 ;
        RECT 66.220 195.225 66.750 195.590 ;
        RECT 67.175 195.055 67.505 195.455 ;
        RECT 67.675 195.225 67.930 195.795 ;
        RECT 68.690 195.775 68.860 196.030 ;
        RECT 68.195 195.605 68.860 195.775 ;
        RECT 69.145 195.730 69.315 196.530 ;
        RECT 72.000 195.920 72.350 197.170 ;
        RECT 75.925 196.440 76.215 197.605 ;
        RECT 77.305 196.515 80.815 197.605 ;
        RECT 68.195 195.225 68.365 195.605 ;
        RECT 68.545 195.055 68.875 195.435 ;
        RECT 69.055 195.225 69.315 195.730 ;
        RECT 73.830 195.600 74.170 196.430 ;
        RECT 77.305 195.995 78.995 196.515 ;
        RECT 79.165 195.825 80.815 196.345 ;
        RECT 70.410 195.055 75.755 195.600 ;
        RECT 75.925 195.055 76.215 195.780 ;
        RECT 77.305 195.055 80.815 195.825 ;
        RECT 80.985 195.225 81.245 197.435 ;
        RECT 81.415 197.225 81.745 197.605 ;
        RECT 82.170 197.055 82.340 197.435 ;
        RECT 82.600 197.225 82.930 197.605 ;
        RECT 83.125 197.055 83.295 197.435 ;
        RECT 83.505 197.225 83.835 197.605 ;
        RECT 84.085 197.055 84.275 197.435 ;
        RECT 84.515 197.225 84.845 197.605 ;
        RECT 85.155 197.105 85.415 197.435 ;
        RECT 81.415 196.885 83.365 197.055 ;
        RECT 81.415 195.965 81.585 196.885 ;
        RECT 81.955 196.295 82.150 196.605 ;
        RECT 82.420 196.295 82.605 196.605 ;
        RECT 81.895 195.965 82.150 196.295 ;
        RECT 82.375 195.965 82.605 196.295 ;
        RECT 81.415 195.055 81.745 195.435 ;
        RECT 81.955 195.390 82.150 195.965 ;
        RECT 82.420 195.385 82.605 195.965 ;
        RECT 82.855 195.395 83.025 196.295 ;
        RECT 83.195 195.895 83.365 196.885 ;
        RECT 83.535 196.885 84.275 197.055 ;
        RECT 83.535 196.375 83.705 196.885 ;
        RECT 83.875 196.545 84.455 196.715 ;
        RECT 84.725 196.595 85.075 196.925 ;
        RECT 84.285 196.425 84.455 196.545 ;
        RECT 85.245 196.425 85.415 197.105 ;
        RECT 85.585 197.050 86.190 197.605 ;
        RECT 86.365 197.095 86.845 197.435 ;
        RECT 87.015 197.060 87.270 197.605 ;
        RECT 85.585 196.950 86.200 197.050 ;
        RECT 86.015 196.925 86.200 196.950 ;
        RECT 83.535 196.205 84.105 196.375 ;
        RECT 84.285 196.255 85.415 196.425 ;
        RECT 83.195 195.565 83.745 195.895 ;
        RECT 83.935 195.725 84.105 196.205 ;
        RECT 84.275 195.915 84.895 196.085 ;
        RECT 84.685 195.735 84.895 195.915 ;
        RECT 83.935 195.395 84.335 195.725 ;
        RECT 85.245 195.555 85.415 196.255 ;
        RECT 85.585 196.330 85.845 196.780 ;
        RECT 86.015 196.680 86.345 196.925 ;
        RECT 86.515 196.605 87.270 196.855 ;
        RECT 87.440 196.735 87.715 197.435 ;
        RECT 86.500 196.570 87.270 196.605 ;
        RECT 86.485 196.560 87.270 196.570 ;
        RECT 86.480 196.545 87.375 196.560 ;
        RECT 86.460 196.530 87.375 196.545 ;
        RECT 86.440 196.520 87.375 196.530 ;
        RECT 86.415 196.510 87.375 196.520 ;
        RECT 86.345 196.480 87.375 196.510 ;
        RECT 86.325 196.450 87.375 196.480 ;
        RECT 86.305 196.420 87.375 196.450 ;
        RECT 86.275 196.395 87.375 196.420 ;
        RECT 86.240 196.360 87.375 196.395 ;
        RECT 86.210 196.355 87.375 196.360 ;
        RECT 86.210 196.350 86.600 196.355 ;
        RECT 86.210 196.340 86.575 196.350 ;
        RECT 86.210 196.335 86.560 196.340 ;
        RECT 86.210 196.330 86.545 196.335 ;
        RECT 85.585 196.325 86.545 196.330 ;
        RECT 85.585 196.315 86.535 196.325 ;
        RECT 85.585 196.310 86.525 196.315 ;
        RECT 85.585 196.300 86.515 196.310 ;
        RECT 85.585 196.290 86.510 196.300 ;
        RECT 85.585 196.285 86.505 196.290 ;
        RECT 85.585 196.270 86.495 196.285 ;
        RECT 85.585 196.255 86.490 196.270 ;
        RECT 85.585 196.230 86.480 196.255 ;
        RECT 85.585 196.160 86.475 196.230 ;
        RECT 85.585 195.605 86.135 195.990 ;
        RECT 82.855 195.225 84.335 195.395 ;
        RECT 84.515 195.055 84.845 195.435 ;
        RECT 85.155 195.225 85.415 195.555 ;
        RECT 86.305 195.435 86.475 196.160 ;
        RECT 85.585 195.265 86.475 195.435 ;
        RECT 86.645 195.760 86.975 196.185 ;
        RECT 87.145 195.960 87.375 196.355 ;
        RECT 86.645 195.275 86.865 195.760 ;
        RECT 87.545 195.705 87.715 196.735 ;
        RECT 87.035 195.055 87.285 195.595 ;
        RECT 87.455 195.225 87.715 195.705 ;
        RECT 87.885 196.635 88.155 197.405 ;
        RECT 88.325 196.825 88.655 197.605 ;
        RECT 88.860 197.000 89.045 197.405 ;
        RECT 89.215 197.180 89.550 197.605 ;
        RECT 88.860 196.825 89.525 197.000 ;
        RECT 87.885 196.465 89.015 196.635 ;
        RECT 87.885 195.555 88.055 196.465 ;
        RECT 88.225 195.715 88.585 196.295 ;
        RECT 88.765 195.965 89.015 196.465 ;
        RECT 89.185 195.795 89.525 196.825 ;
        RECT 89.725 196.515 92.315 197.605 ;
        RECT 89.725 195.995 90.935 196.515 ;
        RECT 92.525 196.465 92.755 197.605 ;
        RECT 92.925 196.455 93.255 197.435 ;
        RECT 93.425 196.465 93.635 197.605 ;
        RECT 93.980 196.975 94.265 197.435 ;
        RECT 94.435 197.145 94.705 197.605 ;
        RECT 93.980 196.755 94.935 196.975 ;
        RECT 91.105 195.825 92.315 196.345 ;
        RECT 92.505 196.045 92.835 196.295 ;
        RECT 88.840 195.625 89.525 195.795 ;
        RECT 87.885 195.225 88.145 195.555 ;
        RECT 88.355 195.055 88.630 195.535 ;
        RECT 88.840 195.225 89.045 195.625 ;
        RECT 89.215 195.055 89.550 195.455 ;
        RECT 89.725 195.055 92.315 195.825 ;
        RECT 92.525 195.055 92.755 195.875 ;
        RECT 93.005 195.855 93.255 196.455 ;
        RECT 93.865 196.025 94.555 196.585 ;
        RECT 92.925 195.225 93.255 195.855 ;
        RECT 93.425 195.055 93.635 195.875 ;
        RECT 94.725 195.855 94.935 196.755 ;
        RECT 93.980 195.685 94.935 195.855 ;
        RECT 95.105 196.585 95.505 197.435 ;
        RECT 95.695 196.975 95.975 197.435 ;
        RECT 96.495 197.145 96.820 197.605 ;
        RECT 95.695 196.755 96.820 196.975 ;
        RECT 95.105 196.025 96.200 196.585 ;
        RECT 96.370 196.295 96.820 196.755 ;
        RECT 96.990 196.465 97.375 197.435 ;
        RECT 93.980 195.225 94.265 195.685 ;
        RECT 94.435 195.055 94.705 195.515 ;
        RECT 95.105 195.225 95.505 196.025 ;
        RECT 96.370 195.965 96.925 196.295 ;
        RECT 96.370 195.855 96.820 195.965 ;
        RECT 95.695 195.685 96.820 195.855 ;
        RECT 97.095 195.795 97.375 196.465 ;
        RECT 97.545 196.845 98.060 197.255 ;
        RECT 98.295 196.845 98.465 197.605 ;
        RECT 98.635 197.265 100.665 197.435 ;
        RECT 97.545 196.035 97.885 196.845 ;
        RECT 98.635 196.600 98.805 197.265 ;
        RECT 99.200 196.925 100.325 197.095 ;
        RECT 98.055 196.410 98.805 196.600 ;
        RECT 98.975 196.585 99.985 196.755 ;
        RECT 97.545 195.865 98.775 196.035 ;
        RECT 95.695 195.225 95.975 195.685 ;
        RECT 96.495 195.055 96.820 195.515 ;
        RECT 96.990 195.225 97.375 195.795 ;
        RECT 97.820 195.260 98.065 195.865 ;
        RECT 98.285 195.055 98.795 195.590 ;
        RECT 98.975 195.225 99.165 196.585 ;
        RECT 99.335 195.565 99.610 196.385 ;
        RECT 99.815 195.785 99.985 196.585 ;
        RECT 100.155 195.795 100.325 196.925 ;
        RECT 100.495 196.295 100.665 197.265 ;
        RECT 100.835 196.465 101.005 197.605 ;
        RECT 101.175 196.465 101.510 197.435 ;
        RECT 100.495 195.965 100.690 196.295 ;
        RECT 100.915 195.965 101.170 196.295 ;
        RECT 100.915 195.795 101.085 195.965 ;
        RECT 101.340 195.795 101.510 196.465 ;
        RECT 101.685 196.440 101.975 197.605 ;
        RECT 102.145 196.515 105.655 197.605 ;
        RECT 105.915 196.675 106.085 197.435 ;
        RECT 106.265 196.845 106.595 197.605 ;
        RECT 102.145 195.995 103.835 196.515 ;
        RECT 105.915 196.505 106.580 196.675 ;
        RECT 106.765 196.530 107.035 197.435 ;
        RECT 106.410 196.360 106.580 196.505 ;
        RECT 104.005 195.825 105.655 196.345 ;
        RECT 105.845 195.955 106.175 196.325 ;
        RECT 106.410 196.030 106.695 196.360 ;
        RECT 100.155 195.625 101.085 195.795 ;
        RECT 100.155 195.590 100.330 195.625 ;
        RECT 99.335 195.395 99.615 195.565 ;
        RECT 99.335 195.225 99.610 195.395 ;
        RECT 99.800 195.225 100.330 195.590 ;
        RECT 100.755 195.055 101.085 195.455 ;
        RECT 101.255 195.225 101.510 195.795 ;
        RECT 101.685 195.055 101.975 195.780 ;
        RECT 102.145 195.055 105.655 195.825 ;
        RECT 106.410 195.775 106.580 196.030 ;
        RECT 105.915 195.605 106.580 195.775 ;
        RECT 106.865 195.730 107.035 196.530 ;
        RECT 107.205 196.515 108.415 197.605 ;
        RECT 108.675 196.675 108.845 197.435 ;
        RECT 109.025 196.845 109.355 197.605 ;
        RECT 107.205 195.975 107.725 196.515 ;
        RECT 108.675 196.505 109.340 196.675 ;
        RECT 109.525 196.530 109.795 197.435 ;
        RECT 109.170 196.360 109.340 196.505 ;
        RECT 107.895 195.805 108.415 196.345 ;
        RECT 108.605 195.955 108.935 196.325 ;
        RECT 109.170 196.030 109.455 196.360 ;
        RECT 105.915 195.225 106.085 195.605 ;
        RECT 106.265 195.055 106.595 195.435 ;
        RECT 106.775 195.225 107.035 195.730 ;
        RECT 107.205 195.055 108.415 195.805 ;
        RECT 109.170 195.775 109.340 196.030 ;
        RECT 108.675 195.605 109.340 195.775 ;
        RECT 109.625 195.730 109.795 196.530 ;
        RECT 109.965 196.845 110.480 197.255 ;
        RECT 110.715 196.845 110.885 197.605 ;
        RECT 111.055 197.265 113.085 197.435 ;
        RECT 109.965 196.035 110.305 196.845 ;
        RECT 111.055 196.600 111.225 197.265 ;
        RECT 111.620 196.925 112.745 197.095 ;
        RECT 110.475 196.410 111.225 196.600 ;
        RECT 111.395 196.585 112.405 196.755 ;
        RECT 109.965 195.865 111.195 196.035 ;
        RECT 108.675 195.225 108.845 195.605 ;
        RECT 109.025 195.055 109.355 195.435 ;
        RECT 109.535 195.225 109.795 195.730 ;
        RECT 110.240 195.260 110.485 195.865 ;
        RECT 110.705 195.055 111.215 195.590 ;
        RECT 111.395 195.225 111.585 196.585 ;
        RECT 111.755 195.905 112.030 196.385 ;
        RECT 111.755 195.735 112.035 195.905 ;
        RECT 112.235 195.785 112.405 196.585 ;
        RECT 112.575 195.795 112.745 196.925 ;
        RECT 112.915 196.295 113.085 197.265 ;
        RECT 113.255 196.465 113.425 197.605 ;
        RECT 113.595 196.465 113.930 197.435 ;
        RECT 112.915 195.965 113.110 196.295 ;
        RECT 113.335 195.965 113.590 196.295 ;
        RECT 113.335 195.795 113.505 195.965 ;
        RECT 113.760 195.795 113.930 196.465 ;
        RECT 111.755 195.225 112.030 195.735 ;
        RECT 112.575 195.625 113.505 195.795 ;
        RECT 112.575 195.590 112.750 195.625 ;
        RECT 112.220 195.225 112.750 195.590 ;
        RECT 113.175 195.055 113.505 195.455 ;
        RECT 113.675 195.225 113.930 195.795 ;
        RECT 114.110 196.415 114.365 197.295 ;
        RECT 114.535 196.465 114.840 197.605 ;
        RECT 115.180 197.225 115.510 197.605 ;
        RECT 115.690 197.055 115.860 197.345 ;
        RECT 116.030 197.145 116.280 197.605 ;
        RECT 115.060 196.885 115.860 197.055 ;
        RECT 116.450 197.095 117.320 197.435 ;
        RECT 114.110 195.765 114.320 196.415 ;
        RECT 115.060 196.295 115.230 196.885 ;
        RECT 116.450 196.715 116.620 197.095 ;
        RECT 117.555 196.975 117.725 197.435 ;
        RECT 117.895 197.145 118.265 197.605 ;
        RECT 118.560 197.005 118.730 197.345 ;
        RECT 118.900 197.175 119.230 197.605 ;
        RECT 119.465 197.005 119.635 197.345 ;
        RECT 115.400 196.545 116.620 196.715 ;
        RECT 116.790 196.635 117.250 196.925 ;
        RECT 117.555 196.805 118.115 196.975 ;
        RECT 118.560 196.835 119.635 197.005 ;
        RECT 119.805 197.105 120.485 197.435 ;
        RECT 120.700 197.105 120.950 197.435 ;
        RECT 121.120 197.145 121.370 197.605 ;
        RECT 117.945 196.665 118.115 196.805 ;
        RECT 116.790 196.625 117.755 196.635 ;
        RECT 116.450 196.455 116.620 196.545 ;
        RECT 117.080 196.465 117.755 196.625 ;
        RECT 114.490 196.265 115.230 196.295 ;
        RECT 114.490 195.965 115.405 196.265 ;
        RECT 115.080 195.790 115.405 195.965 ;
        RECT 114.110 195.235 114.365 195.765 ;
        RECT 114.535 195.055 114.840 195.515 ;
        RECT 115.085 195.435 115.405 195.790 ;
        RECT 115.575 196.005 116.115 196.375 ;
        RECT 116.450 196.285 116.855 196.455 ;
        RECT 115.575 195.605 115.815 196.005 ;
        RECT 116.295 195.835 116.515 196.115 ;
        RECT 115.985 195.665 116.515 195.835 ;
        RECT 115.985 195.435 116.155 195.665 ;
        RECT 116.685 195.505 116.855 196.285 ;
        RECT 117.025 195.675 117.375 196.295 ;
        RECT 117.545 195.675 117.755 196.465 ;
        RECT 117.945 196.495 119.445 196.665 ;
        RECT 117.945 195.805 118.115 196.495 ;
        RECT 119.805 196.325 119.975 197.105 ;
        RECT 120.780 196.975 120.950 197.105 ;
        RECT 118.285 196.155 119.975 196.325 ;
        RECT 120.145 196.545 120.610 196.935 ;
        RECT 120.780 196.805 121.175 196.975 ;
        RECT 118.285 195.975 118.455 196.155 ;
        RECT 115.085 195.265 116.155 195.435 ;
        RECT 116.325 195.055 116.515 195.495 ;
        RECT 116.685 195.225 117.635 195.505 ;
        RECT 117.945 195.415 118.205 195.805 ;
        RECT 118.625 195.735 119.415 195.985 ;
        RECT 117.855 195.245 118.205 195.415 ;
        RECT 118.415 195.055 118.745 195.515 ;
        RECT 119.620 195.445 119.790 196.155 ;
        RECT 120.145 195.955 120.315 196.545 ;
        RECT 119.960 195.735 120.315 195.955 ;
        RECT 120.485 195.735 120.835 196.355 ;
        RECT 121.005 195.445 121.175 196.805 ;
        RECT 121.540 196.635 121.865 197.420 ;
        RECT 121.345 195.585 121.805 196.635 ;
        RECT 119.620 195.275 120.475 195.445 ;
        RECT 120.680 195.275 121.175 195.445 ;
        RECT 121.345 195.055 121.675 195.415 ;
        RECT 122.035 195.315 122.205 197.435 ;
        RECT 122.375 197.105 122.705 197.605 ;
        RECT 122.875 196.935 123.130 197.435 ;
        RECT 122.380 196.765 123.130 196.935 ;
        RECT 122.380 195.775 122.610 196.765 ;
        RECT 122.780 195.945 123.130 196.595 ;
        RECT 123.765 196.515 126.355 197.605 ;
        RECT 126.525 196.515 127.735 197.605 ;
        RECT 123.765 195.995 124.975 196.515 ;
        RECT 125.145 195.825 126.355 196.345 ;
        RECT 126.525 195.975 127.045 196.515 ;
        RECT 122.380 195.605 123.130 195.775 ;
        RECT 122.375 195.055 122.705 195.435 ;
        RECT 122.875 195.315 123.130 195.605 ;
        RECT 123.765 195.055 126.355 195.825 ;
        RECT 127.215 195.805 127.735 196.345 ;
        RECT 126.525 195.055 127.735 195.805 ;
        RECT 29.840 194.885 127.820 195.055 ;
        RECT 29.925 194.135 31.135 194.885 ;
        RECT 31.770 194.340 37.115 194.885 ;
        RECT 29.925 193.595 30.445 194.135 ;
        RECT 30.615 193.425 31.135 193.965 ;
        RECT 29.925 192.335 31.135 193.425 ;
        RECT 33.360 192.770 33.710 194.020 ;
        RECT 35.190 193.510 35.530 194.340 ;
        RECT 37.285 194.160 37.575 194.885 ;
        RECT 37.750 194.340 43.095 194.885 ;
        RECT 31.770 192.335 37.115 192.770 ;
        RECT 37.285 192.335 37.575 193.500 ;
        RECT 39.340 192.770 39.690 194.020 ;
        RECT 41.170 193.510 41.510 194.340 ;
        RECT 43.305 194.065 43.535 194.885 ;
        RECT 43.705 194.085 44.035 194.715 ;
        RECT 43.285 193.645 43.615 193.895 ;
        RECT 43.785 193.485 44.035 194.085 ;
        RECT 44.205 194.065 44.415 194.885 ;
        RECT 44.650 194.335 44.905 194.625 ;
        RECT 45.075 194.505 45.405 194.885 ;
        RECT 44.650 194.165 45.400 194.335 ;
        RECT 37.750 192.335 43.095 192.770 ;
        RECT 43.305 192.335 43.535 193.475 ;
        RECT 43.705 192.505 44.035 193.485 ;
        RECT 44.205 192.335 44.415 193.475 ;
        RECT 44.650 193.345 45.000 193.995 ;
        RECT 45.170 193.175 45.400 194.165 ;
        RECT 44.650 193.005 45.400 193.175 ;
        RECT 44.650 192.505 44.905 193.005 ;
        RECT 45.075 192.335 45.405 192.835 ;
        RECT 45.575 192.505 45.745 194.625 ;
        RECT 46.105 194.525 46.435 194.885 ;
        RECT 46.605 194.495 47.100 194.665 ;
        RECT 47.305 194.495 48.160 194.665 ;
        RECT 45.975 193.305 46.435 194.355 ;
        RECT 45.915 192.520 46.240 193.305 ;
        RECT 46.605 193.135 46.775 194.495 ;
        RECT 46.945 193.585 47.295 194.205 ;
        RECT 47.465 193.985 47.820 194.205 ;
        RECT 47.465 193.395 47.635 193.985 ;
        RECT 47.990 193.785 48.160 194.495 ;
        RECT 49.035 194.425 49.365 194.885 ;
        RECT 49.575 194.525 49.925 194.695 ;
        RECT 48.365 193.955 49.155 194.205 ;
        RECT 49.575 194.135 49.835 194.525 ;
        RECT 50.145 194.435 51.095 194.715 ;
        RECT 51.265 194.445 51.455 194.885 ;
        RECT 51.625 194.505 52.695 194.675 ;
        RECT 49.325 193.785 49.495 193.965 ;
        RECT 46.605 192.965 47.000 193.135 ;
        RECT 47.170 193.005 47.635 193.395 ;
        RECT 47.805 193.615 49.495 193.785 ;
        RECT 46.830 192.835 47.000 192.965 ;
        RECT 47.805 192.835 47.975 193.615 ;
        RECT 49.665 193.445 49.835 194.135 ;
        RECT 48.335 193.275 49.835 193.445 ;
        RECT 50.025 193.475 50.235 194.265 ;
        RECT 50.405 193.645 50.755 194.265 ;
        RECT 50.925 193.655 51.095 194.435 ;
        RECT 51.625 194.275 51.795 194.505 ;
        RECT 51.265 194.105 51.795 194.275 ;
        RECT 51.265 193.825 51.485 194.105 ;
        RECT 51.965 193.935 52.205 194.335 ;
        RECT 50.925 193.485 51.330 193.655 ;
        RECT 51.665 193.565 52.205 193.935 ;
        RECT 52.375 194.150 52.695 194.505 ;
        RECT 52.940 194.425 53.245 194.885 ;
        RECT 53.415 194.175 53.670 194.705 ;
        RECT 52.375 193.975 52.700 194.150 ;
        RECT 52.375 193.675 53.290 193.975 ;
        RECT 52.550 193.645 53.290 193.675 ;
        RECT 50.025 193.315 50.700 193.475 ;
        RECT 51.160 193.395 51.330 193.485 ;
        RECT 50.025 193.305 50.990 193.315 ;
        RECT 49.665 193.135 49.835 193.275 ;
        RECT 46.410 192.335 46.660 192.795 ;
        RECT 46.830 192.505 47.080 192.835 ;
        RECT 47.295 192.505 47.975 192.835 ;
        RECT 48.145 192.935 49.220 193.105 ;
        RECT 49.665 192.965 50.225 193.135 ;
        RECT 50.530 193.015 50.990 193.305 ;
        RECT 51.160 193.225 52.380 193.395 ;
        RECT 48.145 192.595 48.315 192.935 ;
        RECT 48.550 192.335 48.880 192.765 ;
        RECT 49.050 192.595 49.220 192.935 ;
        RECT 49.515 192.335 49.885 192.795 ;
        RECT 50.055 192.505 50.225 192.965 ;
        RECT 51.160 192.845 51.330 193.225 ;
        RECT 52.550 193.055 52.720 193.645 ;
        RECT 53.460 193.525 53.670 194.175 ;
        RECT 50.460 192.505 51.330 192.845 ;
        RECT 51.920 192.885 52.720 193.055 ;
        RECT 51.500 192.335 51.750 192.795 ;
        RECT 51.920 192.595 52.090 192.885 ;
        RECT 52.270 192.335 52.600 192.715 ;
        RECT 52.940 192.335 53.245 193.475 ;
        RECT 53.415 192.645 53.670 193.525 ;
        RECT 53.850 194.175 54.105 194.705 ;
        RECT 54.275 194.425 54.580 194.885 ;
        RECT 54.825 194.505 55.895 194.675 ;
        RECT 53.850 193.525 54.060 194.175 ;
        RECT 54.825 194.150 55.145 194.505 ;
        RECT 54.820 193.975 55.145 194.150 ;
        RECT 54.230 193.675 55.145 193.975 ;
        RECT 55.315 193.935 55.555 194.335 ;
        RECT 55.725 194.275 55.895 194.505 ;
        RECT 56.065 194.445 56.255 194.885 ;
        RECT 56.425 194.435 57.375 194.715 ;
        RECT 57.595 194.525 57.945 194.695 ;
        RECT 55.725 194.105 56.255 194.275 ;
        RECT 54.230 193.645 54.970 193.675 ;
        RECT 53.850 192.645 54.105 193.525 ;
        RECT 54.275 192.335 54.580 193.475 ;
        RECT 54.800 193.055 54.970 193.645 ;
        RECT 55.315 193.565 55.855 193.935 ;
        RECT 56.035 193.825 56.255 194.105 ;
        RECT 56.425 193.655 56.595 194.435 ;
        RECT 56.190 193.485 56.595 193.655 ;
        RECT 56.765 193.645 57.115 194.265 ;
        RECT 56.190 193.395 56.360 193.485 ;
        RECT 57.285 193.475 57.495 194.265 ;
        RECT 55.140 193.225 56.360 193.395 ;
        RECT 56.820 193.315 57.495 193.475 ;
        RECT 54.800 192.885 55.600 193.055 ;
        RECT 54.920 192.335 55.250 192.715 ;
        RECT 55.430 192.595 55.600 192.885 ;
        RECT 56.190 192.845 56.360 193.225 ;
        RECT 56.530 193.305 57.495 193.315 ;
        RECT 57.685 194.135 57.945 194.525 ;
        RECT 58.155 194.425 58.485 194.885 ;
        RECT 59.360 194.495 60.215 194.665 ;
        RECT 60.420 194.495 60.915 194.665 ;
        RECT 61.085 194.525 61.415 194.885 ;
        RECT 57.685 193.445 57.855 194.135 ;
        RECT 58.025 193.785 58.195 193.965 ;
        RECT 58.365 193.955 59.155 194.205 ;
        RECT 59.360 193.785 59.530 194.495 ;
        RECT 59.700 193.985 60.055 194.205 ;
        RECT 58.025 193.615 59.715 193.785 ;
        RECT 56.530 193.015 56.990 193.305 ;
        RECT 57.685 193.275 59.185 193.445 ;
        RECT 57.685 193.135 57.855 193.275 ;
        RECT 57.295 192.965 57.855 193.135 ;
        RECT 55.770 192.335 56.020 192.795 ;
        RECT 56.190 192.505 57.060 192.845 ;
        RECT 57.295 192.505 57.465 192.965 ;
        RECT 58.300 192.935 59.375 193.105 ;
        RECT 57.635 192.335 58.005 192.795 ;
        RECT 58.300 192.595 58.470 192.935 ;
        RECT 58.640 192.335 58.970 192.765 ;
        RECT 59.205 192.595 59.375 192.935 ;
        RECT 59.545 192.835 59.715 193.615 ;
        RECT 59.885 193.395 60.055 193.985 ;
        RECT 60.225 193.585 60.575 194.205 ;
        RECT 59.885 193.005 60.350 193.395 ;
        RECT 60.745 193.135 60.915 194.495 ;
        RECT 61.085 193.305 61.545 194.355 ;
        RECT 60.520 192.965 60.915 193.135 ;
        RECT 60.520 192.835 60.690 192.965 ;
        RECT 59.545 192.505 60.225 192.835 ;
        RECT 60.440 192.505 60.690 192.835 ;
        RECT 60.860 192.335 61.110 192.795 ;
        RECT 61.280 192.520 61.605 193.305 ;
        RECT 61.775 192.505 61.945 194.625 ;
        RECT 62.115 194.505 62.445 194.885 ;
        RECT 62.615 194.335 62.870 194.625 ;
        RECT 62.120 194.165 62.870 194.335 ;
        RECT 62.120 193.175 62.350 194.165 ;
        RECT 63.045 194.160 63.335 194.885 ;
        RECT 63.510 194.175 63.765 194.705 ;
        RECT 63.935 194.425 64.240 194.885 ;
        RECT 64.485 194.505 65.555 194.675 ;
        RECT 62.520 193.345 62.870 193.995 ;
        RECT 63.510 193.525 63.720 194.175 ;
        RECT 64.485 194.150 64.805 194.505 ;
        RECT 64.480 193.975 64.805 194.150 ;
        RECT 63.890 193.675 64.805 193.975 ;
        RECT 64.975 193.935 65.215 194.335 ;
        RECT 65.385 194.275 65.555 194.505 ;
        RECT 65.725 194.445 65.915 194.885 ;
        RECT 66.085 194.435 67.035 194.715 ;
        RECT 67.255 194.525 67.605 194.695 ;
        RECT 65.385 194.105 65.915 194.275 ;
        RECT 63.890 193.645 64.630 193.675 ;
        RECT 62.120 193.005 62.870 193.175 ;
        RECT 62.115 192.335 62.445 192.835 ;
        RECT 62.615 192.505 62.870 193.005 ;
        RECT 63.045 192.335 63.335 193.500 ;
        RECT 63.510 192.645 63.765 193.525 ;
        RECT 63.935 192.335 64.240 193.475 ;
        RECT 64.460 193.055 64.630 193.645 ;
        RECT 64.975 193.565 65.515 193.935 ;
        RECT 65.695 193.825 65.915 194.105 ;
        RECT 66.085 193.655 66.255 194.435 ;
        RECT 65.850 193.485 66.255 193.655 ;
        RECT 66.425 193.645 66.775 194.265 ;
        RECT 65.850 193.395 66.020 193.485 ;
        RECT 66.945 193.475 67.155 194.265 ;
        RECT 64.800 193.225 66.020 193.395 ;
        RECT 66.480 193.315 67.155 193.475 ;
        RECT 64.460 192.885 65.260 193.055 ;
        RECT 64.580 192.335 64.910 192.715 ;
        RECT 65.090 192.595 65.260 192.885 ;
        RECT 65.850 192.845 66.020 193.225 ;
        RECT 66.190 193.305 67.155 193.315 ;
        RECT 67.345 194.135 67.605 194.525 ;
        RECT 67.815 194.425 68.145 194.885 ;
        RECT 69.020 194.495 69.875 194.665 ;
        RECT 70.080 194.495 70.575 194.665 ;
        RECT 70.745 194.525 71.075 194.885 ;
        RECT 67.345 193.445 67.515 194.135 ;
        RECT 67.685 193.785 67.855 193.965 ;
        RECT 68.025 193.955 68.815 194.205 ;
        RECT 69.020 193.785 69.190 194.495 ;
        RECT 69.360 193.985 69.715 194.205 ;
        RECT 67.685 193.615 69.375 193.785 ;
        RECT 66.190 193.015 66.650 193.305 ;
        RECT 67.345 193.275 68.845 193.445 ;
        RECT 67.345 193.135 67.515 193.275 ;
        RECT 66.955 192.965 67.515 193.135 ;
        RECT 65.430 192.335 65.680 192.795 ;
        RECT 65.850 192.505 66.720 192.845 ;
        RECT 66.955 192.505 67.125 192.965 ;
        RECT 67.960 192.935 69.035 193.105 ;
        RECT 67.295 192.335 67.665 192.795 ;
        RECT 67.960 192.595 68.130 192.935 ;
        RECT 68.300 192.335 68.630 192.765 ;
        RECT 68.865 192.595 69.035 192.935 ;
        RECT 69.205 192.835 69.375 193.615 ;
        RECT 69.545 193.395 69.715 193.985 ;
        RECT 69.885 193.585 70.235 194.205 ;
        RECT 69.545 193.005 70.010 193.395 ;
        RECT 70.405 193.135 70.575 194.495 ;
        RECT 70.745 193.305 71.205 194.355 ;
        RECT 70.180 192.965 70.575 193.135 ;
        RECT 70.180 192.835 70.350 192.965 ;
        RECT 69.205 192.505 69.885 192.835 ;
        RECT 70.100 192.505 70.350 192.835 ;
        RECT 70.520 192.335 70.770 192.795 ;
        RECT 70.940 192.520 71.265 193.305 ;
        RECT 71.435 192.505 71.605 194.625 ;
        RECT 71.775 194.505 72.105 194.885 ;
        RECT 72.275 194.335 72.530 194.625 ;
        RECT 71.780 194.165 72.530 194.335 ;
        RECT 73.715 194.335 73.885 194.715 ;
        RECT 74.100 194.505 74.430 194.885 ;
        RECT 73.715 194.165 74.430 194.335 ;
        RECT 71.780 193.175 72.010 194.165 ;
        RECT 72.180 193.345 72.530 193.995 ;
        RECT 73.625 193.615 73.980 193.985 ;
        RECT 74.260 193.975 74.430 194.165 ;
        RECT 74.600 194.140 74.855 194.715 ;
        RECT 74.260 193.645 74.515 193.975 ;
        RECT 74.260 193.435 74.430 193.645 ;
        RECT 73.715 193.265 74.430 193.435 ;
        RECT 74.685 193.410 74.855 194.140 ;
        RECT 75.030 194.045 75.290 194.885 ;
        RECT 75.735 194.490 76.065 194.885 ;
        RECT 76.235 194.315 76.435 194.670 ;
        RECT 76.605 194.485 76.935 194.885 ;
        RECT 77.105 194.315 77.305 194.660 ;
        RECT 75.465 194.145 77.305 194.315 ;
        RECT 77.475 194.145 77.805 194.885 ;
        RECT 78.040 194.315 78.210 194.565 ;
        RECT 78.955 194.490 79.285 194.885 ;
        RECT 79.455 194.315 79.655 194.670 ;
        RECT 79.825 194.485 80.155 194.885 ;
        RECT 80.325 194.315 80.525 194.660 ;
        RECT 78.040 194.145 78.515 194.315 ;
        RECT 71.780 193.005 72.530 193.175 ;
        RECT 71.775 192.335 72.105 192.835 ;
        RECT 72.275 192.505 72.530 193.005 ;
        RECT 73.715 192.505 73.885 193.265 ;
        RECT 74.100 192.335 74.430 193.095 ;
        RECT 74.600 192.505 74.855 193.410 ;
        RECT 75.030 192.335 75.290 193.485 ;
        RECT 75.465 192.520 75.725 194.145 ;
        RECT 75.905 193.175 76.125 193.975 ;
        RECT 76.365 193.355 76.665 193.975 ;
        RECT 76.835 193.355 77.165 193.975 ;
        RECT 77.335 193.355 77.655 193.975 ;
        RECT 77.825 193.355 78.175 193.975 ;
        RECT 78.345 193.175 78.515 194.145 ;
        RECT 75.905 192.965 78.515 193.175 ;
        RECT 78.685 194.145 80.525 194.315 ;
        RECT 80.695 194.145 81.025 194.885 ;
        RECT 81.260 194.315 81.430 194.565 ;
        RECT 82.175 194.490 82.505 194.885 ;
        RECT 82.675 194.315 82.875 194.670 ;
        RECT 83.045 194.485 83.375 194.885 ;
        RECT 83.545 194.315 83.745 194.660 ;
        RECT 81.260 194.145 81.735 194.315 ;
        RECT 77.475 192.335 77.805 192.785 ;
        RECT 78.685 192.520 78.945 194.145 ;
        RECT 79.125 193.175 79.345 193.975 ;
        RECT 79.585 193.355 79.885 193.975 ;
        RECT 80.055 193.355 80.385 193.975 ;
        RECT 80.555 193.355 80.875 193.975 ;
        RECT 81.045 193.355 81.395 193.975 ;
        RECT 81.565 193.175 81.735 194.145 ;
        RECT 79.125 192.965 81.735 193.175 ;
        RECT 81.905 194.145 83.745 194.315 ;
        RECT 83.915 194.145 84.245 194.885 ;
        RECT 84.480 194.315 84.650 194.565 ;
        RECT 84.480 194.145 84.955 194.315 ;
        RECT 80.695 192.335 81.025 192.785 ;
        RECT 81.905 192.520 82.165 194.145 ;
        RECT 82.345 193.175 82.565 193.975 ;
        RECT 82.805 193.355 83.105 193.975 ;
        RECT 83.275 193.355 83.605 193.975 ;
        RECT 83.775 193.355 84.095 193.975 ;
        RECT 84.265 193.355 84.615 193.975 ;
        RECT 84.785 193.175 84.955 194.145 ;
        RECT 85.125 194.115 88.635 194.885 ;
        RECT 88.805 194.160 89.095 194.885 ;
        RECT 82.345 192.965 84.955 193.175 ;
        RECT 85.125 193.425 86.815 193.945 ;
        RECT 86.985 193.595 88.635 194.115 ;
        RECT 89.305 194.065 89.535 194.885 ;
        RECT 89.705 194.085 90.035 194.715 ;
        RECT 89.285 193.645 89.615 193.895 ;
        RECT 83.915 192.335 84.245 192.785 ;
        RECT 85.125 192.335 88.635 193.425 ;
        RECT 88.805 192.335 89.095 193.500 ;
        RECT 89.785 193.485 90.035 194.085 ;
        RECT 90.205 194.065 90.415 194.885 ;
        RECT 91.020 194.175 91.275 194.705 ;
        RECT 91.455 194.425 91.740 194.885 ;
        RECT 89.305 192.335 89.535 193.475 ;
        RECT 89.705 192.505 90.035 193.485 ;
        RECT 90.205 192.335 90.415 193.475 ;
        RECT 91.020 193.315 91.200 194.175 ;
        RECT 91.920 193.975 92.170 194.625 ;
        RECT 91.370 193.645 92.170 193.975 ;
        RECT 91.020 193.185 91.275 193.315 ;
        RECT 90.935 193.015 91.275 193.185 ;
        RECT 91.020 192.645 91.275 193.015 ;
        RECT 91.455 192.335 91.740 193.135 ;
        RECT 91.920 193.055 92.170 193.645 ;
        RECT 92.370 194.290 92.690 194.620 ;
        RECT 92.870 194.405 93.530 194.885 ;
        RECT 93.730 194.495 94.580 194.665 ;
        RECT 92.370 193.395 92.560 194.290 ;
        RECT 92.880 193.965 93.540 194.235 ;
        RECT 93.210 193.905 93.540 193.965 ;
        RECT 92.730 193.735 93.060 193.795 ;
        RECT 93.730 193.735 93.900 194.495 ;
        RECT 95.140 194.425 95.460 194.885 ;
        RECT 95.660 194.245 95.910 194.675 ;
        RECT 96.200 194.445 96.610 194.885 ;
        RECT 96.780 194.505 97.795 194.705 ;
        RECT 94.070 194.075 95.320 194.245 ;
        RECT 94.070 193.955 94.400 194.075 ;
        RECT 92.730 193.565 94.630 193.735 ;
        RECT 92.370 193.225 94.290 193.395 ;
        RECT 92.370 193.205 92.690 193.225 ;
        RECT 91.920 192.545 92.250 193.055 ;
        RECT 92.520 192.595 92.690 193.205 ;
        RECT 94.460 193.055 94.630 193.565 ;
        RECT 94.800 193.495 94.980 193.905 ;
        RECT 95.150 193.315 95.320 194.075 ;
        RECT 92.860 192.335 93.190 193.025 ;
        RECT 93.420 192.885 94.630 193.055 ;
        RECT 94.800 193.005 95.320 193.315 ;
        RECT 95.490 193.905 95.910 194.245 ;
        RECT 96.200 193.905 96.610 194.235 ;
        RECT 95.490 193.135 95.680 193.905 ;
        RECT 96.780 193.775 96.950 194.505 ;
        RECT 98.095 194.335 98.265 194.665 ;
        RECT 98.435 194.505 98.765 194.885 ;
        RECT 97.120 193.955 97.470 194.325 ;
        RECT 96.780 193.735 97.200 193.775 ;
        RECT 95.850 193.565 97.200 193.735 ;
        RECT 95.850 193.405 96.100 193.565 ;
        RECT 96.610 193.135 96.860 193.395 ;
        RECT 95.490 192.885 96.860 193.135 ;
        RECT 93.420 192.595 93.660 192.885 ;
        RECT 94.460 192.805 94.630 192.885 ;
        RECT 93.860 192.335 94.280 192.715 ;
        RECT 94.460 192.555 95.090 192.805 ;
        RECT 95.560 192.335 95.890 192.715 ;
        RECT 96.060 192.595 96.230 192.885 ;
        RECT 97.030 192.720 97.200 193.565 ;
        RECT 97.650 193.395 97.870 194.265 ;
        RECT 98.095 194.145 98.790 194.335 ;
        RECT 97.370 193.015 97.870 193.395 ;
        RECT 98.040 193.345 98.450 193.965 ;
        RECT 98.620 193.175 98.790 194.145 ;
        RECT 98.095 193.005 98.790 193.175 ;
        RECT 96.410 192.335 96.790 192.715 ;
        RECT 97.030 192.550 97.860 192.720 ;
        RECT 98.095 192.505 98.265 193.005 ;
        RECT 98.435 192.335 98.765 192.835 ;
        RECT 98.980 192.505 99.205 194.625 ;
        RECT 99.375 194.505 99.705 194.885 ;
        RECT 99.875 194.335 100.045 194.625 ;
        RECT 99.380 194.165 100.045 194.335 ;
        RECT 99.380 193.175 99.610 194.165 ;
        RECT 100.765 194.115 104.275 194.885 ;
        RECT 99.780 193.345 100.130 193.995 ;
        RECT 100.765 193.425 102.455 193.945 ;
        RECT 102.625 193.595 104.275 194.115 ;
        RECT 104.485 194.065 104.715 194.885 ;
        RECT 104.885 194.085 105.215 194.715 ;
        RECT 104.465 193.645 104.795 193.895 ;
        RECT 104.965 193.485 105.215 194.085 ;
        RECT 105.385 194.065 105.595 194.885 ;
        RECT 105.940 194.255 106.225 194.715 ;
        RECT 106.395 194.425 106.665 194.885 ;
        RECT 105.940 194.085 106.895 194.255 ;
        RECT 99.380 193.005 100.045 193.175 ;
        RECT 99.375 192.335 99.705 192.835 ;
        RECT 99.875 192.505 100.045 193.005 ;
        RECT 100.765 192.335 104.275 193.425 ;
        RECT 104.485 192.335 104.715 193.475 ;
        RECT 104.885 192.505 105.215 193.485 ;
        RECT 105.385 192.335 105.595 193.475 ;
        RECT 105.825 193.355 106.515 193.915 ;
        RECT 106.685 193.185 106.895 194.085 ;
        RECT 105.940 192.965 106.895 193.185 ;
        RECT 107.065 193.915 107.465 194.715 ;
        RECT 107.655 194.255 107.935 194.715 ;
        RECT 108.455 194.425 108.780 194.885 ;
        RECT 107.655 194.085 108.780 194.255 ;
        RECT 108.950 194.145 109.335 194.715 ;
        RECT 108.330 193.975 108.780 194.085 ;
        RECT 107.065 193.355 108.160 193.915 ;
        RECT 108.330 193.645 108.885 193.975 ;
        RECT 105.940 192.505 106.225 192.965 ;
        RECT 106.395 192.335 106.665 192.795 ;
        RECT 107.065 192.505 107.465 193.355 ;
        RECT 108.330 193.185 108.780 193.645 ;
        RECT 109.055 193.475 109.335 194.145 ;
        RECT 107.655 192.965 108.780 193.185 ;
        RECT 107.655 192.505 107.935 192.965 ;
        RECT 108.455 192.335 108.780 192.795 ;
        RECT 108.950 192.505 109.335 193.475 ;
        RECT 109.505 194.145 109.890 194.715 ;
        RECT 110.060 194.425 110.385 194.885 ;
        RECT 110.905 194.255 111.185 194.715 ;
        RECT 109.505 193.475 109.785 194.145 ;
        RECT 110.060 194.085 111.185 194.255 ;
        RECT 110.060 193.975 110.510 194.085 ;
        RECT 109.955 193.645 110.510 193.975 ;
        RECT 111.375 193.915 111.775 194.715 ;
        RECT 112.175 194.425 112.445 194.885 ;
        RECT 112.615 194.255 112.900 194.715 ;
        RECT 109.505 192.505 109.890 193.475 ;
        RECT 110.060 193.185 110.510 193.645 ;
        RECT 110.680 193.355 111.775 193.915 ;
        RECT 110.060 192.965 111.185 193.185 ;
        RECT 110.060 192.335 110.385 192.795 ;
        RECT 110.905 192.505 111.185 192.965 ;
        RECT 111.375 192.505 111.775 193.355 ;
        RECT 111.945 194.085 112.900 194.255 ;
        RECT 113.275 194.335 113.445 194.715 ;
        RECT 113.625 194.505 113.955 194.885 ;
        RECT 113.275 194.165 113.940 194.335 ;
        RECT 114.135 194.210 114.395 194.715 ;
        RECT 111.945 193.185 112.155 194.085 ;
        RECT 112.325 193.355 113.015 193.915 ;
        RECT 113.205 193.615 113.535 193.985 ;
        RECT 113.770 193.910 113.940 194.165 ;
        RECT 113.770 193.580 114.055 193.910 ;
        RECT 113.770 193.435 113.940 193.580 ;
        RECT 113.275 193.265 113.940 193.435 ;
        RECT 114.225 193.410 114.395 194.210 ;
        RECT 114.565 194.160 114.855 194.885 ;
        RECT 115.025 194.145 115.410 194.715 ;
        RECT 115.580 194.425 115.905 194.885 ;
        RECT 116.425 194.255 116.705 194.715 ;
        RECT 111.945 192.965 112.900 193.185 ;
        RECT 112.175 192.335 112.445 192.795 ;
        RECT 112.615 192.505 112.900 192.965 ;
        RECT 113.275 192.505 113.445 193.265 ;
        RECT 113.625 192.335 113.955 193.095 ;
        RECT 114.125 192.505 114.395 193.410 ;
        RECT 114.565 192.335 114.855 193.500 ;
        RECT 115.025 193.475 115.305 194.145 ;
        RECT 115.580 194.085 116.705 194.255 ;
        RECT 115.580 193.975 116.030 194.085 ;
        RECT 115.475 193.645 116.030 193.975 ;
        RECT 116.895 193.915 117.295 194.715 ;
        RECT 117.695 194.425 117.965 194.885 ;
        RECT 118.135 194.255 118.420 194.715 ;
        RECT 115.025 192.505 115.410 193.475 ;
        RECT 115.580 193.185 116.030 193.645 ;
        RECT 116.200 193.355 117.295 193.915 ;
        RECT 115.580 192.965 116.705 193.185 ;
        RECT 115.580 192.335 115.905 192.795 ;
        RECT 116.425 192.505 116.705 192.965 ;
        RECT 116.895 192.505 117.295 193.355 ;
        RECT 117.465 194.085 118.420 194.255 ;
        RECT 119.165 194.115 120.835 194.885 ;
        RECT 121.010 194.340 126.355 194.885 ;
        RECT 117.465 193.185 117.675 194.085 ;
        RECT 117.845 193.355 118.535 193.915 ;
        RECT 119.165 193.425 119.915 193.945 ;
        RECT 120.085 193.595 120.835 194.115 ;
        RECT 117.465 192.965 118.420 193.185 ;
        RECT 117.695 192.335 117.965 192.795 ;
        RECT 118.135 192.505 118.420 192.965 ;
        RECT 119.165 192.335 120.835 193.425 ;
        RECT 122.600 192.770 122.950 194.020 ;
        RECT 124.430 193.510 124.770 194.340 ;
        RECT 126.525 194.135 127.735 194.885 ;
        RECT 126.525 193.425 127.045 193.965 ;
        RECT 127.215 193.595 127.735 194.135 ;
        RECT 121.010 192.335 126.355 192.770 ;
        RECT 126.525 192.335 127.735 193.425 ;
        RECT 29.840 192.165 127.820 192.335 ;
        RECT 29.925 191.075 31.135 192.165 ;
        RECT 31.310 191.730 36.655 192.165 ;
        RECT 29.925 190.365 30.445 190.905 ;
        RECT 30.615 190.535 31.135 191.075 ;
        RECT 32.900 190.480 33.250 191.730 ;
        RECT 36.940 191.535 37.225 191.995 ;
        RECT 37.395 191.705 37.665 192.165 ;
        RECT 36.940 191.315 37.895 191.535 ;
        RECT 29.925 189.615 31.135 190.365 ;
        RECT 34.730 190.160 35.070 190.990 ;
        RECT 36.825 190.585 37.515 191.145 ;
        RECT 37.685 190.415 37.895 191.315 ;
        RECT 36.940 190.245 37.895 190.415 ;
        RECT 38.065 191.145 38.465 191.995 ;
        RECT 38.655 191.535 38.935 191.995 ;
        RECT 39.455 191.705 39.780 192.165 ;
        RECT 38.655 191.315 39.780 191.535 ;
        RECT 38.065 190.585 39.160 191.145 ;
        RECT 39.330 190.855 39.780 191.315 ;
        RECT 39.950 191.025 40.335 191.995 ;
        RECT 31.310 189.615 36.655 190.160 ;
        RECT 36.940 189.785 37.225 190.245 ;
        RECT 37.395 189.615 37.665 190.075 ;
        RECT 38.065 189.785 38.465 190.585 ;
        RECT 39.330 190.525 39.885 190.855 ;
        RECT 39.330 190.415 39.780 190.525 ;
        RECT 38.655 190.245 39.780 190.415 ;
        RECT 40.055 190.355 40.335 191.025 ;
        RECT 40.880 191.185 41.135 191.855 ;
        RECT 41.315 191.365 41.600 192.165 ;
        RECT 41.780 191.445 42.110 191.955 ;
        RECT 40.880 190.465 41.060 191.185 ;
        RECT 41.780 190.855 42.030 191.445 ;
        RECT 42.380 191.295 42.550 191.905 ;
        RECT 42.720 191.475 43.050 192.165 ;
        RECT 43.280 191.615 43.520 191.905 ;
        RECT 43.720 191.785 44.140 192.165 ;
        RECT 44.320 191.695 44.950 191.945 ;
        RECT 45.420 191.785 45.750 192.165 ;
        RECT 44.320 191.615 44.490 191.695 ;
        RECT 45.920 191.615 46.090 191.905 ;
        RECT 46.270 191.785 46.650 192.165 ;
        RECT 46.890 191.780 47.720 191.950 ;
        RECT 43.280 191.445 44.490 191.615 ;
        RECT 41.230 190.525 42.030 190.855 ;
        RECT 38.655 189.785 38.935 190.245 ;
        RECT 39.455 189.615 39.780 190.075 ;
        RECT 39.950 189.785 40.335 190.355 ;
        RECT 40.795 190.325 41.060 190.465 ;
        RECT 40.795 190.295 41.135 190.325 ;
        RECT 40.880 189.795 41.135 190.295 ;
        RECT 41.315 189.615 41.600 190.075 ;
        RECT 41.780 189.875 42.030 190.525 ;
        RECT 42.230 191.275 42.550 191.295 ;
        RECT 42.230 191.105 44.150 191.275 ;
        RECT 42.230 190.210 42.420 191.105 ;
        RECT 44.320 190.935 44.490 191.445 ;
        RECT 44.660 191.185 45.180 191.495 ;
        RECT 42.590 190.765 44.490 190.935 ;
        RECT 42.590 190.705 42.920 190.765 ;
        RECT 43.070 190.535 43.400 190.595 ;
        RECT 42.740 190.265 43.400 190.535 ;
        RECT 42.230 189.880 42.550 190.210 ;
        RECT 42.730 189.615 43.390 190.095 ;
        RECT 43.590 190.005 43.760 190.765 ;
        RECT 44.660 190.595 44.840 191.005 ;
        RECT 43.930 190.425 44.260 190.545 ;
        RECT 45.010 190.425 45.180 191.185 ;
        RECT 43.930 190.255 45.180 190.425 ;
        RECT 45.350 191.365 46.720 191.615 ;
        RECT 45.350 190.595 45.540 191.365 ;
        RECT 46.470 191.105 46.720 191.365 ;
        RECT 45.710 190.935 45.960 191.095 ;
        RECT 46.890 190.935 47.060 191.780 ;
        RECT 47.955 191.495 48.125 191.995 ;
        RECT 48.295 191.665 48.625 192.165 ;
        RECT 47.230 191.105 47.730 191.485 ;
        RECT 47.955 191.325 48.650 191.495 ;
        RECT 45.710 190.765 47.060 190.935 ;
        RECT 46.640 190.725 47.060 190.765 ;
        RECT 45.350 190.255 45.770 190.595 ;
        RECT 46.060 190.265 46.470 190.595 ;
        RECT 43.590 189.835 44.440 190.005 ;
        RECT 45.000 189.615 45.320 190.075 ;
        RECT 45.520 189.825 45.770 190.255 ;
        RECT 46.060 189.615 46.470 190.055 ;
        RECT 46.640 189.995 46.810 190.725 ;
        RECT 46.980 190.175 47.330 190.545 ;
        RECT 47.510 190.235 47.730 191.105 ;
        RECT 47.900 190.535 48.310 191.155 ;
        RECT 48.480 190.355 48.650 191.325 ;
        RECT 47.955 190.165 48.650 190.355 ;
        RECT 46.640 189.795 47.655 189.995 ;
        RECT 47.955 189.835 48.125 190.165 ;
        RECT 48.295 189.615 48.625 189.995 ;
        RECT 48.840 189.875 49.065 191.995 ;
        RECT 49.235 191.665 49.565 192.165 ;
        RECT 49.735 191.495 49.905 191.995 ;
        RECT 49.240 191.325 49.905 191.495 ;
        RECT 49.240 190.335 49.470 191.325 ;
        RECT 49.640 190.505 49.990 191.155 ;
        RECT 50.165 191.000 50.455 192.165 ;
        RECT 50.630 191.025 50.965 191.995 ;
        RECT 51.135 191.025 51.305 192.165 ;
        RECT 51.475 191.825 53.505 191.995 ;
        RECT 50.630 190.355 50.800 191.025 ;
        RECT 51.475 190.855 51.645 191.825 ;
        RECT 50.970 190.525 51.225 190.855 ;
        RECT 51.450 190.525 51.645 190.855 ;
        RECT 51.815 191.485 52.940 191.655 ;
        RECT 51.055 190.355 51.225 190.525 ;
        RECT 51.815 190.355 51.985 191.485 ;
        RECT 49.240 190.165 49.905 190.335 ;
        RECT 49.235 189.615 49.565 189.995 ;
        RECT 49.735 189.875 49.905 190.165 ;
        RECT 50.165 189.615 50.455 190.340 ;
        RECT 50.630 189.785 50.885 190.355 ;
        RECT 51.055 190.185 51.985 190.355 ;
        RECT 52.155 191.145 53.165 191.315 ;
        RECT 52.155 190.345 52.325 191.145 ;
        RECT 51.810 190.150 51.985 190.185 ;
        RECT 51.055 189.615 51.385 190.015 ;
        RECT 51.810 189.785 52.340 190.150 ;
        RECT 52.530 190.125 52.805 190.945 ;
        RECT 52.525 189.955 52.805 190.125 ;
        RECT 52.530 189.785 52.805 189.955 ;
        RECT 52.975 189.785 53.165 191.145 ;
        RECT 53.335 191.160 53.505 191.825 ;
        RECT 53.675 191.405 53.845 192.165 ;
        RECT 54.080 191.405 54.595 191.815 ;
        RECT 53.335 190.970 54.085 191.160 ;
        RECT 54.255 190.595 54.595 191.405 ;
        RECT 55.265 191.025 55.495 192.165 ;
        RECT 55.665 191.015 55.995 191.995 ;
        RECT 56.165 191.025 56.375 192.165 ;
        RECT 56.610 191.025 56.945 191.995 ;
        RECT 57.115 191.025 57.285 192.165 ;
        RECT 57.455 191.825 59.485 191.995 ;
        RECT 55.245 190.605 55.575 190.855 ;
        RECT 53.365 190.425 54.595 190.595 ;
        RECT 53.345 189.615 53.855 190.150 ;
        RECT 54.075 189.820 54.320 190.425 ;
        RECT 55.265 189.615 55.495 190.435 ;
        RECT 55.745 190.415 55.995 191.015 ;
        RECT 55.665 189.785 55.995 190.415 ;
        RECT 56.165 189.615 56.375 190.435 ;
        RECT 56.610 190.355 56.780 191.025 ;
        RECT 57.455 190.855 57.625 191.825 ;
        RECT 56.950 190.525 57.205 190.855 ;
        RECT 57.430 190.525 57.625 190.855 ;
        RECT 57.795 191.485 58.920 191.655 ;
        RECT 57.035 190.355 57.205 190.525 ;
        RECT 57.795 190.355 57.965 191.485 ;
        RECT 56.610 189.785 56.865 190.355 ;
        RECT 57.035 190.185 57.965 190.355 ;
        RECT 58.135 191.145 59.145 191.315 ;
        RECT 58.135 190.345 58.305 191.145 ;
        RECT 58.510 190.805 58.785 190.945 ;
        RECT 58.505 190.635 58.785 190.805 ;
        RECT 57.790 190.150 57.965 190.185 ;
        RECT 57.035 189.615 57.365 190.015 ;
        RECT 57.790 189.785 58.320 190.150 ;
        RECT 58.510 189.785 58.785 190.635 ;
        RECT 58.955 189.785 59.145 191.145 ;
        RECT 59.315 191.160 59.485 191.825 ;
        RECT 59.655 191.405 59.825 192.165 ;
        RECT 60.060 191.405 60.575 191.815 ;
        RECT 59.315 190.970 60.065 191.160 ;
        RECT 60.235 190.595 60.575 191.405 ;
        RECT 59.345 190.425 60.575 190.595 ;
        RECT 60.745 191.405 61.260 191.815 ;
        RECT 61.495 191.405 61.665 192.165 ;
        RECT 61.835 191.825 63.865 191.995 ;
        RECT 60.745 190.595 61.085 191.405 ;
        RECT 61.835 191.160 62.005 191.825 ;
        RECT 62.400 191.485 63.525 191.655 ;
        RECT 61.255 190.970 62.005 191.160 ;
        RECT 62.175 191.145 63.185 191.315 ;
        RECT 60.745 190.425 61.975 190.595 ;
        RECT 59.325 189.615 59.835 190.150 ;
        RECT 60.055 189.820 60.300 190.425 ;
        RECT 61.020 189.820 61.265 190.425 ;
        RECT 61.485 189.615 61.995 190.150 ;
        RECT 62.175 189.785 62.365 191.145 ;
        RECT 62.535 190.125 62.810 190.945 ;
        RECT 63.015 190.345 63.185 191.145 ;
        RECT 63.355 190.355 63.525 191.485 ;
        RECT 63.695 190.855 63.865 191.825 ;
        RECT 64.035 191.025 64.205 192.165 ;
        RECT 64.375 191.025 64.710 191.995 ;
        RECT 63.695 190.525 63.890 190.855 ;
        RECT 64.115 190.525 64.370 190.855 ;
        RECT 64.115 190.355 64.285 190.525 ;
        RECT 64.540 190.355 64.710 191.025 ;
        RECT 63.355 190.185 64.285 190.355 ;
        RECT 63.355 190.150 63.530 190.185 ;
        RECT 62.535 189.955 62.815 190.125 ;
        RECT 62.535 189.785 62.810 189.955 ;
        RECT 63.000 189.785 63.530 190.150 ;
        RECT 63.955 189.615 64.285 190.015 ;
        RECT 64.455 189.785 64.710 190.355 ;
        RECT 64.890 190.975 65.145 191.855 ;
        RECT 65.315 191.025 65.620 192.165 ;
        RECT 65.960 191.785 66.290 192.165 ;
        RECT 66.470 191.615 66.640 191.905 ;
        RECT 66.810 191.705 67.060 192.165 ;
        RECT 65.840 191.445 66.640 191.615 ;
        RECT 67.230 191.655 68.100 191.995 ;
        RECT 64.890 190.325 65.100 190.975 ;
        RECT 65.840 190.855 66.010 191.445 ;
        RECT 67.230 191.275 67.400 191.655 ;
        RECT 68.335 191.535 68.505 191.995 ;
        RECT 68.675 191.705 69.045 192.165 ;
        RECT 69.340 191.565 69.510 191.905 ;
        RECT 69.680 191.735 70.010 192.165 ;
        RECT 70.245 191.565 70.415 191.905 ;
        RECT 66.180 191.105 67.400 191.275 ;
        RECT 67.570 191.195 68.030 191.485 ;
        RECT 68.335 191.365 68.895 191.535 ;
        RECT 69.340 191.395 70.415 191.565 ;
        RECT 70.585 191.665 71.265 191.995 ;
        RECT 71.480 191.665 71.730 191.995 ;
        RECT 71.900 191.705 72.150 192.165 ;
        RECT 68.725 191.225 68.895 191.365 ;
        RECT 67.570 191.185 68.535 191.195 ;
        RECT 67.230 191.015 67.400 191.105 ;
        RECT 67.860 191.025 68.535 191.185 ;
        RECT 65.270 190.825 66.010 190.855 ;
        RECT 65.270 190.525 66.185 190.825 ;
        RECT 65.860 190.350 66.185 190.525 ;
        RECT 64.890 189.795 65.145 190.325 ;
        RECT 65.315 189.615 65.620 190.075 ;
        RECT 65.865 189.995 66.185 190.350 ;
        RECT 66.355 190.565 66.895 190.935 ;
        RECT 67.230 190.845 67.635 191.015 ;
        RECT 66.355 190.165 66.595 190.565 ;
        RECT 67.075 190.395 67.295 190.675 ;
        RECT 66.765 190.225 67.295 190.395 ;
        RECT 66.765 189.995 66.935 190.225 ;
        RECT 67.465 190.065 67.635 190.845 ;
        RECT 67.805 190.235 68.155 190.855 ;
        RECT 68.325 190.235 68.535 191.025 ;
        RECT 68.725 191.055 70.225 191.225 ;
        RECT 68.725 190.365 68.895 191.055 ;
        RECT 70.585 190.885 70.755 191.665 ;
        RECT 71.560 191.535 71.730 191.665 ;
        RECT 69.065 190.715 70.755 190.885 ;
        RECT 70.925 191.105 71.390 191.495 ;
        RECT 71.560 191.365 71.955 191.535 ;
        RECT 69.065 190.535 69.235 190.715 ;
        RECT 65.865 189.825 66.935 189.995 ;
        RECT 67.105 189.615 67.295 190.055 ;
        RECT 67.465 189.785 68.415 190.065 ;
        RECT 68.725 189.975 68.985 190.365 ;
        RECT 69.405 190.295 70.195 190.545 ;
        RECT 68.635 189.805 68.985 189.975 ;
        RECT 69.195 189.615 69.525 190.075 ;
        RECT 70.400 190.005 70.570 190.715 ;
        RECT 70.925 190.515 71.095 191.105 ;
        RECT 70.740 190.295 71.095 190.515 ;
        RECT 71.265 190.295 71.615 190.915 ;
        RECT 71.785 190.005 71.955 191.365 ;
        RECT 72.320 191.195 72.645 191.980 ;
        RECT 72.125 190.145 72.585 191.195 ;
        RECT 70.400 189.835 71.255 190.005 ;
        RECT 71.460 189.835 71.955 190.005 ;
        RECT 72.125 189.615 72.455 189.975 ;
        RECT 72.815 189.875 72.985 191.995 ;
        RECT 73.155 191.665 73.485 192.165 ;
        RECT 73.655 191.495 73.910 191.995 ;
        RECT 73.160 191.325 73.910 191.495 ;
        RECT 73.160 190.335 73.390 191.325 ;
        RECT 74.175 191.235 74.345 191.995 ;
        RECT 74.560 191.405 74.890 192.165 ;
        RECT 73.560 190.505 73.910 191.155 ;
        RECT 74.175 191.065 74.890 191.235 ;
        RECT 75.060 191.090 75.315 191.995 ;
        RECT 74.085 190.515 74.440 190.885 ;
        RECT 74.720 190.855 74.890 191.065 ;
        RECT 74.720 190.525 74.975 190.855 ;
        RECT 74.720 190.335 74.890 190.525 ;
        RECT 75.145 190.360 75.315 191.090 ;
        RECT 75.490 191.015 75.750 192.165 ;
        RECT 75.925 191.000 76.215 192.165 ;
        RECT 77.305 191.665 77.565 191.995 ;
        RECT 77.875 191.785 78.205 192.165 ;
        RECT 77.305 190.985 77.475 191.665 ;
        RECT 78.445 191.615 78.635 191.995 ;
        RECT 78.885 191.785 79.215 192.165 ;
        RECT 79.425 191.615 79.595 191.995 ;
        RECT 79.790 191.785 80.120 192.165 ;
        RECT 80.380 191.615 80.550 191.995 ;
        RECT 80.975 191.785 81.305 192.165 ;
        RECT 77.645 191.155 77.995 191.485 ;
        RECT 78.445 191.445 79.185 191.615 ;
        RECT 78.265 191.105 78.845 191.275 ;
        RECT 78.265 190.985 78.435 191.105 ;
        RECT 77.305 190.815 78.435 190.985 ;
        RECT 79.015 190.935 79.185 191.445 ;
        RECT 73.160 190.165 73.910 190.335 ;
        RECT 73.155 189.615 73.485 189.995 ;
        RECT 73.655 189.875 73.910 190.165 ;
        RECT 74.175 190.165 74.890 190.335 ;
        RECT 74.175 189.785 74.345 190.165 ;
        RECT 74.560 189.615 74.890 189.995 ;
        RECT 75.060 189.785 75.315 190.360 ;
        RECT 75.490 189.615 75.750 190.455 ;
        RECT 75.925 189.615 76.215 190.340 ;
        RECT 77.305 190.115 77.475 190.815 ;
        RECT 78.615 190.765 79.185 190.935 ;
        RECT 79.355 191.445 81.305 191.615 ;
        RECT 77.825 190.475 78.445 190.645 ;
        RECT 77.825 190.295 78.035 190.475 ;
        RECT 78.615 190.285 78.785 190.765 ;
        RECT 79.355 190.455 79.525 191.445 ;
        RECT 80.115 190.855 80.300 191.165 ;
        RECT 80.570 190.855 80.765 191.165 ;
        RECT 77.305 189.785 77.565 190.115 ;
        RECT 77.875 189.615 78.205 189.995 ;
        RECT 78.385 189.955 78.785 190.285 ;
        RECT 78.975 190.125 79.525 190.455 ;
        RECT 79.695 189.955 79.865 190.855 ;
        RECT 78.385 189.785 79.865 189.955 ;
        RECT 80.115 190.525 80.345 190.855 ;
        RECT 80.570 190.525 80.825 190.855 ;
        RECT 81.135 190.525 81.305 191.445 ;
        RECT 80.115 189.945 80.300 190.525 ;
        RECT 80.570 189.950 80.765 190.525 ;
        RECT 80.975 189.615 81.305 189.995 ;
        RECT 81.475 189.785 81.735 191.995 ;
        RECT 81.905 191.075 83.115 192.165 ;
        RECT 83.285 191.405 83.800 191.815 ;
        RECT 84.035 191.405 84.205 192.165 ;
        RECT 84.375 191.825 86.405 191.995 ;
        RECT 81.905 190.535 82.425 191.075 ;
        RECT 82.595 190.365 83.115 190.905 ;
        RECT 83.285 190.595 83.625 191.405 ;
        RECT 84.375 191.160 84.545 191.825 ;
        RECT 84.940 191.485 86.065 191.655 ;
        RECT 83.795 190.970 84.545 191.160 ;
        RECT 84.715 191.145 85.725 191.315 ;
        RECT 83.285 190.425 84.515 190.595 ;
        RECT 81.905 189.615 83.115 190.365 ;
        RECT 83.560 189.820 83.805 190.425 ;
        RECT 84.025 189.615 84.535 190.150 ;
        RECT 84.715 189.785 84.905 191.145 ;
        RECT 85.075 190.125 85.350 190.945 ;
        RECT 85.555 190.345 85.725 191.145 ;
        RECT 85.895 190.355 86.065 191.485 ;
        RECT 86.235 190.855 86.405 191.825 ;
        RECT 86.575 191.025 86.745 192.165 ;
        RECT 86.915 191.025 87.250 191.995 ;
        RECT 86.235 190.525 86.430 190.855 ;
        RECT 86.655 190.525 86.910 190.855 ;
        RECT 86.655 190.355 86.825 190.525 ;
        RECT 87.080 190.355 87.250 191.025 ;
        RECT 85.895 190.185 86.825 190.355 ;
        RECT 85.895 190.150 86.070 190.185 ;
        RECT 85.075 189.955 85.355 190.125 ;
        RECT 85.075 189.785 85.350 189.955 ;
        RECT 85.540 189.785 86.070 190.150 ;
        RECT 86.495 189.615 86.825 190.015 ;
        RECT 86.995 189.785 87.250 190.355 ;
        RECT 87.800 191.185 88.055 191.855 ;
        RECT 88.235 191.365 88.520 192.165 ;
        RECT 88.700 191.445 89.030 191.955 ;
        RECT 87.800 190.325 87.980 191.185 ;
        RECT 88.700 190.855 88.950 191.445 ;
        RECT 89.300 191.295 89.470 191.905 ;
        RECT 89.640 191.475 89.970 192.165 ;
        RECT 90.200 191.615 90.440 191.905 ;
        RECT 90.640 191.785 91.060 192.165 ;
        RECT 91.240 191.695 91.870 191.945 ;
        RECT 92.340 191.785 92.670 192.165 ;
        RECT 91.240 191.615 91.410 191.695 ;
        RECT 92.840 191.615 93.010 191.905 ;
        RECT 93.190 191.785 93.570 192.165 ;
        RECT 93.810 191.780 94.640 191.950 ;
        RECT 90.200 191.445 91.410 191.615 ;
        RECT 88.150 190.525 88.950 190.855 ;
        RECT 87.800 190.125 88.055 190.325 ;
        RECT 87.715 189.955 88.055 190.125 ;
        RECT 87.800 189.795 88.055 189.955 ;
        RECT 88.235 189.615 88.520 190.075 ;
        RECT 88.700 189.875 88.950 190.525 ;
        RECT 89.150 191.275 89.470 191.295 ;
        RECT 89.150 191.105 91.070 191.275 ;
        RECT 89.150 190.210 89.340 191.105 ;
        RECT 91.240 190.935 91.410 191.445 ;
        RECT 91.580 191.185 92.100 191.495 ;
        RECT 89.510 190.765 91.410 190.935 ;
        RECT 89.510 190.705 89.840 190.765 ;
        RECT 89.990 190.535 90.320 190.595 ;
        RECT 89.660 190.265 90.320 190.535 ;
        RECT 89.150 189.880 89.470 190.210 ;
        RECT 89.650 189.615 90.310 190.095 ;
        RECT 90.510 190.005 90.680 190.765 ;
        RECT 91.580 190.595 91.760 191.005 ;
        RECT 90.850 190.425 91.180 190.545 ;
        RECT 91.930 190.425 92.100 191.185 ;
        RECT 90.850 190.255 92.100 190.425 ;
        RECT 92.270 191.365 93.640 191.615 ;
        RECT 92.270 190.595 92.460 191.365 ;
        RECT 93.390 191.105 93.640 191.365 ;
        RECT 92.630 190.935 92.880 191.095 ;
        RECT 93.810 190.935 93.980 191.780 ;
        RECT 94.875 191.495 95.045 191.995 ;
        RECT 95.215 191.665 95.545 192.165 ;
        RECT 94.150 191.105 94.650 191.485 ;
        RECT 94.875 191.325 95.570 191.495 ;
        RECT 92.630 190.765 93.980 190.935 ;
        RECT 93.560 190.725 93.980 190.765 ;
        RECT 92.270 190.255 92.690 190.595 ;
        RECT 92.980 190.265 93.390 190.595 ;
        RECT 90.510 189.835 91.360 190.005 ;
        RECT 91.920 189.615 92.240 190.075 ;
        RECT 92.440 189.825 92.690 190.255 ;
        RECT 92.980 189.615 93.390 190.055 ;
        RECT 93.560 189.995 93.730 190.725 ;
        RECT 93.900 190.175 94.250 190.545 ;
        RECT 94.430 190.235 94.650 191.105 ;
        RECT 94.820 190.535 95.230 191.155 ;
        RECT 95.400 190.355 95.570 191.325 ;
        RECT 94.875 190.165 95.570 190.355 ;
        RECT 93.560 189.795 94.575 189.995 ;
        RECT 94.875 189.835 95.045 190.165 ;
        RECT 95.215 189.615 95.545 189.995 ;
        RECT 95.760 189.875 95.985 191.995 ;
        RECT 96.155 191.665 96.485 192.165 ;
        RECT 96.655 191.495 96.825 191.995 ;
        RECT 96.160 191.325 96.825 191.495 ;
        RECT 96.160 190.335 96.390 191.325 ;
        RECT 96.560 190.505 96.910 191.155 ;
        RECT 97.085 191.090 97.355 191.995 ;
        RECT 97.525 191.405 97.855 192.165 ;
        RECT 98.035 191.235 98.205 191.995 ;
        RECT 96.160 190.165 96.825 190.335 ;
        RECT 96.155 189.615 96.485 189.995 ;
        RECT 96.655 189.875 96.825 190.165 ;
        RECT 97.085 190.290 97.255 191.090 ;
        RECT 97.540 191.065 98.205 191.235 ;
        RECT 97.540 190.920 97.710 191.065 ;
        RECT 98.505 191.025 98.735 192.165 ;
        RECT 98.905 191.015 99.235 191.995 ;
        RECT 99.405 191.025 99.615 192.165 ;
        RECT 99.845 191.075 101.515 192.165 ;
        RECT 97.425 190.590 97.710 190.920 ;
        RECT 97.540 190.335 97.710 190.590 ;
        RECT 97.945 190.515 98.275 190.885 ;
        RECT 98.485 190.605 98.815 190.855 ;
        RECT 97.085 189.785 97.345 190.290 ;
        RECT 97.540 190.165 98.205 190.335 ;
        RECT 97.525 189.615 97.855 189.995 ;
        RECT 98.035 189.785 98.205 190.165 ;
        RECT 98.505 189.615 98.735 190.435 ;
        RECT 98.985 190.415 99.235 191.015 ;
        RECT 99.845 190.555 100.595 191.075 ;
        RECT 101.685 191.000 101.975 192.165 ;
        RECT 102.610 190.975 102.865 191.855 ;
        RECT 103.035 191.025 103.340 192.165 ;
        RECT 103.680 191.785 104.010 192.165 ;
        RECT 104.190 191.615 104.360 191.905 ;
        RECT 104.530 191.705 104.780 192.165 ;
        RECT 103.560 191.445 104.360 191.615 ;
        RECT 104.950 191.655 105.820 191.995 ;
        RECT 98.905 189.785 99.235 190.415 ;
        RECT 99.405 189.615 99.615 190.435 ;
        RECT 100.765 190.385 101.515 190.905 ;
        RECT 99.845 189.615 101.515 190.385 ;
        RECT 101.685 189.615 101.975 190.340 ;
        RECT 102.610 190.325 102.820 190.975 ;
        RECT 103.560 190.855 103.730 191.445 ;
        RECT 104.950 191.275 105.120 191.655 ;
        RECT 106.055 191.535 106.225 191.995 ;
        RECT 106.395 191.705 106.765 192.165 ;
        RECT 107.060 191.565 107.230 191.905 ;
        RECT 107.400 191.735 107.730 192.165 ;
        RECT 107.965 191.565 108.135 191.905 ;
        RECT 103.900 191.105 105.120 191.275 ;
        RECT 105.290 191.195 105.750 191.485 ;
        RECT 106.055 191.365 106.615 191.535 ;
        RECT 107.060 191.395 108.135 191.565 ;
        RECT 108.305 191.665 108.985 191.995 ;
        RECT 109.200 191.665 109.450 191.995 ;
        RECT 109.620 191.705 109.870 192.165 ;
        RECT 106.445 191.225 106.615 191.365 ;
        RECT 105.290 191.185 106.255 191.195 ;
        RECT 104.950 191.015 105.120 191.105 ;
        RECT 105.580 191.025 106.255 191.185 ;
        RECT 102.990 190.825 103.730 190.855 ;
        RECT 102.990 190.525 103.905 190.825 ;
        RECT 103.580 190.350 103.905 190.525 ;
        RECT 102.610 189.795 102.865 190.325 ;
        RECT 103.035 189.615 103.340 190.075 ;
        RECT 103.585 189.995 103.905 190.350 ;
        RECT 104.075 190.565 104.615 190.935 ;
        RECT 104.950 190.845 105.355 191.015 ;
        RECT 104.075 190.165 104.315 190.565 ;
        RECT 104.795 190.395 105.015 190.675 ;
        RECT 104.485 190.225 105.015 190.395 ;
        RECT 104.485 189.995 104.655 190.225 ;
        RECT 105.185 190.065 105.355 190.845 ;
        RECT 105.525 190.235 105.875 190.855 ;
        RECT 106.045 190.235 106.255 191.025 ;
        RECT 106.445 191.055 107.945 191.225 ;
        RECT 106.445 190.365 106.615 191.055 ;
        RECT 108.305 190.885 108.475 191.665 ;
        RECT 109.280 191.535 109.450 191.665 ;
        RECT 106.785 190.715 108.475 190.885 ;
        RECT 108.645 191.105 109.110 191.495 ;
        RECT 109.280 191.365 109.675 191.535 ;
        RECT 106.785 190.535 106.955 190.715 ;
        RECT 103.585 189.825 104.655 189.995 ;
        RECT 104.825 189.615 105.015 190.055 ;
        RECT 105.185 189.785 106.135 190.065 ;
        RECT 106.445 189.975 106.705 190.365 ;
        RECT 107.125 190.295 107.915 190.545 ;
        RECT 106.355 189.805 106.705 189.975 ;
        RECT 106.915 189.615 107.245 190.075 ;
        RECT 108.120 190.005 108.290 190.715 ;
        RECT 108.645 190.515 108.815 191.105 ;
        RECT 108.460 190.295 108.815 190.515 ;
        RECT 108.985 190.295 109.335 190.915 ;
        RECT 109.505 190.005 109.675 191.365 ;
        RECT 110.040 191.195 110.365 191.980 ;
        RECT 109.845 190.145 110.305 191.195 ;
        RECT 108.120 189.835 108.975 190.005 ;
        RECT 109.180 189.835 109.675 190.005 ;
        RECT 109.845 189.615 110.175 189.975 ;
        RECT 110.535 189.875 110.705 191.995 ;
        RECT 110.875 191.665 111.205 192.165 ;
        RECT 111.375 191.495 111.630 191.995 ;
        RECT 110.880 191.325 111.630 191.495 ;
        RECT 112.725 191.405 113.240 191.815 ;
        RECT 113.475 191.405 113.645 192.165 ;
        RECT 113.815 191.825 115.845 191.995 ;
        RECT 110.880 190.335 111.110 191.325 ;
        RECT 111.280 190.505 111.630 191.155 ;
        RECT 112.725 190.595 113.065 191.405 ;
        RECT 113.815 191.160 113.985 191.825 ;
        RECT 114.380 191.485 115.505 191.655 ;
        RECT 113.235 190.970 113.985 191.160 ;
        RECT 114.155 191.145 115.165 191.315 ;
        RECT 112.725 190.425 113.955 190.595 ;
        RECT 110.880 190.165 111.630 190.335 ;
        RECT 110.875 189.615 111.205 189.995 ;
        RECT 111.375 189.875 111.630 190.165 ;
        RECT 113.000 189.820 113.245 190.425 ;
        RECT 113.465 189.615 113.975 190.150 ;
        RECT 114.155 189.785 114.345 191.145 ;
        RECT 114.515 190.805 114.790 190.945 ;
        RECT 114.515 190.635 114.795 190.805 ;
        RECT 114.515 189.785 114.790 190.635 ;
        RECT 114.995 190.345 115.165 191.145 ;
        RECT 115.335 190.355 115.505 191.485 ;
        RECT 115.675 190.855 115.845 191.825 ;
        RECT 116.015 191.025 116.185 192.165 ;
        RECT 116.355 191.025 116.690 191.995 ;
        RECT 115.675 190.525 115.870 190.855 ;
        RECT 116.095 190.525 116.350 190.855 ;
        RECT 116.095 190.355 116.265 190.525 ;
        RECT 116.520 190.355 116.690 191.025 ;
        RECT 115.335 190.185 116.265 190.355 ;
        RECT 115.335 190.150 115.510 190.185 ;
        RECT 114.980 189.785 115.510 190.150 ;
        RECT 115.935 189.615 116.265 190.015 ;
        RECT 116.435 189.785 116.690 190.355 ;
        RECT 116.870 190.975 117.125 191.855 ;
        RECT 117.295 191.025 117.600 192.165 ;
        RECT 117.940 191.785 118.270 192.165 ;
        RECT 118.450 191.615 118.620 191.905 ;
        RECT 118.790 191.705 119.040 192.165 ;
        RECT 117.820 191.445 118.620 191.615 ;
        RECT 119.210 191.655 120.080 191.995 ;
        RECT 116.870 190.325 117.080 190.975 ;
        RECT 117.820 190.855 117.990 191.445 ;
        RECT 119.210 191.275 119.380 191.655 ;
        RECT 120.315 191.535 120.485 191.995 ;
        RECT 120.655 191.705 121.025 192.165 ;
        RECT 121.320 191.565 121.490 191.905 ;
        RECT 121.660 191.735 121.990 192.165 ;
        RECT 122.225 191.565 122.395 191.905 ;
        RECT 118.160 191.105 119.380 191.275 ;
        RECT 119.550 191.195 120.010 191.485 ;
        RECT 120.315 191.365 120.875 191.535 ;
        RECT 121.320 191.395 122.395 191.565 ;
        RECT 122.565 191.665 123.245 191.995 ;
        RECT 123.460 191.665 123.710 191.995 ;
        RECT 123.880 191.705 124.130 192.165 ;
        RECT 120.705 191.225 120.875 191.365 ;
        RECT 119.550 191.185 120.515 191.195 ;
        RECT 119.210 191.015 119.380 191.105 ;
        RECT 119.840 191.025 120.515 191.185 ;
        RECT 117.250 190.825 117.990 190.855 ;
        RECT 117.250 190.525 118.165 190.825 ;
        RECT 117.840 190.350 118.165 190.525 ;
        RECT 116.870 189.795 117.125 190.325 ;
        RECT 117.295 189.615 117.600 190.075 ;
        RECT 117.845 189.995 118.165 190.350 ;
        RECT 118.335 190.565 118.875 190.935 ;
        RECT 119.210 190.845 119.615 191.015 ;
        RECT 118.335 190.165 118.575 190.565 ;
        RECT 119.055 190.395 119.275 190.675 ;
        RECT 118.745 190.225 119.275 190.395 ;
        RECT 118.745 189.995 118.915 190.225 ;
        RECT 119.445 190.065 119.615 190.845 ;
        RECT 119.785 190.235 120.135 190.855 ;
        RECT 120.305 190.235 120.515 191.025 ;
        RECT 120.705 191.055 122.205 191.225 ;
        RECT 120.705 190.365 120.875 191.055 ;
        RECT 122.565 190.885 122.735 191.665 ;
        RECT 123.540 191.535 123.710 191.665 ;
        RECT 121.045 190.715 122.735 190.885 ;
        RECT 122.905 191.105 123.370 191.495 ;
        RECT 123.540 191.365 123.935 191.535 ;
        RECT 121.045 190.535 121.215 190.715 ;
        RECT 117.845 189.825 118.915 189.995 ;
        RECT 119.085 189.615 119.275 190.055 ;
        RECT 119.445 189.785 120.395 190.065 ;
        RECT 120.705 189.975 120.965 190.365 ;
        RECT 121.385 190.295 122.175 190.545 ;
        RECT 120.615 189.805 120.965 189.975 ;
        RECT 121.175 189.615 121.505 190.075 ;
        RECT 122.380 190.005 122.550 190.715 ;
        RECT 122.905 190.515 123.075 191.105 ;
        RECT 122.720 190.295 123.075 190.515 ;
        RECT 123.245 190.295 123.595 190.915 ;
        RECT 123.765 190.005 123.935 191.365 ;
        RECT 124.300 191.195 124.625 191.980 ;
        RECT 124.105 190.145 124.565 191.195 ;
        RECT 122.380 189.835 123.235 190.005 ;
        RECT 123.440 189.835 123.935 190.005 ;
        RECT 124.105 189.615 124.435 189.975 ;
        RECT 124.795 189.875 124.965 191.995 ;
        RECT 125.135 191.665 125.465 192.165 ;
        RECT 125.635 191.495 125.890 191.995 ;
        RECT 125.140 191.325 125.890 191.495 ;
        RECT 125.140 190.335 125.370 191.325 ;
        RECT 125.540 190.505 125.890 191.155 ;
        RECT 126.525 191.075 127.735 192.165 ;
        RECT 126.525 190.535 127.045 191.075 ;
        RECT 127.215 190.365 127.735 190.905 ;
        RECT 125.140 190.165 125.890 190.335 ;
        RECT 125.135 189.615 125.465 189.995 ;
        RECT 125.635 189.875 125.890 190.165 ;
        RECT 126.525 189.615 127.735 190.365 ;
        RECT 29.840 189.445 127.820 189.615 ;
        RECT 29.925 188.695 31.135 189.445 ;
        RECT 29.925 188.155 30.445 188.695 ;
        RECT 31.765 188.675 34.355 189.445 ;
        RECT 30.615 187.985 31.135 188.525 ;
        RECT 29.925 186.895 31.135 187.985 ;
        RECT 31.765 187.985 32.975 188.505 ;
        RECT 33.145 188.155 34.355 188.675 ;
        RECT 34.565 188.625 34.795 189.445 ;
        RECT 34.965 188.645 35.295 189.275 ;
        RECT 34.545 188.205 34.875 188.455 ;
        RECT 35.045 188.045 35.295 188.645 ;
        RECT 35.465 188.625 35.675 189.445 ;
        RECT 35.945 188.625 36.175 189.445 ;
        RECT 36.345 188.645 36.675 189.275 ;
        RECT 35.925 188.205 36.255 188.455 ;
        RECT 36.425 188.045 36.675 188.645 ;
        RECT 36.845 188.625 37.055 189.445 ;
        RECT 37.285 188.720 37.575 189.445 ;
        RECT 37.750 188.735 38.005 189.265 ;
        RECT 38.175 188.985 38.480 189.445 ;
        RECT 38.725 189.065 39.795 189.235 ;
        RECT 37.750 188.085 37.960 188.735 ;
        RECT 38.725 188.710 39.045 189.065 ;
        RECT 38.720 188.535 39.045 188.710 ;
        RECT 38.130 188.235 39.045 188.535 ;
        RECT 39.215 188.495 39.455 188.895 ;
        RECT 39.625 188.835 39.795 189.065 ;
        RECT 39.965 189.005 40.155 189.445 ;
        RECT 40.325 188.995 41.275 189.275 ;
        RECT 41.495 189.085 41.845 189.255 ;
        RECT 39.625 188.665 40.155 188.835 ;
        RECT 38.130 188.205 38.870 188.235 ;
        RECT 31.765 186.895 34.355 187.985 ;
        RECT 34.565 186.895 34.795 188.035 ;
        RECT 34.965 187.065 35.295 188.045 ;
        RECT 35.465 186.895 35.675 188.035 ;
        RECT 35.945 186.895 36.175 188.035 ;
        RECT 36.345 187.065 36.675 188.045 ;
        RECT 36.845 186.895 37.055 188.035 ;
        RECT 37.285 186.895 37.575 188.060 ;
        RECT 37.750 187.205 38.005 188.085 ;
        RECT 38.175 186.895 38.480 188.035 ;
        RECT 38.700 187.615 38.870 188.205 ;
        RECT 39.215 188.125 39.755 188.495 ;
        RECT 39.935 188.385 40.155 188.665 ;
        RECT 40.325 188.215 40.495 188.995 ;
        RECT 40.090 188.045 40.495 188.215 ;
        RECT 40.665 188.205 41.015 188.825 ;
        RECT 40.090 187.955 40.260 188.045 ;
        RECT 41.185 188.035 41.395 188.825 ;
        RECT 39.040 187.785 40.260 187.955 ;
        RECT 40.720 187.875 41.395 188.035 ;
        RECT 38.700 187.445 39.500 187.615 ;
        RECT 38.820 186.895 39.150 187.275 ;
        RECT 39.330 187.155 39.500 187.445 ;
        RECT 40.090 187.405 40.260 187.785 ;
        RECT 40.430 187.865 41.395 187.875 ;
        RECT 41.585 188.695 41.845 189.085 ;
        RECT 42.055 188.985 42.385 189.445 ;
        RECT 43.260 189.055 44.115 189.225 ;
        RECT 44.320 189.055 44.815 189.225 ;
        RECT 44.985 189.085 45.315 189.445 ;
        RECT 41.585 188.005 41.755 188.695 ;
        RECT 41.925 188.345 42.095 188.525 ;
        RECT 42.265 188.515 43.055 188.765 ;
        RECT 43.260 188.345 43.430 189.055 ;
        RECT 43.600 188.545 43.955 188.765 ;
        RECT 41.925 188.175 43.615 188.345 ;
        RECT 40.430 187.575 40.890 187.865 ;
        RECT 41.585 187.835 43.085 188.005 ;
        RECT 41.585 187.695 41.755 187.835 ;
        RECT 41.195 187.525 41.755 187.695 ;
        RECT 39.670 186.895 39.920 187.355 ;
        RECT 40.090 187.065 40.960 187.405 ;
        RECT 41.195 187.065 41.365 187.525 ;
        RECT 42.200 187.495 43.275 187.665 ;
        RECT 41.535 186.895 41.905 187.355 ;
        RECT 42.200 187.155 42.370 187.495 ;
        RECT 42.540 186.895 42.870 187.325 ;
        RECT 43.105 187.155 43.275 187.495 ;
        RECT 43.445 187.395 43.615 188.175 ;
        RECT 43.785 187.955 43.955 188.545 ;
        RECT 44.125 188.145 44.475 188.765 ;
        RECT 43.785 187.565 44.250 187.955 ;
        RECT 44.645 187.695 44.815 189.055 ;
        RECT 44.985 187.865 45.445 188.915 ;
        RECT 44.420 187.525 44.815 187.695 ;
        RECT 44.420 187.395 44.590 187.525 ;
        RECT 43.445 187.065 44.125 187.395 ;
        RECT 44.340 187.065 44.590 187.395 ;
        RECT 44.760 186.895 45.010 187.355 ;
        RECT 45.180 187.080 45.505 187.865 ;
        RECT 45.675 187.065 45.845 189.185 ;
        RECT 46.015 189.065 46.345 189.445 ;
        RECT 46.515 188.895 46.770 189.185 ;
        RECT 46.020 188.725 46.770 188.895 ;
        RECT 46.020 187.735 46.250 188.725 ;
        RECT 47.220 188.635 47.465 189.240 ;
        RECT 47.685 188.910 48.195 189.445 ;
        RECT 46.420 187.905 46.770 188.555 ;
        RECT 46.945 188.465 48.175 188.635 ;
        RECT 46.020 187.565 46.770 187.735 ;
        RECT 46.015 186.895 46.345 187.395 ;
        RECT 46.515 187.065 46.770 187.565 ;
        RECT 46.945 187.655 47.285 188.465 ;
        RECT 47.455 187.900 48.205 188.090 ;
        RECT 46.945 187.245 47.460 187.655 ;
        RECT 47.695 186.895 47.865 187.655 ;
        RECT 48.035 187.235 48.205 187.900 ;
        RECT 48.375 187.915 48.565 189.275 ;
        RECT 48.735 188.765 49.010 189.275 ;
        RECT 49.200 188.910 49.730 189.275 ;
        RECT 50.155 189.045 50.485 189.445 ;
        RECT 49.555 188.875 49.730 188.910 ;
        RECT 48.735 188.595 49.015 188.765 ;
        RECT 48.735 188.115 49.010 188.595 ;
        RECT 49.215 187.915 49.385 188.715 ;
        RECT 48.375 187.745 49.385 187.915 ;
        RECT 49.555 188.705 50.485 188.875 ;
        RECT 50.655 188.705 50.910 189.275 ;
        RECT 51.175 188.895 51.345 189.275 ;
        RECT 51.525 189.065 51.855 189.445 ;
        RECT 51.175 188.725 51.840 188.895 ;
        RECT 52.035 188.770 52.295 189.275 ;
        RECT 49.555 187.575 49.725 188.705 ;
        RECT 50.315 188.535 50.485 188.705 ;
        RECT 48.600 187.405 49.725 187.575 ;
        RECT 49.895 188.205 50.090 188.535 ;
        RECT 50.315 188.205 50.570 188.535 ;
        RECT 49.895 187.235 50.065 188.205 ;
        RECT 50.740 188.035 50.910 188.705 ;
        RECT 51.105 188.175 51.435 188.545 ;
        RECT 51.670 188.470 51.840 188.725 ;
        RECT 48.035 187.065 50.065 187.235 ;
        RECT 50.235 186.895 50.405 188.035 ;
        RECT 50.575 187.065 50.910 188.035 ;
        RECT 51.670 188.140 51.955 188.470 ;
        RECT 51.670 187.995 51.840 188.140 ;
        RECT 51.175 187.825 51.840 187.995 ;
        RECT 52.125 187.970 52.295 188.770 ;
        RECT 51.175 187.065 51.345 187.825 ;
        RECT 51.525 186.895 51.855 187.655 ;
        RECT 52.025 187.065 52.295 187.970 ;
        RECT 52.470 188.735 52.725 189.265 ;
        RECT 52.895 188.985 53.200 189.445 ;
        RECT 53.445 189.065 54.515 189.235 ;
        RECT 52.470 188.085 52.680 188.735 ;
        RECT 53.445 188.710 53.765 189.065 ;
        RECT 53.440 188.535 53.765 188.710 ;
        RECT 52.850 188.235 53.765 188.535 ;
        RECT 53.935 188.495 54.175 188.895 ;
        RECT 54.345 188.835 54.515 189.065 ;
        RECT 54.685 189.005 54.875 189.445 ;
        RECT 55.045 188.995 55.995 189.275 ;
        RECT 56.215 189.085 56.565 189.255 ;
        RECT 54.345 188.665 54.875 188.835 ;
        RECT 52.850 188.205 53.590 188.235 ;
        RECT 52.470 187.205 52.725 188.085 ;
        RECT 52.895 186.895 53.200 188.035 ;
        RECT 53.420 187.615 53.590 188.205 ;
        RECT 53.935 188.125 54.475 188.495 ;
        RECT 54.655 188.385 54.875 188.665 ;
        RECT 55.045 188.215 55.215 188.995 ;
        RECT 54.810 188.045 55.215 188.215 ;
        RECT 55.385 188.205 55.735 188.825 ;
        RECT 54.810 187.955 54.980 188.045 ;
        RECT 55.905 188.035 56.115 188.825 ;
        RECT 53.760 187.785 54.980 187.955 ;
        RECT 55.440 187.875 56.115 188.035 ;
        RECT 53.420 187.445 54.220 187.615 ;
        RECT 53.540 186.895 53.870 187.275 ;
        RECT 54.050 187.155 54.220 187.445 ;
        RECT 54.810 187.405 54.980 187.785 ;
        RECT 55.150 187.865 56.115 187.875 ;
        RECT 56.305 188.695 56.565 189.085 ;
        RECT 56.775 188.985 57.105 189.445 ;
        RECT 57.980 189.055 58.835 189.225 ;
        RECT 59.040 189.055 59.535 189.225 ;
        RECT 59.705 189.085 60.035 189.445 ;
        RECT 56.305 188.005 56.475 188.695 ;
        RECT 56.645 188.345 56.815 188.525 ;
        RECT 56.985 188.515 57.775 188.765 ;
        RECT 57.980 188.345 58.150 189.055 ;
        RECT 58.320 188.545 58.675 188.765 ;
        RECT 56.645 188.175 58.335 188.345 ;
        RECT 55.150 187.575 55.610 187.865 ;
        RECT 56.305 187.835 57.805 188.005 ;
        RECT 56.305 187.695 56.475 187.835 ;
        RECT 55.915 187.525 56.475 187.695 ;
        RECT 54.390 186.895 54.640 187.355 ;
        RECT 54.810 187.065 55.680 187.405 ;
        RECT 55.915 187.065 56.085 187.525 ;
        RECT 56.920 187.495 57.995 187.665 ;
        RECT 56.255 186.895 56.625 187.355 ;
        RECT 56.920 187.155 57.090 187.495 ;
        RECT 57.260 186.895 57.590 187.325 ;
        RECT 57.825 187.155 57.995 187.495 ;
        RECT 58.165 187.395 58.335 188.175 ;
        RECT 58.505 187.955 58.675 188.545 ;
        RECT 58.845 188.145 59.195 188.765 ;
        RECT 58.505 187.565 58.970 187.955 ;
        RECT 59.365 187.695 59.535 189.055 ;
        RECT 59.705 187.865 60.165 188.915 ;
        RECT 59.140 187.525 59.535 187.695 ;
        RECT 59.140 187.395 59.310 187.525 ;
        RECT 58.165 187.065 58.845 187.395 ;
        RECT 59.060 187.065 59.310 187.395 ;
        RECT 59.480 186.895 59.730 187.355 ;
        RECT 59.900 187.080 60.225 187.865 ;
        RECT 60.395 187.065 60.565 189.185 ;
        RECT 60.735 189.065 61.065 189.445 ;
        RECT 61.235 188.895 61.490 189.185 ;
        RECT 60.740 188.725 61.490 188.895 ;
        RECT 60.740 187.735 60.970 188.725 ;
        RECT 61.725 188.625 61.935 189.445 ;
        RECT 62.105 188.645 62.435 189.275 ;
        RECT 61.140 187.905 61.490 188.555 ;
        RECT 62.105 188.045 62.355 188.645 ;
        RECT 62.605 188.625 62.835 189.445 ;
        RECT 63.045 188.720 63.335 189.445 ;
        RECT 64.055 188.895 64.225 189.275 ;
        RECT 64.405 189.065 64.735 189.445 ;
        RECT 64.055 188.725 64.720 188.895 ;
        RECT 64.915 188.770 65.175 189.275 ;
        RECT 62.525 188.205 62.855 188.455 ;
        RECT 63.985 188.175 64.315 188.545 ;
        RECT 64.550 188.470 64.720 188.725 ;
        RECT 64.550 188.140 64.835 188.470 ;
        RECT 60.740 187.565 61.490 187.735 ;
        RECT 60.735 186.895 61.065 187.395 ;
        RECT 61.235 187.065 61.490 187.565 ;
        RECT 61.725 186.895 61.935 188.035 ;
        RECT 62.105 187.065 62.435 188.045 ;
        RECT 62.605 186.895 62.835 188.035 ;
        RECT 63.045 186.895 63.335 188.060 ;
        RECT 64.550 187.995 64.720 188.140 ;
        RECT 64.055 187.825 64.720 187.995 ;
        RECT 65.005 187.970 65.175 188.770 ;
        RECT 64.055 187.065 64.225 187.825 ;
        RECT 64.405 186.895 64.735 187.655 ;
        RECT 64.905 187.065 65.175 187.970 ;
        RECT 65.345 188.705 65.730 189.275 ;
        RECT 65.900 188.985 66.225 189.445 ;
        RECT 66.745 188.815 67.025 189.275 ;
        RECT 65.345 188.035 65.625 188.705 ;
        RECT 65.900 188.645 67.025 188.815 ;
        RECT 65.900 188.535 66.350 188.645 ;
        RECT 65.795 188.205 66.350 188.535 ;
        RECT 67.215 188.475 67.615 189.275 ;
        RECT 68.015 188.985 68.285 189.445 ;
        RECT 68.455 188.815 68.740 189.275 ;
        RECT 65.345 187.065 65.730 188.035 ;
        RECT 65.900 187.745 66.350 188.205 ;
        RECT 66.520 187.915 67.615 188.475 ;
        RECT 65.900 187.525 67.025 187.745 ;
        RECT 65.900 186.895 66.225 187.355 ;
        RECT 66.745 187.065 67.025 187.525 ;
        RECT 67.215 187.065 67.615 187.915 ;
        RECT 67.785 188.645 68.740 188.815 ;
        RECT 69.025 188.705 69.410 189.275 ;
        RECT 69.580 188.985 69.905 189.445 ;
        RECT 70.425 188.815 70.705 189.275 ;
        RECT 67.785 187.745 67.995 188.645 ;
        RECT 68.165 187.915 68.855 188.475 ;
        RECT 69.025 188.035 69.305 188.705 ;
        RECT 69.580 188.645 70.705 188.815 ;
        RECT 69.580 188.535 70.030 188.645 ;
        RECT 69.475 188.205 70.030 188.535 ;
        RECT 70.895 188.475 71.295 189.275 ;
        RECT 71.695 188.985 71.965 189.445 ;
        RECT 72.135 188.815 72.420 189.275 ;
        RECT 73.225 188.975 73.525 189.445 ;
        RECT 67.785 187.525 68.740 187.745 ;
        RECT 68.015 186.895 68.285 187.355 ;
        RECT 68.455 187.065 68.740 187.525 ;
        RECT 69.025 187.065 69.410 188.035 ;
        RECT 69.580 187.745 70.030 188.205 ;
        RECT 70.200 187.915 71.295 188.475 ;
        RECT 69.580 187.525 70.705 187.745 ;
        RECT 69.580 186.895 69.905 187.355 ;
        RECT 70.425 187.065 70.705 187.525 ;
        RECT 70.895 187.065 71.295 187.915 ;
        RECT 71.465 188.645 72.420 188.815 ;
        RECT 73.695 188.805 73.950 189.250 ;
        RECT 74.120 188.975 74.380 189.445 ;
        RECT 74.550 188.805 74.810 189.250 ;
        RECT 74.980 188.975 75.275 189.445 ;
        RECT 75.985 188.965 76.265 189.445 ;
        RECT 71.465 187.745 71.675 188.645 ;
        RECT 72.705 188.635 75.735 188.805 ;
        RECT 76.435 188.795 76.695 189.185 ;
        RECT 76.870 188.965 77.125 189.445 ;
        RECT 77.295 188.795 77.590 189.185 ;
        RECT 77.770 188.965 78.045 189.445 ;
        RECT 78.215 188.945 78.515 189.275 ;
        RECT 78.955 189.050 79.285 189.445 ;
        RECT 71.845 187.915 72.535 188.475 ;
        RECT 72.705 188.070 73.005 188.635 ;
        RECT 73.180 188.240 75.395 188.465 ;
        RECT 75.565 188.070 75.735 188.635 ;
        RECT 72.705 187.900 75.735 188.070 ;
        RECT 75.940 188.625 77.590 188.795 ;
        RECT 75.940 188.115 76.345 188.625 ;
        RECT 76.515 188.285 77.655 188.455 ;
        RECT 75.940 187.945 76.695 188.115 ;
        RECT 71.465 187.525 72.420 187.745 ;
        RECT 71.695 186.895 71.965 187.355 ;
        RECT 72.135 187.065 72.420 187.525 ;
        RECT 72.705 186.895 73.090 187.730 ;
        RECT 73.260 187.095 73.520 187.900 ;
        RECT 73.690 186.895 73.950 187.730 ;
        RECT 74.120 187.095 74.375 187.900 ;
        RECT 74.550 186.895 74.810 187.730 ;
        RECT 74.980 187.095 75.235 187.900 ;
        RECT 75.410 186.895 75.755 187.730 ;
        RECT 75.980 186.895 76.265 187.765 ;
        RECT 76.435 187.695 76.695 187.945 ;
        RECT 77.485 188.035 77.655 188.285 ;
        RECT 77.825 188.205 78.175 188.775 ;
        RECT 78.345 188.035 78.515 188.945 ;
        RECT 79.455 188.875 79.655 189.230 ;
        RECT 79.825 189.045 80.155 189.445 ;
        RECT 80.325 188.875 80.525 189.220 ;
        RECT 77.485 187.865 78.515 188.035 ;
        RECT 76.435 187.525 77.555 187.695 ;
        RECT 76.435 187.065 76.695 187.525 ;
        RECT 76.870 186.895 77.125 187.355 ;
        RECT 77.295 187.065 77.555 187.525 ;
        RECT 77.725 186.895 78.035 187.695 ;
        RECT 78.205 187.065 78.515 187.865 ;
        RECT 78.685 188.705 80.525 188.875 ;
        RECT 80.695 188.705 81.025 189.445 ;
        RECT 81.260 188.875 81.430 189.125 ;
        RECT 81.260 188.705 81.735 188.875 ;
        RECT 78.685 187.080 78.945 188.705 ;
        RECT 79.125 187.735 79.345 188.535 ;
        RECT 79.585 187.915 79.885 188.535 ;
        RECT 80.055 187.915 80.385 188.535 ;
        RECT 80.555 187.915 80.875 188.535 ;
        RECT 81.045 187.915 81.395 188.535 ;
        RECT 81.565 187.735 81.735 188.705 ;
        RECT 81.995 188.795 82.165 189.275 ;
        RECT 82.345 188.965 82.585 189.445 ;
        RECT 82.835 188.795 83.005 189.275 ;
        RECT 83.175 188.965 83.505 189.445 ;
        RECT 83.675 188.795 83.845 189.275 ;
        RECT 81.995 188.625 82.630 188.795 ;
        RECT 82.835 188.625 83.845 188.795 ;
        RECT 84.015 188.645 84.345 189.445 ;
        RECT 84.940 188.635 85.185 189.240 ;
        RECT 85.405 188.910 85.915 189.445 ;
        RECT 82.460 188.455 82.630 188.625 ;
        RECT 83.345 188.595 83.845 188.625 ;
        RECT 81.910 188.215 82.290 188.455 ;
        RECT 82.460 188.285 82.960 188.455 ;
        RECT 82.460 188.045 82.630 188.285 ;
        RECT 83.350 188.085 83.845 188.595 ;
        RECT 79.125 187.525 81.735 187.735 ;
        RECT 81.915 187.875 82.630 188.045 ;
        RECT 82.835 187.915 83.845 188.085 ;
        RECT 84.665 188.465 85.895 188.635 ;
        RECT 80.695 186.895 81.025 187.345 ;
        RECT 81.915 187.065 82.245 187.875 ;
        RECT 82.415 186.895 82.655 187.695 ;
        RECT 82.835 187.065 83.005 187.915 ;
        RECT 83.175 186.895 83.505 187.695 ;
        RECT 83.675 187.065 83.845 187.915 ;
        RECT 84.015 186.895 84.345 188.045 ;
        RECT 84.665 187.655 85.005 188.465 ;
        RECT 85.175 187.900 85.925 188.090 ;
        RECT 84.665 187.245 85.180 187.655 ;
        RECT 85.415 186.895 85.585 187.655 ;
        RECT 85.755 187.235 85.925 187.900 ;
        RECT 86.095 187.915 86.285 189.275 ;
        RECT 86.455 188.765 86.730 189.275 ;
        RECT 86.920 188.910 87.450 189.275 ;
        RECT 87.875 189.045 88.205 189.445 ;
        RECT 87.275 188.875 87.450 188.910 ;
        RECT 86.455 188.595 86.735 188.765 ;
        RECT 86.455 188.115 86.730 188.595 ;
        RECT 86.935 187.915 87.105 188.715 ;
        RECT 86.095 187.745 87.105 187.915 ;
        RECT 87.275 188.705 88.205 188.875 ;
        RECT 88.375 188.705 88.630 189.275 ;
        RECT 88.805 188.720 89.095 189.445 ;
        RECT 90.185 188.935 90.490 189.445 ;
        RECT 87.275 187.575 87.445 188.705 ;
        RECT 88.035 188.535 88.205 188.705 ;
        RECT 86.320 187.405 87.445 187.575 ;
        RECT 87.615 188.205 87.810 188.535 ;
        RECT 88.035 188.205 88.290 188.535 ;
        RECT 87.615 187.235 87.785 188.205 ;
        RECT 88.460 188.035 88.630 188.705 ;
        RECT 90.185 188.205 90.500 188.765 ;
        RECT 90.670 188.455 90.920 189.265 ;
        RECT 91.090 188.920 91.350 189.445 ;
        RECT 91.530 188.455 91.780 189.265 ;
        RECT 91.950 188.885 92.210 189.445 ;
        RECT 92.380 188.795 92.640 189.250 ;
        RECT 92.810 188.965 93.070 189.445 ;
        RECT 93.240 188.795 93.500 189.250 ;
        RECT 93.670 188.965 93.930 189.445 ;
        RECT 94.100 188.795 94.360 189.250 ;
        RECT 94.530 188.965 94.775 189.445 ;
        RECT 94.945 188.795 95.220 189.250 ;
        RECT 95.390 188.965 95.635 189.445 ;
        RECT 95.805 188.795 96.065 189.250 ;
        RECT 96.245 188.965 96.495 189.445 ;
        RECT 96.665 188.795 96.925 189.250 ;
        RECT 97.105 188.965 97.355 189.445 ;
        RECT 97.525 188.795 97.785 189.250 ;
        RECT 97.965 188.965 98.225 189.445 ;
        RECT 98.395 188.795 98.655 189.250 ;
        RECT 98.825 188.965 99.125 189.445 ;
        RECT 92.380 188.625 99.125 188.795 ;
        RECT 90.670 188.205 97.790 188.455 ;
        RECT 85.755 187.065 87.785 187.235 ;
        RECT 87.955 186.895 88.125 188.035 ;
        RECT 88.295 187.065 88.630 188.035 ;
        RECT 88.805 186.895 89.095 188.060 ;
        RECT 90.195 186.895 90.490 187.705 ;
        RECT 90.670 187.065 90.915 188.205 ;
        RECT 91.090 186.895 91.350 187.705 ;
        RECT 91.530 187.070 91.780 188.205 ;
        RECT 97.960 188.035 99.125 188.625 ;
        RECT 92.380 187.810 99.125 188.035 ;
        RECT 99.390 188.735 99.645 189.265 ;
        RECT 99.815 188.985 100.120 189.445 ;
        RECT 100.365 189.065 101.435 189.235 ;
        RECT 99.390 188.085 99.600 188.735 ;
        RECT 100.365 188.710 100.685 189.065 ;
        RECT 100.360 188.535 100.685 188.710 ;
        RECT 99.770 188.235 100.685 188.535 ;
        RECT 100.855 188.495 101.095 188.895 ;
        RECT 101.265 188.835 101.435 189.065 ;
        RECT 101.605 189.005 101.795 189.445 ;
        RECT 101.965 188.995 102.915 189.275 ;
        RECT 103.135 189.085 103.485 189.255 ;
        RECT 101.265 188.665 101.795 188.835 ;
        RECT 99.770 188.205 100.510 188.235 ;
        RECT 92.380 187.795 97.785 187.810 ;
        RECT 91.950 186.900 92.210 187.695 ;
        RECT 92.380 187.070 92.640 187.795 ;
        RECT 92.810 186.900 93.070 187.625 ;
        RECT 93.240 187.070 93.500 187.795 ;
        RECT 93.670 186.900 93.930 187.625 ;
        RECT 94.100 187.070 94.360 187.795 ;
        RECT 94.530 186.900 94.790 187.625 ;
        RECT 94.960 187.070 95.220 187.795 ;
        RECT 95.390 186.900 95.635 187.625 ;
        RECT 95.805 187.070 96.065 187.795 ;
        RECT 96.250 186.900 96.495 187.625 ;
        RECT 96.665 187.070 96.925 187.795 ;
        RECT 97.110 186.900 97.355 187.625 ;
        RECT 97.525 187.070 97.785 187.795 ;
        RECT 97.970 186.900 98.225 187.625 ;
        RECT 98.395 187.070 98.685 187.810 ;
        RECT 91.950 186.895 98.225 186.900 ;
        RECT 98.855 186.895 99.125 187.640 ;
        RECT 99.390 187.205 99.645 188.085 ;
        RECT 99.815 186.895 100.120 188.035 ;
        RECT 100.340 187.615 100.510 188.205 ;
        RECT 100.855 188.125 101.395 188.495 ;
        RECT 101.575 188.385 101.795 188.665 ;
        RECT 101.965 188.215 102.135 188.995 ;
        RECT 101.730 188.045 102.135 188.215 ;
        RECT 102.305 188.205 102.655 188.825 ;
        RECT 101.730 187.955 101.900 188.045 ;
        RECT 102.825 188.035 103.035 188.825 ;
        RECT 100.680 187.785 101.900 187.955 ;
        RECT 102.360 187.875 103.035 188.035 ;
        RECT 100.340 187.445 101.140 187.615 ;
        RECT 100.460 186.895 100.790 187.275 ;
        RECT 100.970 187.155 101.140 187.445 ;
        RECT 101.730 187.405 101.900 187.785 ;
        RECT 102.070 187.865 103.035 187.875 ;
        RECT 103.225 188.695 103.485 189.085 ;
        RECT 103.695 188.985 104.025 189.445 ;
        RECT 104.900 189.055 105.755 189.225 ;
        RECT 105.960 189.055 106.455 189.225 ;
        RECT 106.625 189.085 106.955 189.445 ;
        RECT 103.225 188.005 103.395 188.695 ;
        RECT 103.565 188.345 103.735 188.525 ;
        RECT 103.905 188.515 104.695 188.765 ;
        RECT 104.900 188.345 105.070 189.055 ;
        RECT 105.240 188.545 105.595 188.765 ;
        RECT 103.565 188.175 105.255 188.345 ;
        RECT 102.070 187.575 102.530 187.865 ;
        RECT 103.225 187.835 104.725 188.005 ;
        RECT 103.225 187.695 103.395 187.835 ;
        RECT 102.835 187.525 103.395 187.695 ;
        RECT 101.310 186.895 101.560 187.355 ;
        RECT 101.730 187.065 102.600 187.405 ;
        RECT 102.835 187.065 103.005 187.525 ;
        RECT 103.840 187.495 104.915 187.665 ;
        RECT 103.175 186.895 103.545 187.355 ;
        RECT 103.840 187.155 104.010 187.495 ;
        RECT 104.180 186.895 104.510 187.325 ;
        RECT 104.745 187.155 104.915 187.495 ;
        RECT 105.085 187.395 105.255 188.175 ;
        RECT 105.425 187.955 105.595 188.545 ;
        RECT 105.765 188.145 106.115 188.765 ;
        RECT 105.425 187.565 105.890 187.955 ;
        RECT 106.285 187.695 106.455 189.055 ;
        RECT 106.625 187.865 107.085 188.915 ;
        RECT 106.060 187.525 106.455 187.695 ;
        RECT 106.060 187.395 106.230 187.525 ;
        RECT 105.085 187.065 105.765 187.395 ;
        RECT 105.980 187.065 106.230 187.395 ;
        RECT 106.400 186.895 106.650 187.355 ;
        RECT 106.820 187.080 107.145 187.865 ;
        RECT 107.315 187.065 107.485 189.185 ;
        RECT 107.655 189.065 107.985 189.445 ;
        RECT 108.155 188.895 108.410 189.185 ;
        RECT 107.660 188.725 108.410 188.895 ;
        RECT 107.660 187.735 107.890 188.725 ;
        RECT 108.590 188.705 108.845 189.275 ;
        RECT 109.015 189.045 109.345 189.445 ;
        RECT 109.770 188.910 110.300 189.275 ;
        RECT 110.490 189.105 110.765 189.275 ;
        RECT 110.485 188.935 110.765 189.105 ;
        RECT 109.770 188.875 109.945 188.910 ;
        RECT 109.015 188.705 109.945 188.875 ;
        RECT 108.060 187.905 108.410 188.555 ;
        RECT 108.590 188.035 108.760 188.705 ;
        RECT 109.015 188.535 109.185 188.705 ;
        RECT 108.930 188.205 109.185 188.535 ;
        RECT 109.410 188.205 109.605 188.535 ;
        RECT 107.660 187.565 108.410 187.735 ;
        RECT 107.655 186.895 107.985 187.395 ;
        RECT 108.155 187.065 108.410 187.565 ;
        RECT 108.590 187.065 108.925 188.035 ;
        RECT 109.095 186.895 109.265 188.035 ;
        RECT 109.435 187.235 109.605 188.205 ;
        RECT 109.775 187.575 109.945 188.705 ;
        RECT 110.115 187.915 110.285 188.715 ;
        RECT 110.490 188.115 110.765 188.935 ;
        RECT 110.935 187.915 111.125 189.275 ;
        RECT 111.305 188.910 111.815 189.445 ;
        RECT 112.035 188.635 112.280 189.240 ;
        RECT 111.325 188.465 112.555 188.635 ;
        RECT 112.765 188.625 112.995 189.445 ;
        RECT 113.165 188.645 113.495 189.275 ;
        RECT 110.115 187.745 111.125 187.915 ;
        RECT 111.295 187.900 112.045 188.090 ;
        RECT 109.775 187.405 110.900 187.575 ;
        RECT 111.295 187.235 111.465 187.900 ;
        RECT 112.215 187.655 112.555 188.465 ;
        RECT 112.745 188.205 113.075 188.455 ;
        RECT 113.245 188.045 113.495 188.645 ;
        RECT 113.665 188.625 113.875 189.445 ;
        RECT 114.565 188.720 114.855 189.445 ;
        RECT 115.030 188.735 115.285 189.265 ;
        RECT 115.455 188.985 115.760 189.445 ;
        RECT 116.005 189.065 117.075 189.235 ;
        RECT 115.030 188.085 115.240 188.735 ;
        RECT 116.005 188.710 116.325 189.065 ;
        RECT 116.000 188.535 116.325 188.710 ;
        RECT 115.410 188.235 116.325 188.535 ;
        RECT 116.495 188.495 116.735 188.895 ;
        RECT 116.905 188.835 117.075 189.065 ;
        RECT 117.245 189.005 117.435 189.445 ;
        RECT 117.605 188.995 118.555 189.275 ;
        RECT 118.775 189.085 119.125 189.255 ;
        RECT 116.905 188.665 117.435 188.835 ;
        RECT 115.410 188.205 116.150 188.235 ;
        RECT 109.435 187.065 111.465 187.235 ;
        RECT 111.635 186.895 111.805 187.655 ;
        RECT 112.040 187.245 112.555 187.655 ;
        RECT 112.765 186.895 112.995 188.035 ;
        RECT 113.165 187.065 113.495 188.045 ;
        RECT 113.665 186.895 113.875 188.035 ;
        RECT 114.565 186.895 114.855 188.060 ;
        RECT 115.030 187.205 115.285 188.085 ;
        RECT 115.455 186.895 115.760 188.035 ;
        RECT 115.980 187.615 116.150 188.205 ;
        RECT 116.495 188.125 117.035 188.495 ;
        RECT 117.215 188.385 117.435 188.665 ;
        RECT 117.605 188.215 117.775 188.995 ;
        RECT 117.370 188.045 117.775 188.215 ;
        RECT 117.945 188.205 118.295 188.825 ;
        RECT 117.370 187.955 117.540 188.045 ;
        RECT 118.465 188.035 118.675 188.825 ;
        RECT 116.320 187.785 117.540 187.955 ;
        RECT 118.000 187.875 118.675 188.035 ;
        RECT 115.980 187.445 116.780 187.615 ;
        RECT 116.100 186.895 116.430 187.275 ;
        RECT 116.610 187.155 116.780 187.445 ;
        RECT 117.370 187.405 117.540 187.785 ;
        RECT 117.710 187.865 118.675 187.875 ;
        RECT 118.865 188.695 119.125 189.085 ;
        RECT 119.335 188.985 119.665 189.445 ;
        RECT 120.540 189.055 121.395 189.225 ;
        RECT 121.600 189.055 122.095 189.225 ;
        RECT 122.265 189.085 122.595 189.445 ;
        RECT 118.865 188.005 119.035 188.695 ;
        RECT 119.205 188.345 119.375 188.525 ;
        RECT 119.545 188.515 120.335 188.765 ;
        RECT 120.540 188.345 120.710 189.055 ;
        RECT 120.880 188.545 121.235 188.765 ;
        RECT 119.205 188.175 120.895 188.345 ;
        RECT 117.710 187.575 118.170 187.865 ;
        RECT 118.865 187.835 120.365 188.005 ;
        RECT 118.865 187.695 119.035 187.835 ;
        RECT 118.475 187.525 119.035 187.695 ;
        RECT 116.950 186.895 117.200 187.355 ;
        RECT 117.370 187.065 118.240 187.405 ;
        RECT 118.475 187.065 118.645 187.525 ;
        RECT 119.480 187.495 120.555 187.665 ;
        RECT 118.815 186.895 119.185 187.355 ;
        RECT 119.480 187.155 119.650 187.495 ;
        RECT 119.820 186.895 120.150 187.325 ;
        RECT 120.385 187.155 120.555 187.495 ;
        RECT 120.725 187.395 120.895 188.175 ;
        RECT 121.065 187.955 121.235 188.545 ;
        RECT 121.405 188.145 121.755 188.765 ;
        RECT 121.065 187.565 121.530 187.955 ;
        RECT 121.925 187.695 122.095 189.055 ;
        RECT 122.265 187.865 122.725 188.915 ;
        RECT 121.700 187.525 122.095 187.695 ;
        RECT 121.700 187.395 121.870 187.525 ;
        RECT 120.725 187.065 121.405 187.395 ;
        RECT 121.620 187.065 121.870 187.395 ;
        RECT 122.040 186.895 122.290 187.355 ;
        RECT 122.460 187.080 122.785 187.865 ;
        RECT 122.955 187.065 123.125 189.185 ;
        RECT 123.295 189.065 123.625 189.445 ;
        RECT 123.795 188.895 124.050 189.185 ;
        RECT 123.300 188.725 124.050 188.895 ;
        RECT 123.300 187.735 123.530 188.725 ;
        RECT 124.685 188.675 126.355 189.445 ;
        RECT 126.525 188.695 127.735 189.445 ;
        RECT 123.700 187.905 124.050 188.555 ;
        RECT 124.685 187.985 125.435 188.505 ;
        RECT 125.605 188.155 126.355 188.675 ;
        RECT 126.525 187.985 127.045 188.525 ;
        RECT 127.215 188.155 127.735 188.695 ;
        RECT 123.300 187.565 124.050 187.735 ;
        RECT 123.295 186.895 123.625 187.395 ;
        RECT 123.795 187.065 124.050 187.565 ;
        RECT 124.685 186.895 126.355 187.985 ;
        RECT 126.525 186.895 127.735 187.985 ;
        RECT 29.840 186.725 127.820 186.895 ;
        RECT 29.925 185.635 31.135 186.725 ;
        RECT 31.420 186.095 31.705 186.555 ;
        RECT 31.875 186.265 32.145 186.725 ;
        RECT 31.420 185.875 32.375 186.095 ;
        RECT 29.925 184.925 30.445 185.465 ;
        RECT 30.615 185.095 31.135 185.635 ;
        RECT 31.305 185.145 31.995 185.705 ;
        RECT 32.165 184.975 32.375 185.875 ;
        RECT 29.925 184.175 31.135 184.925 ;
        RECT 31.420 184.805 32.375 184.975 ;
        RECT 32.545 185.705 32.945 186.555 ;
        RECT 33.135 186.095 33.415 186.555 ;
        RECT 33.935 186.265 34.260 186.725 ;
        RECT 33.135 185.875 34.260 186.095 ;
        RECT 32.545 185.145 33.640 185.705 ;
        RECT 33.810 185.415 34.260 185.875 ;
        RECT 34.430 185.585 34.815 186.555 ;
        RECT 31.420 184.345 31.705 184.805 ;
        RECT 31.875 184.175 32.145 184.635 ;
        RECT 32.545 184.345 32.945 185.145 ;
        RECT 33.810 185.085 34.365 185.415 ;
        RECT 33.810 184.975 34.260 185.085 ;
        RECT 33.135 184.805 34.260 184.975 ;
        RECT 34.535 184.915 34.815 185.585 ;
        RECT 33.135 184.345 33.415 184.805 ;
        RECT 33.935 184.175 34.260 184.635 ;
        RECT 34.430 184.345 34.815 184.915 ;
        RECT 34.990 185.535 35.245 186.415 ;
        RECT 35.415 185.585 35.720 186.725 ;
        RECT 36.060 186.345 36.390 186.725 ;
        RECT 36.570 186.175 36.740 186.465 ;
        RECT 36.910 186.265 37.160 186.725 ;
        RECT 35.940 186.005 36.740 186.175 ;
        RECT 37.330 186.215 38.200 186.555 ;
        RECT 34.990 184.885 35.200 185.535 ;
        RECT 35.940 185.415 36.110 186.005 ;
        RECT 37.330 185.835 37.500 186.215 ;
        RECT 38.435 186.095 38.605 186.555 ;
        RECT 38.775 186.265 39.145 186.725 ;
        RECT 39.440 186.125 39.610 186.465 ;
        RECT 39.780 186.295 40.110 186.725 ;
        RECT 40.345 186.125 40.515 186.465 ;
        RECT 36.280 185.665 37.500 185.835 ;
        RECT 37.670 185.755 38.130 186.045 ;
        RECT 38.435 185.925 38.995 186.095 ;
        RECT 39.440 185.955 40.515 186.125 ;
        RECT 40.685 186.225 41.365 186.555 ;
        RECT 41.580 186.225 41.830 186.555 ;
        RECT 42.000 186.265 42.250 186.725 ;
        RECT 38.825 185.785 38.995 185.925 ;
        RECT 37.670 185.745 38.635 185.755 ;
        RECT 37.330 185.575 37.500 185.665 ;
        RECT 37.960 185.585 38.635 185.745 ;
        RECT 35.370 185.385 36.110 185.415 ;
        RECT 35.370 185.085 36.285 185.385 ;
        RECT 35.960 184.910 36.285 185.085 ;
        RECT 34.990 184.355 35.245 184.885 ;
        RECT 35.415 184.175 35.720 184.635 ;
        RECT 35.965 184.555 36.285 184.910 ;
        RECT 36.455 185.125 36.995 185.495 ;
        RECT 37.330 185.405 37.735 185.575 ;
        RECT 36.455 184.725 36.695 185.125 ;
        RECT 37.175 184.955 37.395 185.235 ;
        RECT 36.865 184.785 37.395 184.955 ;
        RECT 36.865 184.555 37.035 184.785 ;
        RECT 37.565 184.625 37.735 185.405 ;
        RECT 37.905 184.795 38.255 185.415 ;
        RECT 38.425 184.795 38.635 185.585 ;
        RECT 38.825 185.615 40.325 185.785 ;
        RECT 38.825 184.925 38.995 185.615 ;
        RECT 40.685 185.445 40.855 186.225 ;
        RECT 41.660 186.095 41.830 186.225 ;
        RECT 39.165 185.275 40.855 185.445 ;
        RECT 41.025 185.665 41.490 186.055 ;
        RECT 41.660 185.925 42.055 186.095 ;
        RECT 39.165 185.095 39.335 185.275 ;
        RECT 35.965 184.385 37.035 184.555 ;
        RECT 37.205 184.175 37.395 184.615 ;
        RECT 37.565 184.345 38.515 184.625 ;
        RECT 38.825 184.535 39.085 184.925 ;
        RECT 39.505 184.855 40.295 185.105 ;
        RECT 38.735 184.365 39.085 184.535 ;
        RECT 39.295 184.175 39.625 184.635 ;
        RECT 40.500 184.565 40.670 185.275 ;
        RECT 41.025 185.075 41.195 185.665 ;
        RECT 40.840 184.855 41.195 185.075 ;
        RECT 41.365 184.855 41.715 185.475 ;
        RECT 41.885 184.565 42.055 185.925 ;
        RECT 42.420 185.755 42.745 186.540 ;
        RECT 42.225 184.705 42.685 185.755 ;
        RECT 40.500 184.395 41.355 184.565 ;
        RECT 41.560 184.395 42.055 184.565 ;
        RECT 42.225 184.175 42.555 184.535 ;
        RECT 42.915 184.435 43.085 186.555 ;
        RECT 43.255 186.225 43.585 186.725 ;
        RECT 43.755 186.055 44.010 186.555 ;
        RECT 43.260 185.885 44.010 186.055 ;
        RECT 44.185 185.965 44.700 186.375 ;
        RECT 44.935 185.965 45.105 186.725 ;
        RECT 45.275 186.385 47.305 186.555 ;
        RECT 43.260 184.895 43.490 185.885 ;
        RECT 43.660 185.065 44.010 185.715 ;
        RECT 44.185 185.155 44.525 185.965 ;
        RECT 45.275 185.720 45.445 186.385 ;
        RECT 45.840 186.045 46.965 186.215 ;
        RECT 44.695 185.530 45.445 185.720 ;
        RECT 45.615 185.705 46.625 185.875 ;
        RECT 44.185 184.985 45.415 185.155 ;
        RECT 43.260 184.725 44.010 184.895 ;
        RECT 43.255 184.175 43.585 184.555 ;
        RECT 43.755 184.435 44.010 184.725 ;
        RECT 44.460 184.380 44.705 184.985 ;
        RECT 44.925 184.175 45.435 184.710 ;
        RECT 45.615 184.345 45.805 185.705 ;
        RECT 45.975 184.685 46.250 185.505 ;
        RECT 46.455 184.905 46.625 185.705 ;
        RECT 46.795 184.915 46.965 186.045 ;
        RECT 47.135 185.415 47.305 186.385 ;
        RECT 47.475 185.585 47.645 186.725 ;
        RECT 47.815 185.585 48.150 186.555 ;
        RECT 48.825 185.585 49.055 186.725 ;
        RECT 47.135 185.085 47.330 185.415 ;
        RECT 47.555 185.085 47.810 185.415 ;
        RECT 47.555 184.915 47.725 185.085 ;
        RECT 47.980 184.915 48.150 185.585 ;
        RECT 49.225 185.575 49.555 186.555 ;
        RECT 49.725 185.585 49.935 186.725 ;
        RECT 48.805 185.165 49.135 185.415 ;
        RECT 46.795 184.745 47.725 184.915 ;
        RECT 46.795 184.710 46.970 184.745 ;
        RECT 45.975 184.515 46.255 184.685 ;
        RECT 45.975 184.345 46.250 184.515 ;
        RECT 46.440 184.345 46.970 184.710 ;
        RECT 47.395 184.175 47.725 184.575 ;
        RECT 47.895 184.345 48.150 184.915 ;
        RECT 48.825 184.175 49.055 184.995 ;
        RECT 49.305 184.975 49.555 185.575 ;
        RECT 50.165 185.560 50.455 186.725 ;
        RECT 51.660 186.095 51.945 186.555 ;
        RECT 52.115 186.265 52.385 186.725 ;
        RECT 51.660 185.875 52.615 186.095 ;
        RECT 51.545 185.145 52.235 185.705 ;
        RECT 49.225 184.345 49.555 184.975 ;
        RECT 49.725 184.175 49.935 184.995 ;
        RECT 52.405 184.975 52.615 185.875 ;
        RECT 50.165 184.175 50.455 184.900 ;
        RECT 51.660 184.805 52.615 184.975 ;
        RECT 52.785 185.705 53.185 186.555 ;
        RECT 53.375 186.095 53.655 186.555 ;
        RECT 54.175 186.265 54.500 186.725 ;
        RECT 53.375 185.875 54.500 186.095 ;
        RECT 52.785 185.145 53.880 185.705 ;
        RECT 54.050 185.415 54.500 185.875 ;
        RECT 54.670 185.585 55.055 186.555 ;
        RECT 55.430 185.755 55.760 186.555 ;
        RECT 55.930 185.925 56.260 186.725 ;
        RECT 56.560 185.755 56.890 186.555 ;
        RECT 57.535 185.925 57.785 186.725 ;
        RECT 55.430 185.585 57.865 185.755 ;
        RECT 58.055 185.585 58.225 186.725 ;
        RECT 58.395 185.585 58.735 186.555 ;
        RECT 58.995 185.980 59.265 186.725 ;
        RECT 59.895 186.720 66.170 186.725 ;
        RECT 59.435 185.810 59.725 186.550 ;
        RECT 59.895 185.995 60.150 186.720 ;
        RECT 60.335 185.825 60.595 186.550 ;
        RECT 60.765 185.995 61.010 186.720 ;
        RECT 61.195 185.825 61.455 186.550 ;
        RECT 61.625 185.995 61.870 186.720 ;
        RECT 62.055 185.825 62.315 186.550 ;
        RECT 62.485 185.995 62.730 186.720 ;
        RECT 62.900 185.825 63.160 186.550 ;
        RECT 63.330 185.995 63.590 186.720 ;
        RECT 63.760 185.825 64.020 186.550 ;
        RECT 64.190 185.995 64.450 186.720 ;
        RECT 64.620 185.825 64.880 186.550 ;
        RECT 65.050 185.995 65.310 186.720 ;
        RECT 65.480 185.825 65.740 186.550 ;
        RECT 65.910 185.925 66.170 186.720 ;
        RECT 60.335 185.810 65.740 185.825 ;
        RECT 51.660 184.345 51.945 184.805 ;
        RECT 52.115 184.175 52.385 184.635 ;
        RECT 52.785 184.345 53.185 185.145 ;
        RECT 54.050 185.085 54.605 185.415 ;
        RECT 54.050 184.975 54.500 185.085 ;
        RECT 53.375 184.805 54.500 184.975 ;
        RECT 54.775 184.915 55.055 185.585 ;
        RECT 55.225 185.165 55.575 185.415 ;
        RECT 55.760 184.955 55.930 185.585 ;
        RECT 56.100 185.165 56.430 185.365 ;
        RECT 56.600 185.165 56.930 185.365 ;
        RECT 57.100 185.165 57.520 185.365 ;
        RECT 57.695 185.335 57.865 185.585 ;
        RECT 57.695 185.165 58.390 185.335 ;
        RECT 53.375 184.345 53.655 184.805 ;
        RECT 54.175 184.175 54.500 184.635 ;
        RECT 54.670 184.345 55.055 184.915 ;
        RECT 55.430 184.345 55.930 184.955 ;
        RECT 56.560 184.825 57.785 184.995 ;
        RECT 58.560 184.975 58.735 185.585 ;
        RECT 56.560 184.345 56.890 184.825 ;
        RECT 57.060 184.175 57.285 184.635 ;
        RECT 57.455 184.345 57.785 184.825 ;
        RECT 57.975 184.175 58.225 184.975 ;
        RECT 58.395 184.345 58.735 184.975 ;
        RECT 58.995 185.585 65.740 185.810 ;
        RECT 58.995 184.995 60.160 185.585 ;
        RECT 66.340 185.415 66.590 186.550 ;
        RECT 66.770 185.915 67.030 186.725 ;
        RECT 67.205 185.415 67.450 186.555 ;
        RECT 67.630 185.915 67.925 186.725 ;
        RECT 68.105 185.965 68.620 186.375 ;
        RECT 68.855 185.965 69.025 186.725 ;
        RECT 69.195 186.385 71.225 186.555 ;
        RECT 60.330 185.165 67.450 185.415 ;
        RECT 58.995 184.825 65.740 184.995 ;
        RECT 58.995 184.175 59.295 184.655 ;
        RECT 59.465 184.370 59.725 184.825 ;
        RECT 59.895 184.175 60.155 184.655 ;
        RECT 60.335 184.370 60.595 184.825 ;
        RECT 60.765 184.175 61.015 184.655 ;
        RECT 61.195 184.370 61.455 184.825 ;
        RECT 61.625 184.175 61.875 184.655 ;
        RECT 62.055 184.370 62.315 184.825 ;
        RECT 62.485 184.175 62.730 184.655 ;
        RECT 62.900 184.370 63.175 184.825 ;
        RECT 63.345 184.175 63.590 184.655 ;
        RECT 63.760 184.370 64.020 184.825 ;
        RECT 64.190 184.175 64.450 184.655 ;
        RECT 64.620 184.370 64.880 184.825 ;
        RECT 65.050 184.175 65.310 184.655 ;
        RECT 65.480 184.370 65.740 184.825 ;
        RECT 65.910 184.175 66.170 184.735 ;
        RECT 66.340 184.355 66.590 185.165 ;
        RECT 66.770 184.175 67.030 184.700 ;
        RECT 67.200 184.355 67.450 185.165 ;
        RECT 67.620 184.855 67.935 185.415 ;
        RECT 68.105 185.155 68.445 185.965 ;
        RECT 69.195 185.720 69.365 186.385 ;
        RECT 69.760 186.045 70.885 186.215 ;
        RECT 68.615 185.530 69.365 185.720 ;
        RECT 69.535 185.705 70.545 185.875 ;
        RECT 68.105 184.985 69.335 185.155 ;
        RECT 67.630 184.175 67.935 184.685 ;
        RECT 68.380 184.380 68.625 184.985 ;
        RECT 68.845 184.175 69.355 184.710 ;
        RECT 69.535 184.345 69.725 185.705 ;
        RECT 69.895 185.365 70.170 185.505 ;
        RECT 69.895 185.195 70.175 185.365 ;
        RECT 69.895 184.345 70.170 185.195 ;
        RECT 70.375 184.905 70.545 185.705 ;
        RECT 70.715 184.915 70.885 186.045 ;
        RECT 71.055 185.415 71.225 186.385 ;
        RECT 71.395 185.585 71.565 186.725 ;
        RECT 71.735 185.585 72.070 186.555 ;
        RECT 71.055 185.085 71.250 185.415 ;
        RECT 71.475 185.085 71.730 185.415 ;
        RECT 71.475 184.915 71.645 185.085 ;
        RECT 71.900 184.915 72.070 185.585 ;
        RECT 70.715 184.745 71.645 184.915 ;
        RECT 70.715 184.710 70.890 184.745 ;
        RECT 70.360 184.345 70.890 184.710 ;
        RECT 71.315 184.175 71.645 184.575 ;
        RECT 71.815 184.345 72.070 184.915 ;
        RECT 72.245 185.585 72.630 186.555 ;
        RECT 72.800 186.265 73.125 186.725 ;
        RECT 73.645 186.095 73.925 186.555 ;
        RECT 72.800 185.875 73.925 186.095 ;
        RECT 72.245 184.915 72.525 185.585 ;
        RECT 72.800 185.415 73.250 185.875 ;
        RECT 74.115 185.705 74.515 186.555 ;
        RECT 74.915 186.265 75.185 186.725 ;
        RECT 75.355 186.095 75.640 186.555 ;
        RECT 72.695 185.085 73.250 185.415 ;
        RECT 73.420 185.145 74.515 185.705 ;
        RECT 72.800 184.975 73.250 185.085 ;
        RECT 72.245 184.345 72.630 184.915 ;
        RECT 72.800 184.805 73.925 184.975 ;
        RECT 72.800 184.175 73.125 184.635 ;
        RECT 73.645 184.345 73.925 184.805 ;
        RECT 74.115 184.345 74.515 185.145 ;
        RECT 74.685 185.875 75.640 186.095 ;
        RECT 74.685 184.975 74.895 185.875 ;
        RECT 75.065 185.145 75.755 185.705 ;
        RECT 75.925 185.560 76.215 186.725 ;
        RECT 76.440 185.855 76.725 186.725 ;
        RECT 76.895 186.095 77.155 186.555 ;
        RECT 77.330 186.265 77.585 186.725 ;
        RECT 77.755 186.095 78.015 186.555 ;
        RECT 76.895 185.925 78.015 186.095 ;
        RECT 78.185 185.925 78.495 186.725 ;
        RECT 76.895 185.675 77.155 185.925 ;
        RECT 78.665 185.755 78.975 186.555 ;
        RECT 76.400 185.505 77.155 185.675 ;
        RECT 77.945 185.585 78.975 185.755 ;
        RECT 79.235 185.795 79.405 186.555 ;
        RECT 79.620 185.965 79.950 186.725 ;
        RECT 79.235 185.625 79.950 185.795 ;
        RECT 80.120 185.650 80.375 186.555 ;
        RECT 76.400 184.995 76.805 185.505 ;
        RECT 77.945 185.335 78.115 185.585 ;
        RECT 76.975 185.165 78.115 185.335 ;
        RECT 74.685 184.805 75.640 184.975 ;
        RECT 74.915 184.175 75.185 184.635 ;
        RECT 75.355 184.345 75.640 184.805 ;
        RECT 75.925 184.175 76.215 184.900 ;
        RECT 76.400 184.825 78.050 184.995 ;
        RECT 78.285 184.845 78.635 185.415 ;
        RECT 76.445 184.175 76.725 184.655 ;
        RECT 76.895 184.435 77.155 184.825 ;
        RECT 77.330 184.175 77.585 184.655 ;
        RECT 77.755 184.435 78.050 184.825 ;
        RECT 78.805 184.675 78.975 185.585 ;
        RECT 79.145 185.075 79.500 185.445 ;
        RECT 79.780 185.415 79.950 185.625 ;
        RECT 79.780 185.085 80.035 185.415 ;
        RECT 79.780 184.895 79.950 185.085 ;
        RECT 80.205 184.920 80.375 185.650 ;
        RECT 80.550 185.575 80.810 186.725 ;
        RECT 81.445 185.585 81.785 186.555 ;
        RECT 81.955 185.585 82.125 186.725 ;
        RECT 82.395 185.925 82.645 186.725 ;
        RECT 83.290 185.755 83.620 186.555 ;
        RECT 83.920 185.925 84.250 186.725 ;
        RECT 84.420 185.755 84.750 186.555 ;
        RECT 82.315 185.585 84.750 185.755 ;
        RECT 85.125 185.965 85.640 186.375 ;
        RECT 85.875 185.965 86.045 186.725 ;
        RECT 86.215 186.385 88.245 186.555 ;
        RECT 78.230 184.175 78.505 184.655 ;
        RECT 78.675 184.345 78.975 184.675 ;
        RECT 79.235 184.725 79.950 184.895 ;
        RECT 79.235 184.345 79.405 184.725 ;
        RECT 79.620 184.175 79.950 184.555 ;
        RECT 80.120 184.345 80.375 184.920 ;
        RECT 80.550 184.175 80.810 185.015 ;
        RECT 81.445 184.975 81.620 185.585 ;
        RECT 82.315 185.335 82.485 185.585 ;
        RECT 81.790 185.165 82.485 185.335 ;
        RECT 82.660 185.165 83.080 185.365 ;
        RECT 83.250 185.165 83.580 185.365 ;
        RECT 83.750 185.165 84.080 185.365 ;
        RECT 81.445 184.345 81.785 184.975 ;
        RECT 81.955 184.175 82.205 184.975 ;
        RECT 82.395 184.825 83.620 184.995 ;
        RECT 82.395 184.345 82.725 184.825 ;
        RECT 82.895 184.175 83.120 184.635 ;
        RECT 83.290 184.345 83.620 184.825 ;
        RECT 84.250 184.955 84.420 185.585 ;
        RECT 84.605 185.165 84.955 185.415 ;
        RECT 85.125 185.155 85.465 185.965 ;
        RECT 86.215 185.720 86.385 186.385 ;
        RECT 86.780 186.045 87.905 186.215 ;
        RECT 85.635 185.530 86.385 185.720 ;
        RECT 86.555 185.705 87.565 185.875 ;
        RECT 85.125 184.985 86.355 185.155 ;
        RECT 84.250 184.345 84.750 184.955 ;
        RECT 85.400 184.380 85.645 184.985 ;
        RECT 85.865 184.175 86.375 184.710 ;
        RECT 86.555 184.345 86.745 185.705 ;
        RECT 86.915 184.685 87.190 185.505 ;
        RECT 87.395 184.905 87.565 185.705 ;
        RECT 87.735 184.915 87.905 186.045 ;
        RECT 88.075 185.415 88.245 186.385 ;
        RECT 88.415 185.585 88.585 186.725 ;
        RECT 88.755 185.585 89.090 186.555 ;
        RECT 88.075 185.085 88.270 185.415 ;
        RECT 88.495 185.085 88.750 185.415 ;
        RECT 88.495 184.915 88.665 185.085 ;
        RECT 88.920 184.915 89.090 185.585 ;
        RECT 87.735 184.745 88.665 184.915 ;
        RECT 87.735 184.710 87.910 184.745 ;
        RECT 86.915 184.515 87.195 184.685 ;
        RECT 86.915 184.345 87.190 184.515 ;
        RECT 87.380 184.345 87.910 184.710 ;
        RECT 88.335 184.175 88.665 184.575 ;
        RECT 88.835 184.345 89.090 184.915 ;
        RECT 89.270 185.535 89.525 186.415 ;
        RECT 89.695 185.585 90.000 186.725 ;
        RECT 90.340 186.345 90.670 186.725 ;
        RECT 90.850 186.175 91.020 186.465 ;
        RECT 91.190 186.265 91.440 186.725 ;
        RECT 90.220 186.005 91.020 186.175 ;
        RECT 91.610 186.215 92.480 186.555 ;
        RECT 89.270 184.885 89.480 185.535 ;
        RECT 90.220 185.415 90.390 186.005 ;
        RECT 91.610 185.835 91.780 186.215 ;
        RECT 92.715 186.095 92.885 186.555 ;
        RECT 93.055 186.265 93.425 186.725 ;
        RECT 93.720 186.125 93.890 186.465 ;
        RECT 94.060 186.295 94.390 186.725 ;
        RECT 94.625 186.125 94.795 186.465 ;
        RECT 90.560 185.665 91.780 185.835 ;
        RECT 91.950 185.755 92.410 186.045 ;
        RECT 92.715 185.925 93.275 186.095 ;
        RECT 93.720 185.955 94.795 186.125 ;
        RECT 94.965 186.225 95.645 186.555 ;
        RECT 95.860 186.225 96.110 186.555 ;
        RECT 96.280 186.265 96.530 186.725 ;
        RECT 93.105 185.785 93.275 185.925 ;
        RECT 91.950 185.745 92.915 185.755 ;
        RECT 91.610 185.575 91.780 185.665 ;
        RECT 92.240 185.585 92.915 185.745 ;
        RECT 89.650 185.385 90.390 185.415 ;
        RECT 89.650 185.085 90.565 185.385 ;
        RECT 90.240 184.910 90.565 185.085 ;
        RECT 89.270 184.355 89.525 184.885 ;
        RECT 89.695 184.175 90.000 184.635 ;
        RECT 90.245 184.555 90.565 184.910 ;
        RECT 90.735 185.125 91.275 185.495 ;
        RECT 91.610 185.405 92.015 185.575 ;
        RECT 90.735 184.725 90.975 185.125 ;
        RECT 91.455 184.955 91.675 185.235 ;
        RECT 91.145 184.785 91.675 184.955 ;
        RECT 91.145 184.555 91.315 184.785 ;
        RECT 91.845 184.625 92.015 185.405 ;
        RECT 92.185 184.795 92.535 185.415 ;
        RECT 92.705 184.795 92.915 185.585 ;
        RECT 93.105 185.615 94.605 185.785 ;
        RECT 93.105 184.925 93.275 185.615 ;
        RECT 94.965 185.445 95.135 186.225 ;
        RECT 95.940 186.095 96.110 186.225 ;
        RECT 93.445 185.275 95.135 185.445 ;
        RECT 95.305 185.665 95.770 186.055 ;
        RECT 95.940 185.925 96.335 186.095 ;
        RECT 93.445 185.095 93.615 185.275 ;
        RECT 90.245 184.385 91.315 184.555 ;
        RECT 91.485 184.175 91.675 184.615 ;
        RECT 91.845 184.345 92.795 184.625 ;
        RECT 93.105 184.535 93.365 184.925 ;
        RECT 93.785 184.855 94.575 185.105 ;
        RECT 93.015 184.365 93.365 184.535 ;
        RECT 93.575 184.175 93.905 184.635 ;
        RECT 94.780 184.565 94.950 185.275 ;
        RECT 95.305 185.075 95.475 185.665 ;
        RECT 95.120 184.855 95.475 185.075 ;
        RECT 95.645 184.855 95.995 185.475 ;
        RECT 96.165 184.565 96.335 185.925 ;
        RECT 96.700 185.755 97.025 186.540 ;
        RECT 96.505 184.705 96.965 185.755 ;
        RECT 94.780 184.395 95.635 184.565 ;
        RECT 95.840 184.395 96.335 184.565 ;
        RECT 96.505 184.175 96.835 184.535 ;
        RECT 97.195 184.435 97.365 186.555 ;
        RECT 97.535 186.225 97.865 186.725 ;
        RECT 98.035 186.055 98.290 186.555 ;
        RECT 97.540 185.885 98.290 186.055 ;
        RECT 97.540 184.895 97.770 185.885 ;
        RECT 97.940 185.065 98.290 185.715 ;
        RECT 98.465 185.650 98.735 186.555 ;
        RECT 98.905 185.965 99.235 186.725 ;
        RECT 99.415 185.795 99.585 186.555 ;
        RECT 97.540 184.725 98.290 184.895 ;
        RECT 97.535 184.175 97.865 184.555 ;
        RECT 98.035 184.435 98.290 184.725 ;
        RECT 98.465 184.850 98.635 185.650 ;
        RECT 98.920 185.625 99.585 185.795 ;
        RECT 100.395 185.795 100.565 186.555 ;
        RECT 100.745 185.965 101.075 186.725 ;
        RECT 100.395 185.625 101.060 185.795 ;
        RECT 101.245 185.650 101.515 186.555 ;
        RECT 98.920 185.480 99.090 185.625 ;
        RECT 98.805 185.150 99.090 185.480 ;
        RECT 100.890 185.480 101.060 185.625 ;
        RECT 98.920 184.895 99.090 185.150 ;
        RECT 99.325 185.075 99.655 185.445 ;
        RECT 100.325 185.075 100.655 185.445 ;
        RECT 100.890 185.150 101.175 185.480 ;
        RECT 100.890 184.895 101.060 185.150 ;
        RECT 98.465 184.345 98.725 184.850 ;
        RECT 98.920 184.725 99.585 184.895 ;
        RECT 98.905 184.175 99.235 184.555 ;
        RECT 99.415 184.345 99.585 184.725 ;
        RECT 100.395 184.725 101.060 184.895 ;
        RECT 101.345 184.850 101.515 185.650 ;
        RECT 101.685 185.560 101.975 186.725 ;
        RECT 102.150 185.585 102.485 186.555 ;
        RECT 102.655 185.585 102.825 186.725 ;
        RECT 102.995 186.385 105.025 186.555 ;
        RECT 102.150 184.915 102.320 185.585 ;
        RECT 102.995 185.415 103.165 186.385 ;
        RECT 102.490 185.085 102.745 185.415 ;
        RECT 102.970 185.085 103.165 185.415 ;
        RECT 103.335 186.045 104.460 186.215 ;
        RECT 102.575 184.915 102.745 185.085 ;
        RECT 103.335 184.915 103.505 186.045 ;
        RECT 100.395 184.345 100.565 184.725 ;
        RECT 100.745 184.175 101.075 184.555 ;
        RECT 101.255 184.345 101.515 184.850 ;
        RECT 101.685 184.175 101.975 184.900 ;
        RECT 102.150 184.345 102.405 184.915 ;
        RECT 102.575 184.745 103.505 184.915 ;
        RECT 103.675 185.705 104.685 185.875 ;
        RECT 103.675 184.905 103.845 185.705 ;
        RECT 104.050 185.365 104.325 185.505 ;
        RECT 104.045 185.195 104.325 185.365 ;
        RECT 103.330 184.710 103.505 184.745 ;
        RECT 102.575 184.175 102.905 184.575 ;
        RECT 103.330 184.345 103.860 184.710 ;
        RECT 104.050 184.345 104.325 185.195 ;
        RECT 104.495 184.345 104.685 185.705 ;
        RECT 104.855 185.720 105.025 186.385 ;
        RECT 105.195 185.965 105.365 186.725 ;
        RECT 105.600 185.965 106.115 186.375 ;
        RECT 104.855 185.530 105.605 185.720 ;
        RECT 105.775 185.155 106.115 185.965 ;
        RECT 104.885 184.985 106.115 185.155 ;
        RECT 106.285 185.585 106.670 186.555 ;
        RECT 106.840 186.265 107.165 186.725 ;
        RECT 107.685 186.095 107.965 186.555 ;
        RECT 106.840 185.875 107.965 186.095 ;
        RECT 104.865 184.175 105.375 184.710 ;
        RECT 105.595 184.380 105.840 184.985 ;
        RECT 106.285 184.915 106.565 185.585 ;
        RECT 106.840 185.415 107.290 185.875 ;
        RECT 108.155 185.705 108.555 186.555 ;
        RECT 108.955 186.265 109.225 186.725 ;
        RECT 109.395 186.095 109.680 186.555 ;
        RECT 106.735 185.085 107.290 185.415 ;
        RECT 107.460 185.145 108.555 185.705 ;
        RECT 106.840 184.975 107.290 185.085 ;
        RECT 106.285 184.345 106.670 184.915 ;
        RECT 106.840 184.805 107.965 184.975 ;
        RECT 106.840 184.175 107.165 184.635 ;
        RECT 107.685 184.345 107.965 184.805 ;
        RECT 108.155 184.345 108.555 185.145 ;
        RECT 108.725 185.875 109.680 186.095 ;
        RECT 108.725 184.975 108.935 185.875 ;
        RECT 109.105 185.145 109.795 185.705 ;
        RECT 109.965 185.585 110.305 186.555 ;
        RECT 110.475 185.585 110.645 186.725 ;
        RECT 110.915 185.925 111.165 186.725 ;
        RECT 111.810 185.755 112.140 186.555 ;
        RECT 112.440 185.925 112.770 186.725 ;
        RECT 112.940 185.755 113.270 186.555 ;
        RECT 110.835 185.585 113.270 185.755 ;
        RECT 114.105 185.965 114.620 186.375 ;
        RECT 114.855 185.965 115.025 186.725 ;
        RECT 115.195 186.385 117.225 186.555 ;
        RECT 109.965 184.975 110.140 185.585 ;
        RECT 110.835 185.335 111.005 185.585 ;
        RECT 110.310 185.165 111.005 185.335 ;
        RECT 111.180 185.165 111.600 185.365 ;
        RECT 111.770 185.165 112.100 185.365 ;
        RECT 112.270 185.165 112.600 185.365 ;
        RECT 108.725 184.805 109.680 184.975 ;
        RECT 108.955 184.175 109.225 184.635 ;
        RECT 109.395 184.345 109.680 184.805 ;
        RECT 109.965 184.345 110.305 184.975 ;
        RECT 110.475 184.175 110.725 184.975 ;
        RECT 110.915 184.825 112.140 184.995 ;
        RECT 110.915 184.345 111.245 184.825 ;
        RECT 111.415 184.175 111.640 184.635 ;
        RECT 111.810 184.345 112.140 184.825 ;
        RECT 112.770 184.955 112.940 185.585 ;
        RECT 113.125 185.165 113.475 185.415 ;
        RECT 114.105 185.155 114.445 185.965 ;
        RECT 115.195 185.720 115.365 186.385 ;
        RECT 115.760 186.045 116.885 186.215 ;
        RECT 114.615 185.530 115.365 185.720 ;
        RECT 115.535 185.705 116.545 185.875 ;
        RECT 114.105 184.985 115.335 185.155 ;
        RECT 112.770 184.345 113.270 184.955 ;
        RECT 114.380 184.380 114.625 184.985 ;
        RECT 114.845 184.175 115.355 184.710 ;
        RECT 115.535 184.345 115.725 185.705 ;
        RECT 115.895 185.365 116.170 185.505 ;
        RECT 115.895 185.195 116.175 185.365 ;
        RECT 115.895 184.345 116.170 185.195 ;
        RECT 116.375 184.905 116.545 185.705 ;
        RECT 116.715 184.915 116.885 186.045 ;
        RECT 117.055 185.415 117.225 186.385 ;
        RECT 117.395 185.585 117.565 186.725 ;
        RECT 117.735 185.585 118.070 186.555 ;
        RECT 117.055 185.085 117.250 185.415 ;
        RECT 117.475 185.085 117.730 185.415 ;
        RECT 117.475 184.915 117.645 185.085 ;
        RECT 117.900 184.915 118.070 185.585 ;
        RECT 116.715 184.745 117.645 184.915 ;
        RECT 116.715 184.710 116.890 184.745 ;
        RECT 116.360 184.345 116.890 184.710 ;
        RECT 117.315 184.175 117.645 184.575 ;
        RECT 117.815 184.345 118.070 184.915 ;
        RECT 118.245 185.585 118.630 186.555 ;
        RECT 118.800 186.265 119.125 186.725 ;
        RECT 119.645 186.095 119.925 186.555 ;
        RECT 118.800 185.875 119.925 186.095 ;
        RECT 118.245 184.915 118.525 185.585 ;
        RECT 118.800 185.415 119.250 185.875 ;
        RECT 120.115 185.705 120.515 186.555 ;
        RECT 120.915 186.265 121.185 186.725 ;
        RECT 121.355 186.095 121.640 186.555 ;
        RECT 118.695 185.085 119.250 185.415 ;
        RECT 119.420 185.145 120.515 185.705 ;
        RECT 118.800 184.975 119.250 185.085 ;
        RECT 118.245 184.345 118.630 184.915 ;
        RECT 118.800 184.805 119.925 184.975 ;
        RECT 118.800 184.175 119.125 184.635 ;
        RECT 119.645 184.345 119.925 184.805 ;
        RECT 120.115 184.345 120.515 185.145 ;
        RECT 120.685 185.875 121.640 186.095 ;
        RECT 120.685 184.975 120.895 185.875 ;
        RECT 122.015 185.795 122.185 186.555 ;
        RECT 122.365 185.965 122.695 186.725 ;
        RECT 121.065 185.145 121.755 185.705 ;
        RECT 122.015 185.625 122.680 185.795 ;
        RECT 122.865 185.650 123.135 186.555 ;
        RECT 122.510 185.480 122.680 185.625 ;
        RECT 121.945 185.075 122.275 185.445 ;
        RECT 122.510 185.150 122.795 185.480 ;
        RECT 120.685 184.805 121.640 184.975 ;
        RECT 122.510 184.895 122.680 185.150 ;
        RECT 120.915 184.175 121.185 184.635 ;
        RECT 121.355 184.345 121.640 184.805 ;
        RECT 122.015 184.725 122.680 184.895 ;
        RECT 122.965 184.850 123.135 185.650 ;
        RECT 123.395 185.795 123.565 186.555 ;
        RECT 123.745 185.965 124.075 186.725 ;
        RECT 123.395 185.625 124.060 185.795 ;
        RECT 124.245 185.650 124.515 186.555 ;
        RECT 123.890 185.480 124.060 185.625 ;
        RECT 123.325 185.075 123.655 185.445 ;
        RECT 123.890 185.150 124.175 185.480 ;
        RECT 123.890 184.895 124.060 185.150 ;
        RECT 122.015 184.345 122.185 184.725 ;
        RECT 122.365 184.175 122.695 184.555 ;
        RECT 122.875 184.345 123.135 184.850 ;
        RECT 123.395 184.725 124.060 184.895 ;
        RECT 124.345 184.850 124.515 185.650 ;
        RECT 124.685 185.635 126.355 186.725 ;
        RECT 126.525 185.635 127.735 186.725 ;
        RECT 124.685 185.115 125.435 185.635 ;
        RECT 125.605 184.945 126.355 185.465 ;
        RECT 126.525 185.095 127.045 185.635 ;
        RECT 123.395 184.345 123.565 184.725 ;
        RECT 123.745 184.175 124.075 184.555 ;
        RECT 124.255 184.345 124.515 184.850 ;
        RECT 124.685 184.175 126.355 184.945 ;
        RECT 127.215 184.925 127.735 185.465 ;
        RECT 126.525 184.175 127.735 184.925 ;
        RECT 29.840 184.005 127.820 184.175 ;
        RECT 29.925 183.255 31.135 184.005 ;
        RECT 29.925 182.715 30.445 183.255 ;
        RECT 32.285 183.185 32.495 184.005 ;
        RECT 32.665 183.205 32.995 183.835 ;
        RECT 30.615 182.545 31.135 183.085 ;
        RECT 32.665 182.605 32.915 183.205 ;
        RECT 33.165 183.185 33.395 184.005 ;
        RECT 33.720 183.375 34.005 183.835 ;
        RECT 34.175 183.545 34.445 184.005 ;
        RECT 33.720 183.205 34.675 183.375 ;
        RECT 33.085 182.765 33.415 183.015 ;
        RECT 29.925 181.455 31.135 182.545 ;
        RECT 32.285 181.455 32.495 182.595 ;
        RECT 32.665 181.625 32.995 182.605 ;
        RECT 33.165 181.455 33.395 182.595 ;
        RECT 33.605 182.475 34.295 183.035 ;
        RECT 34.465 182.305 34.675 183.205 ;
        RECT 33.720 182.085 34.675 182.305 ;
        RECT 34.845 183.035 35.245 183.835 ;
        RECT 35.435 183.375 35.715 183.835 ;
        RECT 36.235 183.545 36.560 184.005 ;
        RECT 35.435 183.205 36.560 183.375 ;
        RECT 36.730 183.265 37.115 183.835 ;
        RECT 37.285 183.280 37.575 184.005 ;
        RECT 38.755 183.455 38.925 183.835 ;
        RECT 39.105 183.625 39.435 184.005 ;
        RECT 38.755 183.285 39.420 183.455 ;
        RECT 39.615 183.330 39.875 183.835 ;
        RECT 36.110 183.095 36.560 183.205 ;
        RECT 34.845 182.475 35.940 183.035 ;
        RECT 36.110 182.765 36.665 183.095 ;
        RECT 33.720 181.625 34.005 182.085 ;
        RECT 34.175 181.455 34.445 181.915 ;
        RECT 34.845 181.625 35.245 182.475 ;
        RECT 36.110 182.305 36.560 182.765 ;
        RECT 36.835 182.595 37.115 183.265 ;
        RECT 38.685 182.735 39.015 183.105 ;
        RECT 39.250 183.030 39.420 183.285 ;
        RECT 39.250 182.700 39.535 183.030 ;
        RECT 35.435 182.085 36.560 182.305 ;
        RECT 35.435 181.625 35.715 182.085 ;
        RECT 36.235 181.455 36.560 181.915 ;
        RECT 36.730 181.625 37.115 182.595 ;
        RECT 37.285 181.455 37.575 182.620 ;
        RECT 39.250 182.555 39.420 182.700 ;
        RECT 38.755 182.385 39.420 182.555 ;
        RECT 39.705 182.530 39.875 183.330 ;
        RECT 38.755 181.625 38.925 182.385 ;
        RECT 39.105 181.455 39.435 182.215 ;
        RECT 39.605 181.625 39.875 182.530 ;
        RECT 40.050 183.265 40.305 183.835 ;
        RECT 40.475 183.605 40.805 184.005 ;
        RECT 41.230 183.470 41.760 183.835 ;
        RECT 41.230 183.435 41.405 183.470 ;
        RECT 40.475 183.265 41.405 183.435 ;
        RECT 40.050 182.595 40.220 183.265 ;
        RECT 40.475 183.095 40.645 183.265 ;
        RECT 40.390 182.765 40.645 183.095 ;
        RECT 40.870 182.765 41.065 183.095 ;
        RECT 40.050 181.625 40.385 182.595 ;
        RECT 40.555 181.455 40.725 182.595 ;
        RECT 40.895 181.795 41.065 182.765 ;
        RECT 41.235 182.135 41.405 183.265 ;
        RECT 41.575 182.475 41.745 183.275 ;
        RECT 41.950 182.985 42.225 183.835 ;
        RECT 41.945 182.815 42.225 182.985 ;
        RECT 41.950 182.675 42.225 182.815 ;
        RECT 42.395 182.475 42.585 183.835 ;
        RECT 42.765 183.470 43.275 184.005 ;
        RECT 43.495 183.195 43.740 183.800 ;
        RECT 44.190 183.295 44.445 183.825 ;
        RECT 44.615 183.545 44.920 184.005 ;
        RECT 45.165 183.625 46.235 183.795 ;
        RECT 42.785 183.025 44.015 183.195 ;
        RECT 41.575 182.305 42.585 182.475 ;
        RECT 42.755 182.460 43.505 182.650 ;
        RECT 41.235 181.965 42.360 182.135 ;
        RECT 42.755 181.795 42.925 182.460 ;
        RECT 43.675 182.215 44.015 183.025 ;
        RECT 40.895 181.625 42.925 181.795 ;
        RECT 43.095 181.455 43.265 182.215 ;
        RECT 43.500 181.805 44.015 182.215 ;
        RECT 44.190 182.645 44.400 183.295 ;
        RECT 45.165 183.270 45.485 183.625 ;
        RECT 45.160 183.095 45.485 183.270 ;
        RECT 44.570 182.795 45.485 183.095 ;
        RECT 45.655 183.055 45.895 183.455 ;
        RECT 46.065 183.395 46.235 183.625 ;
        RECT 46.405 183.565 46.595 184.005 ;
        RECT 46.765 183.555 47.715 183.835 ;
        RECT 47.935 183.645 48.285 183.815 ;
        RECT 46.065 183.225 46.595 183.395 ;
        RECT 44.570 182.765 45.310 182.795 ;
        RECT 44.190 181.765 44.445 182.645 ;
        RECT 44.615 181.455 44.920 182.595 ;
        RECT 45.140 182.175 45.310 182.765 ;
        RECT 45.655 182.685 46.195 183.055 ;
        RECT 46.375 182.945 46.595 183.225 ;
        RECT 46.765 182.775 46.935 183.555 ;
        RECT 46.530 182.605 46.935 182.775 ;
        RECT 47.105 182.765 47.455 183.385 ;
        RECT 46.530 182.515 46.700 182.605 ;
        RECT 47.625 182.595 47.835 183.385 ;
        RECT 45.480 182.345 46.700 182.515 ;
        RECT 47.160 182.435 47.835 182.595 ;
        RECT 45.140 182.005 45.940 182.175 ;
        RECT 45.260 181.455 45.590 181.835 ;
        RECT 45.770 181.715 45.940 182.005 ;
        RECT 46.530 181.965 46.700 182.345 ;
        RECT 46.870 182.425 47.835 182.435 ;
        RECT 48.025 183.255 48.285 183.645 ;
        RECT 48.495 183.545 48.825 184.005 ;
        RECT 49.700 183.615 50.555 183.785 ;
        RECT 50.760 183.615 51.255 183.785 ;
        RECT 51.425 183.645 51.755 184.005 ;
        RECT 48.025 182.565 48.195 183.255 ;
        RECT 48.365 182.905 48.535 183.085 ;
        RECT 48.705 183.075 49.495 183.325 ;
        RECT 49.700 182.905 49.870 183.615 ;
        RECT 50.040 183.105 50.395 183.325 ;
        RECT 48.365 182.735 50.055 182.905 ;
        RECT 46.870 182.135 47.330 182.425 ;
        RECT 48.025 182.395 49.525 182.565 ;
        RECT 48.025 182.255 48.195 182.395 ;
        RECT 47.635 182.085 48.195 182.255 ;
        RECT 46.110 181.455 46.360 181.915 ;
        RECT 46.530 181.625 47.400 181.965 ;
        RECT 47.635 181.625 47.805 182.085 ;
        RECT 48.640 182.055 49.715 182.225 ;
        RECT 47.975 181.455 48.345 181.915 ;
        RECT 48.640 181.715 48.810 182.055 ;
        RECT 48.980 181.455 49.310 181.885 ;
        RECT 49.545 181.715 49.715 182.055 ;
        RECT 49.885 181.955 50.055 182.735 ;
        RECT 50.225 182.515 50.395 183.105 ;
        RECT 50.565 182.705 50.915 183.325 ;
        RECT 50.225 182.125 50.690 182.515 ;
        RECT 51.085 182.255 51.255 183.615 ;
        RECT 51.425 182.425 51.885 183.475 ;
        RECT 50.860 182.085 51.255 182.255 ;
        RECT 50.860 181.955 51.030 182.085 ;
        RECT 49.885 181.625 50.565 181.955 ;
        RECT 50.780 181.625 51.030 181.955 ;
        RECT 51.200 181.455 51.450 181.915 ;
        RECT 51.620 181.640 51.945 182.425 ;
        RECT 52.115 181.625 52.285 183.745 ;
        RECT 52.455 183.625 52.785 184.005 ;
        RECT 52.955 183.455 53.210 183.745 ;
        RECT 52.460 183.285 53.210 183.455 ;
        RECT 52.460 182.295 52.690 183.285 ;
        RECT 53.390 183.265 53.645 183.835 ;
        RECT 53.815 183.605 54.145 184.005 ;
        RECT 54.570 183.470 55.100 183.835 ;
        RECT 55.290 183.665 55.565 183.835 ;
        RECT 55.285 183.495 55.565 183.665 ;
        RECT 54.570 183.435 54.745 183.470 ;
        RECT 53.815 183.265 54.745 183.435 ;
        RECT 52.860 182.465 53.210 183.115 ;
        RECT 53.390 182.595 53.560 183.265 ;
        RECT 53.815 183.095 53.985 183.265 ;
        RECT 53.730 182.765 53.985 183.095 ;
        RECT 54.210 182.765 54.405 183.095 ;
        RECT 52.460 182.125 53.210 182.295 ;
        RECT 52.455 181.455 52.785 181.955 ;
        RECT 52.955 181.625 53.210 182.125 ;
        RECT 53.390 181.625 53.725 182.595 ;
        RECT 53.895 181.455 54.065 182.595 ;
        RECT 54.235 181.795 54.405 182.765 ;
        RECT 54.575 182.135 54.745 183.265 ;
        RECT 54.915 182.475 55.085 183.275 ;
        RECT 55.290 182.675 55.565 183.495 ;
        RECT 55.735 182.475 55.925 183.835 ;
        RECT 56.105 183.470 56.615 184.005 ;
        RECT 56.835 183.195 57.080 183.800 ;
        RECT 57.615 183.455 57.785 183.835 ;
        RECT 57.965 183.625 58.295 184.005 ;
        RECT 57.615 183.285 58.280 183.455 ;
        RECT 58.475 183.330 58.735 183.835 ;
        RECT 56.125 183.025 57.355 183.195 ;
        RECT 54.915 182.305 55.925 182.475 ;
        RECT 56.095 182.460 56.845 182.650 ;
        RECT 54.575 181.965 55.700 182.135 ;
        RECT 56.095 181.795 56.265 182.460 ;
        RECT 57.015 182.215 57.355 183.025 ;
        RECT 57.545 182.735 57.875 183.105 ;
        RECT 58.110 183.030 58.280 183.285 ;
        RECT 58.110 182.700 58.395 183.030 ;
        RECT 58.110 182.555 58.280 182.700 ;
        RECT 54.235 181.625 56.265 181.795 ;
        RECT 56.435 181.455 56.605 182.215 ;
        RECT 56.840 181.805 57.355 182.215 ;
        RECT 57.615 182.385 58.280 182.555 ;
        RECT 58.565 182.530 58.735 183.330 ;
        RECT 59.570 183.225 60.070 183.835 ;
        RECT 59.365 182.765 59.715 183.015 ;
        RECT 59.900 182.595 60.070 183.225 ;
        RECT 60.700 183.355 61.030 183.835 ;
        RECT 61.200 183.545 61.425 184.005 ;
        RECT 61.595 183.355 61.925 183.835 ;
        RECT 60.700 183.185 61.925 183.355 ;
        RECT 62.115 183.205 62.365 184.005 ;
        RECT 62.535 183.205 62.875 183.835 ;
        RECT 63.045 183.280 63.335 184.005 ;
        RECT 60.240 182.815 60.570 183.015 ;
        RECT 60.740 182.815 61.070 183.015 ;
        RECT 61.240 182.815 61.660 183.015 ;
        RECT 61.835 182.845 62.530 183.015 ;
        RECT 61.835 182.595 62.005 182.845 ;
        RECT 62.700 182.595 62.875 183.205 ;
        RECT 64.240 183.195 64.485 183.800 ;
        RECT 64.705 183.470 65.215 184.005 ;
        RECT 63.965 183.025 65.195 183.195 ;
        RECT 57.615 181.625 57.785 182.385 ;
        RECT 57.965 181.455 58.295 182.215 ;
        RECT 58.465 181.625 58.735 182.530 ;
        RECT 59.570 182.425 62.005 182.595 ;
        RECT 59.570 181.625 59.900 182.425 ;
        RECT 60.070 181.455 60.400 182.255 ;
        RECT 60.700 181.625 61.030 182.425 ;
        RECT 61.675 181.455 61.925 182.255 ;
        RECT 62.195 181.455 62.365 182.595 ;
        RECT 62.535 181.625 62.875 182.595 ;
        RECT 63.045 181.455 63.335 182.620 ;
        RECT 63.965 182.215 64.305 183.025 ;
        RECT 64.475 182.460 65.225 182.650 ;
        RECT 63.965 181.805 64.480 182.215 ;
        RECT 64.715 181.455 64.885 182.215 ;
        RECT 65.055 181.795 65.225 182.460 ;
        RECT 65.395 182.475 65.585 183.835 ;
        RECT 65.755 183.665 66.030 183.835 ;
        RECT 65.755 183.495 66.035 183.665 ;
        RECT 65.755 182.675 66.030 183.495 ;
        RECT 66.220 183.470 66.750 183.835 ;
        RECT 67.175 183.605 67.505 184.005 ;
        RECT 66.575 183.435 66.750 183.470 ;
        RECT 66.235 182.475 66.405 183.275 ;
        RECT 65.395 182.305 66.405 182.475 ;
        RECT 66.575 183.265 67.505 183.435 ;
        RECT 67.675 183.265 67.930 183.835 ;
        RECT 66.575 182.135 66.745 183.265 ;
        RECT 67.335 183.095 67.505 183.265 ;
        RECT 65.620 181.965 66.745 182.135 ;
        RECT 66.915 182.765 67.110 183.095 ;
        RECT 67.335 182.765 67.590 183.095 ;
        RECT 66.915 181.795 67.085 182.765 ;
        RECT 67.760 182.595 67.930 183.265 ;
        RECT 65.055 181.625 67.085 181.795 ;
        RECT 67.255 181.455 67.425 182.595 ;
        RECT 67.595 181.625 67.930 182.595 ;
        RECT 68.110 183.295 68.365 183.825 ;
        RECT 68.535 183.545 68.840 184.005 ;
        RECT 69.085 183.625 70.155 183.795 ;
        RECT 68.110 182.645 68.320 183.295 ;
        RECT 69.085 183.270 69.405 183.625 ;
        RECT 69.080 183.095 69.405 183.270 ;
        RECT 68.490 182.795 69.405 183.095 ;
        RECT 69.575 183.055 69.815 183.455 ;
        RECT 69.985 183.395 70.155 183.625 ;
        RECT 70.325 183.565 70.515 184.005 ;
        RECT 70.685 183.555 71.635 183.835 ;
        RECT 71.855 183.645 72.205 183.815 ;
        RECT 69.985 183.225 70.515 183.395 ;
        RECT 68.490 182.765 69.230 182.795 ;
        RECT 68.110 181.765 68.365 182.645 ;
        RECT 68.535 181.455 68.840 182.595 ;
        RECT 69.060 182.175 69.230 182.765 ;
        RECT 69.575 182.685 70.115 183.055 ;
        RECT 70.295 182.945 70.515 183.225 ;
        RECT 70.685 182.775 70.855 183.555 ;
        RECT 70.450 182.605 70.855 182.775 ;
        RECT 71.025 182.765 71.375 183.385 ;
        RECT 70.450 182.515 70.620 182.605 ;
        RECT 71.545 182.595 71.755 183.385 ;
        RECT 69.400 182.345 70.620 182.515 ;
        RECT 71.080 182.435 71.755 182.595 ;
        RECT 69.060 182.005 69.860 182.175 ;
        RECT 69.180 181.455 69.510 181.835 ;
        RECT 69.690 181.715 69.860 182.005 ;
        RECT 70.450 181.965 70.620 182.345 ;
        RECT 70.790 182.425 71.755 182.435 ;
        RECT 71.945 183.255 72.205 183.645 ;
        RECT 72.415 183.545 72.745 184.005 ;
        RECT 73.620 183.615 74.475 183.785 ;
        RECT 74.680 183.615 75.175 183.785 ;
        RECT 75.345 183.645 75.675 184.005 ;
        RECT 71.945 182.565 72.115 183.255 ;
        RECT 72.285 182.905 72.455 183.085 ;
        RECT 72.625 183.075 73.415 183.325 ;
        RECT 73.620 182.905 73.790 183.615 ;
        RECT 73.960 183.105 74.315 183.325 ;
        RECT 72.285 182.735 73.975 182.905 ;
        RECT 70.790 182.135 71.250 182.425 ;
        RECT 71.945 182.395 73.445 182.565 ;
        RECT 71.945 182.255 72.115 182.395 ;
        RECT 71.555 182.085 72.115 182.255 ;
        RECT 70.030 181.455 70.280 181.915 ;
        RECT 70.450 181.625 71.320 181.965 ;
        RECT 71.555 181.625 71.725 182.085 ;
        RECT 72.560 182.055 73.635 182.225 ;
        RECT 71.895 181.455 72.265 181.915 ;
        RECT 72.560 181.715 72.730 182.055 ;
        RECT 72.900 181.455 73.230 181.885 ;
        RECT 73.465 181.715 73.635 182.055 ;
        RECT 73.805 181.955 73.975 182.735 ;
        RECT 74.145 182.515 74.315 183.105 ;
        RECT 74.485 182.705 74.835 183.325 ;
        RECT 74.145 182.125 74.610 182.515 ;
        RECT 75.005 182.255 75.175 183.615 ;
        RECT 75.345 182.425 75.805 183.475 ;
        RECT 74.780 182.085 75.175 182.255 ;
        RECT 74.780 181.955 74.950 182.085 ;
        RECT 73.805 181.625 74.485 181.955 ;
        RECT 74.700 181.625 74.950 181.955 ;
        RECT 75.120 181.455 75.370 181.915 ;
        RECT 75.540 181.640 75.865 182.425 ;
        RECT 76.035 181.625 76.205 183.745 ;
        RECT 76.375 183.625 76.705 184.005 ;
        RECT 76.875 183.455 77.130 183.745 ;
        RECT 76.380 183.285 77.130 183.455 ;
        RECT 77.315 183.475 77.645 183.835 ;
        RECT 77.815 183.645 78.145 184.005 ;
        RECT 78.345 183.475 78.675 183.835 ;
        RECT 76.380 182.295 76.610 183.285 ;
        RECT 77.315 183.265 78.675 183.475 ;
        RECT 79.185 183.245 79.895 183.835 ;
        RECT 76.780 182.465 77.130 183.115 ;
        RECT 77.305 182.765 77.615 183.095 ;
        RECT 77.825 182.765 78.200 183.095 ;
        RECT 78.520 182.765 79.015 183.095 ;
        RECT 76.380 182.125 77.130 182.295 ;
        RECT 76.375 181.455 76.705 181.955 ;
        RECT 76.875 181.625 77.130 182.125 ;
        RECT 77.315 181.455 77.645 182.515 ;
        RECT 77.825 181.795 77.995 182.765 ;
        RECT 78.165 182.275 78.495 182.495 ;
        RECT 78.690 182.475 79.015 182.765 ;
        RECT 79.190 182.475 79.520 183.015 ;
        RECT 79.690 182.275 79.895 183.245 ;
        RECT 78.165 182.045 79.895 182.275 ;
        RECT 78.165 181.645 78.495 182.045 ;
        RECT 78.665 181.455 78.995 181.815 ;
        RECT 79.195 181.625 79.895 182.045 ;
        RECT 80.065 183.205 80.405 183.835 ;
        RECT 80.575 183.205 80.825 184.005 ;
        RECT 81.015 183.355 81.345 183.835 ;
        RECT 81.515 183.545 81.740 184.005 ;
        RECT 81.910 183.355 82.240 183.835 ;
        RECT 80.065 182.595 80.240 183.205 ;
        RECT 81.015 183.185 82.240 183.355 ;
        RECT 82.870 183.225 83.370 183.835 ;
        RECT 80.410 182.845 81.105 183.015 ;
        RECT 80.935 182.595 81.105 182.845 ;
        RECT 81.280 182.815 81.700 183.015 ;
        RECT 81.870 182.815 82.200 183.015 ;
        RECT 82.370 182.815 82.700 183.015 ;
        RECT 82.870 182.595 83.040 183.225 ;
        RECT 83.745 183.205 84.085 183.835 ;
        RECT 84.255 183.205 84.505 184.005 ;
        RECT 84.695 183.355 85.025 183.835 ;
        RECT 85.195 183.545 85.420 184.005 ;
        RECT 85.590 183.355 85.920 183.835 ;
        RECT 83.225 182.765 83.575 183.015 ;
        RECT 83.745 182.595 83.920 183.205 ;
        RECT 84.695 183.185 85.920 183.355 ;
        RECT 86.550 183.225 87.050 183.835 ;
        RECT 84.090 182.845 84.785 183.015 ;
        RECT 84.615 182.595 84.785 182.845 ;
        RECT 84.960 182.815 85.380 183.015 ;
        RECT 85.550 182.815 85.880 183.015 ;
        RECT 86.050 182.815 86.380 183.015 ;
        RECT 86.550 182.595 86.720 183.225 ;
        RECT 87.465 183.185 87.695 184.005 ;
        RECT 87.865 183.205 88.195 183.835 ;
        RECT 86.905 182.765 87.255 183.015 ;
        RECT 87.445 182.765 87.775 183.015 ;
        RECT 87.945 182.605 88.195 183.205 ;
        RECT 88.365 183.185 88.575 184.005 ;
        RECT 88.805 183.280 89.095 184.005 ;
        RECT 89.375 183.525 89.545 184.005 ;
        RECT 89.715 183.355 90.045 183.830 ;
        RECT 90.215 183.525 90.385 184.005 ;
        RECT 90.555 183.355 90.885 183.830 ;
        RECT 91.055 183.525 91.225 184.005 ;
        RECT 91.395 183.355 91.725 183.830 ;
        RECT 91.895 183.525 92.065 184.005 ;
        RECT 92.235 183.355 92.565 183.830 ;
        RECT 92.735 183.525 92.905 184.005 ;
        RECT 93.075 183.355 93.405 183.830 ;
        RECT 93.575 183.525 93.745 184.005 ;
        RECT 93.995 183.830 94.165 183.835 ;
        RECT 93.915 183.355 94.245 183.830 ;
        RECT 94.415 183.525 94.585 184.005 ;
        RECT 94.835 183.830 95.005 183.835 ;
        RECT 94.755 183.355 95.085 183.830 ;
        RECT 95.255 183.525 95.425 184.005 ;
        RECT 95.675 183.830 95.925 183.835 ;
        RECT 95.595 183.355 95.925 183.830 ;
        RECT 96.095 183.525 96.265 184.005 ;
        RECT 96.435 183.355 96.765 183.830 ;
        RECT 96.935 183.525 97.105 184.005 ;
        RECT 97.275 183.355 97.605 183.830 ;
        RECT 97.775 183.525 97.945 184.005 ;
        RECT 98.115 183.355 98.445 183.830 ;
        RECT 98.615 183.525 98.785 184.005 ;
        RECT 98.955 183.355 99.285 183.830 ;
        RECT 99.455 183.525 99.625 184.005 ;
        RECT 99.795 183.355 100.125 183.830 ;
        RECT 89.265 183.185 95.925 183.355 ;
        RECT 96.095 183.185 98.445 183.355 ;
        RECT 98.615 183.185 100.125 183.355 ;
        RECT 100.305 183.265 100.690 183.835 ;
        RECT 100.860 183.545 101.185 184.005 ;
        RECT 101.705 183.375 101.985 183.835 ;
        RECT 89.265 182.645 89.540 183.185 ;
        RECT 96.095 183.015 96.270 183.185 ;
        RECT 98.615 183.015 98.785 183.185 ;
        RECT 89.710 182.815 96.270 183.015 ;
        RECT 96.475 182.815 98.785 183.015 ;
        RECT 98.955 182.815 100.130 183.015 ;
        RECT 96.095 182.645 96.270 182.815 ;
        RECT 98.615 182.645 98.785 182.815 ;
        RECT 80.065 181.625 80.405 182.595 ;
        RECT 80.575 181.455 80.745 182.595 ;
        RECT 80.935 182.425 83.370 182.595 ;
        RECT 81.015 181.455 81.265 182.255 ;
        RECT 81.910 181.625 82.240 182.425 ;
        RECT 82.540 181.455 82.870 182.255 ;
        RECT 83.040 181.625 83.370 182.425 ;
        RECT 83.745 181.625 84.085 182.595 ;
        RECT 84.255 181.455 84.425 182.595 ;
        RECT 84.615 182.425 87.050 182.595 ;
        RECT 84.695 181.455 84.945 182.255 ;
        RECT 85.590 181.625 85.920 182.425 ;
        RECT 86.220 181.455 86.550 182.255 ;
        RECT 86.720 181.625 87.050 182.425 ;
        RECT 87.465 181.455 87.695 182.595 ;
        RECT 87.865 181.625 88.195 182.605 ;
        RECT 88.365 181.455 88.575 182.595 ;
        RECT 88.805 181.455 89.095 182.620 ;
        RECT 89.265 182.475 95.925 182.645 ;
        RECT 96.095 182.475 98.445 182.645 ;
        RECT 98.615 182.475 100.125 182.645 ;
        RECT 89.375 181.455 89.545 182.255 ;
        RECT 89.715 181.625 90.045 182.475 ;
        RECT 90.215 181.455 90.385 182.255 ;
        RECT 90.555 181.625 90.885 182.475 ;
        RECT 91.055 181.455 91.225 182.255 ;
        RECT 91.395 181.625 91.725 182.475 ;
        RECT 91.895 181.455 92.065 182.255 ;
        RECT 92.235 181.625 92.565 182.475 ;
        RECT 92.735 181.455 92.905 182.255 ;
        RECT 93.075 181.625 93.405 182.475 ;
        RECT 93.575 181.455 93.745 182.255 ;
        RECT 93.915 181.625 94.245 182.475 ;
        RECT 94.415 181.455 94.585 182.255 ;
        RECT 94.755 181.625 95.085 182.475 ;
        RECT 95.255 181.455 95.425 182.255 ;
        RECT 95.595 181.625 95.925 182.475 ;
        RECT 96.095 181.455 96.265 182.255 ;
        RECT 96.435 181.625 96.765 182.475 ;
        RECT 96.935 181.455 97.105 182.255 ;
        RECT 97.275 181.625 97.605 182.475 ;
        RECT 97.775 181.455 97.945 182.255 ;
        RECT 98.115 181.625 98.445 182.475 ;
        RECT 98.615 181.455 98.785 182.305 ;
        RECT 98.955 181.625 99.285 182.475 ;
        RECT 99.455 181.455 99.625 182.305 ;
        RECT 99.795 181.625 100.125 182.475 ;
        RECT 100.305 182.595 100.585 183.265 ;
        RECT 100.860 183.205 101.985 183.375 ;
        RECT 100.860 183.095 101.310 183.205 ;
        RECT 100.755 182.765 101.310 183.095 ;
        RECT 102.175 183.035 102.575 183.835 ;
        RECT 102.975 183.545 103.245 184.005 ;
        RECT 103.415 183.375 103.700 183.835 ;
        RECT 100.305 181.625 100.690 182.595 ;
        RECT 100.860 182.305 101.310 182.765 ;
        RECT 101.480 182.475 102.575 183.035 ;
        RECT 100.860 182.085 101.985 182.305 ;
        RECT 100.860 181.455 101.185 181.915 ;
        RECT 101.705 181.625 101.985 182.085 ;
        RECT 102.175 181.625 102.575 182.475 ;
        RECT 102.745 183.205 103.700 183.375 ;
        RECT 103.985 183.205 104.325 183.835 ;
        RECT 104.495 183.205 104.745 184.005 ;
        RECT 104.935 183.355 105.265 183.835 ;
        RECT 105.435 183.545 105.660 184.005 ;
        RECT 105.830 183.355 106.160 183.835 ;
        RECT 102.745 182.305 102.955 183.205 ;
        RECT 103.125 182.475 103.815 183.035 ;
        RECT 103.985 182.595 104.160 183.205 ;
        RECT 104.935 183.185 106.160 183.355 ;
        RECT 106.790 183.225 107.290 183.835 ;
        RECT 104.330 182.845 105.025 183.015 ;
        RECT 104.855 182.595 105.025 182.845 ;
        RECT 105.200 182.815 105.620 183.015 ;
        RECT 105.790 182.815 106.120 183.015 ;
        RECT 106.290 182.815 106.620 183.015 ;
        RECT 106.790 182.595 106.960 183.225 ;
        RECT 107.665 183.205 108.005 183.835 ;
        RECT 108.175 183.205 108.425 184.005 ;
        RECT 108.615 183.355 108.945 183.835 ;
        RECT 109.115 183.545 109.340 184.005 ;
        RECT 109.510 183.355 109.840 183.835 ;
        RECT 107.145 182.765 107.495 183.015 ;
        RECT 107.665 182.595 107.840 183.205 ;
        RECT 108.615 183.185 109.840 183.355 ;
        RECT 110.470 183.225 110.970 183.835 ;
        RECT 108.010 182.845 108.705 183.015 ;
        RECT 108.535 182.595 108.705 182.845 ;
        RECT 108.880 182.815 109.300 183.015 ;
        RECT 109.470 182.815 109.800 183.015 ;
        RECT 109.970 182.815 110.300 183.015 ;
        RECT 110.470 182.595 110.640 183.225 ;
        RECT 111.845 183.185 112.075 184.005 ;
        RECT 112.245 183.205 112.575 183.835 ;
        RECT 110.825 182.765 111.175 183.015 ;
        RECT 111.825 182.765 112.155 183.015 ;
        RECT 112.325 182.605 112.575 183.205 ;
        RECT 112.745 183.185 112.955 184.005 ;
        RECT 113.225 183.185 113.455 184.005 ;
        RECT 113.625 183.205 113.955 183.835 ;
        RECT 113.205 182.765 113.535 183.015 ;
        RECT 113.705 182.605 113.955 183.205 ;
        RECT 114.125 183.185 114.335 184.005 ;
        RECT 114.565 183.280 114.855 184.005 ;
        RECT 115.025 183.205 115.365 183.835 ;
        RECT 115.535 183.205 115.785 184.005 ;
        RECT 115.975 183.355 116.305 183.835 ;
        RECT 116.475 183.545 116.700 184.005 ;
        RECT 116.870 183.355 117.200 183.835 ;
        RECT 102.745 182.085 103.700 182.305 ;
        RECT 102.975 181.455 103.245 181.915 ;
        RECT 103.415 181.625 103.700 182.085 ;
        RECT 103.985 181.625 104.325 182.595 ;
        RECT 104.495 181.455 104.665 182.595 ;
        RECT 104.855 182.425 107.290 182.595 ;
        RECT 104.935 181.455 105.185 182.255 ;
        RECT 105.830 181.625 106.160 182.425 ;
        RECT 106.460 181.455 106.790 182.255 ;
        RECT 106.960 181.625 107.290 182.425 ;
        RECT 107.665 181.625 108.005 182.595 ;
        RECT 108.175 181.455 108.345 182.595 ;
        RECT 108.535 182.425 110.970 182.595 ;
        RECT 108.615 181.455 108.865 182.255 ;
        RECT 109.510 181.625 109.840 182.425 ;
        RECT 110.140 181.455 110.470 182.255 ;
        RECT 110.640 181.625 110.970 182.425 ;
        RECT 111.845 181.455 112.075 182.595 ;
        RECT 112.245 181.625 112.575 182.605 ;
        RECT 112.745 181.455 112.955 182.595 ;
        RECT 113.225 181.455 113.455 182.595 ;
        RECT 113.625 181.625 113.955 182.605 ;
        RECT 114.125 181.455 114.335 182.595 ;
        RECT 114.565 181.455 114.855 182.620 ;
        RECT 115.025 182.595 115.200 183.205 ;
        RECT 115.975 183.185 117.200 183.355 ;
        RECT 117.830 183.225 118.330 183.835 ;
        RECT 118.820 183.375 119.105 183.835 ;
        RECT 119.275 183.545 119.545 184.005 ;
        RECT 115.370 182.845 116.065 183.015 ;
        RECT 115.895 182.595 116.065 182.845 ;
        RECT 116.240 182.815 116.660 183.015 ;
        RECT 116.830 182.815 117.160 183.015 ;
        RECT 117.330 182.815 117.660 183.015 ;
        RECT 117.830 182.595 118.000 183.225 ;
        RECT 118.820 183.205 119.775 183.375 ;
        RECT 118.185 182.765 118.535 183.015 ;
        RECT 115.025 181.625 115.365 182.595 ;
        RECT 115.535 181.455 115.705 182.595 ;
        RECT 115.895 182.425 118.330 182.595 ;
        RECT 118.705 182.475 119.395 183.035 ;
        RECT 115.975 181.455 116.225 182.255 ;
        RECT 116.870 181.625 117.200 182.425 ;
        RECT 117.500 181.455 117.830 182.255 ;
        RECT 118.000 181.625 118.330 182.425 ;
        RECT 119.565 182.305 119.775 183.205 ;
        RECT 118.820 182.085 119.775 182.305 ;
        RECT 119.945 183.035 120.345 183.835 ;
        RECT 120.535 183.375 120.815 183.835 ;
        RECT 121.335 183.545 121.660 184.005 ;
        RECT 120.535 183.205 121.660 183.375 ;
        RECT 121.830 183.265 122.215 183.835 ;
        RECT 122.475 183.455 122.645 183.835 ;
        RECT 122.825 183.625 123.155 184.005 ;
        RECT 122.475 183.285 123.140 183.455 ;
        RECT 123.335 183.330 123.595 183.835 ;
        RECT 121.210 183.095 121.660 183.205 ;
        RECT 119.945 182.475 121.040 183.035 ;
        RECT 121.210 182.765 121.765 183.095 ;
        RECT 118.820 181.625 119.105 182.085 ;
        RECT 119.275 181.455 119.545 181.915 ;
        RECT 119.945 181.625 120.345 182.475 ;
        RECT 121.210 182.305 121.660 182.765 ;
        RECT 121.935 182.595 122.215 183.265 ;
        RECT 122.405 182.735 122.735 183.105 ;
        RECT 122.970 183.030 123.140 183.285 ;
        RECT 120.535 182.085 121.660 182.305 ;
        RECT 120.535 181.625 120.815 182.085 ;
        RECT 121.335 181.455 121.660 181.915 ;
        RECT 121.830 181.625 122.215 182.595 ;
        RECT 122.970 182.700 123.255 183.030 ;
        RECT 122.970 182.555 123.140 182.700 ;
        RECT 122.475 182.385 123.140 182.555 ;
        RECT 123.425 182.530 123.595 183.330 ;
        RECT 123.765 183.235 126.355 184.005 ;
        RECT 126.525 183.255 127.735 184.005 ;
        RECT 122.475 181.625 122.645 182.385 ;
        RECT 122.825 181.455 123.155 182.215 ;
        RECT 123.325 181.625 123.595 182.530 ;
        RECT 123.765 182.545 124.975 183.065 ;
        RECT 125.145 182.715 126.355 183.235 ;
        RECT 126.525 182.545 127.045 183.085 ;
        RECT 127.215 182.715 127.735 183.255 ;
        RECT 123.765 181.455 126.355 182.545 ;
        RECT 126.525 181.455 127.735 182.545 ;
        RECT 29.840 181.285 127.820 181.455 ;
        RECT 29.925 180.195 31.135 181.285 ;
        RECT 29.925 179.485 30.445 180.025 ;
        RECT 30.615 179.655 31.135 180.195 ;
        RECT 31.765 180.145 32.105 181.115 ;
        RECT 32.275 180.145 32.445 181.285 ;
        RECT 32.715 180.485 32.965 181.285 ;
        RECT 33.610 180.315 33.940 181.115 ;
        RECT 34.240 180.485 34.570 181.285 ;
        RECT 34.740 180.315 35.070 181.115 ;
        RECT 32.635 180.145 35.070 180.315 ;
        RECT 35.650 180.315 35.980 181.115 ;
        RECT 36.150 180.485 36.480 181.285 ;
        RECT 36.780 180.315 37.110 181.115 ;
        RECT 37.755 180.485 38.005 181.285 ;
        RECT 35.650 180.145 38.085 180.315 ;
        RECT 38.275 180.145 38.445 181.285 ;
        RECT 38.615 180.145 38.955 181.115 ;
        RECT 31.765 179.535 31.940 180.145 ;
        RECT 32.635 179.895 32.805 180.145 ;
        RECT 32.110 179.725 32.805 179.895 ;
        RECT 32.980 179.725 33.400 179.925 ;
        RECT 33.570 179.725 33.900 179.925 ;
        RECT 34.070 179.725 34.400 179.925 ;
        RECT 29.925 178.735 31.135 179.485 ;
        RECT 31.765 178.905 32.105 179.535 ;
        RECT 32.275 178.735 32.525 179.535 ;
        RECT 32.715 179.385 33.940 179.555 ;
        RECT 32.715 178.905 33.045 179.385 ;
        RECT 33.215 178.735 33.440 179.195 ;
        RECT 33.610 178.905 33.940 179.385 ;
        RECT 34.570 179.515 34.740 180.145 ;
        RECT 34.925 179.725 35.275 179.975 ;
        RECT 35.445 179.725 35.795 179.975 ;
        RECT 35.980 179.515 36.150 180.145 ;
        RECT 36.320 179.725 36.650 179.925 ;
        RECT 36.820 179.725 37.150 179.925 ;
        RECT 37.320 179.725 37.740 179.925 ;
        RECT 37.915 179.895 38.085 180.145 ;
        RECT 37.915 179.725 38.610 179.895 ;
        RECT 38.780 179.585 38.955 180.145 ;
        RECT 34.570 178.905 35.070 179.515 ;
        RECT 35.650 178.905 36.150 179.515 ;
        RECT 36.780 179.385 38.005 179.555 ;
        RECT 38.725 179.535 38.955 179.585 ;
        RECT 36.780 178.905 37.110 179.385 ;
        RECT 37.280 178.735 37.505 179.195 ;
        RECT 37.675 178.905 38.005 179.385 ;
        RECT 38.195 178.735 38.445 179.535 ;
        RECT 38.615 178.905 38.955 179.535 ;
        RECT 39.125 180.145 39.465 181.115 ;
        RECT 39.635 180.145 39.805 181.285 ;
        RECT 40.075 180.485 40.325 181.285 ;
        RECT 40.970 180.315 41.300 181.115 ;
        RECT 41.600 180.485 41.930 181.285 ;
        RECT 42.100 180.315 42.430 181.115 ;
        RECT 42.920 180.655 43.205 181.115 ;
        RECT 43.375 180.825 43.645 181.285 ;
        RECT 42.920 180.435 43.875 180.655 ;
        RECT 39.995 180.145 42.430 180.315 ;
        RECT 39.125 179.535 39.300 180.145 ;
        RECT 39.995 179.895 40.165 180.145 ;
        RECT 39.470 179.725 40.165 179.895 ;
        RECT 40.340 179.725 40.760 179.925 ;
        RECT 40.930 179.725 41.260 179.925 ;
        RECT 41.430 179.725 41.760 179.925 ;
        RECT 39.125 178.905 39.465 179.535 ;
        RECT 39.635 178.735 39.885 179.535 ;
        RECT 40.075 179.385 41.300 179.555 ;
        RECT 40.075 178.905 40.405 179.385 ;
        RECT 40.575 178.735 40.800 179.195 ;
        RECT 40.970 178.905 41.300 179.385 ;
        RECT 41.930 179.515 42.100 180.145 ;
        RECT 42.285 179.725 42.635 179.975 ;
        RECT 42.805 179.705 43.495 180.265 ;
        RECT 43.665 179.535 43.875 180.435 ;
        RECT 41.930 178.905 42.430 179.515 ;
        RECT 42.920 179.365 43.875 179.535 ;
        RECT 44.045 180.265 44.445 181.115 ;
        RECT 44.635 180.655 44.915 181.115 ;
        RECT 45.435 180.825 45.760 181.285 ;
        RECT 44.635 180.435 45.760 180.655 ;
        RECT 44.045 179.705 45.140 180.265 ;
        RECT 45.310 179.975 45.760 180.435 ;
        RECT 45.930 180.145 46.315 181.115 ;
        RECT 46.690 180.315 47.020 181.115 ;
        RECT 47.190 180.485 47.520 181.285 ;
        RECT 47.820 180.315 48.150 181.115 ;
        RECT 48.795 180.485 49.045 181.285 ;
        RECT 46.690 180.145 49.125 180.315 ;
        RECT 49.315 180.145 49.485 181.285 ;
        RECT 49.655 180.145 49.995 181.115 ;
        RECT 42.920 178.905 43.205 179.365 ;
        RECT 43.375 178.735 43.645 179.195 ;
        RECT 44.045 178.905 44.445 179.705 ;
        RECT 45.310 179.645 45.865 179.975 ;
        RECT 45.310 179.535 45.760 179.645 ;
        RECT 44.635 179.365 45.760 179.535 ;
        RECT 46.035 179.475 46.315 180.145 ;
        RECT 46.485 179.725 46.835 179.975 ;
        RECT 47.020 179.515 47.190 180.145 ;
        RECT 47.360 179.725 47.690 179.925 ;
        RECT 47.860 179.725 48.190 179.925 ;
        RECT 48.360 179.725 48.780 179.925 ;
        RECT 48.955 179.895 49.125 180.145 ;
        RECT 48.955 179.725 49.650 179.895 ;
        RECT 44.635 178.905 44.915 179.365 ;
        RECT 45.435 178.735 45.760 179.195 ;
        RECT 45.930 178.905 46.315 179.475 ;
        RECT 46.690 178.905 47.190 179.515 ;
        RECT 47.820 179.385 49.045 179.555 ;
        RECT 49.820 179.535 49.995 180.145 ;
        RECT 50.165 180.120 50.455 181.285 ;
        RECT 50.830 180.315 51.160 181.115 ;
        RECT 51.330 180.485 51.660 181.285 ;
        RECT 51.960 180.315 52.290 181.115 ;
        RECT 52.935 180.485 53.185 181.285 ;
        RECT 50.830 180.145 53.265 180.315 ;
        RECT 53.455 180.145 53.625 181.285 ;
        RECT 53.795 180.145 54.135 181.115 ;
        RECT 50.625 179.725 50.975 179.975 ;
        RECT 47.820 178.905 48.150 179.385 ;
        RECT 48.320 178.735 48.545 179.195 ;
        RECT 48.715 178.905 49.045 179.385 ;
        RECT 49.235 178.735 49.485 179.535 ;
        RECT 49.655 178.905 49.995 179.535 ;
        RECT 51.160 179.515 51.330 180.145 ;
        RECT 51.500 179.725 51.830 179.925 ;
        RECT 52.000 179.725 52.330 179.925 ;
        RECT 52.500 179.725 52.920 179.925 ;
        RECT 53.095 179.895 53.265 180.145 ;
        RECT 53.095 179.725 53.790 179.895 ;
        RECT 50.165 178.735 50.455 179.460 ;
        RECT 50.830 178.905 51.330 179.515 ;
        RECT 51.960 179.385 53.185 179.555 ;
        RECT 53.960 179.535 54.135 180.145 ;
        RECT 51.960 178.905 52.290 179.385 ;
        RECT 52.460 178.735 52.685 179.195 ;
        RECT 52.855 178.905 53.185 179.385 ;
        RECT 53.375 178.735 53.625 179.535 ;
        RECT 53.795 178.905 54.135 179.535 ;
        RECT 54.305 180.145 54.645 181.115 ;
        RECT 54.815 180.145 54.985 181.285 ;
        RECT 55.255 180.485 55.505 181.285 ;
        RECT 56.150 180.315 56.480 181.115 ;
        RECT 56.780 180.485 57.110 181.285 ;
        RECT 57.280 180.315 57.610 181.115 ;
        RECT 55.175 180.145 57.610 180.315 ;
        RECT 57.985 180.145 58.370 181.115 ;
        RECT 58.540 180.825 58.865 181.285 ;
        RECT 59.385 180.655 59.665 181.115 ;
        RECT 58.540 180.435 59.665 180.655 ;
        RECT 54.305 179.535 54.480 180.145 ;
        RECT 55.175 179.895 55.345 180.145 ;
        RECT 54.650 179.725 55.345 179.895 ;
        RECT 55.520 179.725 55.940 179.925 ;
        RECT 56.110 179.725 56.440 179.925 ;
        RECT 56.610 179.725 56.940 179.925 ;
        RECT 54.305 178.905 54.645 179.535 ;
        RECT 54.815 178.735 55.065 179.535 ;
        RECT 55.255 179.385 56.480 179.555 ;
        RECT 55.255 178.905 55.585 179.385 ;
        RECT 55.755 178.735 55.980 179.195 ;
        RECT 56.150 178.905 56.480 179.385 ;
        RECT 57.110 179.515 57.280 180.145 ;
        RECT 57.465 179.725 57.815 179.975 ;
        RECT 57.110 178.905 57.610 179.515 ;
        RECT 57.985 179.475 58.265 180.145 ;
        RECT 58.540 179.975 58.990 180.435 ;
        RECT 59.855 180.265 60.255 181.115 ;
        RECT 60.655 180.825 60.925 181.285 ;
        RECT 61.095 180.655 61.380 181.115 ;
        RECT 58.435 179.645 58.990 179.975 ;
        RECT 59.160 179.705 60.255 180.265 ;
        RECT 58.540 179.535 58.990 179.645 ;
        RECT 57.985 178.905 58.370 179.475 ;
        RECT 58.540 179.365 59.665 179.535 ;
        RECT 58.540 178.735 58.865 179.195 ;
        RECT 59.385 178.905 59.665 179.365 ;
        RECT 59.855 178.905 60.255 179.705 ;
        RECT 60.425 180.435 61.380 180.655 ;
        RECT 61.780 180.655 62.065 181.115 ;
        RECT 62.235 180.825 62.505 181.285 ;
        RECT 61.780 180.435 62.735 180.655 ;
        RECT 60.425 179.535 60.635 180.435 ;
        RECT 60.805 179.705 61.495 180.265 ;
        RECT 61.665 179.705 62.355 180.265 ;
        RECT 62.525 179.535 62.735 180.435 ;
        RECT 60.425 179.365 61.380 179.535 ;
        RECT 60.655 178.735 60.925 179.195 ;
        RECT 61.095 178.905 61.380 179.365 ;
        RECT 61.780 179.365 62.735 179.535 ;
        RECT 62.905 180.265 63.305 181.115 ;
        RECT 63.495 180.655 63.775 181.115 ;
        RECT 64.295 180.825 64.620 181.285 ;
        RECT 63.495 180.435 64.620 180.655 ;
        RECT 62.905 179.705 64.000 180.265 ;
        RECT 64.170 179.975 64.620 180.435 ;
        RECT 64.790 180.145 65.175 181.115 ;
        RECT 61.780 178.905 62.065 179.365 ;
        RECT 62.235 178.735 62.505 179.195 ;
        RECT 62.905 178.905 63.305 179.705 ;
        RECT 64.170 179.645 64.725 179.975 ;
        RECT 64.170 179.535 64.620 179.645 ;
        RECT 63.495 179.365 64.620 179.535 ;
        RECT 64.895 179.475 65.175 180.145 ;
        RECT 65.345 180.195 67.015 181.285 ;
        RECT 65.345 179.675 66.095 180.195 ;
        RECT 67.185 180.145 67.525 181.115 ;
        RECT 67.695 180.145 67.865 181.285 ;
        RECT 68.135 180.485 68.385 181.285 ;
        RECT 69.030 180.315 69.360 181.115 ;
        RECT 69.660 180.485 69.990 181.285 ;
        RECT 70.160 180.315 70.490 181.115 ;
        RECT 68.055 180.145 70.490 180.315 ;
        RECT 70.955 180.355 71.125 181.115 ;
        RECT 71.305 180.525 71.635 181.285 ;
        RECT 70.955 180.185 71.620 180.355 ;
        RECT 71.805 180.210 72.075 181.115 ;
        RECT 66.265 179.505 67.015 180.025 ;
        RECT 63.495 178.905 63.775 179.365 ;
        RECT 64.295 178.735 64.620 179.195 ;
        RECT 64.790 178.905 65.175 179.475 ;
        RECT 65.345 178.735 67.015 179.505 ;
        RECT 67.185 179.535 67.360 180.145 ;
        RECT 68.055 179.895 68.225 180.145 ;
        RECT 67.530 179.725 68.225 179.895 ;
        RECT 68.400 179.725 68.820 179.925 ;
        RECT 68.990 179.725 69.320 179.925 ;
        RECT 69.490 179.725 69.820 179.925 ;
        RECT 67.185 178.905 67.525 179.535 ;
        RECT 67.695 178.735 67.945 179.535 ;
        RECT 68.135 179.385 69.360 179.555 ;
        RECT 68.135 178.905 68.465 179.385 ;
        RECT 68.635 178.735 68.860 179.195 ;
        RECT 69.030 178.905 69.360 179.385 ;
        RECT 69.990 179.515 70.160 180.145 ;
        RECT 71.450 180.040 71.620 180.185 ;
        RECT 70.345 179.725 70.695 179.975 ;
        RECT 70.885 179.635 71.215 180.005 ;
        RECT 71.450 179.710 71.735 180.040 ;
        RECT 69.990 178.905 70.490 179.515 ;
        RECT 71.450 179.455 71.620 179.710 ;
        RECT 70.955 179.285 71.620 179.455 ;
        RECT 71.905 179.410 72.075 180.210 ;
        RECT 72.250 180.135 72.510 181.285 ;
        RECT 72.685 180.210 72.940 181.115 ;
        RECT 73.110 180.525 73.440 181.285 ;
        RECT 73.655 180.355 73.825 181.115 ;
        RECT 70.955 178.905 71.125 179.285 ;
        RECT 71.305 178.735 71.635 179.115 ;
        RECT 71.815 178.905 72.075 179.410 ;
        RECT 72.250 178.735 72.510 179.575 ;
        RECT 72.685 179.480 72.855 180.210 ;
        RECT 73.110 180.185 73.825 180.355 ;
        RECT 73.110 179.975 73.280 180.185 ;
        RECT 74.090 180.135 74.350 181.285 ;
        RECT 74.525 180.210 74.780 181.115 ;
        RECT 74.950 180.525 75.280 181.285 ;
        RECT 75.495 180.355 75.665 181.115 ;
        RECT 73.025 179.645 73.280 179.975 ;
        RECT 72.685 178.905 72.940 179.480 ;
        RECT 73.110 179.455 73.280 179.645 ;
        RECT 73.560 179.635 73.915 180.005 ;
        RECT 73.110 179.285 73.825 179.455 ;
        RECT 73.110 178.735 73.440 179.115 ;
        RECT 73.655 178.905 73.825 179.285 ;
        RECT 74.090 178.735 74.350 179.575 ;
        RECT 74.525 179.480 74.695 180.210 ;
        RECT 74.950 180.185 75.665 180.355 ;
        RECT 74.950 179.975 75.120 180.185 ;
        RECT 75.925 180.120 76.215 181.285 ;
        RECT 76.390 180.135 76.650 181.285 ;
        RECT 76.825 180.210 77.080 181.115 ;
        RECT 77.250 180.525 77.580 181.285 ;
        RECT 77.795 180.355 77.965 181.115 ;
        RECT 74.865 179.645 75.120 179.975 ;
        RECT 74.525 178.905 74.780 179.480 ;
        RECT 74.950 179.455 75.120 179.645 ;
        RECT 75.400 179.635 75.755 180.005 ;
        RECT 74.950 179.285 75.665 179.455 ;
        RECT 74.950 178.735 75.280 179.115 ;
        RECT 75.495 178.905 75.665 179.285 ;
        RECT 75.925 178.735 76.215 179.460 ;
        RECT 76.390 178.735 76.650 179.575 ;
        RECT 76.825 179.480 76.995 180.210 ;
        RECT 77.250 180.185 77.965 180.355 ;
        RECT 78.225 180.195 79.435 181.285 ;
        RECT 79.615 180.305 79.945 181.115 ;
        RECT 80.115 180.485 80.355 181.285 ;
        RECT 77.250 179.975 77.420 180.185 ;
        RECT 77.165 179.645 77.420 179.975 ;
        RECT 76.825 178.905 77.080 179.480 ;
        RECT 77.250 179.455 77.420 179.645 ;
        RECT 77.700 179.635 78.055 180.005 ;
        RECT 78.225 179.655 78.745 180.195 ;
        RECT 79.615 180.135 80.330 180.305 ;
        RECT 78.915 179.485 79.435 180.025 ;
        RECT 79.610 179.725 79.990 179.965 ;
        RECT 80.160 179.895 80.330 180.135 ;
        RECT 80.535 180.265 80.705 181.115 ;
        RECT 80.875 180.485 81.205 181.285 ;
        RECT 81.375 180.265 81.545 181.115 ;
        RECT 80.535 180.095 81.545 180.265 ;
        RECT 81.715 180.135 82.045 181.285 ;
        RECT 82.570 180.315 82.900 181.115 ;
        RECT 83.070 180.485 83.400 181.285 ;
        RECT 83.700 180.315 84.030 181.115 ;
        RECT 84.675 180.485 84.925 181.285 ;
        RECT 82.570 180.145 85.005 180.315 ;
        RECT 85.195 180.145 85.365 181.285 ;
        RECT 85.535 180.145 85.875 181.115 ;
        RECT 80.160 179.725 80.660 179.895 ;
        RECT 80.160 179.555 80.330 179.725 ;
        RECT 81.050 179.555 81.545 180.095 ;
        RECT 82.365 179.725 82.715 179.975 ;
        RECT 77.250 179.285 77.965 179.455 ;
        RECT 77.250 178.735 77.580 179.115 ;
        RECT 77.795 178.905 77.965 179.285 ;
        RECT 78.225 178.735 79.435 179.485 ;
        RECT 79.695 179.385 80.330 179.555 ;
        RECT 80.535 179.385 81.545 179.555 ;
        RECT 79.695 178.905 79.865 179.385 ;
        RECT 80.045 178.735 80.285 179.215 ;
        RECT 80.535 178.905 80.705 179.385 ;
        RECT 80.875 178.735 81.205 179.215 ;
        RECT 81.375 178.905 81.545 179.385 ;
        RECT 81.715 178.735 82.045 179.535 ;
        RECT 82.900 179.515 83.070 180.145 ;
        RECT 83.240 179.725 83.570 179.925 ;
        RECT 83.740 179.725 84.070 179.925 ;
        RECT 84.240 179.725 84.660 179.925 ;
        RECT 84.835 179.895 85.005 180.145 ;
        RECT 84.835 179.725 85.530 179.895 ;
        RECT 82.570 178.905 83.070 179.515 ;
        RECT 83.700 179.385 84.925 179.555 ;
        RECT 85.700 179.535 85.875 180.145 ;
        RECT 83.700 178.905 84.030 179.385 ;
        RECT 84.200 178.735 84.425 179.195 ;
        RECT 84.595 178.905 84.925 179.385 ;
        RECT 85.115 178.735 85.365 179.535 ;
        RECT 85.535 178.905 85.875 179.535 ;
        RECT 86.420 180.305 86.675 180.975 ;
        RECT 86.855 180.485 87.140 181.285 ;
        RECT 87.320 180.565 87.650 181.075 ;
        RECT 86.420 179.445 86.600 180.305 ;
        RECT 87.320 179.975 87.570 180.565 ;
        RECT 87.920 180.415 88.090 181.025 ;
        RECT 88.260 180.595 88.590 181.285 ;
        RECT 88.820 180.735 89.060 181.025 ;
        RECT 89.260 180.905 89.680 181.285 ;
        RECT 89.860 180.815 90.490 181.065 ;
        RECT 90.960 180.905 91.290 181.285 ;
        RECT 89.860 180.735 90.030 180.815 ;
        RECT 91.460 180.735 91.630 181.025 ;
        RECT 91.810 180.905 92.190 181.285 ;
        RECT 92.430 180.900 93.260 181.070 ;
        RECT 88.820 180.565 90.030 180.735 ;
        RECT 86.770 179.645 87.570 179.975 ;
        RECT 86.420 179.245 86.675 179.445 ;
        RECT 86.335 179.075 86.675 179.245 ;
        RECT 86.420 178.915 86.675 179.075 ;
        RECT 86.855 178.735 87.140 179.195 ;
        RECT 87.320 178.995 87.570 179.645 ;
        RECT 87.770 180.395 88.090 180.415 ;
        RECT 87.770 180.225 89.690 180.395 ;
        RECT 87.770 179.330 87.960 180.225 ;
        RECT 89.860 180.055 90.030 180.565 ;
        RECT 90.200 180.305 90.720 180.615 ;
        RECT 88.130 179.885 90.030 180.055 ;
        RECT 88.130 179.825 88.460 179.885 ;
        RECT 88.610 179.655 88.940 179.715 ;
        RECT 88.280 179.385 88.940 179.655 ;
        RECT 87.770 179.000 88.090 179.330 ;
        RECT 88.270 178.735 88.930 179.215 ;
        RECT 89.130 179.125 89.300 179.885 ;
        RECT 90.200 179.715 90.380 180.125 ;
        RECT 89.470 179.545 89.800 179.665 ;
        RECT 90.550 179.545 90.720 180.305 ;
        RECT 89.470 179.375 90.720 179.545 ;
        RECT 90.890 180.485 92.260 180.735 ;
        RECT 90.890 179.715 91.080 180.485 ;
        RECT 92.010 180.225 92.260 180.485 ;
        RECT 91.250 180.055 91.500 180.215 ;
        RECT 92.430 180.055 92.600 180.900 ;
        RECT 93.495 180.615 93.665 181.115 ;
        RECT 93.835 180.785 94.165 181.285 ;
        RECT 92.770 180.225 93.270 180.605 ;
        RECT 93.495 180.445 94.190 180.615 ;
        RECT 91.250 179.885 92.600 180.055 ;
        RECT 92.180 179.845 92.600 179.885 ;
        RECT 90.890 179.375 91.310 179.715 ;
        RECT 91.600 179.385 92.010 179.715 ;
        RECT 89.130 178.955 89.980 179.125 ;
        RECT 90.540 178.735 90.860 179.195 ;
        RECT 91.060 178.945 91.310 179.375 ;
        RECT 91.600 178.735 92.010 179.175 ;
        RECT 92.180 179.115 92.350 179.845 ;
        RECT 92.520 179.295 92.870 179.665 ;
        RECT 93.050 179.355 93.270 180.225 ;
        RECT 93.440 179.655 93.850 180.275 ;
        RECT 94.020 179.475 94.190 180.445 ;
        RECT 93.495 179.285 94.190 179.475 ;
        RECT 92.180 178.915 93.195 179.115 ;
        RECT 93.495 178.955 93.665 179.285 ;
        RECT 93.835 178.735 94.165 179.115 ;
        RECT 94.380 178.995 94.605 181.115 ;
        RECT 94.775 180.785 95.105 181.285 ;
        RECT 95.275 180.615 95.445 181.115 ;
        RECT 94.780 180.445 95.445 180.615 ;
        RECT 94.780 179.455 95.010 180.445 ;
        RECT 95.180 179.625 95.530 180.275 ;
        RECT 95.745 180.145 95.975 181.285 ;
        RECT 96.145 180.135 96.475 181.115 ;
        RECT 96.645 180.145 96.855 181.285 ;
        RECT 98.120 180.655 98.405 181.115 ;
        RECT 98.575 180.825 98.845 181.285 ;
        RECT 98.120 180.435 99.075 180.655 ;
        RECT 95.725 179.725 96.055 179.975 ;
        RECT 94.780 179.285 95.445 179.455 ;
        RECT 94.775 178.735 95.105 179.115 ;
        RECT 95.275 178.995 95.445 179.285 ;
        RECT 95.745 178.735 95.975 179.555 ;
        RECT 96.225 179.535 96.475 180.135 ;
        RECT 98.005 179.705 98.695 180.265 ;
        RECT 96.145 178.905 96.475 179.535 ;
        RECT 96.645 178.735 96.855 179.555 ;
        RECT 98.865 179.535 99.075 180.435 ;
        RECT 98.120 179.365 99.075 179.535 ;
        RECT 99.245 180.265 99.645 181.115 ;
        RECT 99.835 180.655 100.115 181.115 ;
        RECT 100.635 180.825 100.960 181.285 ;
        RECT 99.835 180.435 100.960 180.655 ;
        RECT 99.245 179.705 100.340 180.265 ;
        RECT 100.510 179.975 100.960 180.435 ;
        RECT 101.130 180.145 101.515 181.115 ;
        RECT 98.120 178.905 98.405 179.365 ;
        RECT 98.575 178.735 98.845 179.195 ;
        RECT 99.245 178.905 99.645 179.705 ;
        RECT 100.510 179.645 101.065 179.975 ;
        RECT 100.510 179.535 100.960 179.645 ;
        RECT 99.835 179.365 100.960 179.535 ;
        RECT 101.235 179.475 101.515 180.145 ;
        RECT 101.685 180.120 101.975 181.285 ;
        RECT 102.235 180.355 102.405 181.115 ;
        RECT 102.585 180.525 102.915 181.285 ;
        RECT 102.235 180.185 102.900 180.355 ;
        RECT 103.085 180.210 103.355 181.115 ;
        RECT 102.730 180.040 102.900 180.185 ;
        RECT 102.165 179.635 102.495 180.005 ;
        RECT 102.730 179.710 103.015 180.040 ;
        RECT 99.835 178.905 100.115 179.365 ;
        RECT 100.635 178.735 100.960 179.195 ;
        RECT 101.130 178.905 101.515 179.475 ;
        RECT 101.685 178.735 101.975 179.460 ;
        RECT 102.730 179.455 102.900 179.710 ;
        RECT 102.235 179.285 102.900 179.455 ;
        RECT 103.185 179.410 103.355 180.210 ;
        RECT 103.985 180.195 105.655 181.285 ;
        RECT 106.030 180.315 106.360 181.115 ;
        RECT 106.530 180.485 106.860 181.285 ;
        RECT 107.160 180.315 107.490 181.115 ;
        RECT 108.135 180.485 108.385 181.285 ;
        RECT 103.985 179.675 104.735 180.195 ;
        RECT 106.030 180.145 108.465 180.315 ;
        RECT 108.655 180.145 108.825 181.285 ;
        RECT 108.995 180.145 109.335 181.115 ;
        RECT 104.905 179.505 105.655 180.025 ;
        RECT 105.825 179.725 106.175 179.975 ;
        RECT 106.360 179.515 106.530 180.145 ;
        RECT 106.700 179.725 107.030 179.925 ;
        RECT 107.200 179.725 107.530 179.925 ;
        RECT 107.700 179.725 108.120 179.925 ;
        RECT 108.295 179.895 108.465 180.145 ;
        RECT 108.295 179.725 108.990 179.895 ;
        RECT 102.235 178.905 102.405 179.285 ;
        RECT 102.585 178.735 102.915 179.115 ;
        RECT 103.095 178.905 103.355 179.410 ;
        RECT 103.985 178.735 105.655 179.505 ;
        RECT 106.030 178.905 106.530 179.515 ;
        RECT 107.160 179.385 108.385 179.555 ;
        RECT 109.160 179.535 109.335 180.145 ;
        RECT 107.160 178.905 107.490 179.385 ;
        RECT 107.660 178.735 107.885 179.195 ;
        RECT 108.055 178.905 108.385 179.385 ;
        RECT 108.575 178.735 108.825 179.535 ;
        RECT 108.995 178.905 109.335 179.535 ;
        RECT 109.505 180.145 109.845 181.115 ;
        RECT 110.015 180.145 110.185 181.285 ;
        RECT 110.455 180.485 110.705 181.285 ;
        RECT 111.350 180.315 111.680 181.115 ;
        RECT 111.980 180.485 112.310 181.285 ;
        RECT 112.480 180.315 112.810 181.115 ;
        RECT 113.300 180.655 113.585 181.115 ;
        RECT 113.755 180.825 114.025 181.285 ;
        RECT 113.300 180.435 114.255 180.655 ;
        RECT 110.375 180.145 112.810 180.315 ;
        RECT 109.505 179.535 109.680 180.145 ;
        RECT 110.375 179.895 110.545 180.145 ;
        RECT 109.850 179.725 110.545 179.895 ;
        RECT 110.720 179.725 111.140 179.925 ;
        RECT 111.310 179.725 111.640 179.925 ;
        RECT 111.810 179.725 112.140 179.925 ;
        RECT 109.505 178.905 109.845 179.535 ;
        RECT 110.015 178.735 110.265 179.535 ;
        RECT 110.455 179.385 111.680 179.555 ;
        RECT 110.455 178.905 110.785 179.385 ;
        RECT 110.955 178.735 111.180 179.195 ;
        RECT 111.350 178.905 111.680 179.385 ;
        RECT 112.310 179.515 112.480 180.145 ;
        RECT 112.665 179.725 113.015 179.975 ;
        RECT 113.185 179.705 113.875 180.265 ;
        RECT 114.045 179.535 114.255 180.435 ;
        RECT 112.310 178.905 112.810 179.515 ;
        RECT 113.300 179.365 114.255 179.535 ;
        RECT 114.425 180.265 114.825 181.115 ;
        RECT 115.015 180.655 115.295 181.115 ;
        RECT 115.815 180.825 116.140 181.285 ;
        RECT 115.015 180.435 116.140 180.655 ;
        RECT 114.425 179.705 115.520 180.265 ;
        RECT 115.690 179.975 116.140 180.435 ;
        RECT 116.310 180.145 116.695 181.115 ;
        RECT 113.300 178.905 113.585 179.365 ;
        RECT 113.755 178.735 114.025 179.195 ;
        RECT 114.425 178.905 114.825 179.705 ;
        RECT 115.690 179.645 116.245 179.975 ;
        RECT 115.690 179.535 116.140 179.645 ;
        RECT 115.015 179.365 116.140 179.535 ;
        RECT 116.415 179.475 116.695 180.145 ;
        RECT 115.015 178.905 115.295 179.365 ;
        RECT 115.815 178.735 116.140 179.195 ;
        RECT 116.310 178.905 116.695 179.475 ;
        RECT 116.870 180.095 117.125 180.975 ;
        RECT 117.295 180.145 117.600 181.285 ;
        RECT 117.940 180.905 118.270 181.285 ;
        RECT 118.450 180.735 118.620 181.025 ;
        RECT 118.790 180.825 119.040 181.285 ;
        RECT 117.820 180.565 118.620 180.735 ;
        RECT 119.210 180.775 120.080 181.115 ;
        RECT 116.870 179.445 117.080 180.095 ;
        RECT 117.820 179.975 117.990 180.565 ;
        RECT 119.210 180.395 119.380 180.775 ;
        RECT 120.315 180.655 120.485 181.115 ;
        RECT 120.655 180.825 121.025 181.285 ;
        RECT 121.320 180.685 121.490 181.025 ;
        RECT 121.660 180.855 121.990 181.285 ;
        RECT 122.225 180.685 122.395 181.025 ;
        RECT 118.160 180.225 119.380 180.395 ;
        RECT 119.550 180.315 120.010 180.605 ;
        RECT 120.315 180.485 120.875 180.655 ;
        RECT 121.320 180.515 122.395 180.685 ;
        RECT 122.565 180.785 123.245 181.115 ;
        RECT 123.460 180.785 123.710 181.115 ;
        RECT 123.880 180.825 124.130 181.285 ;
        RECT 120.705 180.345 120.875 180.485 ;
        RECT 119.550 180.305 120.515 180.315 ;
        RECT 119.210 180.135 119.380 180.225 ;
        RECT 119.840 180.145 120.515 180.305 ;
        RECT 117.250 179.945 117.990 179.975 ;
        RECT 117.250 179.645 118.165 179.945 ;
        RECT 117.840 179.470 118.165 179.645 ;
        RECT 116.870 178.915 117.125 179.445 ;
        RECT 117.295 178.735 117.600 179.195 ;
        RECT 117.845 179.115 118.165 179.470 ;
        RECT 118.335 179.685 118.875 180.055 ;
        RECT 119.210 179.965 119.615 180.135 ;
        RECT 118.335 179.285 118.575 179.685 ;
        RECT 119.055 179.515 119.275 179.795 ;
        RECT 118.745 179.345 119.275 179.515 ;
        RECT 118.745 179.115 118.915 179.345 ;
        RECT 119.445 179.185 119.615 179.965 ;
        RECT 119.785 179.355 120.135 179.975 ;
        RECT 120.305 179.355 120.515 180.145 ;
        RECT 120.705 180.175 122.205 180.345 ;
        RECT 120.705 179.485 120.875 180.175 ;
        RECT 122.565 180.005 122.735 180.785 ;
        RECT 123.540 180.655 123.710 180.785 ;
        RECT 121.045 179.835 122.735 180.005 ;
        RECT 122.905 180.225 123.370 180.615 ;
        RECT 123.540 180.485 123.935 180.655 ;
        RECT 121.045 179.655 121.215 179.835 ;
        RECT 117.845 178.945 118.915 179.115 ;
        RECT 119.085 178.735 119.275 179.175 ;
        RECT 119.445 178.905 120.395 179.185 ;
        RECT 120.705 179.095 120.965 179.485 ;
        RECT 121.385 179.415 122.175 179.665 ;
        RECT 120.615 178.925 120.965 179.095 ;
        RECT 121.175 178.735 121.505 179.195 ;
        RECT 122.380 179.125 122.550 179.835 ;
        RECT 122.905 179.635 123.075 180.225 ;
        RECT 122.720 179.415 123.075 179.635 ;
        RECT 123.245 179.415 123.595 180.035 ;
        RECT 123.765 179.125 123.935 180.485 ;
        RECT 124.300 180.315 124.625 181.100 ;
        RECT 124.105 179.265 124.565 180.315 ;
        RECT 122.380 178.955 123.235 179.125 ;
        RECT 123.440 178.955 123.935 179.125 ;
        RECT 124.105 178.735 124.435 179.095 ;
        RECT 124.795 178.995 124.965 181.115 ;
        RECT 125.135 180.785 125.465 181.285 ;
        RECT 125.635 180.615 125.890 181.115 ;
        RECT 125.140 180.445 125.890 180.615 ;
        RECT 125.140 179.455 125.370 180.445 ;
        RECT 125.540 179.625 125.890 180.275 ;
        RECT 126.525 180.195 127.735 181.285 ;
        RECT 126.525 179.655 127.045 180.195 ;
        RECT 127.215 179.485 127.735 180.025 ;
        RECT 125.140 179.285 125.890 179.455 ;
        RECT 125.135 178.735 125.465 179.115 ;
        RECT 125.635 178.995 125.890 179.285 ;
        RECT 126.525 178.735 127.735 179.485 ;
        RECT 29.840 178.565 127.820 178.735 ;
        RECT 29.925 177.815 31.135 178.565 ;
        RECT 29.925 177.275 30.445 177.815 ;
        RECT 31.765 177.795 34.355 178.565 ;
        RECT 34.615 178.015 34.785 178.395 ;
        RECT 34.965 178.185 35.295 178.565 ;
        RECT 34.615 177.845 35.280 178.015 ;
        RECT 35.475 177.890 35.735 178.395 ;
        RECT 30.615 177.105 31.135 177.645 ;
        RECT 29.925 176.015 31.135 177.105 ;
        RECT 31.765 177.105 32.975 177.625 ;
        RECT 33.145 177.275 34.355 177.795 ;
        RECT 34.545 177.295 34.875 177.665 ;
        RECT 35.110 177.590 35.280 177.845 ;
        RECT 35.110 177.260 35.395 177.590 ;
        RECT 35.110 177.115 35.280 177.260 ;
        RECT 31.765 176.015 34.355 177.105 ;
        RECT 34.615 176.945 35.280 177.115 ;
        RECT 35.565 177.090 35.735 177.890 ;
        RECT 35.945 177.745 36.175 178.565 ;
        RECT 36.345 177.765 36.675 178.395 ;
        RECT 35.925 177.325 36.255 177.575 ;
        RECT 36.425 177.165 36.675 177.765 ;
        RECT 36.845 177.745 37.055 178.565 ;
        RECT 37.285 177.840 37.575 178.565 ;
        RECT 37.750 178.015 38.005 178.305 ;
        RECT 38.175 178.185 38.505 178.565 ;
        RECT 37.750 177.845 38.500 178.015 ;
        RECT 34.615 176.185 34.785 176.945 ;
        RECT 34.965 176.015 35.295 176.775 ;
        RECT 35.465 176.185 35.735 177.090 ;
        RECT 35.945 176.015 36.175 177.155 ;
        RECT 36.345 176.185 36.675 177.165 ;
        RECT 36.845 176.015 37.055 177.155 ;
        RECT 37.285 176.015 37.575 177.180 ;
        RECT 37.750 177.025 38.100 177.675 ;
        RECT 38.270 176.855 38.500 177.845 ;
        RECT 37.750 176.685 38.500 176.855 ;
        RECT 37.750 176.185 38.005 176.685 ;
        RECT 38.175 176.015 38.505 176.515 ;
        RECT 38.675 176.185 38.845 178.305 ;
        RECT 39.205 178.205 39.535 178.565 ;
        RECT 39.705 178.175 40.200 178.345 ;
        RECT 40.405 178.175 41.260 178.345 ;
        RECT 39.075 176.985 39.535 178.035 ;
        RECT 39.015 176.200 39.340 176.985 ;
        RECT 39.705 176.815 39.875 178.175 ;
        RECT 40.045 177.265 40.395 177.885 ;
        RECT 40.565 177.665 40.920 177.885 ;
        RECT 40.565 177.075 40.735 177.665 ;
        RECT 41.090 177.465 41.260 178.175 ;
        RECT 42.135 178.105 42.465 178.565 ;
        RECT 42.675 178.205 43.025 178.375 ;
        RECT 41.465 177.635 42.255 177.885 ;
        RECT 42.675 177.815 42.935 178.205 ;
        RECT 43.245 178.115 44.195 178.395 ;
        RECT 44.365 178.125 44.555 178.565 ;
        RECT 44.725 178.185 45.795 178.355 ;
        RECT 42.425 177.465 42.595 177.645 ;
        RECT 39.705 176.645 40.100 176.815 ;
        RECT 40.270 176.685 40.735 177.075 ;
        RECT 40.905 177.295 42.595 177.465 ;
        RECT 39.930 176.515 40.100 176.645 ;
        RECT 40.905 176.515 41.075 177.295 ;
        RECT 42.765 177.125 42.935 177.815 ;
        RECT 41.435 176.955 42.935 177.125 ;
        RECT 43.125 177.155 43.335 177.945 ;
        RECT 43.505 177.325 43.855 177.945 ;
        RECT 44.025 177.335 44.195 178.115 ;
        RECT 44.725 177.955 44.895 178.185 ;
        RECT 44.365 177.785 44.895 177.955 ;
        RECT 44.365 177.505 44.585 177.785 ;
        RECT 45.065 177.615 45.305 178.015 ;
        RECT 44.025 177.165 44.430 177.335 ;
        RECT 44.765 177.245 45.305 177.615 ;
        RECT 45.475 177.830 45.795 178.185 ;
        RECT 46.040 178.105 46.345 178.565 ;
        RECT 46.515 177.855 46.770 178.385 ;
        RECT 45.475 177.655 45.800 177.830 ;
        RECT 45.475 177.355 46.390 177.655 ;
        RECT 45.650 177.325 46.390 177.355 ;
        RECT 43.125 176.995 43.800 177.155 ;
        RECT 44.260 177.075 44.430 177.165 ;
        RECT 43.125 176.985 44.090 176.995 ;
        RECT 42.765 176.815 42.935 176.955 ;
        RECT 39.510 176.015 39.760 176.475 ;
        RECT 39.930 176.185 40.180 176.515 ;
        RECT 40.395 176.185 41.075 176.515 ;
        RECT 41.245 176.615 42.320 176.785 ;
        RECT 42.765 176.645 43.325 176.815 ;
        RECT 43.630 176.695 44.090 176.985 ;
        RECT 44.260 176.905 45.480 177.075 ;
        RECT 41.245 176.275 41.415 176.615 ;
        RECT 41.650 176.015 41.980 176.445 ;
        RECT 42.150 176.275 42.320 176.615 ;
        RECT 42.615 176.015 42.985 176.475 ;
        RECT 43.155 176.185 43.325 176.645 ;
        RECT 44.260 176.525 44.430 176.905 ;
        RECT 45.650 176.735 45.820 177.325 ;
        RECT 46.560 177.205 46.770 177.855 ;
        RECT 43.560 176.185 44.430 176.525 ;
        RECT 45.020 176.565 45.820 176.735 ;
        RECT 44.600 176.015 44.850 176.475 ;
        RECT 45.020 176.275 45.190 176.565 ;
        RECT 45.370 176.015 45.700 176.395 ;
        RECT 46.040 176.015 46.345 177.155 ;
        RECT 46.515 176.325 46.770 177.205 ;
        RECT 46.945 177.765 47.285 178.395 ;
        RECT 47.455 177.765 47.705 178.565 ;
        RECT 47.895 177.915 48.225 178.395 ;
        RECT 48.395 178.105 48.620 178.565 ;
        RECT 48.790 177.915 49.120 178.395 ;
        RECT 46.945 177.155 47.120 177.765 ;
        RECT 47.895 177.745 49.120 177.915 ;
        RECT 49.750 177.785 50.250 178.395 ;
        RECT 50.630 178.015 50.885 178.305 ;
        RECT 51.055 178.185 51.385 178.565 ;
        RECT 50.630 177.845 51.380 178.015 ;
        RECT 47.290 177.405 47.985 177.575 ;
        RECT 47.815 177.155 47.985 177.405 ;
        RECT 48.160 177.375 48.580 177.575 ;
        RECT 48.750 177.375 49.080 177.575 ;
        RECT 49.250 177.375 49.580 177.575 ;
        RECT 49.750 177.155 49.920 177.785 ;
        RECT 50.105 177.325 50.455 177.575 ;
        RECT 46.945 176.185 47.285 177.155 ;
        RECT 47.455 176.015 47.625 177.155 ;
        RECT 47.815 176.985 50.250 177.155 ;
        RECT 50.630 177.025 50.980 177.675 ;
        RECT 47.895 176.015 48.145 176.815 ;
        RECT 48.790 176.185 49.120 176.985 ;
        RECT 49.420 176.015 49.750 176.815 ;
        RECT 49.920 176.185 50.250 176.985 ;
        RECT 51.150 176.855 51.380 177.845 ;
        RECT 50.630 176.685 51.380 176.855 ;
        RECT 50.630 176.185 50.885 176.685 ;
        RECT 51.055 176.015 51.385 176.515 ;
        RECT 51.555 176.185 51.725 178.305 ;
        RECT 52.085 178.205 52.415 178.565 ;
        RECT 52.585 178.175 53.080 178.345 ;
        RECT 53.285 178.175 54.140 178.345 ;
        RECT 51.955 176.985 52.415 178.035 ;
        RECT 51.895 176.200 52.220 176.985 ;
        RECT 52.585 176.815 52.755 178.175 ;
        RECT 52.925 177.265 53.275 177.885 ;
        RECT 53.445 177.665 53.800 177.885 ;
        RECT 53.445 177.075 53.615 177.665 ;
        RECT 53.970 177.465 54.140 178.175 ;
        RECT 55.015 178.105 55.345 178.565 ;
        RECT 55.555 178.205 55.905 178.375 ;
        RECT 54.345 177.635 55.135 177.885 ;
        RECT 55.555 177.815 55.815 178.205 ;
        RECT 56.125 178.115 57.075 178.395 ;
        RECT 57.245 178.125 57.435 178.565 ;
        RECT 57.605 178.185 58.675 178.355 ;
        RECT 55.305 177.465 55.475 177.645 ;
        RECT 52.585 176.645 52.980 176.815 ;
        RECT 53.150 176.685 53.615 177.075 ;
        RECT 53.785 177.295 55.475 177.465 ;
        RECT 52.810 176.515 52.980 176.645 ;
        RECT 53.785 176.515 53.955 177.295 ;
        RECT 55.645 177.125 55.815 177.815 ;
        RECT 54.315 176.955 55.815 177.125 ;
        RECT 56.005 177.155 56.215 177.945 ;
        RECT 56.385 177.325 56.735 177.945 ;
        RECT 56.905 177.335 57.075 178.115 ;
        RECT 57.605 177.955 57.775 178.185 ;
        RECT 57.245 177.785 57.775 177.955 ;
        RECT 57.245 177.505 57.465 177.785 ;
        RECT 57.945 177.615 58.185 178.015 ;
        RECT 56.905 177.165 57.310 177.335 ;
        RECT 57.645 177.245 58.185 177.615 ;
        RECT 58.355 177.830 58.675 178.185 ;
        RECT 58.920 178.105 59.225 178.565 ;
        RECT 59.395 177.855 59.650 178.385 ;
        RECT 58.355 177.655 58.680 177.830 ;
        RECT 58.355 177.355 59.270 177.655 ;
        RECT 58.530 177.325 59.270 177.355 ;
        RECT 56.005 176.995 56.680 177.155 ;
        RECT 57.140 177.075 57.310 177.165 ;
        RECT 56.005 176.985 56.970 176.995 ;
        RECT 55.645 176.815 55.815 176.955 ;
        RECT 52.390 176.015 52.640 176.475 ;
        RECT 52.810 176.185 53.060 176.515 ;
        RECT 53.275 176.185 53.955 176.515 ;
        RECT 54.125 176.615 55.200 176.785 ;
        RECT 55.645 176.645 56.205 176.815 ;
        RECT 56.510 176.695 56.970 176.985 ;
        RECT 57.140 176.905 58.360 177.075 ;
        RECT 54.125 176.275 54.295 176.615 ;
        RECT 54.530 176.015 54.860 176.445 ;
        RECT 55.030 176.275 55.200 176.615 ;
        RECT 55.495 176.015 55.865 176.475 ;
        RECT 56.035 176.185 56.205 176.645 ;
        RECT 57.140 176.525 57.310 176.905 ;
        RECT 58.530 176.735 58.700 177.325 ;
        RECT 59.440 177.205 59.650 177.855 ;
        RECT 60.375 178.015 60.545 178.395 ;
        RECT 60.725 178.185 61.055 178.565 ;
        RECT 60.375 177.845 61.040 178.015 ;
        RECT 61.235 177.890 61.495 178.395 ;
        RECT 60.305 177.295 60.635 177.665 ;
        RECT 60.870 177.590 61.040 177.845 ;
        RECT 56.440 176.185 57.310 176.525 ;
        RECT 57.900 176.565 58.700 176.735 ;
        RECT 57.480 176.015 57.730 176.475 ;
        RECT 57.900 176.275 58.070 176.565 ;
        RECT 58.250 176.015 58.580 176.395 ;
        RECT 58.920 176.015 59.225 177.155 ;
        RECT 59.395 176.325 59.650 177.205 ;
        RECT 60.870 177.260 61.155 177.590 ;
        RECT 60.870 177.115 61.040 177.260 ;
        RECT 60.375 176.945 61.040 177.115 ;
        RECT 61.325 177.090 61.495 177.890 ;
        RECT 61.665 177.815 62.875 178.565 ;
        RECT 63.045 177.840 63.335 178.565 ;
        RECT 63.620 177.935 63.905 178.395 ;
        RECT 64.075 178.105 64.345 178.565 ;
        RECT 60.375 176.185 60.545 176.945 ;
        RECT 60.725 176.015 61.055 176.775 ;
        RECT 61.225 176.185 61.495 177.090 ;
        RECT 61.665 177.105 62.185 177.645 ;
        RECT 62.355 177.275 62.875 177.815 ;
        RECT 63.620 177.765 64.575 177.935 ;
        RECT 61.665 176.015 62.875 177.105 ;
        RECT 63.045 176.015 63.335 177.180 ;
        RECT 63.505 177.035 64.195 177.595 ;
        RECT 64.365 176.865 64.575 177.765 ;
        RECT 63.620 176.645 64.575 176.865 ;
        RECT 64.745 177.595 65.145 178.395 ;
        RECT 65.335 177.935 65.615 178.395 ;
        RECT 66.135 178.105 66.460 178.565 ;
        RECT 65.335 177.765 66.460 177.935 ;
        RECT 66.630 177.825 67.015 178.395 ;
        RECT 66.010 177.655 66.460 177.765 ;
        RECT 64.745 177.035 65.840 177.595 ;
        RECT 66.010 177.325 66.565 177.655 ;
        RECT 63.620 176.185 63.905 176.645 ;
        RECT 64.075 176.015 64.345 176.475 ;
        RECT 64.745 176.185 65.145 177.035 ;
        RECT 66.010 176.865 66.460 177.325 ;
        RECT 66.735 177.155 67.015 177.825 ;
        RECT 67.185 177.795 70.695 178.565 ;
        RECT 65.335 176.645 66.460 176.865 ;
        RECT 65.335 176.185 65.615 176.645 ;
        RECT 66.135 176.015 66.460 176.475 ;
        RECT 66.630 176.185 67.015 177.155 ;
        RECT 67.185 177.105 68.875 177.625 ;
        RECT 69.045 177.275 70.695 177.795 ;
        RECT 70.925 177.745 71.135 178.565 ;
        RECT 71.305 177.765 71.635 178.395 ;
        RECT 71.305 177.165 71.555 177.765 ;
        RECT 71.805 177.745 72.035 178.565 ;
        RECT 72.245 177.795 74.835 178.565 ;
        RECT 71.725 177.325 72.055 177.575 ;
        RECT 67.185 176.015 70.695 177.105 ;
        RECT 70.925 176.015 71.135 177.155 ;
        RECT 71.305 176.185 71.635 177.165 ;
        RECT 71.805 176.015 72.035 177.155 ;
        RECT 72.245 177.105 73.455 177.625 ;
        RECT 73.625 177.275 74.835 177.795 ;
        RECT 75.010 177.725 75.270 178.565 ;
        RECT 75.445 177.820 75.700 178.395 ;
        RECT 75.870 178.185 76.200 178.565 ;
        RECT 76.415 178.015 76.585 178.395 ;
        RECT 75.870 177.845 76.585 178.015 ;
        RECT 76.845 178.065 77.145 178.395 ;
        RECT 77.315 178.085 77.590 178.565 ;
        RECT 72.245 176.015 74.835 177.105 ;
        RECT 75.010 176.015 75.270 177.165 ;
        RECT 75.445 177.090 75.615 177.820 ;
        RECT 75.870 177.655 76.040 177.845 ;
        RECT 75.785 177.325 76.040 177.655 ;
        RECT 75.870 177.115 76.040 177.325 ;
        RECT 76.320 177.295 76.675 177.665 ;
        RECT 76.845 177.155 77.015 178.065 ;
        RECT 77.770 177.915 78.065 178.305 ;
        RECT 78.235 178.085 78.490 178.565 ;
        RECT 78.665 177.915 78.925 178.305 ;
        RECT 79.095 178.085 79.375 178.565 ;
        RECT 79.615 178.035 79.945 178.395 ;
        RECT 80.115 178.205 80.445 178.565 ;
        RECT 80.645 178.035 80.975 178.395 ;
        RECT 77.185 177.325 77.535 177.895 ;
        RECT 77.770 177.745 79.420 177.915 ;
        RECT 79.615 177.825 80.975 178.035 ;
        RECT 81.485 177.805 82.195 178.395 ;
        RECT 77.705 177.405 78.845 177.575 ;
        RECT 77.705 177.155 77.875 177.405 ;
        RECT 79.015 177.235 79.420 177.745 ;
        RECT 79.605 177.325 79.915 177.655 ;
        RECT 80.125 177.325 80.500 177.655 ;
        RECT 80.820 177.325 81.315 177.655 ;
        RECT 75.445 176.185 75.700 177.090 ;
        RECT 75.870 176.945 76.585 177.115 ;
        RECT 75.870 176.015 76.200 176.775 ;
        RECT 76.415 176.185 76.585 176.945 ;
        RECT 76.845 176.985 77.875 177.155 ;
        RECT 78.665 177.065 79.420 177.235 ;
        RECT 76.845 176.185 77.155 176.985 ;
        RECT 78.665 176.815 78.925 177.065 ;
        RECT 77.325 176.015 77.635 176.815 ;
        RECT 77.805 176.645 78.925 176.815 ;
        RECT 77.805 176.185 78.065 176.645 ;
        RECT 78.235 176.015 78.490 176.475 ;
        RECT 78.665 176.185 78.925 176.645 ;
        RECT 79.095 176.015 79.380 176.885 ;
        RECT 79.615 176.015 79.945 177.075 ;
        RECT 80.125 176.400 80.295 177.325 ;
        RECT 80.465 176.835 80.795 177.055 ;
        RECT 80.990 177.035 81.315 177.325 ;
        RECT 81.490 177.035 81.820 177.575 ;
        RECT 81.990 176.835 82.195 177.805 ;
        RECT 82.825 177.795 84.495 178.565 ;
        RECT 80.465 176.605 82.195 176.835 ;
        RECT 80.465 176.205 80.795 176.605 ;
        RECT 80.965 176.015 81.295 176.375 ;
        RECT 81.495 176.185 82.195 176.605 ;
        RECT 82.825 177.105 83.575 177.625 ;
        RECT 83.745 177.275 84.495 177.795 ;
        RECT 84.665 177.825 85.050 178.395 ;
        RECT 85.220 178.105 85.545 178.565 ;
        RECT 86.065 177.935 86.345 178.395 ;
        RECT 84.665 177.155 84.945 177.825 ;
        RECT 85.220 177.765 86.345 177.935 ;
        RECT 85.220 177.655 85.670 177.765 ;
        RECT 85.115 177.325 85.670 177.655 ;
        RECT 86.535 177.595 86.935 178.395 ;
        RECT 87.335 178.105 87.605 178.565 ;
        RECT 87.775 177.935 88.060 178.395 ;
        RECT 82.825 176.015 84.495 177.105 ;
        RECT 84.665 176.185 85.050 177.155 ;
        RECT 85.220 176.865 85.670 177.325 ;
        RECT 85.840 177.035 86.935 177.595 ;
        RECT 85.220 176.645 86.345 176.865 ;
        RECT 85.220 176.015 85.545 176.475 ;
        RECT 86.065 176.185 86.345 176.645 ;
        RECT 86.535 176.185 86.935 177.035 ;
        RECT 87.105 177.765 88.060 177.935 ;
        RECT 88.805 177.840 89.095 178.565 ;
        RECT 87.105 176.865 87.315 177.765 ;
        RECT 89.305 177.745 89.535 178.565 ;
        RECT 89.705 177.765 90.035 178.395 ;
        RECT 87.485 177.035 88.175 177.595 ;
        RECT 89.285 177.325 89.615 177.575 ;
        RECT 87.105 176.645 88.060 176.865 ;
        RECT 87.335 176.015 87.605 176.475 ;
        RECT 87.775 176.185 88.060 176.645 ;
        RECT 88.805 176.015 89.095 177.180 ;
        RECT 89.785 177.165 90.035 177.765 ;
        RECT 90.205 177.745 90.415 178.565 ;
        RECT 90.760 177.935 91.045 178.395 ;
        RECT 91.215 178.105 91.485 178.565 ;
        RECT 90.760 177.765 91.715 177.935 ;
        RECT 89.305 176.015 89.535 177.155 ;
        RECT 89.705 176.185 90.035 177.165 ;
        RECT 90.205 176.015 90.415 177.155 ;
        RECT 90.645 177.035 91.335 177.595 ;
        RECT 91.505 176.865 91.715 177.765 ;
        RECT 90.760 176.645 91.715 176.865 ;
        RECT 91.885 177.595 92.285 178.395 ;
        RECT 92.475 177.935 92.755 178.395 ;
        RECT 93.275 178.105 93.600 178.565 ;
        RECT 92.475 177.765 93.600 177.935 ;
        RECT 93.770 177.825 94.155 178.395 ;
        RECT 93.150 177.655 93.600 177.765 ;
        RECT 91.885 177.035 92.980 177.595 ;
        RECT 93.150 177.325 93.705 177.655 ;
        RECT 90.760 176.185 91.045 176.645 ;
        RECT 91.215 176.015 91.485 176.475 ;
        RECT 91.885 176.185 92.285 177.035 ;
        RECT 93.150 176.865 93.600 177.325 ;
        RECT 93.875 177.155 94.155 177.825 ;
        RECT 92.475 176.645 93.600 176.865 ;
        RECT 92.475 176.185 92.755 176.645 ;
        RECT 93.275 176.015 93.600 176.475 ;
        RECT 93.770 176.185 94.155 177.155 ;
        RECT 94.325 177.890 94.585 178.395 ;
        RECT 94.765 178.185 95.095 178.565 ;
        RECT 95.275 178.015 95.445 178.395 ;
        RECT 94.325 177.090 94.495 177.890 ;
        RECT 94.780 177.845 95.445 178.015 ;
        RECT 96.630 177.855 96.885 178.385 ;
        RECT 97.055 178.105 97.360 178.565 ;
        RECT 97.605 178.185 98.675 178.355 ;
        RECT 94.780 177.590 94.950 177.845 ;
        RECT 94.665 177.260 94.950 177.590 ;
        RECT 95.185 177.295 95.515 177.665 ;
        RECT 94.780 177.115 94.950 177.260 ;
        RECT 96.630 177.205 96.840 177.855 ;
        RECT 97.605 177.830 97.925 178.185 ;
        RECT 97.600 177.655 97.925 177.830 ;
        RECT 97.010 177.355 97.925 177.655 ;
        RECT 98.095 177.615 98.335 178.015 ;
        RECT 98.505 177.955 98.675 178.185 ;
        RECT 98.845 178.125 99.035 178.565 ;
        RECT 99.205 178.115 100.155 178.395 ;
        RECT 100.375 178.205 100.725 178.375 ;
        RECT 98.505 177.785 99.035 177.955 ;
        RECT 97.010 177.325 97.750 177.355 ;
        RECT 94.325 176.185 94.595 177.090 ;
        RECT 94.780 176.945 95.445 177.115 ;
        RECT 94.765 176.015 95.095 176.775 ;
        RECT 95.275 176.185 95.445 176.945 ;
        RECT 96.630 176.325 96.885 177.205 ;
        RECT 97.055 176.015 97.360 177.155 ;
        RECT 97.580 176.735 97.750 177.325 ;
        RECT 98.095 177.245 98.635 177.615 ;
        RECT 98.815 177.505 99.035 177.785 ;
        RECT 99.205 177.335 99.375 178.115 ;
        RECT 98.970 177.165 99.375 177.335 ;
        RECT 99.545 177.325 99.895 177.945 ;
        RECT 98.970 177.075 99.140 177.165 ;
        RECT 100.065 177.155 100.275 177.945 ;
        RECT 97.920 176.905 99.140 177.075 ;
        RECT 99.600 176.995 100.275 177.155 ;
        RECT 97.580 176.565 98.380 176.735 ;
        RECT 97.700 176.015 98.030 176.395 ;
        RECT 98.210 176.275 98.380 176.565 ;
        RECT 98.970 176.525 99.140 176.905 ;
        RECT 99.310 176.985 100.275 176.995 ;
        RECT 100.465 177.815 100.725 178.205 ;
        RECT 100.935 178.105 101.265 178.565 ;
        RECT 102.140 178.175 102.995 178.345 ;
        RECT 103.200 178.175 103.695 178.345 ;
        RECT 103.865 178.205 104.195 178.565 ;
        RECT 100.465 177.125 100.635 177.815 ;
        RECT 100.805 177.465 100.975 177.645 ;
        RECT 101.145 177.635 101.935 177.885 ;
        RECT 102.140 177.465 102.310 178.175 ;
        RECT 102.480 177.665 102.835 177.885 ;
        RECT 100.805 177.295 102.495 177.465 ;
        RECT 99.310 176.695 99.770 176.985 ;
        RECT 100.465 176.955 101.965 177.125 ;
        RECT 100.465 176.815 100.635 176.955 ;
        RECT 100.075 176.645 100.635 176.815 ;
        RECT 98.550 176.015 98.800 176.475 ;
        RECT 98.970 176.185 99.840 176.525 ;
        RECT 100.075 176.185 100.245 176.645 ;
        RECT 101.080 176.615 102.155 176.785 ;
        RECT 100.415 176.015 100.785 176.475 ;
        RECT 101.080 176.275 101.250 176.615 ;
        RECT 101.420 176.015 101.750 176.445 ;
        RECT 101.985 176.275 102.155 176.615 ;
        RECT 102.325 176.515 102.495 177.295 ;
        RECT 102.665 177.075 102.835 177.665 ;
        RECT 103.005 177.265 103.355 177.885 ;
        RECT 102.665 176.685 103.130 177.075 ;
        RECT 103.525 176.815 103.695 178.175 ;
        RECT 103.865 176.985 104.325 178.035 ;
        RECT 103.300 176.645 103.695 176.815 ;
        RECT 103.300 176.515 103.470 176.645 ;
        RECT 102.325 176.185 103.005 176.515 ;
        RECT 103.220 176.185 103.470 176.515 ;
        RECT 103.640 176.015 103.890 176.475 ;
        RECT 104.060 176.200 104.385 176.985 ;
        RECT 104.555 176.185 104.725 178.305 ;
        RECT 104.895 178.185 105.225 178.565 ;
        RECT 105.395 178.015 105.650 178.305 ;
        RECT 104.900 177.845 105.650 178.015 ;
        RECT 104.900 176.855 105.130 177.845 ;
        RECT 105.865 177.745 106.095 178.565 ;
        RECT 106.265 177.765 106.595 178.395 ;
        RECT 105.300 177.025 105.650 177.675 ;
        RECT 105.845 177.325 106.175 177.575 ;
        RECT 106.345 177.165 106.595 177.765 ;
        RECT 106.765 177.745 106.975 178.565 ;
        RECT 107.665 177.795 110.255 178.565 ;
        RECT 104.900 176.685 105.650 176.855 ;
        RECT 104.895 176.015 105.225 176.515 ;
        RECT 105.395 176.185 105.650 176.685 ;
        RECT 105.865 176.015 106.095 177.155 ;
        RECT 106.265 176.185 106.595 177.165 ;
        RECT 106.765 176.015 106.975 177.155 ;
        RECT 107.665 177.105 108.875 177.625 ;
        RECT 109.045 177.275 110.255 177.795 ;
        RECT 110.700 177.755 110.945 178.360 ;
        RECT 111.165 178.030 111.675 178.565 ;
        RECT 110.425 177.585 111.655 177.755 ;
        RECT 107.665 176.015 110.255 177.105 ;
        RECT 110.425 176.775 110.765 177.585 ;
        RECT 110.935 177.020 111.685 177.210 ;
        RECT 110.425 176.365 110.940 176.775 ;
        RECT 111.175 176.015 111.345 176.775 ;
        RECT 111.515 176.355 111.685 177.020 ;
        RECT 111.855 177.035 112.045 178.395 ;
        RECT 112.215 178.225 112.490 178.395 ;
        RECT 112.215 178.055 112.495 178.225 ;
        RECT 112.215 177.235 112.490 178.055 ;
        RECT 112.680 178.030 113.210 178.395 ;
        RECT 113.635 178.165 113.965 178.565 ;
        RECT 113.035 177.995 113.210 178.030 ;
        RECT 112.695 177.035 112.865 177.835 ;
        RECT 111.855 176.865 112.865 177.035 ;
        RECT 113.035 177.825 113.965 177.995 ;
        RECT 114.135 177.825 114.390 178.395 ;
        RECT 114.565 177.840 114.855 178.565 ;
        RECT 113.035 176.695 113.205 177.825 ;
        RECT 113.795 177.655 113.965 177.825 ;
        RECT 112.080 176.525 113.205 176.695 ;
        RECT 113.375 177.325 113.570 177.655 ;
        RECT 113.795 177.325 114.050 177.655 ;
        RECT 113.375 176.355 113.545 177.325 ;
        RECT 114.220 177.155 114.390 177.825 ;
        RECT 115.065 177.745 115.295 178.565 ;
        RECT 115.465 177.765 115.795 178.395 ;
        RECT 115.045 177.325 115.375 177.575 ;
        RECT 111.515 176.185 113.545 176.355 ;
        RECT 113.715 176.015 113.885 177.155 ;
        RECT 114.055 176.185 114.390 177.155 ;
        RECT 114.565 176.015 114.855 177.180 ;
        RECT 115.545 177.165 115.795 177.765 ;
        RECT 115.965 177.745 116.175 178.565 ;
        RECT 116.410 177.855 116.665 178.385 ;
        RECT 116.835 178.105 117.140 178.565 ;
        RECT 117.385 178.185 118.455 178.355 ;
        RECT 115.065 176.015 115.295 177.155 ;
        RECT 115.465 176.185 115.795 177.165 ;
        RECT 116.410 177.205 116.620 177.855 ;
        RECT 117.385 177.830 117.705 178.185 ;
        RECT 117.380 177.655 117.705 177.830 ;
        RECT 116.790 177.355 117.705 177.655 ;
        RECT 117.875 177.615 118.115 178.015 ;
        RECT 118.285 177.955 118.455 178.185 ;
        RECT 118.625 178.125 118.815 178.565 ;
        RECT 118.985 178.115 119.935 178.395 ;
        RECT 120.155 178.205 120.505 178.375 ;
        RECT 118.285 177.785 118.815 177.955 ;
        RECT 116.790 177.325 117.530 177.355 ;
        RECT 115.965 176.015 116.175 177.155 ;
        RECT 116.410 176.325 116.665 177.205 ;
        RECT 116.835 176.015 117.140 177.155 ;
        RECT 117.360 176.735 117.530 177.325 ;
        RECT 117.875 177.245 118.415 177.615 ;
        RECT 118.595 177.505 118.815 177.785 ;
        RECT 118.985 177.335 119.155 178.115 ;
        RECT 118.750 177.165 119.155 177.335 ;
        RECT 119.325 177.325 119.675 177.945 ;
        RECT 118.750 177.075 118.920 177.165 ;
        RECT 119.845 177.155 120.055 177.945 ;
        RECT 117.700 176.905 118.920 177.075 ;
        RECT 119.380 176.995 120.055 177.155 ;
        RECT 117.360 176.565 118.160 176.735 ;
        RECT 117.480 176.015 117.810 176.395 ;
        RECT 117.990 176.275 118.160 176.565 ;
        RECT 118.750 176.525 118.920 176.905 ;
        RECT 119.090 176.985 120.055 176.995 ;
        RECT 120.245 177.815 120.505 178.205 ;
        RECT 120.715 178.105 121.045 178.565 ;
        RECT 121.920 178.175 122.775 178.345 ;
        RECT 122.980 178.175 123.475 178.345 ;
        RECT 123.645 178.205 123.975 178.565 ;
        RECT 120.245 177.125 120.415 177.815 ;
        RECT 120.585 177.465 120.755 177.645 ;
        RECT 120.925 177.635 121.715 177.885 ;
        RECT 121.920 177.465 122.090 178.175 ;
        RECT 122.260 177.665 122.615 177.885 ;
        RECT 120.585 177.295 122.275 177.465 ;
        RECT 119.090 176.695 119.550 176.985 ;
        RECT 120.245 176.955 121.745 177.125 ;
        RECT 120.245 176.815 120.415 176.955 ;
        RECT 119.855 176.645 120.415 176.815 ;
        RECT 118.330 176.015 118.580 176.475 ;
        RECT 118.750 176.185 119.620 176.525 ;
        RECT 119.855 176.185 120.025 176.645 ;
        RECT 120.860 176.615 121.935 176.785 ;
        RECT 120.195 176.015 120.565 176.475 ;
        RECT 120.860 176.275 121.030 176.615 ;
        RECT 121.200 176.015 121.530 176.445 ;
        RECT 121.765 176.275 121.935 176.615 ;
        RECT 122.105 176.515 122.275 177.295 ;
        RECT 122.445 177.075 122.615 177.665 ;
        RECT 122.785 177.265 123.135 177.885 ;
        RECT 122.445 176.685 122.910 177.075 ;
        RECT 123.305 176.815 123.475 178.175 ;
        RECT 123.645 176.985 124.105 178.035 ;
        RECT 123.080 176.645 123.475 176.815 ;
        RECT 123.080 176.515 123.250 176.645 ;
        RECT 122.105 176.185 122.785 176.515 ;
        RECT 123.000 176.185 123.250 176.515 ;
        RECT 123.420 176.015 123.670 176.475 ;
        RECT 123.840 176.200 124.165 176.985 ;
        RECT 124.335 176.185 124.505 178.305 ;
        RECT 124.675 178.185 125.005 178.565 ;
        RECT 125.175 178.015 125.430 178.305 ;
        RECT 124.680 177.845 125.430 178.015 ;
        RECT 124.680 176.855 124.910 177.845 ;
        RECT 126.525 177.815 127.735 178.565 ;
        RECT 125.080 177.025 125.430 177.675 ;
        RECT 126.525 177.105 127.045 177.645 ;
        RECT 127.215 177.275 127.735 177.815 ;
        RECT 124.680 176.685 125.430 176.855 ;
        RECT 124.675 176.015 125.005 176.515 ;
        RECT 125.175 176.185 125.430 176.685 ;
        RECT 126.525 176.015 127.735 177.105 ;
        RECT 29.840 175.845 127.820 176.015 ;
        RECT 29.925 174.755 31.135 175.845 ;
        RECT 29.925 174.045 30.445 174.585 ;
        RECT 30.615 174.215 31.135 174.755 ;
        RECT 31.680 174.865 31.935 175.535 ;
        RECT 32.115 175.045 32.400 175.845 ;
        RECT 32.580 175.125 32.910 175.635 ;
        RECT 29.925 173.295 31.135 174.045 ;
        RECT 31.680 174.005 31.860 174.865 ;
        RECT 32.580 174.535 32.830 175.125 ;
        RECT 33.180 174.975 33.350 175.585 ;
        RECT 33.520 175.155 33.850 175.845 ;
        RECT 34.080 175.295 34.320 175.585 ;
        RECT 34.520 175.465 34.940 175.845 ;
        RECT 35.120 175.375 35.750 175.625 ;
        RECT 36.220 175.465 36.550 175.845 ;
        RECT 35.120 175.295 35.290 175.375 ;
        RECT 36.720 175.295 36.890 175.585 ;
        RECT 37.070 175.465 37.450 175.845 ;
        RECT 37.690 175.460 38.520 175.630 ;
        RECT 34.080 175.125 35.290 175.295 ;
        RECT 32.030 174.205 32.830 174.535 ;
        RECT 31.680 173.805 31.935 174.005 ;
        RECT 31.595 173.635 31.935 173.805 ;
        RECT 31.680 173.475 31.935 173.635 ;
        RECT 32.115 173.295 32.400 173.755 ;
        RECT 32.580 173.555 32.830 174.205 ;
        RECT 33.030 174.955 33.350 174.975 ;
        RECT 33.030 174.785 34.950 174.955 ;
        RECT 33.030 173.890 33.220 174.785 ;
        RECT 35.120 174.615 35.290 175.125 ;
        RECT 35.460 174.865 35.980 175.175 ;
        RECT 33.390 174.445 35.290 174.615 ;
        RECT 33.390 174.385 33.720 174.445 ;
        RECT 33.870 174.215 34.200 174.275 ;
        RECT 33.540 173.945 34.200 174.215 ;
        RECT 33.030 173.560 33.350 173.890 ;
        RECT 33.530 173.295 34.190 173.775 ;
        RECT 34.390 173.685 34.560 174.445 ;
        RECT 35.460 174.275 35.640 174.685 ;
        RECT 34.730 174.105 35.060 174.225 ;
        RECT 35.810 174.105 35.980 174.865 ;
        RECT 34.730 173.935 35.980 174.105 ;
        RECT 36.150 175.045 37.520 175.295 ;
        RECT 36.150 174.275 36.340 175.045 ;
        RECT 37.270 174.785 37.520 175.045 ;
        RECT 36.510 174.615 36.760 174.775 ;
        RECT 37.690 174.615 37.860 175.460 ;
        RECT 38.755 175.175 38.925 175.675 ;
        RECT 39.095 175.345 39.425 175.845 ;
        RECT 38.030 174.785 38.530 175.165 ;
        RECT 38.755 175.005 39.450 175.175 ;
        RECT 36.510 174.445 37.860 174.615 ;
        RECT 37.440 174.405 37.860 174.445 ;
        RECT 36.150 173.935 36.570 174.275 ;
        RECT 36.860 173.945 37.270 174.275 ;
        RECT 34.390 173.515 35.240 173.685 ;
        RECT 35.800 173.295 36.120 173.755 ;
        RECT 36.320 173.505 36.570 173.935 ;
        RECT 36.860 173.295 37.270 173.735 ;
        RECT 37.440 173.675 37.610 174.405 ;
        RECT 37.780 173.855 38.130 174.225 ;
        RECT 38.310 173.915 38.530 174.785 ;
        RECT 38.700 174.215 39.110 174.835 ;
        RECT 39.280 174.035 39.450 175.005 ;
        RECT 38.755 173.845 39.450 174.035 ;
        RECT 37.440 173.475 38.455 173.675 ;
        RECT 38.755 173.515 38.925 173.845 ;
        RECT 39.095 173.295 39.425 173.675 ;
        RECT 39.640 173.555 39.865 175.675 ;
        RECT 40.035 175.345 40.365 175.845 ;
        RECT 40.535 175.175 40.705 175.675 ;
        RECT 40.040 175.005 40.705 175.175 ;
        RECT 40.040 174.015 40.270 175.005 ;
        RECT 40.440 174.185 40.790 174.835 ;
        RECT 41.425 174.705 41.810 175.675 ;
        RECT 41.980 175.385 42.305 175.845 ;
        RECT 42.825 175.215 43.105 175.675 ;
        RECT 41.980 174.995 43.105 175.215 ;
        RECT 41.425 174.035 41.705 174.705 ;
        RECT 41.980 174.535 42.430 174.995 ;
        RECT 43.295 174.825 43.695 175.675 ;
        RECT 44.095 175.385 44.365 175.845 ;
        RECT 44.535 175.215 44.820 175.675 ;
        RECT 41.875 174.205 42.430 174.535 ;
        RECT 42.600 174.265 43.695 174.825 ;
        RECT 41.980 174.095 42.430 174.205 ;
        RECT 40.040 173.845 40.705 174.015 ;
        RECT 40.035 173.295 40.365 173.675 ;
        RECT 40.535 173.555 40.705 173.845 ;
        RECT 41.425 173.465 41.810 174.035 ;
        RECT 41.980 173.925 43.105 174.095 ;
        RECT 41.980 173.295 42.305 173.755 ;
        RECT 42.825 173.465 43.105 173.925 ;
        RECT 43.295 173.465 43.695 174.265 ;
        RECT 43.865 174.995 44.820 175.215 ;
        RECT 43.865 174.095 44.075 174.995 ;
        RECT 44.245 174.265 44.935 174.825 ;
        RECT 45.105 174.705 45.490 175.675 ;
        RECT 45.660 175.385 45.985 175.845 ;
        RECT 46.505 175.215 46.785 175.675 ;
        RECT 45.660 174.995 46.785 175.215 ;
        RECT 43.865 173.925 44.820 174.095 ;
        RECT 44.095 173.295 44.365 173.755 ;
        RECT 44.535 173.465 44.820 173.925 ;
        RECT 45.105 174.035 45.385 174.705 ;
        RECT 45.660 174.535 46.110 174.995 ;
        RECT 46.975 174.825 47.375 175.675 ;
        RECT 47.775 175.385 48.045 175.845 ;
        RECT 48.215 175.215 48.500 175.675 ;
        RECT 45.555 174.205 46.110 174.535 ;
        RECT 46.280 174.265 47.375 174.825 ;
        RECT 45.660 174.095 46.110 174.205 ;
        RECT 45.105 173.465 45.490 174.035 ;
        RECT 45.660 173.925 46.785 174.095 ;
        RECT 45.660 173.295 45.985 173.755 ;
        RECT 46.505 173.465 46.785 173.925 ;
        RECT 46.975 173.465 47.375 174.265 ;
        RECT 47.545 174.995 48.500 175.215 ;
        RECT 47.545 174.095 47.755 174.995 ;
        RECT 47.925 174.265 48.615 174.825 ;
        RECT 48.825 174.705 49.055 175.845 ;
        RECT 49.225 174.695 49.555 175.675 ;
        RECT 49.725 174.705 49.935 175.845 ;
        RECT 48.805 174.285 49.135 174.535 ;
        RECT 47.545 173.925 48.500 174.095 ;
        RECT 47.775 173.295 48.045 173.755 ;
        RECT 48.215 173.465 48.500 173.925 ;
        RECT 48.825 173.295 49.055 174.115 ;
        RECT 49.305 174.095 49.555 174.695 ;
        RECT 50.165 174.680 50.455 175.845 ;
        RECT 50.625 174.755 52.295 175.845 ;
        RECT 50.625 174.235 51.375 174.755 ;
        RECT 52.505 174.705 52.735 175.845 ;
        RECT 52.905 174.695 53.235 175.675 ;
        RECT 53.405 174.705 53.615 175.845 ;
        RECT 49.225 173.465 49.555 174.095 ;
        RECT 49.725 173.295 49.935 174.115 ;
        RECT 51.545 174.065 52.295 174.585 ;
        RECT 52.485 174.285 52.815 174.535 ;
        RECT 50.165 173.295 50.455 174.020 ;
        RECT 50.625 173.295 52.295 174.065 ;
        RECT 52.505 173.295 52.735 174.115 ;
        RECT 52.985 174.095 53.235 174.695 ;
        RECT 53.850 174.655 54.105 175.535 ;
        RECT 54.275 174.705 54.580 175.845 ;
        RECT 54.920 175.465 55.250 175.845 ;
        RECT 55.430 175.295 55.600 175.585 ;
        RECT 55.770 175.385 56.020 175.845 ;
        RECT 54.800 175.125 55.600 175.295 ;
        RECT 56.190 175.335 57.060 175.675 ;
        RECT 52.905 173.465 53.235 174.095 ;
        RECT 53.405 173.295 53.615 174.115 ;
        RECT 53.850 174.005 54.060 174.655 ;
        RECT 54.800 174.535 54.970 175.125 ;
        RECT 56.190 174.955 56.360 175.335 ;
        RECT 57.295 175.215 57.465 175.675 ;
        RECT 57.635 175.385 58.005 175.845 ;
        RECT 58.300 175.245 58.470 175.585 ;
        RECT 58.640 175.415 58.970 175.845 ;
        RECT 59.205 175.245 59.375 175.585 ;
        RECT 55.140 174.785 56.360 174.955 ;
        RECT 56.530 174.875 56.990 175.165 ;
        RECT 57.295 175.045 57.855 175.215 ;
        RECT 58.300 175.075 59.375 175.245 ;
        RECT 59.545 175.345 60.225 175.675 ;
        RECT 60.440 175.345 60.690 175.675 ;
        RECT 60.860 175.385 61.110 175.845 ;
        RECT 57.685 174.905 57.855 175.045 ;
        RECT 56.530 174.865 57.495 174.875 ;
        RECT 56.190 174.695 56.360 174.785 ;
        RECT 56.820 174.705 57.495 174.865 ;
        RECT 54.230 174.505 54.970 174.535 ;
        RECT 54.230 174.205 55.145 174.505 ;
        RECT 54.820 174.030 55.145 174.205 ;
        RECT 53.850 173.475 54.105 174.005 ;
        RECT 54.275 173.295 54.580 173.755 ;
        RECT 54.825 173.675 55.145 174.030 ;
        RECT 55.315 174.245 55.855 174.615 ;
        RECT 56.190 174.525 56.595 174.695 ;
        RECT 55.315 173.845 55.555 174.245 ;
        RECT 56.035 174.075 56.255 174.355 ;
        RECT 55.725 173.905 56.255 174.075 ;
        RECT 55.725 173.675 55.895 173.905 ;
        RECT 56.425 173.745 56.595 174.525 ;
        RECT 56.765 173.915 57.115 174.535 ;
        RECT 57.285 173.915 57.495 174.705 ;
        RECT 57.685 174.735 59.185 174.905 ;
        RECT 57.685 174.045 57.855 174.735 ;
        RECT 59.545 174.565 59.715 175.345 ;
        RECT 60.520 175.215 60.690 175.345 ;
        RECT 58.025 174.395 59.715 174.565 ;
        RECT 59.885 174.785 60.350 175.175 ;
        RECT 60.520 175.045 60.915 175.215 ;
        RECT 58.025 174.215 58.195 174.395 ;
        RECT 54.825 173.505 55.895 173.675 ;
        RECT 56.065 173.295 56.255 173.735 ;
        RECT 56.425 173.465 57.375 173.745 ;
        RECT 57.685 173.655 57.945 174.045 ;
        RECT 58.365 173.975 59.155 174.225 ;
        RECT 57.595 173.485 57.945 173.655 ;
        RECT 58.155 173.295 58.485 173.755 ;
        RECT 59.360 173.685 59.530 174.395 ;
        RECT 59.885 174.195 60.055 174.785 ;
        RECT 59.700 173.975 60.055 174.195 ;
        RECT 60.225 173.975 60.575 174.595 ;
        RECT 60.745 173.685 60.915 175.045 ;
        RECT 61.280 174.875 61.605 175.660 ;
        RECT 61.085 173.825 61.545 174.875 ;
        RECT 59.360 173.515 60.215 173.685 ;
        RECT 60.420 173.515 60.915 173.685 ;
        RECT 61.085 173.295 61.415 173.655 ;
        RECT 61.775 173.555 61.945 175.675 ;
        RECT 62.115 175.345 62.445 175.845 ;
        RECT 62.615 175.175 62.870 175.675 ;
        RECT 62.120 175.005 62.870 175.175 ;
        RECT 62.120 174.015 62.350 175.005 ;
        RECT 62.520 174.185 62.870 174.835 ;
        RECT 63.050 174.705 63.385 175.675 ;
        RECT 63.555 174.705 63.725 175.845 ;
        RECT 63.895 175.505 65.925 175.675 ;
        RECT 63.050 174.035 63.220 174.705 ;
        RECT 63.895 174.535 64.065 175.505 ;
        RECT 63.390 174.205 63.645 174.535 ;
        RECT 63.870 174.205 64.065 174.535 ;
        RECT 64.235 175.165 65.360 175.335 ;
        RECT 63.475 174.035 63.645 174.205 ;
        RECT 64.235 174.035 64.405 175.165 ;
        RECT 62.120 173.845 62.870 174.015 ;
        RECT 62.115 173.295 62.445 173.675 ;
        RECT 62.615 173.555 62.870 173.845 ;
        RECT 63.050 173.465 63.305 174.035 ;
        RECT 63.475 173.865 64.405 174.035 ;
        RECT 64.575 174.825 65.585 174.995 ;
        RECT 64.575 174.025 64.745 174.825 ;
        RECT 64.950 174.485 65.225 174.625 ;
        RECT 64.945 174.315 65.225 174.485 ;
        RECT 64.230 173.830 64.405 173.865 ;
        RECT 63.475 173.295 63.805 173.695 ;
        RECT 64.230 173.465 64.760 173.830 ;
        RECT 64.950 173.465 65.225 174.315 ;
        RECT 65.395 173.465 65.585 174.825 ;
        RECT 65.755 174.840 65.925 175.505 ;
        RECT 66.095 175.085 66.265 175.845 ;
        RECT 66.500 175.085 67.015 175.495 ;
        RECT 65.755 174.650 66.505 174.840 ;
        RECT 66.675 174.275 67.015 175.085 ;
        RECT 65.785 174.105 67.015 174.275 ;
        RECT 67.185 174.755 69.775 175.845 ;
        RECT 67.185 174.235 68.395 174.755 ;
        RECT 70.005 174.705 70.215 175.845 ;
        RECT 70.385 174.695 70.715 175.675 ;
        RECT 70.885 174.705 71.115 175.845 ;
        RECT 71.415 174.915 71.585 175.675 ;
        RECT 71.765 175.085 72.095 175.845 ;
        RECT 71.415 174.745 72.080 174.915 ;
        RECT 72.265 174.770 72.535 175.675 ;
        RECT 65.765 173.295 66.275 173.830 ;
        RECT 66.495 173.500 66.740 174.105 ;
        RECT 68.565 174.065 69.775 174.585 ;
        RECT 67.185 173.295 69.775 174.065 ;
        RECT 70.005 173.295 70.215 174.115 ;
        RECT 70.385 174.095 70.635 174.695 ;
        RECT 71.910 174.600 72.080 174.745 ;
        RECT 70.805 174.285 71.135 174.535 ;
        RECT 71.345 174.195 71.675 174.565 ;
        RECT 71.910 174.270 72.195 174.600 ;
        RECT 70.385 173.465 70.715 174.095 ;
        RECT 70.885 173.295 71.115 174.115 ;
        RECT 71.910 174.015 72.080 174.270 ;
        RECT 71.415 173.845 72.080 174.015 ;
        RECT 72.365 173.970 72.535 174.770 ;
        RECT 73.315 174.695 73.645 175.845 ;
        RECT 73.815 174.825 73.985 175.675 ;
        RECT 74.155 175.045 74.485 175.845 ;
        RECT 74.655 174.825 74.825 175.675 ;
        RECT 75.005 175.045 75.245 175.845 ;
        RECT 75.415 174.865 75.745 175.675 ;
        RECT 73.815 174.655 74.825 174.825 ;
        RECT 75.030 174.695 75.745 174.865 ;
        RECT 73.815 174.115 74.310 174.655 ;
        RECT 75.030 174.455 75.200 174.695 ;
        RECT 75.925 174.680 76.215 175.845 ;
        RECT 76.995 174.695 77.325 175.845 ;
        RECT 77.495 174.825 77.665 175.675 ;
        RECT 77.835 175.045 78.165 175.845 ;
        RECT 78.335 174.825 78.505 175.675 ;
        RECT 78.685 175.045 78.925 175.845 ;
        RECT 79.095 174.865 79.425 175.675 ;
        RECT 77.495 174.655 78.505 174.825 ;
        RECT 78.710 174.695 79.425 174.865 ;
        RECT 80.525 174.875 80.835 175.675 ;
        RECT 81.005 175.045 81.315 175.845 ;
        RECT 81.485 175.215 81.745 175.675 ;
        RECT 81.915 175.385 82.170 175.845 ;
        RECT 82.345 175.215 82.605 175.675 ;
        RECT 81.485 175.045 82.605 175.215 ;
        RECT 80.525 174.705 81.555 174.875 ;
        RECT 74.700 174.285 75.200 174.455 ;
        RECT 75.370 174.285 75.750 174.525 ;
        RECT 75.030 174.115 75.200 174.285 ;
        RECT 77.495 174.115 77.990 174.655 ;
        RECT 78.710 174.455 78.880 174.695 ;
        RECT 78.380 174.285 78.880 174.455 ;
        RECT 79.050 174.285 79.430 174.525 ;
        RECT 78.710 174.115 78.880 174.285 ;
        RECT 71.415 173.465 71.585 173.845 ;
        RECT 71.765 173.295 72.095 173.675 ;
        RECT 72.275 173.465 72.535 173.970 ;
        RECT 73.315 173.295 73.645 174.095 ;
        RECT 73.815 173.945 74.825 174.115 ;
        RECT 75.030 173.945 75.665 174.115 ;
        RECT 73.815 173.465 73.985 173.945 ;
        RECT 74.155 173.295 74.485 173.775 ;
        RECT 74.655 173.465 74.825 173.945 ;
        RECT 75.075 173.295 75.315 173.775 ;
        RECT 75.495 173.465 75.665 173.945 ;
        RECT 75.925 173.295 76.215 174.020 ;
        RECT 76.995 173.295 77.325 174.095 ;
        RECT 77.495 173.945 78.505 174.115 ;
        RECT 78.710 173.945 79.345 174.115 ;
        RECT 77.495 173.465 77.665 173.945 ;
        RECT 77.835 173.295 78.165 173.775 ;
        RECT 78.335 173.465 78.505 173.945 ;
        RECT 78.755 173.295 78.995 173.775 ;
        RECT 79.175 173.465 79.345 173.945 ;
        RECT 80.525 173.795 80.695 174.705 ;
        RECT 80.865 173.965 81.215 174.535 ;
        RECT 81.385 174.455 81.555 174.705 ;
        RECT 82.345 174.795 82.605 175.045 ;
        RECT 82.775 174.975 83.060 175.845 ;
        RECT 82.345 174.625 83.100 174.795 ;
        RECT 81.385 174.285 82.525 174.455 ;
        RECT 82.695 174.115 83.100 174.625 ;
        RECT 83.285 174.755 84.955 175.845 ;
        RECT 85.500 174.865 85.755 175.535 ;
        RECT 85.935 175.045 86.220 175.845 ;
        RECT 86.400 175.125 86.730 175.635 ;
        RECT 83.285 174.235 84.035 174.755 ;
        RECT 81.450 173.945 83.100 174.115 ;
        RECT 84.205 174.065 84.955 174.585 ;
        RECT 80.525 173.465 80.825 173.795 ;
        RECT 80.995 173.295 81.270 173.775 ;
        RECT 81.450 173.555 81.745 173.945 ;
        RECT 81.915 173.295 82.170 173.775 ;
        RECT 82.345 173.555 82.605 173.945 ;
        RECT 82.775 173.295 83.055 173.775 ;
        RECT 83.285 173.295 84.955 174.065 ;
        RECT 85.500 174.005 85.680 174.865 ;
        RECT 86.400 174.535 86.650 175.125 ;
        RECT 87.000 174.975 87.170 175.585 ;
        RECT 87.340 175.155 87.670 175.845 ;
        RECT 87.900 175.295 88.140 175.585 ;
        RECT 88.340 175.465 88.760 175.845 ;
        RECT 88.940 175.375 89.570 175.625 ;
        RECT 90.040 175.465 90.370 175.845 ;
        RECT 88.940 175.295 89.110 175.375 ;
        RECT 90.540 175.295 90.710 175.585 ;
        RECT 90.890 175.465 91.270 175.845 ;
        RECT 91.510 175.460 92.340 175.630 ;
        RECT 87.900 175.125 89.110 175.295 ;
        RECT 85.850 174.205 86.650 174.535 ;
        RECT 85.500 173.805 85.755 174.005 ;
        RECT 85.415 173.635 85.755 173.805 ;
        RECT 85.500 173.475 85.755 173.635 ;
        RECT 85.935 173.295 86.220 173.755 ;
        RECT 86.400 173.555 86.650 174.205 ;
        RECT 86.850 174.955 87.170 174.975 ;
        RECT 86.850 174.785 88.770 174.955 ;
        RECT 86.850 173.890 87.040 174.785 ;
        RECT 88.940 174.615 89.110 175.125 ;
        RECT 89.280 174.865 89.800 175.175 ;
        RECT 87.210 174.445 89.110 174.615 ;
        RECT 87.210 174.385 87.540 174.445 ;
        RECT 87.690 174.215 88.020 174.275 ;
        RECT 87.360 173.945 88.020 174.215 ;
        RECT 86.850 173.560 87.170 173.890 ;
        RECT 87.350 173.295 88.010 173.775 ;
        RECT 88.210 173.685 88.380 174.445 ;
        RECT 89.280 174.275 89.460 174.685 ;
        RECT 88.550 174.105 88.880 174.225 ;
        RECT 89.630 174.105 89.800 174.865 ;
        RECT 88.550 173.935 89.800 174.105 ;
        RECT 89.970 175.045 91.340 175.295 ;
        RECT 89.970 174.275 90.160 175.045 ;
        RECT 91.090 174.785 91.340 175.045 ;
        RECT 90.330 174.615 90.580 174.775 ;
        RECT 91.510 174.615 91.680 175.460 ;
        RECT 92.575 175.175 92.745 175.675 ;
        RECT 92.915 175.345 93.245 175.845 ;
        RECT 91.850 174.785 92.350 175.165 ;
        RECT 92.575 175.005 93.270 175.175 ;
        RECT 90.330 174.445 91.680 174.615 ;
        RECT 91.260 174.405 91.680 174.445 ;
        RECT 89.970 173.935 90.390 174.275 ;
        RECT 90.680 173.945 91.090 174.275 ;
        RECT 88.210 173.515 89.060 173.685 ;
        RECT 89.620 173.295 89.940 173.755 ;
        RECT 90.140 173.505 90.390 173.935 ;
        RECT 90.680 173.295 91.090 173.735 ;
        RECT 91.260 173.675 91.430 174.405 ;
        RECT 91.600 173.855 91.950 174.225 ;
        RECT 92.130 173.915 92.350 174.785 ;
        RECT 92.520 174.215 92.930 174.835 ;
        RECT 93.100 174.035 93.270 175.005 ;
        RECT 92.575 173.845 93.270 174.035 ;
        RECT 91.260 173.475 92.275 173.675 ;
        RECT 92.575 173.515 92.745 173.845 ;
        RECT 92.915 173.295 93.245 173.675 ;
        RECT 93.460 173.555 93.685 175.675 ;
        RECT 93.855 175.345 94.185 175.845 ;
        RECT 94.355 175.175 94.525 175.675 ;
        RECT 93.860 175.005 94.525 175.175 ;
        RECT 93.860 174.015 94.090 175.005 ;
        RECT 94.260 174.185 94.610 174.835 ;
        RECT 95.745 174.705 95.975 175.845 ;
        RECT 96.145 174.695 96.475 175.675 ;
        RECT 96.645 174.705 96.855 175.845 ;
        RECT 97.085 175.085 97.600 175.495 ;
        RECT 97.835 175.085 98.005 175.845 ;
        RECT 98.175 175.505 100.205 175.675 ;
        RECT 95.725 174.285 96.055 174.535 ;
        RECT 93.860 173.845 94.525 174.015 ;
        RECT 93.855 173.295 94.185 173.675 ;
        RECT 94.355 173.555 94.525 173.845 ;
        RECT 95.745 173.295 95.975 174.115 ;
        RECT 96.225 174.095 96.475 174.695 ;
        RECT 97.085 174.275 97.425 175.085 ;
        RECT 98.175 174.840 98.345 175.505 ;
        RECT 98.740 175.165 99.865 175.335 ;
        RECT 97.595 174.650 98.345 174.840 ;
        RECT 98.515 174.825 99.525 174.995 ;
        RECT 96.145 173.465 96.475 174.095 ;
        RECT 96.645 173.295 96.855 174.115 ;
        RECT 97.085 174.105 98.315 174.275 ;
        RECT 97.360 173.500 97.605 174.105 ;
        RECT 97.825 173.295 98.335 173.830 ;
        RECT 98.515 173.465 98.705 174.825 ;
        RECT 98.875 174.485 99.150 174.625 ;
        RECT 98.875 174.315 99.155 174.485 ;
        RECT 98.875 173.465 99.150 174.315 ;
        RECT 99.355 174.025 99.525 174.825 ;
        RECT 99.695 174.035 99.865 175.165 ;
        RECT 100.035 174.535 100.205 175.505 ;
        RECT 100.375 174.705 100.545 175.845 ;
        RECT 100.715 174.705 101.050 175.675 ;
        RECT 100.035 174.205 100.230 174.535 ;
        RECT 100.455 174.205 100.710 174.535 ;
        RECT 100.455 174.035 100.625 174.205 ;
        RECT 100.880 174.035 101.050 174.705 ;
        RECT 101.685 174.680 101.975 175.845 ;
        RECT 102.245 175.385 102.415 175.845 ;
        RECT 102.585 174.895 102.915 175.675 ;
        RECT 103.085 175.045 103.255 175.845 ;
        RECT 102.145 174.875 102.915 174.895 ;
        RECT 103.425 174.875 103.755 175.675 ;
        RECT 103.925 175.045 104.095 175.845 ;
        RECT 104.265 174.875 104.595 175.675 ;
        RECT 102.145 174.705 104.595 174.875 ;
        RECT 104.855 174.705 105.150 175.845 ;
        RECT 99.695 173.865 100.625 174.035 ;
        RECT 99.695 173.830 99.870 173.865 ;
        RECT 99.340 173.465 99.870 173.830 ;
        RECT 100.295 173.295 100.625 173.695 ;
        RECT 100.795 173.465 101.050 174.035 ;
        RECT 102.145 174.115 102.495 174.705 ;
        RECT 106.290 174.655 106.545 175.535 ;
        RECT 106.715 174.705 107.020 175.845 ;
        RECT 107.360 175.465 107.690 175.845 ;
        RECT 107.870 175.295 108.040 175.585 ;
        RECT 108.210 175.385 108.460 175.845 ;
        RECT 107.240 175.125 108.040 175.295 ;
        RECT 108.630 175.335 109.500 175.675 ;
        RECT 102.665 174.285 105.175 174.535 ;
        RECT 101.685 173.295 101.975 174.020 ;
        RECT 102.145 173.935 104.515 174.115 ;
        RECT 102.245 173.295 102.495 173.760 ;
        RECT 102.665 173.465 102.835 173.935 ;
        RECT 103.085 173.295 103.255 173.755 ;
        RECT 103.505 173.465 103.675 173.935 ;
        RECT 103.925 173.295 104.095 173.755 ;
        RECT 104.345 173.465 104.515 173.935 ;
        RECT 106.290 174.005 106.500 174.655 ;
        RECT 107.240 174.535 107.410 175.125 ;
        RECT 108.630 174.955 108.800 175.335 ;
        RECT 109.735 175.215 109.905 175.675 ;
        RECT 110.075 175.385 110.445 175.845 ;
        RECT 110.740 175.245 110.910 175.585 ;
        RECT 111.080 175.415 111.410 175.845 ;
        RECT 111.645 175.245 111.815 175.585 ;
        RECT 107.580 174.785 108.800 174.955 ;
        RECT 108.970 174.875 109.430 175.165 ;
        RECT 109.735 175.045 110.295 175.215 ;
        RECT 110.740 175.075 111.815 175.245 ;
        RECT 111.985 175.345 112.665 175.675 ;
        RECT 112.880 175.345 113.130 175.675 ;
        RECT 113.300 175.385 113.550 175.845 ;
        RECT 110.125 174.905 110.295 175.045 ;
        RECT 108.970 174.865 109.935 174.875 ;
        RECT 108.630 174.695 108.800 174.785 ;
        RECT 109.260 174.705 109.935 174.865 ;
        RECT 106.670 174.505 107.410 174.535 ;
        RECT 106.670 174.205 107.585 174.505 ;
        RECT 107.260 174.030 107.585 174.205 ;
        RECT 104.885 173.295 105.150 173.755 ;
        RECT 106.290 173.475 106.545 174.005 ;
        RECT 106.715 173.295 107.020 173.755 ;
        RECT 107.265 173.675 107.585 174.030 ;
        RECT 107.755 174.245 108.295 174.615 ;
        RECT 108.630 174.525 109.035 174.695 ;
        RECT 107.755 173.845 107.995 174.245 ;
        RECT 108.475 174.075 108.695 174.355 ;
        RECT 108.165 173.905 108.695 174.075 ;
        RECT 108.165 173.675 108.335 173.905 ;
        RECT 108.865 173.745 109.035 174.525 ;
        RECT 109.205 173.915 109.555 174.535 ;
        RECT 109.725 173.915 109.935 174.705 ;
        RECT 110.125 174.735 111.625 174.905 ;
        RECT 110.125 174.045 110.295 174.735 ;
        RECT 111.985 174.565 112.155 175.345 ;
        RECT 112.960 175.215 113.130 175.345 ;
        RECT 110.465 174.395 112.155 174.565 ;
        RECT 112.325 174.785 112.790 175.175 ;
        RECT 112.960 175.045 113.355 175.215 ;
        RECT 110.465 174.215 110.635 174.395 ;
        RECT 107.265 173.505 108.335 173.675 ;
        RECT 108.505 173.295 108.695 173.735 ;
        RECT 108.865 173.465 109.815 173.745 ;
        RECT 110.125 173.655 110.385 174.045 ;
        RECT 110.805 173.975 111.595 174.225 ;
        RECT 110.035 173.485 110.385 173.655 ;
        RECT 110.595 173.295 110.925 173.755 ;
        RECT 111.800 173.685 111.970 174.395 ;
        RECT 112.325 174.195 112.495 174.785 ;
        RECT 112.140 173.975 112.495 174.195 ;
        RECT 112.665 173.975 113.015 174.595 ;
        RECT 113.185 173.685 113.355 175.045 ;
        RECT 113.720 174.875 114.045 175.660 ;
        RECT 113.525 173.825 113.985 174.875 ;
        RECT 111.800 173.515 112.655 173.685 ;
        RECT 112.860 173.515 113.355 173.685 ;
        RECT 113.525 173.295 113.855 173.655 ;
        RECT 114.215 173.555 114.385 175.675 ;
        RECT 114.555 175.345 114.885 175.845 ;
        RECT 115.055 175.175 115.310 175.675 ;
        RECT 114.560 175.005 115.310 175.175 ;
        RECT 115.945 175.085 116.460 175.495 ;
        RECT 116.695 175.085 116.865 175.845 ;
        RECT 117.035 175.505 119.065 175.675 ;
        RECT 114.560 174.015 114.790 175.005 ;
        RECT 114.960 174.185 115.310 174.835 ;
        RECT 115.945 174.275 116.285 175.085 ;
        RECT 117.035 174.840 117.205 175.505 ;
        RECT 117.600 175.165 118.725 175.335 ;
        RECT 116.455 174.650 117.205 174.840 ;
        RECT 117.375 174.825 118.385 174.995 ;
        RECT 115.945 174.105 117.175 174.275 ;
        RECT 114.560 173.845 115.310 174.015 ;
        RECT 114.555 173.295 114.885 173.675 ;
        RECT 115.055 173.555 115.310 173.845 ;
        RECT 116.220 173.500 116.465 174.105 ;
        RECT 116.685 173.295 117.195 173.830 ;
        RECT 117.375 173.465 117.565 174.825 ;
        RECT 117.735 174.485 118.010 174.625 ;
        RECT 117.735 174.315 118.015 174.485 ;
        RECT 117.735 173.465 118.010 174.315 ;
        RECT 118.215 174.025 118.385 174.825 ;
        RECT 118.555 174.035 118.725 175.165 ;
        RECT 118.895 174.535 119.065 175.505 ;
        RECT 119.235 174.705 119.405 175.845 ;
        RECT 119.575 174.705 119.910 175.675 ;
        RECT 118.895 174.205 119.090 174.535 ;
        RECT 119.315 174.205 119.570 174.535 ;
        RECT 119.315 174.035 119.485 174.205 ;
        RECT 119.740 174.035 119.910 174.705 ;
        RECT 118.555 173.865 119.485 174.035 ;
        RECT 118.555 173.830 118.730 173.865 ;
        RECT 118.200 173.465 118.730 173.830 ;
        RECT 119.155 173.295 119.485 173.695 ;
        RECT 119.655 173.465 119.910 174.035 ;
        RECT 120.085 174.705 120.470 175.675 ;
        RECT 120.640 175.385 120.965 175.845 ;
        RECT 121.485 175.215 121.765 175.675 ;
        RECT 120.640 174.995 121.765 175.215 ;
        RECT 120.085 174.035 120.365 174.705 ;
        RECT 120.640 174.535 121.090 174.995 ;
        RECT 121.955 174.825 122.355 175.675 ;
        RECT 122.755 175.385 123.025 175.845 ;
        RECT 123.195 175.215 123.480 175.675 ;
        RECT 123.770 175.420 124.105 175.845 ;
        RECT 124.275 175.240 124.460 175.645 ;
        RECT 120.535 174.205 121.090 174.535 ;
        RECT 121.260 174.265 122.355 174.825 ;
        RECT 120.640 174.095 121.090 174.205 ;
        RECT 120.085 173.465 120.470 174.035 ;
        RECT 120.640 173.925 121.765 174.095 ;
        RECT 120.640 173.295 120.965 173.755 ;
        RECT 121.485 173.465 121.765 173.925 ;
        RECT 121.955 173.465 122.355 174.265 ;
        RECT 122.525 174.995 123.480 175.215 ;
        RECT 123.795 175.065 124.460 175.240 ;
        RECT 124.665 175.065 124.995 175.845 ;
        RECT 122.525 174.095 122.735 174.995 ;
        RECT 122.905 174.265 123.595 174.825 ;
        RECT 122.525 173.925 123.480 174.095 ;
        RECT 122.755 173.295 123.025 173.755 ;
        RECT 123.195 173.465 123.480 173.925 ;
        RECT 123.795 174.035 124.135 175.065 ;
        RECT 125.165 174.875 125.435 175.645 ;
        RECT 124.305 174.705 125.435 174.875 ;
        RECT 124.305 174.205 124.555 174.705 ;
        RECT 123.795 173.865 124.480 174.035 ;
        RECT 124.735 173.955 125.095 174.535 ;
        RECT 123.770 173.295 124.105 173.695 ;
        RECT 124.275 173.465 124.480 173.865 ;
        RECT 125.265 173.795 125.435 174.705 ;
        RECT 126.525 174.755 127.735 175.845 ;
        RECT 126.525 174.215 127.045 174.755 ;
        RECT 127.215 174.045 127.735 174.585 ;
        RECT 124.690 173.295 124.965 173.775 ;
        RECT 125.175 173.465 125.435 173.795 ;
        RECT 126.525 173.295 127.735 174.045 ;
        RECT 29.840 173.125 127.820 173.295 ;
        RECT 29.925 172.375 31.135 173.125 ;
        RECT 29.925 171.835 30.445 172.375 ;
        RECT 31.305 172.355 34.815 173.125 ;
        RECT 30.615 171.665 31.135 172.205 ;
        RECT 29.925 170.575 31.135 171.665 ;
        RECT 31.305 171.665 32.995 172.185 ;
        RECT 33.165 171.835 34.815 172.355 ;
        RECT 35.045 172.305 35.255 173.125 ;
        RECT 35.425 172.325 35.755 172.955 ;
        RECT 35.425 171.725 35.675 172.325 ;
        RECT 35.925 172.305 36.155 173.125 ;
        RECT 37.285 172.400 37.575 173.125 ;
        RECT 38.665 172.450 38.925 172.955 ;
        RECT 39.105 172.745 39.435 173.125 ;
        RECT 39.615 172.575 39.785 172.955 ;
        RECT 35.845 171.885 36.175 172.135 ;
        RECT 31.305 170.575 34.815 171.665 ;
        RECT 35.045 170.575 35.255 171.715 ;
        RECT 35.425 170.745 35.755 171.725 ;
        RECT 35.925 170.575 36.155 171.715 ;
        RECT 37.285 170.575 37.575 171.740 ;
        RECT 38.665 171.650 38.835 172.450 ;
        RECT 39.120 172.405 39.785 172.575 ;
        RECT 40.045 172.450 40.305 172.955 ;
        RECT 40.485 172.745 40.815 173.125 ;
        RECT 40.995 172.575 41.165 172.955 ;
        RECT 39.120 172.150 39.290 172.405 ;
        RECT 39.005 171.820 39.290 172.150 ;
        RECT 39.525 171.855 39.855 172.225 ;
        RECT 39.120 171.675 39.290 171.820 ;
        RECT 38.665 170.745 38.935 171.650 ;
        RECT 39.120 171.505 39.785 171.675 ;
        RECT 39.105 170.575 39.435 171.335 ;
        RECT 39.615 170.745 39.785 171.505 ;
        RECT 40.045 171.650 40.215 172.450 ;
        RECT 40.500 172.405 41.165 172.575 ;
        RECT 40.500 172.150 40.670 172.405 ;
        RECT 41.430 172.385 41.685 172.955 ;
        RECT 41.855 172.725 42.185 173.125 ;
        RECT 42.610 172.590 43.140 172.955 ;
        RECT 42.610 172.555 42.785 172.590 ;
        RECT 41.855 172.385 42.785 172.555 ;
        RECT 40.385 171.820 40.670 172.150 ;
        RECT 40.905 171.855 41.235 172.225 ;
        RECT 40.500 171.675 40.670 171.820 ;
        RECT 41.430 171.715 41.600 172.385 ;
        RECT 41.855 172.215 42.025 172.385 ;
        RECT 41.770 171.885 42.025 172.215 ;
        RECT 42.250 171.885 42.445 172.215 ;
        RECT 40.045 170.745 40.315 171.650 ;
        RECT 40.500 171.505 41.165 171.675 ;
        RECT 40.485 170.575 40.815 171.335 ;
        RECT 40.995 170.745 41.165 171.505 ;
        RECT 41.430 170.745 41.765 171.715 ;
        RECT 41.935 170.575 42.105 171.715 ;
        RECT 42.275 170.915 42.445 171.885 ;
        RECT 42.615 171.255 42.785 172.385 ;
        RECT 42.955 171.595 43.125 172.395 ;
        RECT 43.330 172.105 43.605 172.955 ;
        RECT 43.325 171.935 43.605 172.105 ;
        RECT 43.330 171.795 43.605 171.935 ;
        RECT 43.775 171.595 43.965 172.955 ;
        RECT 44.145 172.590 44.655 173.125 ;
        RECT 44.875 172.315 45.120 172.920 ;
        RECT 46.140 172.495 46.425 172.955 ;
        RECT 46.595 172.665 46.865 173.125 ;
        RECT 46.140 172.325 47.095 172.495 ;
        RECT 44.165 172.145 45.395 172.315 ;
        RECT 42.955 171.425 43.965 171.595 ;
        RECT 44.135 171.580 44.885 171.770 ;
        RECT 42.615 171.085 43.740 171.255 ;
        RECT 44.135 170.915 44.305 171.580 ;
        RECT 45.055 171.335 45.395 172.145 ;
        RECT 46.025 171.595 46.715 172.155 ;
        RECT 46.885 171.425 47.095 172.325 ;
        RECT 42.275 170.745 44.305 170.915 ;
        RECT 44.475 170.575 44.645 171.335 ;
        RECT 44.880 170.925 45.395 171.335 ;
        RECT 46.140 171.205 47.095 171.425 ;
        RECT 47.265 172.155 47.665 172.955 ;
        RECT 47.855 172.495 48.135 172.955 ;
        RECT 48.655 172.665 48.980 173.125 ;
        RECT 47.855 172.325 48.980 172.495 ;
        RECT 49.150 172.385 49.535 172.955 ;
        RECT 48.530 172.215 48.980 172.325 ;
        RECT 47.265 171.595 48.360 172.155 ;
        RECT 48.530 171.885 49.085 172.215 ;
        RECT 46.140 170.745 46.425 171.205 ;
        RECT 46.595 170.575 46.865 171.035 ;
        RECT 47.265 170.745 47.665 171.595 ;
        RECT 48.530 171.425 48.980 171.885 ;
        RECT 49.255 171.715 49.535 172.385 ;
        RECT 47.855 171.205 48.980 171.425 ;
        RECT 47.855 170.745 48.135 171.205 ;
        RECT 48.655 170.575 48.980 171.035 ;
        RECT 49.150 170.745 49.535 171.715 ;
        RECT 49.710 172.385 49.965 172.955 ;
        RECT 50.135 172.725 50.465 173.125 ;
        RECT 50.890 172.590 51.420 172.955 ;
        RECT 50.890 172.555 51.065 172.590 ;
        RECT 50.135 172.385 51.065 172.555 ;
        RECT 51.610 172.445 51.885 172.955 ;
        RECT 49.710 171.715 49.880 172.385 ;
        RECT 50.135 172.215 50.305 172.385 ;
        RECT 50.050 171.885 50.305 172.215 ;
        RECT 50.530 171.885 50.725 172.215 ;
        RECT 49.710 170.745 50.045 171.715 ;
        RECT 50.215 170.575 50.385 171.715 ;
        RECT 50.555 170.915 50.725 171.885 ;
        RECT 50.895 171.255 51.065 172.385 ;
        RECT 51.235 171.595 51.405 172.395 ;
        RECT 51.605 172.275 51.885 172.445 ;
        RECT 51.610 171.795 51.885 172.275 ;
        RECT 52.055 171.595 52.245 172.955 ;
        RECT 52.425 172.590 52.935 173.125 ;
        RECT 53.155 172.315 53.400 172.920 ;
        RECT 53.935 172.645 54.235 173.125 ;
        RECT 54.405 172.475 54.665 172.930 ;
        RECT 54.835 172.645 55.095 173.125 ;
        RECT 55.275 172.475 55.535 172.930 ;
        RECT 55.705 172.645 55.955 173.125 ;
        RECT 56.135 172.475 56.395 172.930 ;
        RECT 56.565 172.645 56.815 173.125 ;
        RECT 56.995 172.475 57.255 172.930 ;
        RECT 57.425 172.645 57.670 173.125 ;
        RECT 57.840 172.475 58.115 172.930 ;
        RECT 58.285 172.645 58.530 173.125 ;
        RECT 58.700 172.475 58.960 172.930 ;
        RECT 59.130 172.645 59.390 173.125 ;
        RECT 59.560 172.475 59.820 172.930 ;
        RECT 59.990 172.645 60.250 173.125 ;
        RECT 60.420 172.475 60.680 172.930 ;
        RECT 60.850 172.565 61.110 173.125 ;
        RECT 52.445 172.145 53.675 172.315 ;
        RECT 51.235 171.425 52.245 171.595 ;
        RECT 52.415 171.580 53.165 171.770 ;
        RECT 50.895 171.085 52.020 171.255 ;
        RECT 52.415 170.915 52.585 171.580 ;
        RECT 53.335 171.335 53.675 172.145 ;
        RECT 53.935 172.305 60.680 172.475 ;
        RECT 53.935 171.715 55.100 172.305 ;
        RECT 61.280 172.135 61.530 172.945 ;
        RECT 61.710 172.600 61.970 173.125 ;
        RECT 62.140 172.135 62.390 172.945 ;
        RECT 62.570 172.615 62.875 173.125 ;
        RECT 55.270 171.885 62.390 172.135 ;
        RECT 62.560 171.885 62.875 172.445 ;
        RECT 63.045 172.400 63.335 173.125 ;
        RECT 63.545 172.305 63.775 173.125 ;
        RECT 63.945 172.325 64.275 172.955 ;
        RECT 63.525 171.885 63.855 172.135 ;
        RECT 53.935 171.490 60.680 171.715 ;
        RECT 50.555 170.745 52.585 170.915 ;
        RECT 52.755 170.575 52.925 171.335 ;
        RECT 53.160 170.925 53.675 171.335 ;
        RECT 53.935 170.575 54.205 171.320 ;
        RECT 54.375 170.750 54.665 171.490 ;
        RECT 55.275 171.475 60.680 171.490 ;
        RECT 54.835 170.580 55.090 171.305 ;
        RECT 55.275 170.750 55.535 171.475 ;
        RECT 55.705 170.580 55.950 171.305 ;
        RECT 56.135 170.750 56.395 171.475 ;
        RECT 56.565 170.580 56.810 171.305 ;
        RECT 56.995 170.750 57.255 171.475 ;
        RECT 57.425 170.580 57.670 171.305 ;
        RECT 57.840 170.750 58.100 171.475 ;
        RECT 58.270 170.580 58.530 171.305 ;
        RECT 58.700 170.750 58.960 171.475 ;
        RECT 59.130 170.580 59.390 171.305 ;
        RECT 59.560 170.750 59.820 171.475 ;
        RECT 59.990 170.580 60.250 171.305 ;
        RECT 60.420 170.750 60.680 171.475 ;
        RECT 60.850 170.580 61.110 171.375 ;
        RECT 61.280 170.750 61.530 171.885 ;
        RECT 54.835 170.575 61.110 170.580 ;
        RECT 61.710 170.575 61.970 171.385 ;
        RECT 62.145 170.745 62.390 171.885 ;
        RECT 62.570 170.575 62.865 171.385 ;
        RECT 63.045 170.575 63.335 171.740 ;
        RECT 64.025 171.725 64.275 172.325 ;
        RECT 64.445 172.305 64.655 173.125 ;
        RECT 64.890 172.415 65.145 172.945 ;
        RECT 65.315 172.665 65.620 173.125 ;
        RECT 65.865 172.745 66.935 172.915 ;
        RECT 63.545 170.575 63.775 171.715 ;
        RECT 63.945 170.745 64.275 171.725 ;
        RECT 64.890 171.765 65.100 172.415 ;
        RECT 65.865 172.390 66.185 172.745 ;
        RECT 65.860 172.215 66.185 172.390 ;
        RECT 65.270 171.915 66.185 172.215 ;
        RECT 66.355 172.175 66.595 172.575 ;
        RECT 66.765 172.515 66.935 172.745 ;
        RECT 67.105 172.685 67.295 173.125 ;
        RECT 67.465 172.675 68.415 172.955 ;
        RECT 68.635 172.765 68.985 172.935 ;
        RECT 66.765 172.345 67.295 172.515 ;
        RECT 65.270 171.885 66.010 171.915 ;
        RECT 64.445 170.575 64.655 171.715 ;
        RECT 64.890 170.885 65.145 171.765 ;
        RECT 65.315 170.575 65.620 171.715 ;
        RECT 65.840 171.295 66.010 171.885 ;
        RECT 66.355 171.805 66.895 172.175 ;
        RECT 67.075 172.065 67.295 172.345 ;
        RECT 67.465 171.895 67.635 172.675 ;
        RECT 67.230 171.725 67.635 171.895 ;
        RECT 67.805 171.885 68.155 172.505 ;
        RECT 67.230 171.635 67.400 171.725 ;
        RECT 68.325 171.715 68.535 172.505 ;
        RECT 66.180 171.465 67.400 171.635 ;
        RECT 67.860 171.555 68.535 171.715 ;
        RECT 65.840 171.125 66.640 171.295 ;
        RECT 65.960 170.575 66.290 170.955 ;
        RECT 66.470 170.835 66.640 171.125 ;
        RECT 67.230 171.085 67.400 171.465 ;
        RECT 67.570 171.545 68.535 171.555 ;
        RECT 68.725 172.375 68.985 172.765 ;
        RECT 69.195 172.665 69.525 173.125 ;
        RECT 70.400 172.735 71.255 172.905 ;
        RECT 71.460 172.735 71.955 172.905 ;
        RECT 72.125 172.765 72.455 173.125 ;
        RECT 68.725 171.685 68.895 172.375 ;
        RECT 69.065 172.025 69.235 172.205 ;
        RECT 69.405 172.195 70.195 172.445 ;
        RECT 70.400 172.025 70.570 172.735 ;
        RECT 70.740 172.225 71.095 172.445 ;
        RECT 69.065 171.855 70.755 172.025 ;
        RECT 67.570 171.255 68.030 171.545 ;
        RECT 68.725 171.515 70.225 171.685 ;
        RECT 68.725 171.375 68.895 171.515 ;
        RECT 68.335 171.205 68.895 171.375 ;
        RECT 66.810 170.575 67.060 171.035 ;
        RECT 67.230 170.745 68.100 171.085 ;
        RECT 68.335 170.745 68.505 171.205 ;
        RECT 69.340 171.175 70.415 171.345 ;
        RECT 68.675 170.575 69.045 171.035 ;
        RECT 69.340 170.835 69.510 171.175 ;
        RECT 69.680 170.575 70.010 171.005 ;
        RECT 70.245 170.835 70.415 171.175 ;
        RECT 70.585 171.075 70.755 171.855 ;
        RECT 70.925 171.635 71.095 172.225 ;
        RECT 71.265 171.825 71.615 172.445 ;
        RECT 70.925 171.245 71.390 171.635 ;
        RECT 71.785 171.375 71.955 172.735 ;
        RECT 72.125 171.545 72.585 172.595 ;
        RECT 71.560 171.205 71.955 171.375 ;
        RECT 71.560 171.075 71.730 171.205 ;
        RECT 70.585 170.745 71.265 171.075 ;
        RECT 71.480 170.745 71.730 171.075 ;
        RECT 71.900 170.575 72.150 171.035 ;
        RECT 72.320 170.760 72.645 171.545 ;
        RECT 72.815 170.745 72.985 172.865 ;
        RECT 73.155 172.745 73.485 173.125 ;
        RECT 73.655 172.575 73.910 172.865 ;
        RECT 75.065 172.645 75.345 173.125 ;
        RECT 73.160 172.405 73.910 172.575 ;
        RECT 75.515 172.475 75.775 172.865 ;
        RECT 75.950 172.645 76.205 173.125 ;
        RECT 76.375 172.475 76.670 172.865 ;
        RECT 76.850 172.645 77.125 173.125 ;
        RECT 77.295 172.625 77.595 172.955 ;
        RECT 73.160 171.415 73.390 172.405 ;
        RECT 75.020 172.305 76.670 172.475 ;
        RECT 73.560 171.585 73.910 172.235 ;
        RECT 75.020 171.795 75.425 172.305 ;
        RECT 75.595 171.965 76.735 172.135 ;
        RECT 75.020 171.625 75.775 171.795 ;
        RECT 73.160 171.245 73.910 171.415 ;
        RECT 73.155 170.575 73.485 171.075 ;
        RECT 73.655 170.745 73.910 171.245 ;
        RECT 75.060 170.575 75.345 171.445 ;
        RECT 75.515 171.375 75.775 171.625 ;
        RECT 76.565 171.715 76.735 171.965 ;
        RECT 76.905 171.885 77.255 172.455 ;
        RECT 77.425 171.715 77.595 172.625 ;
        RECT 78.230 172.285 78.490 173.125 ;
        RECT 78.665 172.380 78.920 172.955 ;
        RECT 79.090 172.745 79.420 173.125 ;
        RECT 79.635 172.575 79.805 172.955 ;
        RECT 79.090 172.405 79.805 172.575 ;
        RECT 76.565 171.545 77.595 171.715 ;
        RECT 75.515 171.205 76.635 171.375 ;
        RECT 75.515 170.745 75.775 171.205 ;
        RECT 75.950 170.575 76.205 171.035 ;
        RECT 76.375 170.745 76.635 171.205 ;
        RECT 76.805 170.575 77.115 171.375 ;
        RECT 77.285 170.745 77.595 171.545 ;
        RECT 78.230 170.575 78.490 171.725 ;
        RECT 78.665 171.650 78.835 172.380 ;
        RECT 79.090 172.215 79.260 172.405 ;
        RECT 80.525 172.355 83.115 173.125 ;
        RECT 79.005 171.885 79.260 172.215 ;
        RECT 79.090 171.675 79.260 171.885 ;
        RECT 79.540 171.855 79.895 172.225 ;
        RECT 78.665 170.745 78.920 171.650 ;
        RECT 79.090 171.505 79.805 171.675 ;
        RECT 79.090 170.575 79.420 171.335 ;
        RECT 79.635 170.745 79.805 171.505 ;
        RECT 80.525 171.665 81.735 172.185 ;
        RECT 81.905 171.835 83.115 172.355 ;
        RECT 83.345 172.305 83.555 173.125 ;
        RECT 83.725 172.325 84.055 172.955 ;
        RECT 83.725 171.725 83.975 172.325 ;
        RECT 84.225 172.305 84.455 173.125 ;
        RECT 84.940 172.315 85.185 172.920 ;
        RECT 85.405 172.590 85.915 173.125 ;
        RECT 84.665 172.145 85.895 172.315 ;
        RECT 84.145 171.885 84.475 172.135 ;
        RECT 80.525 170.575 83.115 171.665 ;
        RECT 83.345 170.575 83.555 171.715 ;
        RECT 83.725 170.745 84.055 171.725 ;
        RECT 84.225 170.575 84.455 171.715 ;
        RECT 84.665 171.335 85.005 172.145 ;
        RECT 85.175 171.580 85.925 171.770 ;
        RECT 84.665 170.925 85.180 171.335 ;
        RECT 85.415 170.575 85.585 171.335 ;
        RECT 85.755 170.915 85.925 171.580 ;
        RECT 86.095 171.595 86.285 172.955 ;
        RECT 86.455 172.105 86.730 172.955 ;
        RECT 86.920 172.590 87.450 172.955 ;
        RECT 87.875 172.725 88.205 173.125 ;
        RECT 87.275 172.555 87.450 172.590 ;
        RECT 86.455 171.935 86.735 172.105 ;
        RECT 86.455 171.795 86.730 171.935 ;
        RECT 86.935 171.595 87.105 172.395 ;
        RECT 86.095 171.425 87.105 171.595 ;
        RECT 87.275 172.385 88.205 172.555 ;
        RECT 88.375 172.385 88.630 172.955 ;
        RECT 88.805 172.400 89.095 173.125 ;
        RECT 90.185 172.615 90.490 173.125 ;
        RECT 87.275 171.255 87.445 172.385 ;
        RECT 88.035 172.215 88.205 172.385 ;
        RECT 86.320 171.085 87.445 171.255 ;
        RECT 87.615 171.885 87.810 172.215 ;
        RECT 88.035 171.885 88.290 172.215 ;
        RECT 87.615 170.915 87.785 171.885 ;
        RECT 88.460 171.715 88.630 172.385 ;
        RECT 90.185 171.885 90.500 172.445 ;
        RECT 90.670 172.135 90.920 172.945 ;
        RECT 91.090 172.600 91.350 173.125 ;
        RECT 91.530 172.135 91.780 172.945 ;
        RECT 91.950 172.565 92.210 173.125 ;
        RECT 92.380 172.475 92.640 172.930 ;
        RECT 92.810 172.645 93.070 173.125 ;
        RECT 93.240 172.475 93.500 172.930 ;
        RECT 93.670 172.645 93.930 173.125 ;
        RECT 94.100 172.475 94.360 172.930 ;
        RECT 94.530 172.645 94.775 173.125 ;
        RECT 94.945 172.475 95.220 172.930 ;
        RECT 95.390 172.645 95.635 173.125 ;
        RECT 95.805 172.475 96.065 172.930 ;
        RECT 96.245 172.645 96.495 173.125 ;
        RECT 96.665 172.475 96.925 172.930 ;
        RECT 97.105 172.645 97.355 173.125 ;
        RECT 97.525 172.475 97.785 172.930 ;
        RECT 97.965 172.645 98.225 173.125 ;
        RECT 98.395 172.475 98.655 172.930 ;
        RECT 98.825 172.645 99.125 173.125 ;
        RECT 92.380 172.305 99.125 172.475 ;
        RECT 90.670 171.885 97.790 172.135 ;
        RECT 85.755 170.745 87.785 170.915 ;
        RECT 87.955 170.575 88.125 171.715 ;
        RECT 88.295 170.745 88.630 171.715 ;
        RECT 88.805 170.575 89.095 171.740 ;
        RECT 90.195 170.575 90.490 171.385 ;
        RECT 90.670 170.745 90.915 171.885 ;
        RECT 91.090 170.575 91.350 171.385 ;
        RECT 91.530 170.750 91.780 171.885 ;
        RECT 97.960 171.715 99.125 172.305 ;
        RECT 92.380 171.490 99.125 171.715 ;
        RECT 99.760 172.415 100.015 172.945 ;
        RECT 100.195 172.665 100.480 173.125 ;
        RECT 99.760 171.555 99.940 172.415 ;
        RECT 100.660 172.215 100.910 172.865 ;
        RECT 100.110 171.885 100.910 172.215 ;
        RECT 92.380 171.475 97.785 171.490 ;
        RECT 91.950 170.580 92.210 171.375 ;
        RECT 92.380 170.750 92.640 171.475 ;
        RECT 92.810 170.580 93.070 171.305 ;
        RECT 93.240 170.750 93.500 171.475 ;
        RECT 93.670 170.580 93.930 171.305 ;
        RECT 94.100 170.750 94.360 171.475 ;
        RECT 94.530 170.580 94.790 171.305 ;
        RECT 94.960 170.750 95.220 171.475 ;
        RECT 95.390 170.580 95.635 171.305 ;
        RECT 95.805 170.750 96.065 171.475 ;
        RECT 96.250 170.580 96.495 171.305 ;
        RECT 96.665 170.750 96.925 171.475 ;
        RECT 97.110 170.580 97.355 171.305 ;
        RECT 97.525 170.750 97.785 171.475 ;
        RECT 97.970 170.580 98.225 171.305 ;
        RECT 98.395 170.750 98.685 171.490 ;
        RECT 91.950 170.575 98.225 170.580 ;
        RECT 98.855 170.575 99.125 171.320 ;
        RECT 99.760 171.085 100.015 171.555 ;
        RECT 99.675 170.915 100.015 171.085 ;
        RECT 99.760 170.885 100.015 170.915 ;
        RECT 100.195 170.575 100.480 171.375 ;
        RECT 100.660 171.295 100.910 171.885 ;
        RECT 101.110 172.530 101.430 172.860 ;
        RECT 101.610 172.645 102.270 173.125 ;
        RECT 102.470 172.735 103.320 172.905 ;
        RECT 101.110 171.635 101.300 172.530 ;
        RECT 101.620 172.205 102.280 172.475 ;
        RECT 101.950 172.145 102.280 172.205 ;
        RECT 101.470 171.975 101.800 172.035 ;
        RECT 102.470 171.975 102.640 172.735 ;
        RECT 103.880 172.665 104.200 173.125 ;
        RECT 104.400 172.485 104.650 172.915 ;
        RECT 104.940 172.685 105.350 173.125 ;
        RECT 105.520 172.745 106.535 172.945 ;
        RECT 102.810 172.315 104.060 172.485 ;
        RECT 102.810 172.195 103.140 172.315 ;
        RECT 101.470 171.805 103.370 171.975 ;
        RECT 101.110 171.465 103.030 171.635 ;
        RECT 101.110 171.445 101.430 171.465 ;
        RECT 100.660 170.785 100.990 171.295 ;
        RECT 101.260 170.835 101.430 171.445 ;
        RECT 103.200 171.295 103.370 171.805 ;
        RECT 103.540 171.735 103.720 172.145 ;
        RECT 103.890 171.555 104.060 172.315 ;
        RECT 101.600 170.575 101.930 171.265 ;
        RECT 102.160 171.125 103.370 171.295 ;
        RECT 103.540 171.245 104.060 171.555 ;
        RECT 104.230 172.145 104.650 172.485 ;
        RECT 104.940 172.145 105.350 172.475 ;
        RECT 104.230 171.375 104.420 172.145 ;
        RECT 105.520 172.015 105.690 172.745 ;
        RECT 106.835 172.575 107.005 172.905 ;
        RECT 107.175 172.745 107.505 173.125 ;
        RECT 105.860 172.195 106.210 172.565 ;
        RECT 105.520 171.975 105.940 172.015 ;
        RECT 104.590 171.805 105.940 171.975 ;
        RECT 104.590 171.645 104.840 171.805 ;
        RECT 105.350 171.375 105.600 171.635 ;
        RECT 104.230 171.125 105.600 171.375 ;
        RECT 102.160 170.835 102.400 171.125 ;
        RECT 103.200 171.045 103.370 171.125 ;
        RECT 102.600 170.575 103.020 170.955 ;
        RECT 103.200 170.795 103.830 171.045 ;
        RECT 104.300 170.575 104.630 170.955 ;
        RECT 104.800 170.835 104.970 171.125 ;
        RECT 105.770 170.960 105.940 171.805 ;
        RECT 106.390 171.635 106.610 172.505 ;
        RECT 106.835 172.385 107.530 172.575 ;
        RECT 106.110 171.255 106.610 171.635 ;
        RECT 106.780 171.585 107.190 172.205 ;
        RECT 107.360 171.415 107.530 172.385 ;
        RECT 106.835 171.245 107.530 171.415 ;
        RECT 105.150 170.575 105.530 170.955 ;
        RECT 105.770 170.790 106.600 170.960 ;
        RECT 106.835 170.745 107.005 171.245 ;
        RECT 107.175 170.575 107.505 171.075 ;
        RECT 107.720 170.745 107.945 172.865 ;
        RECT 108.115 172.745 108.445 173.125 ;
        RECT 108.615 172.575 108.785 172.865 ;
        RECT 108.120 172.405 108.785 172.575 ;
        RECT 109.045 172.450 109.305 172.955 ;
        RECT 109.485 172.745 109.815 173.125 ;
        RECT 109.995 172.575 110.165 172.955 ;
        RECT 108.120 171.415 108.350 172.405 ;
        RECT 108.520 171.585 108.870 172.235 ;
        RECT 109.045 171.650 109.215 172.450 ;
        RECT 109.500 172.405 110.165 172.575 ;
        RECT 109.500 172.150 109.670 172.405 ;
        RECT 110.425 172.385 110.810 172.955 ;
        RECT 110.980 172.665 111.305 173.125 ;
        RECT 111.825 172.495 112.105 172.955 ;
        RECT 109.385 171.820 109.670 172.150 ;
        RECT 109.905 171.855 110.235 172.225 ;
        RECT 109.500 171.675 109.670 171.820 ;
        RECT 110.425 171.715 110.705 172.385 ;
        RECT 110.980 172.325 112.105 172.495 ;
        RECT 110.980 172.215 111.430 172.325 ;
        RECT 110.875 171.885 111.430 172.215 ;
        RECT 112.295 172.155 112.695 172.955 ;
        RECT 113.095 172.665 113.365 173.125 ;
        RECT 113.535 172.495 113.820 172.955 ;
        RECT 108.120 171.245 108.785 171.415 ;
        RECT 108.115 170.575 108.445 171.075 ;
        RECT 108.615 170.745 108.785 171.245 ;
        RECT 109.045 170.745 109.315 171.650 ;
        RECT 109.500 171.505 110.165 171.675 ;
        RECT 109.485 170.575 109.815 171.335 ;
        RECT 109.995 170.745 110.165 171.505 ;
        RECT 110.425 170.745 110.810 171.715 ;
        RECT 110.980 171.425 111.430 171.885 ;
        RECT 111.600 171.595 112.695 172.155 ;
        RECT 110.980 171.205 112.105 171.425 ;
        RECT 110.980 170.575 111.305 171.035 ;
        RECT 111.825 170.745 112.105 171.205 ;
        RECT 112.295 170.745 112.695 171.595 ;
        RECT 112.865 172.325 113.820 172.495 ;
        RECT 114.565 172.400 114.855 173.125 ;
        RECT 112.865 171.425 113.075 172.325 ;
        RECT 116.220 172.315 116.465 172.920 ;
        RECT 116.685 172.590 117.195 173.125 ;
        RECT 113.245 171.595 113.935 172.155 ;
        RECT 115.945 172.145 117.175 172.315 ;
        RECT 112.865 171.205 113.820 171.425 ;
        RECT 113.095 170.575 113.365 171.035 ;
        RECT 113.535 170.745 113.820 171.205 ;
        RECT 114.565 170.575 114.855 171.740 ;
        RECT 115.945 171.335 116.285 172.145 ;
        RECT 116.455 171.580 117.205 171.770 ;
        RECT 115.945 170.925 116.460 171.335 ;
        RECT 116.695 170.575 116.865 171.335 ;
        RECT 117.035 170.915 117.205 171.580 ;
        RECT 117.375 171.595 117.565 172.955 ;
        RECT 117.735 172.785 118.010 172.955 ;
        RECT 117.735 172.615 118.015 172.785 ;
        RECT 117.735 171.795 118.010 172.615 ;
        RECT 118.200 172.590 118.730 172.955 ;
        RECT 119.155 172.725 119.485 173.125 ;
        RECT 118.555 172.555 118.730 172.590 ;
        RECT 118.215 171.595 118.385 172.395 ;
        RECT 117.375 171.425 118.385 171.595 ;
        RECT 118.555 172.385 119.485 172.555 ;
        RECT 119.655 172.385 119.910 172.955 ;
        RECT 118.555 171.255 118.725 172.385 ;
        RECT 119.315 172.215 119.485 172.385 ;
        RECT 117.600 171.085 118.725 171.255 ;
        RECT 118.895 171.885 119.090 172.215 ;
        RECT 119.315 171.885 119.570 172.215 ;
        RECT 118.895 170.915 119.065 171.885 ;
        RECT 119.740 171.715 119.910 172.385 ;
        RECT 120.125 172.305 120.355 173.125 ;
        RECT 120.525 172.325 120.855 172.955 ;
        RECT 120.105 171.885 120.435 172.135 ;
        RECT 120.605 171.725 120.855 172.325 ;
        RECT 121.025 172.305 121.235 173.125 ;
        RECT 121.555 172.575 121.725 172.955 ;
        RECT 121.905 172.745 122.235 173.125 ;
        RECT 121.555 172.405 122.220 172.575 ;
        RECT 122.415 172.450 122.675 172.955 ;
        RECT 121.485 171.855 121.815 172.225 ;
        RECT 122.050 172.150 122.220 172.405 ;
        RECT 117.035 170.745 119.065 170.915 ;
        RECT 119.235 170.575 119.405 171.715 ;
        RECT 119.575 170.745 119.910 171.715 ;
        RECT 120.125 170.575 120.355 171.715 ;
        RECT 120.525 170.745 120.855 171.725 ;
        RECT 122.050 171.820 122.335 172.150 ;
        RECT 121.025 170.575 121.235 171.715 ;
        RECT 122.050 171.675 122.220 171.820 ;
        RECT 121.555 171.505 122.220 171.675 ;
        RECT 122.505 171.650 122.675 172.450 ;
        RECT 122.935 172.575 123.105 172.955 ;
        RECT 123.285 172.745 123.615 173.125 ;
        RECT 122.935 172.405 123.600 172.575 ;
        RECT 123.795 172.450 124.055 172.955 ;
        RECT 122.865 171.855 123.195 172.225 ;
        RECT 123.430 172.150 123.600 172.405 ;
        RECT 123.430 171.820 123.715 172.150 ;
        RECT 123.430 171.675 123.600 171.820 ;
        RECT 121.555 170.745 121.725 171.505 ;
        RECT 121.905 170.575 122.235 171.335 ;
        RECT 122.405 170.745 122.675 171.650 ;
        RECT 122.935 171.505 123.600 171.675 ;
        RECT 123.885 171.650 124.055 172.450 ;
        RECT 124.685 172.355 126.355 173.125 ;
        RECT 126.525 172.375 127.735 173.125 ;
        RECT 122.935 170.745 123.105 171.505 ;
        RECT 123.285 170.575 123.615 171.335 ;
        RECT 123.785 170.745 124.055 171.650 ;
        RECT 124.685 171.665 125.435 172.185 ;
        RECT 125.605 171.835 126.355 172.355 ;
        RECT 126.525 171.665 127.045 172.205 ;
        RECT 127.215 171.835 127.735 172.375 ;
        RECT 124.685 170.575 126.355 171.665 ;
        RECT 126.525 170.575 127.735 171.665 ;
        RECT 29.840 170.405 127.820 170.575 ;
        RECT 29.925 169.315 31.135 170.405 ;
        RECT 29.925 168.605 30.445 169.145 ;
        RECT 30.615 168.775 31.135 169.315 ;
        RECT 31.680 169.425 31.935 170.095 ;
        RECT 32.115 169.605 32.400 170.405 ;
        RECT 32.580 169.685 32.910 170.195 ;
        RECT 29.925 167.855 31.135 168.605 ;
        RECT 31.680 168.565 31.860 169.425 ;
        RECT 32.580 169.095 32.830 169.685 ;
        RECT 33.180 169.535 33.350 170.145 ;
        RECT 33.520 169.715 33.850 170.405 ;
        RECT 34.080 169.855 34.320 170.145 ;
        RECT 34.520 170.025 34.940 170.405 ;
        RECT 35.120 169.935 35.750 170.185 ;
        RECT 36.220 170.025 36.550 170.405 ;
        RECT 35.120 169.855 35.290 169.935 ;
        RECT 36.720 169.855 36.890 170.145 ;
        RECT 37.070 170.025 37.450 170.405 ;
        RECT 37.690 170.020 38.520 170.190 ;
        RECT 34.080 169.685 35.290 169.855 ;
        RECT 32.030 168.765 32.830 169.095 ;
        RECT 31.680 168.365 31.935 168.565 ;
        RECT 31.595 168.195 31.935 168.365 ;
        RECT 31.680 168.035 31.935 168.195 ;
        RECT 32.115 167.855 32.400 168.315 ;
        RECT 32.580 168.115 32.830 168.765 ;
        RECT 33.030 169.515 33.350 169.535 ;
        RECT 33.030 169.345 34.950 169.515 ;
        RECT 33.030 168.450 33.220 169.345 ;
        RECT 35.120 169.175 35.290 169.685 ;
        RECT 35.460 169.425 35.980 169.735 ;
        RECT 33.390 169.005 35.290 169.175 ;
        RECT 33.390 168.945 33.720 169.005 ;
        RECT 33.870 168.775 34.200 168.835 ;
        RECT 33.540 168.505 34.200 168.775 ;
        RECT 33.030 168.120 33.350 168.450 ;
        RECT 33.530 167.855 34.190 168.335 ;
        RECT 34.390 168.245 34.560 169.005 ;
        RECT 35.460 168.835 35.640 169.245 ;
        RECT 34.730 168.665 35.060 168.785 ;
        RECT 35.810 168.665 35.980 169.425 ;
        RECT 34.730 168.495 35.980 168.665 ;
        RECT 36.150 169.605 37.520 169.855 ;
        RECT 36.150 168.835 36.340 169.605 ;
        RECT 37.270 169.345 37.520 169.605 ;
        RECT 36.510 169.175 36.760 169.335 ;
        RECT 37.690 169.175 37.860 170.020 ;
        RECT 38.755 169.735 38.925 170.235 ;
        RECT 39.095 169.905 39.425 170.405 ;
        RECT 38.030 169.345 38.530 169.725 ;
        RECT 38.755 169.565 39.450 169.735 ;
        RECT 36.510 169.005 37.860 169.175 ;
        RECT 37.440 168.965 37.860 169.005 ;
        RECT 36.150 168.495 36.570 168.835 ;
        RECT 36.860 168.505 37.270 168.835 ;
        RECT 34.390 168.075 35.240 168.245 ;
        RECT 35.800 167.855 36.120 168.315 ;
        RECT 36.320 168.065 36.570 168.495 ;
        RECT 36.860 167.855 37.270 168.295 ;
        RECT 37.440 168.235 37.610 168.965 ;
        RECT 37.780 168.415 38.130 168.785 ;
        RECT 38.310 168.475 38.530 169.345 ;
        RECT 38.700 168.775 39.110 169.395 ;
        RECT 39.280 168.595 39.450 169.565 ;
        RECT 38.755 168.405 39.450 168.595 ;
        RECT 37.440 168.035 38.455 168.235 ;
        RECT 38.755 168.075 38.925 168.405 ;
        RECT 39.095 167.855 39.425 168.235 ;
        RECT 39.640 168.115 39.865 170.235 ;
        RECT 40.035 169.905 40.365 170.405 ;
        RECT 40.535 169.735 40.705 170.235 ;
        RECT 40.040 169.565 40.705 169.735 ;
        RECT 40.040 168.575 40.270 169.565 ;
        RECT 40.440 168.745 40.790 169.395 ;
        RECT 40.970 169.265 41.305 170.235 ;
        RECT 41.475 169.265 41.645 170.405 ;
        RECT 41.815 170.065 43.845 170.235 ;
        RECT 40.970 168.595 41.140 169.265 ;
        RECT 41.815 169.095 41.985 170.065 ;
        RECT 41.310 168.765 41.565 169.095 ;
        RECT 41.790 168.765 41.985 169.095 ;
        RECT 42.155 169.725 43.280 169.895 ;
        RECT 41.395 168.595 41.565 168.765 ;
        RECT 42.155 168.595 42.325 169.725 ;
        RECT 40.040 168.405 40.705 168.575 ;
        RECT 40.035 167.855 40.365 168.235 ;
        RECT 40.535 168.115 40.705 168.405 ;
        RECT 40.970 168.025 41.225 168.595 ;
        RECT 41.395 168.425 42.325 168.595 ;
        RECT 42.495 169.385 43.505 169.555 ;
        RECT 42.495 168.585 42.665 169.385 ;
        RECT 42.150 168.390 42.325 168.425 ;
        RECT 41.395 167.855 41.725 168.255 ;
        RECT 42.150 168.025 42.680 168.390 ;
        RECT 42.870 168.365 43.145 169.185 ;
        RECT 42.865 168.195 43.145 168.365 ;
        RECT 42.870 168.025 43.145 168.195 ;
        RECT 43.315 168.025 43.505 169.385 ;
        RECT 43.675 169.400 43.845 170.065 ;
        RECT 44.015 169.645 44.185 170.405 ;
        RECT 44.420 169.645 44.935 170.055 ;
        RECT 43.675 169.210 44.425 169.400 ;
        RECT 44.595 168.835 44.935 169.645 ;
        RECT 43.705 168.665 44.935 168.835 ;
        RECT 45.105 169.315 46.315 170.405 ;
        RECT 46.690 169.435 47.020 170.235 ;
        RECT 47.190 169.605 47.520 170.405 ;
        RECT 47.820 169.435 48.150 170.235 ;
        RECT 48.795 169.605 49.045 170.405 ;
        RECT 45.105 168.775 45.625 169.315 ;
        RECT 46.690 169.265 49.125 169.435 ;
        RECT 49.315 169.265 49.485 170.405 ;
        RECT 49.655 169.265 49.995 170.235 ;
        RECT 43.685 167.855 44.195 168.390 ;
        RECT 44.415 168.060 44.660 168.665 ;
        RECT 45.795 168.605 46.315 169.145 ;
        RECT 46.485 168.845 46.835 169.095 ;
        RECT 47.020 168.635 47.190 169.265 ;
        RECT 47.360 168.845 47.690 169.045 ;
        RECT 47.860 168.845 48.190 169.045 ;
        RECT 48.360 168.845 48.780 169.045 ;
        RECT 48.955 169.015 49.125 169.265 ;
        RECT 48.955 168.845 49.650 169.015 ;
        RECT 45.105 167.855 46.315 168.605 ;
        RECT 46.690 168.025 47.190 168.635 ;
        RECT 47.820 168.505 49.045 168.675 ;
        RECT 49.820 168.655 49.995 169.265 ;
        RECT 50.165 169.240 50.455 170.405 ;
        RECT 51.175 169.475 51.345 170.235 ;
        RECT 51.525 169.645 51.855 170.405 ;
        RECT 51.175 169.305 51.840 169.475 ;
        RECT 52.025 169.330 52.295 170.235 ;
        RECT 51.670 169.160 51.840 169.305 ;
        RECT 51.105 168.755 51.435 169.125 ;
        RECT 51.670 168.830 51.955 169.160 ;
        RECT 47.820 168.025 48.150 168.505 ;
        RECT 48.320 167.855 48.545 168.315 ;
        RECT 48.715 168.025 49.045 168.505 ;
        RECT 49.235 167.855 49.485 168.655 ;
        RECT 49.655 168.025 49.995 168.655 ;
        RECT 50.165 167.855 50.455 168.580 ;
        RECT 51.670 168.575 51.840 168.830 ;
        RECT 51.175 168.405 51.840 168.575 ;
        RECT 52.125 168.530 52.295 169.330 ;
        RECT 52.670 169.435 53.000 170.235 ;
        RECT 53.170 169.605 53.500 170.405 ;
        RECT 53.800 169.435 54.130 170.235 ;
        RECT 54.775 169.605 55.025 170.405 ;
        RECT 52.670 169.265 55.105 169.435 ;
        RECT 55.295 169.265 55.465 170.405 ;
        RECT 55.635 169.265 55.975 170.235 ;
        RECT 56.260 169.775 56.545 170.235 ;
        RECT 56.715 169.945 56.985 170.405 ;
        RECT 56.260 169.555 57.215 169.775 ;
        RECT 52.465 168.845 52.815 169.095 ;
        RECT 53.000 168.635 53.170 169.265 ;
        RECT 53.340 168.845 53.670 169.045 ;
        RECT 53.840 168.845 54.170 169.045 ;
        RECT 54.340 168.845 54.760 169.045 ;
        RECT 54.935 169.015 55.105 169.265 ;
        RECT 54.935 168.845 55.630 169.015 ;
        RECT 51.175 168.025 51.345 168.405 ;
        RECT 51.525 167.855 51.855 168.235 ;
        RECT 52.035 168.025 52.295 168.530 ;
        RECT 52.670 168.025 53.170 168.635 ;
        RECT 53.800 168.505 55.025 168.675 ;
        RECT 55.800 168.655 55.975 169.265 ;
        RECT 56.145 168.825 56.835 169.385 ;
        RECT 57.005 168.655 57.215 169.555 ;
        RECT 53.800 168.025 54.130 168.505 ;
        RECT 54.300 167.855 54.525 168.315 ;
        RECT 54.695 168.025 55.025 168.505 ;
        RECT 55.215 167.855 55.465 168.655 ;
        RECT 55.635 168.025 55.975 168.655 ;
        RECT 56.260 168.485 57.215 168.655 ;
        RECT 57.385 169.385 57.785 170.235 ;
        RECT 57.975 169.775 58.255 170.235 ;
        RECT 58.775 169.945 59.100 170.405 ;
        RECT 57.975 169.555 59.100 169.775 ;
        RECT 57.385 168.825 58.480 169.385 ;
        RECT 58.650 169.095 59.100 169.555 ;
        RECT 59.270 169.265 59.655 170.235 ;
        RECT 59.880 169.605 60.180 170.405 ;
        RECT 60.350 169.435 60.680 170.235 ;
        RECT 60.850 169.605 61.020 170.405 ;
        RECT 61.190 169.435 61.520 170.235 ;
        RECT 61.690 169.605 61.860 170.405 ;
        RECT 62.030 169.435 62.360 170.235 ;
        RECT 62.530 169.605 62.700 170.405 ;
        RECT 62.870 169.435 63.200 170.235 ;
        RECT 63.370 169.605 63.625 170.405 ;
        RECT 56.260 168.025 56.545 168.485 ;
        RECT 56.715 167.855 56.985 168.315 ;
        RECT 57.385 168.025 57.785 168.825 ;
        RECT 58.650 168.765 59.205 169.095 ;
        RECT 58.650 168.655 59.100 168.765 ;
        RECT 57.975 168.485 59.100 168.655 ;
        RECT 59.375 168.595 59.655 169.265 ;
        RECT 57.975 168.025 58.255 168.485 ;
        RECT 58.775 167.855 59.100 168.315 ;
        RECT 59.270 168.025 59.655 168.595 ;
        RECT 59.825 169.265 63.795 169.435 ;
        RECT 59.825 168.675 60.145 169.265 ;
        RECT 60.345 168.845 63.200 169.095 ;
        RECT 63.450 168.675 63.795 169.265 ;
        RECT 63.965 169.315 66.555 170.405 ;
        RECT 63.965 168.795 65.175 169.315 ;
        RECT 66.730 169.215 66.985 170.095 ;
        RECT 67.155 169.265 67.460 170.405 ;
        RECT 67.800 170.025 68.130 170.405 ;
        RECT 68.310 169.855 68.480 170.145 ;
        RECT 68.650 169.945 68.900 170.405 ;
        RECT 67.680 169.685 68.480 169.855 ;
        RECT 69.070 169.895 69.940 170.235 ;
        RECT 59.825 168.485 63.795 168.675 ;
        RECT 65.345 168.625 66.555 169.145 ;
        RECT 59.875 167.855 60.180 168.315 ;
        RECT 60.350 168.025 60.680 168.485 ;
        RECT 60.850 167.855 61.020 168.315 ;
        RECT 61.190 168.025 61.520 168.485 ;
        RECT 61.690 167.855 61.860 168.315 ;
        RECT 62.030 168.025 62.360 168.485 ;
        RECT 62.530 167.855 62.700 168.315 ;
        RECT 62.870 168.025 63.200 168.485 ;
        RECT 63.370 167.855 63.625 168.315 ;
        RECT 63.965 167.855 66.555 168.625 ;
        RECT 66.730 168.565 66.940 169.215 ;
        RECT 67.680 169.095 67.850 169.685 ;
        RECT 69.070 169.515 69.240 169.895 ;
        RECT 70.175 169.775 70.345 170.235 ;
        RECT 70.515 169.945 70.885 170.405 ;
        RECT 71.180 169.805 71.350 170.145 ;
        RECT 71.520 169.975 71.850 170.405 ;
        RECT 72.085 169.805 72.255 170.145 ;
        RECT 68.020 169.345 69.240 169.515 ;
        RECT 69.410 169.435 69.870 169.725 ;
        RECT 70.175 169.605 70.735 169.775 ;
        RECT 71.180 169.635 72.255 169.805 ;
        RECT 72.425 169.905 73.105 170.235 ;
        RECT 73.320 169.905 73.570 170.235 ;
        RECT 73.740 169.945 73.990 170.405 ;
        RECT 70.565 169.465 70.735 169.605 ;
        RECT 69.410 169.425 70.375 169.435 ;
        RECT 69.070 169.255 69.240 169.345 ;
        RECT 69.700 169.265 70.375 169.425 ;
        RECT 67.110 169.065 67.850 169.095 ;
        RECT 67.110 168.765 68.025 169.065 ;
        RECT 67.700 168.590 68.025 168.765 ;
        RECT 66.730 168.035 66.985 168.565 ;
        RECT 67.155 167.855 67.460 168.315 ;
        RECT 67.705 168.235 68.025 168.590 ;
        RECT 68.195 168.805 68.735 169.175 ;
        RECT 69.070 169.085 69.475 169.255 ;
        RECT 68.195 168.405 68.435 168.805 ;
        RECT 68.915 168.635 69.135 168.915 ;
        RECT 68.605 168.465 69.135 168.635 ;
        RECT 68.605 168.235 68.775 168.465 ;
        RECT 69.305 168.305 69.475 169.085 ;
        RECT 69.645 168.475 69.995 169.095 ;
        RECT 70.165 168.475 70.375 169.265 ;
        RECT 70.565 169.295 72.065 169.465 ;
        RECT 70.565 168.605 70.735 169.295 ;
        RECT 72.425 169.125 72.595 169.905 ;
        RECT 73.400 169.775 73.570 169.905 ;
        RECT 70.905 168.955 72.595 169.125 ;
        RECT 72.765 169.345 73.230 169.735 ;
        RECT 73.400 169.605 73.795 169.775 ;
        RECT 70.905 168.775 71.075 168.955 ;
        RECT 67.705 168.065 68.775 168.235 ;
        RECT 68.945 167.855 69.135 168.295 ;
        RECT 69.305 168.025 70.255 168.305 ;
        RECT 70.565 168.215 70.825 168.605 ;
        RECT 71.245 168.535 72.035 168.785 ;
        RECT 70.475 168.045 70.825 168.215 ;
        RECT 71.035 167.855 71.365 168.315 ;
        RECT 72.240 168.245 72.410 168.955 ;
        RECT 72.765 168.755 72.935 169.345 ;
        RECT 72.580 168.535 72.935 168.755 ;
        RECT 73.105 168.535 73.455 169.155 ;
        RECT 73.625 168.245 73.795 169.605 ;
        RECT 74.160 169.435 74.485 170.220 ;
        RECT 73.965 168.385 74.425 169.435 ;
        RECT 72.240 168.075 73.095 168.245 ;
        RECT 73.300 168.075 73.795 168.245 ;
        RECT 73.965 167.855 74.295 168.215 ;
        RECT 74.655 168.115 74.825 170.235 ;
        RECT 74.995 169.905 75.325 170.405 ;
        RECT 75.495 169.735 75.750 170.235 ;
        RECT 75.000 169.565 75.750 169.735 ;
        RECT 75.000 168.575 75.230 169.565 ;
        RECT 75.400 168.745 75.750 169.395 ;
        RECT 75.925 169.240 76.215 170.405 ;
        RECT 77.310 169.255 77.570 170.405 ;
        RECT 77.745 169.330 78.000 170.235 ;
        RECT 78.170 169.645 78.500 170.405 ;
        RECT 78.715 169.475 78.885 170.235 ;
        RECT 75.000 168.405 75.750 168.575 ;
        RECT 74.995 167.855 75.325 168.235 ;
        RECT 75.495 168.115 75.750 168.405 ;
        RECT 75.925 167.855 76.215 168.580 ;
        RECT 77.310 167.855 77.570 168.695 ;
        RECT 77.745 168.600 77.915 169.330 ;
        RECT 78.170 169.305 78.885 169.475 ;
        RECT 78.170 169.095 78.340 169.305 ;
        RECT 79.150 169.255 79.410 170.405 ;
        RECT 79.585 169.330 79.840 170.235 ;
        RECT 80.010 169.645 80.340 170.405 ;
        RECT 80.555 169.475 80.725 170.235 ;
        RECT 78.085 168.765 78.340 169.095 ;
        RECT 77.745 168.025 78.000 168.600 ;
        RECT 78.170 168.575 78.340 168.765 ;
        RECT 78.620 168.755 78.975 169.125 ;
        RECT 78.170 168.405 78.885 168.575 ;
        RECT 78.170 167.855 78.500 168.235 ;
        RECT 78.715 168.025 78.885 168.405 ;
        RECT 79.150 167.855 79.410 168.695 ;
        RECT 79.585 168.600 79.755 169.330 ;
        RECT 80.010 169.305 80.725 169.475 ;
        RECT 80.985 169.315 82.195 170.405 ;
        RECT 80.010 169.095 80.180 169.305 ;
        RECT 79.925 168.765 80.180 169.095 ;
        RECT 79.585 168.025 79.840 168.600 ;
        RECT 80.010 168.575 80.180 168.765 ;
        RECT 80.460 168.755 80.815 169.125 ;
        RECT 80.985 168.775 81.505 169.315 ;
        RECT 82.365 169.265 82.705 170.235 ;
        RECT 82.875 169.265 83.045 170.405 ;
        RECT 83.315 169.605 83.565 170.405 ;
        RECT 84.210 169.435 84.540 170.235 ;
        RECT 84.840 169.605 85.170 170.405 ;
        RECT 85.340 169.435 85.670 170.235 ;
        RECT 83.235 169.265 85.670 169.435 ;
        RECT 86.045 169.645 86.560 170.055 ;
        RECT 86.795 169.645 86.965 170.405 ;
        RECT 87.135 170.065 89.165 170.235 ;
        RECT 81.675 168.605 82.195 169.145 ;
        RECT 80.010 168.405 80.725 168.575 ;
        RECT 80.010 167.855 80.340 168.235 ;
        RECT 80.555 168.025 80.725 168.405 ;
        RECT 80.985 167.855 82.195 168.605 ;
        RECT 82.365 168.655 82.540 169.265 ;
        RECT 83.235 169.015 83.405 169.265 ;
        RECT 82.710 168.845 83.405 169.015 ;
        RECT 83.580 168.845 84.000 169.045 ;
        RECT 84.170 168.845 84.500 169.045 ;
        RECT 84.670 168.845 85.000 169.045 ;
        RECT 82.365 168.025 82.705 168.655 ;
        RECT 82.875 167.855 83.125 168.655 ;
        RECT 83.315 168.505 84.540 168.675 ;
        RECT 83.315 168.025 83.645 168.505 ;
        RECT 83.815 167.855 84.040 168.315 ;
        RECT 84.210 168.025 84.540 168.505 ;
        RECT 85.170 168.635 85.340 169.265 ;
        RECT 85.525 168.845 85.875 169.095 ;
        RECT 86.045 168.835 86.385 169.645 ;
        RECT 87.135 169.400 87.305 170.065 ;
        RECT 87.700 169.725 88.825 169.895 ;
        RECT 86.555 169.210 87.305 169.400 ;
        RECT 87.475 169.385 88.485 169.555 ;
        RECT 86.045 168.665 87.275 168.835 ;
        RECT 85.170 168.025 85.670 168.635 ;
        RECT 86.320 168.060 86.565 168.665 ;
        RECT 86.785 167.855 87.295 168.390 ;
        RECT 87.475 168.025 87.665 169.385 ;
        RECT 87.835 168.365 88.110 169.185 ;
        RECT 88.315 168.585 88.485 169.385 ;
        RECT 88.655 168.595 88.825 169.725 ;
        RECT 88.995 169.095 89.165 170.065 ;
        RECT 89.335 169.265 89.505 170.405 ;
        RECT 89.675 169.265 90.010 170.235 ;
        RECT 90.735 169.475 90.905 170.235 ;
        RECT 91.085 169.645 91.415 170.405 ;
        RECT 90.735 169.305 91.400 169.475 ;
        RECT 91.585 169.330 91.855 170.235 ;
        RECT 88.995 168.765 89.190 169.095 ;
        RECT 89.415 168.765 89.670 169.095 ;
        RECT 89.415 168.595 89.585 168.765 ;
        RECT 89.840 168.595 90.010 169.265 ;
        RECT 91.230 169.160 91.400 169.305 ;
        RECT 90.665 168.755 90.995 169.125 ;
        RECT 91.230 168.830 91.515 169.160 ;
        RECT 88.655 168.425 89.585 168.595 ;
        RECT 88.655 168.390 88.830 168.425 ;
        RECT 87.835 168.195 88.115 168.365 ;
        RECT 87.835 168.025 88.110 168.195 ;
        RECT 88.300 168.025 88.830 168.390 ;
        RECT 89.255 167.855 89.585 168.255 ;
        RECT 89.755 168.025 90.010 168.595 ;
        RECT 91.230 168.575 91.400 168.830 ;
        RECT 90.735 168.405 91.400 168.575 ;
        RECT 91.685 168.530 91.855 169.330 ;
        RECT 92.025 169.315 93.235 170.405 ;
        RECT 93.520 169.775 93.805 170.235 ;
        RECT 93.975 169.945 94.245 170.405 ;
        RECT 93.520 169.555 94.475 169.775 ;
        RECT 92.025 168.775 92.545 169.315 ;
        RECT 92.715 168.605 93.235 169.145 ;
        RECT 93.405 168.825 94.095 169.385 ;
        RECT 94.265 168.655 94.475 169.555 ;
        RECT 90.735 168.025 90.905 168.405 ;
        RECT 91.085 167.855 91.415 168.235 ;
        RECT 91.595 168.025 91.855 168.530 ;
        RECT 92.025 167.855 93.235 168.605 ;
        RECT 93.520 168.485 94.475 168.655 ;
        RECT 94.645 169.385 95.045 170.235 ;
        RECT 95.235 169.775 95.515 170.235 ;
        RECT 96.035 169.945 96.360 170.405 ;
        RECT 95.235 169.555 96.360 169.775 ;
        RECT 94.645 168.825 95.740 169.385 ;
        RECT 95.910 169.095 96.360 169.555 ;
        RECT 96.530 169.265 96.915 170.235 ;
        RECT 93.520 168.025 93.805 168.485 ;
        RECT 93.975 167.855 94.245 168.315 ;
        RECT 94.645 168.025 95.045 168.825 ;
        RECT 95.910 168.765 96.465 169.095 ;
        RECT 95.910 168.655 96.360 168.765 ;
        RECT 95.235 168.485 96.360 168.655 ;
        RECT 96.635 168.595 96.915 169.265 ;
        RECT 97.085 169.645 97.600 170.055 ;
        RECT 97.835 169.645 98.005 170.405 ;
        RECT 98.175 170.065 100.205 170.235 ;
        RECT 97.085 168.835 97.425 169.645 ;
        RECT 98.175 169.400 98.345 170.065 ;
        RECT 98.740 169.725 99.865 169.895 ;
        RECT 97.595 169.210 98.345 169.400 ;
        RECT 98.515 169.385 99.525 169.555 ;
        RECT 97.085 168.665 98.315 168.835 ;
        RECT 95.235 168.025 95.515 168.485 ;
        RECT 96.035 167.855 96.360 168.315 ;
        RECT 96.530 168.025 96.915 168.595 ;
        RECT 97.360 168.060 97.605 168.665 ;
        RECT 97.825 167.855 98.335 168.390 ;
        RECT 98.515 168.025 98.705 169.385 ;
        RECT 98.875 168.365 99.150 169.185 ;
        RECT 99.355 168.585 99.525 169.385 ;
        RECT 99.695 168.595 99.865 169.725 ;
        RECT 100.035 169.095 100.205 170.065 ;
        RECT 100.375 169.265 100.545 170.405 ;
        RECT 100.715 169.265 101.050 170.235 ;
        RECT 100.035 168.765 100.230 169.095 ;
        RECT 100.455 168.765 100.710 169.095 ;
        RECT 100.455 168.595 100.625 168.765 ;
        RECT 100.880 168.595 101.050 169.265 ;
        RECT 101.685 169.240 101.975 170.405 ;
        RECT 102.145 169.315 103.355 170.405 ;
        RECT 103.525 169.645 104.040 170.055 ;
        RECT 104.275 169.645 104.445 170.405 ;
        RECT 104.615 170.065 106.645 170.235 ;
        RECT 102.145 168.775 102.665 169.315 ;
        RECT 102.835 168.605 103.355 169.145 ;
        RECT 103.525 168.835 103.865 169.645 ;
        RECT 104.615 169.400 104.785 170.065 ;
        RECT 105.180 169.725 106.305 169.895 ;
        RECT 104.035 169.210 104.785 169.400 ;
        RECT 104.955 169.385 105.965 169.555 ;
        RECT 103.525 168.665 104.755 168.835 ;
        RECT 99.695 168.425 100.625 168.595 ;
        RECT 99.695 168.390 99.870 168.425 ;
        RECT 98.875 168.195 99.155 168.365 ;
        RECT 98.875 168.025 99.150 168.195 ;
        RECT 99.340 168.025 99.870 168.390 ;
        RECT 100.295 167.855 100.625 168.255 ;
        RECT 100.795 168.025 101.050 168.595 ;
        RECT 101.685 167.855 101.975 168.580 ;
        RECT 102.145 167.855 103.355 168.605 ;
        RECT 103.800 168.060 104.045 168.665 ;
        RECT 104.265 167.855 104.775 168.390 ;
        RECT 104.955 168.025 105.145 169.385 ;
        RECT 105.315 168.705 105.590 169.185 ;
        RECT 105.315 168.535 105.595 168.705 ;
        RECT 105.795 168.585 105.965 169.385 ;
        RECT 106.135 168.595 106.305 169.725 ;
        RECT 106.475 169.095 106.645 170.065 ;
        RECT 106.815 169.265 106.985 170.405 ;
        RECT 107.155 169.265 107.490 170.235 ;
        RECT 106.475 168.765 106.670 169.095 ;
        RECT 106.895 168.765 107.150 169.095 ;
        RECT 106.895 168.595 107.065 168.765 ;
        RECT 107.320 168.595 107.490 169.265 ;
        RECT 107.665 169.315 108.875 170.405 ;
        RECT 109.135 169.475 109.305 170.235 ;
        RECT 109.485 169.645 109.815 170.405 ;
        RECT 107.665 168.775 108.185 169.315 ;
        RECT 109.135 169.305 109.800 169.475 ;
        RECT 109.985 169.330 110.255 170.235 ;
        RECT 109.630 169.160 109.800 169.305 ;
        RECT 108.355 168.605 108.875 169.145 ;
        RECT 109.065 168.755 109.395 169.125 ;
        RECT 109.630 168.830 109.915 169.160 ;
        RECT 105.315 168.025 105.590 168.535 ;
        RECT 106.135 168.425 107.065 168.595 ;
        RECT 106.135 168.390 106.310 168.425 ;
        RECT 105.780 168.025 106.310 168.390 ;
        RECT 106.735 167.855 107.065 168.255 ;
        RECT 107.235 168.025 107.490 168.595 ;
        RECT 107.665 167.855 108.875 168.605 ;
        RECT 109.630 168.575 109.800 168.830 ;
        RECT 109.135 168.405 109.800 168.575 ;
        RECT 110.085 168.530 110.255 169.330 ;
        RECT 110.425 169.645 110.940 170.055 ;
        RECT 111.175 169.645 111.345 170.405 ;
        RECT 111.515 170.065 113.545 170.235 ;
        RECT 110.425 168.835 110.765 169.645 ;
        RECT 111.515 169.400 111.685 170.065 ;
        RECT 112.080 169.725 113.205 169.895 ;
        RECT 110.935 169.210 111.685 169.400 ;
        RECT 111.855 169.385 112.865 169.555 ;
        RECT 110.425 168.665 111.655 168.835 ;
        RECT 109.135 168.025 109.305 168.405 ;
        RECT 109.485 167.855 109.815 168.235 ;
        RECT 109.995 168.025 110.255 168.530 ;
        RECT 110.700 168.060 110.945 168.665 ;
        RECT 111.165 167.855 111.675 168.390 ;
        RECT 111.855 168.025 112.045 169.385 ;
        RECT 112.215 169.045 112.490 169.185 ;
        RECT 112.215 168.875 112.495 169.045 ;
        RECT 112.215 168.025 112.490 168.875 ;
        RECT 112.695 168.585 112.865 169.385 ;
        RECT 113.035 168.595 113.205 169.725 ;
        RECT 113.375 169.095 113.545 170.065 ;
        RECT 113.715 169.265 113.885 170.405 ;
        RECT 114.055 169.265 114.390 170.235 ;
        RECT 113.375 168.765 113.570 169.095 ;
        RECT 113.795 168.765 114.050 169.095 ;
        RECT 113.795 168.595 113.965 168.765 ;
        RECT 114.220 168.595 114.390 169.265 ;
        RECT 115.025 169.315 116.695 170.405 ;
        RECT 115.025 168.795 115.775 169.315 ;
        RECT 116.870 169.215 117.125 170.095 ;
        RECT 117.295 169.265 117.600 170.405 ;
        RECT 117.940 170.025 118.270 170.405 ;
        RECT 118.450 169.855 118.620 170.145 ;
        RECT 118.790 169.945 119.040 170.405 ;
        RECT 117.820 169.685 118.620 169.855 ;
        RECT 119.210 169.895 120.080 170.235 ;
        RECT 115.945 168.625 116.695 169.145 ;
        RECT 113.035 168.425 113.965 168.595 ;
        RECT 113.035 168.390 113.210 168.425 ;
        RECT 112.680 168.025 113.210 168.390 ;
        RECT 113.635 167.855 113.965 168.255 ;
        RECT 114.135 168.025 114.390 168.595 ;
        RECT 115.025 167.855 116.695 168.625 ;
        RECT 116.870 168.565 117.080 169.215 ;
        RECT 117.820 169.095 117.990 169.685 ;
        RECT 119.210 169.515 119.380 169.895 ;
        RECT 120.315 169.775 120.485 170.235 ;
        RECT 120.655 169.945 121.025 170.405 ;
        RECT 121.320 169.805 121.490 170.145 ;
        RECT 121.660 169.975 121.990 170.405 ;
        RECT 122.225 169.805 122.395 170.145 ;
        RECT 118.160 169.345 119.380 169.515 ;
        RECT 119.550 169.435 120.010 169.725 ;
        RECT 120.315 169.605 120.875 169.775 ;
        RECT 121.320 169.635 122.395 169.805 ;
        RECT 122.565 169.905 123.245 170.235 ;
        RECT 123.460 169.905 123.710 170.235 ;
        RECT 123.880 169.945 124.130 170.405 ;
        RECT 120.705 169.465 120.875 169.605 ;
        RECT 119.550 169.425 120.515 169.435 ;
        RECT 119.210 169.255 119.380 169.345 ;
        RECT 119.840 169.265 120.515 169.425 ;
        RECT 117.250 169.065 117.990 169.095 ;
        RECT 117.250 168.765 118.165 169.065 ;
        RECT 117.840 168.590 118.165 168.765 ;
        RECT 116.870 168.035 117.125 168.565 ;
        RECT 117.295 167.855 117.600 168.315 ;
        RECT 117.845 168.235 118.165 168.590 ;
        RECT 118.335 168.805 118.875 169.175 ;
        RECT 119.210 169.085 119.615 169.255 ;
        RECT 118.335 168.405 118.575 168.805 ;
        RECT 119.055 168.635 119.275 168.915 ;
        RECT 118.745 168.465 119.275 168.635 ;
        RECT 118.745 168.235 118.915 168.465 ;
        RECT 119.445 168.305 119.615 169.085 ;
        RECT 119.785 168.475 120.135 169.095 ;
        RECT 120.305 168.475 120.515 169.265 ;
        RECT 120.705 169.295 122.205 169.465 ;
        RECT 120.705 168.605 120.875 169.295 ;
        RECT 122.565 169.125 122.735 169.905 ;
        RECT 123.540 169.775 123.710 169.905 ;
        RECT 121.045 168.955 122.735 169.125 ;
        RECT 122.905 169.345 123.370 169.735 ;
        RECT 123.540 169.605 123.935 169.775 ;
        RECT 121.045 168.775 121.215 168.955 ;
        RECT 117.845 168.065 118.915 168.235 ;
        RECT 119.085 167.855 119.275 168.295 ;
        RECT 119.445 168.025 120.395 168.305 ;
        RECT 120.705 168.215 120.965 168.605 ;
        RECT 121.385 168.535 122.175 168.785 ;
        RECT 120.615 168.045 120.965 168.215 ;
        RECT 121.175 167.855 121.505 168.315 ;
        RECT 122.380 168.245 122.550 168.955 ;
        RECT 122.905 168.755 123.075 169.345 ;
        RECT 122.720 168.535 123.075 168.755 ;
        RECT 123.245 168.535 123.595 169.155 ;
        RECT 123.765 168.245 123.935 169.605 ;
        RECT 124.300 169.435 124.625 170.220 ;
        RECT 124.105 168.385 124.565 169.435 ;
        RECT 122.380 168.075 123.235 168.245 ;
        RECT 123.440 168.075 123.935 168.245 ;
        RECT 124.105 167.855 124.435 168.215 ;
        RECT 124.795 168.115 124.965 170.235 ;
        RECT 125.135 169.905 125.465 170.405 ;
        RECT 125.635 169.735 125.890 170.235 ;
        RECT 125.140 169.565 125.890 169.735 ;
        RECT 125.140 168.575 125.370 169.565 ;
        RECT 125.540 168.745 125.890 169.395 ;
        RECT 126.525 169.315 127.735 170.405 ;
        RECT 126.525 168.775 127.045 169.315 ;
        RECT 127.215 168.605 127.735 169.145 ;
        RECT 125.140 168.405 125.890 168.575 ;
        RECT 125.135 167.855 125.465 168.235 ;
        RECT 125.635 168.115 125.890 168.405 ;
        RECT 126.525 167.855 127.735 168.605 ;
        RECT 29.840 167.685 127.820 167.855 ;
        RECT 29.925 166.935 31.135 167.685 ;
        RECT 29.925 166.395 30.445 166.935 ;
        RECT 31.765 166.915 34.355 167.685 ;
        RECT 30.615 166.225 31.135 166.765 ;
        RECT 29.925 165.135 31.135 166.225 ;
        RECT 31.765 166.225 32.975 166.745 ;
        RECT 33.145 166.395 34.355 166.915 ;
        RECT 34.585 166.865 34.795 167.685 ;
        RECT 34.965 166.885 35.295 167.515 ;
        RECT 34.965 166.285 35.215 166.885 ;
        RECT 35.465 166.865 35.695 167.685 ;
        RECT 35.905 166.935 37.115 167.685 ;
        RECT 37.285 166.960 37.575 167.685 ;
        RECT 37.835 167.135 38.005 167.515 ;
        RECT 38.185 167.305 38.515 167.685 ;
        RECT 37.835 166.965 38.500 167.135 ;
        RECT 38.695 167.010 38.955 167.515 ;
        RECT 35.385 166.445 35.715 166.695 ;
        RECT 31.765 165.135 34.355 166.225 ;
        RECT 34.585 165.135 34.795 166.275 ;
        RECT 34.965 165.305 35.295 166.285 ;
        RECT 35.465 165.135 35.695 166.275 ;
        RECT 35.905 166.225 36.425 166.765 ;
        RECT 36.595 166.395 37.115 166.935 ;
        RECT 37.765 166.415 38.095 166.785 ;
        RECT 38.330 166.710 38.500 166.965 ;
        RECT 38.330 166.380 38.615 166.710 ;
        RECT 35.905 165.135 37.115 166.225 ;
        RECT 37.285 165.135 37.575 166.300 ;
        RECT 38.330 166.235 38.500 166.380 ;
        RECT 37.835 166.065 38.500 166.235 ;
        RECT 38.785 166.210 38.955 167.010 ;
        RECT 39.125 166.915 42.635 167.685 ;
        RECT 37.835 165.305 38.005 166.065 ;
        RECT 38.185 165.135 38.515 165.895 ;
        RECT 38.685 165.305 38.955 166.210 ;
        RECT 39.125 166.225 40.815 166.745 ;
        RECT 40.985 166.395 42.635 166.915 ;
        RECT 43.010 166.905 43.510 167.515 ;
        RECT 42.805 166.445 43.155 166.695 ;
        RECT 43.340 166.275 43.510 166.905 ;
        RECT 44.140 167.035 44.470 167.515 ;
        RECT 44.640 167.225 44.865 167.685 ;
        RECT 45.035 167.035 45.365 167.515 ;
        RECT 44.140 166.865 45.365 167.035 ;
        RECT 45.555 166.885 45.805 167.685 ;
        RECT 45.975 166.885 46.315 167.515 ;
        RECT 43.680 166.495 44.010 166.695 ;
        RECT 44.180 166.495 44.510 166.695 ;
        RECT 44.680 166.495 45.100 166.695 ;
        RECT 45.275 166.525 45.970 166.695 ;
        RECT 45.275 166.275 45.445 166.525 ;
        RECT 46.140 166.275 46.315 166.885 ;
        RECT 46.760 166.875 47.005 167.480 ;
        RECT 47.225 167.150 47.735 167.685 ;
        RECT 39.125 165.135 42.635 166.225 ;
        RECT 43.010 166.105 45.445 166.275 ;
        RECT 43.010 165.305 43.340 166.105 ;
        RECT 43.510 165.135 43.840 165.935 ;
        RECT 44.140 165.305 44.470 166.105 ;
        RECT 45.115 165.135 45.365 165.935 ;
        RECT 45.635 165.135 45.805 166.275 ;
        RECT 45.975 165.305 46.315 166.275 ;
        RECT 46.485 166.705 47.715 166.875 ;
        RECT 46.485 165.895 46.825 166.705 ;
        RECT 46.995 166.140 47.745 166.330 ;
        RECT 46.485 165.485 47.000 165.895 ;
        RECT 47.235 165.135 47.405 165.895 ;
        RECT 47.575 165.475 47.745 166.140 ;
        RECT 47.915 166.155 48.105 167.515 ;
        RECT 48.275 166.665 48.550 167.515 ;
        RECT 48.740 167.150 49.270 167.515 ;
        RECT 49.695 167.285 50.025 167.685 ;
        RECT 49.095 167.115 49.270 167.150 ;
        RECT 48.275 166.495 48.555 166.665 ;
        RECT 48.275 166.355 48.550 166.495 ;
        RECT 48.755 166.155 48.925 166.955 ;
        RECT 47.915 165.985 48.925 166.155 ;
        RECT 49.095 166.945 50.025 167.115 ;
        RECT 50.195 166.945 50.450 167.515 ;
        RECT 49.095 165.815 49.265 166.945 ;
        RECT 49.855 166.775 50.025 166.945 ;
        RECT 48.140 165.645 49.265 165.815 ;
        RECT 49.435 166.445 49.630 166.775 ;
        RECT 49.855 166.445 50.110 166.775 ;
        RECT 49.435 165.475 49.605 166.445 ;
        RECT 50.280 166.275 50.450 166.945 ;
        RECT 50.665 166.865 50.895 167.685 ;
        RECT 51.065 166.885 51.395 167.515 ;
        RECT 50.645 166.445 50.975 166.695 ;
        RECT 51.145 166.285 51.395 166.885 ;
        RECT 51.565 166.865 51.775 167.685 ;
        RECT 52.210 166.905 52.710 167.515 ;
        RECT 52.005 166.445 52.355 166.695 ;
        RECT 47.575 165.305 49.605 165.475 ;
        RECT 49.775 165.135 49.945 166.275 ;
        RECT 50.115 165.305 50.450 166.275 ;
        RECT 50.665 165.135 50.895 166.275 ;
        RECT 51.065 165.305 51.395 166.285 ;
        RECT 52.540 166.275 52.710 166.905 ;
        RECT 53.340 167.035 53.670 167.515 ;
        RECT 53.840 167.225 54.065 167.685 ;
        RECT 54.235 167.035 54.565 167.515 ;
        RECT 53.340 166.865 54.565 167.035 ;
        RECT 54.755 166.885 55.005 167.685 ;
        RECT 55.175 166.885 55.515 167.515 ;
        RECT 52.880 166.495 53.210 166.695 ;
        RECT 53.380 166.495 53.710 166.695 ;
        RECT 53.880 166.495 54.300 166.695 ;
        RECT 54.475 166.525 55.170 166.695 ;
        RECT 54.475 166.275 54.645 166.525 ;
        RECT 55.340 166.275 55.515 166.885 ;
        RECT 51.565 165.135 51.775 166.275 ;
        RECT 52.210 166.105 54.645 166.275 ;
        RECT 52.210 165.305 52.540 166.105 ;
        RECT 52.710 165.135 53.040 165.935 ;
        RECT 53.340 165.305 53.670 166.105 ;
        RECT 54.315 165.135 54.565 165.935 ;
        RECT 54.835 165.135 55.005 166.275 ;
        RECT 55.175 165.305 55.515 166.275 ;
        RECT 55.690 166.945 55.945 167.515 ;
        RECT 56.115 167.285 56.445 167.685 ;
        RECT 56.870 167.150 57.400 167.515 ;
        RECT 56.870 167.115 57.045 167.150 ;
        RECT 56.115 166.945 57.045 167.115 ;
        RECT 57.590 167.005 57.865 167.515 ;
        RECT 55.690 166.275 55.860 166.945 ;
        RECT 56.115 166.775 56.285 166.945 ;
        RECT 56.030 166.445 56.285 166.775 ;
        RECT 56.510 166.445 56.705 166.775 ;
        RECT 55.690 165.305 56.025 166.275 ;
        RECT 56.195 165.135 56.365 166.275 ;
        RECT 56.535 165.475 56.705 166.445 ;
        RECT 56.875 165.815 57.045 166.945 ;
        RECT 57.215 166.155 57.385 166.955 ;
        RECT 57.585 166.835 57.865 167.005 ;
        RECT 57.590 166.355 57.865 166.835 ;
        RECT 58.035 166.155 58.225 167.515 ;
        RECT 58.405 167.150 58.915 167.685 ;
        RECT 59.135 166.875 59.380 167.480 ;
        RECT 60.285 166.915 62.875 167.685 ;
        RECT 63.045 166.960 63.335 167.685 ;
        RECT 63.505 166.915 65.175 167.685 ;
        RECT 58.425 166.705 59.655 166.875 ;
        RECT 57.215 165.985 58.225 166.155 ;
        RECT 58.395 166.140 59.145 166.330 ;
        RECT 56.875 165.645 58.000 165.815 ;
        RECT 58.395 165.475 58.565 166.140 ;
        RECT 59.315 165.895 59.655 166.705 ;
        RECT 56.535 165.305 58.565 165.475 ;
        RECT 58.735 165.135 58.905 165.895 ;
        RECT 59.140 165.485 59.655 165.895 ;
        RECT 60.285 166.225 61.495 166.745 ;
        RECT 61.665 166.395 62.875 166.915 ;
        RECT 60.285 165.135 62.875 166.225 ;
        RECT 63.045 165.135 63.335 166.300 ;
        RECT 63.505 166.225 64.255 166.745 ;
        RECT 64.425 166.395 65.175 166.915 ;
        RECT 65.350 166.945 65.605 167.515 ;
        RECT 65.775 167.285 66.105 167.685 ;
        RECT 66.530 167.150 67.060 167.515 ;
        RECT 66.530 167.115 66.705 167.150 ;
        RECT 65.775 166.945 66.705 167.115 ;
        RECT 65.350 166.275 65.520 166.945 ;
        RECT 65.775 166.775 65.945 166.945 ;
        RECT 65.690 166.445 65.945 166.775 ;
        RECT 66.170 166.445 66.365 166.775 ;
        RECT 63.505 165.135 65.175 166.225 ;
        RECT 65.350 165.305 65.685 166.275 ;
        RECT 65.855 165.135 66.025 166.275 ;
        RECT 66.195 165.475 66.365 166.445 ;
        RECT 66.535 165.815 66.705 166.945 ;
        RECT 66.875 166.155 67.045 166.955 ;
        RECT 67.250 166.665 67.525 167.515 ;
        RECT 67.245 166.495 67.525 166.665 ;
        RECT 67.250 166.355 67.525 166.495 ;
        RECT 67.695 166.155 67.885 167.515 ;
        RECT 68.065 167.150 68.575 167.685 ;
        RECT 68.795 166.875 69.040 167.480 ;
        RECT 69.760 166.875 70.005 167.480 ;
        RECT 70.225 167.150 70.735 167.685 ;
        RECT 68.085 166.705 69.315 166.875 ;
        RECT 66.875 165.985 67.885 166.155 ;
        RECT 68.055 166.140 68.805 166.330 ;
        RECT 66.535 165.645 67.660 165.815 ;
        RECT 68.055 165.475 68.225 166.140 ;
        RECT 68.975 165.895 69.315 166.705 ;
        RECT 66.195 165.305 68.225 165.475 ;
        RECT 68.395 165.135 68.565 165.895 ;
        RECT 68.800 165.485 69.315 165.895 ;
        RECT 69.485 166.705 70.715 166.875 ;
        RECT 69.485 165.895 69.825 166.705 ;
        RECT 69.995 166.140 70.745 166.330 ;
        RECT 69.485 165.485 70.000 165.895 ;
        RECT 70.235 165.135 70.405 165.895 ;
        RECT 70.575 165.475 70.745 166.140 ;
        RECT 70.915 166.155 71.105 167.515 ;
        RECT 71.275 167.005 71.550 167.515 ;
        RECT 71.740 167.150 72.270 167.515 ;
        RECT 72.695 167.285 73.025 167.685 ;
        RECT 72.095 167.115 72.270 167.150 ;
        RECT 71.275 166.835 71.555 167.005 ;
        RECT 71.275 166.355 71.550 166.835 ;
        RECT 71.755 166.155 71.925 166.955 ;
        RECT 70.915 165.985 71.925 166.155 ;
        RECT 72.095 166.945 73.025 167.115 ;
        RECT 73.195 166.945 73.450 167.515 ;
        RECT 72.095 165.815 72.265 166.945 ;
        RECT 72.855 166.775 73.025 166.945 ;
        RECT 71.140 165.645 72.265 165.815 ;
        RECT 72.435 166.445 72.630 166.775 ;
        RECT 72.855 166.445 73.110 166.775 ;
        RECT 72.435 165.475 72.605 166.445 ;
        RECT 73.280 166.275 73.450 166.945 ;
        RECT 74.235 166.885 74.565 167.685 ;
        RECT 74.735 167.035 74.905 167.515 ;
        RECT 75.075 167.205 75.405 167.685 ;
        RECT 75.575 167.035 75.745 167.515 ;
        RECT 75.995 167.205 76.235 167.685 ;
        RECT 76.415 167.035 76.585 167.515 ;
        RECT 74.735 166.865 75.745 167.035 ;
        RECT 75.950 166.865 76.585 167.035 ;
        RECT 74.735 166.325 75.230 166.865 ;
        RECT 75.950 166.695 76.120 166.865 ;
        RECT 77.310 166.845 77.570 167.685 ;
        RECT 77.745 166.940 78.000 167.515 ;
        RECT 78.170 167.305 78.500 167.685 ;
        RECT 78.715 167.135 78.885 167.515 ;
        RECT 78.170 166.965 78.885 167.135 ;
        RECT 75.620 166.525 76.120 166.695 ;
        RECT 70.575 165.305 72.605 165.475 ;
        RECT 72.775 165.135 72.945 166.275 ;
        RECT 73.115 165.305 73.450 166.275 ;
        RECT 74.235 165.135 74.565 166.285 ;
        RECT 74.735 166.155 75.745 166.325 ;
        RECT 74.735 165.305 74.905 166.155 ;
        RECT 75.075 165.135 75.405 165.935 ;
        RECT 75.575 165.305 75.745 166.155 ;
        RECT 75.950 166.285 76.120 166.525 ;
        RECT 76.290 166.455 76.670 166.695 ;
        RECT 75.950 166.115 76.665 166.285 ;
        RECT 75.925 165.135 76.165 165.935 ;
        RECT 76.335 165.305 76.665 166.115 ;
        RECT 77.310 165.135 77.570 166.285 ;
        RECT 77.745 166.210 77.915 166.940 ;
        RECT 78.170 166.775 78.340 166.965 ;
        RECT 79.145 166.915 80.815 167.685 ;
        RECT 78.085 166.445 78.340 166.775 ;
        RECT 78.170 166.235 78.340 166.445 ;
        RECT 78.620 166.415 78.975 166.785 ;
        RECT 77.745 165.305 78.000 166.210 ;
        RECT 78.170 166.065 78.885 166.235 ;
        RECT 78.170 165.135 78.500 165.895 ;
        RECT 78.715 165.305 78.885 166.065 ;
        RECT 79.145 166.225 79.895 166.745 ;
        RECT 80.065 166.395 80.815 166.915 ;
        RECT 80.985 166.885 81.325 167.515 ;
        RECT 81.495 166.885 81.745 167.685 ;
        RECT 81.935 167.035 82.265 167.515 ;
        RECT 82.435 167.225 82.660 167.685 ;
        RECT 82.830 167.035 83.160 167.515 ;
        RECT 80.985 166.275 81.160 166.885 ;
        RECT 81.935 166.865 83.160 167.035 ;
        RECT 83.790 166.905 84.290 167.515 ;
        RECT 81.330 166.525 82.025 166.695 ;
        RECT 81.855 166.275 82.025 166.525 ;
        RECT 82.200 166.495 82.620 166.695 ;
        RECT 82.790 166.495 83.120 166.695 ;
        RECT 83.290 166.495 83.620 166.695 ;
        RECT 83.790 166.275 83.960 166.905 ;
        RECT 84.940 166.875 85.185 167.480 ;
        RECT 85.405 167.150 85.915 167.685 ;
        RECT 84.665 166.705 85.895 166.875 ;
        RECT 84.145 166.445 84.495 166.695 ;
        RECT 79.145 165.135 80.815 166.225 ;
        RECT 80.985 165.305 81.325 166.275 ;
        RECT 81.495 165.135 81.665 166.275 ;
        RECT 81.855 166.105 84.290 166.275 ;
        RECT 81.935 165.135 82.185 165.935 ;
        RECT 82.830 165.305 83.160 166.105 ;
        RECT 83.460 165.135 83.790 165.935 ;
        RECT 83.960 165.305 84.290 166.105 ;
        RECT 84.665 165.895 85.005 166.705 ;
        RECT 85.175 166.140 85.925 166.330 ;
        RECT 84.665 165.485 85.180 165.895 ;
        RECT 85.415 165.135 85.585 165.895 ;
        RECT 85.755 165.475 85.925 166.140 ;
        RECT 86.095 166.155 86.285 167.515 ;
        RECT 86.455 166.665 86.730 167.515 ;
        RECT 86.920 167.150 87.450 167.515 ;
        RECT 87.875 167.285 88.205 167.685 ;
        RECT 87.275 167.115 87.450 167.150 ;
        RECT 86.455 166.495 86.735 166.665 ;
        RECT 86.455 166.355 86.730 166.495 ;
        RECT 86.935 166.155 87.105 166.955 ;
        RECT 86.095 165.985 87.105 166.155 ;
        RECT 87.275 166.945 88.205 167.115 ;
        RECT 88.375 166.945 88.630 167.515 ;
        RECT 88.805 166.960 89.095 167.685 ;
        RECT 87.275 165.815 87.445 166.945 ;
        RECT 88.035 166.775 88.205 166.945 ;
        RECT 86.320 165.645 87.445 165.815 ;
        RECT 87.615 166.445 87.810 166.775 ;
        RECT 88.035 166.445 88.290 166.775 ;
        RECT 87.615 165.475 87.785 166.445 ;
        RECT 88.460 166.275 88.630 166.945 ;
        RECT 90.245 166.865 90.455 167.685 ;
        RECT 90.625 166.885 90.955 167.515 ;
        RECT 85.755 165.305 87.785 165.475 ;
        RECT 87.955 165.135 88.125 166.275 ;
        RECT 88.295 165.305 88.630 166.275 ;
        RECT 88.805 165.135 89.095 166.300 ;
        RECT 90.625 166.285 90.875 166.885 ;
        RECT 91.125 166.865 91.355 167.685 ;
        RECT 91.655 167.135 91.825 167.515 ;
        RECT 92.005 167.305 92.335 167.685 ;
        RECT 91.655 166.965 92.320 167.135 ;
        RECT 92.515 167.010 92.775 167.515 ;
        RECT 91.045 166.445 91.375 166.695 ;
        RECT 91.585 166.415 91.915 166.785 ;
        RECT 92.150 166.710 92.320 166.965 ;
        RECT 92.150 166.380 92.435 166.710 ;
        RECT 90.245 165.135 90.455 166.275 ;
        RECT 90.625 165.305 90.955 166.285 ;
        RECT 91.125 165.135 91.355 166.275 ;
        RECT 92.150 166.235 92.320 166.380 ;
        RECT 91.655 166.065 92.320 166.235 ;
        RECT 92.605 166.210 92.775 167.010 ;
        RECT 91.655 165.305 91.825 166.065 ;
        RECT 92.005 165.135 92.335 165.895 ;
        RECT 92.505 165.305 92.775 166.210 ;
        RECT 93.780 166.975 94.035 167.505 ;
        RECT 94.215 167.225 94.500 167.685 ;
        RECT 93.780 166.115 93.960 166.975 ;
        RECT 94.680 166.775 94.930 167.425 ;
        RECT 94.130 166.445 94.930 166.775 ;
        RECT 93.780 165.985 94.035 166.115 ;
        RECT 93.695 165.815 94.035 165.985 ;
        RECT 93.780 165.445 94.035 165.815 ;
        RECT 94.215 165.135 94.500 165.935 ;
        RECT 94.680 165.855 94.930 166.445 ;
        RECT 95.130 167.090 95.450 167.420 ;
        RECT 95.630 167.205 96.290 167.685 ;
        RECT 96.490 167.295 97.340 167.465 ;
        RECT 95.130 166.195 95.320 167.090 ;
        RECT 95.640 166.765 96.300 167.035 ;
        RECT 95.970 166.705 96.300 166.765 ;
        RECT 95.490 166.535 95.820 166.595 ;
        RECT 96.490 166.535 96.660 167.295 ;
        RECT 97.900 167.225 98.220 167.685 ;
        RECT 98.420 167.045 98.670 167.475 ;
        RECT 98.960 167.245 99.370 167.685 ;
        RECT 99.540 167.305 100.555 167.505 ;
        RECT 96.830 166.875 98.080 167.045 ;
        RECT 96.830 166.755 97.160 166.875 ;
        RECT 95.490 166.365 97.390 166.535 ;
        RECT 95.130 166.025 97.050 166.195 ;
        RECT 95.130 166.005 95.450 166.025 ;
        RECT 94.680 165.345 95.010 165.855 ;
        RECT 95.280 165.395 95.450 166.005 ;
        RECT 97.220 165.855 97.390 166.365 ;
        RECT 97.560 166.295 97.740 166.705 ;
        RECT 97.910 166.115 98.080 166.875 ;
        RECT 95.620 165.135 95.950 165.825 ;
        RECT 96.180 165.685 97.390 165.855 ;
        RECT 97.560 165.805 98.080 166.115 ;
        RECT 98.250 166.705 98.670 167.045 ;
        RECT 98.960 166.705 99.370 167.035 ;
        RECT 98.250 165.935 98.440 166.705 ;
        RECT 99.540 166.575 99.710 167.305 ;
        RECT 100.855 167.135 101.025 167.465 ;
        RECT 101.195 167.305 101.525 167.685 ;
        RECT 99.880 166.755 100.230 167.125 ;
        RECT 99.540 166.535 99.960 166.575 ;
        RECT 98.610 166.365 99.960 166.535 ;
        RECT 98.610 166.205 98.860 166.365 ;
        RECT 99.370 165.935 99.620 166.195 ;
        RECT 98.250 165.685 99.620 165.935 ;
        RECT 96.180 165.395 96.420 165.685 ;
        RECT 97.220 165.605 97.390 165.685 ;
        RECT 96.620 165.135 97.040 165.515 ;
        RECT 97.220 165.355 97.850 165.605 ;
        RECT 98.320 165.135 98.650 165.515 ;
        RECT 98.820 165.395 98.990 165.685 ;
        RECT 99.790 165.520 99.960 166.365 ;
        RECT 100.410 166.195 100.630 167.065 ;
        RECT 100.855 166.945 101.550 167.135 ;
        RECT 100.130 165.815 100.630 166.195 ;
        RECT 100.800 166.145 101.210 166.765 ;
        RECT 101.380 165.975 101.550 166.945 ;
        RECT 100.855 165.805 101.550 165.975 ;
        RECT 99.170 165.135 99.550 165.515 ;
        RECT 99.790 165.350 100.620 165.520 ;
        RECT 100.855 165.305 101.025 165.805 ;
        RECT 101.195 165.135 101.525 165.635 ;
        RECT 101.740 165.305 101.965 167.425 ;
        RECT 102.135 167.305 102.465 167.685 ;
        RECT 102.635 167.135 102.805 167.425 ;
        RECT 102.140 166.965 102.805 167.135 ;
        RECT 103.065 167.010 103.325 167.515 ;
        RECT 103.505 167.305 103.835 167.685 ;
        RECT 104.015 167.135 104.185 167.515 ;
        RECT 102.140 165.975 102.370 166.965 ;
        RECT 102.540 166.145 102.890 166.795 ;
        RECT 103.065 166.210 103.235 167.010 ;
        RECT 103.520 166.965 104.185 167.135 ;
        RECT 103.520 166.710 103.690 166.965 ;
        RECT 104.905 166.915 106.575 167.685 ;
        RECT 103.405 166.380 103.690 166.710 ;
        RECT 103.925 166.415 104.255 166.785 ;
        RECT 103.520 166.235 103.690 166.380 ;
        RECT 102.140 165.805 102.805 165.975 ;
        RECT 102.135 165.135 102.465 165.635 ;
        RECT 102.635 165.305 102.805 165.805 ;
        RECT 103.065 165.305 103.335 166.210 ;
        RECT 103.520 166.065 104.185 166.235 ;
        RECT 103.505 165.135 103.835 165.895 ;
        RECT 104.015 165.305 104.185 166.065 ;
        RECT 104.905 166.225 105.655 166.745 ;
        RECT 105.825 166.395 106.575 166.915 ;
        RECT 106.745 167.010 107.015 167.355 ;
        RECT 107.205 167.285 107.585 167.685 ;
        RECT 107.755 167.115 107.925 167.465 ;
        RECT 108.095 167.285 108.425 167.685 ;
        RECT 108.625 167.115 108.795 167.465 ;
        RECT 108.995 167.185 109.325 167.685 ;
        RECT 106.745 166.275 106.915 167.010 ;
        RECT 107.185 166.945 108.795 167.115 ;
        RECT 107.185 166.775 107.355 166.945 ;
        RECT 107.085 166.445 107.355 166.775 ;
        RECT 107.525 166.445 107.930 166.775 ;
        RECT 107.185 166.275 107.355 166.445 ;
        RECT 104.905 165.135 106.575 166.225 ;
        RECT 106.745 165.305 107.015 166.275 ;
        RECT 107.185 166.105 107.910 166.275 ;
        RECT 108.100 166.155 108.810 166.775 ;
        RECT 108.980 166.445 109.330 167.015 ;
        RECT 109.505 166.885 109.845 167.515 ;
        RECT 110.015 166.885 110.265 167.685 ;
        RECT 110.455 167.035 110.785 167.515 ;
        RECT 110.955 167.225 111.180 167.685 ;
        RECT 111.350 167.035 111.680 167.515 ;
        RECT 109.505 166.275 109.680 166.885 ;
        RECT 110.455 166.865 111.680 167.035 ;
        RECT 112.310 166.905 112.810 167.515 ;
        RECT 113.185 166.935 114.395 167.685 ;
        RECT 114.565 166.960 114.855 167.685 ;
        RECT 115.140 167.055 115.425 167.515 ;
        RECT 115.595 167.225 115.865 167.685 ;
        RECT 109.850 166.525 110.545 166.695 ;
        RECT 110.375 166.275 110.545 166.525 ;
        RECT 110.720 166.495 111.140 166.695 ;
        RECT 111.310 166.495 111.640 166.695 ;
        RECT 111.810 166.495 112.140 166.695 ;
        RECT 112.310 166.275 112.480 166.905 ;
        RECT 112.665 166.445 113.015 166.695 ;
        RECT 107.740 165.985 107.910 166.105 ;
        RECT 109.010 165.985 109.330 166.275 ;
        RECT 107.225 165.135 107.505 165.935 ;
        RECT 107.740 165.815 109.330 165.985 ;
        RECT 107.675 165.355 109.330 165.645 ;
        RECT 109.505 165.305 109.845 166.275 ;
        RECT 110.015 165.135 110.185 166.275 ;
        RECT 110.375 166.105 112.810 166.275 ;
        RECT 110.455 165.135 110.705 165.935 ;
        RECT 111.350 165.305 111.680 166.105 ;
        RECT 111.980 165.135 112.310 165.935 ;
        RECT 112.480 165.305 112.810 166.105 ;
        RECT 113.185 166.225 113.705 166.765 ;
        RECT 113.875 166.395 114.395 166.935 ;
        RECT 115.140 166.885 116.095 167.055 ;
        RECT 113.185 165.135 114.395 166.225 ;
        RECT 114.565 165.135 114.855 166.300 ;
        RECT 115.025 166.155 115.715 166.715 ;
        RECT 115.885 165.985 116.095 166.885 ;
        RECT 115.140 165.765 116.095 165.985 ;
        RECT 116.265 166.715 116.665 167.515 ;
        RECT 116.855 167.055 117.135 167.515 ;
        RECT 117.655 167.225 117.980 167.685 ;
        RECT 116.855 166.885 117.980 167.055 ;
        RECT 118.150 166.945 118.535 167.515 ;
        RECT 117.530 166.775 117.980 166.885 ;
        RECT 116.265 166.155 117.360 166.715 ;
        RECT 117.530 166.445 118.085 166.775 ;
        RECT 115.140 165.305 115.425 165.765 ;
        RECT 115.595 165.135 115.865 165.595 ;
        RECT 116.265 165.305 116.665 166.155 ;
        RECT 117.530 165.985 117.980 166.445 ;
        RECT 118.255 166.275 118.535 166.945 ;
        RECT 118.855 166.885 119.185 167.685 ;
        RECT 119.355 167.035 119.525 167.515 ;
        RECT 119.695 167.205 120.025 167.685 ;
        RECT 120.195 167.035 120.365 167.515 ;
        RECT 120.615 167.205 120.855 167.685 ;
        RECT 121.035 167.035 121.205 167.515 ;
        RECT 119.355 166.865 120.365 167.035 ;
        RECT 120.570 166.865 121.205 167.035 ;
        RECT 121.615 166.885 121.945 167.685 ;
        RECT 122.115 167.035 122.285 167.515 ;
        RECT 122.455 167.205 122.785 167.685 ;
        RECT 122.955 167.035 123.125 167.515 ;
        RECT 123.375 167.205 123.615 167.685 ;
        RECT 123.795 167.035 123.965 167.515 ;
        RECT 122.115 166.865 123.125 167.035 ;
        RECT 123.330 166.865 123.965 167.035 ;
        RECT 124.685 166.915 126.355 167.685 ;
        RECT 126.525 166.935 127.735 167.685 ;
        RECT 119.355 166.325 119.850 166.865 ;
        RECT 120.570 166.695 120.740 166.865 ;
        RECT 120.240 166.525 120.740 166.695 ;
        RECT 116.855 165.765 117.980 165.985 ;
        RECT 116.855 165.305 117.135 165.765 ;
        RECT 117.655 165.135 117.980 165.595 ;
        RECT 118.150 165.305 118.535 166.275 ;
        RECT 118.855 165.135 119.185 166.285 ;
        RECT 119.355 166.155 120.365 166.325 ;
        RECT 119.355 165.305 119.525 166.155 ;
        RECT 119.695 165.135 120.025 165.935 ;
        RECT 120.195 165.305 120.365 166.155 ;
        RECT 120.570 166.285 120.740 166.525 ;
        RECT 120.910 166.455 121.290 166.695 ;
        RECT 122.115 166.325 122.610 166.865 ;
        RECT 123.330 166.695 123.500 166.865 ;
        RECT 123.000 166.525 123.500 166.695 ;
        RECT 120.570 166.115 121.285 166.285 ;
        RECT 120.545 165.135 120.785 165.935 ;
        RECT 120.955 165.305 121.285 166.115 ;
        RECT 121.615 165.135 121.945 166.285 ;
        RECT 122.115 166.155 123.125 166.325 ;
        RECT 122.115 165.305 122.285 166.155 ;
        RECT 122.455 165.135 122.785 165.935 ;
        RECT 122.955 165.305 123.125 166.155 ;
        RECT 123.330 166.285 123.500 166.525 ;
        RECT 123.670 166.455 124.050 166.695 ;
        RECT 123.330 166.115 124.045 166.285 ;
        RECT 123.305 165.135 123.545 165.935 ;
        RECT 123.715 165.305 124.045 166.115 ;
        RECT 124.685 166.225 125.435 166.745 ;
        RECT 125.605 166.395 126.355 166.915 ;
        RECT 126.525 166.225 127.045 166.765 ;
        RECT 127.215 166.395 127.735 166.935 ;
        RECT 124.685 165.135 126.355 166.225 ;
        RECT 126.525 165.135 127.735 166.225 ;
        RECT 29.840 164.965 127.820 165.135 ;
        RECT 29.925 163.875 31.135 164.965 ;
        RECT 29.925 163.165 30.445 163.705 ;
        RECT 30.615 163.335 31.135 163.875 ;
        RECT 32.225 164.205 32.740 164.615 ;
        RECT 32.975 164.205 33.145 164.965 ;
        RECT 33.315 164.625 35.345 164.795 ;
        RECT 32.225 163.395 32.565 164.205 ;
        RECT 33.315 163.960 33.485 164.625 ;
        RECT 33.880 164.285 35.005 164.455 ;
        RECT 32.735 163.770 33.485 163.960 ;
        RECT 33.655 163.945 34.665 164.115 ;
        RECT 32.225 163.225 33.455 163.395 ;
        RECT 29.925 162.415 31.135 163.165 ;
        RECT 32.500 162.620 32.745 163.225 ;
        RECT 32.965 162.415 33.475 162.950 ;
        RECT 33.655 162.585 33.845 163.945 ;
        RECT 34.015 162.925 34.290 163.745 ;
        RECT 34.495 163.145 34.665 163.945 ;
        RECT 34.835 163.155 35.005 164.285 ;
        RECT 35.175 163.655 35.345 164.625 ;
        RECT 35.515 163.825 35.685 164.965 ;
        RECT 35.855 163.825 36.190 164.795 ;
        RECT 35.175 163.325 35.370 163.655 ;
        RECT 35.595 163.325 35.850 163.655 ;
        RECT 35.595 163.155 35.765 163.325 ;
        RECT 36.020 163.155 36.190 163.825 ;
        RECT 36.365 164.205 36.880 164.615 ;
        RECT 37.115 164.205 37.285 164.965 ;
        RECT 37.455 164.625 39.485 164.795 ;
        RECT 36.365 163.395 36.705 164.205 ;
        RECT 37.455 163.960 37.625 164.625 ;
        RECT 38.020 164.285 39.145 164.455 ;
        RECT 36.875 163.770 37.625 163.960 ;
        RECT 37.795 163.945 38.805 164.115 ;
        RECT 36.365 163.225 37.595 163.395 ;
        RECT 34.835 162.985 35.765 163.155 ;
        RECT 34.835 162.950 35.010 162.985 ;
        RECT 34.015 162.755 34.295 162.925 ;
        RECT 34.015 162.585 34.290 162.755 ;
        RECT 34.480 162.585 35.010 162.950 ;
        RECT 35.435 162.415 35.765 162.815 ;
        RECT 35.935 162.585 36.190 163.155 ;
        RECT 36.640 162.620 36.885 163.225 ;
        RECT 37.105 162.415 37.615 162.950 ;
        RECT 37.795 162.585 37.985 163.945 ;
        RECT 38.155 163.265 38.430 163.745 ;
        RECT 38.155 163.095 38.435 163.265 ;
        RECT 38.635 163.145 38.805 163.945 ;
        RECT 38.975 163.155 39.145 164.285 ;
        RECT 39.315 163.655 39.485 164.625 ;
        RECT 39.655 163.825 39.825 164.965 ;
        RECT 39.995 163.825 40.330 164.795 ;
        RECT 39.315 163.325 39.510 163.655 ;
        RECT 39.735 163.325 39.990 163.655 ;
        RECT 39.735 163.155 39.905 163.325 ;
        RECT 40.160 163.155 40.330 163.825 ;
        RECT 38.155 162.585 38.430 163.095 ;
        RECT 38.975 162.985 39.905 163.155 ;
        RECT 38.975 162.950 39.150 162.985 ;
        RECT 38.620 162.585 39.150 162.950 ;
        RECT 39.575 162.415 39.905 162.815 ;
        RECT 40.075 162.585 40.330 163.155 ;
        RECT 40.880 163.985 41.135 164.655 ;
        RECT 41.315 164.165 41.600 164.965 ;
        RECT 41.780 164.245 42.110 164.755 ;
        RECT 40.880 163.125 41.060 163.985 ;
        RECT 41.780 163.655 42.030 164.245 ;
        RECT 42.380 164.095 42.550 164.705 ;
        RECT 42.720 164.275 43.050 164.965 ;
        RECT 43.280 164.415 43.520 164.705 ;
        RECT 43.720 164.585 44.140 164.965 ;
        RECT 44.320 164.495 44.950 164.745 ;
        RECT 45.420 164.585 45.750 164.965 ;
        RECT 44.320 164.415 44.490 164.495 ;
        RECT 45.920 164.415 46.090 164.705 ;
        RECT 46.270 164.585 46.650 164.965 ;
        RECT 46.890 164.580 47.720 164.750 ;
        RECT 43.280 164.245 44.490 164.415 ;
        RECT 41.230 163.325 42.030 163.655 ;
        RECT 40.880 162.925 41.135 163.125 ;
        RECT 40.795 162.755 41.135 162.925 ;
        RECT 40.880 162.595 41.135 162.755 ;
        RECT 41.315 162.415 41.600 162.875 ;
        RECT 41.780 162.675 42.030 163.325 ;
        RECT 42.230 164.075 42.550 164.095 ;
        RECT 42.230 163.905 44.150 164.075 ;
        RECT 42.230 163.010 42.420 163.905 ;
        RECT 44.320 163.735 44.490 164.245 ;
        RECT 44.660 163.985 45.180 164.295 ;
        RECT 42.590 163.565 44.490 163.735 ;
        RECT 42.590 163.505 42.920 163.565 ;
        RECT 43.070 163.335 43.400 163.395 ;
        RECT 42.740 163.065 43.400 163.335 ;
        RECT 42.230 162.680 42.550 163.010 ;
        RECT 42.730 162.415 43.390 162.895 ;
        RECT 43.590 162.805 43.760 163.565 ;
        RECT 44.660 163.395 44.840 163.805 ;
        RECT 43.930 163.225 44.260 163.345 ;
        RECT 45.010 163.225 45.180 163.985 ;
        RECT 43.930 163.055 45.180 163.225 ;
        RECT 45.350 164.165 46.720 164.415 ;
        RECT 45.350 163.395 45.540 164.165 ;
        RECT 46.470 163.905 46.720 164.165 ;
        RECT 45.710 163.735 45.960 163.895 ;
        RECT 46.890 163.735 47.060 164.580 ;
        RECT 47.955 164.295 48.125 164.795 ;
        RECT 48.295 164.465 48.625 164.965 ;
        RECT 47.230 163.905 47.730 164.285 ;
        RECT 47.955 164.125 48.650 164.295 ;
        RECT 45.710 163.565 47.060 163.735 ;
        RECT 46.640 163.525 47.060 163.565 ;
        RECT 45.350 163.055 45.770 163.395 ;
        RECT 46.060 163.065 46.470 163.395 ;
        RECT 43.590 162.635 44.440 162.805 ;
        RECT 45.000 162.415 45.320 162.875 ;
        RECT 45.520 162.625 45.770 163.055 ;
        RECT 46.060 162.415 46.470 162.855 ;
        RECT 46.640 162.795 46.810 163.525 ;
        RECT 46.980 162.975 47.330 163.345 ;
        RECT 47.510 163.035 47.730 163.905 ;
        RECT 47.900 163.335 48.310 163.955 ;
        RECT 48.480 163.155 48.650 164.125 ;
        RECT 47.955 162.965 48.650 163.155 ;
        RECT 46.640 162.595 47.655 162.795 ;
        RECT 47.955 162.635 48.125 162.965 ;
        RECT 48.295 162.415 48.625 162.795 ;
        RECT 48.840 162.675 49.065 164.795 ;
        RECT 49.235 164.465 49.565 164.965 ;
        RECT 49.735 164.295 49.905 164.795 ;
        RECT 49.240 164.125 49.905 164.295 ;
        RECT 49.240 163.135 49.470 164.125 ;
        RECT 49.640 163.305 49.990 163.955 ;
        RECT 50.165 163.800 50.455 164.965 ;
        RECT 51.000 164.625 51.255 164.655 ;
        RECT 50.915 164.455 51.255 164.625 ;
        RECT 51.000 163.985 51.255 164.455 ;
        RECT 51.435 164.165 51.720 164.965 ;
        RECT 51.900 164.245 52.230 164.755 ;
        RECT 49.240 162.965 49.905 163.135 ;
        RECT 49.235 162.415 49.565 162.795 ;
        RECT 49.735 162.675 49.905 162.965 ;
        RECT 50.165 162.415 50.455 163.140 ;
        RECT 51.000 163.125 51.180 163.985 ;
        RECT 51.900 163.655 52.150 164.245 ;
        RECT 52.500 164.095 52.670 164.705 ;
        RECT 52.840 164.275 53.170 164.965 ;
        RECT 53.400 164.415 53.640 164.705 ;
        RECT 53.840 164.585 54.260 164.965 ;
        RECT 54.440 164.495 55.070 164.745 ;
        RECT 55.540 164.585 55.870 164.965 ;
        RECT 54.440 164.415 54.610 164.495 ;
        RECT 56.040 164.415 56.210 164.705 ;
        RECT 56.390 164.585 56.770 164.965 ;
        RECT 57.010 164.580 57.840 164.750 ;
        RECT 53.400 164.245 54.610 164.415 ;
        RECT 51.350 163.325 52.150 163.655 ;
        RECT 51.000 162.595 51.255 163.125 ;
        RECT 51.435 162.415 51.720 162.875 ;
        RECT 51.900 162.675 52.150 163.325 ;
        RECT 52.350 164.075 52.670 164.095 ;
        RECT 52.350 163.905 54.270 164.075 ;
        RECT 52.350 163.010 52.540 163.905 ;
        RECT 54.440 163.735 54.610 164.245 ;
        RECT 54.780 163.985 55.300 164.295 ;
        RECT 52.710 163.565 54.610 163.735 ;
        RECT 52.710 163.505 53.040 163.565 ;
        RECT 53.190 163.335 53.520 163.395 ;
        RECT 52.860 163.065 53.520 163.335 ;
        RECT 52.350 162.680 52.670 163.010 ;
        RECT 52.850 162.415 53.510 162.895 ;
        RECT 53.710 162.805 53.880 163.565 ;
        RECT 54.780 163.395 54.960 163.805 ;
        RECT 54.050 163.225 54.380 163.345 ;
        RECT 55.130 163.225 55.300 163.985 ;
        RECT 54.050 163.055 55.300 163.225 ;
        RECT 55.470 164.165 56.840 164.415 ;
        RECT 55.470 163.395 55.660 164.165 ;
        RECT 56.590 163.905 56.840 164.165 ;
        RECT 55.830 163.735 56.080 163.895 ;
        RECT 57.010 163.735 57.180 164.580 ;
        RECT 58.075 164.295 58.245 164.795 ;
        RECT 58.415 164.465 58.745 164.965 ;
        RECT 57.350 163.905 57.850 164.285 ;
        RECT 58.075 164.125 58.770 164.295 ;
        RECT 55.830 163.565 57.180 163.735 ;
        RECT 56.760 163.525 57.180 163.565 ;
        RECT 55.470 163.055 55.890 163.395 ;
        RECT 56.180 163.065 56.590 163.395 ;
        RECT 53.710 162.635 54.560 162.805 ;
        RECT 55.120 162.415 55.440 162.875 ;
        RECT 55.640 162.625 55.890 163.055 ;
        RECT 56.180 162.415 56.590 162.855 ;
        RECT 56.760 162.795 56.930 163.525 ;
        RECT 57.100 162.975 57.450 163.345 ;
        RECT 57.630 163.035 57.850 163.905 ;
        RECT 58.020 163.335 58.430 163.955 ;
        RECT 58.600 163.155 58.770 164.125 ;
        RECT 58.075 162.965 58.770 163.155 ;
        RECT 56.760 162.595 57.775 162.795 ;
        RECT 58.075 162.635 58.245 162.965 ;
        RECT 58.415 162.415 58.745 162.795 ;
        RECT 58.960 162.675 59.185 164.795 ;
        RECT 59.355 164.465 59.685 164.965 ;
        RECT 59.855 164.295 60.025 164.795 ;
        RECT 59.360 164.125 60.025 164.295 ;
        RECT 60.400 164.335 60.685 164.795 ;
        RECT 60.855 164.505 61.125 164.965 ;
        RECT 59.360 163.135 59.590 164.125 ;
        RECT 60.400 164.115 61.355 164.335 ;
        RECT 59.760 163.305 60.110 163.955 ;
        RECT 60.285 163.385 60.975 163.945 ;
        RECT 61.145 163.215 61.355 164.115 ;
        RECT 59.360 162.965 60.025 163.135 ;
        RECT 59.355 162.415 59.685 162.795 ;
        RECT 59.855 162.675 60.025 162.965 ;
        RECT 60.400 163.045 61.355 163.215 ;
        RECT 61.525 163.945 61.925 164.795 ;
        RECT 62.115 164.335 62.395 164.795 ;
        RECT 62.915 164.505 63.240 164.965 ;
        RECT 62.115 164.115 63.240 164.335 ;
        RECT 61.525 163.385 62.620 163.945 ;
        RECT 62.790 163.655 63.240 164.115 ;
        RECT 63.410 163.825 63.795 164.795 ;
        RECT 60.400 162.585 60.685 163.045 ;
        RECT 60.855 162.415 61.125 162.875 ;
        RECT 61.525 162.585 61.925 163.385 ;
        RECT 62.790 163.325 63.345 163.655 ;
        RECT 62.790 163.215 63.240 163.325 ;
        RECT 62.115 163.045 63.240 163.215 ;
        RECT 63.515 163.155 63.795 163.825 ;
        RECT 62.115 162.585 62.395 163.045 ;
        RECT 62.915 162.415 63.240 162.875 ;
        RECT 63.410 162.585 63.795 163.155 ;
        RECT 63.965 163.825 64.305 164.795 ;
        RECT 64.475 163.825 64.645 164.965 ;
        RECT 64.915 164.165 65.165 164.965 ;
        RECT 65.810 163.995 66.140 164.795 ;
        RECT 66.440 164.165 66.770 164.965 ;
        RECT 66.940 163.995 67.270 164.795 ;
        RECT 64.835 163.825 67.270 163.995 ;
        RECT 67.645 163.825 67.985 164.795 ;
        RECT 68.155 163.825 68.325 164.965 ;
        RECT 68.595 164.165 68.845 164.965 ;
        RECT 69.490 163.995 69.820 164.795 ;
        RECT 70.120 164.165 70.450 164.965 ;
        RECT 70.620 163.995 70.950 164.795 ;
        RECT 68.515 163.825 70.950 163.995 ;
        RECT 71.325 163.875 72.535 164.965 ;
        RECT 72.795 164.035 72.965 164.795 ;
        RECT 73.145 164.205 73.475 164.965 ;
        RECT 63.965 163.215 64.140 163.825 ;
        RECT 64.835 163.575 65.005 163.825 ;
        RECT 64.310 163.405 65.005 163.575 ;
        RECT 65.180 163.405 65.600 163.605 ;
        RECT 65.770 163.405 66.100 163.605 ;
        RECT 66.270 163.405 66.600 163.605 ;
        RECT 63.965 162.585 64.305 163.215 ;
        RECT 64.475 162.415 64.725 163.215 ;
        RECT 64.915 163.065 66.140 163.235 ;
        RECT 64.915 162.585 65.245 163.065 ;
        RECT 65.415 162.415 65.640 162.875 ;
        RECT 65.810 162.585 66.140 163.065 ;
        RECT 66.770 163.195 66.940 163.825 ;
        RECT 67.125 163.405 67.475 163.655 ;
        RECT 67.645 163.215 67.820 163.825 ;
        RECT 68.515 163.575 68.685 163.825 ;
        RECT 67.990 163.405 68.685 163.575 ;
        RECT 68.860 163.405 69.280 163.605 ;
        RECT 69.450 163.405 69.780 163.605 ;
        RECT 69.950 163.405 70.280 163.605 ;
        RECT 66.770 162.585 67.270 163.195 ;
        RECT 67.645 162.585 67.985 163.215 ;
        RECT 68.155 162.415 68.405 163.215 ;
        RECT 68.595 163.065 69.820 163.235 ;
        RECT 68.595 162.585 68.925 163.065 ;
        RECT 69.095 162.415 69.320 162.875 ;
        RECT 69.490 162.585 69.820 163.065 ;
        RECT 70.450 163.195 70.620 163.825 ;
        RECT 70.805 163.405 71.155 163.655 ;
        RECT 71.325 163.335 71.845 163.875 ;
        RECT 72.795 163.865 73.460 164.035 ;
        RECT 73.645 163.890 73.915 164.795 ;
        RECT 73.290 163.720 73.460 163.865 ;
        RECT 70.450 162.585 70.950 163.195 ;
        RECT 72.015 163.165 72.535 163.705 ;
        RECT 72.725 163.315 73.055 163.685 ;
        RECT 73.290 163.390 73.575 163.720 ;
        RECT 71.325 162.415 72.535 163.165 ;
        RECT 73.290 163.135 73.460 163.390 ;
        RECT 72.795 162.965 73.460 163.135 ;
        RECT 73.745 163.090 73.915 163.890 ;
        RECT 74.090 163.815 74.350 164.965 ;
        RECT 74.525 163.890 74.780 164.795 ;
        RECT 74.950 164.205 75.280 164.965 ;
        RECT 75.495 164.035 75.665 164.795 ;
        RECT 72.795 162.585 72.965 162.965 ;
        RECT 73.145 162.415 73.475 162.795 ;
        RECT 73.655 162.585 73.915 163.090 ;
        RECT 74.090 162.415 74.350 163.255 ;
        RECT 74.525 163.160 74.695 163.890 ;
        RECT 74.950 163.865 75.665 164.035 ;
        RECT 74.950 163.655 75.120 163.865 ;
        RECT 75.925 163.800 76.215 164.965 ;
        RECT 76.850 163.815 77.110 164.965 ;
        RECT 77.285 163.890 77.540 164.795 ;
        RECT 77.710 164.205 78.040 164.965 ;
        RECT 78.255 164.035 78.425 164.795 ;
        RECT 74.865 163.325 75.120 163.655 ;
        RECT 74.525 162.585 74.780 163.160 ;
        RECT 74.950 163.135 75.120 163.325 ;
        RECT 75.400 163.315 75.755 163.685 ;
        RECT 74.950 162.965 75.665 163.135 ;
        RECT 74.950 162.415 75.280 162.795 ;
        RECT 75.495 162.585 75.665 162.965 ;
        RECT 75.925 162.415 76.215 163.140 ;
        RECT 76.850 162.415 77.110 163.255 ;
        RECT 77.285 163.160 77.455 163.890 ;
        RECT 77.710 163.865 78.425 164.035 ;
        RECT 78.775 164.035 78.945 164.795 ;
        RECT 79.160 164.205 79.490 164.965 ;
        RECT 78.775 163.865 79.490 164.035 ;
        RECT 79.660 163.890 79.915 164.795 ;
        RECT 77.710 163.655 77.880 163.865 ;
        RECT 77.625 163.325 77.880 163.655 ;
        RECT 77.285 162.585 77.540 163.160 ;
        RECT 77.710 163.135 77.880 163.325 ;
        RECT 78.160 163.315 78.515 163.685 ;
        RECT 78.685 163.315 79.040 163.685 ;
        RECT 79.320 163.655 79.490 163.865 ;
        RECT 79.320 163.325 79.575 163.655 ;
        RECT 79.320 163.135 79.490 163.325 ;
        RECT 79.745 163.160 79.915 163.890 ;
        RECT 80.090 163.815 80.350 164.965 ;
        RECT 80.525 163.875 81.735 164.965 ;
        RECT 80.525 163.335 81.045 163.875 ;
        RECT 81.905 163.825 82.245 164.795 ;
        RECT 82.415 163.825 82.585 164.965 ;
        RECT 82.855 164.165 83.105 164.965 ;
        RECT 83.750 163.995 84.080 164.795 ;
        RECT 84.380 164.165 84.710 164.965 ;
        RECT 84.880 163.995 85.210 164.795 ;
        RECT 82.775 163.825 85.210 163.995 ;
        RECT 85.960 163.985 86.215 164.655 ;
        RECT 86.395 164.165 86.680 164.965 ;
        RECT 86.860 164.245 87.190 164.755 ;
        RECT 85.960 163.945 86.140 163.985 ;
        RECT 77.710 162.965 78.425 163.135 ;
        RECT 77.710 162.415 78.040 162.795 ;
        RECT 78.255 162.585 78.425 162.965 ;
        RECT 78.775 162.965 79.490 163.135 ;
        RECT 78.775 162.585 78.945 162.965 ;
        RECT 79.160 162.415 79.490 162.795 ;
        RECT 79.660 162.585 79.915 163.160 ;
        RECT 80.090 162.415 80.350 163.255 ;
        RECT 81.215 163.165 81.735 163.705 ;
        RECT 80.525 162.415 81.735 163.165 ;
        RECT 81.905 163.215 82.080 163.825 ;
        RECT 82.775 163.575 82.945 163.825 ;
        RECT 82.250 163.405 82.945 163.575 ;
        RECT 83.120 163.405 83.540 163.605 ;
        RECT 83.710 163.405 84.040 163.605 ;
        RECT 84.210 163.405 84.540 163.605 ;
        RECT 81.905 162.585 82.245 163.215 ;
        RECT 82.415 162.415 82.665 163.215 ;
        RECT 82.855 163.065 84.080 163.235 ;
        RECT 82.855 162.585 83.185 163.065 ;
        RECT 83.355 162.415 83.580 162.875 ;
        RECT 83.750 162.585 84.080 163.065 ;
        RECT 84.710 163.195 84.880 163.825 ;
        RECT 85.875 163.775 86.140 163.945 ;
        RECT 85.065 163.405 85.415 163.655 ;
        RECT 84.710 162.585 85.210 163.195 ;
        RECT 85.960 163.125 86.140 163.775 ;
        RECT 86.860 163.655 87.110 164.245 ;
        RECT 87.460 164.095 87.630 164.705 ;
        RECT 87.800 164.275 88.130 164.965 ;
        RECT 88.360 164.415 88.600 164.705 ;
        RECT 88.800 164.585 89.220 164.965 ;
        RECT 89.400 164.495 90.030 164.745 ;
        RECT 90.500 164.585 90.830 164.965 ;
        RECT 89.400 164.415 89.570 164.495 ;
        RECT 91.000 164.415 91.170 164.705 ;
        RECT 91.350 164.585 91.730 164.965 ;
        RECT 91.970 164.580 92.800 164.750 ;
        RECT 88.360 164.245 89.570 164.415 ;
        RECT 86.310 163.325 87.110 163.655 ;
        RECT 85.960 162.595 86.215 163.125 ;
        RECT 86.395 162.415 86.680 162.875 ;
        RECT 86.860 162.675 87.110 163.325 ;
        RECT 87.310 164.075 87.630 164.095 ;
        RECT 87.310 163.905 89.230 164.075 ;
        RECT 87.310 163.010 87.500 163.905 ;
        RECT 89.400 163.735 89.570 164.245 ;
        RECT 89.740 163.985 90.260 164.295 ;
        RECT 87.670 163.565 89.570 163.735 ;
        RECT 87.670 163.505 88.000 163.565 ;
        RECT 88.150 163.335 88.480 163.395 ;
        RECT 87.820 163.065 88.480 163.335 ;
        RECT 87.310 162.680 87.630 163.010 ;
        RECT 87.810 162.415 88.470 162.895 ;
        RECT 88.670 162.805 88.840 163.565 ;
        RECT 89.740 163.395 89.920 163.805 ;
        RECT 89.010 163.225 89.340 163.345 ;
        RECT 90.090 163.225 90.260 163.985 ;
        RECT 89.010 163.055 90.260 163.225 ;
        RECT 90.430 164.165 91.800 164.415 ;
        RECT 90.430 163.395 90.620 164.165 ;
        RECT 91.550 163.905 91.800 164.165 ;
        RECT 90.790 163.735 91.040 163.895 ;
        RECT 91.970 163.735 92.140 164.580 ;
        RECT 93.035 164.295 93.205 164.795 ;
        RECT 93.375 164.465 93.705 164.965 ;
        RECT 92.310 163.905 92.810 164.285 ;
        RECT 93.035 164.125 93.730 164.295 ;
        RECT 90.790 163.565 92.140 163.735 ;
        RECT 91.720 163.525 92.140 163.565 ;
        RECT 90.430 163.055 90.850 163.395 ;
        RECT 91.140 163.065 91.550 163.395 ;
        RECT 88.670 162.635 89.520 162.805 ;
        RECT 90.080 162.415 90.400 162.875 ;
        RECT 90.600 162.625 90.850 163.055 ;
        RECT 91.140 162.415 91.550 162.855 ;
        RECT 91.720 162.795 91.890 163.525 ;
        RECT 92.060 162.975 92.410 163.345 ;
        RECT 92.590 163.035 92.810 163.905 ;
        RECT 92.980 163.335 93.390 163.955 ;
        RECT 93.560 163.155 93.730 164.125 ;
        RECT 93.035 162.965 93.730 163.155 ;
        RECT 91.720 162.595 92.735 162.795 ;
        RECT 93.035 162.635 93.205 162.965 ;
        RECT 93.375 162.415 93.705 162.795 ;
        RECT 93.920 162.675 94.145 164.795 ;
        RECT 94.315 164.465 94.645 164.965 ;
        RECT 94.815 164.295 94.985 164.795 ;
        RECT 94.320 164.125 94.985 164.295 ;
        RECT 94.320 163.135 94.550 164.125 ;
        RECT 94.720 163.305 95.070 163.955 ;
        RECT 95.245 163.875 96.455 164.965 ;
        RECT 95.245 163.335 95.765 163.875 ;
        RECT 96.665 163.825 96.895 164.965 ;
        RECT 97.065 163.815 97.395 164.795 ;
        RECT 97.565 163.825 97.775 164.965 ;
        RECT 98.210 163.995 98.540 164.795 ;
        RECT 98.710 164.165 99.040 164.965 ;
        RECT 99.340 163.995 99.670 164.795 ;
        RECT 100.315 164.165 100.565 164.965 ;
        RECT 98.210 163.825 100.645 163.995 ;
        RECT 100.835 163.825 101.005 164.965 ;
        RECT 101.175 163.825 101.515 164.795 ;
        RECT 95.935 163.165 96.455 163.705 ;
        RECT 96.645 163.405 96.975 163.655 ;
        RECT 94.320 162.965 94.985 163.135 ;
        RECT 94.315 162.415 94.645 162.795 ;
        RECT 94.815 162.675 94.985 162.965 ;
        RECT 95.245 162.415 96.455 163.165 ;
        RECT 96.665 162.415 96.895 163.235 ;
        RECT 97.145 163.215 97.395 163.815 ;
        RECT 98.005 163.405 98.355 163.655 ;
        RECT 97.065 162.585 97.395 163.215 ;
        RECT 97.565 162.415 97.775 163.235 ;
        RECT 98.540 163.195 98.710 163.825 ;
        RECT 98.880 163.405 99.210 163.605 ;
        RECT 99.380 163.405 99.710 163.605 ;
        RECT 99.880 163.405 100.300 163.605 ;
        RECT 100.475 163.575 100.645 163.825 ;
        RECT 100.475 163.405 101.170 163.575 ;
        RECT 98.210 162.585 98.710 163.195 ;
        RECT 99.340 163.065 100.565 163.235 ;
        RECT 101.340 163.215 101.515 163.825 ;
        RECT 101.685 163.800 101.975 164.965 ;
        RECT 102.145 163.875 103.815 164.965 ;
        RECT 104.190 163.995 104.520 164.795 ;
        RECT 104.690 164.165 105.020 164.965 ;
        RECT 105.320 163.995 105.650 164.795 ;
        RECT 106.295 164.165 106.545 164.965 ;
        RECT 102.145 163.355 102.895 163.875 ;
        RECT 104.190 163.825 106.625 163.995 ;
        RECT 106.815 163.825 106.985 164.965 ;
        RECT 107.155 163.825 107.495 164.795 ;
        RECT 99.340 162.585 99.670 163.065 ;
        RECT 99.840 162.415 100.065 162.875 ;
        RECT 100.235 162.585 100.565 163.065 ;
        RECT 100.755 162.415 101.005 163.215 ;
        RECT 101.175 162.585 101.515 163.215 ;
        RECT 103.065 163.185 103.815 163.705 ;
        RECT 103.985 163.405 104.335 163.655 ;
        RECT 104.520 163.195 104.690 163.825 ;
        RECT 104.860 163.405 105.190 163.605 ;
        RECT 105.360 163.405 105.690 163.605 ;
        RECT 105.860 163.435 106.285 163.605 ;
        RECT 106.455 163.575 106.625 163.825 ;
        RECT 105.860 163.405 106.280 163.435 ;
        RECT 106.455 163.405 107.150 163.575 ;
        RECT 107.320 163.265 107.495 163.825 ;
        RECT 101.685 162.415 101.975 163.140 ;
        RECT 102.145 162.415 103.815 163.185 ;
        RECT 104.190 162.585 104.690 163.195 ;
        RECT 105.320 163.065 106.545 163.235 ;
        RECT 107.265 163.215 107.495 163.265 ;
        RECT 105.320 162.585 105.650 163.065 ;
        RECT 105.820 162.415 106.045 162.875 ;
        RECT 106.215 162.585 106.545 163.065 ;
        RECT 106.735 162.415 106.985 163.215 ;
        RECT 107.155 162.585 107.495 163.215 ;
        RECT 107.665 163.825 108.005 164.795 ;
        RECT 108.175 163.825 108.345 164.965 ;
        RECT 108.615 164.165 108.865 164.965 ;
        RECT 109.510 163.995 109.840 164.795 ;
        RECT 110.140 164.165 110.470 164.965 ;
        RECT 110.640 163.995 110.970 164.795 ;
        RECT 108.535 163.825 110.970 163.995 ;
        RECT 111.345 163.825 111.685 164.795 ;
        RECT 111.855 163.825 112.025 164.965 ;
        RECT 112.295 164.165 112.545 164.965 ;
        RECT 113.190 163.995 113.520 164.795 ;
        RECT 113.820 164.165 114.150 164.965 ;
        RECT 114.320 163.995 114.650 164.795 ;
        RECT 112.215 163.825 114.650 163.995 ;
        RECT 115.230 163.995 115.560 164.795 ;
        RECT 115.730 164.165 116.060 164.965 ;
        RECT 116.360 163.995 116.690 164.795 ;
        RECT 117.335 164.165 117.585 164.965 ;
        RECT 115.230 163.825 117.665 163.995 ;
        RECT 117.855 163.825 118.025 164.965 ;
        RECT 118.195 163.825 118.535 164.795 ;
        RECT 107.665 163.215 107.840 163.825 ;
        RECT 108.535 163.575 108.705 163.825 ;
        RECT 108.010 163.405 108.705 163.575 ;
        RECT 108.880 163.405 109.300 163.605 ;
        RECT 109.470 163.405 109.800 163.605 ;
        RECT 109.970 163.405 110.300 163.605 ;
        RECT 107.665 162.585 108.005 163.215 ;
        RECT 108.175 162.415 108.425 163.215 ;
        RECT 108.615 163.065 109.840 163.235 ;
        RECT 108.615 162.585 108.945 163.065 ;
        RECT 109.115 162.415 109.340 162.875 ;
        RECT 109.510 162.585 109.840 163.065 ;
        RECT 110.470 163.195 110.640 163.825 ;
        RECT 110.825 163.405 111.175 163.655 ;
        RECT 111.345 163.215 111.520 163.825 ;
        RECT 112.215 163.575 112.385 163.825 ;
        RECT 111.690 163.405 112.385 163.575 ;
        RECT 112.560 163.405 112.980 163.605 ;
        RECT 113.150 163.405 113.480 163.605 ;
        RECT 113.650 163.405 113.980 163.605 ;
        RECT 110.470 162.585 110.970 163.195 ;
        RECT 111.345 162.585 111.685 163.215 ;
        RECT 111.855 162.415 112.105 163.215 ;
        RECT 112.295 163.065 113.520 163.235 ;
        RECT 112.295 162.585 112.625 163.065 ;
        RECT 112.795 162.415 113.020 162.875 ;
        RECT 113.190 162.585 113.520 163.065 ;
        RECT 114.150 163.195 114.320 163.825 ;
        RECT 114.505 163.405 114.855 163.655 ;
        RECT 115.025 163.405 115.375 163.655 ;
        RECT 115.560 163.195 115.730 163.825 ;
        RECT 115.900 163.405 116.230 163.605 ;
        RECT 116.400 163.405 116.730 163.605 ;
        RECT 116.900 163.405 117.320 163.605 ;
        RECT 117.495 163.575 117.665 163.825 ;
        RECT 117.495 163.405 118.190 163.575 ;
        RECT 114.150 162.585 114.650 163.195 ;
        RECT 115.230 162.585 115.730 163.195 ;
        RECT 116.360 163.065 117.585 163.235 ;
        RECT 118.360 163.215 118.535 163.825 ;
        RECT 119.165 163.875 120.835 164.965 ;
        RECT 121.010 164.530 126.355 164.965 ;
        RECT 119.165 163.355 119.915 163.875 ;
        RECT 116.360 162.585 116.690 163.065 ;
        RECT 116.860 162.415 117.085 162.875 ;
        RECT 117.255 162.585 117.585 163.065 ;
        RECT 117.775 162.415 118.025 163.215 ;
        RECT 118.195 162.585 118.535 163.215 ;
        RECT 120.085 163.185 120.835 163.705 ;
        RECT 122.600 163.280 122.950 164.530 ;
        RECT 126.525 163.875 127.735 164.965 ;
        RECT 119.165 162.415 120.835 163.185 ;
        RECT 124.430 162.960 124.770 163.790 ;
        RECT 126.525 163.335 127.045 163.875 ;
        RECT 127.215 163.165 127.735 163.705 ;
        RECT 121.010 162.415 126.355 162.960 ;
        RECT 126.525 162.415 127.735 163.165 ;
        RECT 29.840 162.245 127.820 162.415 ;
        RECT 29.925 161.495 31.135 162.245 ;
        RECT 29.925 160.955 30.445 161.495 ;
        RECT 32.225 161.475 35.735 162.245 ;
        RECT 30.615 160.785 31.135 161.325 ;
        RECT 29.925 159.695 31.135 160.785 ;
        RECT 32.225 160.785 33.915 161.305 ;
        RECT 34.085 160.955 35.735 161.475 ;
        RECT 35.965 161.425 36.175 162.245 ;
        RECT 36.345 161.445 36.675 162.075 ;
        RECT 36.345 160.845 36.595 161.445 ;
        RECT 36.845 161.425 37.075 162.245 ;
        RECT 37.285 161.520 37.575 162.245 ;
        RECT 37.745 161.475 40.335 162.245 ;
        RECT 36.765 161.005 37.095 161.255 ;
        RECT 32.225 159.695 35.735 160.785 ;
        RECT 35.965 159.695 36.175 160.835 ;
        RECT 36.345 159.865 36.675 160.845 ;
        RECT 36.845 159.695 37.075 160.835 ;
        RECT 37.285 159.695 37.575 160.860 ;
        RECT 37.745 160.785 38.955 161.305 ;
        RECT 39.125 160.955 40.335 161.475 ;
        RECT 40.505 161.570 40.765 162.075 ;
        RECT 40.945 161.865 41.275 162.245 ;
        RECT 41.455 161.695 41.625 162.075 ;
        RECT 37.745 159.695 40.335 160.785 ;
        RECT 40.505 160.770 40.675 161.570 ;
        RECT 40.960 161.525 41.625 161.695 ;
        RECT 40.960 161.270 41.130 161.525 ;
        RECT 41.925 161.425 42.155 162.245 ;
        RECT 42.325 161.445 42.655 162.075 ;
        RECT 40.845 160.940 41.130 161.270 ;
        RECT 41.365 160.975 41.695 161.345 ;
        RECT 41.905 161.005 42.235 161.255 ;
        RECT 40.960 160.795 41.130 160.940 ;
        RECT 42.405 160.845 42.655 161.445 ;
        RECT 42.825 161.425 43.035 162.245 ;
        RECT 43.470 161.465 43.970 162.075 ;
        RECT 43.265 161.005 43.615 161.255 ;
        RECT 40.505 159.865 40.775 160.770 ;
        RECT 40.960 160.625 41.625 160.795 ;
        RECT 40.945 159.695 41.275 160.455 ;
        RECT 41.455 159.865 41.625 160.625 ;
        RECT 41.925 159.695 42.155 160.835 ;
        RECT 42.325 159.865 42.655 160.845 ;
        RECT 43.800 160.835 43.970 161.465 ;
        RECT 44.600 161.595 44.930 162.075 ;
        RECT 45.100 161.785 45.325 162.245 ;
        RECT 45.495 161.595 45.825 162.075 ;
        RECT 44.600 161.425 45.825 161.595 ;
        RECT 46.015 161.445 46.265 162.245 ;
        RECT 46.435 161.445 46.775 162.075 ;
        RECT 47.150 161.465 47.650 162.075 ;
        RECT 44.140 161.055 44.470 161.255 ;
        RECT 44.640 161.055 44.970 161.255 ;
        RECT 45.140 161.055 45.560 161.255 ;
        RECT 45.735 161.085 46.430 161.255 ;
        RECT 45.735 160.835 45.905 161.085 ;
        RECT 46.600 160.835 46.775 161.445 ;
        RECT 46.945 161.005 47.295 161.255 ;
        RECT 47.480 160.835 47.650 161.465 ;
        RECT 48.280 161.595 48.610 162.075 ;
        RECT 48.780 161.785 49.005 162.245 ;
        RECT 49.175 161.595 49.505 162.075 ;
        RECT 48.280 161.425 49.505 161.595 ;
        RECT 49.695 161.445 49.945 162.245 ;
        RECT 50.115 161.445 50.455 162.075 ;
        RECT 47.820 161.055 48.150 161.255 ;
        RECT 48.320 161.055 48.650 161.255 ;
        RECT 48.820 161.055 49.240 161.255 ;
        RECT 49.415 161.085 50.110 161.255 ;
        RECT 49.415 160.835 49.585 161.085 ;
        RECT 50.280 160.835 50.455 161.445 ;
        RECT 42.825 159.695 43.035 160.835 ;
        RECT 43.470 160.665 45.905 160.835 ;
        RECT 43.470 159.865 43.800 160.665 ;
        RECT 43.970 159.695 44.300 160.495 ;
        RECT 44.600 159.865 44.930 160.665 ;
        RECT 45.575 159.695 45.825 160.495 ;
        RECT 46.095 159.695 46.265 160.835 ;
        RECT 46.435 159.865 46.775 160.835 ;
        RECT 47.150 160.665 49.585 160.835 ;
        RECT 47.150 159.865 47.480 160.665 ;
        RECT 47.650 159.695 47.980 160.495 ;
        RECT 48.280 159.865 48.610 160.665 ;
        RECT 49.255 159.695 49.505 160.495 ;
        RECT 49.775 159.695 49.945 160.835 ;
        RECT 50.115 159.865 50.455 160.835 ;
        RECT 50.625 161.570 50.885 162.075 ;
        RECT 51.065 161.865 51.395 162.245 ;
        RECT 51.575 161.695 51.745 162.075 ;
        RECT 50.625 160.770 50.795 161.570 ;
        RECT 51.080 161.525 51.745 161.695 ;
        RECT 51.080 161.270 51.250 161.525 ;
        RECT 52.465 161.475 54.135 162.245 ;
        RECT 54.395 161.695 54.565 162.075 ;
        RECT 54.745 161.865 55.075 162.245 ;
        RECT 54.395 161.525 55.060 161.695 ;
        RECT 55.255 161.570 55.515 162.075 ;
        RECT 50.965 160.940 51.250 161.270 ;
        RECT 51.485 160.975 51.815 161.345 ;
        RECT 51.080 160.795 51.250 160.940 ;
        RECT 50.625 159.865 50.895 160.770 ;
        RECT 51.080 160.625 51.745 160.795 ;
        RECT 51.065 159.695 51.395 160.455 ;
        RECT 51.575 159.865 51.745 160.625 ;
        RECT 52.465 160.785 53.215 161.305 ;
        RECT 53.385 160.955 54.135 161.475 ;
        RECT 54.325 160.975 54.655 161.345 ;
        RECT 54.890 161.270 55.060 161.525 ;
        RECT 54.890 160.940 55.175 161.270 ;
        RECT 54.890 160.795 55.060 160.940 ;
        RECT 52.465 159.695 54.135 160.785 ;
        RECT 54.395 160.625 55.060 160.795 ;
        RECT 55.345 160.770 55.515 161.570 ;
        RECT 54.395 159.865 54.565 160.625 ;
        RECT 54.745 159.695 55.075 160.455 ;
        RECT 55.245 159.865 55.515 160.770 ;
        RECT 55.685 161.445 56.025 162.075 ;
        RECT 56.195 161.445 56.445 162.245 ;
        RECT 56.635 161.595 56.965 162.075 ;
        RECT 57.135 161.785 57.360 162.245 ;
        RECT 57.530 161.595 57.860 162.075 ;
        RECT 55.685 160.835 55.860 161.445 ;
        RECT 56.635 161.425 57.860 161.595 ;
        RECT 58.490 161.465 58.990 162.075 ;
        RECT 56.030 161.085 56.725 161.255 ;
        RECT 56.555 160.835 56.725 161.085 ;
        RECT 56.900 161.055 57.320 161.255 ;
        RECT 57.490 161.055 57.820 161.255 ;
        RECT 57.990 161.055 58.320 161.255 ;
        RECT 58.490 160.835 58.660 161.465 ;
        RECT 59.365 161.445 59.705 162.075 ;
        RECT 59.875 161.445 60.125 162.245 ;
        RECT 60.315 161.595 60.645 162.075 ;
        RECT 60.815 161.785 61.040 162.245 ;
        RECT 61.210 161.595 61.540 162.075 ;
        RECT 58.845 161.005 59.195 161.255 ;
        RECT 59.365 160.835 59.540 161.445 ;
        RECT 60.315 161.425 61.540 161.595 ;
        RECT 62.170 161.465 62.670 162.075 ;
        RECT 63.045 161.520 63.335 162.245 ;
        RECT 63.965 161.475 66.555 162.245 ;
        RECT 59.710 161.085 60.405 161.255 ;
        RECT 60.235 160.835 60.405 161.085 ;
        RECT 60.580 161.055 61.000 161.255 ;
        RECT 61.170 161.055 61.500 161.255 ;
        RECT 61.670 161.055 62.000 161.255 ;
        RECT 62.170 160.835 62.340 161.465 ;
        RECT 62.525 161.005 62.875 161.255 ;
        RECT 55.685 159.865 56.025 160.835 ;
        RECT 56.195 159.695 56.365 160.835 ;
        RECT 56.555 160.665 58.990 160.835 ;
        RECT 56.635 159.695 56.885 160.495 ;
        RECT 57.530 159.865 57.860 160.665 ;
        RECT 58.160 159.695 58.490 160.495 ;
        RECT 58.660 159.865 58.990 160.665 ;
        RECT 59.365 159.865 59.705 160.835 ;
        RECT 59.875 159.695 60.045 160.835 ;
        RECT 60.235 160.665 62.670 160.835 ;
        RECT 60.315 159.695 60.565 160.495 ;
        RECT 61.210 159.865 61.540 160.665 ;
        RECT 61.840 159.695 62.170 160.495 ;
        RECT 62.340 159.865 62.670 160.665 ;
        RECT 63.045 159.695 63.335 160.860 ;
        RECT 63.965 160.785 65.175 161.305 ;
        RECT 65.345 160.955 66.555 161.475 ;
        RECT 66.785 161.425 66.995 162.245 ;
        RECT 67.165 161.445 67.495 162.075 ;
        RECT 67.165 160.845 67.415 161.445 ;
        RECT 67.665 161.425 67.895 162.245 ;
        RECT 68.195 161.695 68.365 162.075 ;
        RECT 68.545 161.865 68.875 162.245 ;
        RECT 68.195 161.525 68.860 161.695 ;
        RECT 69.055 161.570 69.315 162.075 ;
        RECT 67.585 161.005 67.915 161.255 ;
        RECT 68.125 160.975 68.455 161.345 ;
        RECT 68.690 161.270 68.860 161.525 ;
        RECT 68.690 160.940 68.975 161.270 ;
        RECT 63.965 159.695 66.555 160.785 ;
        RECT 66.785 159.695 66.995 160.835 ;
        RECT 67.165 159.865 67.495 160.845 ;
        RECT 67.665 159.695 67.895 160.835 ;
        RECT 68.690 160.795 68.860 160.940 ;
        RECT 68.195 160.625 68.860 160.795 ;
        RECT 69.145 160.770 69.315 161.570 ;
        RECT 69.485 161.475 71.155 162.245 ;
        RECT 68.195 159.865 68.365 160.625 ;
        RECT 68.545 159.695 68.875 160.455 ;
        RECT 69.045 159.865 69.315 160.770 ;
        RECT 69.485 160.785 70.235 161.305 ;
        RECT 70.405 160.955 71.155 161.475 ;
        RECT 71.330 161.405 71.590 162.245 ;
        RECT 71.765 161.500 72.020 162.075 ;
        RECT 72.190 161.865 72.520 162.245 ;
        RECT 72.735 161.695 72.905 162.075 ;
        RECT 73.255 161.765 73.555 162.245 ;
        RECT 72.190 161.525 72.905 161.695 ;
        RECT 73.725 161.595 73.985 162.050 ;
        RECT 74.155 161.765 74.415 162.245 ;
        RECT 74.595 161.595 74.855 162.050 ;
        RECT 75.025 161.765 75.275 162.245 ;
        RECT 75.455 161.595 75.715 162.050 ;
        RECT 75.885 161.765 76.135 162.245 ;
        RECT 76.315 161.595 76.575 162.050 ;
        RECT 76.745 161.765 76.990 162.245 ;
        RECT 77.160 161.595 77.435 162.050 ;
        RECT 77.605 161.765 77.850 162.245 ;
        RECT 78.020 161.595 78.280 162.050 ;
        RECT 78.450 161.765 78.710 162.245 ;
        RECT 78.880 161.595 79.140 162.050 ;
        RECT 79.310 161.765 79.570 162.245 ;
        RECT 79.740 161.595 80.000 162.050 ;
        RECT 80.170 161.685 80.430 162.245 ;
        RECT 73.255 161.565 80.000 161.595 ;
        RECT 69.485 159.695 71.155 160.785 ;
        RECT 71.330 159.695 71.590 160.845 ;
        RECT 71.765 160.770 71.935 161.500 ;
        RECT 72.190 161.335 72.360 161.525 ;
        RECT 73.225 161.425 80.000 161.565 ;
        RECT 73.225 161.395 74.420 161.425 ;
        RECT 72.105 161.005 72.360 161.335 ;
        RECT 72.190 160.795 72.360 161.005 ;
        RECT 72.640 160.975 72.995 161.345 ;
        RECT 73.255 160.835 74.420 161.395 ;
        RECT 80.600 161.255 80.850 162.065 ;
        RECT 81.030 161.720 81.290 162.245 ;
        RECT 81.460 161.255 81.710 162.065 ;
        RECT 81.890 161.735 82.195 162.245 ;
        RECT 74.590 161.005 81.710 161.255 ;
        RECT 81.880 161.005 82.195 161.565 ;
        RECT 82.825 161.445 83.165 162.075 ;
        RECT 83.335 161.445 83.585 162.245 ;
        RECT 83.775 161.595 84.105 162.075 ;
        RECT 84.275 161.785 84.500 162.245 ;
        RECT 84.670 161.595 85.000 162.075 ;
        RECT 71.765 159.865 72.020 160.770 ;
        RECT 72.190 160.625 72.905 160.795 ;
        RECT 72.190 159.695 72.520 160.455 ;
        RECT 72.735 159.865 72.905 160.625 ;
        RECT 73.255 160.610 80.000 160.835 ;
        RECT 73.255 159.695 73.525 160.440 ;
        RECT 73.695 159.870 73.985 160.610 ;
        RECT 74.595 160.595 80.000 160.610 ;
        RECT 74.155 159.700 74.410 160.425 ;
        RECT 74.595 159.870 74.855 160.595 ;
        RECT 75.025 159.700 75.270 160.425 ;
        RECT 75.455 159.870 75.715 160.595 ;
        RECT 75.885 159.700 76.130 160.425 ;
        RECT 76.315 159.870 76.575 160.595 ;
        RECT 76.745 159.700 76.990 160.425 ;
        RECT 77.160 159.870 77.420 160.595 ;
        RECT 77.590 159.700 77.850 160.425 ;
        RECT 78.020 159.870 78.280 160.595 ;
        RECT 78.450 159.700 78.710 160.425 ;
        RECT 78.880 159.870 79.140 160.595 ;
        RECT 79.310 159.700 79.570 160.425 ;
        RECT 79.740 159.870 80.000 160.595 ;
        RECT 80.170 159.700 80.430 160.495 ;
        RECT 80.600 159.870 80.850 161.005 ;
        RECT 74.155 159.695 80.430 159.700 ;
        RECT 81.030 159.695 81.290 160.505 ;
        RECT 81.465 159.865 81.710 161.005 ;
        RECT 82.825 160.835 83.000 161.445 ;
        RECT 83.775 161.425 85.000 161.595 ;
        RECT 85.630 161.465 86.130 162.075 ;
        RECT 86.965 161.475 88.635 162.245 ;
        RECT 88.805 161.520 89.095 162.245 ;
        RECT 89.265 161.475 91.855 162.245 ;
        RECT 83.170 161.085 83.865 161.255 ;
        RECT 83.695 160.835 83.865 161.085 ;
        RECT 84.040 161.055 84.460 161.255 ;
        RECT 84.630 161.055 84.960 161.255 ;
        RECT 85.130 161.055 85.460 161.255 ;
        RECT 85.630 160.835 85.800 161.465 ;
        RECT 85.985 161.005 86.335 161.255 ;
        RECT 81.890 159.695 82.185 160.505 ;
        RECT 82.825 159.865 83.165 160.835 ;
        RECT 83.335 159.695 83.505 160.835 ;
        RECT 83.695 160.665 86.130 160.835 ;
        RECT 83.775 159.695 84.025 160.495 ;
        RECT 84.670 159.865 85.000 160.665 ;
        RECT 85.300 159.695 85.630 160.495 ;
        RECT 85.800 159.865 86.130 160.665 ;
        RECT 86.965 160.785 87.715 161.305 ;
        RECT 87.885 160.955 88.635 161.475 ;
        RECT 86.965 159.695 88.635 160.785 ;
        RECT 88.805 159.695 89.095 160.860 ;
        RECT 89.265 160.785 90.475 161.305 ;
        RECT 90.645 160.955 91.855 161.475 ;
        RECT 92.085 161.425 92.295 162.245 ;
        RECT 92.465 161.445 92.795 162.075 ;
        RECT 92.465 160.845 92.715 161.445 ;
        RECT 92.965 161.425 93.195 162.245 ;
        RECT 93.865 161.475 96.455 162.245 ;
        RECT 92.885 161.005 93.215 161.255 ;
        RECT 89.265 159.695 91.855 160.785 ;
        RECT 92.085 159.695 92.295 160.835 ;
        RECT 92.465 159.865 92.795 160.845 ;
        RECT 92.965 159.695 93.195 160.835 ;
        RECT 93.865 160.785 95.075 161.305 ;
        RECT 95.245 160.955 96.455 161.475 ;
        RECT 96.630 161.535 96.885 162.065 ;
        RECT 97.055 161.785 97.360 162.245 ;
        RECT 97.605 161.865 98.675 162.035 ;
        RECT 96.630 160.885 96.840 161.535 ;
        RECT 97.605 161.510 97.925 161.865 ;
        RECT 97.600 161.335 97.925 161.510 ;
        RECT 97.010 161.035 97.925 161.335 ;
        RECT 98.095 161.295 98.335 161.695 ;
        RECT 98.505 161.635 98.675 161.865 ;
        RECT 98.845 161.805 99.035 162.245 ;
        RECT 99.205 161.795 100.155 162.075 ;
        RECT 100.375 161.885 100.725 162.055 ;
        RECT 98.505 161.465 99.035 161.635 ;
        RECT 97.010 161.005 97.750 161.035 ;
        RECT 93.865 159.695 96.455 160.785 ;
        RECT 96.630 160.005 96.885 160.885 ;
        RECT 97.055 159.695 97.360 160.835 ;
        RECT 97.580 160.415 97.750 161.005 ;
        RECT 98.095 160.925 98.635 161.295 ;
        RECT 98.815 161.185 99.035 161.465 ;
        RECT 99.205 161.015 99.375 161.795 ;
        RECT 98.970 160.845 99.375 161.015 ;
        RECT 99.545 161.005 99.895 161.625 ;
        RECT 98.970 160.755 99.140 160.845 ;
        RECT 100.065 160.835 100.275 161.625 ;
        RECT 97.920 160.585 99.140 160.755 ;
        RECT 99.600 160.675 100.275 160.835 ;
        RECT 97.580 160.245 98.380 160.415 ;
        RECT 97.700 159.695 98.030 160.075 ;
        RECT 98.210 159.955 98.380 160.245 ;
        RECT 98.970 160.205 99.140 160.585 ;
        RECT 99.310 160.665 100.275 160.675 ;
        RECT 100.465 161.495 100.725 161.885 ;
        RECT 100.935 161.785 101.265 162.245 ;
        RECT 102.140 161.855 102.995 162.025 ;
        RECT 103.200 161.855 103.695 162.025 ;
        RECT 103.865 161.885 104.195 162.245 ;
        RECT 100.465 160.805 100.635 161.495 ;
        RECT 100.805 161.145 100.975 161.325 ;
        RECT 101.145 161.315 101.935 161.565 ;
        RECT 102.140 161.145 102.310 161.855 ;
        RECT 102.480 161.345 102.835 161.565 ;
        RECT 100.805 160.975 102.495 161.145 ;
        RECT 99.310 160.375 99.770 160.665 ;
        RECT 100.465 160.635 101.965 160.805 ;
        RECT 100.465 160.495 100.635 160.635 ;
        RECT 100.075 160.325 100.635 160.495 ;
        RECT 98.550 159.695 98.800 160.155 ;
        RECT 98.970 159.865 99.840 160.205 ;
        RECT 100.075 159.865 100.245 160.325 ;
        RECT 101.080 160.295 102.155 160.465 ;
        RECT 100.415 159.695 100.785 160.155 ;
        RECT 101.080 159.955 101.250 160.295 ;
        RECT 101.420 159.695 101.750 160.125 ;
        RECT 101.985 159.955 102.155 160.295 ;
        RECT 102.325 160.195 102.495 160.975 ;
        RECT 102.665 160.755 102.835 161.345 ;
        RECT 103.005 160.945 103.355 161.565 ;
        RECT 102.665 160.365 103.130 160.755 ;
        RECT 103.525 160.495 103.695 161.855 ;
        RECT 103.865 160.665 104.325 161.715 ;
        RECT 103.300 160.325 103.695 160.495 ;
        RECT 103.300 160.195 103.470 160.325 ;
        RECT 102.325 159.865 103.005 160.195 ;
        RECT 103.220 159.865 103.470 160.195 ;
        RECT 103.640 159.695 103.890 160.155 ;
        RECT 104.060 159.880 104.385 160.665 ;
        RECT 104.555 159.865 104.725 161.985 ;
        RECT 104.895 161.865 105.225 162.245 ;
        RECT 105.395 161.695 105.650 161.985 ;
        RECT 104.900 161.525 105.650 161.695 ;
        RECT 104.900 160.535 105.130 161.525 ;
        RECT 105.825 161.495 107.035 162.245 ;
        RECT 105.300 160.705 105.650 161.355 ;
        RECT 105.825 160.785 106.345 161.325 ;
        RECT 106.515 160.955 107.035 161.495 ;
        RECT 107.205 161.445 107.545 162.075 ;
        RECT 107.715 161.445 107.965 162.245 ;
        RECT 108.155 161.595 108.485 162.075 ;
        RECT 108.655 161.785 108.880 162.245 ;
        RECT 109.050 161.595 109.380 162.075 ;
        RECT 107.205 160.835 107.380 161.445 ;
        RECT 108.155 161.425 109.380 161.595 ;
        RECT 110.010 161.465 110.510 162.075 ;
        RECT 111.000 161.615 111.285 162.075 ;
        RECT 111.455 161.785 111.725 162.245 ;
        RECT 107.550 161.085 108.245 161.255 ;
        RECT 108.075 160.835 108.245 161.085 ;
        RECT 108.420 161.055 108.840 161.255 ;
        RECT 109.010 161.055 109.340 161.255 ;
        RECT 109.510 161.055 109.840 161.255 ;
        RECT 110.010 160.835 110.180 161.465 ;
        RECT 111.000 161.445 111.955 161.615 ;
        RECT 110.365 161.005 110.715 161.255 ;
        RECT 104.900 160.365 105.650 160.535 ;
        RECT 104.895 159.695 105.225 160.195 ;
        RECT 105.395 159.865 105.650 160.365 ;
        RECT 105.825 159.695 107.035 160.785 ;
        RECT 107.205 159.865 107.545 160.835 ;
        RECT 107.715 159.695 107.885 160.835 ;
        RECT 108.075 160.665 110.510 160.835 ;
        RECT 110.885 160.715 111.575 161.275 ;
        RECT 108.155 159.695 108.405 160.495 ;
        RECT 109.050 159.865 109.380 160.665 ;
        RECT 109.680 159.695 110.010 160.495 ;
        RECT 110.180 159.865 110.510 160.665 ;
        RECT 111.745 160.545 111.955 161.445 ;
        RECT 111.000 160.325 111.955 160.545 ;
        RECT 112.125 161.275 112.525 162.075 ;
        RECT 112.715 161.615 112.995 162.075 ;
        RECT 113.515 161.785 113.840 162.245 ;
        RECT 112.715 161.445 113.840 161.615 ;
        RECT 114.010 161.505 114.395 162.075 ;
        RECT 114.565 161.520 114.855 162.245 ;
        RECT 113.390 161.335 113.840 161.445 ;
        RECT 112.125 160.715 113.220 161.275 ;
        RECT 113.390 161.005 113.945 161.335 ;
        RECT 111.000 159.865 111.285 160.325 ;
        RECT 111.455 159.695 111.725 160.155 ;
        RECT 112.125 159.865 112.525 160.715 ;
        RECT 113.390 160.545 113.840 161.005 ;
        RECT 114.115 160.835 114.395 161.505 ;
        RECT 115.985 161.425 116.215 162.245 ;
        RECT 116.385 161.445 116.715 162.075 ;
        RECT 115.965 161.005 116.295 161.255 ;
        RECT 112.715 160.325 113.840 160.545 ;
        RECT 112.715 159.865 112.995 160.325 ;
        RECT 113.515 159.695 113.840 160.155 ;
        RECT 114.010 159.865 114.395 160.835 ;
        RECT 114.565 159.695 114.855 160.860 ;
        RECT 116.465 160.845 116.715 161.445 ;
        RECT 116.885 161.425 117.095 162.245 ;
        RECT 117.330 161.535 117.585 162.065 ;
        RECT 117.755 161.785 118.060 162.245 ;
        RECT 118.305 161.865 119.375 162.035 ;
        RECT 115.985 159.695 116.215 160.835 ;
        RECT 116.385 159.865 116.715 160.845 ;
        RECT 117.330 160.885 117.540 161.535 ;
        RECT 118.305 161.510 118.625 161.865 ;
        RECT 118.300 161.335 118.625 161.510 ;
        RECT 117.710 161.035 118.625 161.335 ;
        RECT 118.795 161.295 119.035 161.695 ;
        RECT 119.205 161.635 119.375 161.865 ;
        RECT 119.545 161.805 119.735 162.245 ;
        RECT 119.905 161.795 120.855 162.075 ;
        RECT 121.075 161.885 121.425 162.055 ;
        RECT 119.205 161.465 119.735 161.635 ;
        RECT 117.710 161.005 118.450 161.035 ;
        RECT 116.885 159.695 117.095 160.835 ;
        RECT 117.330 160.005 117.585 160.885 ;
        RECT 117.755 159.695 118.060 160.835 ;
        RECT 118.280 160.415 118.450 161.005 ;
        RECT 118.795 160.925 119.335 161.295 ;
        RECT 119.515 161.185 119.735 161.465 ;
        RECT 119.905 161.015 120.075 161.795 ;
        RECT 119.670 160.845 120.075 161.015 ;
        RECT 120.245 161.005 120.595 161.625 ;
        RECT 119.670 160.755 119.840 160.845 ;
        RECT 120.765 160.835 120.975 161.625 ;
        RECT 118.620 160.585 119.840 160.755 ;
        RECT 120.300 160.675 120.975 160.835 ;
        RECT 118.280 160.245 119.080 160.415 ;
        RECT 118.400 159.695 118.730 160.075 ;
        RECT 118.910 159.955 119.080 160.245 ;
        RECT 119.670 160.205 119.840 160.585 ;
        RECT 120.010 160.665 120.975 160.675 ;
        RECT 121.165 161.495 121.425 161.885 ;
        RECT 121.635 161.785 121.965 162.245 ;
        RECT 122.840 161.855 123.695 162.025 ;
        RECT 123.900 161.855 124.395 162.025 ;
        RECT 124.565 161.885 124.895 162.245 ;
        RECT 121.165 160.805 121.335 161.495 ;
        RECT 121.505 161.145 121.675 161.325 ;
        RECT 121.845 161.315 122.635 161.565 ;
        RECT 122.840 161.145 123.010 161.855 ;
        RECT 123.180 161.345 123.535 161.565 ;
        RECT 121.505 160.975 123.195 161.145 ;
        RECT 120.010 160.375 120.470 160.665 ;
        RECT 121.165 160.635 122.665 160.805 ;
        RECT 121.165 160.495 121.335 160.635 ;
        RECT 120.775 160.325 121.335 160.495 ;
        RECT 119.250 159.695 119.500 160.155 ;
        RECT 119.670 159.865 120.540 160.205 ;
        RECT 120.775 159.865 120.945 160.325 ;
        RECT 121.780 160.295 122.855 160.465 ;
        RECT 121.115 159.695 121.485 160.155 ;
        RECT 121.780 159.955 121.950 160.295 ;
        RECT 122.120 159.695 122.450 160.125 ;
        RECT 122.685 159.955 122.855 160.295 ;
        RECT 123.025 160.195 123.195 160.975 ;
        RECT 123.365 160.755 123.535 161.345 ;
        RECT 123.705 160.945 124.055 161.565 ;
        RECT 123.365 160.365 123.830 160.755 ;
        RECT 124.225 160.495 124.395 161.855 ;
        RECT 124.565 160.665 125.025 161.715 ;
        RECT 124.000 160.325 124.395 160.495 ;
        RECT 124.000 160.195 124.170 160.325 ;
        RECT 123.025 159.865 123.705 160.195 ;
        RECT 123.920 159.865 124.170 160.195 ;
        RECT 124.340 159.695 124.590 160.155 ;
        RECT 124.760 159.880 125.085 160.665 ;
        RECT 125.255 159.865 125.425 161.985 ;
        RECT 125.595 161.865 125.925 162.245 ;
        RECT 126.095 161.695 126.350 161.985 ;
        RECT 125.600 161.525 126.350 161.695 ;
        RECT 125.600 160.535 125.830 161.525 ;
        RECT 126.525 161.495 127.735 162.245 ;
        RECT 126.000 160.705 126.350 161.355 ;
        RECT 126.525 160.785 127.045 161.325 ;
        RECT 127.215 160.955 127.735 161.495 ;
        RECT 125.600 160.365 126.350 160.535 ;
        RECT 125.595 159.695 125.925 160.195 ;
        RECT 126.095 159.865 126.350 160.365 ;
        RECT 126.525 159.695 127.735 160.785 ;
        RECT 29.840 159.525 127.820 159.695 ;
        RECT 29.925 158.435 31.135 159.525 ;
        RECT 32.600 159.185 32.855 159.215 ;
        RECT 32.515 159.015 32.855 159.185 ;
        RECT 29.925 157.725 30.445 158.265 ;
        RECT 30.615 157.895 31.135 158.435 ;
        RECT 32.600 158.545 32.855 159.015 ;
        RECT 33.035 158.725 33.320 159.525 ;
        RECT 33.500 158.805 33.830 159.315 ;
        RECT 29.925 156.975 31.135 157.725 ;
        RECT 32.600 157.685 32.780 158.545 ;
        RECT 33.500 158.215 33.750 158.805 ;
        RECT 34.100 158.655 34.270 159.265 ;
        RECT 34.440 158.835 34.770 159.525 ;
        RECT 35.000 158.975 35.240 159.265 ;
        RECT 35.440 159.145 35.860 159.525 ;
        RECT 36.040 159.055 36.670 159.305 ;
        RECT 37.140 159.145 37.470 159.525 ;
        RECT 36.040 158.975 36.210 159.055 ;
        RECT 37.640 158.975 37.810 159.265 ;
        RECT 37.990 159.145 38.370 159.525 ;
        RECT 38.610 159.140 39.440 159.310 ;
        RECT 35.000 158.805 36.210 158.975 ;
        RECT 32.950 157.885 33.750 158.215 ;
        RECT 32.600 157.155 32.855 157.685 ;
        RECT 33.035 156.975 33.320 157.435 ;
        RECT 33.500 157.235 33.750 157.885 ;
        RECT 33.950 158.635 34.270 158.655 ;
        RECT 33.950 158.465 35.870 158.635 ;
        RECT 33.950 157.570 34.140 158.465 ;
        RECT 36.040 158.295 36.210 158.805 ;
        RECT 36.380 158.545 36.900 158.855 ;
        RECT 34.310 158.125 36.210 158.295 ;
        RECT 34.310 158.065 34.640 158.125 ;
        RECT 34.790 157.895 35.120 157.955 ;
        RECT 34.460 157.625 35.120 157.895 ;
        RECT 33.950 157.240 34.270 157.570 ;
        RECT 34.450 156.975 35.110 157.455 ;
        RECT 35.310 157.365 35.480 158.125 ;
        RECT 36.380 157.955 36.560 158.365 ;
        RECT 35.650 157.785 35.980 157.905 ;
        RECT 36.730 157.785 36.900 158.545 ;
        RECT 35.650 157.615 36.900 157.785 ;
        RECT 37.070 158.725 38.440 158.975 ;
        RECT 37.070 157.955 37.260 158.725 ;
        RECT 38.190 158.465 38.440 158.725 ;
        RECT 37.430 158.295 37.680 158.455 ;
        RECT 38.610 158.295 38.780 159.140 ;
        RECT 39.675 158.855 39.845 159.355 ;
        RECT 40.015 159.025 40.345 159.525 ;
        RECT 38.950 158.465 39.450 158.845 ;
        RECT 39.675 158.685 40.370 158.855 ;
        RECT 37.430 158.125 38.780 158.295 ;
        RECT 38.360 158.085 38.780 158.125 ;
        RECT 37.070 157.615 37.490 157.955 ;
        RECT 37.780 157.625 38.190 157.955 ;
        RECT 35.310 157.195 36.160 157.365 ;
        RECT 36.720 156.975 37.040 157.435 ;
        RECT 37.240 157.185 37.490 157.615 ;
        RECT 37.780 156.975 38.190 157.415 ;
        RECT 38.360 157.355 38.530 158.085 ;
        RECT 38.700 157.535 39.050 157.905 ;
        RECT 39.230 157.595 39.450 158.465 ;
        RECT 39.620 157.895 40.030 158.515 ;
        RECT 40.200 157.715 40.370 158.685 ;
        RECT 39.675 157.525 40.370 157.715 ;
        RECT 38.360 157.155 39.375 157.355 ;
        RECT 39.675 157.195 39.845 157.525 ;
        RECT 40.015 156.975 40.345 157.355 ;
        RECT 40.560 157.235 40.785 159.355 ;
        RECT 40.955 159.025 41.285 159.525 ;
        RECT 41.455 158.855 41.625 159.355 ;
        RECT 40.960 158.685 41.625 158.855 ;
        RECT 40.960 157.695 41.190 158.685 ;
        RECT 41.360 157.865 41.710 158.515 ;
        RECT 41.885 158.435 44.475 159.525 ;
        RECT 44.650 159.090 49.995 159.525 ;
        RECT 41.885 157.915 43.095 158.435 ;
        RECT 43.265 157.745 44.475 158.265 ;
        RECT 46.240 157.840 46.590 159.090 ;
        RECT 50.165 158.360 50.455 159.525 ;
        RECT 51.085 158.435 52.755 159.525 ;
        RECT 40.960 157.525 41.625 157.695 ;
        RECT 40.955 156.975 41.285 157.355 ;
        RECT 41.455 157.235 41.625 157.525 ;
        RECT 41.885 156.975 44.475 157.745 ;
        RECT 48.070 157.520 48.410 158.350 ;
        RECT 51.085 157.915 51.835 158.435 ;
        RECT 52.925 158.385 53.195 159.355 ;
        RECT 53.405 158.725 53.685 159.525 ;
        RECT 53.855 159.015 55.510 159.305 ;
        RECT 53.920 158.675 55.510 158.845 ;
        RECT 53.920 158.555 54.090 158.675 ;
        RECT 53.365 158.385 54.090 158.555 ;
        RECT 52.005 157.745 52.755 158.265 ;
        RECT 44.650 156.975 49.995 157.520 ;
        RECT 50.165 156.975 50.455 157.700 ;
        RECT 51.085 156.975 52.755 157.745 ;
        RECT 52.925 157.650 53.095 158.385 ;
        RECT 53.365 158.215 53.535 158.385 ;
        RECT 54.280 158.335 54.995 158.505 ;
        RECT 55.190 158.385 55.510 158.675 ;
        RECT 55.685 158.435 59.195 159.525 ;
        RECT 53.265 157.885 53.535 158.215 ;
        RECT 53.705 157.885 54.110 158.215 ;
        RECT 54.280 157.885 54.990 158.335 ;
        RECT 53.365 157.715 53.535 157.885 ;
        RECT 52.925 157.305 53.195 157.650 ;
        RECT 53.365 157.545 54.975 157.715 ;
        RECT 55.160 157.645 55.510 158.215 ;
        RECT 55.685 157.915 57.375 158.435 ;
        RECT 59.365 158.385 59.705 159.355 ;
        RECT 59.875 158.385 60.045 159.525 ;
        RECT 60.315 158.725 60.565 159.525 ;
        RECT 61.210 158.555 61.540 159.355 ;
        RECT 61.840 158.725 62.170 159.525 ;
        RECT 62.340 158.555 62.670 159.355 ;
        RECT 60.235 158.385 62.670 158.555 ;
        RECT 63.420 158.545 63.675 159.215 ;
        RECT 63.855 158.725 64.140 159.525 ;
        RECT 64.320 158.805 64.650 159.315 ;
        RECT 57.545 157.745 59.195 158.265 ;
        RECT 53.385 156.975 53.765 157.375 ;
        RECT 53.935 157.195 54.105 157.545 ;
        RECT 54.275 156.975 54.605 157.375 ;
        RECT 54.805 157.195 54.975 157.545 ;
        RECT 55.175 156.975 55.505 157.475 ;
        RECT 55.685 156.975 59.195 157.745 ;
        RECT 59.365 157.775 59.540 158.385 ;
        RECT 60.235 158.135 60.405 158.385 ;
        RECT 59.710 157.965 60.405 158.135 ;
        RECT 60.580 157.965 61.000 158.165 ;
        RECT 61.170 157.965 61.500 158.165 ;
        RECT 61.670 157.965 62.000 158.165 ;
        RECT 59.365 157.145 59.705 157.775 ;
        RECT 59.875 156.975 60.125 157.775 ;
        RECT 60.315 157.625 61.540 157.795 ;
        RECT 60.315 157.145 60.645 157.625 ;
        RECT 60.815 156.975 61.040 157.435 ;
        RECT 61.210 157.145 61.540 157.625 ;
        RECT 62.170 157.755 62.340 158.385 ;
        RECT 62.525 157.965 62.875 158.215 ;
        RECT 63.420 157.825 63.600 158.545 ;
        RECT 64.320 158.215 64.570 158.805 ;
        RECT 64.920 158.655 65.090 159.265 ;
        RECT 65.260 158.835 65.590 159.525 ;
        RECT 65.820 158.975 66.060 159.265 ;
        RECT 66.260 159.145 66.680 159.525 ;
        RECT 66.860 159.055 67.490 159.305 ;
        RECT 67.960 159.145 68.290 159.525 ;
        RECT 66.860 158.975 67.030 159.055 ;
        RECT 68.460 158.975 68.630 159.265 ;
        RECT 68.810 159.145 69.190 159.525 ;
        RECT 69.430 159.140 70.260 159.310 ;
        RECT 65.820 158.805 67.030 158.975 ;
        RECT 63.770 157.885 64.570 158.215 ;
        RECT 62.170 157.145 62.670 157.755 ;
        RECT 63.335 157.685 63.600 157.825 ;
        RECT 63.335 157.655 63.675 157.685 ;
        RECT 63.420 157.155 63.675 157.655 ;
        RECT 63.855 156.975 64.140 157.435 ;
        RECT 64.320 157.235 64.570 157.885 ;
        RECT 64.770 158.635 65.090 158.655 ;
        RECT 64.770 158.465 66.690 158.635 ;
        RECT 64.770 157.570 64.960 158.465 ;
        RECT 66.860 158.295 67.030 158.805 ;
        RECT 67.200 158.545 67.720 158.855 ;
        RECT 65.130 158.125 67.030 158.295 ;
        RECT 65.130 158.065 65.460 158.125 ;
        RECT 65.610 157.895 65.940 157.955 ;
        RECT 65.280 157.625 65.940 157.895 ;
        RECT 64.770 157.240 65.090 157.570 ;
        RECT 65.270 156.975 65.930 157.455 ;
        RECT 66.130 157.365 66.300 158.125 ;
        RECT 67.200 157.955 67.380 158.365 ;
        RECT 66.470 157.785 66.800 157.905 ;
        RECT 67.550 157.785 67.720 158.545 ;
        RECT 66.470 157.615 67.720 157.785 ;
        RECT 67.890 158.725 69.260 158.975 ;
        RECT 67.890 157.955 68.080 158.725 ;
        RECT 69.010 158.465 69.260 158.725 ;
        RECT 68.250 158.295 68.500 158.455 ;
        RECT 69.430 158.295 69.600 159.140 ;
        RECT 70.495 158.855 70.665 159.355 ;
        RECT 70.835 159.025 71.165 159.525 ;
        RECT 69.770 158.465 70.270 158.845 ;
        RECT 70.495 158.685 71.190 158.855 ;
        RECT 68.250 158.125 69.600 158.295 ;
        RECT 69.180 158.085 69.600 158.125 ;
        RECT 67.890 157.615 68.310 157.955 ;
        RECT 68.600 157.625 69.010 157.955 ;
        RECT 66.130 157.195 66.980 157.365 ;
        RECT 67.540 156.975 67.860 157.435 ;
        RECT 68.060 157.185 68.310 157.615 ;
        RECT 68.600 156.975 69.010 157.415 ;
        RECT 69.180 157.355 69.350 158.085 ;
        RECT 69.520 157.535 69.870 157.905 ;
        RECT 70.050 157.595 70.270 158.465 ;
        RECT 70.440 157.895 70.850 158.515 ;
        RECT 71.020 157.715 71.190 158.685 ;
        RECT 70.495 157.525 71.190 157.715 ;
        RECT 69.180 157.155 70.195 157.355 ;
        RECT 70.495 157.195 70.665 157.525 ;
        RECT 70.835 156.975 71.165 157.355 ;
        RECT 71.380 157.235 71.605 159.355 ;
        RECT 71.775 159.025 72.105 159.525 ;
        RECT 72.275 158.855 72.445 159.355 ;
        RECT 71.780 158.685 72.445 158.855 ;
        RECT 71.780 157.695 72.010 158.685 ;
        RECT 72.180 157.865 72.530 158.515 ;
        RECT 73.165 158.435 75.755 159.525 ;
        RECT 73.165 157.915 74.375 158.435 ;
        RECT 75.925 158.360 76.215 159.525 ;
        RECT 76.390 158.375 76.650 159.525 ;
        RECT 76.825 158.450 77.080 159.355 ;
        RECT 77.250 158.765 77.580 159.525 ;
        RECT 77.795 158.595 77.965 159.355 ;
        RECT 74.545 157.745 75.755 158.265 ;
        RECT 71.780 157.525 72.445 157.695 ;
        RECT 71.775 156.975 72.105 157.355 ;
        RECT 72.275 157.235 72.445 157.525 ;
        RECT 73.165 156.975 75.755 157.745 ;
        RECT 75.925 156.975 76.215 157.700 ;
        RECT 76.390 156.975 76.650 157.815 ;
        RECT 76.825 157.720 76.995 158.450 ;
        RECT 77.250 158.425 77.965 158.595 ;
        RECT 78.315 158.595 78.485 159.355 ;
        RECT 78.700 158.765 79.030 159.525 ;
        RECT 78.315 158.425 79.030 158.595 ;
        RECT 79.200 158.450 79.455 159.355 ;
        RECT 77.250 158.215 77.420 158.425 ;
        RECT 77.165 157.885 77.420 158.215 ;
        RECT 76.825 157.145 77.080 157.720 ;
        RECT 77.250 157.695 77.420 157.885 ;
        RECT 77.700 157.875 78.055 158.245 ;
        RECT 78.225 157.875 78.580 158.245 ;
        RECT 78.860 158.215 79.030 158.425 ;
        RECT 78.860 157.885 79.115 158.215 ;
        RECT 78.860 157.695 79.030 157.885 ;
        RECT 79.285 157.720 79.455 158.450 ;
        RECT 79.630 158.375 79.890 159.525 ;
        RECT 80.075 158.465 80.405 159.525 ;
        RECT 80.585 158.215 80.755 159.140 ;
        RECT 80.925 158.935 81.255 159.335 ;
        RECT 81.425 159.165 81.755 159.525 ;
        RECT 81.955 158.935 82.655 159.355 ;
        RECT 80.925 158.705 82.655 158.935 ;
        RECT 80.925 158.485 81.255 158.705 ;
        RECT 81.450 158.215 81.775 158.505 ;
        RECT 80.065 157.885 80.375 158.215 ;
        RECT 80.585 157.885 80.960 158.215 ;
        RECT 81.280 157.885 81.775 158.215 ;
        RECT 81.950 157.965 82.280 158.505 ;
        RECT 77.250 157.525 77.965 157.695 ;
        RECT 77.250 156.975 77.580 157.355 ;
        RECT 77.795 157.145 77.965 157.525 ;
        RECT 78.315 157.525 79.030 157.695 ;
        RECT 78.315 157.145 78.485 157.525 ;
        RECT 78.700 156.975 79.030 157.355 ;
        RECT 79.200 157.145 79.455 157.720 ;
        RECT 79.630 156.975 79.890 157.815 ;
        RECT 82.450 157.735 82.655 158.705 ;
        RECT 80.075 157.505 81.435 157.715 ;
        RECT 80.075 157.145 80.405 157.505 ;
        RECT 80.575 156.975 80.905 157.335 ;
        RECT 81.105 157.145 81.435 157.505 ;
        RECT 81.945 157.145 82.655 157.735 ;
        RECT 82.825 158.385 83.095 159.355 ;
        RECT 83.305 158.725 83.585 159.525 ;
        RECT 83.755 159.015 85.410 159.305 ;
        RECT 83.820 158.675 85.410 158.845 ;
        RECT 83.820 158.555 83.990 158.675 ;
        RECT 83.265 158.385 83.990 158.555 ;
        RECT 82.825 157.650 82.995 158.385 ;
        RECT 83.265 158.215 83.435 158.385 ;
        RECT 84.180 158.335 84.895 158.505 ;
        RECT 85.090 158.385 85.410 158.675 ;
        RECT 86.045 158.435 87.715 159.525 ;
        RECT 88.260 158.545 88.515 159.215 ;
        RECT 88.695 158.725 88.980 159.525 ;
        RECT 89.160 158.805 89.490 159.315 ;
        RECT 83.165 157.885 83.435 158.215 ;
        RECT 83.605 157.885 84.010 158.215 ;
        RECT 84.180 157.885 84.890 158.335 ;
        RECT 83.265 157.715 83.435 157.885 ;
        RECT 82.825 157.305 83.095 157.650 ;
        RECT 83.265 157.545 84.875 157.715 ;
        RECT 85.060 157.645 85.410 158.215 ;
        RECT 86.045 157.915 86.795 158.435 ;
        RECT 86.965 157.745 87.715 158.265 ;
        RECT 83.285 156.975 83.665 157.375 ;
        RECT 83.835 157.195 84.005 157.545 ;
        RECT 84.175 156.975 84.505 157.375 ;
        RECT 84.705 157.195 84.875 157.545 ;
        RECT 85.075 156.975 85.405 157.475 ;
        RECT 86.045 156.975 87.715 157.745 ;
        RECT 88.260 157.685 88.440 158.545 ;
        RECT 89.160 158.215 89.410 158.805 ;
        RECT 89.760 158.655 89.930 159.265 ;
        RECT 90.100 158.835 90.430 159.525 ;
        RECT 90.660 158.975 90.900 159.265 ;
        RECT 91.100 159.145 91.520 159.525 ;
        RECT 91.700 159.055 92.330 159.305 ;
        RECT 92.800 159.145 93.130 159.525 ;
        RECT 91.700 158.975 91.870 159.055 ;
        RECT 93.300 158.975 93.470 159.265 ;
        RECT 93.650 159.145 94.030 159.525 ;
        RECT 94.270 159.140 95.100 159.310 ;
        RECT 90.660 158.805 91.870 158.975 ;
        RECT 88.610 157.885 89.410 158.215 ;
        RECT 88.260 157.485 88.515 157.685 ;
        RECT 88.175 157.315 88.515 157.485 ;
        RECT 88.260 157.155 88.515 157.315 ;
        RECT 88.695 156.975 88.980 157.435 ;
        RECT 89.160 157.235 89.410 157.885 ;
        RECT 89.610 158.635 89.930 158.655 ;
        RECT 89.610 158.465 91.530 158.635 ;
        RECT 89.610 157.570 89.800 158.465 ;
        RECT 91.700 158.295 91.870 158.805 ;
        RECT 92.040 158.545 92.560 158.855 ;
        RECT 89.970 158.125 91.870 158.295 ;
        RECT 89.970 158.065 90.300 158.125 ;
        RECT 90.450 157.895 90.780 157.955 ;
        RECT 90.120 157.625 90.780 157.895 ;
        RECT 89.610 157.240 89.930 157.570 ;
        RECT 90.110 156.975 90.770 157.455 ;
        RECT 90.970 157.365 91.140 158.125 ;
        RECT 92.040 157.955 92.220 158.365 ;
        RECT 91.310 157.785 91.640 157.905 ;
        RECT 92.390 157.785 92.560 158.545 ;
        RECT 91.310 157.615 92.560 157.785 ;
        RECT 92.730 158.725 94.100 158.975 ;
        RECT 92.730 157.955 92.920 158.725 ;
        RECT 93.850 158.465 94.100 158.725 ;
        RECT 93.090 158.295 93.340 158.455 ;
        RECT 94.270 158.295 94.440 159.140 ;
        RECT 95.335 158.855 95.505 159.355 ;
        RECT 95.675 159.025 96.005 159.525 ;
        RECT 94.610 158.465 95.110 158.845 ;
        RECT 95.335 158.685 96.030 158.855 ;
        RECT 93.090 158.125 94.440 158.295 ;
        RECT 94.020 158.085 94.440 158.125 ;
        RECT 92.730 157.615 93.150 157.955 ;
        RECT 93.440 157.625 93.850 157.955 ;
        RECT 90.970 157.195 91.820 157.365 ;
        RECT 92.380 156.975 92.700 157.435 ;
        RECT 92.900 157.185 93.150 157.615 ;
        RECT 93.440 156.975 93.850 157.415 ;
        RECT 94.020 157.355 94.190 158.085 ;
        RECT 94.360 157.535 94.710 157.905 ;
        RECT 94.890 157.595 95.110 158.465 ;
        RECT 95.280 157.895 95.690 158.515 ;
        RECT 95.860 157.715 96.030 158.685 ;
        RECT 95.335 157.525 96.030 157.715 ;
        RECT 94.020 157.155 95.035 157.355 ;
        RECT 95.335 157.195 95.505 157.525 ;
        RECT 95.675 156.975 96.005 157.355 ;
        RECT 96.220 157.235 96.445 159.355 ;
        RECT 96.615 159.025 96.945 159.525 ;
        RECT 97.115 158.855 97.285 159.355 ;
        RECT 96.620 158.685 97.285 158.855 ;
        RECT 96.620 157.695 96.850 158.685 ;
        RECT 97.020 157.865 97.370 158.515 ;
        RECT 97.545 158.435 99.215 159.525 ;
        RECT 97.545 157.915 98.295 158.435 ;
        RECT 99.445 158.385 99.655 159.525 ;
        RECT 99.825 158.375 100.155 159.355 ;
        RECT 100.325 158.385 100.555 159.525 ;
        RECT 98.465 157.745 99.215 158.265 ;
        RECT 96.620 157.525 97.285 157.695 ;
        RECT 96.615 156.975 96.945 157.355 ;
        RECT 97.115 157.235 97.285 157.525 ;
        RECT 97.545 156.975 99.215 157.745 ;
        RECT 99.445 156.975 99.655 157.795 ;
        RECT 99.825 157.775 100.075 158.375 ;
        RECT 101.685 158.360 101.975 159.525 ;
        RECT 102.145 158.435 105.655 159.525 ;
        RECT 100.245 157.965 100.575 158.215 ;
        RECT 102.145 157.915 103.835 158.435 ;
        RECT 105.825 158.385 106.095 159.355 ;
        RECT 106.305 158.725 106.585 159.525 ;
        RECT 106.755 159.015 108.410 159.305 ;
        RECT 106.820 158.675 108.410 158.845 ;
        RECT 106.820 158.555 106.990 158.675 ;
        RECT 106.265 158.385 106.990 158.555 ;
        RECT 99.825 157.145 100.155 157.775 ;
        RECT 100.325 156.975 100.555 157.795 ;
        RECT 104.005 157.745 105.655 158.265 ;
        RECT 101.685 156.975 101.975 157.700 ;
        RECT 102.145 156.975 105.655 157.745 ;
        RECT 105.825 157.650 105.995 158.385 ;
        RECT 106.265 158.215 106.435 158.385 ;
        RECT 107.180 158.335 107.895 158.505 ;
        RECT 108.090 158.385 108.410 158.675 ;
        RECT 108.585 158.385 108.925 159.355 ;
        RECT 109.095 158.385 109.265 159.525 ;
        RECT 109.535 158.725 109.785 159.525 ;
        RECT 110.430 158.555 110.760 159.355 ;
        RECT 111.060 158.725 111.390 159.525 ;
        RECT 111.560 158.555 111.890 159.355 ;
        RECT 109.455 158.385 111.890 158.555 ;
        RECT 113.190 158.385 113.525 159.355 ;
        RECT 113.695 158.385 113.865 159.525 ;
        RECT 114.035 159.185 116.065 159.355 ;
        RECT 106.165 157.885 106.435 158.215 ;
        RECT 106.605 157.885 107.010 158.215 ;
        RECT 107.180 157.885 107.890 158.335 ;
        RECT 106.265 157.715 106.435 157.885 ;
        RECT 105.825 157.305 106.095 157.650 ;
        RECT 106.265 157.545 107.875 157.715 ;
        RECT 108.060 157.645 108.410 158.215 ;
        RECT 108.585 157.825 108.760 158.385 ;
        RECT 109.455 158.135 109.625 158.385 ;
        RECT 108.930 157.965 109.625 158.135 ;
        RECT 109.800 157.965 110.220 158.165 ;
        RECT 110.390 157.965 110.720 158.165 ;
        RECT 110.890 157.965 111.220 158.165 ;
        RECT 108.585 157.775 108.815 157.825 ;
        RECT 106.285 156.975 106.665 157.375 ;
        RECT 106.835 157.195 107.005 157.545 ;
        RECT 107.175 156.975 107.505 157.375 ;
        RECT 107.705 157.195 107.875 157.545 ;
        RECT 108.075 156.975 108.405 157.475 ;
        RECT 108.585 157.145 108.925 157.775 ;
        RECT 109.095 156.975 109.345 157.775 ;
        RECT 109.535 157.625 110.760 157.795 ;
        RECT 109.535 157.145 109.865 157.625 ;
        RECT 110.035 156.975 110.260 157.435 ;
        RECT 110.430 157.145 110.760 157.625 ;
        RECT 111.390 157.755 111.560 158.385 ;
        RECT 111.745 157.965 112.095 158.215 ;
        RECT 111.390 157.145 111.890 157.755 ;
        RECT 113.190 157.715 113.360 158.385 ;
        RECT 114.035 158.215 114.205 159.185 ;
        RECT 113.530 157.885 113.785 158.215 ;
        RECT 114.010 157.885 114.205 158.215 ;
        RECT 114.375 158.845 115.500 159.015 ;
        RECT 113.615 157.715 113.785 157.885 ;
        RECT 114.375 157.715 114.545 158.845 ;
        RECT 113.190 157.145 113.445 157.715 ;
        RECT 113.615 157.545 114.545 157.715 ;
        RECT 114.715 158.505 115.725 158.675 ;
        RECT 114.715 157.705 114.885 158.505 ;
        RECT 115.090 158.165 115.365 158.305 ;
        RECT 115.085 157.995 115.365 158.165 ;
        RECT 114.370 157.510 114.545 157.545 ;
        RECT 113.615 156.975 113.945 157.375 ;
        RECT 114.370 157.145 114.900 157.510 ;
        RECT 115.090 157.145 115.365 157.995 ;
        RECT 115.535 157.145 115.725 158.505 ;
        RECT 115.895 158.520 116.065 159.185 ;
        RECT 116.235 158.765 116.405 159.525 ;
        RECT 116.640 158.765 117.155 159.175 ;
        RECT 115.895 158.330 116.645 158.520 ;
        RECT 116.815 157.955 117.155 158.765 ;
        RECT 115.925 157.785 117.155 157.955 ;
        RECT 117.325 158.765 117.840 159.175 ;
        RECT 118.075 158.765 118.245 159.525 ;
        RECT 118.415 159.185 120.445 159.355 ;
        RECT 117.325 157.955 117.665 158.765 ;
        RECT 118.415 158.520 118.585 159.185 ;
        RECT 118.980 158.845 120.105 159.015 ;
        RECT 117.835 158.330 118.585 158.520 ;
        RECT 118.755 158.505 119.765 158.675 ;
        RECT 117.325 157.785 118.555 157.955 ;
        RECT 115.905 156.975 116.415 157.510 ;
        RECT 116.635 157.180 116.880 157.785 ;
        RECT 117.600 157.180 117.845 157.785 ;
        RECT 118.065 156.975 118.575 157.510 ;
        RECT 118.755 157.145 118.945 158.505 ;
        RECT 119.115 158.165 119.390 158.305 ;
        RECT 119.115 157.995 119.395 158.165 ;
        RECT 119.115 157.145 119.390 157.995 ;
        RECT 119.595 157.705 119.765 158.505 ;
        RECT 119.935 157.715 120.105 158.845 ;
        RECT 120.275 158.215 120.445 159.185 ;
        RECT 120.615 158.385 120.785 159.525 ;
        RECT 120.955 158.385 121.290 159.355 ;
        RECT 122.475 158.595 122.645 159.355 ;
        RECT 122.825 158.765 123.155 159.525 ;
        RECT 122.475 158.425 123.140 158.595 ;
        RECT 123.325 158.450 123.595 159.355 ;
        RECT 120.275 157.885 120.470 158.215 ;
        RECT 120.695 157.885 120.950 158.215 ;
        RECT 120.695 157.715 120.865 157.885 ;
        RECT 121.120 157.715 121.290 158.385 ;
        RECT 122.970 158.280 123.140 158.425 ;
        RECT 122.405 157.875 122.735 158.245 ;
        RECT 122.970 157.950 123.255 158.280 ;
        RECT 119.935 157.545 120.865 157.715 ;
        RECT 119.935 157.510 120.110 157.545 ;
        RECT 119.580 157.145 120.110 157.510 ;
        RECT 120.535 156.975 120.865 157.375 ;
        RECT 121.035 157.145 121.290 157.715 ;
        RECT 122.970 157.695 123.140 157.950 ;
        RECT 122.475 157.525 123.140 157.695 ;
        RECT 123.425 157.650 123.595 158.450 ;
        RECT 123.855 158.595 124.025 159.355 ;
        RECT 124.205 158.765 124.535 159.525 ;
        RECT 123.855 158.425 124.520 158.595 ;
        RECT 124.705 158.450 124.975 159.355 ;
        RECT 124.350 158.280 124.520 158.425 ;
        RECT 123.785 157.875 124.115 158.245 ;
        RECT 124.350 157.950 124.635 158.280 ;
        RECT 124.350 157.695 124.520 157.950 ;
        RECT 122.475 157.145 122.645 157.525 ;
        RECT 122.825 156.975 123.155 157.355 ;
        RECT 123.335 157.145 123.595 157.650 ;
        RECT 123.855 157.525 124.520 157.695 ;
        RECT 124.805 157.650 124.975 158.450 ;
        RECT 125.145 158.435 126.355 159.525 ;
        RECT 126.525 158.435 127.735 159.525 ;
        RECT 125.145 157.895 125.665 158.435 ;
        RECT 125.835 157.725 126.355 158.265 ;
        RECT 126.525 157.895 127.045 158.435 ;
        RECT 127.215 157.725 127.735 158.265 ;
        RECT 123.855 157.145 124.025 157.525 ;
        RECT 124.205 156.975 124.535 157.355 ;
        RECT 124.715 157.145 124.975 157.650 ;
        RECT 125.145 156.975 126.355 157.725 ;
        RECT 126.525 156.975 127.735 157.725 ;
        RECT 29.840 156.805 127.820 156.975 ;
        RECT 29.925 156.055 31.135 156.805 ;
        RECT 29.925 155.515 30.445 156.055 ;
        RECT 31.305 156.035 33.895 156.805 ;
        RECT 30.615 155.345 31.135 155.885 ;
        RECT 29.925 154.255 31.135 155.345 ;
        RECT 31.305 155.345 32.515 155.865 ;
        RECT 32.685 155.515 33.895 156.035 ;
        RECT 34.105 155.985 34.335 156.805 ;
        RECT 34.505 156.005 34.835 156.635 ;
        RECT 34.085 155.565 34.415 155.815 ;
        RECT 34.585 155.405 34.835 156.005 ;
        RECT 35.005 155.985 35.215 156.805 ;
        RECT 35.445 156.035 37.115 156.805 ;
        RECT 37.285 156.080 37.575 156.805 ;
        RECT 37.835 156.255 38.005 156.635 ;
        RECT 38.185 156.425 38.515 156.805 ;
        RECT 37.835 156.085 38.500 156.255 ;
        RECT 38.695 156.130 38.955 156.635 ;
        RECT 40.050 156.260 45.395 156.805 ;
        RECT 31.305 154.255 33.895 155.345 ;
        RECT 34.105 154.255 34.335 155.395 ;
        RECT 34.505 154.425 34.835 155.405 ;
        RECT 35.005 154.255 35.215 155.395 ;
        RECT 35.445 155.345 36.195 155.865 ;
        RECT 36.365 155.515 37.115 156.035 ;
        RECT 37.765 155.535 38.095 155.905 ;
        RECT 38.330 155.830 38.500 156.085 ;
        RECT 38.330 155.500 38.615 155.830 ;
        RECT 35.445 154.255 37.115 155.345 ;
        RECT 37.285 154.255 37.575 155.420 ;
        RECT 38.330 155.355 38.500 155.500 ;
        RECT 37.835 155.185 38.500 155.355 ;
        RECT 38.785 155.330 38.955 156.130 ;
        RECT 37.835 154.425 38.005 155.185 ;
        RECT 38.185 154.255 38.515 155.015 ;
        RECT 38.685 154.425 38.955 155.330 ;
        RECT 41.640 154.690 41.990 155.940 ;
        RECT 43.470 155.430 43.810 156.260 ;
        RECT 45.565 156.130 45.835 156.475 ;
        RECT 46.025 156.405 46.405 156.805 ;
        RECT 46.575 156.235 46.745 156.585 ;
        RECT 46.915 156.405 47.245 156.805 ;
        RECT 47.445 156.235 47.615 156.585 ;
        RECT 47.815 156.305 48.145 156.805 ;
        RECT 45.565 155.395 45.735 156.130 ;
        RECT 46.005 156.065 47.615 156.235 ;
        RECT 46.005 155.895 46.175 156.065 ;
        RECT 45.905 155.565 46.175 155.895 ;
        RECT 46.345 155.565 46.750 155.895 ;
        RECT 46.005 155.395 46.175 155.565 ;
        RECT 40.050 154.255 45.395 154.690 ;
        RECT 45.565 154.425 45.835 155.395 ;
        RECT 46.005 155.225 46.730 155.395 ;
        RECT 46.920 155.275 47.630 155.895 ;
        RECT 47.800 155.565 48.150 156.135 ;
        RECT 48.325 156.005 48.665 156.635 ;
        RECT 48.835 156.005 49.085 156.805 ;
        RECT 49.275 156.155 49.605 156.635 ;
        RECT 49.775 156.345 50.000 156.805 ;
        RECT 50.170 156.155 50.500 156.635 ;
        RECT 48.325 155.955 48.555 156.005 ;
        RECT 49.275 155.985 50.500 156.155 ;
        RECT 51.130 156.025 51.630 156.635 ;
        RECT 52.380 156.465 52.635 156.625 ;
        RECT 52.295 156.295 52.635 156.465 ;
        RECT 52.815 156.345 53.100 156.805 ;
        RECT 52.380 156.095 52.635 156.295 ;
        RECT 48.325 155.395 48.500 155.955 ;
        RECT 48.670 155.645 49.365 155.815 ;
        RECT 49.195 155.395 49.365 155.645 ;
        RECT 49.540 155.615 49.960 155.815 ;
        RECT 50.130 155.615 50.460 155.815 ;
        RECT 50.630 155.615 50.960 155.815 ;
        RECT 51.130 155.395 51.300 156.025 ;
        RECT 51.485 155.565 51.835 155.815 ;
        RECT 46.560 155.105 46.730 155.225 ;
        RECT 47.830 155.105 48.150 155.395 ;
        RECT 46.045 154.255 46.325 155.055 ;
        RECT 46.560 154.935 48.150 155.105 ;
        RECT 46.495 154.475 48.150 154.765 ;
        RECT 48.325 154.425 48.665 155.395 ;
        RECT 48.835 154.255 49.005 155.395 ;
        RECT 49.195 155.225 51.630 155.395 ;
        RECT 49.275 154.255 49.525 155.055 ;
        RECT 50.170 154.425 50.500 155.225 ;
        RECT 50.800 154.255 51.130 155.055 ;
        RECT 51.300 154.425 51.630 155.225 ;
        RECT 52.380 155.235 52.560 156.095 ;
        RECT 53.280 155.895 53.530 156.545 ;
        RECT 52.730 155.565 53.530 155.895 ;
        RECT 52.380 154.565 52.635 155.235 ;
        RECT 52.815 154.255 53.100 155.055 ;
        RECT 53.280 154.975 53.530 155.565 ;
        RECT 53.730 156.210 54.050 156.540 ;
        RECT 54.230 156.325 54.890 156.805 ;
        RECT 55.090 156.415 55.940 156.585 ;
        RECT 53.730 155.315 53.920 156.210 ;
        RECT 54.240 155.885 54.900 156.155 ;
        RECT 54.570 155.825 54.900 155.885 ;
        RECT 54.090 155.655 54.420 155.715 ;
        RECT 55.090 155.655 55.260 156.415 ;
        RECT 56.500 156.345 56.820 156.805 ;
        RECT 57.020 156.165 57.270 156.595 ;
        RECT 57.560 156.365 57.970 156.805 ;
        RECT 58.140 156.425 59.155 156.625 ;
        RECT 55.430 155.995 56.680 156.165 ;
        RECT 55.430 155.875 55.760 155.995 ;
        RECT 54.090 155.485 55.990 155.655 ;
        RECT 53.730 155.145 55.650 155.315 ;
        RECT 53.730 155.125 54.050 155.145 ;
        RECT 53.280 154.465 53.610 154.975 ;
        RECT 53.880 154.515 54.050 155.125 ;
        RECT 55.820 154.975 55.990 155.485 ;
        RECT 56.160 155.415 56.340 155.825 ;
        RECT 56.510 155.235 56.680 155.995 ;
        RECT 54.220 154.255 54.550 154.945 ;
        RECT 54.780 154.805 55.990 154.975 ;
        RECT 56.160 154.925 56.680 155.235 ;
        RECT 56.850 155.825 57.270 156.165 ;
        RECT 57.560 155.825 57.970 156.155 ;
        RECT 56.850 155.055 57.040 155.825 ;
        RECT 58.140 155.695 58.310 156.425 ;
        RECT 59.455 156.255 59.625 156.585 ;
        RECT 59.795 156.425 60.125 156.805 ;
        RECT 58.480 155.875 58.830 156.245 ;
        RECT 58.140 155.655 58.560 155.695 ;
        RECT 57.210 155.485 58.560 155.655 ;
        RECT 57.210 155.325 57.460 155.485 ;
        RECT 57.970 155.055 58.220 155.315 ;
        RECT 56.850 154.805 58.220 155.055 ;
        RECT 54.780 154.515 55.020 154.805 ;
        RECT 55.820 154.725 55.990 154.805 ;
        RECT 55.220 154.255 55.640 154.635 ;
        RECT 55.820 154.475 56.450 154.725 ;
        RECT 56.920 154.255 57.250 154.635 ;
        RECT 57.420 154.515 57.590 154.805 ;
        RECT 58.390 154.640 58.560 155.485 ;
        RECT 59.010 155.315 59.230 156.185 ;
        RECT 59.455 156.065 60.150 156.255 ;
        RECT 58.730 154.935 59.230 155.315 ;
        RECT 59.400 155.265 59.810 155.885 ;
        RECT 59.980 155.095 60.150 156.065 ;
        RECT 59.455 154.925 60.150 155.095 ;
        RECT 57.770 154.255 58.150 154.635 ;
        RECT 58.390 154.470 59.220 154.640 ;
        RECT 59.455 154.425 59.625 154.925 ;
        RECT 59.795 154.255 60.125 154.755 ;
        RECT 60.340 154.425 60.565 156.545 ;
        RECT 60.735 156.425 61.065 156.805 ;
        RECT 61.235 156.255 61.405 156.545 ;
        RECT 60.740 156.085 61.405 156.255 ;
        RECT 60.740 155.095 60.970 156.085 ;
        RECT 61.725 155.985 61.935 156.805 ;
        RECT 62.105 156.005 62.435 156.635 ;
        RECT 61.140 155.265 61.490 155.915 ;
        RECT 62.105 155.405 62.355 156.005 ;
        RECT 62.605 155.985 62.835 156.805 ;
        RECT 63.045 156.080 63.335 156.805 ;
        RECT 63.780 155.995 64.025 156.600 ;
        RECT 64.245 156.270 64.755 156.805 ;
        RECT 63.505 155.825 64.735 155.995 ;
        RECT 62.525 155.565 62.855 155.815 ;
        RECT 60.740 154.925 61.405 155.095 ;
        RECT 60.735 154.255 61.065 154.755 ;
        RECT 61.235 154.425 61.405 154.925 ;
        RECT 61.725 154.255 61.935 155.395 ;
        RECT 62.105 154.425 62.435 155.405 ;
        RECT 62.605 154.255 62.835 155.395 ;
        RECT 63.045 154.255 63.335 155.420 ;
        RECT 63.505 155.015 63.845 155.825 ;
        RECT 64.015 155.260 64.765 155.450 ;
        RECT 63.505 154.605 64.020 155.015 ;
        RECT 64.255 154.255 64.425 155.015 ;
        RECT 64.595 154.595 64.765 155.260 ;
        RECT 64.935 155.275 65.125 156.635 ;
        RECT 65.295 156.125 65.570 156.635 ;
        RECT 65.760 156.270 66.290 156.635 ;
        RECT 66.715 156.405 67.045 156.805 ;
        RECT 66.115 156.235 66.290 156.270 ;
        RECT 65.295 155.955 65.575 156.125 ;
        RECT 65.295 155.475 65.570 155.955 ;
        RECT 65.775 155.275 65.945 156.075 ;
        RECT 64.935 155.105 65.945 155.275 ;
        RECT 66.115 156.065 67.045 156.235 ;
        RECT 67.215 156.065 67.470 156.635 ;
        RECT 66.115 154.935 66.285 156.065 ;
        RECT 66.875 155.895 67.045 156.065 ;
        RECT 65.160 154.765 66.285 154.935 ;
        RECT 66.455 155.565 66.650 155.895 ;
        RECT 66.875 155.565 67.130 155.895 ;
        RECT 66.455 154.595 66.625 155.565 ;
        RECT 67.300 155.395 67.470 156.065 ;
        RECT 68.840 155.995 69.085 156.600 ;
        RECT 69.305 156.270 69.815 156.805 ;
        RECT 64.595 154.425 66.625 154.595 ;
        RECT 66.795 154.255 66.965 155.395 ;
        RECT 67.135 154.425 67.470 155.395 ;
        RECT 68.565 155.825 69.795 155.995 ;
        RECT 68.565 155.015 68.905 155.825 ;
        RECT 69.075 155.260 69.825 155.450 ;
        RECT 68.565 154.605 69.080 155.015 ;
        RECT 69.315 154.255 69.485 155.015 ;
        RECT 69.655 154.595 69.825 155.260 ;
        RECT 69.995 155.275 70.185 156.635 ;
        RECT 70.355 156.125 70.630 156.635 ;
        RECT 70.820 156.270 71.350 156.635 ;
        RECT 71.775 156.405 72.105 156.805 ;
        RECT 71.175 156.235 71.350 156.270 ;
        RECT 70.355 155.955 70.635 156.125 ;
        RECT 70.355 155.475 70.630 155.955 ;
        RECT 70.835 155.275 71.005 156.075 ;
        RECT 69.995 155.105 71.005 155.275 ;
        RECT 71.175 156.065 72.105 156.235 ;
        RECT 72.275 156.065 72.530 156.635 ;
        RECT 71.175 154.935 71.345 156.065 ;
        RECT 71.935 155.895 72.105 156.065 ;
        RECT 70.220 154.765 71.345 154.935 ;
        RECT 71.515 155.565 71.710 155.895 ;
        RECT 71.935 155.565 72.190 155.895 ;
        RECT 71.515 154.595 71.685 155.565 ;
        RECT 72.360 155.395 72.530 156.065 ;
        RECT 72.765 155.985 72.975 156.805 ;
        RECT 73.145 156.005 73.475 156.635 ;
        RECT 73.145 155.405 73.395 156.005 ;
        RECT 73.645 155.985 73.875 156.805 ;
        RECT 75.065 156.325 75.345 156.805 ;
        RECT 75.515 156.155 75.775 156.545 ;
        RECT 75.950 156.325 76.205 156.805 ;
        RECT 76.375 156.155 76.670 156.545 ;
        RECT 76.850 156.325 77.125 156.805 ;
        RECT 77.295 156.305 77.595 156.635 ;
        RECT 75.020 155.985 76.670 156.155 ;
        RECT 73.565 155.565 73.895 155.815 ;
        RECT 75.020 155.475 75.425 155.985 ;
        RECT 75.595 155.645 76.735 155.815 ;
        RECT 69.655 154.425 71.685 154.595 ;
        RECT 71.855 154.255 72.025 155.395 ;
        RECT 72.195 154.425 72.530 155.395 ;
        RECT 72.765 154.255 72.975 155.395 ;
        RECT 73.145 154.425 73.475 155.405 ;
        RECT 73.645 154.255 73.875 155.395 ;
        RECT 75.020 155.305 75.775 155.475 ;
        RECT 75.060 154.255 75.345 155.125 ;
        RECT 75.515 155.055 75.775 155.305 ;
        RECT 76.565 155.395 76.735 155.645 ;
        RECT 76.905 155.565 77.255 156.135 ;
        RECT 77.425 155.395 77.595 156.305 ;
        RECT 76.565 155.225 77.595 155.395 ;
        RECT 75.515 154.885 76.635 155.055 ;
        RECT 75.515 154.425 75.775 154.885 ;
        RECT 75.950 154.255 76.205 154.715 ;
        RECT 76.375 154.425 76.635 154.885 ;
        RECT 76.805 154.255 77.115 155.055 ;
        RECT 77.285 154.425 77.595 155.225 ;
        RECT 78.225 156.305 78.525 156.635 ;
        RECT 78.695 156.325 78.970 156.805 ;
        RECT 78.225 155.395 78.395 156.305 ;
        RECT 79.150 156.155 79.445 156.545 ;
        RECT 79.615 156.325 79.870 156.805 ;
        RECT 80.045 156.155 80.305 156.545 ;
        RECT 80.475 156.325 80.755 156.805 ;
        RECT 78.565 155.565 78.915 156.135 ;
        RECT 79.150 155.985 80.800 156.155 ;
        RECT 81.190 156.025 81.690 156.635 ;
        RECT 79.085 155.645 80.225 155.815 ;
        RECT 79.085 155.395 79.255 155.645 ;
        RECT 80.395 155.475 80.800 155.985 ;
        RECT 80.985 155.565 81.335 155.815 ;
        RECT 78.225 155.225 79.255 155.395 ;
        RECT 80.045 155.305 80.800 155.475 ;
        RECT 81.520 155.395 81.690 156.025 ;
        RECT 82.320 156.155 82.650 156.635 ;
        RECT 82.820 156.345 83.045 156.805 ;
        RECT 83.215 156.155 83.545 156.635 ;
        RECT 82.320 155.985 83.545 156.155 ;
        RECT 83.735 156.005 83.985 156.805 ;
        RECT 84.155 156.005 84.495 156.635 ;
        RECT 81.860 155.615 82.190 155.815 ;
        RECT 82.360 155.615 82.690 155.815 ;
        RECT 82.860 155.615 83.280 155.815 ;
        RECT 83.455 155.645 84.150 155.815 ;
        RECT 83.455 155.395 83.625 155.645 ;
        RECT 84.320 155.395 84.495 156.005 ;
        RECT 84.940 155.995 85.185 156.600 ;
        RECT 85.405 156.270 85.915 156.805 ;
        RECT 78.225 154.425 78.535 155.225 ;
        RECT 80.045 155.055 80.305 155.305 ;
        RECT 81.190 155.225 83.625 155.395 ;
        RECT 78.705 154.255 79.015 155.055 ;
        RECT 79.185 154.885 80.305 155.055 ;
        RECT 79.185 154.425 79.445 154.885 ;
        RECT 79.615 154.255 79.870 154.715 ;
        RECT 80.045 154.425 80.305 154.885 ;
        RECT 80.475 154.255 80.760 155.125 ;
        RECT 81.190 154.425 81.520 155.225 ;
        RECT 81.690 154.255 82.020 155.055 ;
        RECT 82.320 154.425 82.650 155.225 ;
        RECT 83.295 154.255 83.545 155.055 ;
        RECT 83.815 154.255 83.985 155.395 ;
        RECT 84.155 154.425 84.495 155.395 ;
        RECT 84.665 155.825 85.895 155.995 ;
        RECT 84.665 155.015 85.005 155.825 ;
        RECT 85.175 155.260 85.925 155.450 ;
        RECT 84.665 154.605 85.180 155.015 ;
        RECT 85.415 154.255 85.585 155.015 ;
        RECT 85.755 154.595 85.925 155.260 ;
        RECT 86.095 155.275 86.285 156.635 ;
        RECT 86.455 155.785 86.730 156.635 ;
        RECT 86.920 156.270 87.450 156.635 ;
        RECT 87.875 156.405 88.205 156.805 ;
        RECT 87.275 156.235 87.450 156.270 ;
        RECT 86.455 155.615 86.735 155.785 ;
        RECT 86.455 155.475 86.730 155.615 ;
        RECT 86.935 155.275 87.105 156.075 ;
        RECT 86.095 155.105 87.105 155.275 ;
        RECT 87.275 156.065 88.205 156.235 ;
        RECT 88.375 156.065 88.630 156.635 ;
        RECT 88.805 156.080 89.095 156.805 ;
        RECT 87.275 154.935 87.445 156.065 ;
        RECT 88.035 155.895 88.205 156.065 ;
        RECT 86.320 154.765 87.445 154.935 ;
        RECT 87.615 155.565 87.810 155.895 ;
        RECT 88.035 155.565 88.290 155.895 ;
        RECT 87.615 154.595 87.785 155.565 ;
        RECT 88.460 155.395 88.630 156.065 ;
        RECT 89.265 156.055 90.475 156.805 ;
        RECT 85.755 154.425 87.785 154.595 ;
        RECT 87.955 154.255 88.125 155.395 ;
        RECT 88.295 154.425 88.630 155.395 ;
        RECT 88.805 154.255 89.095 155.420 ;
        RECT 89.265 155.345 89.785 155.885 ;
        RECT 89.955 155.515 90.475 156.055 ;
        RECT 90.705 155.985 90.915 156.805 ;
        RECT 91.085 156.005 91.415 156.635 ;
        RECT 91.085 155.405 91.335 156.005 ;
        RECT 91.585 155.985 91.815 156.805 ;
        RECT 92.575 156.255 92.745 156.635 ;
        RECT 92.925 156.425 93.255 156.805 ;
        RECT 92.575 156.085 93.240 156.255 ;
        RECT 93.435 156.130 93.695 156.635 ;
        RECT 91.505 155.565 91.835 155.815 ;
        RECT 92.505 155.535 92.835 155.905 ;
        RECT 93.070 155.830 93.240 156.085 ;
        RECT 93.070 155.500 93.355 155.830 ;
        RECT 89.265 154.255 90.475 155.345 ;
        RECT 90.705 154.255 90.915 155.395 ;
        RECT 91.085 154.425 91.415 155.405 ;
        RECT 91.585 154.255 91.815 155.395 ;
        RECT 93.070 155.355 93.240 155.500 ;
        RECT 92.575 155.185 93.240 155.355 ;
        RECT 93.525 155.330 93.695 156.130 ;
        RECT 93.980 156.175 94.265 156.635 ;
        RECT 94.435 156.345 94.705 156.805 ;
        RECT 93.980 156.005 94.935 156.175 ;
        RECT 92.575 154.425 92.745 155.185 ;
        RECT 92.925 154.255 93.255 155.015 ;
        RECT 93.425 154.425 93.695 155.330 ;
        RECT 93.865 155.275 94.555 155.835 ;
        RECT 94.725 155.105 94.935 156.005 ;
        RECT 93.980 154.885 94.935 155.105 ;
        RECT 95.105 155.835 95.505 156.635 ;
        RECT 95.695 156.175 95.975 156.635 ;
        RECT 96.495 156.345 96.820 156.805 ;
        RECT 95.695 156.005 96.820 156.175 ;
        RECT 96.990 156.065 97.375 156.635 ;
        RECT 96.370 155.895 96.820 156.005 ;
        RECT 95.105 155.275 96.200 155.835 ;
        RECT 96.370 155.565 96.925 155.895 ;
        RECT 93.980 154.425 94.265 154.885 ;
        RECT 94.435 154.255 94.705 154.715 ;
        RECT 95.105 154.425 95.505 155.275 ;
        RECT 96.370 155.105 96.820 155.565 ;
        RECT 97.095 155.395 97.375 156.065 ;
        RECT 97.820 155.995 98.065 156.600 ;
        RECT 98.285 156.270 98.795 156.805 ;
        RECT 95.695 154.885 96.820 155.105 ;
        RECT 95.695 154.425 95.975 154.885 ;
        RECT 96.495 154.255 96.820 154.715 ;
        RECT 96.990 154.425 97.375 155.395 ;
        RECT 97.545 155.825 98.775 155.995 ;
        RECT 97.545 155.015 97.885 155.825 ;
        RECT 98.055 155.260 98.805 155.450 ;
        RECT 97.545 154.605 98.060 155.015 ;
        RECT 98.295 154.255 98.465 155.015 ;
        RECT 98.635 154.595 98.805 155.260 ;
        RECT 98.975 155.275 99.165 156.635 ;
        RECT 99.335 156.125 99.610 156.635 ;
        RECT 99.800 156.270 100.330 156.635 ;
        RECT 100.755 156.405 101.085 156.805 ;
        RECT 100.155 156.235 100.330 156.270 ;
        RECT 99.335 155.955 99.615 156.125 ;
        RECT 99.335 155.475 99.610 155.955 ;
        RECT 99.815 155.275 99.985 156.075 ;
        RECT 98.975 155.105 99.985 155.275 ;
        RECT 100.155 156.065 101.085 156.235 ;
        RECT 101.255 156.065 101.510 156.635 ;
        RECT 101.775 156.255 101.945 156.635 ;
        RECT 102.125 156.425 102.455 156.805 ;
        RECT 101.775 156.085 102.440 156.255 ;
        RECT 102.635 156.130 102.895 156.635 ;
        RECT 100.155 154.935 100.325 156.065 ;
        RECT 100.915 155.895 101.085 156.065 ;
        RECT 99.200 154.765 100.325 154.935 ;
        RECT 100.495 155.565 100.690 155.895 ;
        RECT 100.915 155.565 101.170 155.895 ;
        RECT 100.495 154.595 100.665 155.565 ;
        RECT 101.340 155.395 101.510 156.065 ;
        RECT 101.705 155.535 102.035 155.905 ;
        RECT 102.270 155.830 102.440 156.085 ;
        RECT 98.635 154.425 100.665 154.595 ;
        RECT 100.835 154.255 101.005 155.395 ;
        RECT 101.175 154.425 101.510 155.395 ;
        RECT 102.270 155.500 102.555 155.830 ;
        RECT 102.270 155.355 102.440 155.500 ;
        RECT 101.775 155.185 102.440 155.355 ;
        RECT 102.725 155.330 102.895 156.130 ;
        RECT 103.065 156.055 104.275 156.805 ;
        RECT 101.775 154.425 101.945 155.185 ;
        RECT 102.125 154.255 102.455 155.015 ;
        RECT 102.625 154.425 102.895 155.330 ;
        RECT 103.065 155.345 103.585 155.885 ;
        RECT 103.755 155.515 104.275 156.055 ;
        RECT 104.445 156.035 107.955 156.805 ;
        RECT 108.135 156.305 108.465 156.805 ;
        RECT 108.665 156.235 108.835 156.585 ;
        RECT 109.035 156.405 109.365 156.805 ;
        RECT 109.535 156.235 109.705 156.585 ;
        RECT 109.875 156.405 110.255 156.805 ;
        RECT 104.445 155.345 106.135 155.865 ;
        RECT 106.305 155.515 107.955 156.035 ;
        RECT 108.130 155.565 108.480 156.135 ;
        RECT 108.665 156.065 110.275 156.235 ;
        RECT 110.445 156.130 110.715 156.475 ;
        RECT 110.105 155.895 110.275 156.065 ;
        RECT 103.065 154.255 104.275 155.345 ;
        RECT 104.445 154.255 107.955 155.345 ;
        RECT 108.130 155.105 108.450 155.395 ;
        RECT 108.650 155.275 109.360 155.895 ;
        RECT 109.530 155.565 109.935 155.895 ;
        RECT 110.105 155.565 110.375 155.895 ;
        RECT 110.105 155.395 110.275 155.565 ;
        RECT 110.545 155.395 110.715 156.130 ;
        RECT 111.000 156.175 111.285 156.635 ;
        RECT 111.455 156.345 111.725 156.805 ;
        RECT 111.000 156.005 111.955 156.175 ;
        RECT 109.550 155.225 110.275 155.395 ;
        RECT 109.550 155.105 109.720 155.225 ;
        RECT 108.130 154.935 109.720 155.105 ;
        RECT 108.130 154.475 109.785 154.765 ;
        RECT 109.955 154.255 110.235 155.055 ;
        RECT 110.445 154.425 110.715 155.395 ;
        RECT 110.885 155.275 111.575 155.835 ;
        RECT 111.745 155.105 111.955 156.005 ;
        RECT 111.000 154.885 111.955 155.105 ;
        RECT 112.125 155.835 112.525 156.635 ;
        RECT 112.715 156.175 112.995 156.635 ;
        RECT 113.515 156.345 113.840 156.805 ;
        RECT 112.715 156.005 113.840 156.175 ;
        RECT 114.010 156.065 114.395 156.635 ;
        RECT 114.565 156.080 114.855 156.805 ;
        RECT 113.390 155.895 113.840 156.005 ;
        RECT 112.125 155.275 113.220 155.835 ;
        RECT 113.390 155.565 113.945 155.895 ;
        RECT 111.000 154.425 111.285 154.885 ;
        RECT 111.455 154.255 111.725 154.715 ;
        RECT 112.125 154.425 112.525 155.275 ;
        RECT 113.390 155.105 113.840 155.565 ;
        RECT 114.115 155.395 114.395 156.065 ;
        RECT 115.525 155.985 115.755 156.805 ;
        RECT 115.925 156.005 116.255 156.635 ;
        RECT 115.505 155.565 115.835 155.815 ;
        RECT 112.715 154.885 113.840 155.105 ;
        RECT 112.715 154.425 112.995 154.885 ;
        RECT 113.515 154.255 113.840 154.715 ;
        RECT 114.010 154.425 114.395 155.395 ;
        RECT 114.565 154.255 114.855 155.420 ;
        RECT 116.005 155.405 116.255 156.005 ;
        RECT 116.425 155.985 116.635 156.805 ;
        RECT 117.240 156.095 117.495 156.625 ;
        RECT 117.675 156.345 117.960 156.805 ;
        RECT 115.525 154.255 115.755 155.395 ;
        RECT 115.925 154.425 116.255 155.405 ;
        RECT 116.425 154.255 116.635 155.395 ;
        RECT 117.240 155.235 117.420 156.095 ;
        RECT 118.140 155.895 118.390 156.545 ;
        RECT 117.590 155.565 118.390 155.895 ;
        RECT 117.240 155.105 117.495 155.235 ;
        RECT 117.155 154.935 117.495 155.105 ;
        RECT 117.240 154.565 117.495 154.935 ;
        RECT 117.675 154.255 117.960 155.055 ;
        RECT 118.140 154.975 118.390 155.565 ;
        RECT 118.590 156.210 118.910 156.540 ;
        RECT 119.090 156.325 119.750 156.805 ;
        RECT 119.950 156.415 120.800 156.585 ;
        RECT 118.590 155.315 118.780 156.210 ;
        RECT 119.100 155.885 119.760 156.155 ;
        RECT 119.430 155.825 119.760 155.885 ;
        RECT 118.950 155.655 119.280 155.715 ;
        RECT 119.950 155.655 120.120 156.415 ;
        RECT 121.360 156.345 121.680 156.805 ;
        RECT 121.880 156.165 122.130 156.595 ;
        RECT 122.420 156.365 122.830 156.805 ;
        RECT 123.000 156.425 124.015 156.625 ;
        RECT 120.290 155.995 121.540 156.165 ;
        RECT 120.290 155.875 120.620 155.995 ;
        RECT 118.950 155.485 120.850 155.655 ;
        RECT 118.590 155.145 120.510 155.315 ;
        RECT 118.590 155.125 118.910 155.145 ;
        RECT 118.140 154.465 118.470 154.975 ;
        RECT 118.740 154.515 118.910 155.125 ;
        RECT 120.680 154.975 120.850 155.485 ;
        RECT 121.020 155.415 121.200 155.825 ;
        RECT 121.370 155.235 121.540 155.995 ;
        RECT 119.080 154.255 119.410 154.945 ;
        RECT 119.640 154.805 120.850 154.975 ;
        RECT 121.020 154.925 121.540 155.235 ;
        RECT 121.710 155.825 122.130 156.165 ;
        RECT 122.420 155.825 122.830 156.155 ;
        RECT 121.710 155.055 121.900 155.825 ;
        RECT 123.000 155.695 123.170 156.425 ;
        RECT 124.315 156.255 124.485 156.585 ;
        RECT 124.655 156.425 124.985 156.805 ;
        RECT 123.340 155.875 123.690 156.245 ;
        RECT 123.000 155.655 123.420 155.695 ;
        RECT 122.070 155.485 123.420 155.655 ;
        RECT 122.070 155.325 122.320 155.485 ;
        RECT 122.830 155.055 123.080 155.315 ;
        RECT 121.710 154.805 123.080 155.055 ;
        RECT 119.640 154.515 119.880 154.805 ;
        RECT 120.680 154.725 120.850 154.805 ;
        RECT 120.080 154.255 120.500 154.635 ;
        RECT 120.680 154.475 121.310 154.725 ;
        RECT 121.780 154.255 122.110 154.635 ;
        RECT 122.280 154.515 122.450 154.805 ;
        RECT 123.250 154.640 123.420 155.485 ;
        RECT 123.870 155.315 124.090 156.185 ;
        RECT 124.315 156.065 125.010 156.255 ;
        RECT 123.590 154.935 124.090 155.315 ;
        RECT 124.260 155.265 124.670 155.885 ;
        RECT 124.840 155.095 125.010 156.065 ;
        RECT 124.315 154.925 125.010 155.095 ;
        RECT 122.630 154.255 123.010 154.635 ;
        RECT 123.250 154.470 124.080 154.640 ;
        RECT 124.315 154.425 124.485 154.925 ;
        RECT 124.655 154.255 124.985 154.755 ;
        RECT 125.200 154.425 125.425 156.545 ;
        RECT 125.595 156.425 125.925 156.805 ;
        RECT 126.095 156.255 126.265 156.545 ;
        RECT 125.600 156.085 126.265 156.255 ;
        RECT 125.600 155.095 125.830 156.085 ;
        RECT 126.525 156.055 127.735 156.805 ;
        RECT 126.000 155.265 126.350 155.915 ;
        RECT 126.525 155.345 127.045 155.885 ;
        RECT 127.215 155.515 127.735 156.055 ;
        RECT 125.600 154.925 126.265 155.095 ;
        RECT 125.595 154.255 125.925 154.755 ;
        RECT 126.095 154.425 126.265 154.925 ;
        RECT 126.525 154.255 127.735 155.345 ;
        RECT 29.840 154.085 127.820 154.255 ;
        RECT 29.925 152.995 31.135 154.085 ;
        RECT 29.925 152.285 30.445 152.825 ;
        RECT 30.615 152.455 31.135 152.995 ;
        RECT 31.680 153.105 31.935 153.775 ;
        RECT 32.115 153.285 32.400 154.085 ;
        RECT 32.580 153.365 32.910 153.875 ;
        RECT 29.925 151.535 31.135 152.285 ;
        RECT 31.680 152.245 31.860 153.105 ;
        RECT 32.580 152.775 32.830 153.365 ;
        RECT 33.180 153.215 33.350 153.825 ;
        RECT 33.520 153.395 33.850 154.085 ;
        RECT 34.080 153.535 34.320 153.825 ;
        RECT 34.520 153.705 34.940 154.085 ;
        RECT 35.120 153.615 35.750 153.865 ;
        RECT 36.220 153.705 36.550 154.085 ;
        RECT 35.120 153.535 35.290 153.615 ;
        RECT 36.720 153.535 36.890 153.825 ;
        RECT 37.070 153.705 37.450 154.085 ;
        RECT 37.690 153.700 38.520 153.870 ;
        RECT 34.080 153.365 35.290 153.535 ;
        RECT 32.030 152.445 32.830 152.775 ;
        RECT 31.680 152.045 31.935 152.245 ;
        RECT 31.595 151.875 31.935 152.045 ;
        RECT 31.680 151.715 31.935 151.875 ;
        RECT 32.115 151.535 32.400 151.995 ;
        RECT 32.580 151.795 32.830 152.445 ;
        RECT 33.030 153.195 33.350 153.215 ;
        RECT 33.030 153.025 34.950 153.195 ;
        RECT 33.030 152.130 33.220 153.025 ;
        RECT 35.120 152.855 35.290 153.365 ;
        RECT 35.460 153.105 35.980 153.415 ;
        RECT 33.390 152.685 35.290 152.855 ;
        RECT 33.390 152.625 33.720 152.685 ;
        RECT 33.870 152.455 34.200 152.515 ;
        RECT 33.540 152.185 34.200 152.455 ;
        RECT 33.030 151.800 33.350 152.130 ;
        RECT 33.530 151.535 34.190 152.015 ;
        RECT 34.390 151.925 34.560 152.685 ;
        RECT 35.460 152.515 35.640 152.925 ;
        RECT 34.730 152.345 35.060 152.465 ;
        RECT 35.810 152.345 35.980 153.105 ;
        RECT 34.730 152.175 35.980 152.345 ;
        RECT 36.150 153.285 37.520 153.535 ;
        RECT 36.150 152.515 36.340 153.285 ;
        RECT 37.270 153.025 37.520 153.285 ;
        RECT 36.510 152.855 36.760 153.015 ;
        RECT 37.690 152.855 37.860 153.700 ;
        RECT 38.755 153.415 38.925 153.915 ;
        RECT 39.095 153.585 39.425 154.085 ;
        RECT 38.030 153.025 38.530 153.405 ;
        RECT 38.755 153.245 39.450 153.415 ;
        RECT 36.510 152.685 37.860 152.855 ;
        RECT 37.440 152.645 37.860 152.685 ;
        RECT 36.150 152.175 36.570 152.515 ;
        RECT 36.860 152.185 37.270 152.515 ;
        RECT 34.390 151.755 35.240 151.925 ;
        RECT 35.800 151.535 36.120 151.995 ;
        RECT 36.320 151.745 36.570 152.175 ;
        RECT 36.860 151.535 37.270 151.975 ;
        RECT 37.440 151.915 37.610 152.645 ;
        RECT 37.780 152.095 38.130 152.465 ;
        RECT 38.310 152.155 38.530 153.025 ;
        RECT 38.700 152.455 39.110 153.075 ;
        RECT 39.280 152.275 39.450 153.245 ;
        RECT 38.755 152.085 39.450 152.275 ;
        RECT 37.440 151.715 38.455 151.915 ;
        RECT 38.755 151.755 38.925 152.085 ;
        RECT 39.095 151.535 39.425 151.915 ;
        RECT 39.640 151.795 39.865 153.915 ;
        RECT 40.035 153.585 40.365 154.085 ;
        RECT 40.535 153.415 40.705 153.915 ;
        RECT 40.040 153.245 40.705 153.415 ;
        RECT 40.040 152.255 40.270 153.245 ;
        RECT 40.440 152.425 40.790 153.075 ;
        RECT 41.425 152.995 43.095 154.085 ;
        RECT 43.355 153.155 43.525 153.915 ;
        RECT 43.705 153.325 44.035 154.085 ;
        RECT 41.425 152.475 42.175 152.995 ;
        RECT 43.355 152.985 44.020 153.155 ;
        RECT 44.205 153.010 44.475 153.915 ;
        RECT 43.850 152.840 44.020 152.985 ;
        RECT 42.345 152.305 43.095 152.825 ;
        RECT 43.285 152.435 43.615 152.805 ;
        RECT 43.850 152.510 44.135 152.840 ;
        RECT 40.040 152.085 40.705 152.255 ;
        RECT 40.035 151.535 40.365 151.915 ;
        RECT 40.535 151.795 40.705 152.085 ;
        RECT 41.425 151.535 43.095 152.305 ;
        RECT 43.850 152.255 44.020 152.510 ;
        RECT 43.355 152.085 44.020 152.255 ;
        RECT 44.305 152.210 44.475 153.010 ;
        RECT 43.355 151.705 43.525 152.085 ;
        RECT 43.705 151.535 44.035 151.915 ;
        RECT 44.215 151.705 44.475 152.210 ;
        RECT 44.645 152.945 44.915 153.915 ;
        RECT 45.125 153.285 45.405 154.085 ;
        RECT 45.575 153.575 47.230 153.865 ;
        RECT 47.410 153.575 49.065 153.865 ;
        RECT 45.640 153.235 47.230 153.405 ;
        RECT 45.640 153.115 45.810 153.235 ;
        RECT 45.085 152.945 45.810 153.115 ;
        RECT 44.645 152.210 44.815 152.945 ;
        RECT 45.085 152.775 45.255 152.945 ;
        RECT 44.985 152.445 45.255 152.775 ;
        RECT 45.425 152.445 45.830 152.775 ;
        RECT 46.000 152.445 46.710 153.065 ;
        RECT 46.910 152.945 47.230 153.235 ;
        RECT 47.410 153.235 49.000 153.405 ;
        RECT 49.235 153.285 49.515 154.085 ;
        RECT 47.410 152.945 47.730 153.235 ;
        RECT 48.830 153.115 49.000 153.235 ;
        RECT 45.085 152.275 45.255 152.445 ;
        RECT 44.645 151.865 44.915 152.210 ;
        RECT 45.085 152.105 46.695 152.275 ;
        RECT 46.880 152.205 47.230 152.775 ;
        RECT 47.410 152.205 47.760 152.775 ;
        RECT 47.930 152.445 48.640 153.065 ;
        RECT 48.830 152.945 49.555 153.115 ;
        RECT 49.725 152.945 49.995 153.915 ;
        RECT 49.385 152.775 49.555 152.945 ;
        RECT 48.810 152.445 49.215 152.775 ;
        RECT 49.385 152.445 49.655 152.775 ;
        RECT 49.385 152.275 49.555 152.445 ;
        RECT 45.105 151.535 45.485 151.935 ;
        RECT 45.655 151.755 45.825 152.105 ;
        RECT 45.995 151.535 46.325 151.935 ;
        RECT 46.525 151.755 46.695 152.105 ;
        RECT 47.945 152.105 49.555 152.275 ;
        RECT 49.825 152.210 49.995 152.945 ;
        RECT 50.165 152.920 50.455 154.085 ;
        RECT 50.825 153.415 51.105 154.085 ;
        RECT 51.275 153.195 51.575 153.745 ;
        RECT 51.775 153.365 52.105 154.085 ;
        RECT 52.295 153.365 52.755 153.915 ;
        RECT 50.640 152.775 50.905 153.135 ;
        RECT 51.275 153.025 52.215 153.195 ;
        RECT 52.045 152.775 52.215 153.025 ;
        RECT 50.640 152.525 51.315 152.775 ;
        RECT 51.535 152.525 51.875 152.775 ;
        RECT 52.045 152.445 52.335 152.775 ;
        RECT 52.045 152.355 52.215 152.445 ;
        RECT 46.895 151.535 47.225 152.035 ;
        RECT 47.415 151.535 47.745 152.035 ;
        RECT 47.945 151.755 48.115 152.105 ;
        RECT 48.315 151.535 48.645 151.935 ;
        RECT 48.815 151.755 48.985 152.105 ;
        RECT 49.155 151.535 49.535 151.935 ;
        RECT 49.725 151.865 49.995 152.210 ;
        RECT 50.165 151.535 50.455 152.260 ;
        RECT 50.825 152.165 52.215 152.355 ;
        RECT 50.825 151.805 51.155 152.165 ;
        RECT 52.505 151.995 52.755 153.365 ;
        RECT 51.775 151.535 52.025 151.995 ;
        RECT 52.195 151.705 52.755 151.995 ;
        RECT 52.925 152.945 53.265 153.915 ;
        RECT 53.435 152.945 53.605 154.085 ;
        RECT 53.875 153.285 54.125 154.085 ;
        RECT 54.770 153.115 55.100 153.915 ;
        RECT 55.400 153.285 55.730 154.085 ;
        RECT 55.900 153.115 56.230 153.915 ;
        RECT 56.980 153.745 57.235 153.775 ;
        RECT 56.895 153.575 57.235 153.745 ;
        RECT 53.795 152.945 56.230 153.115 ;
        RECT 56.980 153.105 57.235 153.575 ;
        RECT 57.415 153.285 57.700 154.085 ;
        RECT 57.880 153.365 58.210 153.875 ;
        RECT 52.925 152.895 53.155 152.945 ;
        RECT 52.925 152.335 53.100 152.895 ;
        RECT 53.795 152.695 53.965 152.945 ;
        RECT 53.270 152.525 53.965 152.695 ;
        RECT 54.140 152.525 54.560 152.725 ;
        RECT 54.730 152.525 55.060 152.725 ;
        RECT 55.230 152.525 55.560 152.725 ;
        RECT 52.925 151.705 53.265 152.335 ;
        RECT 53.435 151.535 53.685 152.335 ;
        RECT 53.875 152.185 55.100 152.355 ;
        RECT 53.875 151.705 54.205 152.185 ;
        RECT 54.375 151.535 54.600 151.995 ;
        RECT 54.770 151.705 55.100 152.185 ;
        RECT 55.730 152.315 55.900 152.945 ;
        RECT 56.085 152.525 56.435 152.775 ;
        RECT 55.730 151.705 56.230 152.315 ;
        RECT 56.980 152.245 57.160 153.105 ;
        RECT 57.880 152.775 58.130 153.365 ;
        RECT 58.480 153.215 58.650 153.825 ;
        RECT 58.820 153.395 59.150 154.085 ;
        RECT 59.380 153.535 59.620 153.825 ;
        RECT 59.820 153.705 60.240 154.085 ;
        RECT 60.420 153.615 61.050 153.865 ;
        RECT 61.520 153.705 61.850 154.085 ;
        RECT 60.420 153.535 60.590 153.615 ;
        RECT 62.020 153.535 62.190 153.825 ;
        RECT 62.370 153.705 62.750 154.085 ;
        RECT 62.990 153.700 63.820 153.870 ;
        RECT 59.380 153.365 60.590 153.535 ;
        RECT 57.330 152.445 58.130 152.775 ;
        RECT 56.980 151.715 57.235 152.245 ;
        RECT 57.415 151.535 57.700 151.995 ;
        RECT 57.880 151.795 58.130 152.445 ;
        RECT 58.330 153.195 58.650 153.215 ;
        RECT 58.330 153.025 60.250 153.195 ;
        RECT 58.330 152.130 58.520 153.025 ;
        RECT 60.420 152.855 60.590 153.365 ;
        RECT 60.760 153.105 61.280 153.415 ;
        RECT 58.690 152.685 60.590 152.855 ;
        RECT 58.690 152.625 59.020 152.685 ;
        RECT 59.170 152.455 59.500 152.515 ;
        RECT 58.840 152.185 59.500 152.455 ;
        RECT 58.330 151.800 58.650 152.130 ;
        RECT 58.830 151.535 59.490 152.015 ;
        RECT 59.690 151.925 59.860 152.685 ;
        RECT 60.760 152.515 60.940 152.925 ;
        RECT 60.030 152.345 60.360 152.465 ;
        RECT 61.110 152.345 61.280 153.105 ;
        RECT 60.030 152.175 61.280 152.345 ;
        RECT 61.450 153.285 62.820 153.535 ;
        RECT 61.450 152.515 61.640 153.285 ;
        RECT 62.570 153.025 62.820 153.285 ;
        RECT 61.810 152.855 62.060 153.015 ;
        RECT 62.990 152.855 63.160 153.700 ;
        RECT 64.055 153.415 64.225 153.915 ;
        RECT 64.395 153.585 64.725 154.085 ;
        RECT 63.330 153.025 63.830 153.405 ;
        RECT 64.055 153.245 64.750 153.415 ;
        RECT 61.810 152.685 63.160 152.855 ;
        RECT 62.740 152.645 63.160 152.685 ;
        RECT 61.450 152.175 61.870 152.515 ;
        RECT 62.160 152.185 62.570 152.515 ;
        RECT 59.690 151.755 60.540 151.925 ;
        RECT 61.100 151.535 61.420 151.995 ;
        RECT 61.620 151.745 61.870 152.175 ;
        RECT 62.160 151.535 62.570 151.975 ;
        RECT 62.740 151.915 62.910 152.645 ;
        RECT 63.080 152.095 63.430 152.465 ;
        RECT 63.610 152.155 63.830 153.025 ;
        RECT 64.000 152.455 64.410 153.075 ;
        RECT 64.580 152.275 64.750 153.245 ;
        RECT 64.055 152.085 64.750 152.275 ;
        RECT 62.740 151.715 63.755 151.915 ;
        RECT 64.055 151.755 64.225 152.085 ;
        RECT 64.395 151.535 64.725 151.915 ;
        RECT 64.940 151.795 65.165 153.915 ;
        RECT 65.335 153.585 65.665 154.085 ;
        RECT 65.835 153.415 66.005 153.915 ;
        RECT 65.340 153.245 66.005 153.415 ;
        RECT 65.340 152.255 65.570 153.245 ;
        RECT 65.740 152.425 66.090 153.075 ;
        RECT 66.730 152.895 66.985 153.775 ;
        RECT 67.155 152.945 67.460 154.085 ;
        RECT 67.800 153.705 68.130 154.085 ;
        RECT 68.310 153.535 68.480 153.825 ;
        RECT 68.650 153.625 68.900 154.085 ;
        RECT 67.680 153.365 68.480 153.535 ;
        RECT 69.070 153.575 69.940 153.915 ;
        RECT 65.340 152.085 66.005 152.255 ;
        RECT 65.335 151.535 65.665 151.915 ;
        RECT 65.835 151.795 66.005 152.085 ;
        RECT 66.730 152.245 66.940 152.895 ;
        RECT 67.680 152.775 67.850 153.365 ;
        RECT 69.070 153.195 69.240 153.575 ;
        RECT 70.175 153.455 70.345 153.915 ;
        RECT 70.515 153.625 70.885 154.085 ;
        RECT 71.180 153.485 71.350 153.825 ;
        RECT 71.520 153.655 71.850 154.085 ;
        RECT 72.085 153.485 72.255 153.825 ;
        RECT 68.020 153.025 69.240 153.195 ;
        RECT 69.410 153.115 69.870 153.405 ;
        RECT 70.175 153.285 70.735 153.455 ;
        RECT 71.180 153.315 72.255 153.485 ;
        RECT 72.425 153.585 73.105 153.915 ;
        RECT 73.320 153.585 73.570 153.915 ;
        RECT 73.740 153.625 73.990 154.085 ;
        RECT 70.565 153.145 70.735 153.285 ;
        RECT 69.410 153.105 70.375 153.115 ;
        RECT 69.070 152.935 69.240 153.025 ;
        RECT 69.700 152.945 70.375 153.105 ;
        RECT 67.110 152.745 67.850 152.775 ;
        RECT 67.110 152.445 68.025 152.745 ;
        RECT 67.700 152.270 68.025 152.445 ;
        RECT 66.730 151.715 66.985 152.245 ;
        RECT 67.155 151.535 67.460 151.995 ;
        RECT 67.705 151.915 68.025 152.270 ;
        RECT 68.195 152.485 68.735 152.855 ;
        RECT 69.070 152.765 69.475 152.935 ;
        RECT 68.195 152.085 68.435 152.485 ;
        RECT 68.915 152.315 69.135 152.595 ;
        RECT 68.605 152.145 69.135 152.315 ;
        RECT 68.605 151.915 68.775 152.145 ;
        RECT 69.305 151.985 69.475 152.765 ;
        RECT 69.645 152.155 69.995 152.775 ;
        RECT 70.165 152.155 70.375 152.945 ;
        RECT 70.565 152.975 72.065 153.145 ;
        RECT 70.565 152.285 70.735 152.975 ;
        RECT 72.425 152.805 72.595 153.585 ;
        RECT 73.400 153.455 73.570 153.585 ;
        RECT 70.905 152.635 72.595 152.805 ;
        RECT 72.765 153.025 73.230 153.415 ;
        RECT 73.400 153.285 73.795 153.455 ;
        RECT 70.905 152.455 71.075 152.635 ;
        RECT 67.705 151.745 68.775 151.915 ;
        RECT 68.945 151.535 69.135 151.975 ;
        RECT 69.305 151.705 70.255 151.985 ;
        RECT 70.565 151.895 70.825 152.285 ;
        RECT 71.245 152.215 72.035 152.465 ;
        RECT 70.475 151.725 70.825 151.895 ;
        RECT 71.035 151.535 71.365 151.995 ;
        RECT 72.240 151.925 72.410 152.635 ;
        RECT 72.765 152.435 72.935 153.025 ;
        RECT 72.580 152.215 72.935 152.435 ;
        RECT 73.105 152.215 73.455 152.835 ;
        RECT 73.625 151.925 73.795 153.285 ;
        RECT 74.160 153.115 74.485 153.900 ;
        RECT 73.965 152.065 74.425 153.115 ;
        RECT 72.240 151.755 73.095 151.925 ;
        RECT 73.300 151.755 73.795 151.925 ;
        RECT 73.965 151.535 74.295 151.895 ;
        RECT 74.655 151.795 74.825 153.915 ;
        RECT 74.995 153.585 75.325 154.085 ;
        RECT 75.495 153.415 75.750 153.915 ;
        RECT 75.000 153.245 75.750 153.415 ;
        RECT 75.000 152.255 75.230 153.245 ;
        RECT 75.400 152.425 75.750 153.075 ;
        RECT 75.925 152.920 76.215 154.085 ;
        RECT 76.385 153.010 76.655 153.915 ;
        RECT 76.825 153.325 77.155 154.085 ;
        RECT 77.335 153.155 77.505 153.915 ;
        RECT 75.000 152.085 75.750 152.255 ;
        RECT 74.995 151.535 75.325 151.915 ;
        RECT 75.495 151.795 75.750 152.085 ;
        RECT 75.925 151.535 76.215 152.260 ;
        RECT 76.385 152.210 76.555 153.010 ;
        RECT 76.840 152.985 77.505 153.155 ;
        RECT 77.855 153.155 78.025 153.915 ;
        RECT 78.240 153.325 78.570 154.085 ;
        RECT 77.855 152.985 78.570 153.155 ;
        RECT 78.740 153.010 78.995 153.915 ;
        RECT 76.840 152.840 77.010 152.985 ;
        RECT 76.725 152.510 77.010 152.840 ;
        RECT 76.840 152.255 77.010 152.510 ;
        RECT 77.245 152.435 77.575 152.805 ;
        RECT 77.765 152.435 78.120 152.805 ;
        RECT 78.400 152.775 78.570 152.985 ;
        RECT 78.400 152.445 78.655 152.775 ;
        RECT 78.400 152.255 78.570 152.445 ;
        RECT 78.825 152.280 78.995 153.010 ;
        RECT 79.170 152.935 79.430 154.085 ;
        RECT 79.610 153.575 81.265 153.865 ;
        RECT 79.610 153.235 81.200 153.405 ;
        RECT 81.435 153.285 81.715 154.085 ;
        RECT 79.610 152.945 79.930 153.235 ;
        RECT 81.030 153.115 81.200 153.235 ;
        RECT 76.385 151.705 76.645 152.210 ;
        RECT 76.840 152.085 77.505 152.255 ;
        RECT 76.825 151.535 77.155 151.915 ;
        RECT 77.335 151.705 77.505 152.085 ;
        RECT 77.855 152.085 78.570 152.255 ;
        RECT 77.855 151.705 78.025 152.085 ;
        RECT 78.240 151.535 78.570 151.915 ;
        RECT 78.740 151.705 78.995 152.280 ;
        RECT 79.170 151.535 79.430 152.375 ;
        RECT 79.610 152.205 79.960 152.775 ;
        RECT 80.130 152.445 80.840 153.065 ;
        RECT 81.030 152.945 81.755 153.115 ;
        RECT 81.925 152.945 82.195 153.915 ;
        RECT 81.585 152.775 81.755 152.945 ;
        RECT 81.010 152.445 81.415 152.775 ;
        RECT 81.585 152.445 81.855 152.775 ;
        RECT 81.585 152.275 81.755 152.445 ;
        RECT 80.145 152.105 81.755 152.275 ;
        RECT 82.025 152.210 82.195 152.945 ;
        RECT 79.615 151.535 79.945 152.035 ;
        RECT 80.145 151.755 80.315 152.105 ;
        RECT 80.515 151.535 80.845 151.935 ;
        RECT 81.015 151.755 81.185 152.105 ;
        RECT 81.355 151.535 81.735 151.935 ;
        RECT 81.925 151.865 82.195 152.210 ;
        RECT 82.365 152.945 82.705 153.915 ;
        RECT 82.875 152.945 83.045 154.085 ;
        RECT 83.315 153.285 83.565 154.085 ;
        RECT 84.210 153.115 84.540 153.915 ;
        RECT 84.840 153.285 85.170 154.085 ;
        RECT 85.340 153.115 85.670 153.915 ;
        RECT 83.235 152.945 85.670 153.115 ;
        RECT 86.420 153.105 86.675 153.775 ;
        RECT 86.855 153.285 87.140 154.085 ;
        RECT 87.320 153.365 87.650 153.875 ;
        RECT 86.420 153.065 86.600 153.105 ;
        RECT 82.365 152.385 82.540 152.945 ;
        RECT 83.235 152.695 83.405 152.945 ;
        RECT 82.710 152.525 83.405 152.695 ;
        RECT 83.580 152.525 84.000 152.725 ;
        RECT 84.170 152.525 84.500 152.725 ;
        RECT 84.670 152.525 85.000 152.725 ;
        RECT 82.365 152.335 82.595 152.385 ;
        RECT 82.365 151.705 82.705 152.335 ;
        RECT 82.875 151.535 83.125 152.335 ;
        RECT 83.315 152.185 84.540 152.355 ;
        RECT 83.315 151.705 83.645 152.185 ;
        RECT 83.815 151.535 84.040 151.995 ;
        RECT 84.210 151.705 84.540 152.185 ;
        RECT 85.170 152.315 85.340 152.945 ;
        RECT 86.335 152.895 86.600 153.065 ;
        RECT 85.525 152.525 85.875 152.775 ;
        RECT 85.170 151.705 85.670 152.315 ;
        RECT 86.420 152.245 86.600 152.895 ;
        RECT 87.320 152.775 87.570 153.365 ;
        RECT 87.920 153.215 88.090 153.825 ;
        RECT 88.260 153.395 88.590 154.085 ;
        RECT 88.820 153.535 89.060 153.825 ;
        RECT 89.260 153.705 89.680 154.085 ;
        RECT 89.860 153.615 90.490 153.865 ;
        RECT 90.960 153.705 91.290 154.085 ;
        RECT 89.860 153.535 90.030 153.615 ;
        RECT 91.460 153.535 91.630 153.825 ;
        RECT 91.810 153.705 92.190 154.085 ;
        RECT 92.430 153.700 93.260 153.870 ;
        RECT 88.820 153.365 90.030 153.535 ;
        RECT 86.770 152.445 87.570 152.775 ;
        RECT 86.420 151.715 86.675 152.245 ;
        RECT 86.855 151.535 87.140 151.995 ;
        RECT 87.320 151.795 87.570 152.445 ;
        RECT 87.770 153.195 88.090 153.215 ;
        RECT 87.770 153.025 89.690 153.195 ;
        RECT 87.770 152.130 87.960 153.025 ;
        RECT 89.860 152.855 90.030 153.365 ;
        RECT 90.200 153.105 90.720 153.415 ;
        RECT 88.130 152.685 90.030 152.855 ;
        RECT 88.130 152.625 88.460 152.685 ;
        RECT 88.610 152.455 88.940 152.515 ;
        RECT 88.280 152.185 88.940 152.455 ;
        RECT 87.770 151.800 88.090 152.130 ;
        RECT 88.270 151.535 88.930 152.015 ;
        RECT 89.130 151.925 89.300 152.685 ;
        RECT 90.200 152.515 90.380 152.925 ;
        RECT 89.470 152.345 89.800 152.465 ;
        RECT 90.550 152.345 90.720 153.105 ;
        RECT 89.470 152.175 90.720 152.345 ;
        RECT 90.890 153.285 92.260 153.535 ;
        RECT 90.890 152.515 91.080 153.285 ;
        RECT 92.010 153.025 92.260 153.285 ;
        RECT 91.250 152.855 91.500 153.015 ;
        RECT 92.430 152.855 92.600 153.700 ;
        RECT 93.495 153.415 93.665 153.915 ;
        RECT 93.835 153.585 94.165 154.085 ;
        RECT 92.770 153.025 93.270 153.405 ;
        RECT 93.495 153.245 94.190 153.415 ;
        RECT 91.250 152.685 92.600 152.855 ;
        RECT 92.180 152.645 92.600 152.685 ;
        RECT 90.890 152.175 91.310 152.515 ;
        RECT 91.600 152.185 92.010 152.515 ;
        RECT 89.130 151.755 89.980 151.925 ;
        RECT 90.540 151.535 90.860 151.995 ;
        RECT 91.060 151.745 91.310 152.175 ;
        RECT 91.600 151.535 92.010 151.975 ;
        RECT 92.180 151.915 92.350 152.645 ;
        RECT 92.520 152.095 92.870 152.465 ;
        RECT 93.050 152.155 93.270 153.025 ;
        RECT 93.440 152.455 93.850 153.075 ;
        RECT 94.020 152.275 94.190 153.245 ;
        RECT 93.495 152.085 94.190 152.275 ;
        RECT 92.180 151.715 93.195 151.915 ;
        RECT 93.495 151.755 93.665 152.085 ;
        RECT 93.835 151.535 94.165 151.915 ;
        RECT 94.380 151.795 94.605 153.915 ;
        RECT 94.775 153.585 95.105 154.085 ;
        RECT 95.275 153.415 95.445 153.915 ;
        RECT 94.780 153.245 95.445 153.415 ;
        RECT 94.780 152.255 95.010 153.245 ;
        RECT 95.180 152.425 95.530 153.075 ;
        RECT 96.165 152.995 97.835 154.085 ;
        RECT 96.165 152.475 96.915 152.995 ;
        RECT 98.005 152.945 98.345 153.915 ;
        RECT 98.515 152.945 98.685 154.085 ;
        RECT 98.955 153.285 99.205 154.085 ;
        RECT 99.850 153.115 100.180 153.915 ;
        RECT 100.480 153.285 100.810 154.085 ;
        RECT 100.980 153.115 101.310 153.915 ;
        RECT 98.875 152.945 101.310 153.115 ;
        RECT 97.085 152.305 97.835 152.825 ;
        RECT 94.780 152.085 95.445 152.255 ;
        RECT 94.775 151.535 95.105 151.915 ;
        RECT 95.275 151.795 95.445 152.085 ;
        RECT 96.165 151.535 97.835 152.305 ;
        RECT 98.005 152.335 98.180 152.945 ;
        RECT 98.875 152.695 99.045 152.945 ;
        RECT 98.350 152.525 99.045 152.695 ;
        RECT 99.220 152.525 99.640 152.725 ;
        RECT 99.810 152.525 100.140 152.725 ;
        RECT 100.310 152.525 100.640 152.725 ;
        RECT 98.005 151.705 98.345 152.335 ;
        RECT 98.515 151.535 98.765 152.335 ;
        RECT 98.955 152.185 100.180 152.355 ;
        RECT 98.955 151.705 99.285 152.185 ;
        RECT 99.455 151.535 99.680 151.995 ;
        RECT 99.850 151.705 100.180 152.185 ;
        RECT 100.810 152.315 100.980 152.945 ;
        RECT 101.685 152.920 101.975 154.085 ;
        RECT 102.150 153.650 107.495 154.085 ;
        RECT 101.165 152.525 101.515 152.775 ;
        RECT 103.740 152.400 104.090 153.650 ;
        RECT 107.665 152.945 108.005 153.915 ;
        RECT 108.175 152.945 108.345 154.085 ;
        RECT 108.615 153.285 108.865 154.085 ;
        RECT 109.510 153.115 109.840 153.915 ;
        RECT 110.140 153.285 110.470 154.085 ;
        RECT 110.640 153.115 110.970 153.915 ;
        RECT 108.535 152.945 110.970 153.115 ;
        RECT 111.550 153.115 111.880 153.915 ;
        RECT 112.050 153.285 112.380 154.085 ;
        RECT 112.680 153.115 113.010 153.915 ;
        RECT 113.655 153.285 113.905 154.085 ;
        RECT 111.550 152.945 113.985 153.115 ;
        RECT 114.175 152.945 114.345 154.085 ;
        RECT 114.515 152.945 114.855 153.915 ;
        RECT 100.810 151.705 101.310 152.315 ;
        RECT 101.685 151.535 101.975 152.260 ;
        RECT 105.570 152.080 105.910 152.910 ;
        RECT 107.665 152.335 107.840 152.945 ;
        RECT 108.535 152.695 108.705 152.945 ;
        RECT 108.010 152.525 108.705 152.695 ;
        RECT 108.880 152.525 109.300 152.725 ;
        RECT 109.470 152.525 109.800 152.725 ;
        RECT 109.970 152.525 110.300 152.725 ;
        RECT 102.150 151.535 107.495 152.080 ;
        RECT 107.665 151.705 108.005 152.335 ;
        RECT 108.175 151.535 108.425 152.335 ;
        RECT 108.615 152.185 109.840 152.355 ;
        RECT 108.615 151.705 108.945 152.185 ;
        RECT 109.115 151.535 109.340 151.995 ;
        RECT 109.510 151.705 109.840 152.185 ;
        RECT 110.470 152.315 110.640 152.945 ;
        RECT 110.825 152.525 111.175 152.775 ;
        RECT 111.345 152.525 111.695 152.775 ;
        RECT 111.880 152.315 112.050 152.945 ;
        RECT 112.220 152.525 112.550 152.725 ;
        RECT 112.720 152.525 113.050 152.725 ;
        RECT 113.220 152.525 113.640 152.725 ;
        RECT 113.815 152.695 113.985 152.945 ;
        RECT 113.815 152.525 114.510 152.695 ;
        RECT 110.470 151.705 110.970 152.315 ;
        RECT 111.550 151.705 112.050 152.315 ;
        RECT 112.680 152.185 113.905 152.355 ;
        RECT 114.680 152.335 114.855 152.945 ;
        RECT 115.485 152.995 117.155 154.085 ;
        RECT 117.325 153.325 117.840 153.735 ;
        RECT 118.075 153.325 118.245 154.085 ;
        RECT 118.415 153.745 120.445 153.915 ;
        RECT 115.485 152.475 116.235 152.995 ;
        RECT 112.680 151.705 113.010 152.185 ;
        RECT 113.180 151.535 113.405 151.995 ;
        RECT 113.575 151.705 113.905 152.185 ;
        RECT 114.095 151.535 114.345 152.335 ;
        RECT 114.515 151.705 114.855 152.335 ;
        RECT 116.405 152.305 117.155 152.825 ;
        RECT 117.325 152.515 117.665 153.325 ;
        RECT 118.415 153.080 118.585 153.745 ;
        RECT 118.980 153.405 120.105 153.575 ;
        RECT 117.835 152.890 118.585 153.080 ;
        RECT 118.755 153.065 119.765 153.235 ;
        RECT 117.325 152.345 118.555 152.515 ;
        RECT 115.485 151.535 117.155 152.305 ;
        RECT 117.600 151.740 117.845 152.345 ;
        RECT 118.065 151.535 118.575 152.070 ;
        RECT 118.755 151.705 118.945 153.065 ;
        RECT 119.115 152.725 119.390 152.865 ;
        RECT 119.115 152.555 119.395 152.725 ;
        RECT 119.115 151.705 119.390 152.555 ;
        RECT 119.595 152.265 119.765 153.065 ;
        RECT 119.935 152.275 120.105 153.405 ;
        RECT 120.275 152.775 120.445 153.745 ;
        RECT 120.615 152.945 120.785 154.085 ;
        RECT 120.955 152.945 121.290 153.915 ;
        RECT 120.275 152.445 120.470 152.775 ;
        RECT 120.695 152.445 120.950 152.775 ;
        RECT 120.695 152.275 120.865 152.445 ;
        RECT 121.120 152.275 121.290 152.945 ;
        RECT 121.465 152.995 122.675 154.085 ;
        RECT 122.845 152.995 126.355 154.085 ;
        RECT 126.525 152.995 127.735 154.085 ;
        RECT 121.465 152.455 121.985 152.995 ;
        RECT 122.155 152.285 122.675 152.825 ;
        RECT 122.845 152.475 124.535 152.995 ;
        RECT 124.705 152.305 126.355 152.825 ;
        RECT 126.525 152.455 127.045 152.995 ;
        RECT 119.935 152.105 120.865 152.275 ;
        RECT 119.935 152.070 120.110 152.105 ;
        RECT 119.580 151.705 120.110 152.070 ;
        RECT 120.535 151.535 120.865 151.935 ;
        RECT 121.035 151.705 121.290 152.275 ;
        RECT 121.465 151.535 122.675 152.285 ;
        RECT 122.845 151.535 126.355 152.305 ;
        RECT 127.215 152.285 127.735 152.825 ;
        RECT 126.525 151.535 127.735 152.285 ;
        RECT 29.840 151.365 127.820 151.535 ;
        RECT 29.925 150.615 31.135 151.365 ;
        RECT 29.925 150.075 30.445 150.615 ;
        RECT 31.825 150.545 32.035 151.365 ;
        RECT 32.205 150.565 32.535 151.195 ;
        RECT 30.615 149.905 31.135 150.445 ;
        RECT 32.205 149.965 32.455 150.565 ;
        RECT 32.705 150.545 32.935 151.365 ;
        RECT 33.420 150.555 33.665 151.160 ;
        RECT 33.885 150.830 34.395 151.365 ;
        RECT 33.145 150.385 34.375 150.555 ;
        RECT 32.625 150.125 32.955 150.375 ;
        RECT 29.925 148.815 31.135 149.905 ;
        RECT 31.825 148.815 32.035 149.955 ;
        RECT 32.205 148.985 32.535 149.965 ;
        RECT 32.705 148.815 32.935 149.955 ;
        RECT 33.145 149.575 33.485 150.385 ;
        RECT 33.655 149.820 34.405 150.010 ;
        RECT 33.145 149.165 33.660 149.575 ;
        RECT 33.895 148.815 34.065 149.575 ;
        RECT 34.235 149.155 34.405 149.820 ;
        RECT 34.575 149.835 34.765 151.195 ;
        RECT 34.935 151.025 35.210 151.195 ;
        RECT 34.935 150.855 35.215 151.025 ;
        RECT 34.935 150.035 35.210 150.855 ;
        RECT 35.400 150.830 35.930 151.195 ;
        RECT 36.355 150.965 36.685 151.365 ;
        RECT 35.755 150.795 35.930 150.830 ;
        RECT 35.415 149.835 35.585 150.635 ;
        RECT 34.575 149.665 35.585 149.835 ;
        RECT 35.755 150.625 36.685 150.795 ;
        RECT 36.855 150.625 37.110 151.195 ;
        RECT 37.285 150.640 37.575 151.365 ;
        RECT 38.120 150.655 38.375 151.185 ;
        RECT 38.555 150.905 38.840 151.365 ;
        RECT 35.755 149.495 35.925 150.625 ;
        RECT 36.515 150.455 36.685 150.625 ;
        RECT 34.800 149.325 35.925 149.495 ;
        RECT 36.095 150.125 36.290 150.455 ;
        RECT 36.515 150.125 36.770 150.455 ;
        RECT 36.095 149.155 36.265 150.125 ;
        RECT 36.940 149.955 37.110 150.625 ;
        RECT 34.235 148.985 36.265 149.155 ;
        RECT 36.435 148.815 36.605 149.955 ;
        RECT 36.775 148.985 37.110 149.955 ;
        RECT 37.285 148.815 37.575 149.980 ;
        RECT 38.120 149.795 38.300 150.655 ;
        RECT 39.020 150.455 39.270 151.105 ;
        RECT 38.470 150.125 39.270 150.455 ;
        RECT 38.120 149.325 38.375 149.795 ;
        RECT 38.035 149.155 38.375 149.325 ;
        RECT 38.120 149.125 38.375 149.155 ;
        RECT 38.555 148.815 38.840 149.615 ;
        RECT 39.020 149.535 39.270 150.125 ;
        RECT 39.470 150.770 39.790 151.100 ;
        RECT 39.970 150.885 40.630 151.365 ;
        RECT 40.830 150.975 41.680 151.145 ;
        RECT 39.470 149.875 39.660 150.770 ;
        RECT 39.980 150.445 40.640 150.715 ;
        RECT 40.310 150.385 40.640 150.445 ;
        RECT 39.830 150.215 40.160 150.275 ;
        RECT 40.830 150.215 41.000 150.975 ;
        RECT 42.240 150.905 42.560 151.365 ;
        RECT 42.760 150.725 43.010 151.155 ;
        RECT 43.300 150.925 43.710 151.365 ;
        RECT 43.880 150.985 44.895 151.185 ;
        RECT 41.170 150.555 42.420 150.725 ;
        RECT 41.170 150.435 41.500 150.555 ;
        RECT 39.830 150.045 41.730 150.215 ;
        RECT 39.470 149.705 41.390 149.875 ;
        RECT 39.470 149.685 39.790 149.705 ;
        RECT 39.020 149.025 39.350 149.535 ;
        RECT 39.620 149.075 39.790 149.685 ;
        RECT 41.560 149.535 41.730 150.045 ;
        RECT 41.900 149.975 42.080 150.385 ;
        RECT 42.250 149.795 42.420 150.555 ;
        RECT 39.960 148.815 40.290 149.505 ;
        RECT 40.520 149.365 41.730 149.535 ;
        RECT 41.900 149.485 42.420 149.795 ;
        RECT 42.590 150.385 43.010 150.725 ;
        RECT 43.300 150.385 43.710 150.715 ;
        RECT 42.590 149.615 42.780 150.385 ;
        RECT 43.880 150.255 44.050 150.985 ;
        RECT 45.195 150.815 45.365 151.145 ;
        RECT 45.535 150.985 45.865 151.365 ;
        RECT 44.220 150.435 44.570 150.805 ;
        RECT 43.880 150.215 44.300 150.255 ;
        RECT 42.950 150.045 44.300 150.215 ;
        RECT 42.950 149.885 43.200 150.045 ;
        RECT 43.710 149.615 43.960 149.875 ;
        RECT 42.590 149.365 43.960 149.615 ;
        RECT 40.520 149.075 40.760 149.365 ;
        RECT 41.560 149.285 41.730 149.365 ;
        RECT 40.960 148.815 41.380 149.195 ;
        RECT 41.560 149.035 42.190 149.285 ;
        RECT 42.660 148.815 42.990 149.195 ;
        RECT 43.160 149.075 43.330 149.365 ;
        RECT 44.130 149.200 44.300 150.045 ;
        RECT 44.750 149.875 44.970 150.745 ;
        RECT 45.195 150.625 45.890 150.815 ;
        RECT 44.470 149.495 44.970 149.875 ;
        RECT 45.140 149.825 45.550 150.445 ;
        RECT 45.720 149.655 45.890 150.625 ;
        RECT 45.195 149.485 45.890 149.655 ;
        RECT 43.510 148.815 43.890 149.195 ;
        RECT 44.130 149.030 44.960 149.200 ;
        RECT 45.195 148.985 45.365 149.485 ;
        RECT 45.535 148.815 45.865 149.315 ;
        RECT 46.080 148.985 46.305 151.105 ;
        RECT 46.475 150.985 46.805 151.365 ;
        RECT 46.975 150.815 47.145 151.105 ;
        RECT 46.480 150.645 47.145 150.815 ;
        RECT 47.405 150.905 47.965 151.195 ;
        RECT 48.135 150.905 48.385 151.365 ;
        RECT 46.480 149.655 46.710 150.645 ;
        RECT 46.880 149.825 47.230 150.475 ;
        RECT 46.480 149.485 47.145 149.655 ;
        RECT 46.475 148.815 46.805 149.315 ;
        RECT 46.975 148.985 47.145 149.485 ;
        RECT 47.405 149.535 47.655 150.905 ;
        RECT 49.005 150.735 49.335 151.095 ;
        RECT 47.945 150.545 49.335 150.735 ;
        RECT 49.705 150.905 50.265 151.195 ;
        RECT 50.435 150.905 50.685 151.365 ;
        RECT 47.945 150.455 48.115 150.545 ;
        RECT 47.825 150.125 48.115 150.455 ;
        RECT 48.285 150.125 48.625 150.375 ;
        RECT 48.845 150.125 49.520 150.375 ;
        RECT 47.945 149.875 48.115 150.125 ;
        RECT 47.945 149.705 48.885 149.875 ;
        RECT 49.255 149.765 49.520 150.125 ;
        RECT 47.405 148.985 47.865 149.535 ;
        RECT 48.055 148.815 48.385 149.535 ;
        RECT 48.585 149.155 48.885 149.705 ;
        RECT 49.705 149.535 49.955 150.905 ;
        RECT 51.305 150.735 51.635 151.095 ;
        RECT 50.245 150.545 51.635 150.735 ;
        RECT 52.925 150.565 53.265 151.195 ;
        RECT 53.435 150.565 53.685 151.365 ;
        RECT 53.875 150.715 54.205 151.195 ;
        RECT 54.375 150.905 54.600 151.365 ;
        RECT 54.770 150.715 55.100 151.195 ;
        RECT 50.245 150.455 50.415 150.545 ;
        RECT 50.125 150.125 50.415 150.455 ;
        RECT 50.585 150.125 50.925 150.375 ;
        RECT 51.145 150.125 51.820 150.375 ;
        RECT 50.245 149.875 50.415 150.125 ;
        RECT 50.245 149.705 51.185 149.875 ;
        RECT 51.555 149.765 51.820 150.125 ;
        RECT 52.925 149.955 53.100 150.565 ;
        RECT 53.875 150.545 55.100 150.715 ;
        RECT 55.730 150.585 56.230 151.195 ;
        RECT 53.270 150.205 53.965 150.375 ;
        RECT 53.795 149.955 53.965 150.205 ;
        RECT 54.140 150.175 54.560 150.375 ;
        RECT 54.730 150.175 55.060 150.375 ;
        RECT 55.230 150.175 55.560 150.375 ;
        RECT 55.730 149.955 55.900 150.585 ;
        RECT 57.800 150.555 58.045 151.160 ;
        RECT 58.265 150.830 58.775 151.365 ;
        RECT 57.525 150.385 58.755 150.555 ;
        RECT 56.085 150.125 56.435 150.375 ;
        RECT 49.055 148.815 49.335 149.485 ;
        RECT 49.705 148.985 50.165 149.535 ;
        RECT 50.355 148.815 50.685 149.535 ;
        RECT 50.885 149.155 51.185 149.705 ;
        RECT 51.355 148.815 51.635 149.485 ;
        RECT 52.925 148.985 53.265 149.955 ;
        RECT 53.435 148.815 53.605 149.955 ;
        RECT 53.795 149.785 56.230 149.955 ;
        RECT 53.875 148.815 54.125 149.615 ;
        RECT 54.770 148.985 55.100 149.785 ;
        RECT 55.400 148.815 55.730 149.615 ;
        RECT 55.900 148.985 56.230 149.785 ;
        RECT 57.525 149.575 57.865 150.385 ;
        RECT 58.035 149.820 58.785 150.010 ;
        RECT 57.525 149.165 58.040 149.575 ;
        RECT 58.275 148.815 58.445 149.575 ;
        RECT 58.615 149.155 58.785 149.820 ;
        RECT 58.955 149.835 59.145 151.195 ;
        RECT 59.315 151.025 59.590 151.195 ;
        RECT 59.315 150.855 59.595 151.025 ;
        RECT 59.315 150.035 59.590 150.855 ;
        RECT 59.780 150.830 60.310 151.195 ;
        RECT 60.735 150.965 61.065 151.365 ;
        RECT 60.135 150.795 60.310 150.830 ;
        RECT 59.795 149.835 59.965 150.635 ;
        RECT 58.955 149.665 59.965 149.835 ;
        RECT 60.135 150.625 61.065 150.795 ;
        RECT 61.235 150.625 61.490 151.195 ;
        RECT 60.135 149.495 60.305 150.625 ;
        RECT 60.895 150.455 61.065 150.625 ;
        RECT 59.180 149.325 60.305 149.495 ;
        RECT 60.475 150.125 60.670 150.455 ;
        RECT 60.895 150.125 61.150 150.455 ;
        RECT 60.475 149.155 60.645 150.125 ;
        RECT 61.320 149.955 61.490 150.625 ;
        RECT 58.615 148.985 60.645 149.155 ;
        RECT 60.815 148.815 60.985 149.955 ;
        RECT 61.155 148.985 61.490 149.955 ;
        RECT 61.665 150.690 61.925 151.195 ;
        RECT 62.105 150.985 62.435 151.365 ;
        RECT 62.615 150.815 62.785 151.195 ;
        RECT 61.665 149.890 61.835 150.690 ;
        RECT 62.120 150.645 62.785 150.815 ;
        RECT 62.120 150.390 62.290 150.645 ;
        RECT 63.045 150.640 63.335 151.365 ;
        RECT 63.505 150.615 64.715 151.365 ;
        RECT 62.005 150.060 62.290 150.390 ;
        RECT 62.525 150.095 62.855 150.465 ;
        RECT 62.120 149.915 62.290 150.060 ;
        RECT 61.665 148.985 61.935 149.890 ;
        RECT 62.120 149.745 62.785 149.915 ;
        RECT 62.105 148.815 62.435 149.575 ;
        RECT 62.615 148.985 62.785 149.745 ;
        RECT 63.045 148.815 63.335 149.980 ;
        RECT 63.505 149.905 64.025 150.445 ;
        RECT 64.195 150.075 64.715 150.615 ;
        RECT 64.885 150.565 65.225 151.195 ;
        RECT 65.395 150.565 65.645 151.365 ;
        RECT 65.835 150.715 66.165 151.195 ;
        RECT 66.335 150.905 66.560 151.365 ;
        RECT 66.730 150.715 67.060 151.195 ;
        RECT 64.885 149.955 65.060 150.565 ;
        RECT 65.835 150.545 67.060 150.715 ;
        RECT 67.690 150.585 68.190 151.195 ;
        RECT 65.230 150.205 65.925 150.375 ;
        RECT 65.755 149.955 65.925 150.205 ;
        RECT 66.100 150.175 66.520 150.375 ;
        RECT 66.690 150.175 67.020 150.375 ;
        RECT 67.190 150.175 67.520 150.375 ;
        RECT 67.690 149.955 67.860 150.585 ;
        RECT 68.605 150.545 68.835 151.365 ;
        RECT 69.005 150.565 69.335 151.195 ;
        RECT 68.045 150.125 68.395 150.375 ;
        RECT 68.585 150.125 68.915 150.375 ;
        RECT 69.085 149.965 69.335 150.565 ;
        RECT 69.505 150.545 69.715 151.365 ;
        RECT 70.320 150.655 70.575 151.185 ;
        RECT 70.755 150.905 71.040 151.365 ;
        RECT 63.505 148.815 64.715 149.905 ;
        RECT 64.885 148.985 65.225 149.955 ;
        RECT 65.395 148.815 65.565 149.955 ;
        RECT 65.755 149.785 68.190 149.955 ;
        RECT 65.835 148.815 66.085 149.615 ;
        RECT 66.730 148.985 67.060 149.785 ;
        RECT 67.360 148.815 67.690 149.615 ;
        RECT 67.860 148.985 68.190 149.785 ;
        RECT 68.605 148.815 68.835 149.955 ;
        RECT 69.005 148.985 69.335 149.965 ;
        RECT 69.505 148.815 69.715 149.955 ;
        RECT 70.320 149.795 70.500 150.655 ;
        RECT 71.220 150.455 71.470 151.105 ;
        RECT 70.670 150.125 71.470 150.455 ;
        RECT 70.320 149.325 70.575 149.795 ;
        RECT 70.235 149.155 70.575 149.325 ;
        RECT 70.320 149.125 70.575 149.155 ;
        RECT 70.755 148.815 71.040 149.615 ;
        RECT 71.220 149.535 71.470 150.125 ;
        RECT 71.670 150.770 71.990 151.100 ;
        RECT 72.170 150.885 72.830 151.365 ;
        RECT 73.030 150.975 73.880 151.145 ;
        RECT 71.670 149.875 71.860 150.770 ;
        RECT 72.180 150.445 72.840 150.715 ;
        RECT 72.510 150.385 72.840 150.445 ;
        RECT 72.030 150.215 72.360 150.275 ;
        RECT 73.030 150.215 73.200 150.975 ;
        RECT 74.440 150.905 74.760 151.365 ;
        RECT 74.960 150.725 75.210 151.155 ;
        RECT 75.500 150.925 75.910 151.365 ;
        RECT 76.080 150.985 77.095 151.185 ;
        RECT 73.370 150.555 74.620 150.725 ;
        RECT 73.370 150.435 73.700 150.555 ;
        RECT 72.030 150.045 73.930 150.215 ;
        RECT 71.670 149.705 73.590 149.875 ;
        RECT 71.670 149.685 71.990 149.705 ;
        RECT 71.220 149.025 71.550 149.535 ;
        RECT 71.820 149.075 71.990 149.685 ;
        RECT 73.760 149.535 73.930 150.045 ;
        RECT 74.100 149.975 74.280 150.385 ;
        RECT 74.450 149.795 74.620 150.555 ;
        RECT 72.160 148.815 72.490 149.505 ;
        RECT 72.720 149.365 73.930 149.535 ;
        RECT 74.100 149.485 74.620 149.795 ;
        RECT 74.790 150.385 75.210 150.725 ;
        RECT 75.500 150.385 75.910 150.715 ;
        RECT 74.790 149.615 74.980 150.385 ;
        RECT 76.080 150.255 76.250 150.985 ;
        RECT 77.395 150.815 77.565 151.145 ;
        RECT 77.735 150.985 78.065 151.365 ;
        RECT 76.420 150.435 76.770 150.805 ;
        RECT 76.080 150.215 76.500 150.255 ;
        RECT 75.150 150.045 76.500 150.215 ;
        RECT 75.150 149.885 75.400 150.045 ;
        RECT 75.910 149.615 76.160 149.875 ;
        RECT 74.790 149.365 76.160 149.615 ;
        RECT 72.720 149.075 72.960 149.365 ;
        RECT 73.760 149.285 73.930 149.365 ;
        RECT 73.160 148.815 73.580 149.195 ;
        RECT 73.760 149.035 74.390 149.285 ;
        RECT 74.860 148.815 75.190 149.195 ;
        RECT 75.360 149.075 75.530 149.365 ;
        RECT 76.330 149.200 76.500 150.045 ;
        RECT 76.950 149.875 77.170 150.745 ;
        RECT 77.395 150.625 78.090 150.815 ;
        RECT 76.670 149.495 77.170 149.875 ;
        RECT 77.340 149.825 77.750 150.445 ;
        RECT 77.920 149.655 78.090 150.625 ;
        RECT 77.395 149.485 78.090 149.655 ;
        RECT 75.710 148.815 76.090 149.195 ;
        RECT 76.330 149.030 77.160 149.200 ;
        RECT 77.395 148.985 77.565 149.485 ;
        RECT 77.735 148.815 78.065 149.315 ;
        RECT 78.280 148.985 78.505 151.105 ;
        RECT 78.675 150.985 79.005 151.365 ;
        RECT 79.175 150.815 79.345 151.105 ;
        RECT 78.680 150.645 79.345 150.815 ;
        RECT 79.605 150.690 79.865 151.195 ;
        RECT 80.045 150.985 80.375 151.365 ;
        RECT 80.555 150.815 80.725 151.195 ;
        RECT 78.680 149.655 78.910 150.645 ;
        RECT 79.080 149.825 79.430 150.475 ;
        RECT 79.605 149.890 79.775 150.690 ;
        RECT 80.060 150.645 80.725 150.815 ;
        RECT 80.060 150.390 80.230 150.645 ;
        RECT 80.985 150.595 84.495 151.365 ;
        RECT 79.945 150.060 80.230 150.390 ;
        RECT 80.465 150.095 80.795 150.465 ;
        RECT 80.060 149.915 80.230 150.060 ;
        RECT 78.680 149.485 79.345 149.655 ;
        RECT 78.675 148.815 79.005 149.315 ;
        RECT 79.175 148.985 79.345 149.485 ;
        RECT 79.605 148.985 79.875 149.890 ;
        RECT 80.060 149.745 80.725 149.915 ;
        RECT 80.045 148.815 80.375 149.575 ;
        RECT 80.555 148.985 80.725 149.745 ;
        RECT 80.985 149.905 82.675 150.425 ;
        RECT 82.845 150.075 84.495 150.595 ;
        RECT 84.940 150.555 85.185 151.160 ;
        RECT 85.405 150.830 85.915 151.365 ;
        RECT 84.665 150.385 85.895 150.555 ;
        RECT 80.985 148.815 84.495 149.905 ;
        RECT 84.665 149.575 85.005 150.385 ;
        RECT 85.175 149.820 85.925 150.010 ;
        RECT 84.665 149.165 85.180 149.575 ;
        RECT 85.415 148.815 85.585 149.575 ;
        RECT 85.755 149.155 85.925 149.820 ;
        RECT 86.095 149.835 86.285 151.195 ;
        RECT 86.455 150.345 86.730 151.195 ;
        RECT 86.920 150.830 87.450 151.195 ;
        RECT 87.875 150.965 88.205 151.365 ;
        RECT 87.275 150.795 87.450 150.830 ;
        RECT 86.455 150.175 86.735 150.345 ;
        RECT 86.455 150.035 86.730 150.175 ;
        RECT 86.935 149.835 87.105 150.635 ;
        RECT 86.095 149.665 87.105 149.835 ;
        RECT 87.275 150.625 88.205 150.795 ;
        RECT 88.375 150.625 88.630 151.195 ;
        RECT 88.805 150.640 89.095 151.365 ;
        RECT 87.275 149.495 87.445 150.625 ;
        RECT 88.035 150.455 88.205 150.625 ;
        RECT 86.320 149.325 87.445 149.495 ;
        RECT 87.615 150.125 87.810 150.455 ;
        RECT 88.035 150.125 88.290 150.455 ;
        RECT 87.615 149.155 87.785 150.125 ;
        RECT 88.460 149.955 88.630 150.625 ;
        RECT 89.725 150.595 91.395 151.365 ;
        RECT 91.655 150.815 91.825 151.195 ;
        RECT 92.005 150.985 92.335 151.365 ;
        RECT 91.655 150.645 92.320 150.815 ;
        RECT 92.515 150.690 92.775 151.195 ;
        RECT 85.755 148.985 87.785 149.155 ;
        RECT 87.955 148.815 88.125 149.955 ;
        RECT 88.295 148.985 88.630 149.955 ;
        RECT 88.805 148.815 89.095 149.980 ;
        RECT 89.725 149.905 90.475 150.425 ;
        RECT 90.645 150.075 91.395 150.595 ;
        RECT 91.585 150.095 91.915 150.465 ;
        RECT 92.150 150.390 92.320 150.645 ;
        RECT 92.150 150.060 92.435 150.390 ;
        RECT 92.150 149.915 92.320 150.060 ;
        RECT 89.725 148.815 91.395 149.905 ;
        RECT 91.655 149.745 92.320 149.915 ;
        RECT 92.605 149.890 92.775 150.690 ;
        RECT 93.405 150.595 96.915 151.365 ;
        RECT 91.655 148.985 91.825 149.745 ;
        RECT 92.005 148.815 92.335 149.575 ;
        RECT 92.505 148.985 92.775 149.890 ;
        RECT 93.405 149.905 95.095 150.425 ;
        RECT 95.265 150.075 96.915 150.595 ;
        RECT 97.460 150.655 97.715 151.185 ;
        RECT 97.895 150.905 98.180 151.365 ;
        RECT 93.405 148.815 96.915 149.905 ;
        RECT 97.460 149.795 97.640 150.655 ;
        RECT 98.360 150.455 98.610 151.105 ;
        RECT 97.810 150.125 98.610 150.455 ;
        RECT 97.460 149.325 97.715 149.795 ;
        RECT 97.375 149.155 97.715 149.325 ;
        RECT 97.460 149.125 97.715 149.155 ;
        RECT 97.895 148.815 98.180 149.615 ;
        RECT 98.360 149.535 98.610 150.125 ;
        RECT 98.810 150.770 99.130 151.100 ;
        RECT 99.310 150.885 99.970 151.365 ;
        RECT 100.170 150.975 101.020 151.145 ;
        RECT 98.810 149.875 99.000 150.770 ;
        RECT 99.320 150.445 99.980 150.715 ;
        RECT 99.650 150.385 99.980 150.445 ;
        RECT 99.170 150.215 99.500 150.275 ;
        RECT 100.170 150.215 100.340 150.975 ;
        RECT 101.580 150.905 101.900 151.365 ;
        RECT 102.100 150.725 102.350 151.155 ;
        RECT 102.640 150.925 103.050 151.365 ;
        RECT 103.220 150.985 104.235 151.185 ;
        RECT 100.510 150.555 101.760 150.725 ;
        RECT 100.510 150.435 100.840 150.555 ;
        RECT 99.170 150.045 101.070 150.215 ;
        RECT 98.810 149.705 100.730 149.875 ;
        RECT 98.810 149.685 99.130 149.705 ;
        RECT 98.360 149.025 98.690 149.535 ;
        RECT 98.960 149.075 99.130 149.685 ;
        RECT 100.900 149.535 101.070 150.045 ;
        RECT 101.240 149.975 101.420 150.385 ;
        RECT 101.590 149.795 101.760 150.555 ;
        RECT 99.300 148.815 99.630 149.505 ;
        RECT 99.860 149.365 101.070 149.535 ;
        RECT 101.240 149.485 101.760 149.795 ;
        RECT 101.930 150.385 102.350 150.725 ;
        RECT 102.640 150.385 103.050 150.715 ;
        RECT 101.930 149.615 102.120 150.385 ;
        RECT 103.220 150.255 103.390 150.985 ;
        RECT 104.535 150.815 104.705 151.145 ;
        RECT 104.875 150.985 105.205 151.365 ;
        RECT 103.560 150.435 103.910 150.805 ;
        RECT 103.220 150.215 103.640 150.255 ;
        RECT 102.290 150.045 103.640 150.215 ;
        RECT 102.290 149.885 102.540 150.045 ;
        RECT 103.050 149.615 103.300 149.875 ;
        RECT 101.930 149.365 103.300 149.615 ;
        RECT 99.860 149.075 100.100 149.365 ;
        RECT 100.900 149.285 101.070 149.365 ;
        RECT 100.300 148.815 100.720 149.195 ;
        RECT 100.900 149.035 101.530 149.285 ;
        RECT 102.000 148.815 102.330 149.195 ;
        RECT 102.500 149.075 102.670 149.365 ;
        RECT 103.470 149.200 103.640 150.045 ;
        RECT 104.090 149.875 104.310 150.745 ;
        RECT 104.535 150.625 105.230 150.815 ;
        RECT 103.810 149.495 104.310 149.875 ;
        RECT 104.480 149.825 104.890 150.445 ;
        RECT 105.060 149.655 105.230 150.625 ;
        RECT 104.535 149.485 105.230 149.655 ;
        RECT 102.850 148.815 103.230 149.195 ;
        RECT 103.470 149.030 104.300 149.200 ;
        RECT 104.535 148.985 104.705 149.485 ;
        RECT 104.875 148.815 105.205 149.315 ;
        RECT 105.420 148.985 105.645 151.105 ;
        RECT 105.815 150.985 106.145 151.365 ;
        RECT 106.315 150.815 106.485 151.105 ;
        RECT 105.820 150.645 106.485 150.815 ;
        RECT 105.820 149.655 106.050 150.645 ;
        RECT 106.745 150.615 107.955 151.365 ;
        RECT 106.220 149.825 106.570 150.475 ;
        RECT 106.745 149.905 107.265 150.445 ;
        RECT 107.435 150.075 107.955 150.615 ;
        RECT 108.125 150.565 108.465 151.195 ;
        RECT 108.635 150.565 108.885 151.365 ;
        RECT 109.075 150.715 109.405 151.195 ;
        RECT 109.575 150.905 109.800 151.365 ;
        RECT 109.970 150.715 110.300 151.195 ;
        RECT 108.125 149.955 108.300 150.565 ;
        RECT 109.075 150.545 110.300 150.715 ;
        RECT 110.930 150.585 111.430 151.195 ;
        RECT 111.805 150.615 113.015 151.365 ;
        RECT 108.470 150.205 109.165 150.375 ;
        RECT 108.995 149.955 109.165 150.205 ;
        RECT 109.340 150.175 109.760 150.375 ;
        RECT 109.930 150.175 110.260 150.375 ;
        RECT 110.430 150.175 110.760 150.375 ;
        RECT 110.930 149.955 111.100 150.585 ;
        RECT 111.285 150.125 111.635 150.375 ;
        RECT 105.820 149.485 106.485 149.655 ;
        RECT 105.815 148.815 106.145 149.315 ;
        RECT 106.315 148.985 106.485 149.485 ;
        RECT 106.745 148.815 107.955 149.905 ;
        RECT 108.125 148.985 108.465 149.955 ;
        RECT 108.635 148.815 108.805 149.955 ;
        RECT 108.995 149.785 111.430 149.955 ;
        RECT 109.075 148.815 109.325 149.615 ;
        RECT 109.970 148.985 110.300 149.785 ;
        RECT 110.600 148.815 110.930 149.615 ;
        RECT 111.100 148.985 111.430 149.785 ;
        RECT 111.805 149.905 112.325 150.445 ;
        RECT 112.495 150.075 113.015 150.615 ;
        RECT 113.225 150.545 113.455 151.365 ;
        RECT 113.625 150.565 113.955 151.195 ;
        RECT 113.205 150.125 113.535 150.375 ;
        RECT 113.705 149.965 113.955 150.565 ;
        RECT 114.125 150.545 114.335 151.365 ;
        RECT 114.565 150.640 114.855 151.365 ;
        RECT 115.525 150.545 115.755 151.365 ;
        RECT 115.925 150.565 116.255 151.195 ;
        RECT 115.505 150.125 115.835 150.375 ;
        RECT 111.805 148.815 113.015 149.905 ;
        RECT 113.225 148.815 113.455 149.955 ;
        RECT 113.625 148.985 113.955 149.965 ;
        RECT 114.125 148.815 114.335 149.955 ;
        RECT 114.565 148.815 114.855 149.980 ;
        RECT 116.005 149.965 116.255 150.565 ;
        RECT 116.425 150.545 116.635 151.365 ;
        RECT 117.240 150.655 117.495 151.185 ;
        RECT 117.675 150.905 117.960 151.365 ;
        RECT 117.240 150.345 117.420 150.655 ;
        RECT 118.140 150.455 118.390 151.105 ;
        RECT 117.155 150.175 117.420 150.345 ;
        RECT 115.525 148.815 115.755 149.955 ;
        RECT 115.925 148.985 116.255 149.965 ;
        RECT 116.425 148.815 116.635 149.955 ;
        RECT 117.240 149.795 117.420 150.175 ;
        RECT 117.590 150.125 118.390 150.455 ;
        RECT 117.240 149.125 117.495 149.795 ;
        RECT 117.675 148.815 117.960 149.615 ;
        RECT 118.140 149.535 118.390 150.125 ;
        RECT 118.590 150.770 118.910 151.100 ;
        RECT 119.090 150.885 119.750 151.365 ;
        RECT 119.950 150.975 120.800 151.145 ;
        RECT 118.590 149.875 118.780 150.770 ;
        RECT 119.100 150.445 119.760 150.715 ;
        RECT 119.430 150.385 119.760 150.445 ;
        RECT 118.950 150.215 119.280 150.275 ;
        RECT 119.950 150.215 120.120 150.975 ;
        RECT 121.360 150.905 121.680 151.365 ;
        RECT 121.880 150.725 122.130 151.155 ;
        RECT 122.420 150.925 122.830 151.365 ;
        RECT 123.000 150.985 124.015 151.185 ;
        RECT 120.290 150.555 121.540 150.725 ;
        RECT 120.290 150.435 120.620 150.555 ;
        RECT 118.950 150.045 120.850 150.215 ;
        RECT 118.590 149.705 120.510 149.875 ;
        RECT 118.590 149.685 118.910 149.705 ;
        RECT 118.140 149.025 118.470 149.535 ;
        RECT 118.740 149.075 118.910 149.685 ;
        RECT 120.680 149.535 120.850 150.045 ;
        RECT 121.020 149.975 121.200 150.385 ;
        RECT 121.370 149.795 121.540 150.555 ;
        RECT 119.080 148.815 119.410 149.505 ;
        RECT 119.640 149.365 120.850 149.535 ;
        RECT 121.020 149.485 121.540 149.795 ;
        RECT 121.710 150.385 122.130 150.725 ;
        RECT 122.420 150.385 122.830 150.715 ;
        RECT 121.710 149.615 121.900 150.385 ;
        RECT 123.000 150.255 123.170 150.985 ;
        RECT 124.315 150.815 124.485 151.145 ;
        RECT 124.655 150.985 124.985 151.365 ;
        RECT 123.340 150.435 123.690 150.805 ;
        RECT 123.000 150.215 123.420 150.255 ;
        RECT 122.070 150.045 123.420 150.215 ;
        RECT 122.070 149.885 122.320 150.045 ;
        RECT 122.830 149.615 123.080 149.875 ;
        RECT 121.710 149.365 123.080 149.615 ;
        RECT 119.640 149.075 119.880 149.365 ;
        RECT 120.680 149.285 120.850 149.365 ;
        RECT 120.080 148.815 120.500 149.195 ;
        RECT 120.680 149.035 121.310 149.285 ;
        RECT 121.780 148.815 122.110 149.195 ;
        RECT 122.280 149.075 122.450 149.365 ;
        RECT 123.250 149.200 123.420 150.045 ;
        RECT 123.870 149.875 124.090 150.745 ;
        RECT 124.315 150.625 125.010 150.815 ;
        RECT 123.590 149.495 124.090 149.875 ;
        RECT 124.260 149.825 124.670 150.445 ;
        RECT 124.840 149.655 125.010 150.625 ;
        RECT 124.315 149.485 125.010 149.655 ;
        RECT 122.630 148.815 123.010 149.195 ;
        RECT 123.250 149.030 124.080 149.200 ;
        RECT 124.315 148.985 124.485 149.485 ;
        RECT 124.655 148.815 124.985 149.315 ;
        RECT 125.200 148.985 125.425 151.105 ;
        RECT 125.595 150.985 125.925 151.365 ;
        RECT 126.095 150.815 126.265 151.105 ;
        RECT 125.600 150.645 126.265 150.815 ;
        RECT 125.600 149.655 125.830 150.645 ;
        RECT 126.525 150.615 127.735 151.365 ;
        RECT 126.000 149.825 126.350 150.475 ;
        RECT 126.525 149.905 127.045 150.445 ;
        RECT 127.215 150.075 127.735 150.615 ;
        RECT 125.600 149.485 126.265 149.655 ;
        RECT 125.595 148.815 125.925 149.315 ;
        RECT 126.095 148.985 126.265 149.485 ;
        RECT 126.525 148.815 127.735 149.905 ;
        RECT 29.840 148.645 127.820 148.815 ;
        RECT 29.925 147.555 31.135 148.645 ;
        RECT 29.925 146.845 30.445 147.385 ;
        RECT 30.615 147.015 31.135 147.555 ;
        RECT 31.680 147.665 31.935 148.335 ;
        RECT 32.115 147.845 32.400 148.645 ;
        RECT 32.580 147.925 32.910 148.435 ;
        RECT 29.925 146.095 31.135 146.845 ;
        RECT 31.680 146.805 31.860 147.665 ;
        RECT 32.580 147.335 32.830 147.925 ;
        RECT 33.180 147.775 33.350 148.385 ;
        RECT 33.520 147.955 33.850 148.645 ;
        RECT 34.080 148.095 34.320 148.385 ;
        RECT 34.520 148.265 34.940 148.645 ;
        RECT 35.120 148.175 35.750 148.425 ;
        RECT 36.220 148.265 36.550 148.645 ;
        RECT 35.120 148.095 35.290 148.175 ;
        RECT 36.720 148.095 36.890 148.385 ;
        RECT 37.070 148.265 37.450 148.645 ;
        RECT 37.690 148.260 38.520 148.430 ;
        RECT 34.080 147.925 35.290 148.095 ;
        RECT 32.030 147.005 32.830 147.335 ;
        RECT 31.680 146.605 31.935 146.805 ;
        RECT 31.595 146.435 31.935 146.605 ;
        RECT 31.680 146.275 31.935 146.435 ;
        RECT 32.115 146.095 32.400 146.555 ;
        RECT 32.580 146.355 32.830 147.005 ;
        RECT 33.030 147.755 33.350 147.775 ;
        RECT 33.030 147.585 34.950 147.755 ;
        RECT 33.030 146.690 33.220 147.585 ;
        RECT 35.120 147.415 35.290 147.925 ;
        RECT 35.460 147.665 35.980 147.975 ;
        RECT 33.390 147.245 35.290 147.415 ;
        RECT 33.390 147.185 33.720 147.245 ;
        RECT 33.870 147.015 34.200 147.075 ;
        RECT 33.540 146.745 34.200 147.015 ;
        RECT 33.030 146.360 33.350 146.690 ;
        RECT 33.530 146.095 34.190 146.575 ;
        RECT 34.390 146.485 34.560 147.245 ;
        RECT 35.460 147.075 35.640 147.485 ;
        RECT 34.730 146.905 35.060 147.025 ;
        RECT 35.810 146.905 35.980 147.665 ;
        RECT 34.730 146.735 35.980 146.905 ;
        RECT 36.150 147.845 37.520 148.095 ;
        RECT 36.150 147.075 36.340 147.845 ;
        RECT 37.270 147.585 37.520 147.845 ;
        RECT 36.510 147.415 36.760 147.575 ;
        RECT 37.690 147.415 37.860 148.260 ;
        RECT 38.755 147.975 38.925 148.475 ;
        RECT 39.095 148.145 39.425 148.645 ;
        RECT 38.030 147.585 38.530 147.965 ;
        RECT 38.755 147.805 39.450 147.975 ;
        RECT 36.510 147.245 37.860 147.415 ;
        RECT 37.440 147.205 37.860 147.245 ;
        RECT 36.150 146.735 36.570 147.075 ;
        RECT 36.860 146.745 37.270 147.075 ;
        RECT 34.390 146.315 35.240 146.485 ;
        RECT 35.800 146.095 36.120 146.555 ;
        RECT 36.320 146.305 36.570 146.735 ;
        RECT 36.860 146.095 37.270 146.535 ;
        RECT 37.440 146.475 37.610 147.205 ;
        RECT 37.780 146.655 38.130 147.025 ;
        RECT 38.310 146.715 38.530 147.585 ;
        RECT 38.700 147.015 39.110 147.635 ;
        RECT 39.280 146.835 39.450 147.805 ;
        RECT 38.755 146.645 39.450 146.835 ;
        RECT 37.440 146.275 38.455 146.475 ;
        RECT 38.755 146.315 38.925 146.645 ;
        RECT 39.095 146.095 39.425 146.475 ;
        RECT 39.640 146.355 39.865 148.475 ;
        RECT 40.035 148.145 40.365 148.645 ;
        RECT 40.535 147.975 40.705 148.475 ;
        RECT 40.040 147.805 40.705 147.975 ;
        RECT 40.040 146.815 40.270 147.805 ;
        RECT 40.440 146.985 40.790 147.635 ;
        RECT 40.965 147.555 42.635 148.645 ;
        RECT 40.965 147.035 41.715 147.555 ;
        RECT 42.810 147.505 43.145 148.475 ;
        RECT 43.315 147.505 43.485 148.645 ;
        RECT 43.655 148.305 45.685 148.475 ;
        RECT 41.885 146.865 42.635 147.385 ;
        RECT 40.040 146.645 40.705 146.815 ;
        RECT 40.035 146.095 40.365 146.475 ;
        RECT 40.535 146.355 40.705 146.645 ;
        RECT 40.965 146.095 42.635 146.865 ;
        RECT 42.810 146.835 42.980 147.505 ;
        RECT 43.655 147.335 43.825 148.305 ;
        RECT 43.150 147.005 43.405 147.335 ;
        RECT 43.630 147.005 43.825 147.335 ;
        RECT 43.995 147.965 45.120 148.135 ;
        RECT 43.235 146.835 43.405 147.005 ;
        RECT 43.995 146.835 44.165 147.965 ;
        RECT 42.810 146.265 43.065 146.835 ;
        RECT 43.235 146.665 44.165 146.835 ;
        RECT 44.335 147.625 45.345 147.795 ;
        RECT 44.335 146.825 44.505 147.625 ;
        RECT 44.710 146.945 44.985 147.425 ;
        RECT 44.705 146.775 44.985 146.945 ;
        RECT 43.990 146.630 44.165 146.665 ;
        RECT 43.235 146.095 43.565 146.495 ;
        RECT 43.990 146.265 44.520 146.630 ;
        RECT 44.710 146.265 44.985 146.775 ;
        RECT 45.155 146.265 45.345 147.625 ;
        RECT 45.515 147.640 45.685 148.305 ;
        RECT 45.855 147.885 46.025 148.645 ;
        RECT 46.260 147.885 46.775 148.295 ;
        RECT 45.515 147.450 46.265 147.640 ;
        RECT 46.435 147.075 46.775 147.885 ;
        RECT 45.545 146.905 46.775 147.075 ;
        RECT 46.945 147.925 47.405 148.475 ;
        RECT 47.595 147.925 47.925 148.645 ;
        RECT 45.525 146.095 46.035 146.630 ;
        RECT 46.255 146.300 46.500 146.905 ;
        RECT 46.945 146.555 47.195 147.925 ;
        RECT 48.125 147.755 48.425 148.305 ;
        RECT 48.595 147.975 48.875 148.645 ;
        RECT 47.485 147.585 48.425 147.755 ;
        RECT 47.485 147.335 47.655 147.585 ;
        RECT 48.795 147.335 49.060 147.695 ;
        RECT 50.165 147.480 50.455 148.645 ;
        RECT 51.145 147.505 51.355 148.645 ;
        RECT 51.525 147.495 51.855 148.475 ;
        RECT 52.025 147.505 52.255 148.645 ;
        RECT 52.465 147.505 52.735 148.475 ;
        RECT 52.945 147.845 53.225 148.645 ;
        RECT 53.395 148.135 55.050 148.425 ;
        RECT 53.460 147.795 55.050 147.965 ;
        RECT 55.225 147.810 55.610 148.645 ;
        RECT 53.460 147.675 53.630 147.795 ;
        RECT 52.905 147.505 53.630 147.675 ;
        RECT 47.365 147.005 47.655 147.335 ;
        RECT 47.825 147.085 48.165 147.335 ;
        RECT 48.385 147.085 49.060 147.335 ;
        RECT 47.485 146.915 47.655 147.005 ;
        RECT 47.485 146.725 48.875 146.915 ;
        RECT 46.945 146.265 47.505 146.555 ;
        RECT 47.675 146.095 47.925 146.555 ;
        RECT 48.545 146.365 48.875 146.725 ;
        RECT 50.165 146.095 50.455 146.820 ;
        RECT 51.145 146.095 51.355 146.915 ;
        RECT 51.525 146.895 51.775 147.495 ;
        RECT 51.945 147.085 52.275 147.335 ;
        RECT 51.525 146.265 51.855 146.895 ;
        RECT 52.025 146.095 52.255 146.915 ;
        RECT 52.465 146.770 52.635 147.505 ;
        RECT 52.905 147.335 53.075 147.505 ;
        RECT 53.820 147.455 54.535 147.625 ;
        RECT 54.730 147.505 55.050 147.795 ;
        RECT 55.780 147.640 56.040 148.445 ;
        RECT 56.210 147.810 56.470 148.645 ;
        RECT 56.640 147.640 56.895 148.445 ;
        RECT 57.070 147.810 57.330 148.645 ;
        RECT 57.500 147.640 57.755 148.445 ;
        RECT 57.930 147.810 58.275 148.645 ;
        RECT 58.560 148.015 58.845 148.475 ;
        RECT 59.015 148.185 59.285 148.645 ;
        RECT 58.560 147.795 59.515 148.015 ;
        RECT 55.225 147.470 58.255 147.640 ;
        RECT 52.805 147.005 53.075 147.335 ;
        RECT 53.245 147.005 53.650 147.335 ;
        RECT 53.820 147.005 54.530 147.455 ;
        RECT 52.905 146.835 53.075 147.005 ;
        RECT 52.465 146.425 52.735 146.770 ;
        RECT 52.905 146.665 54.515 146.835 ;
        RECT 54.700 146.765 55.050 147.335 ;
        RECT 55.225 146.905 55.525 147.470 ;
        RECT 55.700 147.075 57.915 147.300 ;
        RECT 58.085 146.905 58.255 147.470 ;
        RECT 58.445 147.065 59.135 147.625 ;
        RECT 55.225 146.735 58.255 146.905 ;
        RECT 59.305 146.895 59.515 147.795 ;
        RECT 52.925 146.095 53.305 146.495 ;
        RECT 53.475 146.315 53.645 146.665 ;
        RECT 53.815 146.095 54.145 146.495 ;
        RECT 54.345 146.315 54.515 146.665 ;
        RECT 54.715 146.095 55.045 146.595 ;
        RECT 55.745 146.095 56.045 146.565 ;
        RECT 56.215 146.290 56.470 146.735 ;
        RECT 56.640 146.095 56.900 146.565 ;
        RECT 57.070 146.290 57.330 146.735 ;
        RECT 58.560 146.725 59.515 146.895 ;
        RECT 59.685 147.625 60.085 148.475 ;
        RECT 60.275 148.015 60.555 148.475 ;
        RECT 61.075 148.185 61.400 148.645 ;
        RECT 60.275 147.795 61.400 148.015 ;
        RECT 59.685 147.065 60.780 147.625 ;
        RECT 60.950 147.335 61.400 147.795 ;
        RECT 61.570 147.505 61.955 148.475 ;
        RECT 57.500 146.095 57.795 146.565 ;
        RECT 58.560 146.265 58.845 146.725 ;
        RECT 59.015 146.095 59.285 146.555 ;
        RECT 59.685 146.265 60.085 147.065 ;
        RECT 60.950 147.005 61.505 147.335 ;
        RECT 60.950 146.895 61.400 147.005 ;
        RECT 60.275 146.725 61.400 146.895 ;
        RECT 61.675 146.835 61.955 147.505 ;
        RECT 62.125 147.555 64.715 148.645 ;
        RECT 65.000 148.015 65.285 148.475 ;
        RECT 65.455 148.185 65.725 148.645 ;
        RECT 65.000 147.795 65.955 148.015 ;
        RECT 62.125 147.035 63.335 147.555 ;
        RECT 63.505 146.865 64.715 147.385 ;
        RECT 64.885 147.065 65.575 147.625 ;
        RECT 65.745 146.895 65.955 147.795 ;
        RECT 60.275 146.265 60.555 146.725 ;
        RECT 61.075 146.095 61.400 146.555 ;
        RECT 61.570 146.265 61.955 146.835 ;
        RECT 62.125 146.095 64.715 146.865 ;
        RECT 65.000 146.725 65.955 146.895 ;
        RECT 66.125 147.625 66.525 148.475 ;
        RECT 66.715 148.015 66.995 148.475 ;
        RECT 67.515 148.185 67.840 148.645 ;
        RECT 66.715 147.795 67.840 148.015 ;
        RECT 66.125 147.065 67.220 147.625 ;
        RECT 67.390 147.335 67.840 147.795 ;
        RECT 68.010 147.505 68.395 148.475 ;
        RECT 65.000 146.265 65.285 146.725 ;
        RECT 65.455 146.095 65.725 146.555 ;
        RECT 66.125 146.265 66.525 147.065 ;
        RECT 67.390 147.005 67.945 147.335 ;
        RECT 67.390 146.895 67.840 147.005 ;
        RECT 66.715 146.725 67.840 146.895 ;
        RECT 68.115 146.835 68.395 147.505 ;
        RECT 69.025 147.555 70.695 148.645 ;
        RECT 70.865 147.885 71.380 148.295 ;
        RECT 71.615 147.885 71.785 148.645 ;
        RECT 71.955 148.305 73.985 148.475 ;
        RECT 69.025 147.035 69.775 147.555 ;
        RECT 69.945 146.865 70.695 147.385 ;
        RECT 70.865 147.075 71.205 147.885 ;
        RECT 71.955 147.640 72.125 148.305 ;
        RECT 72.520 147.965 73.645 148.135 ;
        RECT 71.375 147.450 72.125 147.640 ;
        RECT 72.295 147.625 73.305 147.795 ;
        RECT 70.865 146.905 72.095 147.075 ;
        RECT 66.715 146.265 66.995 146.725 ;
        RECT 67.515 146.095 67.840 146.555 ;
        RECT 68.010 146.265 68.395 146.835 ;
        RECT 69.025 146.095 70.695 146.865 ;
        RECT 71.140 146.300 71.385 146.905 ;
        RECT 71.605 146.095 72.115 146.630 ;
        RECT 72.295 146.265 72.485 147.625 ;
        RECT 72.655 147.285 72.930 147.425 ;
        RECT 72.655 147.115 72.935 147.285 ;
        RECT 72.655 146.265 72.930 147.115 ;
        RECT 73.135 146.825 73.305 147.625 ;
        RECT 73.475 146.835 73.645 147.965 ;
        RECT 73.815 147.335 73.985 148.305 ;
        RECT 74.155 147.505 74.325 148.645 ;
        RECT 74.495 147.505 74.830 148.475 ;
        RECT 73.815 147.005 74.010 147.335 ;
        RECT 74.235 147.005 74.490 147.335 ;
        RECT 74.235 146.835 74.405 147.005 ;
        RECT 74.660 146.835 74.830 147.505 ;
        RECT 75.925 147.480 76.215 148.645 ;
        RECT 77.305 147.555 80.815 148.645 ;
        RECT 80.990 148.210 86.335 148.645 ;
        RECT 77.305 147.035 78.995 147.555 ;
        RECT 79.165 146.865 80.815 147.385 ;
        RECT 82.580 146.960 82.930 148.210 ;
        RECT 86.880 147.665 87.135 148.335 ;
        RECT 87.315 147.845 87.600 148.645 ;
        RECT 87.780 147.925 88.110 148.435 ;
        RECT 73.475 146.665 74.405 146.835 ;
        RECT 73.475 146.630 73.650 146.665 ;
        RECT 73.120 146.265 73.650 146.630 ;
        RECT 74.075 146.095 74.405 146.495 ;
        RECT 74.575 146.265 74.830 146.835 ;
        RECT 75.925 146.095 76.215 146.820 ;
        RECT 77.305 146.095 80.815 146.865 ;
        RECT 84.410 146.640 84.750 147.470 ;
        RECT 86.880 146.805 87.060 147.665 ;
        RECT 87.780 147.335 88.030 147.925 ;
        RECT 88.380 147.775 88.550 148.385 ;
        RECT 88.720 147.955 89.050 148.645 ;
        RECT 89.280 148.095 89.520 148.385 ;
        RECT 89.720 148.265 90.140 148.645 ;
        RECT 90.320 148.175 90.950 148.425 ;
        RECT 91.420 148.265 91.750 148.645 ;
        RECT 90.320 148.095 90.490 148.175 ;
        RECT 91.920 148.095 92.090 148.385 ;
        RECT 92.270 148.265 92.650 148.645 ;
        RECT 92.890 148.260 93.720 148.430 ;
        RECT 89.280 147.925 90.490 148.095 ;
        RECT 87.230 147.005 88.030 147.335 ;
        RECT 80.990 146.095 86.335 146.640 ;
        RECT 86.880 146.605 87.135 146.805 ;
        RECT 86.795 146.435 87.135 146.605 ;
        RECT 86.880 146.275 87.135 146.435 ;
        RECT 87.315 146.095 87.600 146.555 ;
        RECT 87.780 146.355 88.030 147.005 ;
        RECT 88.230 147.755 88.550 147.775 ;
        RECT 88.230 147.585 90.150 147.755 ;
        RECT 88.230 146.690 88.420 147.585 ;
        RECT 90.320 147.415 90.490 147.925 ;
        RECT 90.660 147.665 91.180 147.975 ;
        RECT 88.590 147.245 90.490 147.415 ;
        RECT 88.590 147.185 88.920 147.245 ;
        RECT 89.070 147.015 89.400 147.075 ;
        RECT 88.740 146.745 89.400 147.015 ;
        RECT 88.230 146.360 88.550 146.690 ;
        RECT 88.730 146.095 89.390 146.575 ;
        RECT 89.590 146.485 89.760 147.245 ;
        RECT 90.660 147.075 90.840 147.485 ;
        RECT 89.930 146.905 90.260 147.025 ;
        RECT 91.010 146.905 91.180 147.665 ;
        RECT 89.930 146.735 91.180 146.905 ;
        RECT 91.350 147.845 92.720 148.095 ;
        RECT 91.350 147.075 91.540 147.845 ;
        RECT 92.470 147.585 92.720 147.845 ;
        RECT 91.710 147.415 91.960 147.575 ;
        RECT 92.890 147.415 93.060 148.260 ;
        RECT 93.955 147.975 94.125 148.475 ;
        RECT 94.295 148.145 94.625 148.645 ;
        RECT 93.230 147.585 93.730 147.965 ;
        RECT 93.955 147.805 94.650 147.975 ;
        RECT 91.710 147.245 93.060 147.415 ;
        RECT 92.640 147.205 93.060 147.245 ;
        RECT 91.350 146.735 91.770 147.075 ;
        RECT 92.060 146.745 92.470 147.075 ;
        RECT 89.590 146.315 90.440 146.485 ;
        RECT 91.000 146.095 91.320 146.555 ;
        RECT 91.520 146.305 91.770 146.735 ;
        RECT 92.060 146.095 92.470 146.535 ;
        RECT 92.640 146.475 92.810 147.205 ;
        RECT 92.980 146.655 93.330 147.025 ;
        RECT 93.510 146.715 93.730 147.585 ;
        RECT 93.900 147.015 94.310 147.635 ;
        RECT 94.480 146.835 94.650 147.805 ;
        RECT 93.955 146.645 94.650 146.835 ;
        RECT 92.640 146.275 93.655 146.475 ;
        RECT 93.955 146.315 94.125 146.645 ;
        RECT 94.295 146.095 94.625 146.475 ;
        RECT 94.840 146.355 95.065 148.475 ;
        RECT 95.235 148.145 95.565 148.645 ;
        RECT 95.735 147.975 95.905 148.475 ;
        RECT 95.240 147.805 95.905 147.975 ;
        RECT 95.240 146.815 95.470 147.805 ;
        RECT 95.640 146.985 95.990 147.635 ;
        RECT 96.165 147.555 97.375 148.645 ;
        RECT 96.165 147.015 96.685 147.555 ;
        RECT 97.585 147.505 97.815 148.645 ;
        RECT 97.985 147.495 98.315 148.475 ;
        RECT 98.485 147.505 98.695 148.645 ;
        RECT 98.930 148.135 100.585 148.425 ;
        RECT 98.930 147.795 100.520 147.965 ;
        RECT 100.755 147.845 101.035 148.645 ;
        RECT 98.930 147.505 99.250 147.795 ;
        RECT 100.350 147.675 100.520 147.795 ;
        RECT 96.855 146.845 97.375 147.385 ;
        RECT 97.565 147.085 97.895 147.335 ;
        RECT 95.240 146.645 95.905 146.815 ;
        RECT 95.235 146.095 95.565 146.475 ;
        RECT 95.735 146.355 95.905 146.645 ;
        RECT 96.165 146.095 97.375 146.845 ;
        RECT 97.585 146.095 97.815 146.915 ;
        RECT 98.065 146.895 98.315 147.495 ;
        RECT 97.985 146.265 98.315 146.895 ;
        RECT 98.485 146.095 98.695 146.915 ;
        RECT 98.930 146.765 99.280 147.335 ;
        RECT 99.450 147.005 100.160 147.625 ;
        RECT 100.350 147.505 101.075 147.675 ;
        RECT 101.245 147.505 101.515 148.475 ;
        RECT 100.905 147.335 101.075 147.505 ;
        RECT 100.330 147.005 100.735 147.335 ;
        RECT 100.905 147.005 101.175 147.335 ;
        RECT 100.905 146.835 101.075 147.005 ;
        RECT 99.465 146.665 101.075 146.835 ;
        RECT 101.345 146.770 101.515 147.505 ;
        RECT 101.685 147.480 101.975 148.645 ;
        RECT 103.065 147.885 103.580 148.295 ;
        RECT 103.815 147.885 103.985 148.645 ;
        RECT 104.155 148.305 106.185 148.475 ;
        RECT 103.065 147.075 103.405 147.885 ;
        RECT 104.155 147.640 104.325 148.305 ;
        RECT 104.720 147.965 105.845 148.135 ;
        RECT 103.575 147.450 104.325 147.640 ;
        RECT 104.495 147.625 105.505 147.795 ;
        RECT 103.065 146.905 104.295 147.075 ;
        RECT 98.935 146.095 99.265 146.595 ;
        RECT 99.465 146.315 99.635 146.665 ;
        RECT 99.835 146.095 100.165 146.495 ;
        RECT 100.335 146.315 100.505 146.665 ;
        RECT 100.675 146.095 101.055 146.495 ;
        RECT 101.245 146.425 101.515 146.770 ;
        RECT 101.685 146.095 101.975 146.820 ;
        RECT 103.340 146.300 103.585 146.905 ;
        RECT 103.805 146.095 104.315 146.630 ;
        RECT 104.495 146.265 104.685 147.625 ;
        RECT 104.855 146.945 105.130 147.425 ;
        RECT 104.855 146.775 105.135 146.945 ;
        RECT 105.335 146.825 105.505 147.625 ;
        RECT 105.675 146.835 105.845 147.965 ;
        RECT 106.015 147.335 106.185 148.305 ;
        RECT 106.355 147.505 106.525 148.645 ;
        RECT 106.695 147.505 107.030 148.475 ;
        RECT 107.210 148.135 108.865 148.425 ;
        RECT 107.210 147.795 108.800 147.965 ;
        RECT 109.035 147.845 109.315 148.645 ;
        RECT 107.210 147.505 107.530 147.795 ;
        RECT 108.630 147.675 108.800 147.795 ;
        RECT 106.015 147.005 106.210 147.335 ;
        RECT 106.435 147.005 106.690 147.335 ;
        RECT 106.435 146.835 106.605 147.005 ;
        RECT 106.860 146.835 107.030 147.505 ;
        RECT 104.855 146.265 105.130 146.775 ;
        RECT 105.675 146.665 106.605 146.835 ;
        RECT 105.675 146.630 105.850 146.665 ;
        RECT 105.320 146.265 105.850 146.630 ;
        RECT 106.275 146.095 106.605 146.495 ;
        RECT 106.775 146.265 107.030 146.835 ;
        RECT 107.210 146.765 107.560 147.335 ;
        RECT 107.730 147.005 108.440 147.625 ;
        RECT 108.630 147.505 109.355 147.675 ;
        RECT 109.525 147.505 109.795 148.475 ;
        RECT 109.185 147.335 109.355 147.505 ;
        RECT 108.610 147.005 109.015 147.335 ;
        RECT 109.185 147.005 109.455 147.335 ;
        RECT 109.185 146.835 109.355 147.005 ;
        RECT 107.745 146.665 109.355 146.835 ;
        RECT 109.625 146.770 109.795 147.505 ;
        RECT 107.215 146.095 107.545 146.595 ;
        RECT 107.745 146.315 107.915 146.665 ;
        RECT 108.115 146.095 108.445 146.495 ;
        RECT 108.615 146.315 108.785 146.665 ;
        RECT 108.955 146.095 109.335 146.495 ;
        RECT 109.525 146.425 109.795 146.770 ;
        RECT 109.965 147.505 110.235 148.475 ;
        RECT 110.445 147.845 110.725 148.645 ;
        RECT 110.895 148.135 112.550 148.425 ;
        RECT 110.960 147.795 112.550 147.965 ;
        RECT 110.960 147.675 111.130 147.795 ;
        RECT 110.405 147.505 111.130 147.675 ;
        RECT 109.965 146.770 110.135 147.505 ;
        RECT 110.405 147.335 110.575 147.505 ;
        RECT 111.320 147.455 112.035 147.625 ;
        RECT 112.230 147.505 112.550 147.795 ;
        RECT 114.020 147.665 114.275 148.335 ;
        RECT 114.455 147.845 114.740 148.645 ;
        RECT 114.920 147.925 115.250 148.435 ;
        RECT 110.305 147.005 110.575 147.335 ;
        RECT 110.745 147.005 111.150 147.335 ;
        RECT 111.320 147.005 112.030 147.455 ;
        RECT 110.405 146.835 110.575 147.005 ;
        RECT 109.965 146.425 110.235 146.770 ;
        RECT 110.405 146.665 112.015 146.835 ;
        RECT 112.200 146.765 112.550 147.335 ;
        RECT 114.020 146.805 114.200 147.665 ;
        RECT 114.920 147.335 115.170 147.925 ;
        RECT 115.520 147.775 115.690 148.385 ;
        RECT 115.860 147.955 116.190 148.645 ;
        RECT 116.420 148.095 116.660 148.385 ;
        RECT 116.860 148.265 117.280 148.645 ;
        RECT 117.460 148.175 118.090 148.425 ;
        RECT 118.560 148.265 118.890 148.645 ;
        RECT 117.460 148.095 117.630 148.175 ;
        RECT 119.060 148.095 119.230 148.385 ;
        RECT 119.410 148.265 119.790 148.645 ;
        RECT 120.030 148.260 120.860 148.430 ;
        RECT 116.420 147.925 117.630 148.095 ;
        RECT 114.370 147.005 115.170 147.335 ;
        RECT 110.425 146.095 110.805 146.495 ;
        RECT 110.975 146.315 111.145 146.665 ;
        RECT 111.315 146.095 111.645 146.495 ;
        RECT 111.845 146.315 112.015 146.665 ;
        RECT 114.020 146.605 114.275 146.805 ;
        RECT 112.215 146.095 112.545 146.595 ;
        RECT 113.935 146.435 114.275 146.605 ;
        RECT 114.020 146.275 114.275 146.435 ;
        RECT 114.455 146.095 114.740 146.555 ;
        RECT 114.920 146.355 115.170 147.005 ;
        RECT 115.370 147.755 115.690 147.775 ;
        RECT 115.370 147.585 117.290 147.755 ;
        RECT 115.370 146.690 115.560 147.585 ;
        RECT 117.460 147.415 117.630 147.925 ;
        RECT 117.800 147.665 118.320 147.975 ;
        RECT 115.730 147.245 117.630 147.415 ;
        RECT 115.730 147.185 116.060 147.245 ;
        RECT 116.210 147.015 116.540 147.075 ;
        RECT 115.880 146.745 116.540 147.015 ;
        RECT 115.370 146.360 115.690 146.690 ;
        RECT 115.870 146.095 116.530 146.575 ;
        RECT 116.730 146.485 116.900 147.245 ;
        RECT 117.800 147.075 117.980 147.485 ;
        RECT 117.070 146.905 117.400 147.025 ;
        RECT 118.150 146.905 118.320 147.665 ;
        RECT 117.070 146.735 118.320 146.905 ;
        RECT 118.490 147.845 119.860 148.095 ;
        RECT 118.490 147.075 118.680 147.845 ;
        RECT 119.610 147.585 119.860 147.845 ;
        RECT 118.850 147.415 119.100 147.575 ;
        RECT 120.030 147.415 120.200 148.260 ;
        RECT 121.095 147.975 121.265 148.475 ;
        RECT 121.435 148.145 121.765 148.645 ;
        RECT 120.370 147.585 120.870 147.965 ;
        RECT 121.095 147.805 121.790 147.975 ;
        RECT 118.850 147.245 120.200 147.415 ;
        RECT 119.780 147.205 120.200 147.245 ;
        RECT 118.490 146.735 118.910 147.075 ;
        RECT 119.200 146.745 119.610 147.075 ;
        RECT 116.730 146.315 117.580 146.485 ;
        RECT 118.140 146.095 118.460 146.555 ;
        RECT 118.660 146.305 118.910 146.735 ;
        RECT 119.200 146.095 119.610 146.535 ;
        RECT 119.780 146.475 119.950 147.205 ;
        RECT 120.120 146.655 120.470 147.025 ;
        RECT 120.650 146.715 120.870 147.585 ;
        RECT 121.040 147.015 121.450 147.635 ;
        RECT 121.620 146.835 121.790 147.805 ;
        RECT 121.095 146.645 121.790 146.835 ;
        RECT 119.780 146.275 120.795 146.475 ;
        RECT 121.095 146.315 121.265 146.645 ;
        RECT 121.435 146.095 121.765 146.475 ;
        RECT 121.980 146.355 122.205 148.475 ;
        RECT 122.375 148.145 122.705 148.645 ;
        RECT 122.875 147.975 123.045 148.475 ;
        RECT 122.380 147.805 123.045 147.975 ;
        RECT 122.380 146.815 122.610 147.805 ;
        RECT 123.395 147.715 123.565 148.475 ;
        RECT 123.745 147.885 124.075 148.645 ;
        RECT 122.780 146.985 123.130 147.635 ;
        RECT 123.395 147.545 124.060 147.715 ;
        RECT 124.245 147.570 124.515 148.475 ;
        RECT 123.890 147.400 124.060 147.545 ;
        RECT 123.325 146.995 123.655 147.365 ;
        RECT 123.890 147.070 124.175 147.400 ;
        RECT 123.890 146.815 124.060 147.070 ;
        RECT 122.380 146.645 123.045 146.815 ;
        RECT 122.375 146.095 122.705 146.475 ;
        RECT 122.875 146.355 123.045 146.645 ;
        RECT 123.395 146.645 124.060 146.815 ;
        RECT 124.345 146.770 124.515 147.570 ;
        RECT 124.685 147.555 126.355 148.645 ;
        RECT 126.525 147.555 127.735 148.645 ;
        RECT 124.685 147.035 125.435 147.555 ;
        RECT 125.605 146.865 126.355 147.385 ;
        RECT 126.525 147.015 127.045 147.555 ;
        RECT 123.395 146.265 123.565 146.645 ;
        RECT 123.745 146.095 124.075 146.475 ;
        RECT 124.255 146.265 124.515 146.770 ;
        RECT 124.685 146.095 126.355 146.865 ;
        RECT 127.215 146.845 127.735 147.385 ;
        RECT 126.525 146.095 127.735 146.845 ;
        RECT 29.840 145.925 127.820 146.095 ;
        RECT 29.925 145.175 31.135 145.925 ;
        RECT 29.925 144.635 30.445 145.175 ;
        RECT 31.825 145.105 32.035 145.925 ;
        RECT 32.205 145.125 32.535 145.755 ;
        RECT 30.615 144.465 31.135 145.005 ;
        RECT 32.205 144.525 32.455 145.125 ;
        RECT 32.705 145.105 32.935 145.925 ;
        RECT 33.420 145.115 33.665 145.720 ;
        RECT 33.885 145.390 34.395 145.925 ;
        RECT 33.145 144.945 34.375 145.115 ;
        RECT 32.625 144.685 32.955 144.935 ;
        RECT 29.925 143.375 31.135 144.465 ;
        RECT 31.825 143.375 32.035 144.515 ;
        RECT 32.205 143.545 32.535 144.525 ;
        RECT 32.705 143.375 32.935 144.515 ;
        RECT 33.145 144.135 33.485 144.945 ;
        RECT 33.655 144.380 34.405 144.570 ;
        RECT 33.145 143.725 33.660 144.135 ;
        RECT 33.895 143.375 34.065 144.135 ;
        RECT 34.235 143.715 34.405 144.380 ;
        RECT 34.575 144.395 34.765 145.755 ;
        RECT 34.935 145.585 35.210 145.755 ;
        RECT 34.935 145.415 35.215 145.585 ;
        RECT 34.935 144.595 35.210 145.415 ;
        RECT 35.400 145.390 35.930 145.755 ;
        RECT 36.355 145.525 36.685 145.925 ;
        RECT 35.755 145.355 35.930 145.390 ;
        RECT 35.415 144.395 35.585 145.195 ;
        RECT 34.575 144.225 35.585 144.395 ;
        RECT 35.755 145.185 36.685 145.355 ;
        RECT 36.855 145.185 37.110 145.755 ;
        RECT 37.285 145.200 37.575 145.925 ;
        RECT 37.835 145.375 38.005 145.755 ;
        RECT 38.185 145.545 38.515 145.925 ;
        RECT 37.835 145.205 38.500 145.375 ;
        RECT 38.695 145.250 38.955 145.755 ;
        RECT 35.755 144.055 35.925 145.185 ;
        RECT 36.515 145.015 36.685 145.185 ;
        RECT 34.800 143.885 35.925 144.055 ;
        RECT 36.095 144.685 36.290 145.015 ;
        RECT 36.515 144.685 36.770 145.015 ;
        RECT 36.095 143.715 36.265 144.685 ;
        RECT 36.940 144.515 37.110 145.185 ;
        RECT 37.765 144.655 38.095 145.025 ;
        RECT 38.330 144.950 38.500 145.205 ;
        RECT 38.330 144.620 38.615 144.950 ;
        RECT 34.235 143.545 36.265 143.715 ;
        RECT 36.435 143.375 36.605 144.515 ;
        RECT 36.775 143.545 37.110 144.515 ;
        RECT 37.285 143.375 37.575 144.540 ;
        RECT 38.330 144.475 38.500 144.620 ;
        RECT 37.835 144.305 38.500 144.475 ;
        RECT 38.785 144.450 38.955 145.250 ;
        RECT 39.125 145.155 42.635 145.925 ;
        RECT 42.810 145.380 48.155 145.925 ;
        RECT 48.330 145.380 53.675 145.925 ;
        RECT 53.935 145.445 54.235 145.925 ;
        RECT 37.835 143.545 38.005 144.305 ;
        RECT 38.185 143.375 38.515 144.135 ;
        RECT 38.685 143.545 38.955 144.450 ;
        RECT 39.125 144.465 40.815 144.985 ;
        RECT 40.985 144.635 42.635 145.155 ;
        RECT 39.125 143.375 42.635 144.465 ;
        RECT 44.400 143.810 44.750 145.060 ;
        RECT 46.230 144.550 46.570 145.380 ;
        RECT 49.920 143.810 50.270 145.060 ;
        RECT 51.750 144.550 52.090 145.380 ;
        RECT 54.405 145.275 54.665 145.730 ;
        RECT 54.835 145.445 55.095 145.925 ;
        RECT 55.275 145.275 55.535 145.730 ;
        RECT 55.705 145.445 55.955 145.925 ;
        RECT 56.135 145.275 56.395 145.730 ;
        RECT 56.565 145.445 56.815 145.925 ;
        RECT 56.995 145.275 57.255 145.730 ;
        RECT 57.425 145.445 57.670 145.925 ;
        RECT 57.840 145.275 58.115 145.730 ;
        RECT 58.285 145.445 58.530 145.925 ;
        RECT 58.700 145.275 58.960 145.730 ;
        RECT 59.130 145.445 59.390 145.925 ;
        RECT 59.560 145.275 59.820 145.730 ;
        RECT 59.990 145.445 60.250 145.925 ;
        RECT 60.420 145.275 60.680 145.730 ;
        RECT 60.850 145.365 61.110 145.925 ;
        RECT 53.935 145.105 60.680 145.275 ;
        RECT 53.935 144.515 55.100 145.105 ;
        RECT 61.280 144.935 61.530 145.745 ;
        RECT 61.710 145.400 61.970 145.925 ;
        RECT 62.140 144.935 62.390 145.745 ;
        RECT 62.570 145.415 62.875 145.925 ;
        RECT 55.270 144.685 62.390 144.935 ;
        RECT 62.560 144.685 62.875 145.245 ;
        RECT 63.045 145.200 63.335 145.925 ;
        RECT 63.965 145.425 64.225 145.755 ;
        RECT 64.395 145.565 64.725 145.925 ;
        RECT 64.980 145.545 66.280 145.755 ;
        RECT 63.965 145.415 64.195 145.425 ;
        RECT 53.935 144.290 60.680 144.515 ;
        RECT 42.810 143.375 48.155 143.810 ;
        RECT 48.330 143.375 53.675 143.810 ;
        RECT 53.935 143.375 54.205 144.120 ;
        RECT 54.375 143.550 54.665 144.290 ;
        RECT 55.275 144.275 60.680 144.290 ;
        RECT 54.835 143.380 55.090 144.105 ;
        RECT 55.275 143.550 55.535 144.275 ;
        RECT 55.705 143.380 55.950 144.105 ;
        RECT 56.135 143.550 56.395 144.275 ;
        RECT 56.565 143.380 56.810 144.105 ;
        RECT 56.995 143.550 57.255 144.275 ;
        RECT 57.425 143.380 57.670 144.105 ;
        RECT 57.840 143.550 58.100 144.275 ;
        RECT 58.270 143.380 58.530 144.105 ;
        RECT 58.700 143.550 58.960 144.275 ;
        RECT 59.130 143.380 59.390 144.105 ;
        RECT 59.560 143.550 59.820 144.275 ;
        RECT 59.990 143.380 60.250 144.105 ;
        RECT 60.420 143.550 60.680 144.275 ;
        RECT 60.850 143.380 61.110 144.175 ;
        RECT 61.280 143.550 61.530 144.685 ;
        RECT 54.835 143.375 61.110 143.380 ;
        RECT 61.710 143.375 61.970 144.185 ;
        RECT 62.145 143.545 62.390 144.685 ;
        RECT 62.570 143.375 62.865 144.185 ;
        RECT 63.045 143.375 63.335 144.540 ;
        RECT 63.965 144.225 64.135 145.415 ;
        RECT 64.980 145.395 65.150 145.545 ;
        RECT 64.395 145.270 65.150 145.395 ;
        RECT 64.305 145.225 65.150 145.270 ;
        RECT 64.305 145.105 64.575 145.225 ;
        RECT 64.305 144.530 64.475 145.105 ;
        RECT 64.705 144.665 65.115 144.970 ;
        RECT 65.405 144.935 65.615 145.335 ;
        RECT 65.285 144.725 65.615 144.935 ;
        RECT 65.860 144.935 66.080 145.335 ;
        RECT 66.555 145.160 67.010 145.925 ;
        RECT 67.185 145.125 67.525 145.755 ;
        RECT 67.695 145.125 67.945 145.925 ;
        RECT 68.135 145.275 68.465 145.755 ;
        RECT 68.635 145.465 68.860 145.925 ;
        RECT 69.030 145.275 69.360 145.755 ;
        RECT 65.860 144.725 66.335 144.935 ;
        RECT 66.525 144.735 67.015 144.935 ;
        RECT 64.305 144.495 64.505 144.530 ;
        RECT 65.835 144.495 67.010 144.555 ;
        RECT 64.305 144.385 67.010 144.495 ;
        RECT 64.365 144.325 66.165 144.385 ;
        RECT 65.835 144.295 66.165 144.325 ;
        RECT 63.965 143.545 64.225 144.225 ;
        RECT 64.395 143.375 64.645 144.155 ;
        RECT 64.895 144.125 65.730 144.135 ;
        RECT 66.320 144.125 66.505 144.215 ;
        RECT 64.895 143.925 66.505 144.125 ;
        RECT 64.895 143.545 65.145 143.925 ;
        RECT 66.275 143.885 66.505 143.925 ;
        RECT 66.755 143.765 67.010 144.385 ;
        RECT 65.315 143.375 65.670 143.755 ;
        RECT 66.675 143.545 67.010 143.765 ;
        RECT 67.185 144.515 67.360 145.125 ;
        RECT 68.135 145.105 69.360 145.275 ;
        RECT 69.990 145.145 70.490 145.755 ;
        RECT 71.325 145.155 74.835 145.925 ;
        RECT 75.095 145.375 75.265 145.755 ;
        RECT 75.445 145.545 75.775 145.925 ;
        RECT 75.095 145.205 75.760 145.375 ;
        RECT 75.955 145.250 76.215 145.755 ;
        RECT 76.390 145.525 76.725 145.925 ;
        RECT 76.895 145.355 77.100 145.755 ;
        RECT 77.310 145.445 77.585 145.925 ;
        RECT 77.795 145.425 78.055 145.755 ;
        RECT 67.530 144.765 68.225 144.935 ;
        RECT 68.055 144.515 68.225 144.765 ;
        RECT 68.400 144.735 68.820 144.935 ;
        RECT 68.990 144.735 69.320 144.935 ;
        RECT 69.490 144.735 69.820 144.935 ;
        RECT 69.990 144.515 70.160 145.145 ;
        RECT 70.345 144.685 70.695 144.935 ;
        RECT 67.185 143.545 67.525 144.515 ;
        RECT 67.695 143.375 67.865 144.515 ;
        RECT 68.055 144.345 70.490 144.515 ;
        RECT 68.135 143.375 68.385 144.175 ;
        RECT 69.030 143.545 69.360 144.345 ;
        RECT 69.660 143.375 69.990 144.175 ;
        RECT 70.160 143.545 70.490 144.345 ;
        RECT 71.325 144.465 73.015 144.985 ;
        RECT 73.185 144.635 74.835 145.155 ;
        RECT 75.025 144.655 75.355 145.025 ;
        RECT 75.590 144.950 75.760 145.205 ;
        RECT 75.590 144.620 75.875 144.950 ;
        RECT 75.590 144.475 75.760 144.620 ;
        RECT 71.325 143.375 74.835 144.465 ;
        RECT 75.095 144.305 75.760 144.475 ;
        RECT 76.045 144.450 76.215 145.250 ;
        RECT 75.095 143.545 75.265 144.305 ;
        RECT 75.445 143.375 75.775 144.135 ;
        RECT 75.945 143.545 76.215 144.450 ;
        RECT 76.415 145.185 77.100 145.355 ;
        RECT 76.415 144.155 76.755 145.185 ;
        RECT 76.925 144.515 77.175 145.015 ;
        RECT 77.355 144.685 77.715 145.265 ;
        RECT 77.885 144.515 78.055 145.425 ;
        RECT 76.925 144.345 78.055 144.515 ;
        RECT 76.415 143.980 77.080 144.155 ;
        RECT 76.390 143.375 76.725 143.800 ;
        RECT 76.895 143.575 77.080 143.980 ;
        RECT 77.285 143.375 77.615 144.155 ;
        RECT 77.785 143.575 78.055 144.345 ;
        RECT 78.225 145.250 78.495 145.595 ;
        RECT 78.685 145.525 79.065 145.925 ;
        RECT 79.235 145.355 79.405 145.705 ;
        RECT 79.575 145.525 79.905 145.925 ;
        RECT 80.105 145.355 80.275 145.705 ;
        RECT 80.475 145.425 80.805 145.925 ;
        RECT 78.225 144.515 78.395 145.250 ;
        RECT 78.665 145.185 80.275 145.355 ;
        RECT 78.665 145.015 78.835 145.185 ;
        RECT 78.565 144.685 78.835 145.015 ;
        RECT 79.005 144.685 79.410 145.015 ;
        RECT 78.665 144.515 78.835 144.685 ;
        RECT 79.580 144.565 80.290 145.015 ;
        RECT 80.460 144.685 80.810 145.255 ;
        RECT 80.985 145.125 81.325 145.755 ;
        RECT 81.495 145.125 81.745 145.925 ;
        RECT 81.935 145.275 82.265 145.755 ;
        RECT 82.435 145.465 82.660 145.925 ;
        RECT 82.830 145.275 83.160 145.755 ;
        RECT 80.985 145.075 81.215 145.125 ;
        RECT 81.935 145.105 83.160 145.275 ;
        RECT 83.790 145.145 84.290 145.755 ;
        RECT 78.225 143.545 78.495 144.515 ;
        RECT 78.665 144.345 79.390 144.515 ;
        RECT 79.580 144.395 80.295 144.565 ;
        RECT 80.985 144.515 81.160 145.075 ;
        RECT 81.330 144.765 82.025 144.935 ;
        RECT 81.855 144.515 82.025 144.765 ;
        RECT 82.200 144.735 82.620 144.935 ;
        RECT 82.790 144.735 83.120 144.935 ;
        RECT 83.290 144.735 83.620 144.935 ;
        RECT 83.790 144.515 83.960 145.145 ;
        RECT 84.940 145.115 85.185 145.720 ;
        RECT 85.405 145.390 85.915 145.925 ;
        RECT 84.665 144.945 85.895 145.115 ;
        RECT 84.145 144.685 84.495 144.935 ;
        RECT 79.220 144.225 79.390 144.345 ;
        RECT 80.490 144.225 80.810 144.515 ;
        RECT 78.705 143.375 78.985 144.175 ;
        RECT 79.220 144.055 80.810 144.225 ;
        RECT 79.155 143.595 80.810 143.885 ;
        RECT 80.985 143.545 81.325 144.515 ;
        RECT 81.495 143.375 81.665 144.515 ;
        RECT 81.855 144.345 84.290 144.515 ;
        RECT 81.935 143.375 82.185 144.175 ;
        RECT 82.830 143.545 83.160 144.345 ;
        RECT 83.460 143.375 83.790 144.175 ;
        RECT 83.960 143.545 84.290 144.345 ;
        RECT 84.665 144.135 85.005 144.945 ;
        RECT 85.175 144.380 85.925 144.570 ;
        RECT 84.665 143.725 85.180 144.135 ;
        RECT 85.415 143.375 85.585 144.135 ;
        RECT 85.755 143.715 85.925 144.380 ;
        RECT 86.095 144.395 86.285 145.755 ;
        RECT 86.455 144.905 86.730 145.755 ;
        RECT 86.920 145.390 87.450 145.755 ;
        RECT 87.875 145.525 88.205 145.925 ;
        RECT 87.275 145.355 87.450 145.390 ;
        RECT 86.455 144.735 86.735 144.905 ;
        RECT 86.455 144.595 86.730 144.735 ;
        RECT 86.935 144.395 87.105 145.195 ;
        RECT 86.095 144.225 87.105 144.395 ;
        RECT 87.275 145.185 88.205 145.355 ;
        RECT 88.375 145.185 88.630 145.755 ;
        RECT 88.805 145.200 89.095 145.925 ;
        RECT 87.275 144.055 87.445 145.185 ;
        RECT 88.035 145.015 88.205 145.185 ;
        RECT 86.320 143.885 87.445 144.055 ;
        RECT 87.615 144.685 87.810 145.015 ;
        RECT 88.035 144.685 88.290 145.015 ;
        RECT 87.615 143.715 87.785 144.685 ;
        RECT 88.460 144.515 88.630 145.185 ;
        RECT 89.540 145.115 89.785 145.720 ;
        RECT 90.005 145.390 90.515 145.925 ;
        RECT 89.265 144.945 90.495 145.115 ;
        RECT 85.755 143.545 87.785 143.715 ;
        RECT 87.955 143.375 88.125 144.515 ;
        RECT 88.295 143.545 88.630 144.515 ;
        RECT 88.805 143.375 89.095 144.540 ;
        RECT 89.265 144.135 89.605 144.945 ;
        RECT 89.775 144.380 90.525 144.570 ;
        RECT 89.265 143.725 89.780 144.135 ;
        RECT 90.015 143.375 90.185 144.135 ;
        RECT 90.355 143.715 90.525 144.380 ;
        RECT 90.695 144.395 90.885 145.755 ;
        RECT 91.055 145.585 91.330 145.755 ;
        RECT 91.055 145.415 91.335 145.585 ;
        RECT 91.055 144.595 91.330 145.415 ;
        RECT 91.520 145.390 92.050 145.755 ;
        RECT 92.475 145.525 92.805 145.925 ;
        RECT 91.875 145.355 92.050 145.390 ;
        RECT 91.535 144.395 91.705 145.195 ;
        RECT 90.695 144.225 91.705 144.395 ;
        RECT 91.875 145.185 92.805 145.355 ;
        RECT 92.975 145.185 93.230 145.755 ;
        RECT 93.405 145.415 93.710 145.925 ;
        RECT 91.875 144.055 92.045 145.185 ;
        RECT 92.635 145.015 92.805 145.185 ;
        RECT 90.920 143.885 92.045 144.055 ;
        RECT 92.215 144.685 92.410 145.015 ;
        RECT 92.635 144.685 92.890 145.015 ;
        RECT 92.215 143.715 92.385 144.685 ;
        RECT 93.060 144.515 93.230 145.185 ;
        RECT 93.405 144.685 93.720 145.245 ;
        RECT 93.890 144.935 94.140 145.745 ;
        RECT 94.310 145.400 94.570 145.925 ;
        RECT 94.750 144.935 95.000 145.745 ;
        RECT 95.170 145.365 95.430 145.925 ;
        RECT 95.600 145.275 95.860 145.730 ;
        RECT 96.030 145.445 96.290 145.925 ;
        RECT 96.460 145.275 96.720 145.730 ;
        RECT 96.890 145.445 97.150 145.925 ;
        RECT 97.320 145.275 97.580 145.730 ;
        RECT 97.750 145.445 97.995 145.925 ;
        RECT 98.165 145.275 98.440 145.730 ;
        RECT 98.610 145.445 98.855 145.925 ;
        RECT 99.025 145.275 99.285 145.730 ;
        RECT 99.465 145.445 99.715 145.925 ;
        RECT 99.885 145.275 100.145 145.730 ;
        RECT 100.325 145.445 100.575 145.925 ;
        RECT 100.745 145.275 101.005 145.730 ;
        RECT 101.185 145.445 101.445 145.925 ;
        RECT 101.615 145.275 101.875 145.730 ;
        RECT 102.045 145.445 102.345 145.925 ;
        RECT 95.600 145.245 102.345 145.275 ;
        RECT 95.600 145.105 102.375 145.245 ;
        RECT 103.065 145.155 104.735 145.925 ;
        RECT 101.180 145.075 102.375 145.105 ;
        RECT 93.890 144.685 101.010 144.935 ;
        RECT 90.355 143.545 92.385 143.715 ;
        RECT 92.555 143.375 92.725 144.515 ;
        RECT 92.895 143.545 93.230 144.515 ;
        RECT 93.415 143.375 93.710 144.185 ;
        RECT 93.890 143.545 94.135 144.685 ;
        RECT 94.310 143.375 94.570 144.185 ;
        RECT 94.750 143.550 95.000 144.685 ;
        RECT 101.180 144.515 102.345 145.075 ;
        RECT 95.600 144.290 102.345 144.515 ;
        RECT 103.065 144.465 103.815 144.985 ;
        RECT 103.985 144.635 104.735 145.155 ;
        RECT 104.905 145.250 105.165 145.755 ;
        RECT 105.345 145.545 105.675 145.925 ;
        RECT 105.855 145.375 106.025 145.755 ;
        RECT 95.600 144.275 101.005 144.290 ;
        RECT 95.170 143.380 95.430 144.175 ;
        RECT 95.600 143.550 95.860 144.275 ;
        RECT 96.030 143.380 96.290 144.105 ;
        RECT 96.460 143.550 96.720 144.275 ;
        RECT 96.890 143.380 97.150 144.105 ;
        RECT 97.320 143.550 97.580 144.275 ;
        RECT 97.750 143.380 98.010 144.105 ;
        RECT 98.180 143.550 98.440 144.275 ;
        RECT 98.610 143.380 98.855 144.105 ;
        RECT 99.025 143.550 99.285 144.275 ;
        RECT 99.470 143.380 99.715 144.105 ;
        RECT 99.885 143.550 100.145 144.275 ;
        RECT 100.330 143.380 100.575 144.105 ;
        RECT 100.745 143.550 101.005 144.275 ;
        RECT 101.190 143.380 101.445 144.105 ;
        RECT 101.615 143.550 101.905 144.290 ;
        RECT 95.170 143.375 101.445 143.380 ;
        RECT 102.075 143.375 102.345 144.120 ;
        RECT 103.065 143.375 104.735 144.465 ;
        RECT 104.905 144.450 105.075 145.250 ;
        RECT 105.360 145.205 106.025 145.375 ;
        RECT 105.360 144.950 105.530 145.205 ;
        RECT 106.285 145.155 108.875 145.925 ;
        RECT 109.050 145.380 114.395 145.925 ;
        RECT 105.245 144.620 105.530 144.950 ;
        RECT 105.765 144.655 106.095 145.025 ;
        RECT 105.360 144.475 105.530 144.620 ;
        RECT 104.905 143.545 105.175 144.450 ;
        RECT 105.360 144.305 106.025 144.475 ;
        RECT 105.345 143.375 105.675 144.135 ;
        RECT 105.855 143.545 106.025 144.305 ;
        RECT 106.285 144.465 107.495 144.985 ;
        RECT 107.665 144.635 108.875 145.155 ;
        RECT 106.285 143.375 108.875 144.465 ;
        RECT 110.640 143.810 110.990 145.060 ;
        RECT 112.470 144.550 112.810 145.380 ;
        RECT 114.565 145.200 114.855 145.925 ;
        RECT 115.300 145.115 115.545 145.720 ;
        RECT 115.765 145.390 116.275 145.925 ;
        RECT 115.025 144.945 116.255 145.115 ;
        RECT 109.050 143.375 114.395 143.810 ;
        RECT 114.565 143.375 114.855 144.540 ;
        RECT 115.025 144.135 115.365 144.945 ;
        RECT 115.535 144.380 116.285 144.570 ;
        RECT 115.025 143.725 115.540 144.135 ;
        RECT 115.775 143.375 115.945 144.135 ;
        RECT 116.115 143.715 116.285 144.380 ;
        RECT 116.455 144.395 116.645 145.755 ;
        RECT 116.815 145.585 117.090 145.755 ;
        RECT 116.815 145.415 117.095 145.585 ;
        RECT 116.815 144.595 117.090 145.415 ;
        RECT 117.280 145.390 117.810 145.755 ;
        RECT 118.235 145.525 118.565 145.925 ;
        RECT 117.635 145.355 117.810 145.390 ;
        RECT 117.295 144.395 117.465 145.195 ;
        RECT 116.455 144.225 117.465 144.395 ;
        RECT 117.635 145.185 118.565 145.355 ;
        RECT 118.735 145.185 118.990 145.755 ;
        RECT 119.715 145.375 119.885 145.755 ;
        RECT 120.065 145.545 120.395 145.925 ;
        RECT 119.715 145.205 120.380 145.375 ;
        RECT 120.575 145.250 120.835 145.755 ;
        RECT 121.010 145.380 126.355 145.925 ;
        RECT 117.635 144.055 117.805 145.185 ;
        RECT 118.395 145.015 118.565 145.185 ;
        RECT 116.680 143.885 117.805 144.055 ;
        RECT 117.975 144.685 118.170 145.015 ;
        RECT 118.395 144.685 118.650 145.015 ;
        RECT 117.975 143.715 118.145 144.685 ;
        RECT 118.820 144.515 118.990 145.185 ;
        RECT 119.645 144.655 119.975 145.025 ;
        RECT 120.210 144.950 120.380 145.205 ;
        RECT 116.115 143.545 118.145 143.715 ;
        RECT 118.315 143.375 118.485 144.515 ;
        RECT 118.655 143.545 118.990 144.515 ;
        RECT 120.210 144.620 120.495 144.950 ;
        RECT 120.210 144.475 120.380 144.620 ;
        RECT 119.715 144.305 120.380 144.475 ;
        RECT 120.665 144.450 120.835 145.250 ;
        RECT 119.715 143.545 119.885 144.305 ;
        RECT 120.065 143.375 120.395 144.135 ;
        RECT 120.565 143.545 120.835 144.450 ;
        RECT 122.600 143.810 122.950 145.060 ;
        RECT 124.430 144.550 124.770 145.380 ;
        RECT 126.525 145.175 127.735 145.925 ;
        RECT 126.525 144.465 127.045 145.005 ;
        RECT 127.215 144.635 127.735 145.175 ;
        RECT 121.010 143.375 126.355 143.810 ;
        RECT 126.525 143.375 127.735 144.465 ;
        RECT 29.840 143.205 127.820 143.375 ;
        RECT 29.925 142.115 31.135 143.205 ;
        RECT 32.600 142.225 32.855 142.895 ;
        RECT 33.035 142.405 33.320 143.205 ;
        RECT 33.500 142.485 33.830 142.995 ;
        RECT 32.600 142.185 32.780 142.225 ;
        RECT 29.925 141.405 30.445 141.945 ;
        RECT 30.615 141.575 31.135 142.115 ;
        RECT 32.515 142.015 32.780 142.185 ;
        RECT 29.925 140.655 31.135 141.405 ;
        RECT 32.600 141.365 32.780 142.015 ;
        RECT 33.500 141.895 33.750 142.485 ;
        RECT 34.100 142.335 34.270 142.945 ;
        RECT 34.440 142.515 34.770 143.205 ;
        RECT 35.000 142.655 35.240 142.945 ;
        RECT 35.440 142.825 35.860 143.205 ;
        RECT 36.040 142.735 36.670 142.985 ;
        RECT 37.140 142.825 37.470 143.205 ;
        RECT 36.040 142.655 36.210 142.735 ;
        RECT 37.640 142.655 37.810 142.945 ;
        RECT 37.990 142.825 38.370 143.205 ;
        RECT 38.610 142.820 39.440 142.990 ;
        RECT 35.000 142.485 36.210 142.655 ;
        RECT 32.950 141.565 33.750 141.895 ;
        RECT 32.600 140.835 32.855 141.365 ;
        RECT 33.035 140.655 33.320 141.115 ;
        RECT 33.500 140.915 33.750 141.565 ;
        RECT 33.950 142.315 34.270 142.335 ;
        RECT 33.950 142.145 35.870 142.315 ;
        RECT 33.950 141.250 34.140 142.145 ;
        RECT 36.040 141.975 36.210 142.485 ;
        RECT 36.380 142.225 36.900 142.535 ;
        RECT 34.310 141.805 36.210 141.975 ;
        RECT 34.310 141.745 34.640 141.805 ;
        RECT 34.790 141.575 35.120 141.635 ;
        RECT 34.460 141.305 35.120 141.575 ;
        RECT 33.950 140.920 34.270 141.250 ;
        RECT 34.450 140.655 35.110 141.135 ;
        RECT 35.310 141.045 35.480 141.805 ;
        RECT 36.380 141.635 36.560 142.045 ;
        RECT 35.650 141.465 35.980 141.585 ;
        RECT 36.730 141.465 36.900 142.225 ;
        RECT 35.650 141.295 36.900 141.465 ;
        RECT 37.070 142.405 38.440 142.655 ;
        RECT 37.070 141.635 37.260 142.405 ;
        RECT 38.190 142.145 38.440 142.405 ;
        RECT 37.430 141.975 37.680 142.135 ;
        RECT 38.610 141.975 38.780 142.820 ;
        RECT 39.675 142.535 39.845 143.035 ;
        RECT 40.015 142.705 40.345 143.205 ;
        RECT 38.950 142.145 39.450 142.525 ;
        RECT 39.675 142.365 40.370 142.535 ;
        RECT 37.430 141.805 38.780 141.975 ;
        RECT 38.360 141.765 38.780 141.805 ;
        RECT 37.070 141.295 37.490 141.635 ;
        RECT 37.780 141.305 38.190 141.635 ;
        RECT 35.310 140.875 36.160 141.045 ;
        RECT 36.720 140.655 37.040 141.115 ;
        RECT 37.240 140.865 37.490 141.295 ;
        RECT 37.780 140.655 38.190 141.095 ;
        RECT 38.360 141.035 38.530 141.765 ;
        RECT 38.700 141.215 39.050 141.585 ;
        RECT 39.230 141.275 39.450 142.145 ;
        RECT 39.620 141.575 40.030 142.195 ;
        RECT 40.200 141.395 40.370 142.365 ;
        RECT 39.675 141.205 40.370 141.395 ;
        RECT 38.360 140.835 39.375 141.035 ;
        RECT 39.675 140.875 39.845 141.205 ;
        RECT 40.015 140.655 40.345 141.035 ;
        RECT 40.560 140.915 40.785 143.035 ;
        RECT 40.955 142.705 41.285 143.205 ;
        RECT 41.455 142.535 41.625 143.035 ;
        RECT 40.960 142.365 41.625 142.535 ;
        RECT 40.960 141.375 41.190 142.365 ;
        RECT 41.360 141.545 41.710 142.195 ;
        RECT 41.885 142.115 44.475 143.205 ;
        RECT 41.885 141.595 43.095 142.115 ;
        RECT 44.685 142.065 44.915 143.205 ;
        RECT 45.085 142.055 45.415 143.035 ;
        RECT 45.585 142.065 45.795 143.205 ;
        RECT 46.030 142.065 46.365 143.035 ;
        RECT 46.535 142.065 46.705 143.205 ;
        RECT 46.875 142.865 48.905 143.035 ;
        RECT 43.265 141.425 44.475 141.945 ;
        RECT 44.665 141.645 44.995 141.895 ;
        RECT 40.960 141.205 41.625 141.375 ;
        RECT 40.955 140.655 41.285 141.035 ;
        RECT 41.455 140.915 41.625 141.205 ;
        RECT 41.885 140.655 44.475 141.425 ;
        RECT 44.685 140.655 44.915 141.475 ;
        RECT 45.165 141.455 45.415 142.055 ;
        RECT 45.085 140.825 45.415 141.455 ;
        RECT 45.585 140.655 45.795 141.475 ;
        RECT 46.030 141.395 46.200 142.065 ;
        RECT 46.875 141.895 47.045 142.865 ;
        RECT 46.370 141.565 46.625 141.895 ;
        RECT 46.850 141.565 47.045 141.895 ;
        RECT 47.215 142.525 48.340 142.695 ;
        RECT 46.455 141.395 46.625 141.565 ;
        RECT 47.215 141.395 47.385 142.525 ;
        RECT 46.030 140.825 46.285 141.395 ;
        RECT 46.455 141.225 47.385 141.395 ;
        RECT 47.555 142.185 48.565 142.355 ;
        RECT 47.555 141.385 47.725 142.185 ;
        RECT 47.210 141.190 47.385 141.225 ;
        RECT 46.455 140.655 46.785 141.055 ;
        RECT 47.210 140.825 47.740 141.190 ;
        RECT 47.930 141.165 48.205 141.985 ;
        RECT 47.925 140.995 48.205 141.165 ;
        RECT 47.930 140.825 48.205 140.995 ;
        RECT 48.375 140.825 48.565 142.185 ;
        RECT 48.735 142.200 48.905 142.865 ;
        RECT 49.075 142.445 49.245 143.205 ;
        RECT 49.480 142.445 49.995 142.855 ;
        RECT 48.735 142.010 49.485 142.200 ;
        RECT 49.655 141.635 49.995 142.445 ;
        RECT 50.165 142.040 50.455 143.205 ;
        RECT 51.085 142.115 53.675 143.205 ;
        RECT 54.045 142.535 54.325 143.205 ;
        RECT 54.495 142.315 54.795 142.865 ;
        RECT 54.995 142.485 55.325 143.205 ;
        RECT 55.515 142.485 55.975 143.035 ;
        RECT 48.765 141.465 49.995 141.635 ;
        RECT 51.085 141.595 52.295 142.115 ;
        RECT 48.745 140.655 49.255 141.190 ;
        RECT 49.475 140.860 49.720 141.465 ;
        RECT 52.465 141.425 53.675 141.945 ;
        RECT 53.860 141.895 54.125 142.255 ;
        RECT 54.495 142.145 55.435 142.315 ;
        RECT 55.265 141.895 55.435 142.145 ;
        RECT 53.860 141.645 54.535 141.895 ;
        RECT 54.755 141.645 55.095 141.895 ;
        RECT 55.265 141.565 55.555 141.895 ;
        RECT 55.265 141.475 55.435 141.565 ;
        RECT 50.165 140.655 50.455 141.380 ;
        RECT 51.085 140.655 53.675 141.425 ;
        RECT 54.045 141.285 55.435 141.475 ;
        RECT 54.045 140.925 54.375 141.285 ;
        RECT 55.725 141.115 55.975 142.485 ;
        RECT 54.995 140.655 55.245 141.115 ;
        RECT 55.415 140.825 55.975 141.115 ;
        RECT 56.145 142.065 56.415 143.035 ;
        RECT 56.625 142.405 56.905 143.205 ;
        RECT 57.075 142.695 58.730 142.985 ;
        RECT 57.140 142.355 58.730 142.525 ;
        RECT 57.140 142.235 57.310 142.355 ;
        RECT 56.585 142.065 57.310 142.235 ;
        RECT 56.145 141.330 56.315 142.065 ;
        RECT 56.585 141.895 56.755 142.065 ;
        RECT 56.485 141.565 56.755 141.895 ;
        RECT 56.925 141.565 57.330 141.895 ;
        RECT 57.500 141.565 58.210 142.185 ;
        RECT 58.410 142.065 58.730 142.355 ;
        RECT 59.365 142.115 62.875 143.205 ;
        RECT 63.050 142.695 64.705 142.985 ;
        RECT 63.050 142.355 64.640 142.525 ;
        RECT 64.875 142.405 65.155 143.205 ;
        RECT 56.585 141.395 56.755 141.565 ;
        RECT 56.145 140.985 56.415 141.330 ;
        RECT 56.585 141.225 58.195 141.395 ;
        RECT 58.380 141.325 58.730 141.895 ;
        RECT 59.365 141.595 61.055 142.115 ;
        RECT 63.050 142.065 63.370 142.355 ;
        RECT 64.470 142.235 64.640 142.355 ;
        RECT 63.565 142.015 64.280 142.185 ;
        RECT 64.470 142.065 65.195 142.235 ;
        RECT 65.365 142.065 65.635 143.035 ;
        RECT 61.225 141.425 62.875 141.945 ;
        RECT 56.605 140.655 56.985 141.055 ;
        RECT 57.155 140.875 57.325 141.225 ;
        RECT 57.495 140.655 57.825 141.055 ;
        RECT 58.025 140.875 58.195 141.225 ;
        RECT 58.395 140.655 58.725 141.155 ;
        RECT 59.365 140.655 62.875 141.425 ;
        RECT 63.050 141.325 63.400 141.895 ;
        RECT 63.570 141.565 64.280 142.015 ;
        RECT 65.025 141.895 65.195 142.065 ;
        RECT 64.450 141.565 64.855 141.895 ;
        RECT 65.025 141.565 65.295 141.895 ;
        RECT 65.025 141.395 65.195 141.565 ;
        RECT 63.585 141.225 65.195 141.395 ;
        RECT 65.465 141.330 65.635 142.065 ;
        RECT 63.055 140.655 63.385 141.155 ;
        RECT 63.585 140.875 63.755 141.225 ;
        RECT 63.955 140.655 64.285 141.055 ;
        RECT 64.455 140.875 64.625 141.225 ;
        RECT 64.795 140.655 65.175 141.055 ;
        RECT 65.365 140.985 65.635 141.330 ;
        RECT 65.805 142.065 66.145 143.035 ;
        RECT 66.315 142.065 66.485 143.205 ;
        RECT 66.755 142.405 67.005 143.205 ;
        RECT 67.650 142.235 67.980 143.035 ;
        RECT 68.280 142.405 68.610 143.205 ;
        RECT 68.780 142.235 69.110 143.035 ;
        RECT 66.675 142.065 69.110 142.235 ;
        RECT 70.445 142.065 70.675 143.205 ;
        RECT 65.805 141.455 65.980 142.065 ;
        RECT 66.675 141.815 66.845 142.065 ;
        RECT 66.150 141.645 66.845 141.815 ;
        RECT 67.020 141.645 67.440 141.845 ;
        RECT 67.610 141.645 67.940 141.845 ;
        RECT 68.110 141.645 68.440 141.845 ;
        RECT 65.805 140.825 66.145 141.455 ;
        RECT 66.315 140.655 66.565 141.455 ;
        RECT 66.755 141.305 67.980 141.475 ;
        RECT 66.755 140.825 67.085 141.305 ;
        RECT 67.255 140.655 67.480 141.115 ;
        RECT 67.650 140.825 67.980 141.305 ;
        RECT 68.610 141.435 68.780 142.065 ;
        RECT 70.845 142.055 71.175 143.035 ;
        RECT 71.345 142.065 71.555 143.205 ;
        RECT 71.785 142.445 72.300 142.855 ;
        RECT 72.535 142.445 72.705 143.205 ;
        RECT 72.875 142.865 74.905 143.035 ;
        RECT 68.965 141.645 69.315 141.895 ;
        RECT 70.425 141.645 70.755 141.895 ;
        RECT 68.610 140.825 69.110 141.435 ;
        RECT 70.445 140.655 70.675 141.475 ;
        RECT 70.925 141.455 71.175 142.055 ;
        RECT 71.785 141.635 72.125 142.445 ;
        RECT 72.875 142.200 73.045 142.865 ;
        RECT 73.440 142.525 74.565 142.695 ;
        RECT 72.295 142.010 73.045 142.200 ;
        RECT 73.215 142.185 74.225 142.355 ;
        RECT 70.845 140.825 71.175 141.455 ;
        RECT 71.345 140.655 71.555 141.475 ;
        RECT 71.785 141.465 73.015 141.635 ;
        RECT 72.060 140.860 72.305 141.465 ;
        RECT 72.525 140.655 73.035 141.190 ;
        RECT 73.215 140.825 73.405 142.185 ;
        RECT 73.575 141.845 73.850 141.985 ;
        RECT 73.575 141.675 73.855 141.845 ;
        RECT 73.575 140.825 73.850 141.675 ;
        RECT 74.055 141.385 74.225 142.185 ;
        RECT 74.395 141.395 74.565 142.525 ;
        RECT 74.735 141.895 74.905 142.865 ;
        RECT 75.075 142.065 75.245 143.205 ;
        RECT 75.415 142.065 75.750 143.035 ;
        RECT 74.735 141.565 74.930 141.895 ;
        RECT 75.155 141.565 75.410 141.895 ;
        RECT 75.155 141.395 75.325 141.565 ;
        RECT 75.580 141.395 75.750 142.065 ;
        RECT 75.925 142.040 76.215 143.205 ;
        RECT 76.850 142.780 77.185 143.205 ;
        RECT 77.355 142.600 77.540 143.005 ;
        RECT 76.875 142.425 77.540 142.600 ;
        RECT 77.745 142.425 78.075 143.205 ;
        RECT 74.395 141.225 75.325 141.395 ;
        RECT 74.395 141.190 74.570 141.225 ;
        RECT 74.040 140.825 74.570 141.190 ;
        RECT 74.995 140.655 75.325 141.055 ;
        RECT 75.495 140.825 75.750 141.395 ;
        RECT 76.875 141.395 77.215 142.425 ;
        RECT 78.245 142.235 78.515 143.005 ;
        RECT 77.385 142.065 78.515 142.235 ;
        RECT 77.385 141.565 77.635 142.065 ;
        RECT 75.925 140.655 76.215 141.380 ;
        RECT 76.875 141.225 77.560 141.395 ;
        RECT 77.815 141.315 78.175 141.895 ;
        RECT 76.850 140.655 77.185 141.055 ;
        RECT 77.355 140.825 77.560 141.225 ;
        RECT 78.345 141.155 78.515 142.065 ;
        RECT 77.770 140.655 78.045 141.135 ;
        RECT 78.255 140.825 78.515 141.155 ;
        RECT 78.685 142.485 79.145 143.035 ;
        RECT 79.335 142.485 79.665 143.205 ;
        RECT 78.685 141.115 78.935 142.485 ;
        RECT 79.865 142.315 80.165 142.865 ;
        RECT 80.335 142.535 80.615 143.205 ;
        RECT 79.225 142.145 80.165 142.315 ;
        RECT 79.225 141.895 79.395 142.145 ;
        RECT 80.535 141.895 80.800 142.255 ;
        RECT 79.105 141.565 79.395 141.895 ;
        RECT 79.565 141.645 79.905 141.895 ;
        RECT 80.125 141.645 80.800 141.895 ;
        RECT 81.445 142.065 81.715 143.035 ;
        RECT 81.925 142.405 82.205 143.205 ;
        RECT 82.375 142.695 84.030 142.985 ;
        RECT 82.440 142.355 84.030 142.525 ;
        RECT 82.440 142.235 82.610 142.355 ;
        RECT 81.885 142.065 82.610 142.235 ;
        RECT 79.225 141.475 79.395 141.565 ;
        RECT 79.225 141.285 80.615 141.475 ;
        RECT 78.685 140.825 79.245 141.115 ;
        RECT 79.415 140.655 79.665 141.115 ;
        RECT 80.285 140.925 80.615 141.285 ;
        RECT 81.445 141.330 81.615 142.065 ;
        RECT 81.885 141.895 82.055 142.065 ;
        RECT 82.800 142.015 83.515 142.185 ;
        RECT 83.710 142.065 84.030 142.355 ;
        RECT 84.205 142.065 84.545 143.035 ;
        RECT 84.715 142.065 84.885 143.205 ;
        RECT 85.155 142.405 85.405 143.205 ;
        RECT 86.050 142.235 86.380 143.035 ;
        RECT 86.680 142.405 87.010 143.205 ;
        RECT 87.180 142.235 87.510 143.035 ;
        RECT 85.075 142.065 87.510 142.235 ;
        RECT 88.895 142.275 89.065 143.035 ;
        RECT 89.245 142.445 89.575 143.205 ;
        RECT 88.895 142.105 89.560 142.275 ;
        RECT 89.745 142.130 90.015 143.035 ;
        RECT 81.785 141.565 82.055 141.895 ;
        RECT 82.225 141.565 82.630 141.895 ;
        RECT 82.800 141.565 83.510 142.015 ;
        RECT 81.885 141.395 82.055 141.565 ;
        RECT 81.445 140.985 81.715 141.330 ;
        RECT 81.885 141.225 83.495 141.395 ;
        RECT 83.680 141.325 84.030 141.895 ;
        RECT 84.205 141.505 84.380 142.065 ;
        RECT 85.075 141.815 85.245 142.065 ;
        RECT 84.550 141.645 85.245 141.815 ;
        RECT 85.420 141.645 85.840 141.845 ;
        RECT 86.010 141.645 86.340 141.845 ;
        RECT 86.510 141.645 86.840 141.845 ;
        RECT 84.205 141.455 84.435 141.505 ;
        RECT 81.905 140.655 82.285 141.055 ;
        RECT 82.455 140.875 82.625 141.225 ;
        RECT 82.795 140.655 83.125 141.055 ;
        RECT 83.325 140.875 83.495 141.225 ;
        RECT 83.695 140.655 84.025 141.155 ;
        RECT 84.205 140.825 84.545 141.455 ;
        RECT 84.715 140.655 84.965 141.455 ;
        RECT 85.155 141.305 86.380 141.475 ;
        RECT 85.155 140.825 85.485 141.305 ;
        RECT 85.655 140.655 85.880 141.115 ;
        RECT 86.050 140.825 86.380 141.305 ;
        RECT 87.010 141.435 87.180 142.065 ;
        RECT 89.390 141.960 89.560 142.105 ;
        RECT 87.365 141.645 87.715 141.895 ;
        RECT 88.825 141.555 89.155 141.925 ;
        RECT 89.390 141.630 89.675 141.960 ;
        RECT 87.010 140.825 87.510 141.435 ;
        RECT 89.390 141.375 89.560 141.630 ;
        RECT 88.895 141.205 89.560 141.375 ;
        RECT 89.845 141.330 90.015 142.130 ;
        RECT 90.245 142.065 90.455 143.205 ;
        RECT 90.625 142.055 90.955 143.035 ;
        RECT 91.125 142.065 91.355 143.205 ;
        RECT 91.940 142.225 92.195 142.895 ;
        RECT 92.375 142.405 92.660 143.205 ;
        RECT 92.840 142.485 93.170 142.995 ;
        RECT 91.940 142.185 92.120 142.225 ;
        RECT 88.895 140.825 89.065 141.205 ;
        RECT 89.245 140.655 89.575 141.035 ;
        RECT 89.755 140.825 90.015 141.330 ;
        RECT 90.245 140.655 90.455 141.475 ;
        RECT 90.625 141.455 90.875 142.055 ;
        RECT 91.855 142.015 92.120 142.185 ;
        RECT 91.045 141.645 91.375 141.895 ;
        RECT 90.625 140.825 90.955 141.455 ;
        RECT 91.125 140.655 91.355 141.475 ;
        RECT 91.940 141.365 92.120 142.015 ;
        RECT 92.840 141.895 93.090 142.485 ;
        RECT 93.440 142.335 93.610 142.945 ;
        RECT 93.780 142.515 94.110 143.205 ;
        RECT 94.340 142.655 94.580 142.945 ;
        RECT 94.780 142.825 95.200 143.205 ;
        RECT 95.380 142.735 96.010 142.985 ;
        RECT 96.480 142.825 96.810 143.205 ;
        RECT 95.380 142.655 95.550 142.735 ;
        RECT 96.980 142.655 97.150 142.945 ;
        RECT 97.330 142.825 97.710 143.205 ;
        RECT 97.950 142.820 98.780 142.990 ;
        RECT 94.340 142.485 95.550 142.655 ;
        RECT 92.290 141.565 93.090 141.895 ;
        RECT 91.940 140.835 92.195 141.365 ;
        RECT 92.375 140.655 92.660 141.115 ;
        RECT 92.840 140.915 93.090 141.565 ;
        RECT 93.290 142.315 93.610 142.335 ;
        RECT 93.290 142.145 95.210 142.315 ;
        RECT 93.290 141.250 93.480 142.145 ;
        RECT 95.380 141.975 95.550 142.485 ;
        RECT 95.720 142.225 96.240 142.535 ;
        RECT 93.650 141.805 95.550 141.975 ;
        RECT 93.650 141.745 93.980 141.805 ;
        RECT 94.130 141.575 94.460 141.635 ;
        RECT 93.800 141.305 94.460 141.575 ;
        RECT 93.290 140.920 93.610 141.250 ;
        RECT 93.790 140.655 94.450 141.135 ;
        RECT 94.650 141.045 94.820 141.805 ;
        RECT 95.720 141.635 95.900 142.045 ;
        RECT 94.990 141.465 95.320 141.585 ;
        RECT 96.070 141.465 96.240 142.225 ;
        RECT 94.990 141.295 96.240 141.465 ;
        RECT 96.410 142.405 97.780 142.655 ;
        RECT 96.410 141.635 96.600 142.405 ;
        RECT 97.530 142.145 97.780 142.405 ;
        RECT 96.770 141.975 97.020 142.135 ;
        RECT 97.950 141.975 98.120 142.820 ;
        RECT 99.015 142.535 99.185 143.035 ;
        RECT 99.355 142.705 99.685 143.205 ;
        RECT 98.290 142.145 98.790 142.525 ;
        RECT 99.015 142.365 99.710 142.535 ;
        RECT 96.770 141.805 98.120 141.975 ;
        RECT 97.700 141.765 98.120 141.805 ;
        RECT 96.410 141.295 96.830 141.635 ;
        RECT 97.120 141.305 97.530 141.635 ;
        RECT 94.650 140.875 95.500 141.045 ;
        RECT 96.060 140.655 96.380 141.115 ;
        RECT 96.580 140.865 96.830 141.295 ;
        RECT 97.120 140.655 97.530 141.095 ;
        RECT 97.700 141.035 97.870 141.765 ;
        RECT 98.040 141.215 98.390 141.585 ;
        RECT 98.570 141.275 98.790 142.145 ;
        RECT 98.960 141.575 99.370 142.195 ;
        RECT 99.540 141.395 99.710 142.365 ;
        RECT 99.015 141.205 99.710 141.395 ;
        RECT 97.700 140.835 98.715 141.035 ;
        RECT 99.015 140.875 99.185 141.205 ;
        RECT 99.355 140.655 99.685 141.035 ;
        RECT 99.900 140.915 100.125 143.035 ;
        RECT 100.295 142.705 100.625 143.205 ;
        RECT 100.795 142.535 100.965 143.035 ;
        RECT 100.300 142.365 100.965 142.535 ;
        RECT 100.300 141.375 100.530 142.365 ;
        RECT 100.700 141.545 101.050 142.195 ;
        RECT 101.685 142.040 101.975 143.205 ;
        RECT 103.065 142.115 106.575 143.205 ;
        RECT 106.945 142.535 107.225 143.205 ;
        RECT 107.395 142.315 107.695 142.865 ;
        RECT 107.895 142.485 108.225 143.205 ;
        RECT 108.415 142.485 108.875 143.035 ;
        RECT 103.065 141.595 104.755 142.115 ;
        RECT 104.925 141.425 106.575 141.945 ;
        RECT 106.760 141.895 107.025 142.255 ;
        RECT 107.395 142.145 108.335 142.315 ;
        RECT 108.165 141.895 108.335 142.145 ;
        RECT 106.760 141.645 107.435 141.895 ;
        RECT 107.655 141.645 107.995 141.895 ;
        RECT 108.165 141.565 108.455 141.895 ;
        RECT 108.165 141.475 108.335 141.565 ;
        RECT 100.300 141.205 100.965 141.375 ;
        RECT 100.295 140.655 100.625 141.035 ;
        RECT 100.795 140.915 100.965 141.205 ;
        RECT 101.685 140.655 101.975 141.380 ;
        RECT 103.065 140.655 106.575 141.425 ;
        RECT 106.945 141.285 108.335 141.475 ;
        RECT 106.945 140.925 107.275 141.285 ;
        RECT 108.625 141.115 108.875 142.485 ;
        RECT 109.045 142.115 110.255 143.205 ;
        RECT 110.625 142.535 110.905 143.205 ;
        RECT 111.075 142.315 111.375 142.865 ;
        RECT 111.575 142.485 111.905 143.205 ;
        RECT 112.095 142.485 112.555 143.035 ;
        RECT 109.045 141.575 109.565 142.115 ;
        RECT 109.735 141.405 110.255 141.945 ;
        RECT 110.440 141.895 110.705 142.255 ;
        RECT 111.075 142.145 112.015 142.315 ;
        RECT 111.845 141.895 112.015 142.145 ;
        RECT 110.440 141.645 111.115 141.895 ;
        RECT 111.335 141.645 111.675 141.895 ;
        RECT 111.845 141.565 112.135 141.895 ;
        RECT 111.845 141.475 112.015 141.565 ;
        RECT 107.895 140.655 108.145 141.115 ;
        RECT 108.315 140.825 108.875 141.115 ;
        RECT 109.045 140.655 110.255 141.405 ;
        RECT 110.625 141.285 112.015 141.475 ;
        RECT 110.625 140.925 110.955 141.285 ;
        RECT 112.305 141.115 112.555 142.485 ;
        RECT 111.575 140.655 111.825 141.115 ;
        RECT 111.995 140.825 112.555 141.115 ;
        RECT 112.725 142.485 113.185 143.035 ;
        RECT 113.375 142.485 113.705 143.205 ;
        RECT 112.725 141.115 112.975 142.485 ;
        RECT 113.905 142.315 114.205 142.865 ;
        RECT 114.375 142.535 114.655 143.205 ;
        RECT 113.265 142.145 114.205 142.315 ;
        RECT 115.025 142.445 115.540 142.855 ;
        RECT 115.775 142.445 115.945 143.205 ;
        RECT 116.115 142.865 118.145 143.035 ;
        RECT 113.265 141.895 113.435 142.145 ;
        RECT 114.575 141.895 114.840 142.255 ;
        RECT 113.145 141.565 113.435 141.895 ;
        RECT 113.605 141.645 113.945 141.895 ;
        RECT 114.165 141.645 114.840 141.895 ;
        RECT 113.265 141.475 113.435 141.565 ;
        RECT 115.025 141.635 115.365 142.445 ;
        RECT 116.115 142.200 116.285 142.865 ;
        RECT 116.680 142.525 117.805 142.695 ;
        RECT 115.535 142.010 116.285 142.200 ;
        RECT 116.455 142.185 117.465 142.355 ;
        RECT 113.265 141.285 114.655 141.475 ;
        RECT 115.025 141.465 116.255 141.635 ;
        RECT 112.725 140.825 113.285 141.115 ;
        RECT 113.455 140.655 113.705 141.115 ;
        RECT 114.325 140.925 114.655 141.285 ;
        RECT 115.300 140.860 115.545 141.465 ;
        RECT 115.765 140.655 116.275 141.190 ;
        RECT 116.455 140.825 116.645 142.185 ;
        RECT 116.815 141.165 117.090 141.985 ;
        RECT 117.295 141.385 117.465 142.185 ;
        RECT 117.635 141.395 117.805 142.525 ;
        RECT 117.975 141.895 118.145 142.865 ;
        RECT 118.315 142.065 118.485 143.205 ;
        RECT 118.655 142.065 118.990 143.035 ;
        RECT 117.975 141.565 118.170 141.895 ;
        RECT 118.395 141.565 118.650 141.895 ;
        RECT 118.395 141.395 118.565 141.565 ;
        RECT 118.820 141.395 118.990 142.065 ;
        RECT 119.165 142.115 120.835 143.205 ;
        RECT 121.010 142.770 126.355 143.205 ;
        RECT 119.165 141.595 119.915 142.115 ;
        RECT 120.085 141.425 120.835 141.945 ;
        RECT 122.600 141.520 122.950 142.770 ;
        RECT 126.525 142.115 127.735 143.205 ;
        RECT 117.635 141.225 118.565 141.395 ;
        RECT 117.635 141.190 117.810 141.225 ;
        RECT 116.815 140.995 117.095 141.165 ;
        RECT 116.815 140.825 117.090 140.995 ;
        RECT 117.280 140.825 117.810 141.190 ;
        RECT 118.235 140.655 118.565 141.055 ;
        RECT 118.735 140.825 118.990 141.395 ;
        RECT 119.165 140.655 120.835 141.425 ;
        RECT 124.430 141.200 124.770 142.030 ;
        RECT 126.525 141.575 127.045 142.115 ;
        RECT 127.215 141.405 127.735 141.945 ;
        RECT 121.010 140.655 126.355 141.200 ;
        RECT 126.525 140.655 127.735 141.405 ;
        RECT 29.840 140.485 127.820 140.655 ;
        RECT 29.925 139.735 31.135 140.485 ;
        RECT 29.925 139.195 30.445 139.735 ;
        RECT 31.825 139.665 32.035 140.485 ;
        RECT 32.205 139.685 32.535 140.315 ;
        RECT 30.615 139.025 31.135 139.565 ;
        RECT 32.205 139.085 32.455 139.685 ;
        RECT 32.705 139.665 32.935 140.485 ;
        RECT 33.420 139.675 33.665 140.280 ;
        RECT 33.885 139.950 34.395 140.485 ;
        RECT 33.145 139.505 34.375 139.675 ;
        RECT 32.625 139.245 32.955 139.495 ;
        RECT 29.925 137.935 31.135 139.025 ;
        RECT 31.825 137.935 32.035 139.075 ;
        RECT 32.205 138.105 32.535 139.085 ;
        RECT 32.705 137.935 32.935 139.075 ;
        RECT 33.145 138.695 33.485 139.505 ;
        RECT 33.655 138.940 34.405 139.130 ;
        RECT 33.145 138.285 33.660 138.695 ;
        RECT 33.895 137.935 34.065 138.695 ;
        RECT 34.235 138.275 34.405 138.940 ;
        RECT 34.575 138.955 34.765 140.315 ;
        RECT 34.935 140.145 35.210 140.315 ;
        RECT 34.935 139.975 35.215 140.145 ;
        RECT 34.935 139.155 35.210 139.975 ;
        RECT 35.400 139.950 35.930 140.315 ;
        RECT 36.355 140.085 36.685 140.485 ;
        RECT 35.755 139.915 35.930 139.950 ;
        RECT 35.415 138.955 35.585 139.755 ;
        RECT 34.575 138.785 35.585 138.955 ;
        RECT 35.755 139.745 36.685 139.915 ;
        RECT 36.855 139.745 37.110 140.315 ;
        RECT 37.285 139.760 37.575 140.485 ;
        RECT 35.755 138.615 35.925 139.745 ;
        RECT 36.515 139.575 36.685 139.745 ;
        RECT 34.800 138.445 35.925 138.615 ;
        RECT 36.095 139.245 36.290 139.575 ;
        RECT 36.515 139.245 36.770 139.575 ;
        RECT 36.095 138.275 36.265 139.245 ;
        RECT 36.940 139.075 37.110 139.745 ;
        RECT 37.745 139.735 38.955 140.485 ;
        RECT 39.215 139.935 39.385 140.315 ;
        RECT 39.565 140.105 39.895 140.485 ;
        RECT 39.215 139.765 39.880 139.935 ;
        RECT 40.075 139.810 40.335 140.315 ;
        RECT 34.235 138.105 36.265 138.275 ;
        RECT 36.435 137.935 36.605 139.075 ;
        RECT 36.775 138.105 37.110 139.075 ;
        RECT 37.285 137.935 37.575 139.100 ;
        RECT 37.745 139.025 38.265 139.565 ;
        RECT 38.435 139.195 38.955 139.735 ;
        RECT 39.145 139.215 39.475 139.585 ;
        RECT 39.710 139.510 39.880 139.765 ;
        RECT 39.710 139.180 39.995 139.510 ;
        RECT 39.710 139.035 39.880 139.180 ;
        RECT 37.745 137.935 38.955 139.025 ;
        RECT 39.215 138.865 39.880 139.035 ;
        RECT 40.165 139.010 40.335 139.810 ;
        RECT 41.515 139.935 41.685 140.315 ;
        RECT 41.865 140.105 42.195 140.485 ;
        RECT 41.515 139.765 42.180 139.935 ;
        RECT 42.375 139.810 42.635 140.315 ;
        RECT 41.445 139.215 41.775 139.585 ;
        RECT 42.010 139.510 42.180 139.765 ;
        RECT 42.010 139.180 42.295 139.510 ;
        RECT 42.010 139.035 42.180 139.180 ;
        RECT 39.215 138.105 39.385 138.865 ;
        RECT 39.565 137.935 39.895 138.695 ;
        RECT 40.065 138.105 40.335 139.010 ;
        RECT 41.515 138.865 42.180 139.035 ;
        RECT 42.465 139.010 42.635 139.810 ;
        RECT 42.895 139.935 43.065 140.225 ;
        RECT 43.235 140.105 43.565 140.485 ;
        RECT 42.895 139.765 43.560 139.935 ;
        RECT 41.515 138.105 41.685 138.865 ;
        RECT 41.865 137.935 42.195 138.695 ;
        RECT 42.365 138.105 42.635 139.010 ;
        RECT 42.810 138.945 43.160 139.595 ;
        RECT 43.330 138.775 43.560 139.765 ;
        RECT 42.895 138.605 43.560 138.775 ;
        RECT 42.895 138.105 43.065 138.605 ;
        RECT 43.235 137.935 43.565 138.435 ;
        RECT 43.735 138.105 43.960 140.225 ;
        RECT 44.175 140.105 44.505 140.485 ;
        RECT 44.675 139.935 44.845 140.265 ;
        RECT 45.145 140.105 46.160 140.305 ;
        RECT 44.150 139.745 44.845 139.935 ;
        RECT 44.150 138.775 44.320 139.745 ;
        RECT 44.490 138.945 44.900 139.565 ;
        RECT 45.070 138.995 45.290 139.865 ;
        RECT 45.470 139.555 45.820 139.925 ;
        RECT 45.990 139.375 46.160 140.105 ;
        RECT 46.330 140.045 46.740 140.485 ;
        RECT 47.030 139.845 47.280 140.275 ;
        RECT 47.480 140.025 47.800 140.485 ;
        RECT 48.360 140.095 49.210 140.265 ;
        RECT 46.330 139.505 46.740 139.835 ;
        RECT 47.030 139.505 47.450 139.845 ;
        RECT 45.740 139.335 46.160 139.375 ;
        RECT 45.740 139.165 47.090 139.335 ;
        RECT 44.150 138.605 44.845 138.775 ;
        RECT 45.070 138.615 45.570 138.995 ;
        RECT 44.175 137.935 44.505 138.435 ;
        RECT 44.675 138.105 44.845 138.605 ;
        RECT 45.740 138.320 45.910 139.165 ;
        RECT 46.840 139.005 47.090 139.165 ;
        RECT 46.080 138.735 46.330 138.995 ;
        RECT 47.260 138.735 47.450 139.505 ;
        RECT 46.080 138.485 47.450 138.735 ;
        RECT 47.620 139.675 48.870 139.845 ;
        RECT 47.620 138.915 47.790 139.675 ;
        RECT 48.540 139.555 48.870 139.675 ;
        RECT 47.960 139.095 48.140 139.505 ;
        RECT 49.040 139.335 49.210 140.095 ;
        RECT 49.410 140.005 50.070 140.485 ;
        RECT 50.250 139.890 50.570 140.220 ;
        RECT 49.400 139.565 50.060 139.835 ;
        RECT 49.400 139.505 49.730 139.565 ;
        RECT 49.880 139.335 50.210 139.395 ;
        RECT 48.310 139.165 50.210 139.335 ;
        RECT 47.620 138.605 48.140 138.915 ;
        RECT 48.310 138.655 48.480 139.165 ;
        RECT 50.380 138.995 50.570 139.890 ;
        RECT 48.650 138.825 50.570 138.995 ;
        RECT 50.250 138.805 50.570 138.825 ;
        RECT 50.770 139.575 51.020 140.225 ;
        RECT 51.200 140.025 51.485 140.485 ;
        RECT 51.665 139.775 51.920 140.305 ;
        RECT 52.525 140.005 52.805 140.485 ;
        RECT 52.975 139.835 53.235 140.225 ;
        RECT 53.410 140.005 53.665 140.485 ;
        RECT 53.835 139.835 54.130 140.225 ;
        RECT 54.310 140.005 54.585 140.485 ;
        RECT 54.755 139.985 55.055 140.315 ;
        RECT 50.770 139.245 51.570 139.575 ;
        RECT 48.310 138.485 49.520 138.655 ;
        RECT 45.080 138.150 45.910 138.320 ;
        RECT 46.150 137.935 46.530 138.315 ;
        RECT 46.710 138.195 46.880 138.485 ;
        RECT 48.310 138.405 48.480 138.485 ;
        RECT 47.050 137.935 47.380 138.315 ;
        RECT 47.850 138.155 48.480 138.405 ;
        RECT 48.660 137.935 49.080 138.315 ;
        RECT 49.280 138.195 49.520 138.485 ;
        RECT 49.750 137.935 50.080 138.625 ;
        RECT 50.250 138.195 50.420 138.805 ;
        RECT 50.770 138.655 51.020 139.245 ;
        RECT 51.740 139.125 51.920 139.775 ;
        RECT 52.480 139.665 54.130 139.835 ;
        RECT 52.480 139.155 52.885 139.665 ;
        RECT 53.055 139.325 54.195 139.495 ;
        RECT 51.740 138.955 52.005 139.125 ;
        RECT 52.480 138.985 53.235 139.155 ;
        RECT 51.740 138.915 51.920 138.955 ;
        RECT 50.690 138.145 51.020 138.655 ;
        RECT 51.200 137.935 51.485 138.735 ;
        RECT 51.665 138.245 51.920 138.915 ;
        RECT 52.520 137.935 52.805 138.805 ;
        RECT 52.975 138.735 53.235 138.985 ;
        RECT 54.025 139.075 54.195 139.325 ;
        RECT 54.365 139.245 54.715 139.815 ;
        RECT 54.885 139.075 55.055 139.985 ;
        RECT 54.025 138.905 55.055 139.075 ;
        RECT 52.975 138.565 54.095 138.735 ;
        RECT 52.975 138.105 53.235 138.565 ;
        RECT 53.410 137.935 53.665 138.395 ;
        RECT 53.835 138.105 54.095 138.565 ;
        RECT 54.265 137.935 54.575 138.735 ;
        RECT 54.745 138.105 55.055 138.905 ;
        RECT 55.225 139.810 55.485 140.315 ;
        RECT 55.665 140.105 55.995 140.485 ;
        RECT 56.175 139.935 56.345 140.315 ;
        RECT 55.225 139.010 55.395 139.810 ;
        RECT 55.680 139.765 56.345 139.935 ;
        RECT 56.605 139.810 56.875 140.155 ;
        RECT 57.065 140.085 57.445 140.485 ;
        RECT 57.615 139.915 57.785 140.265 ;
        RECT 57.955 140.085 58.285 140.485 ;
        RECT 58.485 139.915 58.655 140.265 ;
        RECT 58.855 139.985 59.185 140.485 ;
        RECT 55.680 139.510 55.850 139.765 ;
        RECT 55.565 139.180 55.850 139.510 ;
        RECT 56.085 139.215 56.415 139.585 ;
        RECT 55.680 139.035 55.850 139.180 ;
        RECT 56.605 139.075 56.775 139.810 ;
        RECT 57.045 139.745 58.655 139.915 ;
        RECT 57.045 139.575 57.215 139.745 ;
        RECT 56.945 139.245 57.215 139.575 ;
        RECT 57.385 139.245 57.790 139.575 ;
        RECT 57.045 139.075 57.215 139.245 ;
        RECT 55.225 138.105 55.495 139.010 ;
        RECT 55.680 138.865 56.345 139.035 ;
        RECT 55.665 137.935 55.995 138.695 ;
        RECT 56.175 138.105 56.345 138.865 ;
        RECT 56.605 138.105 56.875 139.075 ;
        RECT 57.045 138.905 57.770 139.075 ;
        RECT 57.960 138.955 58.670 139.575 ;
        RECT 58.840 139.245 59.190 139.815 ;
        RECT 59.365 139.685 59.705 140.315 ;
        RECT 59.875 139.685 60.125 140.485 ;
        RECT 60.315 139.835 60.645 140.315 ;
        RECT 60.815 140.025 61.040 140.485 ;
        RECT 61.210 139.835 61.540 140.315 ;
        RECT 59.365 139.075 59.540 139.685 ;
        RECT 60.315 139.665 61.540 139.835 ;
        RECT 62.170 139.705 62.670 140.315 ;
        RECT 63.045 139.760 63.335 140.485 ;
        RECT 63.975 139.985 64.305 140.485 ;
        RECT 64.505 139.915 64.675 140.265 ;
        RECT 64.875 140.085 65.205 140.485 ;
        RECT 65.375 139.915 65.545 140.265 ;
        RECT 65.715 140.085 66.095 140.485 ;
        RECT 59.710 139.325 60.405 139.495 ;
        RECT 60.235 139.075 60.405 139.325 ;
        RECT 60.580 139.295 61.000 139.495 ;
        RECT 61.170 139.295 61.500 139.495 ;
        RECT 61.670 139.295 62.000 139.495 ;
        RECT 62.170 139.075 62.340 139.705 ;
        RECT 62.525 139.245 62.875 139.495 ;
        RECT 63.970 139.245 64.320 139.815 ;
        RECT 64.505 139.745 66.115 139.915 ;
        RECT 66.285 139.810 66.555 140.155 ;
        RECT 65.945 139.575 66.115 139.745 ;
        RECT 57.600 138.785 57.770 138.905 ;
        RECT 58.870 138.785 59.190 139.075 ;
        RECT 57.085 137.935 57.365 138.735 ;
        RECT 57.600 138.615 59.190 138.785 ;
        RECT 57.535 138.155 59.190 138.445 ;
        RECT 59.365 138.105 59.705 139.075 ;
        RECT 59.875 137.935 60.045 139.075 ;
        RECT 60.235 138.905 62.670 139.075 ;
        RECT 60.315 137.935 60.565 138.735 ;
        RECT 61.210 138.105 61.540 138.905 ;
        RECT 61.840 137.935 62.170 138.735 ;
        RECT 62.340 138.105 62.670 138.905 ;
        RECT 63.045 137.935 63.335 139.100 ;
        RECT 63.970 138.785 64.290 139.075 ;
        RECT 64.490 138.955 65.200 139.575 ;
        RECT 65.370 139.245 65.775 139.575 ;
        RECT 65.945 139.245 66.215 139.575 ;
        RECT 65.945 139.075 66.115 139.245 ;
        RECT 66.385 139.075 66.555 139.810 ;
        RECT 65.390 138.905 66.115 139.075 ;
        RECT 65.390 138.785 65.560 138.905 ;
        RECT 63.970 138.615 65.560 138.785 ;
        RECT 63.970 138.155 65.625 138.445 ;
        RECT 65.795 137.935 66.075 138.735 ;
        RECT 66.285 138.105 66.555 139.075 ;
        RECT 66.725 139.685 67.065 140.315 ;
        RECT 67.235 139.685 67.485 140.485 ;
        RECT 67.675 139.835 68.005 140.315 ;
        RECT 68.175 140.025 68.400 140.485 ;
        RECT 68.570 139.835 68.900 140.315 ;
        RECT 66.725 139.635 66.955 139.685 ;
        RECT 67.675 139.665 68.900 139.835 ;
        RECT 69.530 139.705 70.030 140.315 ;
        RECT 70.780 139.775 71.035 140.305 ;
        RECT 71.215 140.025 71.500 140.485 ;
        RECT 66.725 139.075 66.900 139.635 ;
        RECT 67.070 139.325 67.765 139.495 ;
        RECT 67.595 139.075 67.765 139.325 ;
        RECT 67.940 139.295 68.360 139.495 ;
        RECT 68.530 139.295 68.860 139.495 ;
        RECT 69.030 139.295 69.360 139.495 ;
        RECT 69.530 139.075 69.700 139.705 ;
        RECT 69.885 139.245 70.235 139.495 ;
        RECT 66.725 138.105 67.065 139.075 ;
        RECT 67.235 137.935 67.405 139.075 ;
        RECT 67.595 138.905 70.030 139.075 ;
        RECT 67.675 137.935 67.925 138.735 ;
        RECT 68.570 138.105 68.900 138.905 ;
        RECT 69.200 137.935 69.530 138.735 ;
        RECT 69.700 138.105 70.030 138.905 ;
        RECT 70.780 138.915 70.960 139.775 ;
        RECT 71.680 139.575 71.930 140.225 ;
        RECT 71.130 139.245 71.930 139.575 ;
        RECT 70.780 138.445 71.035 138.915 ;
        RECT 70.695 138.275 71.035 138.445 ;
        RECT 70.780 138.245 71.035 138.275 ;
        RECT 71.215 137.935 71.500 138.735 ;
        RECT 71.680 138.655 71.930 139.245 ;
        RECT 72.130 139.890 72.450 140.220 ;
        RECT 72.630 140.005 73.290 140.485 ;
        RECT 73.490 140.095 74.340 140.265 ;
        RECT 72.130 138.995 72.320 139.890 ;
        RECT 72.640 139.565 73.300 139.835 ;
        RECT 72.970 139.505 73.300 139.565 ;
        RECT 72.490 139.335 72.820 139.395 ;
        RECT 73.490 139.335 73.660 140.095 ;
        RECT 74.900 140.025 75.220 140.485 ;
        RECT 75.420 139.845 75.670 140.275 ;
        RECT 75.960 140.045 76.370 140.485 ;
        RECT 76.540 140.105 77.555 140.305 ;
        RECT 73.830 139.675 75.080 139.845 ;
        RECT 73.830 139.555 74.160 139.675 ;
        RECT 72.490 139.165 74.390 139.335 ;
        RECT 72.130 138.825 74.050 138.995 ;
        RECT 72.130 138.805 72.450 138.825 ;
        RECT 71.680 138.145 72.010 138.655 ;
        RECT 72.280 138.195 72.450 138.805 ;
        RECT 74.220 138.655 74.390 139.165 ;
        RECT 74.560 139.095 74.740 139.505 ;
        RECT 74.910 138.915 75.080 139.675 ;
        RECT 72.620 137.935 72.950 138.625 ;
        RECT 73.180 138.485 74.390 138.655 ;
        RECT 74.560 138.605 75.080 138.915 ;
        RECT 75.250 139.505 75.670 139.845 ;
        RECT 75.960 139.505 76.370 139.835 ;
        RECT 75.250 138.735 75.440 139.505 ;
        RECT 76.540 139.375 76.710 140.105 ;
        RECT 77.855 139.935 78.025 140.265 ;
        RECT 78.195 140.105 78.525 140.485 ;
        RECT 76.880 139.555 77.230 139.925 ;
        RECT 76.540 139.335 76.960 139.375 ;
        RECT 75.610 139.165 76.960 139.335 ;
        RECT 75.610 139.005 75.860 139.165 ;
        RECT 76.370 138.735 76.620 138.995 ;
        RECT 75.250 138.485 76.620 138.735 ;
        RECT 73.180 138.195 73.420 138.485 ;
        RECT 74.220 138.405 74.390 138.485 ;
        RECT 73.620 137.935 74.040 138.315 ;
        RECT 74.220 138.155 74.850 138.405 ;
        RECT 75.320 137.935 75.650 138.315 ;
        RECT 75.820 138.195 75.990 138.485 ;
        RECT 76.790 138.320 76.960 139.165 ;
        RECT 77.410 138.995 77.630 139.865 ;
        RECT 77.855 139.745 78.550 139.935 ;
        RECT 77.130 138.615 77.630 138.995 ;
        RECT 77.800 138.945 78.210 139.565 ;
        RECT 78.380 138.775 78.550 139.745 ;
        RECT 77.855 138.605 78.550 138.775 ;
        RECT 76.170 137.935 76.550 138.315 ;
        RECT 76.790 138.150 77.620 138.320 ;
        RECT 77.855 138.105 78.025 138.605 ;
        RECT 78.195 137.935 78.525 138.435 ;
        RECT 78.740 138.105 78.965 140.225 ;
        RECT 79.135 140.105 79.465 140.485 ;
        RECT 79.635 139.935 79.805 140.225 ;
        RECT 79.140 139.765 79.805 139.935 ;
        RECT 80.065 139.985 80.365 140.315 ;
        RECT 80.535 140.005 80.810 140.485 ;
        RECT 79.140 138.775 79.370 139.765 ;
        RECT 79.540 138.945 79.890 139.595 ;
        RECT 80.065 139.075 80.235 139.985 ;
        RECT 80.990 139.835 81.285 140.225 ;
        RECT 81.455 140.005 81.710 140.485 ;
        RECT 81.885 139.835 82.145 140.225 ;
        RECT 82.315 140.005 82.595 140.485 ;
        RECT 80.405 139.245 80.755 139.815 ;
        RECT 80.990 139.665 82.640 139.835 ;
        RECT 82.825 139.715 86.335 140.485 ;
        RECT 80.925 139.325 82.065 139.495 ;
        RECT 80.925 139.075 81.095 139.325 ;
        RECT 82.235 139.155 82.640 139.665 ;
        RECT 80.065 138.905 81.095 139.075 ;
        RECT 81.885 138.985 82.640 139.155 ;
        RECT 82.825 139.025 84.515 139.545 ;
        RECT 84.685 139.195 86.335 139.715 ;
        RECT 86.505 140.025 87.065 140.315 ;
        RECT 87.235 140.025 87.485 140.485 ;
        RECT 79.140 138.605 79.805 138.775 ;
        RECT 79.135 137.935 79.465 138.435 ;
        RECT 79.635 138.105 79.805 138.605 ;
        RECT 80.065 138.105 80.375 138.905 ;
        RECT 81.885 138.735 82.145 138.985 ;
        RECT 80.545 137.935 80.855 138.735 ;
        RECT 81.025 138.565 82.145 138.735 ;
        RECT 81.025 138.105 81.285 138.565 ;
        RECT 81.455 137.935 81.710 138.395 ;
        RECT 81.885 138.105 82.145 138.565 ;
        RECT 82.315 137.935 82.600 138.805 ;
        RECT 82.825 137.935 86.335 139.025 ;
        RECT 86.505 138.655 86.755 140.025 ;
        RECT 88.105 139.855 88.435 140.215 ;
        RECT 87.045 139.665 88.435 139.855 ;
        RECT 88.805 139.760 89.095 140.485 ;
        RECT 89.725 139.715 92.315 140.485 ;
        RECT 92.575 139.935 92.745 140.315 ;
        RECT 92.925 140.105 93.255 140.485 ;
        RECT 92.575 139.765 93.240 139.935 ;
        RECT 93.435 139.810 93.695 140.315 ;
        RECT 87.045 139.575 87.215 139.665 ;
        RECT 86.925 139.245 87.215 139.575 ;
        RECT 87.385 139.245 87.725 139.495 ;
        RECT 87.945 139.245 88.620 139.495 ;
        RECT 87.045 138.995 87.215 139.245 ;
        RECT 87.045 138.825 87.985 138.995 ;
        RECT 88.355 138.885 88.620 139.245 ;
        RECT 86.505 138.105 86.965 138.655 ;
        RECT 87.155 137.935 87.485 138.655 ;
        RECT 87.685 138.275 87.985 138.825 ;
        RECT 88.155 137.935 88.435 138.605 ;
        RECT 88.805 137.935 89.095 139.100 ;
        RECT 89.725 139.025 90.935 139.545 ;
        RECT 91.105 139.195 92.315 139.715 ;
        RECT 92.505 139.215 92.835 139.585 ;
        RECT 93.070 139.510 93.240 139.765 ;
        RECT 93.070 139.180 93.355 139.510 ;
        RECT 93.070 139.035 93.240 139.180 ;
        RECT 89.725 137.935 92.315 139.025 ;
        RECT 92.575 138.865 93.240 139.035 ;
        RECT 93.525 139.010 93.695 139.810 ;
        RECT 93.955 139.935 94.125 140.315 ;
        RECT 94.305 140.105 94.635 140.485 ;
        RECT 93.955 139.765 94.620 139.935 ;
        RECT 94.815 139.810 95.075 140.315 ;
        RECT 93.885 139.215 94.215 139.585 ;
        RECT 94.450 139.510 94.620 139.765 ;
        RECT 94.450 139.180 94.735 139.510 ;
        RECT 94.450 139.035 94.620 139.180 ;
        RECT 92.575 138.105 92.745 138.865 ;
        RECT 92.925 137.935 93.255 138.695 ;
        RECT 93.425 138.105 93.695 139.010 ;
        RECT 93.955 138.865 94.620 139.035 ;
        RECT 94.905 139.010 95.075 139.810 ;
        RECT 95.305 139.665 95.515 140.485 ;
        RECT 95.685 139.685 96.015 140.315 ;
        RECT 95.685 139.085 95.935 139.685 ;
        RECT 96.185 139.665 96.415 140.485 ;
        RECT 97.285 139.855 97.615 140.215 ;
        RECT 98.235 140.025 98.485 140.485 ;
        RECT 98.655 140.025 99.215 140.315 ;
        RECT 97.285 139.665 98.675 139.855 ;
        RECT 98.505 139.575 98.675 139.665 ;
        RECT 96.105 139.245 96.435 139.495 ;
        RECT 97.100 139.245 97.775 139.495 ;
        RECT 97.995 139.245 98.335 139.495 ;
        RECT 98.505 139.245 98.795 139.575 ;
        RECT 93.955 138.105 94.125 138.865 ;
        RECT 94.305 137.935 94.635 138.695 ;
        RECT 94.805 138.105 95.075 139.010 ;
        RECT 95.305 137.935 95.515 139.075 ;
        RECT 95.685 138.105 96.015 139.085 ;
        RECT 96.185 137.935 96.415 139.075 ;
        RECT 97.100 138.885 97.365 139.245 ;
        RECT 98.505 138.995 98.675 139.245 ;
        RECT 97.735 138.825 98.675 138.995 ;
        RECT 97.285 137.935 97.565 138.605 ;
        RECT 97.735 138.275 98.035 138.825 ;
        RECT 98.965 138.655 99.215 140.025 ;
        RECT 99.905 140.015 100.205 140.485 ;
        RECT 100.375 139.845 100.630 140.290 ;
        RECT 100.800 140.015 101.060 140.485 ;
        RECT 101.230 139.845 101.490 140.290 ;
        RECT 101.660 140.015 101.955 140.485 ;
        RECT 99.385 139.675 102.415 139.845 ;
        RECT 102.605 139.735 103.815 140.485 ;
        RECT 99.385 139.110 99.685 139.675 ;
        RECT 99.860 139.280 102.075 139.505 ;
        RECT 102.245 139.110 102.415 139.675 ;
        RECT 99.385 138.940 102.415 139.110 ;
        RECT 102.605 139.025 103.125 139.565 ;
        RECT 103.295 139.195 103.815 139.735 ;
        RECT 104.185 139.855 104.515 140.215 ;
        RECT 105.135 140.025 105.385 140.485 ;
        RECT 105.555 140.025 106.115 140.315 ;
        RECT 104.185 139.665 105.575 139.855 ;
        RECT 105.405 139.575 105.575 139.665 ;
        RECT 104.000 139.245 104.675 139.495 ;
        RECT 104.895 139.245 105.235 139.495 ;
        RECT 105.405 139.245 105.695 139.575 ;
        RECT 98.235 137.935 98.565 138.655 ;
        RECT 98.755 138.105 99.215 138.655 ;
        RECT 99.385 137.935 99.770 138.770 ;
        RECT 99.940 138.135 100.200 138.940 ;
        RECT 100.370 137.935 100.630 138.770 ;
        RECT 100.800 138.135 101.055 138.940 ;
        RECT 101.230 137.935 101.490 138.770 ;
        RECT 101.660 138.135 101.915 138.940 ;
        RECT 102.090 137.935 102.435 138.770 ;
        RECT 102.605 137.935 103.815 139.025 ;
        RECT 104.000 138.885 104.265 139.245 ;
        RECT 105.405 138.995 105.575 139.245 ;
        RECT 104.635 138.825 105.575 138.995 ;
        RECT 104.185 137.935 104.465 138.605 ;
        RECT 104.635 138.275 104.935 138.825 ;
        RECT 105.865 138.655 106.115 140.025 ;
        RECT 106.485 139.855 106.815 140.215 ;
        RECT 107.435 140.025 107.685 140.485 ;
        RECT 107.855 140.025 108.415 140.315 ;
        RECT 106.485 139.665 107.875 139.855 ;
        RECT 107.705 139.575 107.875 139.665 ;
        RECT 106.300 139.245 106.975 139.495 ;
        RECT 107.195 139.245 107.535 139.495 ;
        RECT 107.705 139.245 107.995 139.575 ;
        RECT 106.300 138.885 106.565 139.245 ;
        RECT 107.705 138.995 107.875 139.245 ;
        RECT 105.135 137.935 105.465 138.655 ;
        RECT 105.655 138.105 106.115 138.655 ;
        RECT 106.935 138.825 107.875 138.995 ;
        RECT 106.485 137.935 106.765 138.605 ;
        RECT 106.935 138.275 107.235 138.825 ;
        RECT 108.165 138.655 108.415 140.025 ;
        RECT 108.860 139.675 109.105 140.280 ;
        RECT 109.325 139.950 109.835 140.485 ;
        RECT 107.435 137.935 107.765 138.655 ;
        RECT 107.955 138.105 108.415 138.655 ;
        RECT 108.585 139.505 109.815 139.675 ;
        RECT 108.585 138.695 108.925 139.505 ;
        RECT 109.095 138.940 109.845 139.130 ;
        RECT 108.585 138.285 109.100 138.695 ;
        RECT 109.335 137.935 109.505 138.695 ;
        RECT 109.675 138.275 109.845 138.940 ;
        RECT 110.015 138.955 110.205 140.315 ;
        RECT 110.375 139.805 110.650 140.315 ;
        RECT 110.840 139.950 111.370 140.315 ;
        RECT 111.795 140.085 112.125 140.485 ;
        RECT 111.195 139.915 111.370 139.950 ;
        RECT 110.375 139.635 110.655 139.805 ;
        RECT 110.375 139.155 110.650 139.635 ;
        RECT 110.855 138.955 111.025 139.755 ;
        RECT 110.015 138.785 111.025 138.955 ;
        RECT 111.195 139.745 112.125 139.915 ;
        RECT 112.295 139.745 112.550 140.315 ;
        RECT 111.195 138.615 111.365 139.745 ;
        RECT 111.955 139.575 112.125 139.745 ;
        RECT 110.240 138.445 111.365 138.615 ;
        RECT 111.535 139.245 111.730 139.575 ;
        RECT 111.955 139.245 112.210 139.575 ;
        RECT 111.535 138.275 111.705 139.245 ;
        RECT 112.380 139.075 112.550 139.745 ;
        RECT 112.725 139.715 114.395 140.485 ;
        RECT 114.565 139.760 114.855 140.485 ;
        RECT 115.025 139.715 116.695 140.485 ;
        RECT 109.675 138.105 111.705 138.275 ;
        RECT 111.875 137.935 112.045 139.075 ;
        RECT 112.215 138.105 112.550 139.075 ;
        RECT 112.725 139.025 113.475 139.545 ;
        RECT 113.645 139.195 114.395 139.715 ;
        RECT 112.725 137.935 114.395 139.025 ;
        RECT 114.565 137.935 114.855 139.100 ;
        RECT 115.025 139.025 115.775 139.545 ;
        RECT 115.945 139.195 116.695 139.715 ;
        RECT 117.240 139.775 117.495 140.305 ;
        RECT 117.675 140.025 117.960 140.485 ;
        RECT 115.025 137.935 116.695 139.025 ;
        RECT 117.240 138.915 117.420 139.775 ;
        RECT 118.140 139.575 118.390 140.225 ;
        RECT 117.590 139.245 118.390 139.575 ;
        RECT 117.240 138.785 117.495 138.915 ;
        RECT 117.155 138.615 117.495 138.785 ;
        RECT 117.240 138.245 117.495 138.615 ;
        RECT 117.675 137.935 117.960 138.735 ;
        RECT 118.140 138.655 118.390 139.245 ;
        RECT 118.590 139.890 118.910 140.220 ;
        RECT 119.090 140.005 119.750 140.485 ;
        RECT 119.950 140.095 120.800 140.265 ;
        RECT 118.590 138.995 118.780 139.890 ;
        RECT 119.100 139.565 119.760 139.835 ;
        RECT 119.430 139.505 119.760 139.565 ;
        RECT 118.950 139.335 119.280 139.395 ;
        RECT 119.950 139.335 120.120 140.095 ;
        RECT 121.360 140.025 121.680 140.485 ;
        RECT 121.880 139.845 122.130 140.275 ;
        RECT 122.420 140.045 122.830 140.485 ;
        RECT 123.000 140.105 124.015 140.305 ;
        RECT 120.290 139.675 121.540 139.845 ;
        RECT 120.290 139.555 120.620 139.675 ;
        RECT 118.950 139.165 120.850 139.335 ;
        RECT 118.590 138.825 120.510 138.995 ;
        RECT 118.590 138.805 118.910 138.825 ;
        RECT 118.140 138.145 118.470 138.655 ;
        RECT 118.740 138.195 118.910 138.805 ;
        RECT 120.680 138.655 120.850 139.165 ;
        RECT 121.020 139.095 121.200 139.505 ;
        RECT 121.370 138.915 121.540 139.675 ;
        RECT 119.080 137.935 119.410 138.625 ;
        RECT 119.640 138.485 120.850 138.655 ;
        RECT 121.020 138.605 121.540 138.915 ;
        RECT 121.710 139.505 122.130 139.845 ;
        RECT 122.420 139.505 122.830 139.835 ;
        RECT 121.710 138.735 121.900 139.505 ;
        RECT 123.000 139.375 123.170 140.105 ;
        RECT 124.315 139.935 124.485 140.265 ;
        RECT 124.655 140.105 124.985 140.485 ;
        RECT 123.340 139.555 123.690 139.925 ;
        RECT 123.000 139.335 123.420 139.375 ;
        RECT 122.070 139.165 123.420 139.335 ;
        RECT 122.070 139.005 122.320 139.165 ;
        RECT 122.830 138.735 123.080 138.995 ;
        RECT 121.710 138.485 123.080 138.735 ;
        RECT 119.640 138.195 119.880 138.485 ;
        RECT 120.680 138.405 120.850 138.485 ;
        RECT 120.080 137.935 120.500 138.315 ;
        RECT 120.680 138.155 121.310 138.405 ;
        RECT 121.780 137.935 122.110 138.315 ;
        RECT 122.280 138.195 122.450 138.485 ;
        RECT 123.250 138.320 123.420 139.165 ;
        RECT 123.870 138.995 124.090 139.865 ;
        RECT 124.315 139.745 125.010 139.935 ;
        RECT 123.590 138.615 124.090 138.995 ;
        RECT 124.260 138.945 124.670 139.565 ;
        RECT 124.840 138.775 125.010 139.745 ;
        RECT 124.315 138.605 125.010 138.775 ;
        RECT 122.630 137.935 123.010 138.315 ;
        RECT 123.250 138.150 124.080 138.320 ;
        RECT 124.315 138.105 124.485 138.605 ;
        RECT 124.655 137.935 124.985 138.435 ;
        RECT 125.200 138.105 125.425 140.225 ;
        RECT 125.595 140.105 125.925 140.485 ;
        RECT 126.095 139.935 126.265 140.225 ;
        RECT 125.600 139.765 126.265 139.935 ;
        RECT 125.600 138.775 125.830 139.765 ;
        RECT 126.525 139.735 127.735 140.485 ;
        RECT 126.000 138.945 126.350 139.595 ;
        RECT 126.525 139.025 127.045 139.565 ;
        RECT 127.215 139.195 127.735 139.735 ;
        RECT 125.600 138.605 126.265 138.775 ;
        RECT 125.595 137.935 125.925 138.435 ;
        RECT 126.095 138.105 126.265 138.605 ;
        RECT 126.525 137.935 127.735 139.025 ;
        RECT 29.840 137.765 127.820 137.935 ;
        RECT 29.925 136.675 31.135 137.765 ;
        RECT 29.925 135.965 30.445 136.505 ;
        RECT 30.615 136.135 31.135 136.675 ;
        RECT 31.765 136.675 33.435 137.765 ;
        RECT 33.610 137.330 38.955 137.765 ;
        RECT 31.765 136.155 32.515 136.675 ;
        RECT 32.685 135.985 33.435 136.505 ;
        RECT 35.200 136.080 35.550 137.330 ;
        RECT 39.165 136.625 39.395 137.765 ;
        RECT 39.565 136.615 39.895 137.595 ;
        RECT 40.065 136.625 40.275 137.765 ;
        RECT 40.880 137.425 41.135 137.455 ;
        RECT 40.795 137.255 41.135 137.425 ;
        RECT 40.880 136.785 41.135 137.255 ;
        RECT 41.315 136.965 41.600 137.765 ;
        RECT 41.780 137.045 42.110 137.555 ;
        RECT 29.925 135.215 31.135 135.965 ;
        RECT 31.765 135.215 33.435 135.985 ;
        RECT 37.030 135.760 37.370 136.590 ;
        RECT 39.145 136.205 39.475 136.455 ;
        RECT 33.610 135.215 38.955 135.760 ;
        RECT 39.165 135.215 39.395 136.035 ;
        RECT 39.645 136.015 39.895 136.615 ;
        RECT 39.565 135.385 39.895 136.015 ;
        RECT 40.065 135.215 40.275 136.035 ;
        RECT 40.880 135.925 41.060 136.785 ;
        RECT 41.780 136.455 42.030 137.045 ;
        RECT 42.380 136.895 42.550 137.505 ;
        RECT 42.720 137.075 43.050 137.765 ;
        RECT 43.280 137.215 43.520 137.505 ;
        RECT 43.720 137.385 44.140 137.765 ;
        RECT 44.320 137.295 44.950 137.545 ;
        RECT 45.420 137.385 45.750 137.765 ;
        RECT 44.320 137.215 44.490 137.295 ;
        RECT 45.920 137.215 46.090 137.505 ;
        RECT 46.270 137.385 46.650 137.765 ;
        RECT 46.890 137.380 47.720 137.550 ;
        RECT 43.280 137.045 44.490 137.215 ;
        RECT 41.230 136.125 42.030 136.455 ;
        RECT 40.880 135.395 41.135 135.925 ;
        RECT 41.315 135.215 41.600 135.675 ;
        RECT 41.780 135.475 42.030 136.125 ;
        RECT 42.230 136.875 42.550 136.895 ;
        RECT 42.230 136.705 44.150 136.875 ;
        RECT 42.230 135.810 42.420 136.705 ;
        RECT 44.320 136.535 44.490 137.045 ;
        RECT 44.660 136.785 45.180 137.095 ;
        RECT 42.590 136.365 44.490 136.535 ;
        RECT 42.590 136.305 42.920 136.365 ;
        RECT 43.070 136.135 43.400 136.195 ;
        RECT 42.740 135.865 43.400 136.135 ;
        RECT 42.230 135.480 42.550 135.810 ;
        RECT 42.730 135.215 43.390 135.695 ;
        RECT 43.590 135.605 43.760 136.365 ;
        RECT 44.660 136.195 44.840 136.605 ;
        RECT 43.930 136.025 44.260 136.145 ;
        RECT 45.010 136.025 45.180 136.785 ;
        RECT 43.930 135.855 45.180 136.025 ;
        RECT 45.350 136.965 46.720 137.215 ;
        RECT 45.350 136.195 45.540 136.965 ;
        RECT 46.470 136.705 46.720 136.965 ;
        RECT 45.710 136.535 45.960 136.695 ;
        RECT 46.890 136.535 47.060 137.380 ;
        RECT 47.955 137.095 48.125 137.595 ;
        RECT 48.295 137.265 48.625 137.765 ;
        RECT 47.230 136.705 47.730 137.085 ;
        RECT 47.955 136.925 48.650 137.095 ;
        RECT 45.710 136.365 47.060 136.535 ;
        RECT 46.640 136.325 47.060 136.365 ;
        RECT 45.350 135.855 45.770 136.195 ;
        RECT 46.060 135.865 46.470 136.195 ;
        RECT 43.590 135.435 44.440 135.605 ;
        RECT 45.000 135.215 45.320 135.675 ;
        RECT 45.520 135.425 45.770 135.855 ;
        RECT 46.060 135.215 46.470 135.655 ;
        RECT 46.640 135.595 46.810 136.325 ;
        RECT 46.980 135.775 47.330 136.145 ;
        RECT 47.510 135.835 47.730 136.705 ;
        RECT 47.900 136.135 48.310 136.755 ;
        RECT 48.480 135.955 48.650 136.925 ;
        RECT 47.955 135.765 48.650 135.955 ;
        RECT 46.640 135.395 47.655 135.595 ;
        RECT 47.955 135.435 48.125 135.765 ;
        RECT 48.295 135.215 48.625 135.595 ;
        RECT 48.840 135.475 49.065 137.595 ;
        RECT 49.235 137.265 49.565 137.765 ;
        RECT 49.735 137.095 49.905 137.595 ;
        RECT 49.240 136.925 49.905 137.095 ;
        RECT 49.240 135.935 49.470 136.925 ;
        RECT 49.640 136.105 49.990 136.755 ;
        RECT 50.165 136.600 50.455 137.765 ;
        RECT 50.625 137.005 51.140 137.415 ;
        RECT 51.375 137.005 51.545 137.765 ;
        RECT 51.715 137.425 53.745 137.595 ;
        RECT 50.625 136.195 50.965 137.005 ;
        RECT 51.715 136.760 51.885 137.425 ;
        RECT 52.280 137.085 53.405 137.255 ;
        RECT 51.135 136.570 51.885 136.760 ;
        RECT 52.055 136.745 53.065 136.915 ;
        RECT 50.625 136.025 51.855 136.195 ;
        RECT 49.240 135.765 49.905 135.935 ;
        RECT 49.235 135.215 49.565 135.595 ;
        RECT 49.735 135.475 49.905 135.765 ;
        RECT 50.165 135.215 50.455 135.940 ;
        RECT 50.900 135.420 51.145 136.025 ;
        RECT 51.365 135.215 51.875 135.750 ;
        RECT 52.055 135.385 52.245 136.745 ;
        RECT 52.415 136.405 52.690 136.545 ;
        RECT 52.415 136.235 52.695 136.405 ;
        RECT 52.415 135.385 52.690 136.235 ;
        RECT 52.895 135.945 53.065 136.745 ;
        RECT 53.235 135.955 53.405 137.085 ;
        RECT 53.575 136.455 53.745 137.425 ;
        RECT 53.915 136.625 54.085 137.765 ;
        RECT 54.255 136.625 54.590 137.595 ;
        RECT 55.425 137.095 55.705 137.765 ;
        RECT 55.875 136.875 56.175 137.425 ;
        RECT 56.375 137.045 56.705 137.765 ;
        RECT 56.895 137.045 57.355 137.595 ;
        RECT 53.575 136.125 53.770 136.455 ;
        RECT 53.995 136.125 54.250 136.455 ;
        RECT 53.995 135.955 54.165 136.125 ;
        RECT 54.420 135.955 54.590 136.625 ;
        RECT 55.240 136.455 55.505 136.815 ;
        RECT 55.875 136.705 56.815 136.875 ;
        RECT 56.645 136.455 56.815 136.705 ;
        RECT 55.240 136.205 55.915 136.455 ;
        RECT 56.135 136.205 56.475 136.455 ;
        RECT 56.645 136.125 56.935 136.455 ;
        RECT 56.645 136.035 56.815 136.125 ;
        RECT 53.235 135.785 54.165 135.955 ;
        RECT 53.235 135.750 53.410 135.785 ;
        RECT 52.880 135.385 53.410 135.750 ;
        RECT 53.835 135.215 54.165 135.615 ;
        RECT 54.335 135.385 54.590 135.955 ;
        RECT 55.425 135.845 56.815 136.035 ;
        RECT 55.425 135.485 55.755 135.845 ;
        RECT 57.105 135.675 57.355 137.045 ;
        RECT 57.615 137.020 57.885 137.765 ;
        RECT 58.515 137.760 64.790 137.765 ;
        RECT 58.055 136.850 58.345 137.590 ;
        RECT 58.515 137.035 58.770 137.760 ;
        RECT 58.955 136.865 59.215 137.590 ;
        RECT 59.385 137.035 59.630 137.760 ;
        RECT 59.815 136.865 60.075 137.590 ;
        RECT 60.245 137.035 60.490 137.760 ;
        RECT 60.675 136.865 60.935 137.590 ;
        RECT 61.105 137.035 61.350 137.760 ;
        RECT 61.520 136.865 61.780 137.590 ;
        RECT 61.950 137.035 62.210 137.760 ;
        RECT 62.380 136.865 62.640 137.590 ;
        RECT 62.810 137.035 63.070 137.760 ;
        RECT 63.240 136.865 63.500 137.590 ;
        RECT 63.670 137.035 63.930 137.760 ;
        RECT 64.100 136.865 64.360 137.590 ;
        RECT 64.530 136.965 64.790 137.760 ;
        RECT 58.955 136.850 64.360 136.865 ;
        RECT 57.615 136.625 64.360 136.850 ;
        RECT 57.615 136.065 58.780 136.625 ;
        RECT 64.960 136.455 65.210 137.590 ;
        RECT 65.390 136.955 65.650 137.765 ;
        RECT 65.825 136.455 66.070 137.595 ;
        RECT 66.250 136.955 66.545 137.765 ;
        RECT 66.725 136.675 70.235 137.765 ;
        RECT 70.405 137.005 70.920 137.415 ;
        RECT 71.155 137.005 71.325 137.765 ;
        RECT 71.495 137.425 73.525 137.595 ;
        RECT 58.950 136.205 66.070 136.455 ;
        RECT 57.585 136.035 58.780 136.065 ;
        RECT 57.585 135.895 64.360 136.035 ;
        RECT 57.615 135.865 64.360 135.895 ;
        RECT 56.375 135.215 56.625 135.675 ;
        RECT 56.795 135.385 57.355 135.675 ;
        RECT 57.615 135.215 57.915 135.695 ;
        RECT 58.085 135.410 58.345 135.865 ;
        RECT 58.515 135.215 58.775 135.695 ;
        RECT 58.955 135.410 59.215 135.865 ;
        RECT 59.385 135.215 59.635 135.695 ;
        RECT 59.815 135.410 60.075 135.865 ;
        RECT 60.245 135.215 60.495 135.695 ;
        RECT 60.675 135.410 60.935 135.865 ;
        RECT 61.105 135.215 61.350 135.695 ;
        RECT 61.520 135.410 61.795 135.865 ;
        RECT 61.965 135.215 62.210 135.695 ;
        RECT 62.380 135.410 62.640 135.865 ;
        RECT 62.810 135.215 63.070 135.695 ;
        RECT 63.240 135.410 63.500 135.865 ;
        RECT 63.670 135.215 63.930 135.695 ;
        RECT 64.100 135.410 64.360 135.865 ;
        RECT 64.530 135.215 64.790 135.775 ;
        RECT 64.960 135.395 65.210 136.205 ;
        RECT 65.390 135.215 65.650 135.740 ;
        RECT 65.820 135.395 66.070 136.205 ;
        RECT 66.240 135.895 66.555 136.455 ;
        RECT 66.725 136.155 68.415 136.675 ;
        RECT 68.585 135.985 70.235 136.505 ;
        RECT 70.405 136.195 70.745 137.005 ;
        RECT 71.495 136.760 71.665 137.425 ;
        RECT 72.060 137.085 73.185 137.255 ;
        RECT 70.915 136.570 71.665 136.760 ;
        RECT 71.835 136.745 72.845 136.915 ;
        RECT 70.405 136.025 71.635 136.195 ;
        RECT 66.250 135.215 66.555 135.725 ;
        RECT 66.725 135.215 70.235 135.985 ;
        RECT 70.680 135.420 70.925 136.025 ;
        RECT 71.145 135.215 71.655 135.750 ;
        RECT 71.835 135.385 72.025 136.745 ;
        RECT 72.195 136.405 72.470 136.545 ;
        RECT 72.195 136.235 72.475 136.405 ;
        RECT 72.195 135.385 72.470 136.235 ;
        RECT 72.675 135.945 72.845 136.745 ;
        RECT 73.015 135.955 73.185 137.085 ;
        RECT 73.355 136.455 73.525 137.425 ;
        RECT 73.695 136.625 73.865 137.765 ;
        RECT 74.035 136.625 74.370 137.595 ;
        RECT 73.355 136.125 73.550 136.455 ;
        RECT 73.775 136.125 74.030 136.455 ;
        RECT 73.775 135.955 73.945 136.125 ;
        RECT 74.200 135.955 74.370 136.625 ;
        RECT 74.545 136.675 75.755 137.765 ;
        RECT 74.545 136.135 75.065 136.675 ;
        RECT 75.925 136.600 76.215 137.765 ;
        RECT 76.845 136.675 80.355 137.765 ;
        RECT 80.525 137.045 80.985 137.595 ;
        RECT 81.175 137.045 81.505 137.765 ;
        RECT 75.235 135.965 75.755 136.505 ;
        RECT 76.845 136.155 78.535 136.675 ;
        RECT 78.705 135.985 80.355 136.505 ;
        RECT 73.015 135.785 73.945 135.955 ;
        RECT 73.015 135.750 73.190 135.785 ;
        RECT 72.660 135.385 73.190 135.750 ;
        RECT 73.615 135.215 73.945 135.615 ;
        RECT 74.115 135.385 74.370 135.955 ;
        RECT 74.545 135.215 75.755 135.965 ;
        RECT 75.925 135.215 76.215 135.940 ;
        RECT 76.845 135.215 80.355 135.985 ;
        RECT 80.525 135.675 80.775 137.045 ;
        RECT 81.705 136.875 82.005 137.425 ;
        RECT 82.175 137.095 82.455 137.765 ;
        RECT 81.065 136.705 82.005 136.875 ;
        RECT 82.825 137.045 83.285 137.595 ;
        RECT 83.475 137.045 83.805 137.765 ;
        RECT 81.065 136.455 81.235 136.705 ;
        RECT 82.375 136.455 82.640 136.815 ;
        RECT 80.945 136.125 81.235 136.455 ;
        RECT 81.405 136.205 81.745 136.455 ;
        RECT 81.965 136.205 82.640 136.455 ;
        RECT 81.065 136.035 81.235 136.125 ;
        RECT 81.065 135.845 82.455 136.035 ;
        RECT 80.525 135.385 81.085 135.675 ;
        RECT 81.255 135.215 81.505 135.675 ;
        RECT 82.125 135.485 82.455 135.845 ;
        RECT 82.825 135.675 83.075 137.045 ;
        RECT 84.005 136.875 84.305 137.425 ;
        RECT 84.475 137.095 84.755 137.765 ;
        RECT 83.365 136.705 84.305 136.875 ;
        RECT 85.125 137.045 85.585 137.595 ;
        RECT 85.775 137.045 86.105 137.765 ;
        RECT 83.365 136.455 83.535 136.705 ;
        RECT 84.675 136.455 84.940 136.815 ;
        RECT 83.245 136.125 83.535 136.455 ;
        RECT 83.705 136.205 84.045 136.455 ;
        RECT 84.265 136.205 84.940 136.455 ;
        RECT 83.365 136.035 83.535 136.125 ;
        RECT 83.365 135.845 84.755 136.035 ;
        RECT 82.825 135.385 83.385 135.675 ;
        RECT 83.555 135.215 83.805 135.675 ;
        RECT 84.425 135.485 84.755 135.845 ;
        RECT 85.125 135.675 85.375 137.045 ;
        RECT 86.305 136.875 86.605 137.425 ;
        RECT 86.775 137.095 87.055 137.765 ;
        RECT 87.895 136.955 88.190 137.765 ;
        RECT 85.665 136.705 86.605 136.875 ;
        RECT 85.665 136.455 85.835 136.705 ;
        RECT 86.975 136.455 87.240 136.815 ;
        RECT 88.370 136.455 88.615 137.595 ;
        RECT 88.790 136.955 89.050 137.765 ;
        RECT 89.650 137.760 95.925 137.765 ;
        RECT 89.230 136.455 89.480 137.590 ;
        RECT 89.650 136.965 89.910 137.760 ;
        RECT 90.080 136.865 90.340 137.590 ;
        RECT 90.510 137.035 90.770 137.760 ;
        RECT 90.940 136.865 91.200 137.590 ;
        RECT 91.370 137.035 91.630 137.760 ;
        RECT 91.800 136.865 92.060 137.590 ;
        RECT 92.230 137.035 92.490 137.760 ;
        RECT 92.660 136.865 92.920 137.590 ;
        RECT 93.090 137.035 93.335 137.760 ;
        RECT 93.505 136.865 93.765 137.590 ;
        RECT 93.950 137.035 94.195 137.760 ;
        RECT 94.365 136.865 94.625 137.590 ;
        RECT 94.810 137.035 95.055 137.760 ;
        RECT 95.225 136.865 95.485 137.590 ;
        RECT 95.670 137.035 95.925 137.760 ;
        RECT 90.080 136.850 95.485 136.865 ;
        RECT 96.095 136.850 96.385 137.590 ;
        RECT 96.555 137.020 96.825 137.765 ;
        RECT 97.085 137.005 97.600 137.415 ;
        RECT 97.835 137.005 98.005 137.765 ;
        RECT 98.175 137.425 100.205 137.595 ;
        RECT 90.080 136.625 96.825 136.850 ;
        RECT 85.545 136.125 85.835 136.455 ;
        RECT 86.005 136.205 86.345 136.455 ;
        RECT 86.565 136.205 87.240 136.455 ;
        RECT 85.665 136.035 85.835 136.125 ;
        RECT 85.665 135.845 87.055 136.035 ;
        RECT 87.885 135.895 88.200 136.455 ;
        RECT 88.370 136.205 95.490 136.455 ;
        RECT 85.125 135.385 85.685 135.675 ;
        RECT 85.855 135.215 86.105 135.675 ;
        RECT 86.725 135.485 87.055 135.845 ;
        RECT 87.885 135.215 88.190 135.725 ;
        RECT 88.370 135.395 88.620 136.205 ;
        RECT 88.790 135.215 89.050 135.740 ;
        RECT 89.230 135.395 89.480 136.205 ;
        RECT 95.660 136.035 96.825 136.625 ;
        RECT 90.080 135.865 96.825 136.035 ;
        RECT 97.085 136.195 97.425 137.005 ;
        RECT 98.175 136.760 98.345 137.425 ;
        RECT 98.740 137.085 99.865 137.255 ;
        RECT 97.595 136.570 98.345 136.760 ;
        RECT 98.515 136.745 99.525 136.915 ;
        RECT 97.085 136.025 98.315 136.195 ;
        RECT 89.650 135.215 89.910 135.775 ;
        RECT 90.080 135.410 90.340 135.865 ;
        RECT 90.510 135.215 90.770 135.695 ;
        RECT 90.940 135.410 91.200 135.865 ;
        RECT 91.370 135.215 91.630 135.695 ;
        RECT 91.800 135.410 92.060 135.865 ;
        RECT 92.230 135.215 92.475 135.695 ;
        RECT 92.645 135.410 92.920 135.865 ;
        RECT 93.090 135.215 93.335 135.695 ;
        RECT 93.505 135.410 93.765 135.865 ;
        RECT 93.945 135.215 94.195 135.695 ;
        RECT 94.365 135.410 94.625 135.865 ;
        RECT 94.805 135.215 95.055 135.695 ;
        RECT 95.225 135.410 95.485 135.865 ;
        RECT 95.665 135.215 95.925 135.695 ;
        RECT 96.095 135.410 96.355 135.865 ;
        RECT 96.525 135.215 96.825 135.695 ;
        RECT 97.360 135.420 97.605 136.025 ;
        RECT 97.825 135.215 98.335 135.750 ;
        RECT 98.515 135.385 98.705 136.745 ;
        RECT 98.875 136.405 99.150 136.545 ;
        RECT 98.875 136.235 99.155 136.405 ;
        RECT 98.875 135.385 99.150 136.235 ;
        RECT 99.355 135.945 99.525 136.745 ;
        RECT 99.695 135.955 99.865 137.085 ;
        RECT 100.035 136.455 100.205 137.425 ;
        RECT 100.375 136.625 100.545 137.765 ;
        RECT 100.715 136.625 101.050 137.595 ;
        RECT 100.035 136.125 100.230 136.455 ;
        RECT 100.455 136.125 100.710 136.455 ;
        RECT 100.455 135.955 100.625 136.125 ;
        RECT 100.880 135.955 101.050 136.625 ;
        RECT 101.685 136.600 101.975 137.765 ;
        RECT 102.185 136.625 102.415 137.765 ;
        RECT 102.585 136.615 102.915 137.595 ;
        RECT 103.085 136.625 103.295 137.765 ;
        RECT 103.900 136.785 104.155 137.455 ;
        RECT 104.335 136.965 104.620 137.765 ;
        RECT 104.800 137.045 105.130 137.555 ;
        RECT 102.165 136.205 102.495 136.455 ;
        RECT 99.695 135.785 100.625 135.955 ;
        RECT 99.695 135.750 99.870 135.785 ;
        RECT 99.340 135.385 99.870 135.750 ;
        RECT 100.295 135.215 100.625 135.615 ;
        RECT 100.795 135.385 101.050 135.955 ;
        RECT 101.685 135.215 101.975 135.940 ;
        RECT 102.185 135.215 102.415 136.035 ;
        RECT 102.665 136.015 102.915 136.615 ;
        RECT 102.585 135.385 102.915 136.015 ;
        RECT 103.085 135.215 103.295 136.035 ;
        RECT 103.900 135.925 104.080 136.785 ;
        RECT 104.800 136.455 105.050 137.045 ;
        RECT 105.400 136.895 105.570 137.505 ;
        RECT 105.740 137.075 106.070 137.765 ;
        RECT 106.300 137.215 106.540 137.505 ;
        RECT 106.740 137.385 107.160 137.765 ;
        RECT 107.340 137.295 107.970 137.545 ;
        RECT 108.440 137.385 108.770 137.765 ;
        RECT 107.340 137.215 107.510 137.295 ;
        RECT 108.940 137.215 109.110 137.505 ;
        RECT 109.290 137.385 109.670 137.765 ;
        RECT 109.910 137.380 110.740 137.550 ;
        RECT 106.300 137.045 107.510 137.215 ;
        RECT 104.250 136.125 105.050 136.455 ;
        RECT 103.900 135.725 104.155 135.925 ;
        RECT 103.815 135.555 104.155 135.725 ;
        RECT 103.900 135.395 104.155 135.555 ;
        RECT 104.335 135.215 104.620 135.675 ;
        RECT 104.800 135.475 105.050 136.125 ;
        RECT 105.250 136.875 105.570 136.895 ;
        RECT 105.250 136.705 107.170 136.875 ;
        RECT 105.250 135.810 105.440 136.705 ;
        RECT 107.340 136.535 107.510 137.045 ;
        RECT 107.680 136.785 108.200 137.095 ;
        RECT 105.610 136.365 107.510 136.535 ;
        RECT 105.610 136.305 105.940 136.365 ;
        RECT 106.090 136.135 106.420 136.195 ;
        RECT 105.760 135.865 106.420 136.135 ;
        RECT 105.250 135.480 105.570 135.810 ;
        RECT 105.750 135.215 106.410 135.695 ;
        RECT 106.610 135.605 106.780 136.365 ;
        RECT 107.680 136.195 107.860 136.605 ;
        RECT 106.950 136.025 107.280 136.145 ;
        RECT 108.030 136.025 108.200 136.785 ;
        RECT 106.950 135.855 108.200 136.025 ;
        RECT 108.370 136.965 109.740 137.215 ;
        RECT 108.370 136.195 108.560 136.965 ;
        RECT 109.490 136.705 109.740 136.965 ;
        RECT 108.730 136.535 108.980 136.695 ;
        RECT 109.910 136.535 110.080 137.380 ;
        RECT 110.975 137.095 111.145 137.595 ;
        RECT 111.315 137.265 111.645 137.765 ;
        RECT 110.250 136.705 110.750 137.085 ;
        RECT 110.975 136.925 111.670 137.095 ;
        RECT 108.730 136.365 110.080 136.535 ;
        RECT 109.660 136.325 110.080 136.365 ;
        RECT 108.370 135.855 108.790 136.195 ;
        RECT 109.080 135.865 109.490 136.195 ;
        RECT 106.610 135.435 107.460 135.605 ;
        RECT 108.020 135.215 108.340 135.675 ;
        RECT 108.540 135.425 108.790 135.855 ;
        RECT 109.080 135.215 109.490 135.655 ;
        RECT 109.660 135.595 109.830 136.325 ;
        RECT 110.000 135.775 110.350 136.145 ;
        RECT 110.530 135.835 110.750 136.705 ;
        RECT 110.920 136.135 111.330 136.755 ;
        RECT 111.500 135.955 111.670 136.925 ;
        RECT 110.975 135.765 111.670 135.955 ;
        RECT 109.660 135.395 110.675 135.595 ;
        RECT 110.975 135.435 111.145 135.765 ;
        RECT 111.315 135.215 111.645 135.595 ;
        RECT 111.860 135.475 112.085 137.595 ;
        RECT 112.255 137.265 112.585 137.765 ;
        RECT 112.755 137.095 112.925 137.595 ;
        RECT 112.260 136.925 112.925 137.095 ;
        RECT 112.260 135.935 112.490 136.925 ;
        RECT 112.660 136.105 113.010 136.755 ;
        RECT 113.185 136.690 113.455 137.595 ;
        RECT 113.625 137.005 113.955 137.765 ;
        RECT 114.135 136.835 114.305 137.595 ;
        RECT 112.260 135.765 112.925 135.935 ;
        RECT 112.255 135.215 112.585 135.595 ;
        RECT 112.755 135.475 112.925 135.765 ;
        RECT 113.185 135.890 113.355 136.690 ;
        RECT 113.640 136.665 114.305 136.835 ;
        RECT 113.640 136.520 113.810 136.665 ;
        RECT 114.605 136.625 114.835 137.765 ;
        RECT 115.005 136.615 115.335 137.595 ;
        RECT 115.505 136.625 115.715 137.765 ;
        RECT 116.320 136.785 116.575 137.455 ;
        RECT 116.755 136.965 117.040 137.765 ;
        RECT 117.220 137.045 117.550 137.555 ;
        RECT 113.525 136.190 113.810 136.520 ;
        RECT 113.640 135.935 113.810 136.190 ;
        RECT 114.045 136.115 114.375 136.485 ;
        RECT 114.585 136.205 114.915 136.455 ;
        RECT 113.185 135.385 113.445 135.890 ;
        RECT 113.640 135.765 114.305 135.935 ;
        RECT 113.625 135.215 113.955 135.595 ;
        RECT 114.135 135.385 114.305 135.765 ;
        RECT 114.605 135.215 114.835 136.035 ;
        RECT 115.085 136.015 115.335 136.615 ;
        RECT 115.005 135.385 115.335 136.015 ;
        RECT 115.505 135.215 115.715 136.035 ;
        RECT 116.320 135.925 116.500 136.785 ;
        RECT 117.220 136.455 117.470 137.045 ;
        RECT 117.820 136.895 117.990 137.505 ;
        RECT 118.160 137.075 118.490 137.765 ;
        RECT 118.720 137.215 118.960 137.505 ;
        RECT 119.160 137.385 119.580 137.765 ;
        RECT 119.760 137.295 120.390 137.545 ;
        RECT 120.860 137.385 121.190 137.765 ;
        RECT 119.760 137.215 119.930 137.295 ;
        RECT 121.360 137.215 121.530 137.505 ;
        RECT 121.710 137.385 122.090 137.765 ;
        RECT 122.330 137.380 123.160 137.550 ;
        RECT 118.720 137.045 119.930 137.215 ;
        RECT 116.670 136.125 117.470 136.455 ;
        RECT 116.320 135.725 116.575 135.925 ;
        RECT 116.235 135.555 116.575 135.725 ;
        RECT 116.320 135.395 116.575 135.555 ;
        RECT 116.755 135.215 117.040 135.675 ;
        RECT 117.220 135.475 117.470 136.125 ;
        RECT 117.670 136.875 117.990 136.895 ;
        RECT 117.670 136.705 119.590 136.875 ;
        RECT 117.670 135.810 117.860 136.705 ;
        RECT 119.760 136.535 119.930 137.045 ;
        RECT 120.100 136.785 120.620 137.095 ;
        RECT 118.030 136.365 119.930 136.535 ;
        RECT 118.030 136.305 118.360 136.365 ;
        RECT 118.510 136.135 118.840 136.195 ;
        RECT 118.180 135.865 118.840 136.135 ;
        RECT 117.670 135.480 117.990 135.810 ;
        RECT 118.170 135.215 118.830 135.695 ;
        RECT 119.030 135.605 119.200 136.365 ;
        RECT 120.100 136.195 120.280 136.605 ;
        RECT 119.370 136.025 119.700 136.145 ;
        RECT 120.450 136.025 120.620 136.785 ;
        RECT 119.370 135.855 120.620 136.025 ;
        RECT 120.790 136.965 122.160 137.215 ;
        RECT 120.790 136.195 120.980 136.965 ;
        RECT 121.910 136.705 122.160 136.965 ;
        RECT 121.150 136.535 121.400 136.695 ;
        RECT 122.330 136.535 122.500 137.380 ;
        RECT 123.395 137.095 123.565 137.595 ;
        RECT 123.735 137.265 124.065 137.765 ;
        RECT 122.670 136.705 123.170 137.085 ;
        RECT 123.395 136.925 124.090 137.095 ;
        RECT 121.150 136.365 122.500 136.535 ;
        RECT 122.080 136.325 122.500 136.365 ;
        RECT 120.790 135.855 121.210 136.195 ;
        RECT 121.500 135.865 121.910 136.195 ;
        RECT 119.030 135.435 119.880 135.605 ;
        RECT 120.440 135.215 120.760 135.675 ;
        RECT 120.960 135.425 121.210 135.855 ;
        RECT 121.500 135.215 121.910 135.655 ;
        RECT 122.080 135.595 122.250 136.325 ;
        RECT 122.420 135.775 122.770 136.145 ;
        RECT 122.950 135.835 123.170 136.705 ;
        RECT 123.340 136.135 123.750 136.755 ;
        RECT 123.920 135.955 124.090 136.925 ;
        RECT 123.395 135.765 124.090 135.955 ;
        RECT 122.080 135.395 123.095 135.595 ;
        RECT 123.395 135.435 123.565 135.765 ;
        RECT 123.735 135.215 124.065 135.595 ;
        RECT 124.280 135.475 124.505 137.595 ;
        RECT 124.675 137.265 125.005 137.765 ;
        RECT 125.175 137.095 125.345 137.595 ;
        RECT 124.680 136.925 125.345 137.095 ;
        RECT 124.680 135.935 124.910 136.925 ;
        RECT 125.080 136.105 125.430 136.755 ;
        RECT 126.525 136.675 127.735 137.765 ;
        RECT 126.525 136.135 127.045 136.675 ;
        RECT 127.215 135.965 127.735 136.505 ;
        RECT 124.680 135.765 125.345 135.935 ;
        RECT 124.675 135.215 125.005 135.595 ;
        RECT 125.175 135.475 125.345 135.765 ;
        RECT 126.525 135.215 127.735 135.965 ;
        RECT 29.840 135.045 127.820 135.215 ;
        RECT 29.925 134.295 31.135 135.045 ;
        RECT 29.925 133.755 30.445 134.295 ;
        RECT 31.305 134.275 32.975 135.045 ;
        RECT 30.615 133.585 31.135 134.125 ;
        RECT 29.925 132.495 31.135 133.585 ;
        RECT 31.305 133.585 32.055 134.105 ;
        RECT 32.225 133.755 32.975 134.275 ;
        RECT 33.150 134.305 33.405 134.875 ;
        RECT 33.575 134.645 33.905 135.045 ;
        RECT 34.330 134.510 34.860 134.875 ;
        RECT 35.050 134.705 35.325 134.875 ;
        RECT 35.045 134.535 35.325 134.705 ;
        RECT 34.330 134.475 34.505 134.510 ;
        RECT 33.575 134.305 34.505 134.475 ;
        RECT 33.150 133.635 33.320 134.305 ;
        RECT 33.575 134.135 33.745 134.305 ;
        RECT 33.490 133.805 33.745 134.135 ;
        RECT 33.970 133.805 34.165 134.135 ;
        RECT 31.305 132.495 32.975 133.585 ;
        RECT 33.150 132.665 33.485 133.635 ;
        RECT 33.655 132.495 33.825 133.635 ;
        RECT 33.995 132.835 34.165 133.805 ;
        RECT 34.335 133.175 34.505 134.305 ;
        RECT 34.675 133.515 34.845 134.315 ;
        RECT 35.050 133.715 35.325 134.535 ;
        RECT 35.495 133.515 35.685 134.875 ;
        RECT 35.865 134.510 36.375 135.045 ;
        RECT 36.595 134.235 36.840 134.840 ;
        RECT 37.285 134.320 37.575 135.045 ;
        RECT 37.835 134.495 38.005 134.785 ;
        RECT 38.175 134.665 38.505 135.045 ;
        RECT 37.835 134.325 38.500 134.495 ;
        RECT 35.885 134.065 37.115 134.235 ;
        RECT 34.675 133.345 35.685 133.515 ;
        RECT 35.855 133.500 36.605 133.690 ;
        RECT 34.335 133.005 35.460 133.175 ;
        RECT 35.855 132.835 36.025 133.500 ;
        RECT 36.775 133.255 37.115 134.065 ;
        RECT 33.995 132.665 36.025 132.835 ;
        RECT 36.195 132.495 36.365 133.255 ;
        RECT 36.600 132.845 37.115 133.255 ;
        RECT 37.285 132.495 37.575 133.660 ;
        RECT 37.750 133.505 38.100 134.155 ;
        RECT 38.270 133.335 38.500 134.325 ;
        RECT 37.835 133.165 38.500 133.335 ;
        RECT 37.835 132.665 38.005 133.165 ;
        RECT 38.175 132.495 38.505 132.995 ;
        RECT 38.675 132.665 38.900 134.785 ;
        RECT 39.115 134.665 39.445 135.045 ;
        RECT 39.615 134.495 39.785 134.825 ;
        RECT 40.085 134.665 41.100 134.865 ;
        RECT 39.090 134.305 39.785 134.495 ;
        RECT 39.090 133.335 39.260 134.305 ;
        RECT 39.430 133.505 39.840 134.125 ;
        RECT 40.010 133.555 40.230 134.425 ;
        RECT 40.410 134.115 40.760 134.485 ;
        RECT 40.930 133.935 41.100 134.665 ;
        RECT 41.270 134.605 41.680 135.045 ;
        RECT 41.970 134.405 42.220 134.835 ;
        RECT 42.420 134.585 42.740 135.045 ;
        RECT 43.300 134.655 44.150 134.825 ;
        RECT 41.270 134.065 41.680 134.395 ;
        RECT 41.970 134.065 42.390 134.405 ;
        RECT 40.680 133.895 41.100 133.935 ;
        RECT 40.680 133.725 42.030 133.895 ;
        RECT 39.090 133.165 39.785 133.335 ;
        RECT 40.010 133.175 40.510 133.555 ;
        RECT 39.115 132.495 39.445 132.995 ;
        RECT 39.615 132.665 39.785 133.165 ;
        RECT 40.680 132.880 40.850 133.725 ;
        RECT 41.780 133.565 42.030 133.725 ;
        RECT 41.020 133.295 41.270 133.555 ;
        RECT 42.200 133.295 42.390 134.065 ;
        RECT 41.020 133.045 42.390 133.295 ;
        RECT 42.560 134.235 43.810 134.405 ;
        RECT 42.560 133.475 42.730 134.235 ;
        RECT 43.480 134.115 43.810 134.235 ;
        RECT 42.900 133.655 43.080 134.065 ;
        RECT 43.980 133.895 44.150 134.655 ;
        RECT 44.350 134.565 45.010 135.045 ;
        RECT 45.190 134.450 45.510 134.780 ;
        RECT 44.340 134.125 45.000 134.395 ;
        RECT 44.340 134.065 44.670 134.125 ;
        RECT 44.820 133.895 45.150 133.955 ;
        RECT 43.250 133.725 45.150 133.895 ;
        RECT 42.560 133.165 43.080 133.475 ;
        RECT 43.250 133.215 43.420 133.725 ;
        RECT 45.320 133.555 45.510 134.450 ;
        RECT 43.590 133.385 45.510 133.555 ;
        RECT 45.190 133.365 45.510 133.385 ;
        RECT 45.710 134.135 45.960 134.785 ;
        RECT 46.140 134.585 46.425 135.045 ;
        RECT 46.605 134.705 46.860 134.865 ;
        RECT 46.605 134.535 46.945 134.705 ;
        RECT 46.605 134.335 46.860 134.535 ;
        RECT 45.710 133.805 46.510 134.135 ;
        RECT 43.250 133.045 44.460 133.215 ;
        RECT 40.020 132.710 40.850 132.880 ;
        RECT 41.090 132.495 41.470 132.875 ;
        RECT 41.650 132.755 41.820 133.045 ;
        RECT 43.250 132.965 43.420 133.045 ;
        RECT 41.990 132.495 42.320 132.875 ;
        RECT 42.790 132.715 43.420 132.965 ;
        RECT 43.600 132.495 44.020 132.875 ;
        RECT 44.220 132.755 44.460 133.045 ;
        RECT 44.690 132.495 45.020 133.185 ;
        RECT 45.190 132.755 45.360 133.365 ;
        RECT 45.710 133.215 45.960 133.805 ;
        RECT 46.680 133.475 46.860 134.335 ;
        RECT 47.495 134.495 47.665 134.785 ;
        RECT 47.835 134.665 48.165 135.045 ;
        RECT 47.495 134.325 48.160 134.495 ;
        RECT 47.410 133.505 47.760 134.155 ;
        RECT 45.630 132.705 45.960 133.215 ;
        RECT 46.140 132.495 46.425 133.295 ;
        RECT 46.605 132.805 46.860 133.475 ;
        RECT 47.930 133.335 48.160 134.325 ;
        RECT 47.495 133.165 48.160 133.335 ;
        RECT 47.495 132.665 47.665 133.165 ;
        RECT 47.835 132.495 48.165 132.995 ;
        RECT 48.335 132.665 48.560 134.785 ;
        RECT 48.775 134.665 49.105 135.045 ;
        RECT 49.275 134.495 49.445 134.825 ;
        RECT 49.745 134.665 50.760 134.865 ;
        RECT 48.750 134.305 49.445 134.495 ;
        RECT 48.750 133.335 48.920 134.305 ;
        RECT 49.090 133.505 49.500 134.125 ;
        RECT 49.670 133.555 49.890 134.425 ;
        RECT 50.070 134.115 50.420 134.485 ;
        RECT 50.590 133.935 50.760 134.665 ;
        RECT 50.930 134.605 51.340 135.045 ;
        RECT 51.630 134.405 51.880 134.835 ;
        RECT 52.080 134.585 52.400 135.045 ;
        RECT 52.960 134.655 53.810 134.825 ;
        RECT 50.930 134.065 51.340 134.395 ;
        RECT 51.630 134.065 52.050 134.405 ;
        RECT 50.340 133.895 50.760 133.935 ;
        RECT 50.340 133.725 51.690 133.895 ;
        RECT 48.750 133.165 49.445 133.335 ;
        RECT 49.670 133.175 50.170 133.555 ;
        RECT 48.775 132.495 49.105 132.995 ;
        RECT 49.275 132.665 49.445 133.165 ;
        RECT 50.340 132.880 50.510 133.725 ;
        RECT 51.440 133.565 51.690 133.725 ;
        RECT 50.680 133.295 50.930 133.555 ;
        RECT 51.860 133.295 52.050 134.065 ;
        RECT 50.680 133.045 52.050 133.295 ;
        RECT 52.220 134.235 53.470 134.405 ;
        RECT 52.220 133.475 52.390 134.235 ;
        RECT 53.140 134.115 53.470 134.235 ;
        RECT 52.560 133.655 52.740 134.065 ;
        RECT 53.640 133.895 53.810 134.655 ;
        RECT 54.010 134.565 54.670 135.045 ;
        RECT 54.850 134.450 55.170 134.780 ;
        RECT 54.000 134.125 54.660 134.395 ;
        RECT 54.000 134.065 54.330 134.125 ;
        RECT 54.480 133.895 54.810 133.955 ;
        RECT 52.910 133.725 54.810 133.895 ;
        RECT 52.220 133.165 52.740 133.475 ;
        RECT 52.910 133.215 53.080 133.725 ;
        RECT 54.980 133.555 55.170 134.450 ;
        RECT 53.250 133.385 55.170 133.555 ;
        RECT 54.850 133.365 55.170 133.385 ;
        RECT 55.370 134.135 55.620 134.785 ;
        RECT 55.800 134.585 56.085 135.045 ;
        RECT 56.265 134.705 56.520 134.865 ;
        RECT 56.265 134.535 56.605 134.705 ;
        RECT 56.265 134.335 56.520 134.535 ;
        RECT 55.370 133.805 56.170 134.135 ;
        RECT 52.910 133.045 54.120 133.215 ;
        RECT 49.680 132.710 50.510 132.880 ;
        RECT 50.750 132.495 51.130 132.875 ;
        RECT 51.310 132.755 51.480 133.045 ;
        RECT 52.910 132.965 53.080 133.045 ;
        RECT 51.650 132.495 51.980 132.875 ;
        RECT 52.450 132.715 53.080 132.965 ;
        RECT 53.260 132.495 53.680 132.875 ;
        RECT 53.880 132.755 54.120 133.045 ;
        RECT 54.350 132.495 54.680 133.185 ;
        RECT 54.850 132.755 55.020 133.365 ;
        RECT 55.370 133.215 55.620 133.805 ;
        RECT 56.340 133.475 56.520 134.335 ;
        RECT 58.185 134.415 58.515 134.775 ;
        RECT 59.135 134.585 59.385 135.045 ;
        RECT 59.555 134.585 60.115 134.875 ;
        RECT 58.185 134.225 59.575 134.415 ;
        RECT 59.405 134.135 59.575 134.225 ;
        RECT 55.290 132.705 55.620 133.215 ;
        RECT 55.800 132.495 56.085 133.295 ;
        RECT 56.265 132.805 56.520 133.475 ;
        RECT 58.000 133.805 58.675 134.055 ;
        RECT 58.895 133.805 59.235 134.055 ;
        RECT 59.405 133.805 59.695 134.135 ;
        RECT 58.000 133.445 58.265 133.805 ;
        RECT 59.405 133.555 59.575 133.805 ;
        RECT 58.635 133.385 59.575 133.555 ;
        RECT 58.185 132.495 58.465 133.165 ;
        RECT 58.635 132.835 58.935 133.385 ;
        RECT 59.865 133.215 60.115 134.585 ;
        RECT 60.295 134.545 60.625 135.045 ;
        RECT 60.825 134.475 60.995 134.825 ;
        RECT 61.195 134.645 61.525 135.045 ;
        RECT 61.695 134.475 61.865 134.825 ;
        RECT 62.035 134.645 62.415 135.045 ;
        RECT 60.290 133.805 60.640 134.375 ;
        RECT 60.825 134.305 62.435 134.475 ;
        RECT 62.605 134.370 62.875 134.715 ;
        RECT 62.265 134.135 62.435 134.305 ;
        RECT 60.810 133.685 61.520 134.135 ;
        RECT 61.690 133.805 62.095 134.135 ;
        RECT 62.265 133.805 62.535 134.135 ;
        RECT 59.135 132.495 59.465 133.215 ;
        RECT 59.655 132.665 60.115 133.215 ;
        RECT 60.290 133.345 60.610 133.635 ;
        RECT 60.805 133.515 61.520 133.685 ;
        RECT 62.265 133.635 62.435 133.805 ;
        RECT 62.705 133.635 62.875 134.370 ;
        RECT 63.045 134.320 63.335 135.045 ;
        RECT 63.965 134.245 64.305 134.875 ;
        RECT 64.475 134.245 64.725 135.045 ;
        RECT 64.915 134.395 65.245 134.875 ;
        RECT 65.415 134.585 65.640 135.045 ;
        RECT 65.810 134.395 66.140 134.875 ;
        RECT 61.710 133.465 62.435 133.635 ;
        RECT 61.710 133.345 61.880 133.465 ;
        RECT 60.290 133.175 61.880 133.345 ;
        RECT 60.290 132.715 61.945 133.005 ;
        RECT 62.115 132.495 62.395 133.295 ;
        RECT 62.605 132.665 62.875 133.635 ;
        RECT 63.045 132.495 63.335 133.660 ;
        RECT 63.965 133.635 64.140 134.245 ;
        RECT 64.915 134.225 66.140 134.395 ;
        RECT 66.770 134.265 67.270 134.875 ;
        RECT 64.310 133.885 65.005 134.055 ;
        RECT 64.835 133.635 65.005 133.885 ;
        RECT 65.180 133.855 65.600 134.055 ;
        RECT 65.770 133.855 66.100 134.055 ;
        RECT 66.270 133.855 66.600 134.055 ;
        RECT 66.770 133.635 66.940 134.265 ;
        RECT 67.685 134.225 67.915 135.045 ;
        RECT 68.085 134.245 68.415 134.875 ;
        RECT 67.125 133.805 67.475 134.055 ;
        RECT 67.665 133.805 67.995 134.055 ;
        RECT 68.165 133.645 68.415 134.245 ;
        RECT 68.585 134.225 68.795 135.045 ;
        RECT 69.300 134.235 69.545 134.840 ;
        RECT 69.765 134.510 70.275 135.045 ;
        RECT 63.965 132.665 64.305 133.635 ;
        RECT 64.475 132.495 64.645 133.635 ;
        RECT 64.835 133.465 67.270 133.635 ;
        RECT 64.915 132.495 65.165 133.295 ;
        RECT 65.810 132.665 66.140 133.465 ;
        RECT 66.440 132.495 66.770 133.295 ;
        RECT 66.940 132.665 67.270 133.465 ;
        RECT 67.685 132.495 67.915 133.635 ;
        RECT 68.085 132.665 68.415 133.645 ;
        RECT 69.025 134.065 70.255 134.235 ;
        RECT 68.585 132.495 68.795 133.635 ;
        RECT 69.025 133.255 69.365 134.065 ;
        RECT 69.535 133.500 70.285 133.690 ;
        RECT 69.025 132.845 69.540 133.255 ;
        RECT 69.775 132.495 69.945 133.255 ;
        RECT 70.115 132.835 70.285 133.500 ;
        RECT 70.455 133.515 70.645 134.875 ;
        RECT 70.815 134.025 71.090 134.875 ;
        RECT 71.280 134.510 71.810 134.875 ;
        RECT 72.235 134.645 72.565 135.045 ;
        RECT 71.635 134.475 71.810 134.510 ;
        RECT 70.815 133.855 71.095 134.025 ;
        RECT 70.815 133.715 71.090 133.855 ;
        RECT 71.295 133.515 71.465 134.315 ;
        RECT 70.455 133.345 71.465 133.515 ;
        RECT 71.635 134.305 72.565 134.475 ;
        RECT 72.735 134.305 72.990 134.875 ;
        RECT 71.635 133.175 71.805 134.305 ;
        RECT 72.395 134.135 72.565 134.305 ;
        RECT 70.680 133.005 71.805 133.175 ;
        RECT 71.975 133.805 72.170 134.135 ;
        RECT 72.395 133.805 72.650 134.135 ;
        RECT 71.975 132.835 72.145 133.805 ;
        RECT 72.820 133.635 72.990 134.305 ;
        RECT 73.225 134.225 73.435 135.045 ;
        RECT 73.605 134.245 73.935 134.875 ;
        RECT 73.605 133.645 73.855 134.245 ;
        RECT 74.105 134.225 74.335 135.045 ;
        RECT 74.545 134.370 74.805 134.875 ;
        RECT 74.985 134.665 75.315 135.045 ;
        RECT 75.495 134.495 75.665 134.875 ;
        RECT 74.025 133.805 74.355 134.055 ;
        RECT 70.115 132.665 72.145 132.835 ;
        RECT 72.315 132.495 72.485 133.635 ;
        RECT 72.655 132.665 72.990 133.635 ;
        RECT 73.225 132.495 73.435 133.635 ;
        RECT 73.605 132.665 73.935 133.645 ;
        RECT 74.105 132.495 74.335 133.635 ;
        RECT 74.545 133.570 74.715 134.370 ;
        RECT 75.000 134.325 75.665 134.495 ;
        RECT 75.000 134.070 75.170 134.325 ;
        RECT 76.845 134.275 80.355 135.045 ;
        RECT 74.885 133.740 75.170 134.070 ;
        RECT 75.405 133.775 75.735 134.145 ;
        RECT 75.000 133.595 75.170 133.740 ;
        RECT 74.545 132.665 74.815 133.570 ;
        RECT 75.000 133.425 75.665 133.595 ;
        RECT 74.985 132.495 75.315 133.255 ;
        RECT 75.495 132.665 75.665 133.425 ;
        RECT 76.845 133.585 78.535 134.105 ;
        RECT 78.705 133.755 80.355 134.275 ;
        RECT 80.565 134.225 80.795 135.045 ;
        RECT 80.965 134.245 81.295 134.875 ;
        RECT 80.545 133.805 80.875 134.055 ;
        RECT 81.045 133.645 81.295 134.245 ;
        RECT 81.465 134.225 81.675 135.045 ;
        RECT 81.945 134.225 82.175 135.045 ;
        RECT 82.345 134.245 82.675 134.875 ;
        RECT 81.925 133.805 82.255 134.055 ;
        RECT 82.425 133.645 82.675 134.245 ;
        RECT 82.845 134.225 83.055 135.045 ;
        RECT 83.560 134.235 83.805 134.840 ;
        RECT 84.025 134.510 84.535 135.045 ;
        RECT 76.845 132.495 80.355 133.585 ;
        RECT 80.565 132.495 80.795 133.635 ;
        RECT 80.965 132.665 81.295 133.645 ;
        RECT 81.465 132.495 81.675 133.635 ;
        RECT 81.945 132.495 82.175 133.635 ;
        RECT 82.345 132.665 82.675 133.645 ;
        RECT 83.285 134.065 84.515 134.235 ;
        RECT 82.845 132.495 83.055 133.635 ;
        RECT 83.285 133.255 83.625 134.065 ;
        RECT 83.795 133.500 84.545 133.690 ;
        RECT 83.285 132.845 83.800 133.255 ;
        RECT 84.035 132.495 84.205 133.255 ;
        RECT 84.375 132.835 84.545 133.500 ;
        RECT 84.715 133.515 84.905 134.875 ;
        RECT 85.075 134.705 85.350 134.875 ;
        RECT 85.075 134.535 85.355 134.705 ;
        RECT 85.075 133.715 85.350 134.535 ;
        RECT 85.540 134.510 86.070 134.875 ;
        RECT 86.495 134.645 86.825 135.045 ;
        RECT 85.895 134.475 86.070 134.510 ;
        RECT 85.555 133.515 85.725 134.315 ;
        RECT 84.715 133.345 85.725 133.515 ;
        RECT 85.895 134.305 86.825 134.475 ;
        RECT 86.995 134.305 87.250 134.875 ;
        RECT 85.895 133.175 86.065 134.305 ;
        RECT 86.655 134.135 86.825 134.305 ;
        RECT 84.940 133.005 86.065 133.175 ;
        RECT 86.235 133.805 86.430 134.135 ;
        RECT 86.655 133.805 86.910 134.135 ;
        RECT 86.235 132.835 86.405 133.805 ;
        RECT 87.080 133.635 87.250 134.305 ;
        RECT 87.465 134.225 87.695 135.045 ;
        RECT 87.865 134.245 88.195 134.875 ;
        RECT 87.445 133.805 87.775 134.055 ;
        RECT 87.945 133.645 88.195 134.245 ;
        RECT 88.365 134.225 88.575 135.045 ;
        RECT 88.805 134.320 89.095 135.045 ;
        RECT 89.540 134.235 89.785 134.840 ;
        RECT 90.005 134.510 90.515 135.045 ;
        RECT 89.265 134.065 90.495 134.235 ;
        RECT 84.375 132.665 86.405 132.835 ;
        RECT 86.575 132.495 86.745 133.635 ;
        RECT 86.915 132.665 87.250 133.635 ;
        RECT 87.465 132.495 87.695 133.635 ;
        RECT 87.865 132.665 88.195 133.645 ;
        RECT 88.365 132.495 88.575 133.635 ;
        RECT 88.805 132.495 89.095 133.660 ;
        RECT 89.265 133.255 89.605 134.065 ;
        RECT 89.775 133.500 90.525 133.690 ;
        RECT 89.265 132.845 89.780 133.255 ;
        RECT 90.015 132.495 90.185 133.255 ;
        RECT 90.355 132.835 90.525 133.500 ;
        RECT 90.695 133.515 90.885 134.875 ;
        RECT 91.055 134.025 91.330 134.875 ;
        RECT 91.520 134.510 92.050 134.875 ;
        RECT 92.475 134.645 92.805 135.045 ;
        RECT 91.875 134.475 92.050 134.510 ;
        RECT 91.055 133.855 91.335 134.025 ;
        RECT 91.055 133.715 91.330 133.855 ;
        RECT 91.535 133.515 91.705 134.315 ;
        RECT 90.695 133.345 91.705 133.515 ;
        RECT 91.875 134.305 92.805 134.475 ;
        RECT 92.975 134.305 93.230 134.875 ;
        RECT 93.465 134.565 93.745 135.045 ;
        RECT 93.915 134.395 94.175 134.785 ;
        RECT 94.350 134.565 94.605 135.045 ;
        RECT 94.775 134.395 95.070 134.785 ;
        RECT 95.250 134.565 95.525 135.045 ;
        RECT 95.695 134.545 95.995 134.875 ;
        RECT 96.540 134.705 96.795 134.865 ;
        RECT 91.875 133.175 92.045 134.305 ;
        RECT 92.635 134.135 92.805 134.305 ;
        RECT 90.920 133.005 92.045 133.175 ;
        RECT 92.215 133.805 92.410 134.135 ;
        RECT 92.635 133.805 92.890 134.135 ;
        RECT 92.215 132.835 92.385 133.805 ;
        RECT 93.060 133.635 93.230 134.305 ;
        RECT 90.355 132.665 92.385 132.835 ;
        RECT 92.555 132.495 92.725 133.635 ;
        RECT 92.895 132.665 93.230 133.635 ;
        RECT 93.420 134.225 95.070 134.395 ;
        RECT 93.420 133.715 93.825 134.225 ;
        RECT 93.995 133.885 95.135 134.055 ;
        RECT 93.420 133.545 94.175 133.715 ;
        RECT 93.460 132.495 93.745 133.365 ;
        RECT 93.915 133.295 94.175 133.545 ;
        RECT 94.965 133.635 95.135 133.885 ;
        RECT 95.305 133.805 95.655 134.375 ;
        RECT 95.825 133.635 95.995 134.545 ;
        RECT 96.455 134.535 96.795 134.705 ;
        RECT 96.975 134.585 97.260 135.045 ;
        RECT 94.965 133.465 95.995 133.635 ;
        RECT 93.915 133.125 95.035 133.295 ;
        RECT 93.915 132.665 94.175 133.125 ;
        RECT 94.350 132.495 94.605 132.955 ;
        RECT 94.775 132.665 95.035 133.125 ;
        RECT 95.205 132.495 95.515 133.295 ;
        RECT 95.685 132.665 95.995 133.465 ;
        RECT 96.540 134.335 96.795 134.535 ;
        RECT 96.540 133.475 96.720 134.335 ;
        RECT 97.440 134.135 97.690 134.785 ;
        RECT 96.890 133.805 97.690 134.135 ;
        RECT 96.540 132.805 96.795 133.475 ;
        RECT 96.975 132.495 97.260 133.295 ;
        RECT 97.440 133.215 97.690 133.805 ;
        RECT 97.890 134.450 98.210 134.780 ;
        RECT 98.390 134.565 99.050 135.045 ;
        RECT 99.250 134.655 100.100 134.825 ;
        RECT 97.890 133.555 98.080 134.450 ;
        RECT 98.400 134.125 99.060 134.395 ;
        RECT 98.730 134.065 99.060 134.125 ;
        RECT 98.250 133.895 98.580 133.955 ;
        RECT 99.250 133.895 99.420 134.655 ;
        RECT 100.660 134.585 100.980 135.045 ;
        RECT 101.180 134.405 101.430 134.835 ;
        RECT 101.720 134.605 102.130 135.045 ;
        RECT 102.300 134.665 103.315 134.865 ;
        RECT 99.590 134.235 100.840 134.405 ;
        RECT 99.590 134.115 99.920 134.235 ;
        RECT 98.250 133.725 100.150 133.895 ;
        RECT 97.890 133.385 99.810 133.555 ;
        RECT 97.890 133.365 98.210 133.385 ;
        RECT 97.440 132.705 97.770 133.215 ;
        RECT 98.040 132.755 98.210 133.365 ;
        RECT 99.980 133.215 100.150 133.725 ;
        RECT 100.320 133.655 100.500 134.065 ;
        RECT 100.670 133.475 100.840 134.235 ;
        RECT 98.380 132.495 98.710 133.185 ;
        RECT 98.940 133.045 100.150 133.215 ;
        RECT 100.320 133.165 100.840 133.475 ;
        RECT 101.010 134.065 101.430 134.405 ;
        RECT 101.720 134.065 102.130 134.395 ;
        RECT 101.010 133.295 101.200 134.065 ;
        RECT 102.300 133.935 102.470 134.665 ;
        RECT 103.615 134.495 103.785 134.825 ;
        RECT 103.955 134.665 104.285 135.045 ;
        RECT 102.640 134.115 102.990 134.485 ;
        RECT 102.300 133.895 102.720 133.935 ;
        RECT 101.370 133.725 102.720 133.895 ;
        RECT 101.370 133.565 101.620 133.725 ;
        RECT 102.130 133.295 102.380 133.555 ;
        RECT 101.010 133.045 102.380 133.295 ;
        RECT 98.940 132.755 99.180 133.045 ;
        RECT 99.980 132.965 100.150 133.045 ;
        RECT 99.380 132.495 99.800 132.875 ;
        RECT 99.980 132.715 100.610 132.965 ;
        RECT 101.080 132.495 101.410 132.875 ;
        RECT 101.580 132.755 101.750 133.045 ;
        RECT 102.550 132.880 102.720 133.725 ;
        RECT 103.170 133.555 103.390 134.425 ;
        RECT 103.615 134.305 104.310 134.495 ;
        RECT 102.890 133.175 103.390 133.555 ;
        RECT 103.560 133.505 103.970 134.125 ;
        RECT 104.140 133.335 104.310 134.305 ;
        RECT 103.615 133.165 104.310 133.335 ;
        RECT 101.930 132.495 102.310 132.875 ;
        RECT 102.550 132.710 103.380 132.880 ;
        RECT 103.615 132.665 103.785 133.165 ;
        RECT 103.955 132.495 104.285 132.995 ;
        RECT 104.500 132.665 104.725 134.785 ;
        RECT 104.895 134.665 105.225 135.045 ;
        RECT 105.395 134.495 105.565 134.785 ;
        RECT 104.900 134.325 105.565 134.495 ;
        RECT 104.900 133.335 105.130 134.325 ;
        RECT 105.830 134.305 106.085 134.875 ;
        RECT 106.255 134.645 106.585 135.045 ;
        RECT 107.010 134.510 107.540 134.875 ;
        RECT 107.730 134.705 108.005 134.875 ;
        RECT 107.725 134.535 108.005 134.705 ;
        RECT 107.010 134.475 107.185 134.510 ;
        RECT 106.255 134.305 107.185 134.475 ;
        RECT 105.300 133.505 105.650 134.155 ;
        RECT 105.830 133.635 106.000 134.305 ;
        RECT 106.255 134.135 106.425 134.305 ;
        RECT 106.170 133.805 106.425 134.135 ;
        RECT 106.650 133.805 106.845 134.135 ;
        RECT 104.900 133.165 105.565 133.335 ;
        RECT 104.895 132.495 105.225 132.995 ;
        RECT 105.395 132.665 105.565 133.165 ;
        RECT 105.830 132.665 106.165 133.635 ;
        RECT 106.335 132.495 106.505 133.635 ;
        RECT 106.675 132.835 106.845 133.805 ;
        RECT 107.015 133.175 107.185 134.305 ;
        RECT 107.355 133.515 107.525 134.315 ;
        RECT 107.730 133.715 108.005 134.535 ;
        RECT 108.175 133.515 108.365 134.875 ;
        RECT 108.545 134.510 109.055 135.045 ;
        RECT 109.275 134.235 109.520 134.840 ;
        RECT 110.885 134.275 114.395 135.045 ;
        RECT 114.565 134.320 114.855 135.045 ;
        RECT 108.565 134.065 109.795 134.235 ;
        RECT 107.355 133.345 108.365 133.515 ;
        RECT 108.535 133.500 109.285 133.690 ;
        RECT 107.015 133.005 108.140 133.175 ;
        RECT 108.535 132.835 108.705 133.500 ;
        RECT 109.455 133.255 109.795 134.065 ;
        RECT 106.675 132.665 108.705 132.835 ;
        RECT 108.875 132.495 109.045 133.255 ;
        RECT 109.280 132.845 109.795 133.255 ;
        RECT 110.885 133.585 112.575 134.105 ;
        RECT 112.745 133.755 114.395 134.275 ;
        RECT 115.300 134.235 115.545 134.840 ;
        RECT 115.765 134.510 116.275 135.045 ;
        RECT 115.025 134.065 116.255 134.235 ;
        RECT 110.885 132.495 114.395 133.585 ;
        RECT 114.565 132.495 114.855 133.660 ;
        RECT 115.025 133.255 115.365 134.065 ;
        RECT 115.535 133.500 116.285 133.690 ;
        RECT 115.025 132.845 115.540 133.255 ;
        RECT 115.775 132.495 115.945 133.255 ;
        RECT 116.115 132.835 116.285 133.500 ;
        RECT 116.455 133.515 116.645 134.875 ;
        RECT 116.815 134.705 117.090 134.875 ;
        RECT 116.815 134.535 117.095 134.705 ;
        RECT 116.815 133.715 117.090 134.535 ;
        RECT 117.280 134.510 117.810 134.875 ;
        RECT 118.235 134.645 118.565 135.045 ;
        RECT 117.635 134.475 117.810 134.510 ;
        RECT 117.295 133.515 117.465 134.315 ;
        RECT 116.455 133.345 117.465 133.515 ;
        RECT 117.635 134.305 118.565 134.475 ;
        RECT 118.735 134.305 118.990 134.875 ;
        RECT 117.635 133.175 117.805 134.305 ;
        RECT 118.395 134.135 118.565 134.305 ;
        RECT 116.680 133.005 117.805 133.175 ;
        RECT 117.975 133.805 118.170 134.135 ;
        RECT 118.395 133.805 118.650 134.135 ;
        RECT 117.975 132.835 118.145 133.805 ;
        RECT 118.820 133.635 118.990 134.305 ;
        RECT 119.205 134.225 119.435 135.045 ;
        RECT 119.605 134.245 119.935 134.875 ;
        RECT 119.185 133.805 119.515 134.055 ;
        RECT 119.685 133.645 119.935 134.245 ;
        RECT 120.105 134.225 120.315 135.045 ;
        RECT 121.095 134.495 121.265 134.875 ;
        RECT 121.445 134.665 121.775 135.045 ;
        RECT 121.095 134.325 121.760 134.495 ;
        RECT 121.955 134.370 122.215 134.875 ;
        RECT 121.025 133.775 121.355 134.145 ;
        RECT 121.590 134.070 121.760 134.325 ;
        RECT 116.115 132.665 118.145 132.835 ;
        RECT 118.315 132.495 118.485 133.635 ;
        RECT 118.655 132.665 118.990 133.635 ;
        RECT 119.205 132.495 119.435 133.635 ;
        RECT 119.605 132.665 119.935 133.645 ;
        RECT 121.590 133.740 121.875 134.070 ;
        RECT 120.105 132.495 120.315 133.635 ;
        RECT 121.590 133.595 121.760 133.740 ;
        RECT 121.095 133.425 121.760 133.595 ;
        RECT 122.045 133.570 122.215 134.370 ;
        RECT 122.475 134.495 122.645 134.875 ;
        RECT 122.825 134.665 123.155 135.045 ;
        RECT 122.475 134.325 123.140 134.495 ;
        RECT 123.335 134.370 123.595 134.875 ;
        RECT 122.405 133.775 122.735 134.145 ;
        RECT 122.970 134.070 123.140 134.325 ;
        RECT 122.970 133.740 123.255 134.070 ;
        RECT 122.970 133.595 123.140 133.740 ;
        RECT 121.095 132.665 121.265 133.425 ;
        RECT 121.445 132.495 121.775 133.255 ;
        RECT 121.945 132.665 122.215 133.570 ;
        RECT 122.475 133.425 123.140 133.595 ;
        RECT 123.425 133.570 123.595 134.370 ;
        RECT 123.765 134.275 126.355 135.045 ;
        RECT 126.525 134.295 127.735 135.045 ;
        RECT 122.475 132.665 122.645 133.425 ;
        RECT 122.825 132.495 123.155 133.255 ;
        RECT 123.325 132.665 123.595 133.570 ;
        RECT 123.765 133.585 124.975 134.105 ;
        RECT 125.145 133.755 126.355 134.275 ;
        RECT 126.525 133.585 127.045 134.125 ;
        RECT 127.215 133.755 127.735 134.295 ;
        RECT 123.765 132.495 126.355 133.585 ;
        RECT 126.525 132.495 127.735 133.585 ;
        RECT 29.840 132.325 127.820 132.495 ;
        RECT 29.925 131.235 31.135 132.325 ;
        RECT 29.925 130.525 30.445 131.065 ;
        RECT 30.615 130.695 31.135 131.235 ;
        RECT 32.285 131.185 32.495 132.325 ;
        RECT 32.665 131.175 32.995 132.155 ;
        RECT 33.165 131.185 33.395 132.325 ;
        RECT 33.695 131.395 33.865 132.155 ;
        RECT 34.045 131.565 34.375 132.325 ;
        RECT 33.695 131.225 34.360 131.395 ;
        RECT 34.545 131.250 34.815 132.155 ;
        RECT 29.925 129.775 31.135 130.525 ;
        RECT 32.285 129.775 32.495 130.595 ;
        RECT 32.665 130.575 32.915 131.175 ;
        RECT 34.190 131.080 34.360 131.225 ;
        RECT 33.085 130.765 33.415 131.015 ;
        RECT 33.625 130.675 33.955 131.045 ;
        RECT 34.190 130.750 34.475 131.080 ;
        RECT 32.665 129.945 32.995 130.575 ;
        RECT 33.165 129.775 33.395 130.595 ;
        RECT 34.190 130.495 34.360 130.750 ;
        RECT 33.695 130.325 34.360 130.495 ;
        RECT 34.645 130.450 34.815 131.250 ;
        RECT 34.985 131.565 35.500 131.975 ;
        RECT 35.735 131.565 35.905 132.325 ;
        RECT 36.075 131.985 38.105 132.155 ;
        RECT 34.985 130.755 35.325 131.565 ;
        RECT 36.075 131.320 36.245 131.985 ;
        RECT 36.640 131.645 37.765 131.815 ;
        RECT 35.495 131.130 36.245 131.320 ;
        RECT 36.415 131.305 37.425 131.475 ;
        RECT 34.985 130.585 36.215 130.755 ;
        RECT 33.695 129.945 33.865 130.325 ;
        RECT 34.045 129.775 34.375 130.155 ;
        RECT 34.555 129.945 34.815 130.450 ;
        RECT 35.260 129.980 35.505 130.585 ;
        RECT 35.725 129.775 36.235 130.310 ;
        RECT 36.415 129.945 36.605 131.305 ;
        RECT 36.775 130.285 37.050 131.105 ;
        RECT 37.255 130.505 37.425 131.305 ;
        RECT 37.595 130.515 37.765 131.645 ;
        RECT 37.935 131.015 38.105 131.985 ;
        RECT 38.275 131.185 38.445 132.325 ;
        RECT 38.615 131.185 38.950 132.155 ;
        RECT 39.215 131.655 39.385 132.155 ;
        RECT 39.555 131.825 39.885 132.325 ;
        RECT 39.215 131.485 39.880 131.655 ;
        RECT 37.935 130.685 38.130 131.015 ;
        RECT 38.355 130.685 38.610 131.015 ;
        RECT 38.355 130.515 38.525 130.685 ;
        RECT 38.780 130.515 38.950 131.185 ;
        RECT 39.130 130.665 39.480 131.315 ;
        RECT 37.595 130.345 38.525 130.515 ;
        RECT 37.595 130.310 37.770 130.345 ;
        RECT 36.775 130.115 37.055 130.285 ;
        RECT 36.775 129.945 37.050 130.115 ;
        RECT 37.240 129.945 37.770 130.310 ;
        RECT 38.195 129.775 38.525 130.175 ;
        RECT 38.695 129.945 38.950 130.515 ;
        RECT 39.650 130.495 39.880 131.485 ;
        RECT 39.215 130.325 39.880 130.495 ;
        RECT 39.215 130.035 39.385 130.325 ;
        RECT 39.555 129.775 39.885 130.155 ;
        RECT 40.055 130.035 40.280 132.155 ;
        RECT 40.495 131.825 40.825 132.325 ;
        RECT 40.995 131.655 41.165 132.155 ;
        RECT 41.400 131.940 42.230 132.110 ;
        RECT 42.470 131.945 42.850 132.325 ;
        RECT 40.470 131.485 41.165 131.655 ;
        RECT 40.470 130.515 40.640 131.485 ;
        RECT 40.810 130.695 41.220 131.315 ;
        RECT 41.390 131.265 41.890 131.645 ;
        RECT 40.470 130.325 41.165 130.515 ;
        RECT 41.390 130.395 41.610 131.265 ;
        RECT 42.060 131.095 42.230 131.940 ;
        RECT 43.030 131.775 43.200 132.065 ;
        RECT 43.370 131.945 43.700 132.325 ;
        RECT 44.170 131.855 44.800 132.105 ;
        RECT 44.980 131.945 45.400 132.325 ;
        RECT 44.630 131.775 44.800 131.855 ;
        RECT 45.600 131.775 45.840 132.065 ;
        RECT 42.400 131.525 43.770 131.775 ;
        RECT 42.400 131.265 42.650 131.525 ;
        RECT 43.160 131.095 43.410 131.255 ;
        RECT 42.060 130.925 43.410 131.095 ;
        RECT 42.060 130.885 42.480 130.925 ;
        RECT 41.790 130.335 42.140 130.705 ;
        RECT 40.495 129.775 40.825 130.155 ;
        RECT 40.995 129.995 41.165 130.325 ;
        RECT 42.310 130.155 42.480 130.885 ;
        RECT 43.580 130.755 43.770 131.525 ;
        RECT 42.650 130.425 43.060 130.755 ;
        RECT 43.350 130.415 43.770 130.755 ;
        RECT 43.940 131.345 44.460 131.655 ;
        RECT 44.630 131.605 45.840 131.775 ;
        RECT 46.070 131.635 46.400 132.325 ;
        RECT 43.940 130.585 44.110 131.345 ;
        RECT 44.280 130.755 44.460 131.165 ;
        RECT 44.630 131.095 44.800 131.605 ;
        RECT 46.570 131.455 46.740 132.065 ;
        RECT 47.010 131.605 47.340 132.115 ;
        RECT 46.570 131.435 46.890 131.455 ;
        RECT 44.970 131.265 46.890 131.435 ;
        RECT 44.630 130.925 46.530 131.095 ;
        RECT 44.860 130.585 45.190 130.705 ;
        RECT 43.940 130.415 45.190 130.585 ;
        RECT 41.465 129.955 42.480 130.155 ;
        RECT 42.650 129.775 43.060 130.215 ;
        RECT 43.350 129.985 43.600 130.415 ;
        RECT 43.800 129.775 44.120 130.235 ;
        RECT 45.360 130.165 45.530 130.925 ;
        RECT 46.200 130.865 46.530 130.925 ;
        RECT 45.720 130.695 46.050 130.755 ;
        RECT 45.720 130.425 46.380 130.695 ;
        RECT 46.700 130.370 46.890 131.265 ;
        RECT 44.680 129.995 45.530 130.165 ;
        RECT 45.730 129.775 46.390 130.255 ;
        RECT 46.570 130.040 46.890 130.370 ;
        RECT 47.090 131.015 47.340 131.605 ;
        RECT 47.520 131.525 47.805 132.325 ;
        RECT 47.985 131.985 48.240 132.015 ;
        RECT 47.985 131.815 48.325 131.985 ;
        RECT 47.985 131.345 48.240 131.815 ;
        RECT 47.090 130.685 47.890 131.015 ;
        RECT 47.090 130.035 47.340 130.685 ;
        RECT 48.060 130.485 48.240 131.345 ;
        RECT 48.875 131.395 49.045 132.155 ;
        RECT 49.225 131.565 49.555 132.325 ;
        RECT 48.875 131.225 49.540 131.395 ;
        RECT 49.725 131.250 49.995 132.155 ;
        RECT 49.370 131.080 49.540 131.225 ;
        RECT 48.805 130.675 49.135 131.045 ;
        RECT 49.370 130.750 49.655 131.080 ;
        RECT 49.370 130.495 49.540 130.750 ;
        RECT 47.520 129.775 47.805 130.235 ;
        RECT 47.985 129.955 48.240 130.485 ;
        RECT 48.875 130.325 49.540 130.495 ;
        RECT 49.825 130.450 49.995 131.250 ;
        RECT 50.165 131.160 50.455 132.325 ;
        RECT 50.630 131.185 50.965 132.155 ;
        RECT 51.135 131.185 51.305 132.325 ;
        RECT 51.475 131.985 53.505 132.155 ;
        RECT 50.630 130.515 50.800 131.185 ;
        RECT 51.475 131.015 51.645 131.985 ;
        RECT 50.970 130.685 51.225 131.015 ;
        RECT 51.450 130.685 51.645 131.015 ;
        RECT 51.815 131.645 52.940 131.815 ;
        RECT 51.055 130.515 51.225 130.685 ;
        RECT 51.815 130.515 51.985 131.645 ;
        RECT 48.875 129.945 49.045 130.325 ;
        RECT 49.225 129.775 49.555 130.155 ;
        RECT 49.735 129.945 49.995 130.450 ;
        RECT 50.165 129.775 50.455 130.500 ;
        RECT 50.630 129.945 50.885 130.515 ;
        RECT 51.055 130.345 51.985 130.515 ;
        RECT 52.155 131.305 53.165 131.475 ;
        RECT 52.155 130.505 52.325 131.305 ;
        RECT 52.530 130.625 52.805 131.105 ;
        RECT 52.525 130.455 52.805 130.625 ;
        RECT 51.810 130.310 51.985 130.345 ;
        RECT 51.055 129.775 51.385 130.175 ;
        RECT 51.810 129.945 52.340 130.310 ;
        RECT 52.530 129.945 52.805 130.455 ;
        RECT 52.975 129.945 53.165 131.305 ;
        RECT 53.335 131.320 53.505 131.985 ;
        RECT 53.675 131.565 53.845 132.325 ;
        RECT 54.080 131.565 54.595 131.975 ;
        RECT 55.885 131.655 56.165 132.325 ;
        RECT 53.335 131.130 54.085 131.320 ;
        RECT 54.255 130.755 54.595 131.565 ;
        RECT 56.335 131.435 56.635 131.985 ;
        RECT 56.835 131.605 57.165 132.325 ;
        RECT 57.355 131.605 57.815 132.155 ;
        RECT 55.700 131.015 55.965 131.375 ;
        RECT 56.335 131.265 57.275 131.435 ;
        RECT 57.105 131.015 57.275 131.265 ;
        RECT 55.700 130.765 56.375 131.015 ;
        RECT 56.595 130.765 56.935 131.015 ;
        RECT 53.365 130.585 54.595 130.755 ;
        RECT 57.105 130.685 57.395 131.015 ;
        RECT 57.105 130.595 57.275 130.685 ;
        RECT 53.345 129.775 53.855 130.310 ;
        RECT 54.075 129.980 54.320 130.585 ;
        RECT 55.885 130.405 57.275 130.595 ;
        RECT 55.885 130.045 56.215 130.405 ;
        RECT 57.565 130.235 57.815 131.605 ;
        RECT 57.985 131.565 58.500 131.975 ;
        RECT 58.735 131.565 58.905 132.325 ;
        RECT 59.075 131.985 61.105 132.155 ;
        RECT 57.985 130.755 58.325 131.565 ;
        RECT 59.075 131.320 59.245 131.985 ;
        RECT 59.640 131.645 60.765 131.815 ;
        RECT 58.495 131.130 59.245 131.320 ;
        RECT 59.415 131.305 60.425 131.475 ;
        RECT 57.985 130.585 59.215 130.755 ;
        RECT 56.835 129.775 57.085 130.235 ;
        RECT 57.255 129.945 57.815 130.235 ;
        RECT 58.260 129.980 58.505 130.585 ;
        RECT 58.725 129.775 59.235 130.310 ;
        RECT 59.415 129.945 59.605 131.305 ;
        RECT 59.775 130.285 60.050 131.105 ;
        RECT 60.255 130.505 60.425 131.305 ;
        RECT 60.595 130.515 60.765 131.645 ;
        RECT 60.935 131.015 61.105 131.985 ;
        RECT 61.275 131.185 61.445 132.325 ;
        RECT 61.615 131.185 61.950 132.155 ;
        RECT 60.935 130.685 61.130 131.015 ;
        RECT 61.355 130.685 61.610 131.015 ;
        RECT 61.355 130.515 61.525 130.685 ;
        RECT 61.780 130.515 61.950 131.185 ;
        RECT 62.125 131.565 62.640 131.975 ;
        RECT 62.875 131.565 63.045 132.325 ;
        RECT 63.215 131.985 65.245 132.155 ;
        RECT 62.125 130.755 62.465 131.565 ;
        RECT 63.215 131.320 63.385 131.985 ;
        RECT 63.780 131.645 64.905 131.815 ;
        RECT 62.635 131.130 63.385 131.320 ;
        RECT 63.555 131.305 64.565 131.475 ;
        RECT 62.125 130.585 63.355 130.755 ;
        RECT 60.595 130.345 61.525 130.515 ;
        RECT 60.595 130.310 60.770 130.345 ;
        RECT 59.775 130.115 60.055 130.285 ;
        RECT 59.775 129.945 60.050 130.115 ;
        RECT 60.240 129.945 60.770 130.310 ;
        RECT 61.195 129.775 61.525 130.175 ;
        RECT 61.695 129.945 61.950 130.515 ;
        RECT 62.400 129.980 62.645 130.585 ;
        RECT 62.865 129.775 63.375 130.310 ;
        RECT 63.555 129.945 63.745 131.305 ;
        RECT 63.915 130.625 64.190 131.105 ;
        RECT 63.915 130.455 64.195 130.625 ;
        RECT 64.395 130.505 64.565 131.305 ;
        RECT 64.735 130.515 64.905 131.645 ;
        RECT 65.075 131.015 65.245 131.985 ;
        RECT 65.415 131.185 65.585 132.325 ;
        RECT 65.755 131.185 66.090 132.155 ;
        RECT 66.640 131.985 66.895 132.015 ;
        RECT 66.555 131.815 66.895 131.985 ;
        RECT 65.075 130.685 65.270 131.015 ;
        RECT 65.495 130.685 65.750 131.015 ;
        RECT 65.495 130.515 65.665 130.685 ;
        RECT 65.920 130.515 66.090 131.185 ;
        RECT 63.915 129.945 64.190 130.455 ;
        RECT 64.735 130.345 65.665 130.515 ;
        RECT 64.735 130.310 64.910 130.345 ;
        RECT 64.380 129.945 64.910 130.310 ;
        RECT 65.335 129.775 65.665 130.175 ;
        RECT 65.835 129.945 66.090 130.515 ;
        RECT 66.640 131.345 66.895 131.815 ;
        RECT 67.075 131.525 67.360 132.325 ;
        RECT 67.540 131.605 67.870 132.115 ;
        RECT 66.640 130.485 66.820 131.345 ;
        RECT 67.540 131.015 67.790 131.605 ;
        RECT 68.140 131.455 68.310 132.065 ;
        RECT 68.480 131.635 68.810 132.325 ;
        RECT 69.040 131.775 69.280 132.065 ;
        RECT 69.480 131.945 69.900 132.325 ;
        RECT 70.080 131.855 70.710 132.105 ;
        RECT 71.180 131.945 71.510 132.325 ;
        RECT 70.080 131.775 70.250 131.855 ;
        RECT 71.680 131.775 71.850 132.065 ;
        RECT 72.030 131.945 72.410 132.325 ;
        RECT 72.650 131.940 73.480 132.110 ;
        RECT 69.040 131.605 70.250 131.775 ;
        RECT 66.990 130.685 67.790 131.015 ;
        RECT 66.640 129.955 66.895 130.485 ;
        RECT 67.075 129.775 67.360 130.235 ;
        RECT 67.540 130.035 67.790 130.685 ;
        RECT 67.990 131.435 68.310 131.455 ;
        RECT 67.990 131.265 69.910 131.435 ;
        RECT 67.990 130.370 68.180 131.265 ;
        RECT 70.080 131.095 70.250 131.605 ;
        RECT 70.420 131.345 70.940 131.655 ;
        RECT 68.350 130.925 70.250 131.095 ;
        RECT 68.350 130.865 68.680 130.925 ;
        RECT 68.830 130.695 69.160 130.755 ;
        RECT 68.500 130.425 69.160 130.695 ;
        RECT 67.990 130.040 68.310 130.370 ;
        RECT 68.490 129.775 69.150 130.255 ;
        RECT 69.350 130.165 69.520 130.925 ;
        RECT 70.420 130.755 70.600 131.165 ;
        RECT 69.690 130.585 70.020 130.705 ;
        RECT 70.770 130.585 70.940 131.345 ;
        RECT 69.690 130.415 70.940 130.585 ;
        RECT 71.110 131.525 72.480 131.775 ;
        RECT 71.110 130.755 71.300 131.525 ;
        RECT 72.230 131.265 72.480 131.525 ;
        RECT 71.470 131.095 71.720 131.255 ;
        RECT 72.650 131.095 72.820 131.940 ;
        RECT 73.715 131.655 73.885 132.155 ;
        RECT 74.055 131.825 74.385 132.325 ;
        RECT 72.990 131.265 73.490 131.645 ;
        RECT 73.715 131.485 74.410 131.655 ;
        RECT 71.470 130.925 72.820 131.095 ;
        RECT 72.400 130.885 72.820 130.925 ;
        RECT 71.110 130.415 71.530 130.755 ;
        RECT 71.820 130.425 72.230 130.755 ;
        RECT 69.350 129.995 70.200 130.165 ;
        RECT 70.760 129.775 71.080 130.235 ;
        RECT 71.280 129.985 71.530 130.415 ;
        RECT 71.820 129.775 72.230 130.215 ;
        RECT 72.400 130.155 72.570 130.885 ;
        RECT 72.740 130.335 73.090 130.705 ;
        RECT 73.270 130.395 73.490 131.265 ;
        RECT 73.660 130.695 74.070 131.315 ;
        RECT 74.240 130.515 74.410 131.485 ;
        RECT 73.715 130.325 74.410 130.515 ;
        RECT 72.400 129.955 73.415 130.155 ;
        RECT 73.715 129.995 73.885 130.325 ;
        RECT 74.055 129.775 74.385 130.155 ;
        RECT 74.600 130.035 74.825 132.155 ;
        RECT 74.995 131.825 75.325 132.325 ;
        RECT 75.495 131.655 75.665 132.155 ;
        RECT 75.000 131.485 75.665 131.655 ;
        RECT 75.000 130.495 75.230 131.485 ;
        RECT 75.400 130.665 75.750 131.315 ;
        RECT 75.925 131.160 76.215 132.325 ;
        RECT 76.385 131.565 76.900 131.975 ;
        RECT 77.135 131.565 77.305 132.325 ;
        RECT 77.475 131.985 79.505 132.155 ;
        RECT 76.385 130.755 76.725 131.565 ;
        RECT 77.475 131.320 77.645 131.985 ;
        RECT 78.040 131.645 79.165 131.815 ;
        RECT 76.895 131.130 77.645 131.320 ;
        RECT 77.815 131.305 78.825 131.475 ;
        RECT 76.385 130.585 77.615 130.755 ;
        RECT 75.000 130.325 75.665 130.495 ;
        RECT 74.995 129.775 75.325 130.155 ;
        RECT 75.495 130.035 75.665 130.325 ;
        RECT 75.925 129.775 76.215 130.500 ;
        RECT 76.660 129.980 76.905 130.585 ;
        RECT 77.125 129.775 77.635 130.310 ;
        RECT 77.815 129.945 78.005 131.305 ;
        RECT 78.175 130.965 78.450 131.105 ;
        RECT 78.175 130.795 78.455 130.965 ;
        RECT 78.175 129.945 78.450 130.795 ;
        RECT 78.655 130.505 78.825 131.305 ;
        RECT 78.995 130.515 79.165 131.645 ;
        RECT 79.335 131.015 79.505 131.985 ;
        RECT 79.675 131.185 79.845 132.325 ;
        RECT 80.015 131.185 80.350 132.155 ;
        RECT 80.900 131.345 81.155 132.015 ;
        RECT 81.335 131.525 81.620 132.325 ;
        RECT 81.800 131.605 82.130 132.115 ;
        RECT 80.900 131.305 81.080 131.345 ;
        RECT 79.335 130.685 79.530 131.015 ;
        RECT 79.755 130.685 80.010 131.015 ;
        RECT 79.755 130.515 79.925 130.685 ;
        RECT 80.180 130.515 80.350 131.185 ;
        RECT 80.815 131.135 81.080 131.305 ;
        RECT 78.995 130.345 79.925 130.515 ;
        RECT 78.995 130.310 79.170 130.345 ;
        RECT 78.640 129.945 79.170 130.310 ;
        RECT 79.595 129.775 79.925 130.175 ;
        RECT 80.095 129.945 80.350 130.515 ;
        RECT 80.900 130.485 81.080 131.135 ;
        RECT 81.800 131.015 82.050 131.605 ;
        RECT 82.400 131.455 82.570 132.065 ;
        RECT 82.740 131.635 83.070 132.325 ;
        RECT 83.300 131.775 83.540 132.065 ;
        RECT 83.740 131.945 84.160 132.325 ;
        RECT 84.340 131.855 84.970 132.105 ;
        RECT 85.440 131.945 85.770 132.325 ;
        RECT 84.340 131.775 84.510 131.855 ;
        RECT 85.940 131.775 86.110 132.065 ;
        RECT 86.290 131.945 86.670 132.325 ;
        RECT 86.910 131.940 87.740 132.110 ;
        RECT 83.300 131.605 84.510 131.775 ;
        RECT 81.250 130.685 82.050 131.015 ;
        RECT 80.900 129.955 81.155 130.485 ;
        RECT 81.335 129.775 81.620 130.235 ;
        RECT 81.800 130.035 82.050 130.685 ;
        RECT 82.250 131.435 82.570 131.455 ;
        RECT 82.250 131.265 84.170 131.435 ;
        RECT 82.250 130.370 82.440 131.265 ;
        RECT 84.340 131.095 84.510 131.605 ;
        RECT 84.680 131.345 85.200 131.655 ;
        RECT 82.610 130.925 84.510 131.095 ;
        RECT 82.610 130.865 82.940 130.925 ;
        RECT 83.090 130.695 83.420 130.755 ;
        RECT 82.760 130.425 83.420 130.695 ;
        RECT 82.250 130.040 82.570 130.370 ;
        RECT 82.750 129.775 83.410 130.255 ;
        RECT 83.610 130.165 83.780 130.925 ;
        RECT 84.680 130.755 84.860 131.165 ;
        RECT 83.950 130.585 84.280 130.705 ;
        RECT 85.030 130.585 85.200 131.345 ;
        RECT 83.950 130.415 85.200 130.585 ;
        RECT 85.370 131.525 86.740 131.775 ;
        RECT 85.370 130.755 85.560 131.525 ;
        RECT 86.490 131.265 86.740 131.525 ;
        RECT 85.730 131.095 85.980 131.255 ;
        RECT 86.910 131.095 87.080 131.940 ;
        RECT 87.975 131.655 88.145 132.155 ;
        RECT 88.315 131.825 88.645 132.325 ;
        RECT 87.250 131.265 87.750 131.645 ;
        RECT 87.975 131.485 88.670 131.655 ;
        RECT 85.730 130.925 87.080 131.095 ;
        RECT 86.660 130.885 87.080 130.925 ;
        RECT 85.370 130.415 85.790 130.755 ;
        RECT 86.080 130.425 86.490 130.755 ;
        RECT 83.610 129.995 84.460 130.165 ;
        RECT 85.020 129.775 85.340 130.235 ;
        RECT 85.540 129.985 85.790 130.415 ;
        RECT 86.080 129.775 86.490 130.215 ;
        RECT 86.660 130.155 86.830 130.885 ;
        RECT 87.000 130.335 87.350 130.705 ;
        RECT 87.530 130.395 87.750 131.265 ;
        RECT 87.920 130.695 88.330 131.315 ;
        RECT 88.500 130.515 88.670 131.485 ;
        RECT 87.975 130.325 88.670 130.515 ;
        RECT 86.660 129.955 87.675 130.155 ;
        RECT 87.975 129.995 88.145 130.325 ;
        RECT 88.315 129.775 88.645 130.155 ;
        RECT 88.860 130.035 89.085 132.155 ;
        RECT 89.255 131.825 89.585 132.325 ;
        RECT 89.755 131.655 89.925 132.155 ;
        RECT 89.260 131.485 89.925 131.655 ;
        RECT 89.260 130.495 89.490 131.485 ;
        RECT 89.660 130.665 90.010 131.315 ;
        RECT 90.185 131.250 90.455 132.155 ;
        RECT 90.625 131.565 90.955 132.325 ;
        RECT 91.135 131.395 91.305 132.155 ;
        RECT 92.400 131.985 92.655 132.015 ;
        RECT 92.315 131.815 92.655 131.985 ;
        RECT 89.260 130.325 89.925 130.495 ;
        RECT 89.255 129.775 89.585 130.155 ;
        RECT 89.755 130.035 89.925 130.325 ;
        RECT 90.185 130.450 90.355 131.250 ;
        RECT 90.640 131.225 91.305 131.395 ;
        RECT 92.400 131.345 92.655 131.815 ;
        RECT 92.835 131.525 93.120 132.325 ;
        RECT 93.300 131.605 93.630 132.115 ;
        RECT 90.640 131.080 90.810 131.225 ;
        RECT 90.525 130.750 90.810 131.080 ;
        RECT 90.640 130.495 90.810 130.750 ;
        RECT 91.045 130.675 91.375 131.045 ;
        RECT 90.185 129.945 90.445 130.450 ;
        RECT 90.640 130.325 91.305 130.495 ;
        RECT 90.625 129.775 90.955 130.155 ;
        RECT 91.135 129.945 91.305 130.325 ;
        RECT 92.400 130.485 92.580 131.345 ;
        RECT 93.300 131.015 93.550 131.605 ;
        RECT 93.900 131.455 94.070 132.065 ;
        RECT 94.240 131.635 94.570 132.325 ;
        RECT 94.800 131.775 95.040 132.065 ;
        RECT 95.240 131.945 95.660 132.325 ;
        RECT 95.840 131.855 96.470 132.105 ;
        RECT 96.940 131.945 97.270 132.325 ;
        RECT 95.840 131.775 96.010 131.855 ;
        RECT 97.440 131.775 97.610 132.065 ;
        RECT 97.790 131.945 98.170 132.325 ;
        RECT 98.410 131.940 99.240 132.110 ;
        RECT 94.800 131.605 96.010 131.775 ;
        RECT 92.750 130.685 93.550 131.015 ;
        RECT 92.400 129.955 92.655 130.485 ;
        RECT 92.835 129.775 93.120 130.235 ;
        RECT 93.300 130.035 93.550 130.685 ;
        RECT 93.750 131.435 94.070 131.455 ;
        RECT 93.750 131.265 95.670 131.435 ;
        RECT 93.750 130.370 93.940 131.265 ;
        RECT 95.840 131.095 96.010 131.605 ;
        RECT 96.180 131.345 96.700 131.655 ;
        RECT 94.110 130.925 96.010 131.095 ;
        RECT 94.110 130.865 94.440 130.925 ;
        RECT 94.590 130.695 94.920 130.755 ;
        RECT 94.260 130.425 94.920 130.695 ;
        RECT 93.750 130.040 94.070 130.370 ;
        RECT 94.250 129.775 94.910 130.255 ;
        RECT 95.110 130.165 95.280 130.925 ;
        RECT 96.180 130.755 96.360 131.165 ;
        RECT 95.450 130.585 95.780 130.705 ;
        RECT 96.530 130.585 96.700 131.345 ;
        RECT 95.450 130.415 96.700 130.585 ;
        RECT 96.870 131.525 98.240 131.775 ;
        RECT 96.870 130.755 97.060 131.525 ;
        RECT 97.990 131.265 98.240 131.525 ;
        RECT 97.230 131.095 97.480 131.255 ;
        RECT 98.410 131.095 98.580 131.940 ;
        RECT 99.475 131.655 99.645 132.155 ;
        RECT 99.815 131.825 100.145 132.325 ;
        RECT 98.750 131.265 99.250 131.645 ;
        RECT 99.475 131.485 100.170 131.655 ;
        RECT 97.230 130.925 98.580 131.095 ;
        RECT 98.160 130.885 98.580 130.925 ;
        RECT 96.870 130.415 97.290 130.755 ;
        RECT 97.580 130.425 97.990 130.755 ;
        RECT 95.110 129.995 95.960 130.165 ;
        RECT 96.520 129.775 96.840 130.235 ;
        RECT 97.040 129.985 97.290 130.415 ;
        RECT 97.580 129.775 97.990 130.215 ;
        RECT 98.160 130.155 98.330 130.885 ;
        RECT 98.500 130.335 98.850 130.705 ;
        RECT 99.030 130.395 99.250 131.265 ;
        RECT 99.420 130.695 99.830 131.315 ;
        RECT 100.000 130.515 100.170 131.485 ;
        RECT 99.475 130.325 100.170 130.515 ;
        RECT 98.160 129.955 99.175 130.155 ;
        RECT 99.475 129.995 99.645 130.325 ;
        RECT 99.815 129.775 100.145 130.155 ;
        RECT 100.360 130.035 100.585 132.155 ;
        RECT 100.755 131.825 101.085 132.325 ;
        RECT 101.255 131.655 101.425 132.155 ;
        RECT 100.760 131.485 101.425 131.655 ;
        RECT 100.760 130.495 100.990 131.485 ;
        RECT 101.160 130.665 101.510 131.315 ;
        RECT 101.685 131.160 101.975 132.325 ;
        RECT 102.185 131.185 102.415 132.325 ;
        RECT 102.585 131.175 102.915 132.155 ;
        RECT 103.085 131.185 103.295 132.325 ;
        RECT 103.525 131.250 103.795 132.155 ;
        RECT 103.965 131.565 104.295 132.325 ;
        RECT 104.475 131.395 104.645 132.155 ;
        RECT 102.165 130.765 102.495 131.015 ;
        RECT 100.760 130.325 101.425 130.495 ;
        RECT 100.755 129.775 101.085 130.155 ;
        RECT 101.255 130.035 101.425 130.325 ;
        RECT 101.685 129.775 101.975 130.500 ;
        RECT 102.185 129.775 102.415 130.595 ;
        RECT 102.665 130.575 102.915 131.175 ;
        RECT 102.585 129.945 102.915 130.575 ;
        RECT 103.085 129.775 103.295 130.595 ;
        RECT 103.525 130.450 103.695 131.250 ;
        RECT 103.980 131.225 104.645 131.395 ;
        RECT 104.905 131.235 106.115 132.325 ;
        RECT 106.285 131.565 106.800 131.975 ;
        RECT 107.035 131.565 107.205 132.325 ;
        RECT 107.375 131.985 109.405 132.155 ;
        RECT 103.980 131.080 104.150 131.225 ;
        RECT 103.865 130.750 104.150 131.080 ;
        RECT 103.980 130.495 104.150 130.750 ;
        RECT 104.385 130.675 104.715 131.045 ;
        RECT 104.905 130.695 105.425 131.235 ;
        RECT 105.595 130.525 106.115 131.065 ;
        RECT 106.285 130.755 106.625 131.565 ;
        RECT 107.375 131.320 107.545 131.985 ;
        RECT 107.940 131.645 109.065 131.815 ;
        RECT 106.795 131.130 107.545 131.320 ;
        RECT 107.715 131.305 108.725 131.475 ;
        RECT 106.285 130.585 107.515 130.755 ;
        RECT 103.525 129.945 103.785 130.450 ;
        RECT 103.980 130.325 104.645 130.495 ;
        RECT 103.965 129.775 104.295 130.155 ;
        RECT 104.475 129.945 104.645 130.325 ;
        RECT 104.905 129.775 106.115 130.525 ;
        RECT 106.560 129.980 106.805 130.585 ;
        RECT 107.025 129.775 107.535 130.310 ;
        RECT 107.715 129.945 107.905 131.305 ;
        RECT 108.075 130.965 108.350 131.105 ;
        RECT 108.075 130.795 108.355 130.965 ;
        RECT 108.075 129.945 108.350 130.795 ;
        RECT 108.555 130.505 108.725 131.305 ;
        RECT 108.895 130.515 109.065 131.645 ;
        RECT 109.235 131.015 109.405 131.985 ;
        RECT 109.575 131.185 109.745 132.325 ;
        RECT 109.915 131.185 110.250 132.155 ;
        RECT 110.515 131.395 110.685 132.155 ;
        RECT 110.865 131.565 111.195 132.325 ;
        RECT 110.515 131.225 111.180 131.395 ;
        RECT 111.365 131.250 111.635 132.155 ;
        RECT 109.235 130.685 109.430 131.015 ;
        RECT 109.655 130.685 109.910 131.015 ;
        RECT 109.655 130.515 109.825 130.685 ;
        RECT 110.080 130.515 110.250 131.185 ;
        RECT 111.010 131.080 111.180 131.225 ;
        RECT 110.445 130.675 110.775 131.045 ;
        RECT 111.010 130.750 111.295 131.080 ;
        RECT 108.895 130.345 109.825 130.515 ;
        RECT 108.895 130.310 109.070 130.345 ;
        RECT 108.540 129.945 109.070 130.310 ;
        RECT 109.495 129.775 109.825 130.175 ;
        RECT 109.995 129.945 110.250 130.515 ;
        RECT 111.010 130.495 111.180 130.750 ;
        RECT 110.515 130.325 111.180 130.495 ;
        RECT 111.465 130.450 111.635 131.250 ;
        RECT 112.725 131.565 113.240 131.975 ;
        RECT 113.475 131.565 113.645 132.325 ;
        RECT 113.815 131.985 115.845 132.155 ;
        RECT 112.725 130.755 113.065 131.565 ;
        RECT 113.815 131.320 113.985 131.985 ;
        RECT 114.380 131.645 115.505 131.815 ;
        RECT 113.235 131.130 113.985 131.320 ;
        RECT 114.155 131.305 115.165 131.475 ;
        RECT 112.725 130.585 113.955 130.755 ;
        RECT 110.515 129.945 110.685 130.325 ;
        RECT 110.865 129.775 111.195 130.155 ;
        RECT 111.375 129.945 111.635 130.450 ;
        RECT 113.000 129.980 113.245 130.585 ;
        RECT 113.465 129.775 113.975 130.310 ;
        RECT 114.155 129.945 114.345 131.305 ;
        RECT 114.515 130.285 114.790 131.105 ;
        RECT 114.995 130.505 115.165 131.305 ;
        RECT 115.335 130.515 115.505 131.645 ;
        RECT 115.675 131.015 115.845 131.985 ;
        RECT 116.015 131.185 116.185 132.325 ;
        RECT 116.355 131.185 116.690 132.155 ;
        RECT 117.365 131.185 117.595 132.325 ;
        RECT 115.675 130.685 115.870 131.015 ;
        RECT 116.095 130.685 116.350 131.015 ;
        RECT 116.095 130.515 116.265 130.685 ;
        RECT 116.520 130.515 116.690 131.185 ;
        RECT 117.765 131.175 118.095 132.155 ;
        RECT 118.265 131.185 118.475 132.325 ;
        RECT 118.795 131.395 118.965 132.155 ;
        RECT 119.145 131.565 119.475 132.325 ;
        RECT 118.795 131.225 119.460 131.395 ;
        RECT 119.645 131.250 119.915 132.155 ;
        RECT 121.010 131.890 126.355 132.325 ;
        RECT 117.345 130.765 117.675 131.015 ;
        RECT 115.335 130.345 116.265 130.515 ;
        RECT 115.335 130.310 115.510 130.345 ;
        RECT 114.515 130.115 114.795 130.285 ;
        RECT 114.515 129.945 114.790 130.115 ;
        RECT 114.980 129.945 115.510 130.310 ;
        RECT 115.935 129.775 116.265 130.175 ;
        RECT 116.435 129.945 116.690 130.515 ;
        RECT 117.365 129.775 117.595 130.595 ;
        RECT 117.845 130.575 118.095 131.175 ;
        RECT 119.290 131.080 119.460 131.225 ;
        RECT 118.725 130.675 119.055 131.045 ;
        RECT 119.290 130.750 119.575 131.080 ;
        RECT 117.765 129.945 118.095 130.575 ;
        RECT 118.265 129.775 118.475 130.595 ;
        RECT 119.290 130.495 119.460 130.750 ;
        RECT 118.795 130.325 119.460 130.495 ;
        RECT 119.745 130.450 119.915 131.250 ;
        RECT 122.600 130.640 122.950 131.890 ;
        RECT 126.525 131.235 127.735 132.325 ;
        RECT 118.795 129.945 118.965 130.325 ;
        RECT 119.145 129.775 119.475 130.155 ;
        RECT 119.655 129.945 119.915 130.450 ;
        RECT 124.430 130.320 124.770 131.150 ;
        RECT 126.525 130.695 127.045 131.235 ;
        RECT 127.215 130.525 127.735 131.065 ;
        RECT 121.010 129.775 126.355 130.320 ;
        RECT 126.525 129.775 127.735 130.525 ;
        RECT 29.840 129.605 127.820 129.775 ;
        RECT 29.925 128.855 31.135 129.605 ;
        RECT 29.925 128.315 30.445 128.855 ;
        RECT 31.765 128.835 35.275 129.605 ;
        RECT 30.615 128.145 31.135 128.685 ;
        RECT 29.925 127.055 31.135 128.145 ;
        RECT 31.765 128.145 33.455 128.665 ;
        RECT 33.625 128.315 35.275 128.835 ;
        RECT 35.485 128.785 35.715 129.605 ;
        RECT 35.885 128.805 36.215 129.435 ;
        RECT 35.465 128.365 35.795 128.615 ;
        RECT 35.965 128.205 36.215 128.805 ;
        RECT 36.385 128.785 36.595 129.605 ;
        RECT 37.285 128.880 37.575 129.605 ;
        RECT 38.295 129.055 38.465 129.435 ;
        RECT 38.645 129.225 38.975 129.605 ;
        RECT 38.295 128.885 38.960 129.055 ;
        RECT 39.155 128.930 39.415 129.435 ;
        RECT 38.225 128.335 38.555 128.705 ;
        RECT 38.790 128.630 38.960 128.885 ;
        RECT 38.790 128.300 39.075 128.630 ;
        RECT 31.765 127.055 35.275 128.145 ;
        RECT 35.485 127.055 35.715 128.195 ;
        RECT 35.885 127.225 36.215 128.205 ;
        RECT 36.385 127.055 36.595 128.195 ;
        RECT 37.285 127.055 37.575 128.220 ;
        RECT 38.790 128.155 38.960 128.300 ;
        RECT 38.295 127.985 38.960 128.155 ;
        RECT 39.245 128.130 39.415 128.930 ;
        RECT 39.625 128.785 39.855 129.605 ;
        RECT 40.025 128.805 40.355 129.435 ;
        RECT 39.605 128.365 39.935 128.615 ;
        RECT 40.105 128.205 40.355 128.805 ;
        RECT 40.525 128.785 40.735 129.605 ;
        RECT 41.055 129.055 41.225 129.435 ;
        RECT 41.405 129.225 41.735 129.605 ;
        RECT 41.055 128.885 41.720 129.055 ;
        RECT 41.915 128.930 42.175 129.435 ;
        RECT 40.985 128.335 41.315 128.705 ;
        RECT 41.550 128.630 41.720 128.885 ;
        RECT 38.295 127.225 38.465 127.985 ;
        RECT 38.645 127.055 38.975 127.815 ;
        RECT 39.145 127.225 39.415 128.130 ;
        RECT 39.625 127.055 39.855 128.195 ;
        RECT 40.025 127.225 40.355 128.205 ;
        RECT 41.550 128.300 41.835 128.630 ;
        RECT 40.525 127.055 40.735 128.195 ;
        RECT 41.550 128.155 41.720 128.300 ;
        RECT 41.055 127.985 41.720 128.155 ;
        RECT 42.005 128.130 42.175 128.930 ;
        RECT 42.385 128.785 42.615 129.605 ;
        RECT 42.785 128.805 43.115 129.435 ;
        RECT 42.365 128.365 42.695 128.615 ;
        RECT 42.865 128.205 43.115 128.805 ;
        RECT 43.285 128.785 43.495 129.605 ;
        RECT 44.100 128.895 44.355 129.425 ;
        RECT 44.535 129.145 44.820 129.605 ;
        RECT 41.055 127.225 41.225 127.985 ;
        RECT 41.405 127.055 41.735 127.815 ;
        RECT 41.905 127.225 42.175 128.130 ;
        RECT 42.385 127.055 42.615 128.195 ;
        RECT 42.785 127.225 43.115 128.205 ;
        RECT 43.285 127.055 43.495 128.195 ;
        RECT 44.100 128.035 44.280 128.895 ;
        RECT 45.000 128.695 45.250 129.345 ;
        RECT 44.450 128.365 45.250 128.695 ;
        RECT 44.100 127.565 44.355 128.035 ;
        RECT 44.015 127.395 44.355 127.565 ;
        RECT 44.100 127.365 44.355 127.395 ;
        RECT 44.535 127.055 44.820 127.855 ;
        RECT 45.000 127.775 45.250 128.365 ;
        RECT 45.450 129.010 45.770 129.340 ;
        RECT 45.950 129.125 46.610 129.605 ;
        RECT 46.810 129.215 47.660 129.385 ;
        RECT 45.450 128.115 45.640 129.010 ;
        RECT 45.960 128.685 46.620 128.955 ;
        RECT 46.290 128.625 46.620 128.685 ;
        RECT 45.810 128.455 46.140 128.515 ;
        RECT 46.810 128.455 46.980 129.215 ;
        RECT 48.220 129.145 48.540 129.605 ;
        RECT 48.740 128.965 48.990 129.395 ;
        RECT 49.280 129.165 49.690 129.605 ;
        RECT 49.860 129.225 50.875 129.425 ;
        RECT 47.150 128.795 48.400 128.965 ;
        RECT 47.150 128.675 47.480 128.795 ;
        RECT 45.810 128.285 47.710 128.455 ;
        RECT 45.450 127.945 47.370 128.115 ;
        RECT 45.450 127.925 45.770 127.945 ;
        RECT 45.000 127.265 45.330 127.775 ;
        RECT 45.600 127.315 45.770 127.925 ;
        RECT 47.540 127.775 47.710 128.285 ;
        RECT 47.880 128.215 48.060 128.625 ;
        RECT 48.230 128.035 48.400 128.795 ;
        RECT 45.940 127.055 46.270 127.745 ;
        RECT 46.500 127.605 47.710 127.775 ;
        RECT 47.880 127.725 48.400 128.035 ;
        RECT 48.570 128.625 48.990 128.965 ;
        RECT 49.280 128.625 49.690 128.955 ;
        RECT 48.570 127.855 48.760 128.625 ;
        RECT 49.860 128.495 50.030 129.225 ;
        RECT 51.175 129.055 51.345 129.385 ;
        RECT 51.515 129.225 51.845 129.605 ;
        RECT 50.200 128.675 50.550 129.045 ;
        RECT 49.860 128.455 50.280 128.495 ;
        RECT 48.930 128.285 50.280 128.455 ;
        RECT 48.930 128.125 49.180 128.285 ;
        RECT 49.690 127.855 49.940 128.115 ;
        RECT 48.570 127.605 49.940 127.855 ;
        RECT 46.500 127.315 46.740 127.605 ;
        RECT 47.540 127.525 47.710 127.605 ;
        RECT 46.940 127.055 47.360 127.435 ;
        RECT 47.540 127.275 48.170 127.525 ;
        RECT 48.640 127.055 48.970 127.435 ;
        RECT 49.140 127.315 49.310 127.605 ;
        RECT 50.110 127.440 50.280 128.285 ;
        RECT 50.730 128.115 50.950 128.985 ;
        RECT 51.175 128.865 51.870 129.055 ;
        RECT 50.450 127.735 50.950 128.115 ;
        RECT 51.120 128.065 51.530 128.685 ;
        RECT 51.700 127.895 51.870 128.865 ;
        RECT 51.175 127.725 51.870 127.895 ;
        RECT 49.490 127.055 49.870 127.435 ;
        RECT 50.110 127.270 50.940 127.440 ;
        RECT 51.175 127.225 51.345 127.725 ;
        RECT 51.515 127.055 51.845 127.555 ;
        RECT 52.060 127.225 52.285 129.345 ;
        RECT 52.455 129.225 52.785 129.605 ;
        RECT 52.955 129.055 53.125 129.345 ;
        RECT 53.760 129.265 54.015 129.425 ;
        RECT 53.675 129.095 54.015 129.265 ;
        RECT 54.195 129.145 54.480 129.605 ;
        RECT 52.460 128.885 53.125 129.055 ;
        RECT 53.760 128.895 54.015 129.095 ;
        RECT 52.460 127.895 52.690 128.885 ;
        RECT 52.860 128.065 53.210 128.715 ;
        RECT 53.760 128.035 53.940 128.895 ;
        RECT 54.660 128.695 54.910 129.345 ;
        RECT 54.110 128.365 54.910 128.695 ;
        RECT 52.460 127.725 53.125 127.895 ;
        RECT 52.455 127.055 52.785 127.555 ;
        RECT 52.955 127.225 53.125 127.725 ;
        RECT 53.760 127.365 54.015 128.035 ;
        RECT 54.195 127.055 54.480 127.855 ;
        RECT 54.660 127.775 54.910 128.365 ;
        RECT 55.110 129.010 55.430 129.340 ;
        RECT 55.610 129.125 56.270 129.605 ;
        RECT 56.470 129.215 57.320 129.385 ;
        RECT 55.110 128.115 55.300 129.010 ;
        RECT 55.620 128.685 56.280 128.955 ;
        RECT 55.950 128.625 56.280 128.685 ;
        RECT 55.470 128.455 55.800 128.515 ;
        RECT 56.470 128.455 56.640 129.215 ;
        RECT 57.880 129.145 58.200 129.605 ;
        RECT 58.400 128.965 58.650 129.395 ;
        RECT 58.940 129.165 59.350 129.605 ;
        RECT 59.520 129.225 60.535 129.425 ;
        RECT 56.810 128.795 58.060 128.965 ;
        RECT 56.810 128.675 57.140 128.795 ;
        RECT 55.470 128.285 57.370 128.455 ;
        RECT 55.110 127.945 57.030 128.115 ;
        RECT 55.110 127.925 55.430 127.945 ;
        RECT 54.660 127.265 54.990 127.775 ;
        RECT 55.260 127.315 55.430 127.925 ;
        RECT 57.200 127.775 57.370 128.285 ;
        RECT 57.540 128.215 57.720 128.625 ;
        RECT 57.890 128.035 58.060 128.795 ;
        RECT 55.600 127.055 55.930 127.745 ;
        RECT 56.160 127.605 57.370 127.775 ;
        RECT 57.540 127.725 58.060 128.035 ;
        RECT 58.230 128.625 58.650 128.965 ;
        RECT 58.940 128.625 59.350 128.955 ;
        RECT 58.230 127.855 58.420 128.625 ;
        RECT 59.520 128.495 59.690 129.225 ;
        RECT 60.835 129.055 61.005 129.385 ;
        RECT 61.175 129.225 61.505 129.605 ;
        RECT 59.860 128.675 60.210 129.045 ;
        RECT 59.520 128.455 59.940 128.495 ;
        RECT 58.590 128.285 59.940 128.455 ;
        RECT 58.590 128.125 58.840 128.285 ;
        RECT 59.350 127.855 59.600 128.115 ;
        RECT 58.230 127.605 59.600 127.855 ;
        RECT 56.160 127.315 56.400 127.605 ;
        RECT 57.200 127.525 57.370 127.605 ;
        RECT 56.600 127.055 57.020 127.435 ;
        RECT 57.200 127.275 57.830 127.525 ;
        RECT 58.300 127.055 58.630 127.435 ;
        RECT 58.800 127.315 58.970 127.605 ;
        RECT 59.770 127.440 59.940 128.285 ;
        RECT 60.390 128.115 60.610 128.985 ;
        RECT 60.835 128.865 61.530 129.055 ;
        RECT 60.110 127.735 60.610 128.115 ;
        RECT 60.780 128.065 61.190 128.685 ;
        RECT 61.360 127.895 61.530 128.865 ;
        RECT 60.835 127.725 61.530 127.895 ;
        RECT 59.150 127.055 59.530 127.435 ;
        RECT 59.770 127.270 60.600 127.440 ;
        RECT 60.835 127.225 61.005 127.725 ;
        RECT 61.175 127.055 61.505 127.555 ;
        RECT 61.720 127.225 61.945 129.345 ;
        RECT 62.115 129.225 62.445 129.605 ;
        RECT 62.615 129.055 62.785 129.345 ;
        RECT 62.120 128.885 62.785 129.055 ;
        RECT 62.120 127.895 62.350 128.885 ;
        RECT 63.045 128.880 63.335 129.605 ;
        RECT 63.505 128.930 63.765 129.435 ;
        RECT 63.945 129.225 64.275 129.605 ;
        RECT 64.455 129.055 64.625 129.435 ;
        RECT 62.520 128.065 62.870 128.715 ;
        RECT 62.120 127.725 62.785 127.895 ;
        RECT 62.115 127.055 62.445 127.555 ;
        RECT 62.615 127.225 62.785 127.725 ;
        RECT 63.045 127.055 63.335 128.220 ;
        RECT 63.505 128.130 63.675 128.930 ;
        RECT 63.960 128.885 64.625 129.055 ;
        RECT 63.960 128.630 64.130 128.885 ;
        RECT 64.945 128.785 65.155 129.605 ;
        RECT 65.325 128.805 65.655 129.435 ;
        RECT 63.845 128.300 64.130 128.630 ;
        RECT 64.365 128.335 64.695 128.705 ;
        RECT 63.960 128.155 64.130 128.300 ;
        RECT 65.325 128.205 65.575 128.805 ;
        RECT 65.825 128.785 66.055 129.605 ;
        RECT 66.355 129.055 66.525 129.435 ;
        RECT 66.705 129.225 67.035 129.605 ;
        RECT 66.355 128.885 67.020 129.055 ;
        RECT 67.215 128.930 67.475 129.435 ;
        RECT 68.480 129.265 68.735 129.425 ;
        RECT 68.395 129.095 68.735 129.265 ;
        RECT 68.915 129.145 69.200 129.605 ;
        RECT 65.745 128.365 66.075 128.615 ;
        RECT 66.285 128.335 66.615 128.705 ;
        RECT 66.850 128.630 67.020 128.885 ;
        RECT 66.850 128.300 67.135 128.630 ;
        RECT 63.505 127.225 63.775 128.130 ;
        RECT 63.960 127.985 64.625 128.155 ;
        RECT 63.945 127.055 64.275 127.815 ;
        RECT 64.455 127.225 64.625 127.985 ;
        RECT 64.945 127.055 65.155 128.195 ;
        RECT 65.325 127.225 65.655 128.205 ;
        RECT 65.825 127.055 66.055 128.195 ;
        RECT 66.850 128.155 67.020 128.300 ;
        RECT 66.355 127.985 67.020 128.155 ;
        RECT 67.305 128.130 67.475 128.930 ;
        RECT 66.355 127.225 66.525 127.985 ;
        RECT 66.705 127.055 67.035 127.815 ;
        RECT 67.205 127.225 67.475 128.130 ;
        RECT 68.480 128.895 68.735 129.095 ;
        RECT 68.480 128.035 68.660 128.895 ;
        RECT 69.380 128.695 69.630 129.345 ;
        RECT 68.830 128.365 69.630 128.695 ;
        RECT 68.480 127.365 68.735 128.035 ;
        RECT 68.915 127.055 69.200 127.855 ;
        RECT 69.380 127.775 69.630 128.365 ;
        RECT 69.830 129.010 70.150 129.340 ;
        RECT 70.330 129.125 70.990 129.605 ;
        RECT 71.190 129.215 72.040 129.385 ;
        RECT 69.830 128.115 70.020 129.010 ;
        RECT 70.340 128.685 71.000 128.955 ;
        RECT 70.670 128.625 71.000 128.685 ;
        RECT 70.190 128.455 70.520 128.515 ;
        RECT 71.190 128.455 71.360 129.215 ;
        RECT 72.600 129.145 72.920 129.605 ;
        RECT 73.120 128.965 73.370 129.395 ;
        RECT 73.660 129.165 74.070 129.605 ;
        RECT 74.240 129.225 75.255 129.425 ;
        RECT 71.530 128.795 72.780 128.965 ;
        RECT 71.530 128.675 71.860 128.795 ;
        RECT 70.190 128.285 72.090 128.455 ;
        RECT 69.830 127.945 71.750 128.115 ;
        RECT 69.830 127.925 70.150 127.945 ;
        RECT 69.380 127.265 69.710 127.775 ;
        RECT 69.980 127.315 70.150 127.925 ;
        RECT 71.920 127.775 72.090 128.285 ;
        RECT 72.260 128.215 72.440 128.625 ;
        RECT 72.610 128.035 72.780 128.795 ;
        RECT 70.320 127.055 70.650 127.745 ;
        RECT 70.880 127.605 72.090 127.775 ;
        RECT 72.260 127.725 72.780 128.035 ;
        RECT 72.950 128.625 73.370 128.965 ;
        RECT 73.660 128.625 74.070 128.955 ;
        RECT 72.950 127.855 73.140 128.625 ;
        RECT 74.240 128.495 74.410 129.225 ;
        RECT 75.555 129.055 75.725 129.385 ;
        RECT 75.895 129.225 76.225 129.605 ;
        RECT 74.580 128.675 74.930 129.045 ;
        RECT 74.240 128.455 74.660 128.495 ;
        RECT 73.310 128.285 74.660 128.455 ;
        RECT 73.310 128.125 73.560 128.285 ;
        RECT 74.070 127.855 74.320 128.115 ;
        RECT 72.950 127.605 74.320 127.855 ;
        RECT 70.880 127.315 71.120 127.605 ;
        RECT 71.920 127.525 72.090 127.605 ;
        RECT 71.320 127.055 71.740 127.435 ;
        RECT 71.920 127.275 72.550 127.525 ;
        RECT 73.020 127.055 73.350 127.435 ;
        RECT 73.520 127.315 73.690 127.605 ;
        RECT 74.490 127.440 74.660 128.285 ;
        RECT 75.110 128.115 75.330 128.985 ;
        RECT 75.555 128.865 76.250 129.055 ;
        RECT 74.830 127.735 75.330 128.115 ;
        RECT 75.500 128.065 75.910 128.685 ;
        RECT 76.080 127.895 76.250 128.865 ;
        RECT 75.555 127.725 76.250 127.895 ;
        RECT 73.870 127.055 74.250 127.435 ;
        RECT 74.490 127.270 75.320 127.440 ;
        RECT 75.555 127.225 75.725 127.725 ;
        RECT 75.895 127.055 76.225 127.555 ;
        RECT 76.440 127.225 76.665 129.345 ;
        RECT 76.835 129.225 77.165 129.605 ;
        RECT 77.335 129.055 77.505 129.345 ;
        RECT 76.840 128.885 77.505 129.055 ;
        RECT 76.840 127.895 77.070 128.885 ;
        RECT 77.765 128.855 78.975 129.605 ;
        RECT 79.520 129.265 79.775 129.425 ;
        RECT 79.435 129.095 79.775 129.265 ;
        RECT 79.955 129.145 80.240 129.605 ;
        RECT 77.240 128.065 77.590 128.715 ;
        RECT 77.765 128.145 78.285 128.685 ;
        RECT 78.455 128.315 78.975 128.855 ;
        RECT 79.520 128.895 79.775 129.095 ;
        RECT 76.840 127.725 77.505 127.895 ;
        RECT 76.835 127.055 77.165 127.555 ;
        RECT 77.335 127.225 77.505 127.725 ;
        RECT 77.765 127.055 78.975 128.145 ;
        RECT 79.520 128.035 79.700 128.895 ;
        RECT 80.420 128.695 80.670 129.345 ;
        RECT 79.870 128.365 80.670 128.695 ;
        RECT 79.520 127.365 79.775 128.035 ;
        RECT 79.955 127.055 80.240 127.855 ;
        RECT 80.420 127.775 80.670 128.365 ;
        RECT 80.870 129.010 81.190 129.340 ;
        RECT 81.370 129.125 82.030 129.605 ;
        RECT 82.230 129.215 83.080 129.385 ;
        RECT 80.870 128.115 81.060 129.010 ;
        RECT 81.380 128.685 82.040 128.955 ;
        RECT 81.710 128.625 82.040 128.685 ;
        RECT 81.230 128.455 81.560 128.515 ;
        RECT 82.230 128.455 82.400 129.215 ;
        RECT 83.640 129.145 83.960 129.605 ;
        RECT 84.160 128.965 84.410 129.395 ;
        RECT 84.700 129.165 85.110 129.605 ;
        RECT 85.280 129.225 86.295 129.425 ;
        RECT 82.570 128.795 83.820 128.965 ;
        RECT 82.570 128.675 82.900 128.795 ;
        RECT 81.230 128.285 83.130 128.455 ;
        RECT 80.870 127.945 82.790 128.115 ;
        RECT 80.870 127.925 81.190 127.945 ;
        RECT 80.420 127.265 80.750 127.775 ;
        RECT 81.020 127.315 81.190 127.925 ;
        RECT 82.960 127.775 83.130 128.285 ;
        RECT 83.300 128.215 83.480 128.625 ;
        RECT 83.650 128.035 83.820 128.795 ;
        RECT 81.360 127.055 81.690 127.745 ;
        RECT 81.920 127.605 83.130 127.775 ;
        RECT 83.300 127.725 83.820 128.035 ;
        RECT 83.990 128.625 84.410 128.965 ;
        RECT 84.700 128.625 85.110 128.955 ;
        RECT 83.990 127.855 84.180 128.625 ;
        RECT 85.280 128.495 85.450 129.225 ;
        RECT 86.595 129.055 86.765 129.385 ;
        RECT 86.935 129.225 87.265 129.605 ;
        RECT 85.620 128.675 85.970 129.045 ;
        RECT 85.280 128.455 85.700 128.495 ;
        RECT 84.350 128.285 85.700 128.455 ;
        RECT 84.350 128.125 84.600 128.285 ;
        RECT 85.110 127.855 85.360 128.115 ;
        RECT 83.990 127.605 85.360 127.855 ;
        RECT 81.920 127.315 82.160 127.605 ;
        RECT 82.960 127.525 83.130 127.605 ;
        RECT 82.360 127.055 82.780 127.435 ;
        RECT 82.960 127.275 83.590 127.525 ;
        RECT 84.060 127.055 84.390 127.435 ;
        RECT 84.560 127.315 84.730 127.605 ;
        RECT 85.530 127.440 85.700 128.285 ;
        RECT 86.150 128.115 86.370 128.985 ;
        RECT 86.595 128.865 87.290 129.055 ;
        RECT 85.870 127.735 86.370 128.115 ;
        RECT 86.540 128.065 86.950 128.685 ;
        RECT 87.120 127.895 87.290 128.865 ;
        RECT 86.595 127.725 87.290 127.895 ;
        RECT 84.910 127.055 85.290 127.435 ;
        RECT 85.530 127.270 86.360 127.440 ;
        RECT 86.595 127.225 86.765 127.725 ;
        RECT 86.935 127.055 87.265 127.555 ;
        RECT 87.480 127.225 87.705 129.345 ;
        RECT 87.875 129.225 88.205 129.605 ;
        RECT 88.375 129.055 88.545 129.345 ;
        RECT 87.880 128.885 88.545 129.055 ;
        RECT 87.880 127.895 88.110 128.885 ;
        RECT 88.805 128.880 89.095 129.605 ;
        RECT 89.640 129.265 89.895 129.425 ;
        RECT 89.555 129.095 89.895 129.265 ;
        RECT 90.075 129.145 90.360 129.605 ;
        RECT 89.640 128.895 89.895 129.095 ;
        RECT 88.280 128.065 88.630 128.715 ;
        RECT 87.880 127.725 88.545 127.895 ;
        RECT 87.875 127.055 88.205 127.555 ;
        RECT 88.375 127.225 88.545 127.725 ;
        RECT 88.805 127.055 89.095 128.220 ;
        RECT 89.640 128.035 89.820 128.895 ;
        RECT 90.540 128.695 90.790 129.345 ;
        RECT 89.990 128.365 90.790 128.695 ;
        RECT 89.640 127.365 89.895 128.035 ;
        RECT 90.075 127.055 90.360 127.855 ;
        RECT 90.540 127.775 90.790 128.365 ;
        RECT 90.990 129.010 91.310 129.340 ;
        RECT 91.490 129.125 92.150 129.605 ;
        RECT 92.350 129.215 93.200 129.385 ;
        RECT 90.990 128.115 91.180 129.010 ;
        RECT 91.500 128.685 92.160 128.955 ;
        RECT 91.830 128.625 92.160 128.685 ;
        RECT 91.350 128.455 91.680 128.515 ;
        RECT 92.350 128.455 92.520 129.215 ;
        RECT 93.760 129.145 94.080 129.605 ;
        RECT 94.280 128.965 94.530 129.395 ;
        RECT 94.820 129.165 95.230 129.605 ;
        RECT 95.400 129.225 96.415 129.425 ;
        RECT 92.690 128.795 93.940 128.965 ;
        RECT 92.690 128.675 93.020 128.795 ;
        RECT 91.350 128.285 93.250 128.455 ;
        RECT 90.990 127.945 92.910 128.115 ;
        RECT 90.990 127.925 91.310 127.945 ;
        RECT 90.540 127.265 90.870 127.775 ;
        RECT 91.140 127.315 91.310 127.925 ;
        RECT 93.080 127.775 93.250 128.285 ;
        RECT 93.420 128.215 93.600 128.625 ;
        RECT 93.770 128.035 93.940 128.795 ;
        RECT 91.480 127.055 91.810 127.745 ;
        RECT 92.040 127.605 93.250 127.775 ;
        RECT 93.420 127.725 93.940 128.035 ;
        RECT 94.110 128.625 94.530 128.965 ;
        RECT 94.820 128.625 95.230 128.955 ;
        RECT 94.110 127.855 94.300 128.625 ;
        RECT 95.400 128.495 95.570 129.225 ;
        RECT 96.715 129.055 96.885 129.385 ;
        RECT 97.055 129.225 97.385 129.605 ;
        RECT 95.740 128.675 96.090 129.045 ;
        RECT 95.400 128.455 95.820 128.495 ;
        RECT 94.470 128.285 95.820 128.455 ;
        RECT 94.470 128.125 94.720 128.285 ;
        RECT 95.230 127.855 95.480 128.115 ;
        RECT 94.110 127.605 95.480 127.855 ;
        RECT 92.040 127.315 92.280 127.605 ;
        RECT 93.080 127.525 93.250 127.605 ;
        RECT 92.480 127.055 92.900 127.435 ;
        RECT 93.080 127.275 93.710 127.525 ;
        RECT 94.180 127.055 94.510 127.435 ;
        RECT 94.680 127.315 94.850 127.605 ;
        RECT 95.650 127.440 95.820 128.285 ;
        RECT 96.270 128.115 96.490 128.985 ;
        RECT 96.715 128.865 97.410 129.055 ;
        RECT 95.990 127.735 96.490 128.115 ;
        RECT 96.660 128.065 97.070 128.685 ;
        RECT 97.240 127.895 97.410 128.865 ;
        RECT 96.715 127.725 97.410 127.895 ;
        RECT 95.030 127.055 95.410 127.435 ;
        RECT 95.650 127.270 96.480 127.440 ;
        RECT 96.715 127.225 96.885 127.725 ;
        RECT 97.055 127.055 97.385 127.555 ;
        RECT 97.600 127.225 97.825 129.345 ;
        RECT 97.995 129.225 98.325 129.605 ;
        RECT 98.495 129.055 98.665 129.345 ;
        RECT 98.000 128.885 98.665 129.055 ;
        RECT 99.385 128.930 99.645 129.435 ;
        RECT 99.825 129.225 100.155 129.605 ;
        RECT 100.335 129.055 100.505 129.435 ;
        RECT 98.000 127.895 98.230 128.885 ;
        RECT 98.400 128.065 98.750 128.715 ;
        RECT 99.385 128.130 99.555 128.930 ;
        RECT 99.840 128.885 100.505 129.055 ;
        RECT 99.840 128.630 100.010 128.885 ;
        RECT 101.225 128.835 104.735 129.605 ;
        RECT 105.280 129.265 105.535 129.425 ;
        RECT 105.195 129.095 105.535 129.265 ;
        RECT 105.715 129.145 106.000 129.605 ;
        RECT 99.725 128.300 100.010 128.630 ;
        RECT 100.245 128.335 100.575 128.705 ;
        RECT 99.840 128.155 100.010 128.300 ;
        RECT 98.000 127.725 98.665 127.895 ;
        RECT 97.995 127.055 98.325 127.555 ;
        RECT 98.495 127.225 98.665 127.725 ;
        RECT 99.385 127.225 99.655 128.130 ;
        RECT 99.840 127.985 100.505 128.155 ;
        RECT 99.825 127.055 100.155 127.815 ;
        RECT 100.335 127.225 100.505 127.985 ;
        RECT 101.225 128.145 102.915 128.665 ;
        RECT 103.085 128.315 104.735 128.835 ;
        RECT 105.280 128.895 105.535 129.095 ;
        RECT 101.225 127.055 104.735 128.145 ;
        RECT 105.280 128.035 105.460 128.895 ;
        RECT 106.180 128.695 106.430 129.345 ;
        RECT 105.630 128.365 106.430 128.695 ;
        RECT 105.280 127.365 105.535 128.035 ;
        RECT 105.715 127.055 106.000 127.855 ;
        RECT 106.180 127.775 106.430 128.365 ;
        RECT 106.630 129.010 106.950 129.340 ;
        RECT 107.130 129.125 107.790 129.605 ;
        RECT 107.990 129.215 108.840 129.385 ;
        RECT 106.630 128.115 106.820 129.010 ;
        RECT 107.140 128.685 107.800 128.955 ;
        RECT 107.470 128.625 107.800 128.685 ;
        RECT 106.990 128.455 107.320 128.515 ;
        RECT 107.990 128.455 108.160 129.215 ;
        RECT 109.400 129.145 109.720 129.605 ;
        RECT 109.920 128.965 110.170 129.395 ;
        RECT 110.460 129.165 110.870 129.605 ;
        RECT 111.040 129.225 112.055 129.425 ;
        RECT 108.330 128.795 109.580 128.965 ;
        RECT 108.330 128.675 108.660 128.795 ;
        RECT 106.990 128.285 108.890 128.455 ;
        RECT 106.630 127.945 108.550 128.115 ;
        RECT 106.630 127.925 106.950 127.945 ;
        RECT 106.180 127.265 106.510 127.775 ;
        RECT 106.780 127.315 106.950 127.925 ;
        RECT 108.720 127.775 108.890 128.285 ;
        RECT 109.060 128.215 109.240 128.625 ;
        RECT 109.410 128.035 109.580 128.795 ;
        RECT 107.120 127.055 107.450 127.745 ;
        RECT 107.680 127.605 108.890 127.775 ;
        RECT 109.060 127.725 109.580 128.035 ;
        RECT 109.750 128.625 110.170 128.965 ;
        RECT 110.460 128.625 110.870 128.955 ;
        RECT 109.750 127.855 109.940 128.625 ;
        RECT 111.040 128.495 111.210 129.225 ;
        RECT 112.355 129.055 112.525 129.385 ;
        RECT 112.695 129.225 113.025 129.605 ;
        RECT 111.380 128.675 111.730 129.045 ;
        RECT 111.040 128.455 111.460 128.495 ;
        RECT 110.110 128.285 111.460 128.455 ;
        RECT 110.110 128.125 110.360 128.285 ;
        RECT 110.870 127.855 111.120 128.115 ;
        RECT 109.750 127.605 111.120 127.855 ;
        RECT 107.680 127.315 107.920 127.605 ;
        RECT 108.720 127.525 108.890 127.605 ;
        RECT 108.120 127.055 108.540 127.435 ;
        RECT 108.720 127.275 109.350 127.525 ;
        RECT 109.820 127.055 110.150 127.435 ;
        RECT 110.320 127.315 110.490 127.605 ;
        RECT 111.290 127.440 111.460 128.285 ;
        RECT 111.910 128.115 112.130 128.985 ;
        RECT 112.355 128.865 113.050 129.055 ;
        RECT 111.630 127.735 112.130 128.115 ;
        RECT 112.300 128.065 112.710 128.685 ;
        RECT 112.880 127.895 113.050 128.865 ;
        RECT 112.355 127.725 113.050 127.895 ;
        RECT 110.670 127.055 111.050 127.435 ;
        RECT 111.290 127.270 112.120 127.440 ;
        RECT 112.355 127.225 112.525 127.725 ;
        RECT 112.695 127.055 113.025 127.555 ;
        RECT 113.240 127.225 113.465 129.345 ;
        RECT 113.635 129.225 113.965 129.605 ;
        RECT 114.135 129.055 114.305 129.345 ;
        RECT 113.640 128.885 114.305 129.055 ;
        RECT 113.640 127.895 113.870 128.885 ;
        RECT 114.565 128.880 114.855 129.605 ;
        RECT 115.400 129.265 115.655 129.425 ;
        RECT 115.315 129.095 115.655 129.265 ;
        RECT 115.835 129.145 116.120 129.605 ;
        RECT 115.400 128.895 115.655 129.095 ;
        RECT 114.040 128.065 114.390 128.715 ;
        RECT 113.640 127.725 114.305 127.895 ;
        RECT 113.635 127.055 113.965 127.555 ;
        RECT 114.135 127.225 114.305 127.725 ;
        RECT 114.565 127.055 114.855 128.220 ;
        RECT 115.400 128.035 115.580 128.895 ;
        RECT 116.300 128.695 116.550 129.345 ;
        RECT 115.750 128.365 116.550 128.695 ;
        RECT 115.400 127.365 115.655 128.035 ;
        RECT 115.835 127.055 116.120 127.855 ;
        RECT 116.300 127.775 116.550 128.365 ;
        RECT 116.750 129.010 117.070 129.340 ;
        RECT 117.250 129.125 117.910 129.605 ;
        RECT 118.110 129.215 118.960 129.385 ;
        RECT 116.750 128.115 116.940 129.010 ;
        RECT 117.260 128.685 117.920 128.955 ;
        RECT 117.590 128.625 117.920 128.685 ;
        RECT 117.110 128.455 117.440 128.515 ;
        RECT 118.110 128.455 118.280 129.215 ;
        RECT 119.520 129.145 119.840 129.605 ;
        RECT 120.040 128.965 120.290 129.395 ;
        RECT 120.580 129.165 120.990 129.605 ;
        RECT 121.160 129.225 122.175 129.425 ;
        RECT 118.450 128.795 119.700 128.965 ;
        RECT 118.450 128.675 118.780 128.795 ;
        RECT 117.110 128.285 119.010 128.455 ;
        RECT 116.750 127.945 118.670 128.115 ;
        RECT 116.750 127.925 117.070 127.945 ;
        RECT 116.300 127.265 116.630 127.775 ;
        RECT 116.900 127.315 117.070 127.925 ;
        RECT 118.840 127.775 119.010 128.285 ;
        RECT 119.180 128.215 119.360 128.625 ;
        RECT 119.530 128.035 119.700 128.795 ;
        RECT 117.240 127.055 117.570 127.745 ;
        RECT 117.800 127.605 119.010 127.775 ;
        RECT 119.180 127.725 119.700 128.035 ;
        RECT 119.870 128.625 120.290 128.965 ;
        RECT 120.580 128.625 120.990 128.955 ;
        RECT 119.870 127.855 120.060 128.625 ;
        RECT 121.160 128.495 121.330 129.225 ;
        RECT 122.475 129.055 122.645 129.385 ;
        RECT 122.815 129.225 123.145 129.605 ;
        RECT 121.500 128.675 121.850 129.045 ;
        RECT 121.160 128.455 121.580 128.495 ;
        RECT 120.230 128.285 121.580 128.455 ;
        RECT 120.230 128.125 120.480 128.285 ;
        RECT 120.990 127.855 121.240 128.115 ;
        RECT 119.870 127.605 121.240 127.855 ;
        RECT 117.800 127.315 118.040 127.605 ;
        RECT 118.840 127.525 119.010 127.605 ;
        RECT 118.240 127.055 118.660 127.435 ;
        RECT 118.840 127.275 119.470 127.525 ;
        RECT 119.940 127.055 120.270 127.435 ;
        RECT 120.440 127.315 120.610 127.605 ;
        RECT 121.410 127.440 121.580 128.285 ;
        RECT 122.030 128.115 122.250 128.985 ;
        RECT 122.475 128.865 123.170 129.055 ;
        RECT 121.750 127.735 122.250 128.115 ;
        RECT 122.420 128.065 122.830 128.685 ;
        RECT 123.000 127.895 123.170 128.865 ;
        RECT 122.475 127.725 123.170 127.895 ;
        RECT 120.790 127.055 121.170 127.435 ;
        RECT 121.410 127.270 122.240 127.440 ;
        RECT 122.475 127.225 122.645 127.725 ;
        RECT 122.815 127.055 123.145 127.555 ;
        RECT 123.360 127.225 123.585 129.345 ;
        RECT 123.755 129.225 124.085 129.605 ;
        RECT 124.255 129.055 124.425 129.345 ;
        RECT 123.760 128.885 124.425 129.055 ;
        RECT 123.760 127.895 123.990 128.885 ;
        RECT 124.685 128.835 126.355 129.605 ;
        RECT 126.525 128.855 127.735 129.605 ;
        RECT 124.160 128.065 124.510 128.715 ;
        RECT 124.685 128.145 125.435 128.665 ;
        RECT 125.605 128.315 126.355 128.835 ;
        RECT 126.525 128.145 127.045 128.685 ;
        RECT 127.215 128.315 127.735 128.855 ;
        RECT 123.760 127.725 124.425 127.895 ;
        RECT 123.755 127.055 124.085 127.555 ;
        RECT 124.255 127.225 124.425 127.725 ;
        RECT 124.685 127.055 126.355 128.145 ;
        RECT 126.525 127.055 127.735 128.145 ;
        RECT 29.840 126.885 127.820 127.055 ;
        RECT 29.925 125.795 31.135 126.885 ;
        RECT 29.925 125.085 30.445 125.625 ;
        RECT 30.615 125.255 31.135 125.795 ;
        RECT 31.305 125.795 33.895 126.885 ;
        RECT 34.375 126.045 34.545 126.885 ;
        RECT 34.755 125.875 35.005 126.715 ;
        RECT 35.215 126.045 35.385 126.885 ;
        RECT 35.555 125.875 35.845 126.715 ;
        RECT 31.305 125.275 32.515 125.795 ;
        RECT 34.120 125.705 35.845 125.875 ;
        RECT 36.055 125.825 36.225 126.885 ;
        RECT 36.520 126.505 36.850 126.885 ;
        RECT 37.030 126.335 37.200 126.625 ;
        RECT 37.370 126.425 37.620 126.885 ;
        RECT 36.400 126.165 37.200 126.335 ;
        RECT 37.790 126.375 38.660 126.715 ;
        RECT 32.685 125.105 33.895 125.625 ;
        RECT 29.925 124.335 31.135 125.085 ;
        RECT 31.305 124.335 33.895 125.105 ;
        RECT 34.120 125.155 34.530 125.705 ;
        RECT 36.400 125.545 36.570 126.165 ;
        RECT 37.790 125.995 37.960 126.375 ;
        RECT 38.895 126.255 39.065 126.715 ;
        RECT 39.235 126.425 39.605 126.885 ;
        RECT 39.900 126.285 40.070 126.625 ;
        RECT 40.240 126.455 40.570 126.885 ;
        RECT 40.805 126.285 40.975 126.625 ;
        RECT 36.740 125.825 37.960 125.995 ;
        RECT 38.130 125.915 38.590 126.205 ;
        RECT 38.895 126.085 39.455 126.255 ;
        RECT 39.900 126.115 40.975 126.285 ;
        RECT 41.145 126.385 41.825 126.715 ;
        RECT 42.040 126.385 42.290 126.715 ;
        RECT 42.460 126.425 42.710 126.885 ;
        RECT 39.285 125.945 39.455 126.085 ;
        RECT 38.130 125.905 39.095 125.915 ;
        RECT 37.790 125.735 37.960 125.825 ;
        RECT 38.420 125.745 39.095 125.905 ;
        RECT 36.400 125.535 36.745 125.545 ;
        RECT 34.715 125.325 36.745 125.535 ;
        RECT 34.120 124.985 35.885 125.155 ;
        RECT 34.375 124.335 34.545 124.805 ;
        RECT 34.715 124.505 35.045 124.985 ;
        RECT 35.215 124.335 35.385 124.805 ;
        RECT 35.555 124.505 35.885 124.985 ;
        RECT 36.055 124.335 36.225 125.145 ;
        RECT 36.420 125.070 36.745 125.325 ;
        RECT 36.425 124.715 36.745 125.070 ;
        RECT 36.915 125.285 37.455 125.655 ;
        RECT 37.790 125.565 38.195 125.735 ;
        RECT 36.915 124.885 37.155 125.285 ;
        RECT 37.635 125.115 37.855 125.395 ;
        RECT 37.325 124.945 37.855 125.115 ;
        RECT 37.325 124.715 37.495 124.945 ;
        RECT 38.025 124.785 38.195 125.565 ;
        RECT 38.365 124.955 38.715 125.575 ;
        RECT 38.885 124.955 39.095 125.745 ;
        RECT 39.285 125.775 40.785 125.945 ;
        RECT 39.285 125.085 39.455 125.775 ;
        RECT 41.145 125.605 41.315 126.385 ;
        RECT 42.120 126.255 42.290 126.385 ;
        RECT 39.625 125.435 41.315 125.605 ;
        RECT 41.485 125.825 41.950 126.215 ;
        RECT 42.120 126.085 42.515 126.255 ;
        RECT 39.625 125.255 39.795 125.435 ;
        RECT 36.425 124.545 37.495 124.715 ;
        RECT 37.665 124.335 37.855 124.775 ;
        RECT 38.025 124.505 38.975 124.785 ;
        RECT 39.285 124.695 39.545 125.085 ;
        RECT 39.965 125.015 40.755 125.265 ;
        RECT 39.195 124.525 39.545 124.695 ;
        RECT 39.755 124.335 40.085 124.795 ;
        RECT 40.960 124.725 41.130 125.435 ;
        RECT 41.485 125.235 41.655 125.825 ;
        RECT 41.300 125.015 41.655 125.235 ;
        RECT 41.825 125.015 42.175 125.635 ;
        RECT 42.345 124.725 42.515 126.085 ;
        RECT 42.880 125.915 43.205 126.700 ;
        RECT 42.685 124.865 43.145 125.915 ;
        RECT 40.960 124.555 41.815 124.725 ;
        RECT 42.020 124.555 42.515 124.725 ;
        RECT 42.685 124.335 43.015 124.695 ;
        RECT 43.375 124.595 43.545 126.715 ;
        RECT 43.715 126.385 44.045 126.885 ;
        RECT 44.215 126.215 44.470 126.715 ;
        RECT 43.720 126.045 44.470 126.215 ;
        RECT 43.720 125.055 43.950 126.045 ;
        RECT 44.120 125.225 44.470 125.875 ;
        RECT 45.110 125.745 45.445 126.715 ;
        RECT 45.615 125.745 45.785 126.885 ;
        RECT 45.955 126.545 47.985 126.715 ;
        RECT 45.110 125.075 45.280 125.745 ;
        RECT 45.955 125.575 46.125 126.545 ;
        RECT 45.450 125.245 45.705 125.575 ;
        RECT 45.930 125.245 46.125 125.575 ;
        RECT 46.295 126.205 47.420 126.375 ;
        RECT 45.535 125.075 45.705 125.245 ;
        RECT 46.295 125.075 46.465 126.205 ;
        RECT 43.720 124.885 44.470 125.055 ;
        RECT 43.715 124.335 44.045 124.715 ;
        RECT 44.215 124.595 44.470 124.885 ;
        RECT 45.110 124.505 45.365 125.075 ;
        RECT 45.535 124.905 46.465 125.075 ;
        RECT 46.635 125.865 47.645 126.035 ;
        RECT 46.635 125.065 46.805 125.865 ;
        RECT 47.010 125.525 47.285 125.665 ;
        RECT 47.005 125.355 47.285 125.525 ;
        RECT 46.290 124.870 46.465 124.905 ;
        RECT 45.535 124.335 45.865 124.735 ;
        RECT 46.290 124.505 46.820 124.870 ;
        RECT 47.010 124.505 47.285 125.355 ;
        RECT 47.455 124.505 47.645 125.865 ;
        RECT 47.815 125.880 47.985 126.545 ;
        RECT 48.155 126.125 48.325 126.885 ;
        RECT 48.560 126.125 49.075 126.535 ;
        RECT 47.815 125.690 48.565 125.880 ;
        RECT 48.735 125.315 49.075 126.125 ;
        RECT 50.165 125.720 50.455 126.885 ;
        RECT 51.235 125.735 51.565 126.885 ;
        RECT 51.735 125.865 51.905 126.715 ;
        RECT 52.075 126.085 52.405 126.885 ;
        RECT 52.575 125.865 52.745 126.715 ;
        RECT 52.925 126.085 53.165 126.885 ;
        RECT 53.335 125.905 53.665 126.715 ;
        RECT 54.505 126.215 54.785 126.885 ;
        RECT 54.955 125.995 55.255 126.545 ;
        RECT 55.455 126.165 55.785 126.885 ;
        RECT 55.975 126.165 56.435 126.715 ;
        RECT 56.805 126.215 57.085 126.885 ;
        RECT 47.845 125.145 49.075 125.315 ;
        RECT 51.735 125.695 52.745 125.865 ;
        RECT 52.950 125.735 53.665 125.905 ;
        RECT 51.735 125.185 52.230 125.695 ;
        RECT 52.950 125.495 53.120 125.735 ;
        RECT 54.320 125.575 54.585 125.935 ;
        RECT 54.955 125.825 55.895 125.995 ;
        RECT 55.725 125.575 55.895 125.825 ;
        RECT 52.620 125.325 53.120 125.495 ;
        RECT 53.290 125.325 53.670 125.565 ;
        RECT 54.320 125.325 54.995 125.575 ;
        RECT 55.215 125.325 55.555 125.575 ;
        RECT 51.735 125.155 52.235 125.185 ;
        RECT 52.950 125.155 53.120 125.325 ;
        RECT 55.725 125.245 56.015 125.575 ;
        RECT 55.725 125.155 55.895 125.245 ;
        RECT 47.825 124.335 48.335 124.870 ;
        RECT 48.555 124.540 48.800 125.145 ;
        RECT 50.165 124.335 50.455 125.060 ;
        RECT 51.235 124.335 51.565 125.135 ;
        RECT 51.735 124.985 52.745 125.155 ;
        RECT 52.950 124.985 53.585 125.155 ;
        RECT 51.735 124.505 51.905 124.985 ;
        RECT 52.075 124.335 52.405 124.815 ;
        RECT 52.575 124.505 52.745 124.985 ;
        RECT 52.995 124.335 53.235 124.815 ;
        RECT 53.415 124.505 53.585 124.985 ;
        RECT 54.505 124.965 55.895 125.155 ;
        RECT 54.505 124.605 54.835 124.965 ;
        RECT 56.185 124.795 56.435 126.165 ;
        RECT 57.255 125.995 57.555 126.545 ;
        RECT 57.755 126.165 58.085 126.885 ;
        RECT 58.275 126.165 58.735 126.715 ;
        RECT 59.280 126.545 59.535 126.575 ;
        RECT 59.195 126.375 59.535 126.545 ;
        RECT 56.620 125.575 56.885 125.935 ;
        RECT 57.255 125.825 58.195 125.995 ;
        RECT 58.025 125.575 58.195 125.825 ;
        RECT 56.620 125.325 57.295 125.575 ;
        RECT 57.515 125.325 57.855 125.575 ;
        RECT 58.025 125.245 58.315 125.575 ;
        RECT 58.025 125.155 58.195 125.245 ;
        RECT 55.455 124.335 55.705 124.795 ;
        RECT 55.875 124.505 56.435 124.795 ;
        RECT 56.805 124.965 58.195 125.155 ;
        RECT 56.805 124.605 57.135 124.965 ;
        RECT 58.485 124.795 58.735 126.165 ;
        RECT 57.755 124.335 58.005 124.795 ;
        RECT 58.175 124.505 58.735 124.795 ;
        RECT 59.280 125.905 59.535 126.375 ;
        RECT 59.715 126.085 60.000 126.885 ;
        RECT 60.180 126.165 60.510 126.675 ;
        RECT 59.280 125.045 59.460 125.905 ;
        RECT 60.180 125.575 60.430 126.165 ;
        RECT 60.780 126.015 60.950 126.625 ;
        RECT 61.120 126.195 61.450 126.885 ;
        RECT 61.680 126.335 61.920 126.625 ;
        RECT 62.120 126.505 62.540 126.885 ;
        RECT 62.720 126.415 63.350 126.665 ;
        RECT 63.820 126.505 64.150 126.885 ;
        RECT 62.720 126.335 62.890 126.415 ;
        RECT 64.320 126.335 64.490 126.625 ;
        RECT 64.670 126.505 65.050 126.885 ;
        RECT 65.290 126.500 66.120 126.670 ;
        RECT 61.680 126.165 62.890 126.335 ;
        RECT 59.630 125.245 60.430 125.575 ;
        RECT 59.280 124.515 59.535 125.045 ;
        RECT 59.715 124.335 60.000 124.795 ;
        RECT 60.180 124.595 60.430 125.245 ;
        RECT 60.630 125.995 60.950 126.015 ;
        RECT 60.630 125.825 62.550 125.995 ;
        RECT 60.630 124.930 60.820 125.825 ;
        RECT 62.720 125.655 62.890 126.165 ;
        RECT 63.060 125.905 63.580 126.215 ;
        RECT 60.990 125.485 62.890 125.655 ;
        RECT 60.990 125.425 61.320 125.485 ;
        RECT 61.470 125.255 61.800 125.315 ;
        RECT 61.140 124.985 61.800 125.255 ;
        RECT 60.630 124.600 60.950 124.930 ;
        RECT 61.130 124.335 61.790 124.815 ;
        RECT 61.990 124.725 62.160 125.485 ;
        RECT 63.060 125.315 63.240 125.725 ;
        RECT 62.330 125.145 62.660 125.265 ;
        RECT 63.410 125.145 63.580 125.905 ;
        RECT 62.330 124.975 63.580 125.145 ;
        RECT 63.750 126.085 65.120 126.335 ;
        RECT 63.750 125.315 63.940 126.085 ;
        RECT 64.870 125.825 65.120 126.085 ;
        RECT 64.110 125.655 64.360 125.815 ;
        RECT 65.290 125.655 65.460 126.500 ;
        RECT 66.355 126.215 66.525 126.715 ;
        RECT 66.695 126.385 67.025 126.885 ;
        RECT 65.630 125.825 66.130 126.205 ;
        RECT 66.355 126.045 67.050 126.215 ;
        RECT 64.110 125.485 65.460 125.655 ;
        RECT 65.040 125.445 65.460 125.485 ;
        RECT 63.750 124.975 64.170 125.315 ;
        RECT 64.460 124.985 64.870 125.315 ;
        RECT 61.990 124.555 62.840 124.725 ;
        RECT 63.400 124.335 63.720 124.795 ;
        RECT 63.920 124.545 64.170 124.975 ;
        RECT 64.460 124.335 64.870 124.775 ;
        RECT 65.040 124.715 65.210 125.445 ;
        RECT 65.380 124.895 65.730 125.265 ;
        RECT 65.910 124.955 66.130 125.825 ;
        RECT 66.300 125.255 66.710 125.875 ;
        RECT 66.880 125.075 67.050 126.045 ;
        RECT 66.355 124.885 67.050 125.075 ;
        RECT 65.040 124.515 66.055 124.715 ;
        RECT 66.355 124.555 66.525 124.885 ;
        RECT 66.695 124.335 67.025 124.715 ;
        RECT 67.240 124.595 67.465 126.715 ;
        RECT 67.635 126.385 67.965 126.885 ;
        RECT 68.135 126.215 68.305 126.715 ;
        RECT 67.640 126.045 68.305 126.215 ;
        RECT 67.640 125.055 67.870 126.045 ;
        RECT 68.040 125.225 68.390 125.875 ;
        RECT 68.565 125.795 69.775 126.885 ;
        RECT 69.945 125.795 73.455 126.885 ;
        RECT 73.715 125.955 73.885 126.715 ;
        RECT 74.065 126.125 74.395 126.885 ;
        RECT 68.565 125.255 69.085 125.795 ;
        RECT 69.255 125.085 69.775 125.625 ;
        RECT 69.945 125.275 71.635 125.795 ;
        RECT 73.715 125.785 74.380 125.955 ;
        RECT 74.565 125.810 74.835 126.715 ;
        RECT 74.210 125.640 74.380 125.785 ;
        RECT 71.805 125.105 73.455 125.625 ;
        RECT 73.645 125.235 73.975 125.605 ;
        RECT 74.210 125.310 74.495 125.640 ;
        RECT 67.640 124.885 68.305 125.055 ;
        RECT 67.635 124.335 67.965 124.715 ;
        RECT 68.135 124.595 68.305 124.885 ;
        RECT 68.565 124.335 69.775 125.085 ;
        RECT 69.945 124.335 73.455 125.105 ;
        RECT 74.210 125.055 74.380 125.310 ;
        RECT 73.715 124.885 74.380 125.055 ;
        RECT 74.665 125.010 74.835 125.810 ;
        RECT 75.925 125.720 76.215 126.885 ;
        RECT 76.390 126.450 81.735 126.885 ;
        RECT 81.910 126.450 87.255 126.885 ;
        RECT 77.980 125.200 78.330 126.450 ;
        RECT 73.715 124.505 73.885 124.885 ;
        RECT 74.065 124.335 74.395 124.715 ;
        RECT 74.575 124.505 74.835 125.010 ;
        RECT 75.925 124.335 76.215 125.060 ;
        RECT 79.810 124.880 80.150 125.710 ;
        RECT 83.500 125.200 83.850 126.450 ;
        RECT 87.515 125.955 87.685 126.715 ;
        RECT 87.865 126.125 88.195 126.885 ;
        RECT 87.515 125.785 88.180 125.955 ;
        RECT 88.365 125.810 88.635 126.715 ;
        RECT 85.330 124.880 85.670 125.710 ;
        RECT 88.010 125.640 88.180 125.785 ;
        RECT 87.445 125.235 87.775 125.605 ;
        RECT 88.010 125.310 88.295 125.640 ;
        RECT 88.010 125.055 88.180 125.310 ;
        RECT 87.515 124.885 88.180 125.055 ;
        RECT 88.465 125.010 88.635 125.810 ;
        RECT 88.805 125.795 90.015 126.885 ;
        RECT 90.190 126.450 95.535 126.885 ;
        RECT 88.805 125.255 89.325 125.795 ;
        RECT 89.495 125.085 90.015 125.625 ;
        RECT 91.780 125.200 92.130 126.450 ;
        RECT 95.765 125.745 95.975 126.885 ;
        RECT 96.145 125.735 96.475 126.715 ;
        RECT 96.645 125.745 96.875 126.885 ;
        RECT 98.005 125.795 101.515 126.885 ;
        RECT 76.390 124.335 81.735 124.880 ;
        RECT 81.910 124.335 87.255 124.880 ;
        RECT 87.515 124.505 87.685 124.885 ;
        RECT 87.865 124.335 88.195 124.715 ;
        RECT 88.375 124.505 88.635 125.010 ;
        RECT 88.805 124.335 90.015 125.085 ;
        RECT 93.610 124.880 93.950 125.710 ;
        RECT 90.190 124.335 95.535 124.880 ;
        RECT 95.765 124.335 95.975 125.155 ;
        RECT 96.145 125.135 96.395 125.735 ;
        RECT 96.565 125.325 96.895 125.575 ;
        RECT 98.005 125.275 99.695 125.795 ;
        RECT 101.685 125.720 101.975 126.885 ;
        RECT 103.070 126.450 108.415 126.885 ;
        RECT 96.145 124.505 96.475 125.135 ;
        RECT 96.645 124.335 96.875 125.155 ;
        RECT 99.865 125.105 101.515 125.625 ;
        RECT 104.660 125.200 105.010 126.450 ;
        RECT 108.645 125.745 108.855 126.885 ;
        RECT 109.025 125.735 109.355 126.715 ;
        RECT 109.525 125.745 109.755 126.885 ;
        RECT 110.885 125.795 114.395 126.885 ;
        RECT 114.570 126.450 119.915 126.885 ;
        RECT 98.005 124.335 101.515 125.105 ;
        RECT 101.685 124.335 101.975 125.060 ;
        RECT 106.490 124.880 106.830 125.710 ;
        RECT 103.070 124.335 108.415 124.880 ;
        RECT 108.645 124.335 108.855 125.155 ;
        RECT 109.025 125.135 109.275 125.735 ;
        RECT 109.445 125.325 109.775 125.575 ;
        RECT 110.885 125.275 112.575 125.795 ;
        RECT 109.025 124.505 109.355 125.135 ;
        RECT 109.525 124.335 109.755 125.155 ;
        RECT 112.745 125.105 114.395 125.625 ;
        RECT 116.160 125.200 116.510 126.450 ;
        RECT 120.125 125.745 120.355 126.885 ;
        RECT 120.525 125.735 120.855 126.715 ;
        RECT 121.025 125.745 121.235 126.885 ;
        RECT 121.555 125.955 121.725 126.715 ;
        RECT 121.905 126.125 122.235 126.885 ;
        RECT 121.555 125.785 122.220 125.955 ;
        RECT 122.405 125.810 122.675 126.715 ;
        RECT 110.885 124.335 114.395 125.105 ;
        RECT 117.990 124.880 118.330 125.710 ;
        RECT 120.105 125.325 120.435 125.575 ;
        RECT 114.570 124.335 119.915 124.880 ;
        RECT 120.125 124.335 120.355 125.155 ;
        RECT 120.605 125.135 120.855 125.735 ;
        RECT 122.050 125.640 122.220 125.785 ;
        RECT 121.485 125.235 121.815 125.605 ;
        RECT 122.050 125.310 122.335 125.640 ;
        RECT 120.525 124.505 120.855 125.135 ;
        RECT 121.025 124.335 121.235 125.155 ;
        RECT 122.050 125.055 122.220 125.310 ;
        RECT 121.555 124.885 122.220 125.055 ;
        RECT 122.505 125.010 122.675 125.810 ;
        RECT 121.555 124.505 121.725 124.885 ;
        RECT 121.905 124.335 122.235 124.715 ;
        RECT 122.415 124.505 122.675 125.010 ;
        RECT 122.845 125.810 123.115 126.715 ;
        RECT 123.285 126.125 123.615 126.885 ;
        RECT 123.795 125.955 123.965 126.715 ;
        RECT 122.845 125.010 123.015 125.810 ;
        RECT 123.300 125.785 123.965 125.955 ;
        RECT 124.685 125.795 126.355 126.885 ;
        RECT 126.525 125.795 127.735 126.885 ;
        RECT 123.300 125.640 123.470 125.785 ;
        RECT 123.185 125.310 123.470 125.640 ;
        RECT 123.300 125.055 123.470 125.310 ;
        RECT 123.705 125.235 124.035 125.605 ;
        RECT 124.685 125.275 125.435 125.795 ;
        RECT 125.605 125.105 126.355 125.625 ;
        RECT 126.525 125.255 127.045 125.795 ;
        RECT 122.845 124.505 123.105 125.010 ;
        RECT 123.300 124.885 123.965 125.055 ;
        RECT 123.285 124.335 123.615 124.715 ;
        RECT 123.795 124.505 123.965 124.885 ;
        RECT 124.685 124.335 126.355 125.105 ;
        RECT 127.215 125.085 127.735 125.625 ;
        RECT 126.525 124.335 127.735 125.085 ;
        RECT 29.840 124.165 127.820 124.335 ;
        RECT 29.925 123.415 31.135 124.165 ;
        RECT 31.770 123.620 37.115 124.165 ;
        RECT 29.925 122.875 30.445 123.415 ;
        RECT 30.615 122.705 31.135 123.245 ;
        RECT 29.925 121.615 31.135 122.705 ;
        RECT 33.360 122.050 33.710 123.300 ;
        RECT 35.190 122.790 35.530 123.620 ;
        RECT 37.285 123.440 37.575 124.165 ;
        RECT 38.055 123.695 38.225 124.165 ;
        RECT 38.395 123.515 38.725 123.995 ;
        RECT 38.895 123.695 39.065 124.165 ;
        RECT 39.235 123.515 39.565 123.995 ;
        RECT 37.800 123.345 39.565 123.515 ;
        RECT 39.735 123.355 39.905 124.165 ;
        RECT 40.105 123.785 41.175 123.955 ;
        RECT 40.105 123.430 40.425 123.785 ;
        RECT 37.800 122.795 38.210 123.345 ;
        RECT 40.100 123.175 40.425 123.430 ;
        RECT 38.395 122.965 40.425 123.175 ;
        RECT 40.080 122.955 40.425 122.965 ;
        RECT 40.595 123.215 40.835 123.615 ;
        RECT 41.005 123.555 41.175 123.785 ;
        RECT 41.345 123.725 41.535 124.165 ;
        RECT 41.705 123.715 42.655 123.995 ;
        RECT 42.875 123.805 43.225 123.975 ;
        RECT 41.005 123.385 41.535 123.555 ;
        RECT 31.770 121.615 37.115 122.050 ;
        RECT 37.285 121.615 37.575 122.780 ;
        RECT 37.800 122.625 39.525 122.795 ;
        RECT 38.055 121.615 38.225 122.455 ;
        RECT 38.435 121.785 38.685 122.625 ;
        RECT 38.895 121.615 39.065 122.455 ;
        RECT 39.235 121.785 39.525 122.625 ;
        RECT 39.735 121.615 39.905 122.675 ;
        RECT 40.080 122.335 40.250 122.955 ;
        RECT 40.595 122.845 41.135 123.215 ;
        RECT 41.315 123.105 41.535 123.385 ;
        RECT 41.705 122.935 41.875 123.715 ;
        RECT 41.470 122.765 41.875 122.935 ;
        RECT 42.045 122.925 42.395 123.545 ;
        RECT 41.470 122.675 41.640 122.765 ;
        RECT 42.565 122.755 42.775 123.545 ;
        RECT 40.420 122.505 41.640 122.675 ;
        RECT 42.100 122.595 42.775 122.755 ;
        RECT 40.080 122.165 40.880 122.335 ;
        RECT 40.200 121.615 40.530 121.995 ;
        RECT 40.710 121.875 40.880 122.165 ;
        RECT 41.470 122.125 41.640 122.505 ;
        RECT 41.810 122.585 42.775 122.595 ;
        RECT 42.965 123.415 43.225 123.805 ;
        RECT 43.435 123.705 43.765 124.165 ;
        RECT 44.640 123.775 45.495 123.945 ;
        RECT 45.700 123.775 46.195 123.945 ;
        RECT 46.365 123.805 46.695 124.165 ;
        RECT 42.965 122.725 43.135 123.415 ;
        RECT 43.305 123.065 43.475 123.245 ;
        RECT 43.645 123.235 44.435 123.485 ;
        RECT 44.640 123.065 44.810 123.775 ;
        RECT 44.980 123.265 45.335 123.485 ;
        RECT 43.305 122.895 44.995 123.065 ;
        RECT 41.810 122.295 42.270 122.585 ;
        RECT 42.965 122.555 44.465 122.725 ;
        RECT 42.965 122.415 43.135 122.555 ;
        RECT 42.575 122.245 43.135 122.415 ;
        RECT 41.050 121.615 41.300 122.075 ;
        RECT 41.470 121.785 42.340 122.125 ;
        RECT 42.575 121.785 42.745 122.245 ;
        RECT 43.580 122.215 44.655 122.385 ;
        RECT 42.915 121.615 43.285 122.075 ;
        RECT 43.580 121.875 43.750 122.215 ;
        RECT 43.920 121.615 44.250 122.045 ;
        RECT 44.485 121.875 44.655 122.215 ;
        RECT 44.825 122.115 44.995 122.895 ;
        RECT 45.165 122.675 45.335 123.265 ;
        RECT 45.505 122.865 45.855 123.485 ;
        RECT 45.165 122.285 45.630 122.675 ;
        RECT 46.025 122.415 46.195 123.775 ;
        RECT 46.365 122.585 46.825 123.635 ;
        RECT 45.800 122.245 46.195 122.415 ;
        RECT 45.800 122.115 45.970 122.245 ;
        RECT 44.825 121.785 45.505 122.115 ;
        RECT 45.720 121.785 45.970 122.115 ;
        RECT 46.140 121.615 46.390 122.075 ;
        RECT 46.560 121.800 46.885 122.585 ;
        RECT 47.055 121.785 47.225 123.905 ;
        RECT 47.395 123.785 47.725 124.165 ;
        RECT 47.895 123.615 48.150 123.905 ;
        RECT 47.400 123.445 48.150 123.615 ;
        RECT 48.325 123.490 48.585 123.995 ;
        RECT 48.765 123.785 49.095 124.165 ;
        RECT 49.275 123.615 49.445 123.995 ;
        RECT 47.400 122.455 47.630 123.445 ;
        RECT 47.800 122.625 48.150 123.275 ;
        RECT 48.325 122.690 48.495 123.490 ;
        RECT 48.780 123.445 49.445 123.615 ;
        RECT 48.780 123.190 48.950 123.445 ;
        RECT 50.165 123.395 51.835 124.165 ;
        RECT 52.010 123.620 57.355 124.165 ;
        RECT 48.665 122.860 48.950 123.190 ;
        RECT 49.185 122.895 49.515 123.265 ;
        RECT 48.780 122.715 48.950 122.860 ;
        RECT 47.400 122.285 48.150 122.455 ;
        RECT 47.395 121.615 47.725 122.115 ;
        RECT 47.895 121.785 48.150 122.285 ;
        RECT 48.325 121.785 48.595 122.690 ;
        RECT 48.780 122.545 49.445 122.715 ;
        RECT 48.765 121.615 49.095 122.375 ;
        RECT 49.275 121.785 49.445 122.545 ;
        RECT 50.165 122.705 50.915 123.225 ;
        RECT 51.085 122.875 51.835 123.395 ;
        RECT 50.165 121.615 51.835 122.705 ;
        RECT 53.600 122.050 53.950 123.300 ;
        RECT 55.430 122.790 55.770 123.620 ;
        RECT 57.585 123.345 57.795 124.165 ;
        RECT 57.965 123.365 58.295 123.995 ;
        RECT 57.965 122.765 58.215 123.365 ;
        RECT 58.465 123.345 58.695 124.165 ;
        RECT 59.365 123.395 62.875 124.165 ;
        RECT 63.045 123.440 63.335 124.165 ;
        RECT 64.515 123.615 64.685 123.995 ;
        RECT 64.865 123.785 65.195 124.165 ;
        RECT 64.515 123.445 65.180 123.615 ;
        RECT 65.375 123.490 65.635 123.995 ;
        RECT 58.385 122.925 58.715 123.175 ;
        RECT 52.010 121.615 57.355 122.050 ;
        RECT 57.585 121.615 57.795 122.755 ;
        RECT 57.965 121.785 58.295 122.765 ;
        RECT 58.465 121.615 58.695 122.755 ;
        RECT 59.365 122.705 61.055 123.225 ;
        RECT 61.225 122.875 62.875 123.395 ;
        RECT 64.445 122.895 64.775 123.265 ;
        RECT 65.010 123.190 65.180 123.445 ;
        RECT 65.010 122.860 65.295 123.190 ;
        RECT 59.365 121.615 62.875 122.705 ;
        RECT 63.045 121.615 63.335 122.780 ;
        RECT 65.010 122.715 65.180 122.860 ;
        RECT 64.515 122.545 65.180 122.715 ;
        RECT 65.465 122.690 65.635 123.490 ;
        RECT 65.805 123.415 67.015 124.165 ;
        RECT 64.515 121.785 64.685 122.545 ;
        RECT 64.865 121.615 65.195 122.375 ;
        RECT 65.365 121.785 65.635 122.690 ;
        RECT 65.805 122.705 66.325 123.245 ;
        RECT 66.495 122.875 67.015 123.415 ;
        RECT 67.185 123.395 70.695 124.165 ;
        RECT 67.185 122.705 68.875 123.225 ;
        RECT 69.045 122.875 70.695 123.395 ;
        RECT 70.955 123.515 71.125 123.995 ;
        RECT 71.305 123.685 71.545 124.165 ;
        RECT 71.795 123.515 71.965 123.995 ;
        RECT 72.135 123.685 72.465 124.165 ;
        RECT 72.635 123.515 72.805 123.995 ;
        RECT 70.955 123.345 71.590 123.515 ;
        RECT 71.795 123.345 72.805 123.515 ;
        RECT 72.975 123.365 73.305 124.165 ;
        RECT 73.625 123.415 74.835 124.165 ;
        RECT 71.420 123.175 71.590 123.345 ;
        RECT 70.870 122.935 71.250 123.175 ;
        RECT 71.420 123.005 71.920 123.175 ;
        RECT 72.310 123.145 72.805 123.345 ;
        RECT 71.420 122.765 71.590 123.005 ;
        RECT 72.305 122.975 72.805 123.145 ;
        RECT 72.310 122.805 72.805 122.975 ;
        RECT 65.805 121.615 67.015 122.705 ;
        RECT 67.185 121.615 70.695 122.705 ;
        RECT 70.875 122.595 71.590 122.765 ;
        RECT 71.795 122.635 72.805 122.805 ;
        RECT 70.875 121.785 71.205 122.595 ;
        RECT 71.375 121.615 71.615 122.415 ;
        RECT 71.795 121.785 71.965 122.635 ;
        RECT 72.135 121.615 72.465 122.415 ;
        RECT 72.635 121.785 72.805 122.635 ;
        RECT 72.975 121.615 73.305 122.765 ;
        RECT 73.625 122.705 74.145 123.245 ;
        RECT 74.315 122.875 74.835 123.415 ;
        RECT 75.005 123.395 78.515 124.165 ;
        RECT 78.690 123.620 84.035 124.165 ;
        RECT 75.005 122.705 76.695 123.225 ;
        RECT 76.865 122.875 78.515 123.395 ;
        RECT 73.625 121.615 74.835 122.705 ;
        RECT 75.005 121.615 78.515 122.705 ;
        RECT 80.280 122.050 80.630 123.300 ;
        RECT 82.110 122.790 82.450 123.620 ;
        RECT 84.265 123.345 84.475 124.165 ;
        RECT 84.645 123.365 84.975 123.995 ;
        RECT 84.645 122.765 84.895 123.365 ;
        RECT 85.145 123.345 85.375 124.165 ;
        RECT 86.135 123.515 86.305 123.995 ;
        RECT 86.485 123.685 86.725 124.165 ;
        RECT 86.975 123.515 87.145 123.995 ;
        RECT 87.315 123.685 87.645 124.165 ;
        RECT 87.815 123.515 87.985 123.995 ;
        RECT 86.135 123.345 86.770 123.515 ;
        RECT 86.975 123.345 87.985 123.515 ;
        RECT 88.155 123.365 88.485 124.165 ;
        RECT 88.805 123.440 89.095 124.165 ;
        RECT 89.725 123.395 93.235 124.165 ;
        RECT 86.600 123.175 86.770 123.345 ;
        RECT 85.065 122.925 85.395 123.175 ;
        RECT 86.050 122.935 86.430 123.175 ;
        RECT 86.600 123.005 87.100 123.175 ;
        RECT 87.490 123.145 87.985 123.345 ;
        RECT 86.600 122.765 86.770 123.005 ;
        RECT 87.485 122.975 87.985 123.145 ;
        RECT 87.490 122.805 87.985 122.975 ;
        RECT 78.690 121.615 84.035 122.050 ;
        RECT 84.265 121.615 84.475 122.755 ;
        RECT 84.645 121.785 84.975 122.765 ;
        RECT 85.145 121.615 85.375 122.755 ;
        RECT 86.055 122.595 86.770 122.765 ;
        RECT 86.975 122.635 87.985 122.805 ;
        RECT 86.055 121.785 86.385 122.595 ;
        RECT 86.555 121.615 86.795 122.415 ;
        RECT 86.975 121.785 87.145 122.635 ;
        RECT 87.315 121.615 87.645 122.415 ;
        RECT 87.815 121.785 87.985 122.635 ;
        RECT 88.155 121.615 88.485 122.765 ;
        RECT 88.805 121.615 89.095 122.780 ;
        RECT 89.725 122.705 91.415 123.225 ;
        RECT 91.585 122.875 93.235 123.395 ;
        RECT 93.465 123.345 93.675 124.165 ;
        RECT 93.845 123.365 94.175 123.995 ;
        RECT 93.845 122.765 94.095 123.365 ;
        RECT 94.345 123.345 94.575 124.165 ;
        RECT 94.875 123.615 95.045 123.995 ;
        RECT 95.225 123.785 95.555 124.165 ;
        RECT 94.875 123.445 95.540 123.615 ;
        RECT 95.735 123.490 95.995 123.995 ;
        RECT 94.265 122.925 94.595 123.175 ;
        RECT 94.805 122.895 95.135 123.265 ;
        RECT 95.370 123.190 95.540 123.445 ;
        RECT 95.370 122.860 95.655 123.190 ;
        RECT 89.725 121.615 93.235 122.705 ;
        RECT 93.465 121.615 93.675 122.755 ;
        RECT 93.845 121.785 94.175 122.765 ;
        RECT 94.345 121.615 94.575 122.755 ;
        RECT 95.370 122.715 95.540 122.860 ;
        RECT 94.875 122.545 95.540 122.715 ;
        RECT 95.825 122.690 95.995 123.490 ;
        RECT 96.165 123.395 98.755 124.165 ;
        RECT 99.015 123.615 99.185 123.995 ;
        RECT 99.365 123.785 99.695 124.165 ;
        RECT 99.015 123.445 99.680 123.615 ;
        RECT 99.875 123.490 100.135 123.995 ;
        RECT 94.875 121.785 95.045 122.545 ;
        RECT 95.225 121.615 95.555 122.375 ;
        RECT 95.725 121.785 95.995 122.690 ;
        RECT 96.165 122.705 97.375 123.225 ;
        RECT 97.545 122.875 98.755 123.395 ;
        RECT 98.945 122.895 99.275 123.265 ;
        RECT 99.510 123.190 99.680 123.445 ;
        RECT 99.510 122.860 99.795 123.190 ;
        RECT 99.510 122.715 99.680 122.860 ;
        RECT 96.165 121.615 98.755 122.705 ;
        RECT 99.015 122.545 99.680 122.715 ;
        RECT 99.965 122.690 100.135 123.490 ;
        RECT 100.305 123.395 102.895 124.165 ;
        RECT 103.155 123.615 103.325 123.995 ;
        RECT 103.505 123.785 103.835 124.165 ;
        RECT 103.155 123.445 103.820 123.615 ;
        RECT 104.015 123.490 104.275 123.995 ;
        RECT 99.015 121.785 99.185 122.545 ;
        RECT 99.365 121.615 99.695 122.375 ;
        RECT 99.865 121.785 100.135 122.690 ;
        RECT 100.305 122.705 101.515 123.225 ;
        RECT 101.685 122.875 102.895 123.395 ;
        RECT 103.085 122.895 103.415 123.265 ;
        RECT 103.650 123.190 103.820 123.445 ;
        RECT 103.650 122.860 103.935 123.190 ;
        RECT 103.650 122.715 103.820 122.860 ;
        RECT 100.305 121.615 102.895 122.705 ;
        RECT 103.155 122.545 103.820 122.715 ;
        RECT 104.105 122.690 104.275 123.490 ;
        RECT 104.905 123.395 108.415 124.165 ;
        RECT 108.675 123.615 108.845 123.995 ;
        RECT 109.025 123.785 109.355 124.165 ;
        RECT 108.675 123.445 109.340 123.615 ;
        RECT 109.535 123.490 109.795 123.995 ;
        RECT 103.155 121.785 103.325 122.545 ;
        RECT 103.505 121.615 103.835 122.375 ;
        RECT 104.005 121.785 104.275 122.690 ;
        RECT 104.905 122.705 106.595 123.225 ;
        RECT 106.765 122.875 108.415 123.395 ;
        RECT 108.605 122.895 108.935 123.265 ;
        RECT 109.170 123.190 109.340 123.445 ;
        RECT 109.170 122.860 109.455 123.190 ;
        RECT 109.170 122.715 109.340 122.860 ;
        RECT 104.905 121.615 108.415 122.705 ;
        RECT 108.675 122.545 109.340 122.715 ;
        RECT 109.625 122.690 109.795 123.490 ;
        RECT 110.425 123.395 112.095 124.165 ;
        RECT 112.355 123.615 112.525 123.995 ;
        RECT 112.705 123.785 113.035 124.165 ;
        RECT 112.355 123.445 113.020 123.615 ;
        RECT 113.215 123.490 113.475 123.995 ;
        RECT 108.675 121.785 108.845 122.545 ;
        RECT 109.025 121.615 109.355 122.375 ;
        RECT 109.525 121.785 109.795 122.690 ;
        RECT 110.425 122.705 111.175 123.225 ;
        RECT 111.345 122.875 112.095 123.395 ;
        RECT 112.285 122.895 112.615 123.265 ;
        RECT 112.850 123.190 113.020 123.445 ;
        RECT 112.850 122.860 113.135 123.190 ;
        RECT 112.850 122.715 113.020 122.860 ;
        RECT 110.425 121.615 112.095 122.705 ;
        RECT 112.355 122.545 113.020 122.715 ;
        RECT 113.305 122.690 113.475 123.490 ;
        RECT 114.565 123.440 114.855 124.165 ;
        RECT 115.950 123.615 116.205 123.905 ;
        RECT 116.375 123.785 116.705 124.165 ;
        RECT 115.950 123.445 116.700 123.615 ;
        RECT 112.355 121.785 112.525 122.545 ;
        RECT 112.705 121.615 113.035 122.375 ;
        RECT 113.205 121.785 113.475 122.690 ;
        RECT 114.565 121.615 114.855 122.780 ;
        RECT 115.950 122.625 116.300 123.275 ;
        RECT 116.470 122.455 116.700 123.445 ;
        RECT 115.950 122.285 116.700 122.455 ;
        RECT 115.950 121.785 116.205 122.285 ;
        RECT 116.375 121.615 116.705 122.115 ;
        RECT 116.875 121.785 117.045 123.905 ;
        RECT 117.405 123.805 117.735 124.165 ;
        RECT 117.905 123.775 118.400 123.945 ;
        RECT 118.605 123.775 119.460 123.945 ;
        RECT 117.275 122.585 117.735 123.635 ;
        RECT 117.215 121.800 117.540 122.585 ;
        RECT 117.905 122.415 118.075 123.775 ;
        RECT 118.245 122.865 118.595 123.485 ;
        RECT 118.765 123.265 119.120 123.485 ;
        RECT 118.765 122.675 118.935 123.265 ;
        RECT 119.290 123.065 119.460 123.775 ;
        RECT 120.335 123.705 120.665 124.165 ;
        RECT 120.875 123.805 121.225 123.975 ;
        RECT 119.665 123.235 120.455 123.485 ;
        RECT 120.875 123.415 121.135 123.805 ;
        RECT 121.445 123.715 122.395 123.995 ;
        RECT 122.565 123.725 122.755 124.165 ;
        RECT 122.925 123.785 123.995 123.955 ;
        RECT 120.625 123.065 120.795 123.245 ;
        RECT 117.905 122.245 118.300 122.415 ;
        RECT 118.470 122.285 118.935 122.675 ;
        RECT 119.105 122.895 120.795 123.065 ;
        RECT 118.130 122.115 118.300 122.245 ;
        RECT 119.105 122.115 119.275 122.895 ;
        RECT 120.965 122.725 121.135 123.415 ;
        RECT 119.635 122.555 121.135 122.725 ;
        RECT 121.325 122.755 121.535 123.545 ;
        RECT 121.705 122.925 122.055 123.545 ;
        RECT 122.225 122.935 122.395 123.715 ;
        RECT 122.925 123.555 123.095 123.785 ;
        RECT 122.565 123.385 123.095 123.555 ;
        RECT 122.565 123.105 122.785 123.385 ;
        RECT 123.265 123.215 123.505 123.615 ;
        RECT 122.225 122.765 122.630 122.935 ;
        RECT 122.965 122.845 123.505 123.215 ;
        RECT 123.675 123.430 123.995 123.785 ;
        RECT 123.675 123.175 124.000 123.430 ;
        RECT 124.195 123.355 124.365 124.165 ;
        RECT 124.535 123.515 124.865 123.995 ;
        RECT 125.035 123.695 125.205 124.165 ;
        RECT 125.375 123.515 125.705 123.995 ;
        RECT 125.875 123.695 126.045 124.165 ;
        RECT 124.535 123.345 126.300 123.515 ;
        RECT 126.525 123.415 127.735 124.165 ;
        RECT 123.675 122.965 125.705 123.175 ;
        RECT 123.675 122.955 124.020 122.965 ;
        RECT 121.325 122.595 122.000 122.755 ;
        RECT 122.460 122.675 122.630 122.765 ;
        RECT 121.325 122.585 122.290 122.595 ;
        RECT 120.965 122.415 121.135 122.555 ;
        RECT 117.710 121.615 117.960 122.075 ;
        RECT 118.130 121.785 118.380 122.115 ;
        RECT 118.595 121.785 119.275 122.115 ;
        RECT 119.445 122.215 120.520 122.385 ;
        RECT 120.965 122.245 121.525 122.415 ;
        RECT 121.830 122.295 122.290 122.585 ;
        RECT 122.460 122.505 123.680 122.675 ;
        RECT 119.445 121.875 119.615 122.215 ;
        RECT 119.850 121.615 120.180 122.045 ;
        RECT 120.350 121.875 120.520 122.215 ;
        RECT 120.815 121.615 121.185 122.075 ;
        RECT 121.355 121.785 121.525 122.245 ;
        RECT 122.460 122.125 122.630 122.505 ;
        RECT 123.850 122.335 124.020 122.955 ;
        RECT 125.890 122.795 126.300 123.345 ;
        RECT 121.760 121.785 122.630 122.125 ;
        RECT 123.220 122.165 124.020 122.335 ;
        RECT 122.800 121.615 123.050 122.075 ;
        RECT 123.220 121.875 123.390 122.165 ;
        RECT 123.570 121.615 123.900 121.995 ;
        RECT 124.195 121.615 124.365 122.675 ;
        RECT 124.575 122.625 126.300 122.795 ;
        RECT 126.525 122.705 127.045 123.245 ;
        RECT 127.215 122.875 127.735 123.415 ;
        RECT 124.575 121.785 124.865 122.625 ;
        RECT 125.035 121.615 125.205 122.455 ;
        RECT 125.415 121.785 125.665 122.625 ;
        RECT 125.875 121.615 126.045 122.455 ;
        RECT 126.525 121.615 127.735 122.705 ;
        RECT 29.840 121.445 127.820 121.615 ;
        RECT 29.925 120.355 31.135 121.445 ;
        RECT 31.310 121.010 36.655 121.445 ;
        RECT 29.925 119.645 30.445 120.185 ;
        RECT 30.615 119.815 31.135 120.355 ;
        RECT 32.900 119.760 33.250 121.010 ;
        RECT 36.915 120.515 37.085 121.275 ;
        RECT 37.265 120.685 37.595 121.445 ;
        RECT 36.915 120.345 37.580 120.515 ;
        RECT 37.765 120.370 38.035 121.275 ;
        RECT 29.925 118.895 31.135 119.645 ;
        RECT 34.730 119.440 35.070 120.270 ;
        RECT 37.410 120.200 37.580 120.345 ;
        RECT 36.845 119.795 37.175 120.165 ;
        RECT 37.410 119.870 37.695 120.200 ;
        RECT 37.410 119.615 37.580 119.870 ;
        RECT 36.915 119.445 37.580 119.615 ;
        RECT 37.865 119.570 38.035 120.370 ;
        RECT 38.295 120.515 38.465 121.275 ;
        RECT 38.645 120.685 38.975 121.445 ;
        RECT 38.295 120.345 38.960 120.515 ;
        RECT 39.145 120.370 39.415 121.275 ;
        RECT 39.895 120.605 40.065 121.445 ;
        RECT 40.275 120.435 40.525 121.275 ;
        RECT 40.735 120.605 40.905 121.445 ;
        RECT 41.075 120.435 41.365 121.275 ;
        RECT 38.790 120.200 38.960 120.345 ;
        RECT 38.225 119.795 38.555 120.165 ;
        RECT 38.790 119.870 39.075 120.200 ;
        RECT 38.790 119.615 38.960 119.870 ;
        RECT 31.310 118.895 36.655 119.440 ;
        RECT 36.915 119.065 37.085 119.445 ;
        RECT 37.265 118.895 37.595 119.275 ;
        RECT 37.775 119.065 38.035 119.570 ;
        RECT 38.295 119.445 38.960 119.615 ;
        RECT 39.245 119.570 39.415 120.370 ;
        RECT 38.295 119.065 38.465 119.445 ;
        RECT 38.645 118.895 38.975 119.275 ;
        RECT 39.155 119.065 39.415 119.570 ;
        RECT 39.640 120.265 41.365 120.435 ;
        RECT 41.575 120.385 41.745 121.445 ;
        RECT 42.040 121.065 42.370 121.445 ;
        RECT 42.550 120.895 42.720 121.185 ;
        RECT 42.890 120.985 43.140 121.445 ;
        RECT 41.920 120.725 42.720 120.895 ;
        RECT 43.310 120.935 44.180 121.275 ;
        RECT 39.640 119.715 40.050 120.265 ;
        RECT 41.920 120.105 42.090 120.725 ;
        RECT 43.310 120.555 43.480 120.935 ;
        RECT 44.415 120.815 44.585 121.275 ;
        RECT 44.755 120.985 45.125 121.445 ;
        RECT 45.420 120.845 45.590 121.185 ;
        RECT 45.760 121.015 46.090 121.445 ;
        RECT 46.325 120.845 46.495 121.185 ;
        RECT 42.260 120.385 43.480 120.555 ;
        RECT 43.650 120.475 44.110 120.765 ;
        RECT 44.415 120.645 44.975 120.815 ;
        RECT 45.420 120.675 46.495 120.845 ;
        RECT 46.665 120.945 47.345 121.275 ;
        RECT 47.560 120.945 47.810 121.275 ;
        RECT 47.980 120.985 48.230 121.445 ;
        RECT 44.805 120.505 44.975 120.645 ;
        RECT 43.650 120.465 44.615 120.475 ;
        RECT 43.310 120.295 43.480 120.385 ;
        RECT 43.940 120.305 44.615 120.465 ;
        RECT 41.920 120.095 42.265 120.105 ;
        RECT 40.235 119.885 42.265 120.095 ;
        RECT 39.640 119.545 41.405 119.715 ;
        RECT 39.895 118.895 40.065 119.365 ;
        RECT 40.235 119.065 40.565 119.545 ;
        RECT 40.735 118.895 40.905 119.365 ;
        RECT 41.075 119.065 41.405 119.545 ;
        RECT 41.575 118.895 41.745 119.705 ;
        RECT 41.940 119.630 42.265 119.885 ;
        RECT 41.945 119.275 42.265 119.630 ;
        RECT 42.435 119.845 42.975 120.215 ;
        RECT 43.310 120.125 43.715 120.295 ;
        RECT 42.435 119.445 42.675 119.845 ;
        RECT 43.155 119.675 43.375 119.955 ;
        RECT 42.845 119.505 43.375 119.675 ;
        RECT 42.845 119.275 43.015 119.505 ;
        RECT 43.545 119.345 43.715 120.125 ;
        RECT 43.885 119.515 44.235 120.135 ;
        RECT 44.405 119.515 44.615 120.305 ;
        RECT 44.805 120.335 46.305 120.505 ;
        RECT 44.805 119.645 44.975 120.335 ;
        RECT 46.665 120.165 46.835 120.945 ;
        RECT 47.640 120.815 47.810 120.945 ;
        RECT 45.145 119.995 46.835 120.165 ;
        RECT 47.005 120.385 47.470 120.775 ;
        RECT 47.640 120.645 48.035 120.815 ;
        RECT 45.145 119.815 45.315 119.995 ;
        RECT 41.945 119.105 43.015 119.275 ;
        RECT 43.185 118.895 43.375 119.335 ;
        RECT 43.545 119.065 44.495 119.345 ;
        RECT 44.805 119.255 45.065 119.645 ;
        RECT 45.485 119.575 46.275 119.825 ;
        RECT 44.715 119.085 45.065 119.255 ;
        RECT 45.275 118.895 45.605 119.355 ;
        RECT 46.480 119.285 46.650 119.995 ;
        RECT 47.005 119.795 47.175 120.385 ;
        RECT 46.820 119.575 47.175 119.795 ;
        RECT 47.345 119.575 47.695 120.195 ;
        RECT 47.865 119.285 48.035 120.645 ;
        RECT 48.400 120.475 48.725 121.260 ;
        RECT 48.205 119.425 48.665 120.475 ;
        RECT 46.480 119.115 47.335 119.285 ;
        RECT 47.540 119.115 48.035 119.285 ;
        RECT 48.205 118.895 48.535 119.255 ;
        RECT 48.895 119.155 49.065 121.275 ;
        RECT 49.235 120.945 49.565 121.445 ;
        RECT 49.735 120.775 49.990 121.275 ;
        RECT 49.240 120.605 49.990 120.775 ;
        RECT 49.240 119.615 49.470 120.605 ;
        RECT 49.640 119.785 49.990 120.435 ;
        RECT 50.165 120.280 50.455 121.445 ;
        RECT 50.625 120.370 50.895 121.275 ;
        RECT 51.065 120.685 51.395 121.445 ;
        RECT 51.575 120.515 51.745 121.275 ;
        RECT 49.240 119.445 49.990 119.615 ;
        RECT 49.235 118.895 49.565 119.275 ;
        RECT 49.735 119.155 49.990 119.445 ;
        RECT 50.165 118.895 50.455 119.620 ;
        RECT 50.625 119.570 50.795 120.370 ;
        RECT 51.080 120.345 51.745 120.515 ;
        RECT 51.080 120.200 51.250 120.345 ;
        RECT 52.985 120.305 53.195 121.445 ;
        RECT 50.965 119.870 51.250 120.200 ;
        RECT 53.365 120.295 53.695 121.275 ;
        RECT 53.865 120.305 54.095 121.445 ;
        RECT 54.305 120.355 55.515 121.445 ;
        RECT 55.685 120.370 55.955 121.275 ;
        RECT 56.125 120.685 56.455 121.445 ;
        RECT 56.635 120.515 56.805 121.275 ;
        RECT 51.080 119.615 51.250 119.870 ;
        RECT 51.485 119.795 51.815 120.165 ;
        RECT 50.625 119.065 50.885 119.570 ;
        RECT 51.080 119.445 51.745 119.615 ;
        RECT 51.065 118.895 51.395 119.275 ;
        RECT 51.575 119.065 51.745 119.445 ;
        RECT 52.985 118.895 53.195 119.715 ;
        RECT 53.365 119.695 53.615 120.295 ;
        RECT 53.785 119.885 54.115 120.135 ;
        RECT 54.305 119.815 54.825 120.355 ;
        RECT 53.365 119.065 53.695 119.695 ;
        RECT 53.865 118.895 54.095 119.715 ;
        RECT 54.995 119.645 55.515 120.185 ;
        RECT 54.305 118.895 55.515 119.645 ;
        RECT 55.685 119.570 55.855 120.370 ;
        RECT 56.140 120.345 56.805 120.515 ;
        RECT 57.155 120.515 57.325 121.275 ;
        RECT 57.505 120.685 57.835 121.445 ;
        RECT 57.155 120.345 57.820 120.515 ;
        RECT 58.005 120.370 58.275 121.275 ;
        RECT 58.755 120.605 58.925 121.445 ;
        RECT 59.135 120.435 59.385 121.275 ;
        RECT 59.595 120.605 59.765 121.445 ;
        RECT 59.935 120.435 60.225 121.275 ;
        RECT 56.140 120.200 56.310 120.345 ;
        RECT 56.025 119.870 56.310 120.200 ;
        RECT 57.650 120.200 57.820 120.345 ;
        RECT 56.140 119.615 56.310 119.870 ;
        RECT 56.545 119.795 56.875 120.165 ;
        RECT 57.085 119.795 57.415 120.165 ;
        RECT 57.650 119.870 57.935 120.200 ;
        RECT 57.650 119.615 57.820 119.870 ;
        RECT 55.685 119.065 55.945 119.570 ;
        RECT 56.140 119.445 56.805 119.615 ;
        RECT 56.125 118.895 56.455 119.275 ;
        RECT 56.635 119.065 56.805 119.445 ;
        RECT 57.155 119.445 57.820 119.615 ;
        RECT 58.105 119.570 58.275 120.370 ;
        RECT 57.155 119.065 57.325 119.445 ;
        RECT 57.505 118.895 57.835 119.275 ;
        RECT 58.015 119.065 58.275 119.570 ;
        RECT 58.500 120.265 60.225 120.435 ;
        RECT 60.435 120.385 60.605 121.445 ;
        RECT 60.900 121.065 61.230 121.445 ;
        RECT 61.410 120.895 61.580 121.185 ;
        RECT 61.750 120.985 62.000 121.445 ;
        RECT 60.780 120.725 61.580 120.895 ;
        RECT 62.170 120.935 63.040 121.275 ;
        RECT 58.500 119.715 58.910 120.265 ;
        RECT 60.780 120.105 60.950 120.725 ;
        RECT 62.170 120.555 62.340 120.935 ;
        RECT 63.275 120.815 63.445 121.275 ;
        RECT 63.615 120.985 63.985 121.445 ;
        RECT 64.280 120.845 64.450 121.185 ;
        RECT 64.620 121.015 64.950 121.445 ;
        RECT 65.185 120.845 65.355 121.185 ;
        RECT 61.120 120.385 62.340 120.555 ;
        RECT 62.510 120.475 62.970 120.765 ;
        RECT 63.275 120.645 63.835 120.815 ;
        RECT 64.280 120.675 65.355 120.845 ;
        RECT 65.525 120.945 66.205 121.275 ;
        RECT 66.420 120.945 66.670 121.275 ;
        RECT 66.840 120.985 67.090 121.445 ;
        RECT 63.665 120.505 63.835 120.645 ;
        RECT 62.510 120.465 63.475 120.475 ;
        RECT 62.170 120.295 62.340 120.385 ;
        RECT 62.800 120.305 63.475 120.465 ;
        RECT 60.780 120.095 61.125 120.105 ;
        RECT 59.095 119.885 61.125 120.095 ;
        RECT 58.500 119.545 60.265 119.715 ;
        RECT 58.755 118.895 58.925 119.365 ;
        RECT 59.095 119.065 59.425 119.545 ;
        RECT 59.595 118.895 59.765 119.365 ;
        RECT 59.935 119.065 60.265 119.545 ;
        RECT 60.435 118.895 60.605 119.705 ;
        RECT 60.800 119.630 61.125 119.885 ;
        RECT 60.805 119.275 61.125 119.630 ;
        RECT 61.295 119.845 61.835 120.215 ;
        RECT 62.170 120.125 62.575 120.295 ;
        RECT 61.295 119.445 61.535 119.845 ;
        RECT 62.015 119.675 62.235 119.955 ;
        RECT 61.705 119.505 62.235 119.675 ;
        RECT 61.705 119.275 61.875 119.505 ;
        RECT 62.405 119.345 62.575 120.125 ;
        RECT 62.745 119.515 63.095 120.135 ;
        RECT 63.265 119.515 63.475 120.305 ;
        RECT 63.665 120.335 65.165 120.505 ;
        RECT 63.665 119.645 63.835 120.335 ;
        RECT 65.525 120.165 65.695 120.945 ;
        RECT 66.500 120.815 66.670 120.945 ;
        RECT 64.005 119.995 65.695 120.165 ;
        RECT 65.865 120.385 66.330 120.775 ;
        RECT 66.500 120.645 66.895 120.815 ;
        RECT 64.005 119.815 64.175 119.995 ;
        RECT 60.805 119.105 61.875 119.275 ;
        RECT 62.045 118.895 62.235 119.335 ;
        RECT 62.405 119.065 63.355 119.345 ;
        RECT 63.665 119.255 63.925 119.645 ;
        RECT 64.345 119.575 65.135 119.825 ;
        RECT 63.575 119.085 63.925 119.255 ;
        RECT 64.135 118.895 64.465 119.355 ;
        RECT 65.340 119.285 65.510 119.995 ;
        RECT 65.865 119.795 66.035 120.385 ;
        RECT 65.680 119.575 66.035 119.795 ;
        RECT 66.205 119.575 66.555 120.195 ;
        RECT 66.725 119.285 66.895 120.645 ;
        RECT 67.260 120.475 67.585 121.260 ;
        RECT 67.065 119.425 67.525 120.475 ;
        RECT 65.340 119.115 66.195 119.285 ;
        RECT 66.400 119.115 66.895 119.285 ;
        RECT 67.065 118.895 67.395 119.255 ;
        RECT 67.755 119.155 67.925 121.275 ;
        RECT 68.095 120.945 68.425 121.445 ;
        RECT 68.595 120.775 68.850 121.275 ;
        RECT 68.100 120.605 68.850 120.775 ;
        RECT 68.100 119.615 68.330 120.605 ;
        RECT 69.115 120.515 69.285 121.275 ;
        RECT 69.465 120.685 69.795 121.445 ;
        RECT 68.500 119.785 68.850 120.435 ;
        RECT 69.115 120.345 69.780 120.515 ;
        RECT 69.965 120.370 70.235 121.275 ;
        RECT 69.610 120.200 69.780 120.345 ;
        RECT 69.045 119.795 69.375 120.165 ;
        RECT 69.610 119.870 69.895 120.200 ;
        RECT 69.610 119.615 69.780 119.870 ;
        RECT 68.100 119.445 68.850 119.615 ;
        RECT 68.095 118.895 68.425 119.275 ;
        RECT 68.595 119.155 68.850 119.445 ;
        RECT 69.115 119.445 69.780 119.615 ;
        RECT 70.065 119.570 70.235 120.370 ;
        RECT 70.905 120.305 71.135 121.445 ;
        RECT 71.305 120.295 71.635 121.275 ;
        RECT 71.805 120.305 72.015 121.445 ;
        RECT 72.285 120.305 72.515 121.445 ;
        RECT 72.685 120.295 73.015 121.275 ;
        RECT 73.185 120.305 73.395 121.445 ;
        RECT 73.715 120.515 73.885 121.275 ;
        RECT 74.065 120.685 74.395 121.445 ;
        RECT 73.715 120.345 74.380 120.515 ;
        RECT 74.565 120.370 74.835 121.275 ;
        RECT 70.885 119.885 71.215 120.135 ;
        RECT 69.115 119.065 69.285 119.445 ;
        RECT 69.465 118.895 69.795 119.275 ;
        RECT 69.975 119.065 70.235 119.570 ;
        RECT 70.905 118.895 71.135 119.715 ;
        RECT 71.385 119.695 71.635 120.295 ;
        RECT 72.265 119.885 72.595 120.135 ;
        RECT 71.305 119.065 71.635 119.695 ;
        RECT 71.805 118.895 72.015 119.715 ;
        RECT 72.285 118.895 72.515 119.715 ;
        RECT 72.765 119.695 73.015 120.295 ;
        RECT 74.210 120.200 74.380 120.345 ;
        RECT 73.645 119.795 73.975 120.165 ;
        RECT 74.210 119.870 74.495 120.200 ;
        RECT 72.685 119.065 73.015 119.695 ;
        RECT 73.185 118.895 73.395 119.715 ;
        RECT 74.210 119.615 74.380 119.870 ;
        RECT 73.715 119.445 74.380 119.615 ;
        RECT 74.665 119.570 74.835 120.370 ;
        RECT 75.925 120.280 76.215 121.445 ;
        RECT 76.385 120.355 77.595 121.445 ;
        RECT 77.855 120.515 78.025 121.275 ;
        RECT 78.205 120.685 78.535 121.445 ;
        RECT 76.385 119.815 76.905 120.355 ;
        RECT 77.855 120.345 78.520 120.515 ;
        RECT 78.705 120.370 78.975 121.275 ;
        RECT 79.455 120.605 79.625 121.445 ;
        RECT 79.835 120.435 80.085 121.275 ;
        RECT 80.295 120.605 80.465 121.445 ;
        RECT 80.635 120.435 80.925 121.275 ;
        RECT 78.350 120.200 78.520 120.345 ;
        RECT 77.075 119.645 77.595 120.185 ;
        RECT 77.785 119.795 78.115 120.165 ;
        RECT 78.350 119.870 78.635 120.200 ;
        RECT 73.715 119.065 73.885 119.445 ;
        RECT 74.065 118.895 74.395 119.275 ;
        RECT 74.575 119.065 74.835 119.570 ;
        RECT 75.925 118.895 76.215 119.620 ;
        RECT 76.385 118.895 77.595 119.645 ;
        RECT 78.350 119.615 78.520 119.870 ;
        RECT 77.855 119.445 78.520 119.615 ;
        RECT 78.805 119.570 78.975 120.370 ;
        RECT 77.855 119.065 78.025 119.445 ;
        RECT 78.205 118.895 78.535 119.275 ;
        RECT 78.715 119.065 78.975 119.570 ;
        RECT 79.200 120.265 80.925 120.435 ;
        RECT 81.135 120.385 81.305 121.445 ;
        RECT 81.600 121.065 81.930 121.445 ;
        RECT 82.110 120.895 82.280 121.185 ;
        RECT 82.450 120.985 82.700 121.445 ;
        RECT 81.480 120.725 82.280 120.895 ;
        RECT 82.870 120.935 83.740 121.275 ;
        RECT 79.200 119.715 79.610 120.265 ;
        RECT 81.480 120.105 81.650 120.725 ;
        RECT 82.870 120.555 83.040 120.935 ;
        RECT 83.975 120.815 84.145 121.275 ;
        RECT 84.315 120.985 84.685 121.445 ;
        RECT 84.980 120.845 85.150 121.185 ;
        RECT 85.320 121.015 85.650 121.445 ;
        RECT 85.885 120.845 86.055 121.185 ;
        RECT 81.820 120.385 83.040 120.555 ;
        RECT 83.210 120.475 83.670 120.765 ;
        RECT 83.975 120.645 84.535 120.815 ;
        RECT 84.980 120.675 86.055 120.845 ;
        RECT 86.225 120.945 86.905 121.275 ;
        RECT 87.120 120.945 87.370 121.275 ;
        RECT 87.540 120.985 87.790 121.445 ;
        RECT 84.365 120.505 84.535 120.645 ;
        RECT 83.210 120.465 84.175 120.475 ;
        RECT 82.870 120.295 83.040 120.385 ;
        RECT 83.500 120.305 84.175 120.465 ;
        RECT 81.480 120.095 81.825 120.105 ;
        RECT 79.795 119.885 81.825 120.095 ;
        RECT 79.200 119.545 80.965 119.715 ;
        RECT 79.455 118.895 79.625 119.365 ;
        RECT 79.795 119.065 80.125 119.545 ;
        RECT 80.295 118.895 80.465 119.365 ;
        RECT 80.635 119.065 80.965 119.545 ;
        RECT 81.135 118.895 81.305 119.705 ;
        RECT 81.500 119.630 81.825 119.885 ;
        RECT 81.505 119.275 81.825 119.630 ;
        RECT 81.995 119.845 82.535 120.215 ;
        RECT 82.870 120.125 83.275 120.295 ;
        RECT 81.995 119.445 82.235 119.845 ;
        RECT 82.715 119.675 82.935 119.955 ;
        RECT 82.405 119.505 82.935 119.675 ;
        RECT 82.405 119.275 82.575 119.505 ;
        RECT 83.105 119.345 83.275 120.125 ;
        RECT 83.445 119.515 83.795 120.135 ;
        RECT 83.965 119.515 84.175 120.305 ;
        RECT 84.365 120.335 85.865 120.505 ;
        RECT 84.365 119.645 84.535 120.335 ;
        RECT 86.225 120.165 86.395 120.945 ;
        RECT 87.200 120.815 87.370 120.945 ;
        RECT 84.705 119.995 86.395 120.165 ;
        RECT 86.565 120.385 87.030 120.775 ;
        RECT 87.200 120.645 87.595 120.815 ;
        RECT 84.705 119.815 84.875 119.995 ;
        RECT 81.505 119.105 82.575 119.275 ;
        RECT 82.745 118.895 82.935 119.335 ;
        RECT 83.105 119.065 84.055 119.345 ;
        RECT 84.365 119.255 84.625 119.645 ;
        RECT 85.045 119.575 85.835 119.825 ;
        RECT 84.275 119.085 84.625 119.255 ;
        RECT 84.835 118.895 85.165 119.355 ;
        RECT 86.040 119.285 86.210 119.995 ;
        RECT 86.565 119.795 86.735 120.385 ;
        RECT 86.380 119.575 86.735 119.795 ;
        RECT 86.905 119.575 87.255 120.195 ;
        RECT 87.425 119.285 87.595 120.645 ;
        RECT 87.960 120.475 88.285 121.260 ;
        RECT 87.765 119.425 88.225 120.475 ;
        RECT 86.040 119.115 86.895 119.285 ;
        RECT 87.100 119.115 87.595 119.285 ;
        RECT 87.765 118.895 88.095 119.255 ;
        RECT 88.455 119.155 88.625 121.275 ;
        RECT 88.795 120.945 89.125 121.445 ;
        RECT 89.295 120.775 89.550 121.275 ;
        RECT 88.800 120.605 89.550 120.775 ;
        RECT 88.800 119.615 89.030 120.605 ;
        RECT 89.815 120.515 89.985 121.275 ;
        RECT 90.165 120.685 90.495 121.445 ;
        RECT 89.200 119.785 89.550 120.435 ;
        RECT 89.815 120.345 90.480 120.515 ;
        RECT 90.665 120.370 90.935 121.275 ;
        RECT 91.415 120.605 91.585 121.445 ;
        RECT 91.795 120.435 92.045 121.275 ;
        RECT 92.255 120.605 92.425 121.445 ;
        RECT 92.595 120.435 92.885 121.275 ;
        RECT 90.310 120.200 90.480 120.345 ;
        RECT 89.745 119.795 90.075 120.165 ;
        RECT 90.310 119.870 90.595 120.200 ;
        RECT 90.310 119.615 90.480 119.870 ;
        RECT 88.800 119.445 89.550 119.615 ;
        RECT 88.795 118.895 89.125 119.275 ;
        RECT 89.295 119.155 89.550 119.445 ;
        RECT 89.815 119.445 90.480 119.615 ;
        RECT 90.765 119.570 90.935 120.370 ;
        RECT 89.815 119.065 89.985 119.445 ;
        RECT 90.165 118.895 90.495 119.275 ;
        RECT 90.675 119.065 90.935 119.570 ;
        RECT 91.160 120.265 92.885 120.435 ;
        RECT 93.095 120.385 93.265 121.445 ;
        RECT 93.560 121.065 93.890 121.445 ;
        RECT 94.070 120.895 94.240 121.185 ;
        RECT 94.410 120.985 94.660 121.445 ;
        RECT 93.440 120.725 94.240 120.895 ;
        RECT 94.830 120.935 95.700 121.275 ;
        RECT 91.160 119.715 91.570 120.265 ;
        RECT 93.440 120.105 93.610 120.725 ;
        RECT 94.830 120.555 95.000 120.935 ;
        RECT 95.935 120.815 96.105 121.275 ;
        RECT 96.275 120.985 96.645 121.445 ;
        RECT 96.940 120.845 97.110 121.185 ;
        RECT 97.280 121.015 97.610 121.445 ;
        RECT 97.845 120.845 98.015 121.185 ;
        RECT 93.780 120.385 95.000 120.555 ;
        RECT 95.170 120.475 95.630 120.765 ;
        RECT 95.935 120.645 96.495 120.815 ;
        RECT 96.940 120.675 98.015 120.845 ;
        RECT 98.185 120.945 98.865 121.275 ;
        RECT 99.080 120.945 99.330 121.275 ;
        RECT 99.500 120.985 99.750 121.445 ;
        RECT 96.325 120.505 96.495 120.645 ;
        RECT 95.170 120.465 96.135 120.475 ;
        RECT 94.830 120.295 95.000 120.385 ;
        RECT 95.460 120.305 96.135 120.465 ;
        RECT 93.440 120.095 93.785 120.105 ;
        RECT 91.755 119.885 93.785 120.095 ;
        RECT 91.160 119.545 92.925 119.715 ;
        RECT 91.415 118.895 91.585 119.365 ;
        RECT 91.755 119.065 92.085 119.545 ;
        RECT 92.255 118.895 92.425 119.365 ;
        RECT 92.595 119.065 92.925 119.545 ;
        RECT 93.095 118.895 93.265 119.705 ;
        RECT 93.460 119.630 93.785 119.885 ;
        RECT 93.465 119.275 93.785 119.630 ;
        RECT 93.955 119.845 94.495 120.215 ;
        RECT 94.830 120.125 95.235 120.295 ;
        RECT 93.955 119.445 94.195 119.845 ;
        RECT 94.675 119.675 94.895 119.955 ;
        RECT 94.365 119.505 94.895 119.675 ;
        RECT 94.365 119.275 94.535 119.505 ;
        RECT 95.065 119.345 95.235 120.125 ;
        RECT 95.405 119.515 95.755 120.135 ;
        RECT 95.925 119.515 96.135 120.305 ;
        RECT 96.325 120.335 97.825 120.505 ;
        RECT 96.325 119.645 96.495 120.335 ;
        RECT 98.185 120.165 98.355 120.945 ;
        RECT 99.160 120.815 99.330 120.945 ;
        RECT 96.665 119.995 98.355 120.165 ;
        RECT 98.525 120.385 98.990 120.775 ;
        RECT 99.160 120.645 99.555 120.815 ;
        RECT 96.665 119.815 96.835 119.995 ;
        RECT 93.465 119.105 94.535 119.275 ;
        RECT 94.705 118.895 94.895 119.335 ;
        RECT 95.065 119.065 96.015 119.345 ;
        RECT 96.325 119.255 96.585 119.645 ;
        RECT 97.005 119.575 97.795 119.825 ;
        RECT 96.235 119.085 96.585 119.255 ;
        RECT 96.795 118.895 97.125 119.355 ;
        RECT 98.000 119.285 98.170 119.995 ;
        RECT 98.525 119.795 98.695 120.385 ;
        RECT 98.340 119.575 98.695 119.795 ;
        RECT 98.865 119.575 99.215 120.195 ;
        RECT 99.385 119.285 99.555 120.645 ;
        RECT 99.920 120.475 100.245 121.260 ;
        RECT 99.725 119.425 100.185 120.475 ;
        RECT 98.000 119.115 98.855 119.285 ;
        RECT 99.060 119.115 99.555 119.285 ;
        RECT 99.725 118.895 100.055 119.255 ;
        RECT 100.415 119.155 100.585 121.275 ;
        RECT 100.755 120.945 101.085 121.445 ;
        RECT 101.255 120.775 101.510 121.275 ;
        RECT 100.760 120.605 101.510 120.775 ;
        RECT 100.760 119.615 100.990 120.605 ;
        RECT 101.160 119.785 101.510 120.435 ;
        RECT 101.685 120.280 101.975 121.445 ;
        RECT 103.375 120.605 103.545 121.445 ;
        RECT 103.755 120.435 104.005 121.275 ;
        RECT 104.215 120.605 104.385 121.445 ;
        RECT 104.555 120.435 104.845 121.275 ;
        RECT 103.120 120.265 104.845 120.435 ;
        RECT 105.055 120.385 105.225 121.445 ;
        RECT 105.520 121.065 105.850 121.445 ;
        RECT 106.030 120.895 106.200 121.185 ;
        RECT 106.370 120.985 106.620 121.445 ;
        RECT 105.400 120.725 106.200 120.895 ;
        RECT 106.790 120.935 107.660 121.275 ;
        RECT 103.120 119.715 103.530 120.265 ;
        RECT 105.400 120.105 105.570 120.725 ;
        RECT 106.790 120.555 106.960 120.935 ;
        RECT 107.895 120.815 108.065 121.275 ;
        RECT 108.235 120.985 108.605 121.445 ;
        RECT 108.900 120.845 109.070 121.185 ;
        RECT 109.240 121.015 109.570 121.445 ;
        RECT 109.805 120.845 109.975 121.185 ;
        RECT 105.740 120.385 106.960 120.555 ;
        RECT 107.130 120.475 107.590 120.765 ;
        RECT 107.895 120.645 108.455 120.815 ;
        RECT 108.900 120.675 109.975 120.845 ;
        RECT 110.145 120.945 110.825 121.275 ;
        RECT 111.040 120.945 111.290 121.275 ;
        RECT 111.460 120.985 111.710 121.445 ;
        RECT 108.285 120.505 108.455 120.645 ;
        RECT 107.130 120.465 108.095 120.475 ;
        RECT 106.790 120.295 106.960 120.385 ;
        RECT 107.420 120.305 108.095 120.465 ;
        RECT 105.400 120.095 105.745 120.105 ;
        RECT 103.715 119.885 105.745 120.095 ;
        RECT 100.760 119.445 101.510 119.615 ;
        RECT 100.755 118.895 101.085 119.275 ;
        RECT 101.255 119.155 101.510 119.445 ;
        RECT 101.685 118.895 101.975 119.620 ;
        RECT 103.120 119.545 104.885 119.715 ;
        RECT 103.375 118.895 103.545 119.365 ;
        RECT 103.715 119.065 104.045 119.545 ;
        RECT 104.215 118.895 104.385 119.365 ;
        RECT 104.555 119.065 104.885 119.545 ;
        RECT 105.055 118.895 105.225 119.705 ;
        RECT 105.420 119.630 105.745 119.885 ;
        RECT 105.425 119.275 105.745 119.630 ;
        RECT 105.915 119.845 106.455 120.215 ;
        RECT 106.790 120.125 107.195 120.295 ;
        RECT 105.915 119.445 106.155 119.845 ;
        RECT 106.635 119.675 106.855 119.955 ;
        RECT 106.325 119.505 106.855 119.675 ;
        RECT 106.325 119.275 106.495 119.505 ;
        RECT 107.025 119.345 107.195 120.125 ;
        RECT 107.365 119.515 107.715 120.135 ;
        RECT 107.885 119.515 108.095 120.305 ;
        RECT 108.285 120.335 109.785 120.505 ;
        RECT 108.285 119.645 108.455 120.335 ;
        RECT 110.145 120.165 110.315 120.945 ;
        RECT 111.120 120.815 111.290 120.945 ;
        RECT 108.625 119.995 110.315 120.165 ;
        RECT 110.485 120.385 110.950 120.775 ;
        RECT 111.120 120.645 111.515 120.815 ;
        RECT 108.625 119.815 108.795 119.995 ;
        RECT 105.425 119.105 106.495 119.275 ;
        RECT 106.665 118.895 106.855 119.335 ;
        RECT 107.025 119.065 107.975 119.345 ;
        RECT 108.285 119.255 108.545 119.645 ;
        RECT 108.965 119.575 109.755 119.825 ;
        RECT 108.195 119.085 108.545 119.255 ;
        RECT 108.755 118.895 109.085 119.355 ;
        RECT 109.960 119.285 110.130 119.995 ;
        RECT 110.485 119.795 110.655 120.385 ;
        RECT 110.300 119.575 110.655 119.795 ;
        RECT 110.825 119.575 111.175 120.195 ;
        RECT 111.345 119.285 111.515 120.645 ;
        RECT 111.880 120.475 112.205 121.260 ;
        RECT 111.685 119.425 112.145 120.475 ;
        RECT 109.960 119.115 110.815 119.285 ;
        RECT 111.020 119.115 111.515 119.285 ;
        RECT 111.685 118.895 112.015 119.255 ;
        RECT 112.375 119.155 112.545 121.275 ;
        RECT 112.715 120.945 113.045 121.445 ;
        RECT 113.215 120.775 113.470 121.275 ;
        RECT 112.720 120.605 113.470 120.775 ;
        RECT 112.720 119.615 112.950 120.605 ;
        RECT 113.120 119.785 113.470 120.435 ;
        RECT 113.645 120.370 113.915 121.275 ;
        RECT 114.085 120.685 114.415 121.445 ;
        RECT 114.595 120.515 114.765 121.275 ;
        RECT 116.255 120.605 116.425 121.445 ;
        RECT 112.720 119.445 113.470 119.615 ;
        RECT 112.715 118.895 113.045 119.275 ;
        RECT 113.215 119.155 113.470 119.445 ;
        RECT 113.645 119.570 113.815 120.370 ;
        RECT 114.100 120.345 114.765 120.515 ;
        RECT 116.635 120.435 116.885 121.275 ;
        RECT 117.095 120.605 117.265 121.445 ;
        RECT 117.435 120.435 117.725 121.275 ;
        RECT 114.100 120.200 114.270 120.345 ;
        RECT 113.985 119.870 114.270 120.200 ;
        RECT 116.000 120.265 117.725 120.435 ;
        RECT 117.935 120.385 118.105 121.445 ;
        RECT 118.400 121.065 118.730 121.445 ;
        RECT 118.910 120.895 119.080 121.185 ;
        RECT 119.250 120.985 119.500 121.445 ;
        RECT 118.280 120.725 119.080 120.895 ;
        RECT 119.670 120.935 120.540 121.275 ;
        RECT 114.100 119.615 114.270 119.870 ;
        RECT 114.505 119.795 114.835 120.165 ;
        RECT 116.000 119.715 116.410 120.265 ;
        RECT 118.280 120.105 118.450 120.725 ;
        RECT 119.670 120.555 119.840 120.935 ;
        RECT 120.775 120.815 120.945 121.275 ;
        RECT 121.115 120.985 121.485 121.445 ;
        RECT 121.780 120.845 121.950 121.185 ;
        RECT 122.120 121.015 122.450 121.445 ;
        RECT 122.685 120.845 122.855 121.185 ;
        RECT 118.620 120.385 119.840 120.555 ;
        RECT 120.010 120.475 120.470 120.765 ;
        RECT 120.775 120.645 121.335 120.815 ;
        RECT 121.780 120.675 122.855 120.845 ;
        RECT 123.025 120.945 123.705 121.275 ;
        RECT 123.920 120.945 124.170 121.275 ;
        RECT 124.340 120.985 124.590 121.445 ;
        RECT 121.165 120.505 121.335 120.645 ;
        RECT 120.010 120.465 120.975 120.475 ;
        RECT 119.670 120.295 119.840 120.385 ;
        RECT 120.300 120.305 120.975 120.465 ;
        RECT 118.280 120.095 118.625 120.105 ;
        RECT 116.595 119.885 118.625 120.095 ;
        RECT 113.645 119.065 113.905 119.570 ;
        RECT 114.100 119.445 114.765 119.615 ;
        RECT 116.000 119.545 117.765 119.715 ;
        RECT 114.085 118.895 114.415 119.275 ;
        RECT 114.595 119.065 114.765 119.445 ;
        RECT 116.255 118.895 116.425 119.365 ;
        RECT 116.595 119.065 116.925 119.545 ;
        RECT 117.095 118.895 117.265 119.365 ;
        RECT 117.435 119.065 117.765 119.545 ;
        RECT 117.935 118.895 118.105 119.705 ;
        RECT 118.300 119.630 118.625 119.885 ;
        RECT 118.305 119.275 118.625 119.630 ;
        RECT 118.795 119.845 119.335 120.215 ;
        RECT 119.670 120.125 120.075 120.295 ;
        RECT 118.795 119.445 119.035 119.845 ;
        RECT 119.515 119.675 119.735 119.955 ;
        RECT 119.205 119.505 119.735 119.675 ;
        RECT 119.205 119.275 119.375 119.505 ;
        RECT 119.905 119.345 120.075 120.125 ;
        RECT 120.245 119.515 120.595 120.135 ;
        RECT 120.765 119.515 120.975 120.305 ;
        RECT 121.165 120.335 122.665 120.505 ;
        RECT 121.165 119.645 121.335 120.335 ;
        RECT 123.025 120.165 123.195 120.945 ;
        RECT 124.000 120.815 124.170 120.945 ;
        RECT 121.505 119.995 123.195 120.165 ;
        RECT 123.365 120.385 123.830 120.775 ;
        RECT 124.000 120.645 124.395 120.815 ;
        RECT 121.505 119.815 121.675 119.995 ;
        RECT 118.305 119.105 119.375 119.275 ;
        RECT 119.545 118.895 119.735 119.335 ;
        RECT 119.905 119.065 120.855 119.345 ;
        RECT 121.165 119.255 121.425 119.645 ;
        RECT 121.845 119.575 122.635 119.825 ;
        RECT 121.075 119.085 121.425 119.255 ;
        RECT 121.635 118.895 121.965 119.355 ;
        RECT 122.840 119.285 123.010 119.995 ;
        RECT 123.365 119.795 123.535 120.385 ;
        RECT 123.180 119.575 123.535 119.795 ;
        RECT 123.705 119.575 124.055 120.195 ;
        RECT 124.225 119.285 124.395 120.645 ;
        RECT 124.760 120.475 125.085 121.260 ;
        RECT 124.565 119.425 125.025 120.475 ;
        RECT 122.840 119.115 123.695 119.285 ;
        RECT 123.900 119.115 124.395 119.285 ;
        RECT 124.565 118.895 124.895 119.255 ;
        RECT 125.255 119.155 125.425 121.275 ;
        RECT 125.595 120.945 125.925 121.445 ;
        RECT 126.095 120.775 126.350 121.275 ;
        RECT 125.600 120.605 126.350 120.775 ;
        RECT 125.600 119.615 125.830 120.605 ;
        RECT 126.000 119.785 126.350 120.435 ;
        RECT 126.525 120.355 127.735 121.445 ;
        RECT 126.525 119.815 127.045 120.355 ;
        RECT 127.215 119.645 127.735 120.185 ;
        RECT 125.600 119.445 126.350 119.615 ;
        RECT 125.595 118.895 125.925 119.275 ;
        RECT 126.095 119.155 126.350 119.445 ;
        RECT 126.525 118.895 127.735 119.645 ;
        RECT 29.840 118.725 127.820 118.895 ;
        RECT 29.925 117.975 31.135 118.725 ;
        RECT 29.925 117.435 30.445 117.975 ;
        RECT 31.765 117.955 35.275 118.725 ;
        RECT 30.615 117.265 31.135 117.805 ;
        RECT 29.925 116.175 31.135 117.265 ;
        RECT 31.765 117.265 33.455 117.785 ;
        RECT 33.625 117.435 35.275 117.955 ;
        RECT 35.505 117.905 35.715 118.725 ;
        RECT 35.885 117.925 36.215 118.555 ;
        RECT 35.885 117.325 36.135 117.925 ;
        RECT 36.385 117.905 36.615 118.725 ;
        RECT 37.285 118.000 37.575 118.725 ;
        RECT 37.785 117.905 38.015 118.725 ;
        RECT 38.185 117.925 38.515 118.555 ;
        RECT 36.305 117.485 36.635 117.735 ;
        RECT 37.765 117.485 38.095 117.735 ;
        RECT 31.765 116.175 35.275 117.265 ;
        RECT 35.505 116.175 35.715 117.315 ;
        RECT 35.885 116.345 36.215 117.325 ;
        RECT 36.385 116.175 36.615 117.315 ;
        RECT 37.285 116.175 37.575 117.340 ;
        RECT 38.265 117.325 38.515 117.925 ;
        RECT 38.685 117.905 38.895 118.725 ;
        RECT 39.165 117.905 39.395 118.725 ;
        RECT 39.565 117.925 39.895 118.555 ;
        RECT 39.145 117.485 39.475 117.735 ;
        RECT 39.645 117.325 39.895 117.925 ;
        RECT 40.065 117.905 40.275 118.725 ;
        RECT 40.545 117.905 40.775 118.725 ;
        RECT 40.945 117.925 41.275 118.555 ;
        RECT 40.525 117.485 40.855 117.735 ;
        RECT 41.025 117.325 41.275 117.925 ;
        RECT 41.445 117.905 41.655 118.725 ;
        RECT 41.890 118.175 42.145 118.465 ;
        RECT 42.315 118.345 42.645 118.725 ;
        RECT 41.890 118.005 42.640 118.175 ;
        RECT 37.785 116.175 38.015 117.315 ;
        RECT 38.185 116.345 38.515 117.325 ;
        RECT 38.685 116.175 38.895 117.315 ;
        RECT 39.165 116.175 39.395 117.315 ;
        RECT 39.565 116.345 39.895 117.325 ;
        RECT 40.065 116.175 40.275 117.315 ;
        RECT 40.545 116.175 40.775 117.315 ;
        RECT 40.945 116.345 41.275 117.325 ;
        RECT 41.445 116.175 41.655 117.315 ;
        RECT 41.890 117.185 42.240 117.835 ;
        RECT 42.410 117.015 42.640 118.005 ;
        RECT 41.890 116.845 42.640 117.015 ;
        RECT 41.890 116.345 42.145 116.845 ;
        RECT 42.315 116.175 42.645 116.675 ;
        RECT 42.815 116.345 42.985 118.465 ;
        RECT 43.345 118.365 43.675 118.725 ;
        RECT 43.845 118.335 44.340 118.505 ;
        RECT 44.545 118.335 45.400 118.505 ;
        RECT 43.215 117.145 43.675 118.195 ;
        RECT 43.155 116.360 43.480 117.145 ;
        RECT 43.845 116.975 44.015 118.335 ;
        RECT 44.185 117.425 44.535 118.045 ;
        RECT 44.705 117.825 45.060 118.045 ;
        RECT 44.705 117.235 44.875 117.825 ;
        RECT 45.230 117.625 45.400 118.335 ;
        RECT 46.275 118.265 46.605 118.725 ;
        RECT 46.815 118.365 47.165 118.535 ;
        RECT 45.605 117.795 46.395 118.045 ;
        RECT 46.815 117.975 47.075 118.365 ;
        RECT 47.385 118.275 48.335 118.555 ;
        RECT 48.505 118.285 48.695 118.725 ;
        RECT 48.865 118.345 49.935 118.515 ;
        RECT 46.565 117.625 46.735 117.805 ;
        RECT 43.845 116.805 44.240 116.975 ;
        RECT 44.410 116.845 44.875 117.235 ;
        RECT 45.045 117.455 46.735 117.625 ;
        RECT 44.070 116.675 44.240 116.805 ;
        RECT 45.045 116.675 45.215 117.455 ;
        RECT 46.905 117.285 47.075 117.975 ;
        RECT 45.575 117.115 47.075 117.285 ;
        RECT 47.265 117.315 47.475 118.105 ;
        RECT 47.645 117.485 47.995 118.105 ;
        RECT 48.165 117.495 48.335 118.275 ;
        RECT 48.865 118.115 49.035 118.345 ;
        RECT 48.505 117.945 49.035 118.115 ;
        RECT 48.505 117.665 48.725 117.945 ;
        RECT 49.205 117.775 49.445 118.175 ;
        RECT 48.165 117.325 48.570 117.495 ;
        RECT 48.905 117.405 49.445 117.775 ;
        RECT 49.615 117.990 49.935 118.345 ;
        RECT 49.615 117.735 49.940 117.990 ;
        RECT 50.135 117.915 50.305 118.725 ;
        RECT 50.475 118.075 50.805 118.555 ;
        RECT 50.975 118.255 51.145 118.725 ;
        RECT 51.315 118.075 51.645 118.555 ;
        RECT 51.815 118.255 51.985 118.725 ;
        RECT 52.775 118.255 52.945 118.725 ;
        RECT 53.115 118.075 53.445 118.555 ;
        RECT 53.615 118.255 53.785 118.725 ;
        RECT 53.955 118.075 54.285 118.555 ;
        RECT 50.475 117.905 52.240 118.075 ;
        RECT 49.615 117.525 51.645 117.735 ;
        RECT 49.615 117.515 49.960 117.525 ;
        RECT 47.265 117.155 47.940 117.315 ;
        RECT 48.400 117.235 48.570 117.325 ;
        RECT 47.265 117.145 48.230 117.155 ;
        RECT 46.905 116.975 47.075 117.115 ;
        RECT 43.650 116.175 43.900 116.635 ;
        RECT 44.070 116.345 44.320 116.675 ;
        RECT 44.535 116.345 45.215 116.675 ;
        RECT 45.385 116.775 46.460 116.945 ;
        RECT 46.905 116.805 47.465 116.975 ;
        RECT 47.770 116.855 48.230 117.145 ;
        RECT 48.400 117.065 49.620 117.235 ;
        RECT 45.385 116.435 45.555 116.775 ;
        RECT 45.790 116.175 46.120 116.605 ;
        RECT 46.290 116.435 46.460 116.775 ;
        RECT 46.755 116.175 47.125 116.635 ;
        RECT 47.295 116.345 47.465 116.805 ;
        RECT 48.400 116.685 48.570 117.065 ;
        RECT 49.790 116.895 49.960 117.515 ;
        RECT 51.830 117.355 52.240 117.905 ;
        RECT 47.700 116.345 48.570 116.685 ;
        RECT 49.160 116.725 49.960 116.895 ;
        RECT 48.740 116.175 48.990 116.635 ;
        RECT 49.160 116.435 49.330 116.725 ;
        RECT 49.510 116.175 49.840 116.555 ;
        RECT 50.135 116.175 50.305 117.235 ;
        RECT 50.515 117.185 52.240 117.355 ;
        RECT 52.520 117.905 54.285 118.075 ;
        RECT 54.455 117.915 54.625 118.725 ;
        RECT 54.825 118.345 55.895 118.515 ;
        RECT 54.825 117.990 55.145 118.345 ;
        RECT 52.520 117.355 52.930 117.905 ;
        RECT 54.820 117.735 55.145 117.990 ;
        RECT 53.115 117.525 55.145 117.735 ;
        RECT 54.800 117.515 55.145 117.525 ;
        RECT 55.315 117.775 55.555 118.175 ;
        RECT 55.725 118.115 55.895 118.345 ;
        RECT 56.065 118.285 56.255 118.725 ;
        RECT 56.425 118.275 57.375 118.555 ;
        RECT 57.595 118.365 57.945 118.535 ;
        RECT 55.725 117.945 56.255 118.115 ;
        RECT 52.520 117.185 54.245 117.355 ;
        RECT 50.515 116.345 50.805 117.185 ;
        RECT 50.975 116.175 51.145 117.015 ;
        RECT 51.355 116.345 51.605 117.185 ;
        RECT 51.815 116.175 51.985 117.015 ;
        RECT 52.775 116.175 52.945 117.015 ;
        RECT 53.155 116.345 53.405 117.185 ;
        RECT 53.615 116.175 53.785 117.015 ;
        RECT 53.955 116.345 54.245 117.185 ;
        RECT 54.455 116.175 54.625 117.235 ;
        RECT 54.800 116.895 54.970 117.515 ;
        RECT 55.315 117.405 55.855 117.775 ;
        RECT 56.035 117.665 56.255 117.945 ;
        RECT 56.425 117.495 56.595 118.275 ;
        RECT 56.190 117.325 56.595 117.495 ;
        RECT 56.765 117.485 57.115 118.105 ;
        RECT 56.190 117.235 56.360 117.325 ;
        RECT 57.285 117.315 57.495 118.105 ;
        RECT 55.140 117.065 56.360 117.235 ;
        RECT 56.820 117.155 57.495 117.315 ;
        RECT 54.800 116.725 55.600 116.895 ;
        RECT 54.920 116.175 55.250 116.555 ;
        RECT 55.430 116.435 55.600 116.725 ;
        RECT 56.190 116.685 56.360 117.065 ;
        RECT 56.530 117.145 57.495 117.155 ;
        RECT 57.685 117.975 57.945 118.365 ;
        RECT 58.155 118.265 58.485 118.725 ;
        RECT 59.360 118.335 60.215 118.505 ;
        RECT 60.420 118.335 60.915 118.505 ;
        RECT 61.085 118.365 61.415 118.725 ;
        RECT 57.685 117.285 57.855 117.975 ;
        RECT 58.025 117.625 58.195 117.805 ;
        RECT 58.365 117.795 59.155 118.045 ;
        RECT 59.360 117.625 59.530 118.335 ;
        RECT 59.700 117.825 60.055 118.045 ;
        RECT 58.025 117.455 59.715 117.625 ;
        RECT 56.530 116.855 56.990 117.145 ;
        RECT 57.685 117.115 59.185 117.285 ;
        RECT 57.685 116.975 57.855 117.115 ;
        RECT 57.295 116.805 57.855 116.975 ;
        RECT 55.770 116.175 56.020 116.635 ;
        RECT 56.190 116.345 57.060 116.685 ;
        RECT 57.295 116.345 57.465 116.805 ;
        RECT 58.300 116.775 59.375 116.945 ;
        RECT 57.635 116.175 58.005 116.635 ;
        RECT 58.300 116.435 58.470 116.775 ;
        RECT 58.640 116.175 58.970 116.605 ;
        RECT 59.205 116.435 59.375 116.775 ;
        RECT 59.545 116.675 59.715 117.455 ;
        RECT 59.885 117.235 60.055 117.825 ;
        RECT 60.225 117.425 60.575 118.045 ;
        RECT 59.885 116.845 60.350 117.235 ;
        RECT 60.745 116.975 60.915 118.335 ;
        RECT 61.085 117.145 61.545 118.195 ;
        RECT 60.520 116.805 60.915 116.975 ;
        RECT 60.520 116.675 60.690 116.805 ;
        RECT 59.545 116.345 60.225 116.675 ;
        RECT 60.440 116.345 60.690 116.675 ;
        RECT 60.860 116.175 61.110 116.635 ;
        RECT 61.280 116.360 61.605 117.145 ;
        RECT 61.775 116.345 61.945 118.465 ;
        RECT 62.115 118.345 62.445 118.725 ;
        RECT 62.615 118.175 62.870 118.465 ;
        RECT 62.120 118.005 62.870 118.175 ;
        RECT 62.120 117.015 62.350 118.005 ;
        RECT 63.045 118.000 63.335 118.725 ;
        RECT 63.815 118.255 63.985 118.725 ;
        RECT 64.155 118.075 64.485 118.555 ;
        RECT 64.655 118.255 64.825 118.725 ;
        RECT 64.995 118.075 65.325 118.555 ;
        RECT 63.560 117.905 65.325 118.075 ;
        RECT 65.495 117.915 65.665 118.725 ;
        RECT 65.865 118.345 66.935 118.515 ;
        RECT 65.865 117.990 66.185 118.345 ;
        RECT 62.520 117.185 62.870 117.835 ;
        RECT 63.560 117.355 63.970 117.905 ;
        RECT 65.860 117.735 66.185 117.990 ;
        RECT 64.155 117.525 66.185 117.735 ;
        RECT 65.840 117.515 66.185 117.525 ;
        RECT 66.355 117.775 66.595 118.175 ;
        RECT 66.765 118.115 66.935 118.345 ;
        RECT 67.105 118.285 67.295 118.725 ;
        RECT 67.465 118.275 68.415 118.555 ;
        RECT 68.635 118.365 68.985 118.535 ;
        RECT 66.765 117.945 67.295 118.115 ;
        RECT 62.120 116.845 62.870 117.015 ;
        RECT 62.115 116.175 62.445 116.675 ;
        RECT 62.615 116.345 62.870 116.845 ;
        RECT 63.045 116.175 63.335 117.340 ;
        RECT 63.560 117.185 65.285 117.355 ;
        RECT 63.815 116.175 63.985 117.015 ;
        RECT 64.195 116.345 64.445 117.185 ;
        RECT 64.655 116.175 64.825 117.015 ;
        RECT 64.995 116.345 65.285 117.185 ;
        RECT 65.495 116.175 65.665 117.235 ;
        RECT 65.840 116.895 66.010 117.515 ;
        RECT 66.355 117.405 66.895 117.775 ;
        RECT 67.075 117.665 67.295 117.945 ;
        RECT 67.465 117.495 67.635 118.275 ;
        RECT 67.230 117.325 67.635 117.495 ;
        RECT 67.805 117.485 68.155 118.105 ;
        RECT 67.230 117.235 67.400 117.325 ;
        RECT 68.325 117.315 68.535 118.105 ;
        RECT 66.180 117.065 67.400 117.235 ;
        RECT 67.860 117.155 68.535 117.315 ;
        RECT 65.840 116.725 66.640 116.895 ;
        RECT 65.960 116.175 66.290 116.555 ;
        RECT 66.470 116.435 66.640 116.725 ;
        RECT 67.230 116.685 67.400 117.065 ;
        RECT 67.570 117.145 68.535 117.155 ;
        RECT 68.725 117.975 68.985 118.365 ;
        RECT 69.195 118.265 69.525 118.725 ;
        RECT 70.400 118.335 71.255 118.505 ;
        RECT 71.460 118.335 71.955 118.505 ;
        RECT 72.125 118.365 72.455 118.725 ;
        RECT 68.725 117.285 68.895 117.975 ;
        RECT 69.065 117.625 69.235 117.805 ;
        RECT 69.405 117.795 70.195 118.045 ;
        RECT 70.400 117.625 70.570 118.335 ;
        RECT 70.740 117.825 71.095 118.045 ;
        RECT 69.065 117.455 70.755 117.625 ;
        RECT 67.570 116.855 68.030 117.145 ;
        RECT 68.725 117.115 70.225 117.285 ;
        RECT 68.725 116.975 68.895 117.115 ;
        RECT 68.335 116.805 68.895 116.975 ;
        RECT 66.810 116.175 67.060 116.635 ;
        RECT 67.230 116.345 68.100 116.685 ;
        RECT 68.335 116.345 68.505 116.805 ;
        RECT 69.340 116.775 70.415 116.945 ;
        RECT 68.675 116.175 69.045 116.635 ;
        RECT 69.340 116.435 69.510 116.775 ;
        RECT 69.680 116.175 70.010 116.605 ;
        RECT 70.245 116.435 70.415 116.775 ;
        RECT 70.585 116.675 70.755 117.455 ;
        RECT 70.925 117.235 71.095 117.825 ;
        RECT 71.265 117.425 71.615 118.045 ;
        RECT 70.925 116.845 71.390 117.235 ;
        RECT 71.785 116.975 71.955 118.335 ;
        RECT 72.125 117.145 72.585 118.195 ;
        RECT 71.560 116.805 71.955 116.975 ;
        RECT 71.560 116.675 71.730 116.805 ;
        RECT 70.585 116.345 71.265 116.675 ;
        RECT 71.480 116.345 71.730 116.675 ;
        RECT 71.900 116.175 72.150 116.635 ;
        RECT 72.320 116.360 72.645 117.145 ;
        RECT 72.815 116.345 72.985 118.465 ;
        RECT 73.155 118.345 73.485 118.725 ;
        RECT 73.655 118.175 73.910 118.465 ;
        RECT 74.395 118.255 74.565 118.725 ;
        RECT 73.160 118.005 73.910 118.175 ;
        RECT 74.735 118.075 75.065 118.555 ;
        RECT 75.235 118.255 75.405 118.725 ;
        RECT 75.575 118.075 75.905 118.555 ;
        RECT 73.160 117.015 73.390 118.005 ;
        RECT 74.140 117.905 75.905 118.075 ;
        RECT 76.075 117.915 76.245 118.725 ;
        RECT 76.445 118.345 77.515 118.515 ;
        RECT 76.445 117.990 76.765 118.345 ;
        RECT 73.560 117.185 73.910 117.835 ;
        RECT 74.140 117.355 74.550 117.905 ;
        RECT 76.440 117.735 76.765 117.990 ;
        RECT 74.735 117.525 76.765 117.735 ;
        RECT 76.420 117.515 76.765 117.525 ;
        RECT 76.935 117.775 77.175 118.175 ;
        RECT 77.345 118.115 77.515 118.345 ;
        RECT 77.685 118.285 77.875 118.725 ;
        RECT 78.045 118.275 78.995 118.555 ;
        RECT 79.215 118.365 79.565 118.535 ;
        RECT 77.345 117.945 77.875 118.115 ;
        RECT 74.140 117.185 75.865 117.355 ;
        RECT 73.160 116.845 73.910 117.015 ;
        RECT 73.155 116.175 73.485 116.675 ;
        RECT 73.655 116.345 73.910 116.845 ;
        RECT 74.395 116.175 74.565 117.015 ;
        RECT 74.775 116.345 75.025 117.185 ;
        RECT 75.235 116.175 75.405 117.015 ;
        RECT 75.575 116.345 75.865 117.185 ;
        RECT 76.075 116.175 76.245 117.235 ;
        RECT 76.420 116.895 76.590 117.515 ;
        RECT 76.935 117.405 77.475 117.775 ;
        RECT 77.655 117.665 77.875 117.945 ;
        RECT 78.045 117.495 78.215 118.275 ;
        RECT 77.810 117.325 78.215 117.495 ;
        RECT 78.385 117.485 78.735 118.105 ;
        RECT 77.810 117.235 77.980 117.325 ;
        RECT 78.905 117.315 79.115 118.105 ;
        RECT 76.760 117.065 77.980 117.235 ;
        RECT 78.440 117.155 79.115 117.315 ;
        RECT 76.420 116.725 77.220 116.895 ;
        RECT 76.540 116.175 76.870 116.555 ;
        RECT 77.050 116.435 77.220 116.725 ;
        RECT 77.810 116.685 77.980 117.065 ;
        RECT 78.150 117.145 79.115 117.155 ;
        RECT 79.305 117.975 79.565 118.365 ;
        RECT 79.775 118.265 80.105 118.725 ;
        RECT 80.980 118.335 81.835 118.505 ;
        RECT 82.040 118.335 82.535 118.505 ;
        RECT 82.705 118.365 83.035 118.725 ;
        RECT 79.305 117.285 79.475 117.975 ;
        RECT 79.645 117.625 79.815 117.805 ;
        RECT 79.985 117.795 80.775 118.045 ;
        RECT 80.980 117.625 81.150 118.335 ;
        RECT 81.320 117.825 81.675 118.045 ;
        RECT 79.645 117.455 81.335 117.625 ;
        RECT 78.150 116.855 78.610 117.145 ;
        RECT 79.305 117.115 80.805 117.285 ;
        RECT 79.305 116.975 79.475 117.115 ;
        RECT 78.915 116.805 79.475 116.975 ;
        RECT 77.390 116.175 77.640 116.635 ;
        RECT 77.810 116.345 78.680 116.685 ;
        RECT 78.915 116.345 79.085 116.805 ;
        RECT 79.920 116.775 80.995 116.945 ;
        RECT 79.255 116.175 79.625 116.635 ;
        RECT 79.920 116.435 80.090 116.775 ;
        RECT 80.260 116.175 80.590 116.605 ;
        RECT 80.825 116.435 80.995 116.775 ;
        RECT 81.165 116.675 81.335 117.455 ;
        RECT 81.505 117.235 81.675 117.825 ;
        RECT 81.845 117.425 82.195 118.045 ;
        RECT 81.505 116.845 81.970 117.235 ;
        RECT 82.365 116.975 82.535 118.335 ;
        RECT 82.705 117.145 83.165 118.195 ;
        RECT 82.140 116.805 82.535 116.975 ;
        RECT 82.140 116.675 82.310 116.805 ;
        RECT 81.165 116.345 81.845 116.675 ;
        RECT 82.060 116.345 82.310 116.675 ;
        RECT 82.480 116.175 82.730 116.635 ;
        RECT 82.900 116.360 83.225 117.145 ;
        RECT 83.395 116.345 83.565 118.465 ;
        RECT 83.735 118.345 84.065 118.725 ;
        RECT 84.235 118.175 84.490 118.465 ;
        RECT 83.740 118.005 84.490 118.175 ;
        RECT 85.215 118.175 85.385 118.555 ;
        RECT 85.565 118.345 85.895 118.725 ;
        RECT 85.215 118.005 85.880 118.175 ;
        RECT 86.075 118.050 86.335 118.555 ;
        RECT 83.740 117.015 83.970 118.005 ;
        RECT 84.140 117.185 84.490 117.835 ;
        RECT 85.145 117.455 85.475 117.825 ;
        RECT 85.710 117.750 85.880 118.005 ;
        RECT 85.710 117.420 85.995 117.750 ;
        RECT 85.710 117.275 85.880 117.420 ;
        RECT 85.215 117.105 85.880 117.275 ;
        RECT 86.165 117.250 86.335 118.050 ;
        RECT 86.565 117.905 86.775 118.725 ;
        RECT 86.945 117.925 87.275 118.555 ;
        RECT 86.945 117.325 87.195 117.925 ;
        RECT 87.445 117.905 87.675 118.725 ;
        RECT 88.805 118.000 89.095 118.725 ;
        RECT 89.575 118.255 89.745 118.725 ;
        RECT 89.915 118.075 90.245 118.555 ;
        RECT 90.415 118.255 90.585 118.725 ;
        RECT 90.755 118.075 91.085 118.555 ;
        RECT 89.320 117.905 91.085 118.075 ;
        RECT 91.255 117.915 91.425 118.725 ;
        RECT 91.625 118.345 92.695 118.515 ;
        RECT 91.625 117.990 91.945 118.345 ;
        RECT 87.365 117.485 87.695 117.735 ;
        RECT 89.320 117.355 89.730 117.905 ;
        RECT 91.620 117.735 91.945 117.990 ;
        RECT 89.915 117.525 91.945 117.735 ;
        RECT 91.600 117.515 91.945 117.525 ;
        RECT 92.115 117.775 92.355 118.175 ;
        RECT 92.525 118.115 92.695 118.345 ;
        RECT 92.865 118.285 93.055 118.725 ;
        RECT 93.225 118.275 94.175 118.555 ;
        RECT 94.395 118.365 94.745 118.535 ;
        RECT 92.525 117.945 93.055 118.115 ;
        RECT 83.740 116.845 84.490 117.015 ;
        RECT 83.735 116.175 84.065 116.675 ;
        RECT 84.235 116.345 84.490 116.845 ;
        RECT 85.215 116.345 85.385 117.105 ;
        RECT 85.565 116.175 85.895 116.935 ;
        RECT 86.065 116.345 86.335 117.250 ;
        RECT 86.565 116.175 86.775 117.315 ;
        RECT 86.945 116.345 87.275 117.325 ;
        RECT 87.445 116.175 87.675 117.315 ;
        RECT 88.805 116.175 89.095 117.340 ;
        RECT 89.320 117.185 91.045 117.355 ;
        RECT 89.575 116.175 89.745 117.015 ;
        RECT 89.955 116.345 90.205 117.185 ;
        RECT 90.415 116.175 90.585 117.015 ;
        RECT 90.755 116.345 91.045 117.185 ;
        RECT 91.255 116.175 91.425 117.235 ;
        RECT 91.600 116.895 91.770 117.515 ;
        RECT 92.115 117.405 92.655 117.775 ;
        RECT 92.835 117.665 93.055 117.945 ;
        RECT 93.225 117.495 93.395 118.275 ;
        RECT 92.990 117.325 93.395 117.495 ;
        RECT 93.565 117.485 93.915 118.105 ;
        RECT 92.990 117.235 93.160 117.325 ;
        RECT 94.085 117.315 94.295 118.105 ;
        RECT 91.940 117.065 93.160 117.235 ;
        RECT 93.620 117.155 94.295 117.315 ;
        RECT 91.600 116.725 92.400 116.895 ;
        RECT 91.720 116.175 92.050 116.555 ;
        RECT 92.230 116.435 92.400 116.725 ;
        RECT 92.990 116.685 93.160 117.065 ;
        RECT 93.330 117.145 94.295 117.155 ;
        RECT 94.485 117.975 94.745 118.365 ;
        RECT 94.955 118.265 95.285 118.725 ;
        RECT 96.160 118.335 97.015 118.505 ;
        RECT 97.220 118.335 97.715 118.505 ;
        RECT 97.885 118.365 98.215 118.725 ;
        RECT 94.485 117.285 94.655 117.975 ;
        RECT 94.825 117.625 94.995 117.805 ;
        RECT 95.165 117.795 95.955 118.045 ;
        RECT 96.160 117.625 96.330 118.335 ;
        RECT 96.500 117.825 96.855 118.045 ;
        RECT 94.825 117.455 96.515 117.625 ;
        RECT 93.330 116.855 93.790 117.145 ;
        RECT 94.485 117.115 95.985 117.285 ;
        RECT 94.485 116.975 94.655 117.115 ;
        RECT 94.095 116.805 94.655 116.975 ;
        RECT 92.570 116.175 92.820 116.635 ;
        RECT 92.990 116.345 93.860 116.685 ;
        RECT 94.095 116.345 94.265 116.805 ;
        RECT 95.100 116.775 96.175 116.945 ;
        RECT 94.435 116.175 94.805 116.635 ;
        RECT 95.100 116.435 95.270 116.775 ;
        RECT 95.440 116.175 95.770 116.605 ;
        RECT 96.005 116.435 96.175 116.775 ;
        RECT 96.345 116.675 96.515 117.455 ;
        RECT 96.685 117.235 96.855 117.825 ;
        RECT 97.025 117.425 97.375 118.045 ;
        RECT 96.685 116.845 97.150 117.235 ;
        RECT 97.545 116.975 97.715 118.335 ;
        RECT 97.885 117.145 98.345 118.195 ;
        RECT 97.320 116.805 97.715 116.975 ;
        RECT 97.320 116.675 97.490 116.805 ;
        RECT 96.345 116.345 97.025 116.675 ;
        RECT 97.240 116.345 97.490 116.675 ;
        RECT 97.660 116.175 97.910 116.635 ;
        RECT 98.080 116.360 98.405 117.145 ;
        RECT 98.575 116.345 98.745 118.465 ;
        RECT 98.915 118.345 99.245 118.725 ;
        RECT 99.415 118.175 99.670 118.465 ;
        RECT 100.155 118.255 100.325 118.725 ;
        RECT 98.920 118.005 99.670 118.175 ;
        RECT 100.495 118.075 100.825 118.555 ;
        RECT 100.995 118.255 101.165 118.725 ;
        RECT 101.335 118.075 101.665 118.555 ;
        RECT 98.920 117.015 99.150 118.005 ;
        RECT 99.900 117.905 101.665 118.075 ;
        RECT 101.835 117.915 102.005 118.725 ;
        RECT 102.205 118.345 103.275 118.515 ;
        RECT 102.205 117.990 102.525 118.345 ;
        RECT 99.320 117.185 99.670 117.835 ;
        RECT 99.900 117.355 100.310 117.905 ;
        RECT 102.200 117.735 102.525 117.990 ;
        RECT 100.495 117.525 102.525 117.735 ;
        RECT 102.180 117.515 102.525 117.525 ;
        RECT 102.695 117.775 102.935 118.175 ;
        RECT 103.105 118.115 103.275 118.345 ;
        RECT 103.445 118.285 103.635 118.725 ;
        RECT 103.805 118.275 104.755 118.555 ;
        RECT 104.975 118.365 105.325 118.535 ;
        RECT 103.105 117.945 103.635 118.115 ;
        RECT 99.900 117.185 101.625 117.355 ;
        RECT 98.920 116.845 99.670 117.015 ;
        RECT 98.915 116.175 99.245 116.675 ;
        RECT 99.415 116.345 99.670 116.845 ;
        RECT 100.155 116.175 100.325 117.015 ;
        RECT 100.535 116.345 100.785 117.185 ;
        RECT 100.995 116.175 101.165 117.015 ;
        RECT 101.335 116.345 101.625 117.185 ;
        RECT 101.835 116.175 102.005 117.235 ;
        RECT 102.180 116.895 102.350 117.515 ;
        RECT 102.695 117.405 103.235 117.775 ;
        RECT 103.415 117.665 103.635 117.945 ;
        RECT 103.805 117.495 103.975 118.275 ;
        RECT 103.570 117.325 103.975 117.495 ;
        RECT 104.145 117.485 104.495 118.105 ;
        RECT 103.570 117.235 103.740 117.325 ;
        RECT 104.665 117.315 104.875 118.105 ;
        RECT 102.520 117.065 103.740 117.235 ;
        RECT 104.200 117.155 104.875 117.315 ;
        RECT 102.180 116.725 102.980 116.895 ;
        RECT 102.300 116.175 102.630 116.555 ;
        RECT 102.810 116.435 102.980 116.725 ;
        RECT 103.570 116.685 103.740 117.065 ;
        RECT 103.910 117.145 104.875 117.155 ;
        RECT 105.065 117.975 105.325 118.365 ;
        RECT 105.535 118.265 105.865 118.725 ;
        RECT 106.740 118.335 107.595 118.505 ;
        RECT 107.800 118.335 108.295 118.505 ;
        RECT 108.465 118.365 108.795 118.725 ;
        RECT 105.065 117.285 105.235 117.975 ;
        RECT 105.405 117.625 105.575 117.805 ;
        RECT 105.745 117.795 106.535 118.045 ;
        RECT 106.740 117.625 106.910 118.335 ;
        RECT 107.080 117.825 107.435 118.045 ;
        RECT 105.405 117.455 107.095 117.625 ;
        RECT 103.910 116.855 104.370 117.145 ;
        RECT 105.065 117.115 106.565 117.285 ;
        RECT 105.065 116.975 105.235 117.115 ;
        RECT 104.675 116.805 105.235 116.975 ;
        RECT 103.150 116.175 103.400 116.635 ;
        RECT 103.570 116.345 104.440 116.685 ;
        RECT 104.675 116.345 104.845 116.805 ;
        RECT 105.680 116.775 106.755 116.945 ;
        RECT 105.015 116.175 105.385 116.635 ;
        RECT 105.680 116.435 105.850 116.775 ;
        RECT 106.020 116.175 106.350 116.605 ;
        RECT 106.585 116.435 106.755 116.775 ;
        RECT 106.925 116.675 107.095 117.455 ;
        RECT 107.265 117.235 107.435 117.825 ;
        RECT 107.605 117.425 107.955 118.045 ;
        RECT 107.265 116.845 107.730 117.235 ;
        RECT 108.125 116.975 108.295 118.335 ;
        RECT 108.465 117.145 108.925 118.195 ;
        RECT 107.900 116.805 108.295 116.975 ;
        RECT 107.900 116.675 108.070 116.805 ;
        RECT 106.925 116.345 107.605 116.675 ;
        RECT 107.820 116.345 108.070 116.675 ;
        RECT 108.240 116.175 108.490 116.635 ;
        RECT 108.660 116.360 108.985 117.145 ;
        RECT 109.155 116.345 109.325 118.465 ;
        RECT 109.495 118.345 109.825 118.725 ;
        RECT 109.995 118.175 110.250 118.465 ;
        RECT 109.500 118.005 110.250 118.175 ;
        RECT 109.500 117.015 109.730 118.005 ;
        RECT 110.485 117.905 110.695 118.725 ;
        RECT 110.865 117.925 111.195 118.555 ;
        RECT 109.900 117.185 110.250 117.835 ;
        RECT 110.865 117.325 111.115 117.925 ;
        RECT 111.365 117.905 111.595 118.725 ;
        RECT 111.865 117.905 112.075 118.725 ;
        RECT 112.245 117.925 112.575 118.555 ;
        RECT 111.285 117.485 111.615 117.735 ;
        RECT 112.245 117.325 112.495 117.925 ;
        RECT 112.745 117.905 112.975 118.725 ;
        RECT 113.185 117.975 114.395 118.725 ;
        RECT 114.565 118.000 114.855 118.725 ;
        RECT 115.335 118.255 115.505 118.725 ;
        RECT 115.675 118.075 116.005 118.555 ;
        RECT 116.175 118.255 116.345 118.725 ;
        RECT 116.515 118.075 116.845 118.555 ;
        RECT 112.665 117.485 112.995 117.735 ;
        RECT 109.500 116.845 110.250 117.015 ;
        RECT 109.495 116.175 109.825 116.675 ;
        RECT 109.995 116.345 110.250 116.845 ;
        RECT 110.485 116.175 110.695 117.315 ;
        RECT 110.865 116.345 111.195 117.325 ;
        RECT 111.365 116.175 111.595 117.315 ;
        RECT 111.865 116.175 112.075 117.315 ;
        RECT 112.245 116.345 112.575 117.325 ;
        RECT 112.745 116.175 112.975 117.315 ;
        RECT 113.185 117.265 113.705 117.805 ;
        RECT 113.875 117.435 114.395 117.975 ;
        RECT 115.080 117.905 116.845 118.075 ;
        RECT 117.015 117.915 117.185 118.725 ;
        RECT 117.385 118.345 118.455 118.515 ;
        RECT 117.385 117.990 117.705 118.345 ;
        RECT 115.080 117.355 115.490 117.905 ;
        RECT 117.380 117.735 117.705 117.990 ;
        RECT 115.675 117.525 117.705 117.735 ;
        RECT 117.360 117.515 117.705 117.525 ;
        RECT 117.875 117.775 118.115 118.175 ;
        RECT 118.285 118.115 118.455 118.345 ;
        RECT 118.625 118.285 118.815 118.725 ;
        RECT 118.985 118.275 119.935 118.555 ;
        RECT 120.155 118.365 120.505 118.535 ;
        RECT 118.285 117.945 118.815 118.115 ;
        RECT 113.185 116.175 114.395 117.265 ;
        RECT 114.565 116.175 114.855 117.340 ;
        RECT 115.080 117.185 116.805 117.355 ;
        RECT 115.335 116.175 115.505 117.015 ;
        RECT 115.715 116.345 115.965 117.185 ;
        RECT 116.175 116.175 116.345 117.015 ;
        RECT 116.515 116.345 116.805 117.185 ;
        RECT 117.015 116.175 117.185 117.235 ;
        RECT 117.360 116.895 117.530 117.515 ;
        RECT 117.875 117.405 118.415 117.775 ;
        RECT 118.595 117.665 118.815 117.945 ;
        RECT 118.985 117.495 119.155 118.275 ;
        RECT 118.750 117.325 119.155 117.495 ;
        RECT 119.325 117.485 119.675 118.105 ;
        RECT 118.750 117.235 118.920 117.325 ;
        RECT 119.845 117.315 120.055 118.105 ;
        RECT 117.700 117.065 118.920 117.235 ;
        RECT 119.380 117.155 120.055 117.315 ;
        RECT 117.360 116.725 118.160 116.895 ;
        RECT 117.480 116.175 117.810 116.555 ;
        RECT 117.990 116.435 118.160 116.725 ;
        RECT 118.750 116.685 118.920 117.065 ;
        RECT 119.090 117.145 120.055 117.155 ;
        RECT 120.245 117.975 120.505 118.365 ;
        RECT 120.715 118.265 121.045 118.725 ;
        RECT 121.920 118.335 122.775 118.505 ;
        RECT 122.980 118.335 123.475 118.505 ;
        RECT 123.645 118.365 123.975 118.725 ;
        RECT 120.245 117.285 120.415 117.975 ;
        RECT 120.585 117.625 120.755 117.805 ;
        RECT 120.925 117.795 121.715 118.045 ;
        RECT 121.920 117.625 122.090 118.335 ;
        RECT 122.260 117.825 122.615 118.045 ;
        RECT 120.585 117.455 122.275 117.625 ;
        RECT 119.090 116.855 119.550 117.145 ;
        RECT 120.245 117.115 121.745 117.285 ;
        RECT 120.245 116.975 120.415 117.115 ;
        RECT 119.855 116.805 120.415 116.975 ;
        RECT 118.330 116.175 118.580 116.635 ;
        RECT 118.750 116.345 119.620 116.685 ;
        RECT 119.855 116.345 120.025 116.805 ;
        RECT 120.860 116.775 121.935 116.945 ;
        RECT 120.195 116.175 120.565 116.635 ;
        RECT 120.860 116.435 121.030 116.775 ;
        RECT 121.200 116.175 121.530 116.605 ;
        RECT 121.765 116.435 121.935 116.775 ;
        RECT 122.105 116.675 122.275 117.455 ;
        RECT 122.445 117.235 122.615 117.825 ;
        RECT 122.785 117.425 123.135 118.045 ;
        RECT 122.445 116.845 122.910 117.235 ;
        RECT 123.305 116.975 123.475 118.335 ;
        RECT 123.645 117.145 124.105 118.195 ;
        RECT 123.080 116.805 123.475 116.975 ;
        RECT 123.080 116.675 123.250 116.805 ;
        RECT 122.105 116.345 122.785 116.675 ;
        RECT 123.000 116.345 123.250 116.675 ;
        RECT 123.420 116.175 123.670 116.635 ;
        RECT 123.840 116.360 124.165 117.145 ;
        RECT 124.335 116.345 124.505 118.465 ;
        RECT 124.675 118.345 125.005 118.725 ;
        RECT 125.175 118.175 125.430 118.465 ;
        RECT 124.680 118.005 125.430 118.175 ;
        RECT 124.680 117.015 124.910 118.005 ;
        RECT 126.525 117.975 127.735 118.725 ;
        RECT 125.080 117.185 125.430 117.835 ;
        RECT 126.525 117.265 127.045 117.805 ;
        RECT 127.215 117.435 127.735 117.975 ;
        RECT 124.680 116.845 125.430 117.015 ;
        RECT 124.675 116.175 125.005 116.675 ;
        RECT 125.175 116.345 125.430 116.845 ;
        RECT 126.525 116.175 127.735 117.265 ;
        RECT 29.840 116.005 127.820 116.175 ;
        RECT 29.925 114.915 31.135 116.005 ;
        RECT 31.770 115.570 37.115 116.005 ;
        RECT 29.925 114.205 30.445 114.745 ;
        RECT 30.615 114.375 31.135 114.915 ;
        RECT 33.360 114.320 33.710 115.570 ;
        RECT 37.285 114.840 37.575 116.005 ;
        RECT 38.515 115.165 38.685 116.005 ;
        RECT 38.895 114.995 39.145 115.835 ;
        RECT 39.355 115.165 39.525 116.005 ;
        RECT 39.695 114.995 39.985 115.835 ;
        RECT 29.925 113.455 31.135 114.205 ;
        RECT 35.190 114.000 35.530 114.830 ;
        RECT 38.260 114.825 39.985 114.995 ;
        RECT 40.195 114.945 40.365 116.005 ;
        RECT 40.660 115.625 40.990 116.005 ;
        RECT 41.170 115.455 41.340 115.745 ;
        RECT 41.510 115.545 41.760 116.005 ;
        RECT 40.540 115.285 41.340 115.455 ;
        RECT 41.930 115.495 42.800 115.835 ;
        RECT 38.260 114.275 38.670 114.825 ;
        RECT 40.540 114.665 40.710 115.285 ;
        RECT 41.930 115.115 42.100 115.495 ;
        RECT 43.035 115.375 43.205 115.835 ;
        RECT 43.375 115.545 43.745 116.005 ;
        RECT 44.040 115.405 44.210 115.745 ;
        RECT 44.380 115.575 44.710 116.005 ;
        RECT 44.945 115.405 45.115 115.745 ;
        RECT 40.880 114.945 42.100 115.115 ;
        RECT 42.270 115.035 42.730 115.325 ;
        RECT 43.035 115.205 43.595 115.375 ;
        RECT 44.040 115.235 45.115 115.405 ;
        RECT 45.285 115.505 45.965 115.835 ;
        RECT 46.180 115.505 46.430 115.835 ;
        RECT 46.600 115.545 46.850 116.005 ;
        RECT 43.425 115.065 43.595 115.205 ;
        RECT 42.270 115.025 43.235 115.035 ;
        RECT 41.930 114.855 42.100 114.945 ;
        RECT 42.560 114.865 43.235 115.025 ;
        RECT 40.540 114.655 40.885 114.665 ;
        RECT 38.855 114.445 40.885 114.655 ;
        RECT 31.770 113.455 37.115 114.000 ;
        RECT 37.285 113.455 37.575 114.180 ;
        RECT 38.260 114.105 40.025 114.275 ;
        RECT 38.515 113.455 38.685 113.925 ;
        RECT 38.855 113.625 39.185 114.105 ;
        RECT 39.355 113.455 39.525 113.925 ;
        RECT 39.695 113.625 40.025 114.105 ;
        RECT 40.195 113.455 40.365 114.265 ;
        RECT 40.560 114.190 40.885 114.445 ;
        RECT 40.565 113.835 40.885 114.190 ;
        RECT 41.055 114.405 41.595 114.775 ;
        RECT 41.930 114.685 42.335 114.855 ;
        RECT 41.055 114.005 41.295 114.405 ;
        RECT 41.775 114.235 41.995 114.515 ;
        RECT 41.465 114.065 41.995 114.235 ;
        RECT 41.465 113.835 41.635 114.065 ;
        RECT 42.165 113.905 42.335 114.685 ;
        RECT 42.505 114.075 42.855 114.695 ;
        RECT 43.025 114.075 43.235 114.865 ;
        RECT 43.425 114.895 44.925 115.065 ;
        RECT 43.425 114.205 43.595 114.895 ;
        RECT 45.285 114.725 45.455 115.505 ;
        RECT 46.260 115.375 46.430 115.505 ;
        RECT 43.765 114.555 45.455 114.725 ;
        RECT 45.625 114.945 46.090 115.335 ;
        RECT 46.260 115.205 46.655 115.375 ;
        RECT 43.765 114.375 43.935 114.555 ;
        RECT 40.565 113.665 41.635 113.835 ;
        RECT 41.805 113.455 41.995 113.895 ;
        RECT 42.165 113.625 43.115 113.905 ;
        RECT 43.425 113.815 43.685 114.205 ;
        RECT 44.105 114.135 44.895 114.385 ;
        RECT 43.335 113.645 43.685 113.815 ;
        RECT 43.895 113.455 44.225 113.915 ;
        RECT 45.100 113.845 45.270 114.555 ;
        RECT 45.625 114.355 45.795 114.945 ;
        RECT 45.440 114.135 45.795 114.355 ;
        RECT 45.965 114.135 46.315 114.755 ;
        RECT 46.485 113.845 46.655 115.205 ;
        RECT 47.020 115.035 47.345 115.820 ;
        RECT 46.825 113.985 47.285 115.035 ;
        RECT 45.100 113.675 45.955 113.845 ;
        RECT 46.160 113.675 46.655 113.845 ;
        RECT 46.825 113.455 47.155 113.815 ;
        RECT 47.515 113.715 47.685 115.835 ;
        RECT 47.855 115.505 48.185 116.005 ;
        RECT 48.355 115.335 48.610 115.835 ;
        RECT 47.860 115.165 48.610 115.335 ;
        RECT 47.860 114.175 48.090 115.165 ;
        RECT 48.260 114.345 48.610 114.995 ;
        RECT 48.785 114.915 49.995 116.005 ;
        RECT 48.785 114.375 49.305 114.915 ;
        RECT 50.165 114.840 50.455 116.005 ;
        RECT 50.625 114.915 51.835 116.005 ;
        RECT 52.010 115.570 57.355 116.005 ;
        RECT 49.475 114.205 49.995 114.745 ;
        RECT 50.625 114.375 51.145 114.915 ;
        RECT 51.315 114.205 51.835 114.745 ;
        RECT 53.600 114.320 53.950 115.570 ;
        RECT 57.585 114.865 57.795 116.005 ;
        RECT 57.965 114.855 58.295 115.835 ;
        RECT 58.465 114.865 58.695 116.005 ;
        RECT 58.905 114.915 61.495 116.005 ;
        RECT 47.860 114.005 48.610 114.175 ;
        RECT 47.855 113.455 48.185 113.835 ;
        RECT 48.355 113.715 48.610 114.005 ;
        RECT 48.785 113.455 49.995 114.205 ;
        RECT 50.165 113.455 50.455 114.180 ;
        RECT 50.625 113.455 51.835 114.205 ;
        RECT 55.430 114.000 55.770 114.830 ;
        RECT 52.010 113.455 57.355 114.000 ;
        RECT 57.585 113.455 57.795 114.275 ;
        RECT 57.965 114.255 58.215 114.855 ;
        RECT 58.385 114.445 58.715 114.695 ;
        RECT 58.905 114.395 60.115 114.915 ;
        RECT 61.705 114.865 61.935 116.005 ;
        RECT 62.105 114.855 62.435 115.835 ;
        RECT 62.605 114.865 62.815 116.005 ;
        RECT 57.965 113.625 58.295 114.255 ;
        RECT 58.465 113.455 58.695 114.275 ;
        RECT 60.285 114.225 61.495 114.745 ;
        RECT 61.685 114.445 62.015 114.695 ;
        RECT 58.905 113.455 61.495 114.225 ;
        RECT 61.705 113.455 61.935 114.275 ;
        RECT 62.185 114.255 62.435 114.855 ;
        RECT 63.045 114.840 63.335 116.005 ;
        RECT 64.005 114.865 64.235 116.005 ;
        RECT 64.405 114.855 64.735 115.835 ;
        RECT 64.905 114.865 65.115 116.005 ;
        RECT 65.655 115.165 65.825 116.005 ;
        RECT 66.035 114.995 66.285 115.835 ;
        RECT 66.495 115.165 66.665 116.005 ;
        RECT 66.835 114.995 67.125 115.835 ;
        RECT 63.985 114.445 64.315 114.695 ;
        RECT 62.105 113.625 62.435 114.255 ;
        RECT 62.605 113.455 62.815 114.275 ;
        RECT 63.045 113.455 63.335 114.180 ;
        RECT 64.005 113.455 64.235 114.275 ;
        RECT 64.485 114.255 64.735 114.855 ;
        RECT 65.400 114.825 67.125 114.995 ;
        RECT 67.335 114.945 67.505 116.005 ;
        RECT 67.800 115.625 68.130 116.005 ;
        RECT 68.310 115.455 68.480 115.745 ;
        RECT 68.650 115.545 68.900 116.005 ;
        RECT 67.680 115.285 68.480 115.455 ;
        RECT 69.070 115.495 69.940 115.835 ;
        RECT 65.400 114.275 65.810 114.825 ;
        RECT 67.680 114.665 67.850 115.285 ;
        RECT 69.070 115.115 69.240 115.495 ;
        RECT 70.175 115.375 70.345 115.835 ;
        RECT 70.515 115.545 70.885 116.005 ;
        RECT 71.180 115.405 71.350 115.745 ;
        RECT 71.520 115.575 71.850 116.005 ;
        RECT 72.085 115.405 72.255 115.745 ;
        RECT 68.020 114.945 69.240 115.115 ;
        RECT 69.410 115.035 69.870 115.325 ;
        RECT 70.175 115.205 70.735 115.375 ;
        RECT 71.180 115.235 72.255 115.405 ;
        RECT 72.425 115.505 73.105 115.835 ;
        RECT 73.320 115.505 73.570 115.835 ;
        RECT 73.740 115.545 73.990 116.005 ;
        RECT 70.565 115.065 70.735 115.205 ;
        RECT 69.410 115.025 70.375 115.035 ;
        RECT 69.070 114.855 69.240 114.945 ;
        RECT 69.700 114.865 70.375 115.025 ;
        RECT 67.680 114.655 68.025 114.665 ;
        RECT 65.995 114.445 68.025 114.655 ;
        RECT 64.405 113.625 64.735 114.255 ;
        RECT 64.905 113.455 65.115 114.275 ;
        RECT 65.400 114.105 67.165 114.275 ;
        RECT 65.655 113.455 65.825 113.925 ;
        RECT 65.995 113.625 66.325 114.105 ;
        RECT 66.495 113.455 66.665 113.925 ;
        RECT 66.835 113.625 67.165 114.105 ;
        RECT 67.335 113.455 67.505 114.265 ;
        RECT 67.700 114.190 68.025 114.445 ;
        RECT 67.705 113.835 68.025 114.190 ;
        RECT 68.195 114.405 68.735 114.775 ;
        RECT 69.070 114.685 69.475 114.855 ;
        RECT 68.195 114.005 68.435 114.405 ;
        RECT 68.915 114.235 69.135 114.515 ;
        RECT 68.605 114.065 69.135 114.235 ;
        RECT 68.605 113.835 68.775 114.065 ;
        RECT 69.305 113.905 69.475 114.685 ;
        RECT 69.645 114.075 69.995 114.695 ;
        RECT 70.165 114.075 70.375 114.865 ;
        RECT 70.565 114.895 72.065 115.065 ;
        RECT 70.565 114.205 70.735 114.895 ;
        RECT 72.425 114.725 72.595 115.505 ;
        RECT 73.400 115.375 73.570 115.505 ;
        RECT 70.905 114.555 72.595 114.725 ;
        RECT 72.765 114.945 73.230 115.335 ;
        RECT 73.400 115.205 73.795 115.375 ;
        RECT 70.905 114.375 71.075 114.555 ;
        RECT 67.705 113.665 68.775 113.835 ;
        RECT 68.945 113.455 69.135 113.895 ;
        RECT 69.305 113.625 70.255 113.905 ;
        RECT 70.565 113.815 70.825 114.205 ;
        RECT 71.245 114.135 72.035 114.385 ;
        RECT 70.475 113.645 70.825 113.815 ;
        RECT 71.035 113.455 71.365 113.915 ;
        RECT 72.240 113.845 72.410 114.555 ;
        RECT 72.765 114.355 72.935 114.945 ;
        RECT 72.580 114.135 72.935 114.355 ;
        RECT 73.105 114.135 73.455 114.755 ;
        RECT 73.625 113.845 73.795 115.205 ;
        RECT 74.160 115.035 74.485 115.820 ;
        RECT 73.965 113.985 74.425 115.035 ;
        RECT 72.240 113.675 73.095 113.845 ;
        RECT 73.300 113.675 73.795 113.845 ;
        RECT 73.965 113.455 74.295 113.815 ;
        RECT 74.655 113.715 74.825 115.835 ;
        RECT 74.995 115.505 75.325 116.005 ;
        RECT 75.495 115.335 75.750 115.835 ;
        RECT 75.000 115.165 75.750 115.335 ;
        RECT 75.000 114.175 75.230 115.165 ;
        RECT 75.400 114.345 75.750 114.995 ;
        RECT 75.925 114.840 76.215 116.005 ;
        RECT 76.390 115.570 81.735 116.005 ;
        RECT 81.910 115.570 87.255 116.005 ;
        RECT 77.980 114.320 78.330 115.570 ;
        RECT 75.000 114.005 75.750 114.175 ;
        RECT 74.995 113.455 75.325 113.835 ;
        RECT 75.495 113.715 75.750 114.005 ;
        RECT 75.925 113.455 76.215 114.180 ;
        RECT 79.810 114.000 80.150 114.830 ;
        RECT 83.500 114.320 83.850 115.570 ;
        RECT 87.465 114.865 87.695 116.005 ;
        RECT 87.865 114.855 88.195 115.835 ;
        RECT 88.365 114.865 88.575 116.005 ;
        RECT 85.330 114.000 85.670 114.830 ;
        RECT 87.445 114.445 87.775 114.695 ;
        RECT 76.390 113.455 81.735 114.000 ;
        RECT 81.910 113.455 87.255 114.000 ;
        RECT 87.465 113.455 87.695 114.275 ;
        RECT 87.945 114.255 88.195 114.855 ;
        RECT 88.805 114.840 89.095 116.005 ;
        RECT 89.575 115.165 89.745 116.005 ;
        RECT 89.955 114.995 90.205 115.835 ;
        RECT 90.415 115.165 90.585 116.005 ;
        RECT 90.755 114.995 91.045 115.835 ;
        RECT 89.320 114.825 91.045 114.995 ;
        RECT 91.255 114.945 91.425 116.005 ;
        RECT 91.720 115.625 92.050 116.005 ;
        RECT 92.230 115.455 92.400 115.745 ;
        RECT 92.570 115.545 92.820 116.005 ;
        RECT 91.600 115.285 92.400 115.455 ;
        RECT 92.990 115.495 93.860 115.835 ;
        RECT 89.320 114.275 89.730 114.825 ;
        RECT 91.600 114.665 91.770 115.285 ;
        RECT 92.990 115.115 93.160 115.495 ;
        RECT 94.095 115.375 94.265 115.835 ;
        RECT 94.435 115.545 94.805 116.005 ;
        RECT 95.100 115.405 95.270 115.745 ;
        RECT 95.440 115.575 95.770 116.005 ;
        RECT 96.005 115.405 96.175 115.745 ;
        RECT 91.940 114.945 93.160 115.115 ;
        RECT 93.330 115.035 93.790 115.325 ;
        RECT 94.095 115.205 94.655 115.375 ;
        RECT 95.100 115.235 96.175 115.405 ;
        RECT 96.345 115.505 97.025 115.835 ;
        RECT 97.240 115.505 97.490 115.835 ;
        RECT 97.660 115.545 97.910 116.005 ;
        RECT 94.485 115.065 94.655 115.205 ;
        RECT 93.330 115.025 94.295 115.035 ;
        RECT 92.990 114.855 93.160 114.945 ;
        RECT 93.620 114.865 94.295 115.025 ;
        RECT 91.600 114.655 91.945 114.665 ;
        RECT 89.915 114.445 91.945 114.655 ;
        RECT 87.865 113.625 88.195 114.255 ;
        RECT 88.365 113.455 88.575 114.275 ;
        RECT 88.805 113.455 89.095 114.180 ;
        RECT 89.320 114.105 91.085 114.275 ;
        RECT 89.575 113.455 89.745 113.925 ;
        RECT 89.915 113.625 90.245 114.105 ;
        RECT 90.415 113.455 90.585 113.925 ;
        RECT 90.755 113.625 91.085 114.105 ;
        RECT 91.255 113.455 91.425 114.265 ;
        RECT 91.620 114.190 91.945 114.445 ;
        RECT 91.625 113.835 91.945 114.190 ;
        RECT 92.115 114.405 92.655 114.775 ;
        RECT 92.990 114.685 93.395 114.855 ;
        RECT 92.115 114.005 92.355 114.405 ;
        RECT 92.835 114.235 93.055 114.515 ;
        RECT 92.525 114.065 93.055 114.235 ;
        RECT 92.525 113.835 92.695 114.065 ;
        RECT 93.225 113.905 93.395 114.685 ;
        RECT 93.565 114.075 93.915 114.695 ;
        RECT 94.085 114.075 94.295 114.865 ;
        RECT 94.485 114.895 95.985 115.065 ;
        RECT 94.485 114.205 94.655 114.895 ;
        RECT 96.345 114.725 96.515 115.505 ;
        RECT 97.320 115.375 97.490 115.505 ;
        RECT 94.825 114.555 96.515 114.725 ;
        RECT 96.685 114.945 97.150 115.335 ;
        RECT 97.320 115.205 97.715 115.375 ;
        RECT 94.825 114.375 94.995 114.555 ;
        RECT 91.625 113.665 92.695 113.835 ;
        RECT 92.865 113.455 93.055 113.895 ;
        RECT 93.225 113.625 94.175 113.905 ;
        RECT 94.485 113.815 94.745 114.205 ;
        RECT 95.165 114.135 95.955 114.385 ;
        RECT 94.395 113.645 94.745 113.815 ;
        RECT 94.955 113.455 95.285 113.915 ;
        RECT 96.160 113.845 96.330 114.555 ;
        RECT 96.685 114.355 96.855 114.945 ;
        RECT 96.500 114.135 96.855 114.355 ;
        RECT 97.025 114.135 97.375 114.755 ;
        RECT 97.545 113.845 97.715 115.205 ;
        RECT 98.080 115.035 98.405 115.820 ;
        RECT 97.885 113.985 98.345 115.035 ;
        RECT 96.160 113.675 97.015 113.845 ;
        RECT 97.220 113.675 97.715 113.845 ;
        RECT 97.885 113.455 98.215 113.815 ;
        RECT 98.575 113.715 98.745 115.835 ;
        RECT 98.915 115.505 99.245 116.005 ;
        RECT 99.415 115.335 99.670 115.835 ;
        RECT 98.920 115.165 99.670 115.335 ;
        RECT 98.920 114.175 99.150 115.165 ;
        RECT 99.320 114.345 99.670 114.995 ;
        RECT 99.905 114.865 100.115 116.005 ;
        RECT 100.285 114.855 100.615 115.835 ;
        RECT 100.785 114.865 101.015 116.005 ;
        RECT 98.920 114.005 99.670 114.175 ;
        RECT 98.915 113.455 99.245 113.835 ;
        RECT 99.415 113.715 99.670 114.005 ;
        RECT 99.905 113.455 100.115 114.275 ;
        RECT 100.285 114.255 100.535 114.855 ;
        RECT 101.685 114.840 101.975 116.005 ;
        RECT 102.645 114.865 102.875 116.005 ;
        RECT 103.045 114.855 103.375 115.835 ;
        RECT 103.545 114.865 103.755 116.005 ;
        RECT 104.295 115.165 104.465 116.005 ;
        RECT 104.675 114.995 104.925 115.835 ;
        RECT 105.135 115.165 105.305 116.005 ;
        RECT 105.475 114.995 105.765 115.835 ;
        RECT 100.705 114.445 101.035 114.695 ;
        RECT 102.625 114.445 102.955 114.695 ;
        RECT 100.285 113.625 100.615 114.255 ;
        RECT 100.785 113.455 101.015 114.275 ;
        RECT 101.685 113.455 101.975 114.180 ;
        RECT 102.645 113.455 102.875 114.275 ;
        RECT 103.125 114.255 103.375 114.855 ;
        RECT 104.040 114.825 105.765 114.995 ;
        RECT 105.975 114.945 106.145 116.005 ;
        RECT 106.440 115.625 106.770 116.005 ;
        RECT 106.950 115.455 107.120 115.745 ;
        RECT 107.290 115.545 107.540 116.005 ;
        RECT 106.320 115.285 107.120 115.455 ;
        RECT 107.710 115.495 108.580 115.835 ;
        RECT 104.040 114.275 104.450 114.825 ;
        RECT 106.320 114.665 106.490 115.285 ;
        RECT 107.710 115.115 107.880 115.495 ;
        RECT 108.815 115.375 108.985 115.835 ;
        RECT 109.155 115.545 109.525 116.005 ;
        RECT 109.820 115.405 109.990 115.745 ;
        RECT 110.160 115.575 110.490 116.005 ;
        RECT 110.725 115.405 110.895 115.745 ;
        RECT 106.660 114.945 107.880 115.115 ;
        RECT 108.050 115.035 108.510 115.325 ;
        RECT 108.815 115.205 109.375 115.375 ;
        RECT 109.820 115.235 110.895 115.405 ;
        RECT 111.065 115.505 111.745 115.835 ;
        RECT 111.960 115.505 112.210 115.835 ;
        RECT 112.380 115.545 112.630 116.005 ;
        RECT 109.205 115.065 109.375 115.205 ;
        RECT 108.050 115.025 109.015 115.035 ;
        RECT 107.710 114.855 107.880 114.945 ;
        RECT 108.340 114.865 109.015 115.025 ;
        RECT 106.320 114.655 106.665 114.665 ;
        RECT 104.635 114.445 106.665 114.655 ;
        RECT 103.045 113.625 103.375 114.255 ;
        RECT 103.545 113.455 103.755 114.275 ;
        RECT 104.040 114.105 105.805 114.275 ;
        RECT 104.295 113.455 104.465 113.925 ;
        RECT 104.635 113.625 104.965 114.105 ;
        RECT 105.135 113.455 105.305 113.925 ;
        RECT 105.475 113.625 105.805 114.105 ;
        RECT 105.975 113.455 106.145 114.265 ;
        RECT 106.340 114.190 106.665 114.445 ;
        RECT 106.345 113.835 106.665 114.190 ;
        RECT 106.835 114.405 107.375 114.775 ;
        RECT 107.710 114.685 108.115 114.855 ;
        RECT 106.835 114.005 107.075 114.405 ;
        RECT 107.555 114.235 107.775 114.515 ;
        RECT 107.245 114.065 107.775 114.235 ;
        RECT 107.245 113.835 107.415 114.065 ;
        RECT 107.945 113.905 108.115 114.685 ;
        RECT 108.285 114.075 108.635 114.695 ;
        RECT 108.805 114.075 109.015 114.865 ;
        RECT 109.205 114.895 110.705 115.065 ;
        RECT 109.205 114.205 109.375 114.895 ;
        RECT 111.065 114.725 111.235 115.505 ;
        RECT 112.040 115.375 112.210 115.505 ;
        RECT 109.545 114.555 111.235 114.725 ;
        RECT 111.405 114.945 111.870 115.335 ;
        RECT 112.040 115.205 112.435 115.375 ;
        RECT 109.545 114.375 109.715 114.555 ;
        RECT 106.345 113.665 107.415 113.835 ;
        RECT 107.585 113.455 107.775 113.895 ;
        RECT 107.945 113.625 108.895 113.905 ;
        RECT 109.205 113.815 109.465 114.205 ;
        RECT 109.885 114.135 110.675 114.385 ;
        RECT 109.115 113.645 109.465 113.815 ;
        RECT 109.675 113.455 110.005 113.915 ;
        RECT 110.880 113.845 111.050 114.555 ;
        RECT 111.405 114.355 111.575 114.945 ;
        RECT 111.220 114.135 111.575 114.355 ;
        RECT 111.745 114.135 112.095 114.755 ;
        RECT 112.265 113.845 112.435 115.205 ;
        RECT 112.800 115.035 113.125 115.820 ;
        RECT 112.605 113.985 113.065 115.035 ;
        RECT 110.880 113.675 111.735 113.845 ;
        RECT 111.940 113.675 112.435 113.845 ;
        RECT 112.605 113.455 112.935 113.815 ;
        RECT 113.295 113.715 113.465 115.835 ;
        RECT 113.635 115.505 113.965 116.005 ;
        RECT 114.135 115.335 114.390 115.835 ;
        RECT 113.640 115.165 114.390 115.335 ;
        RECT 113.640 114.175 113.870 115.165 ;
        RECT 114.040 114.345 114.390 114.995 ;
        RECT 114.565 114.840 114.855 116.005 ;
        RECT 115.025 114.915 117.615 116.005 ;
        RECT 115.025 114.395 116.235 114.915 ;
        RECT 117.825 114.865 118.055 116.005 ;
        RECT 118.225 114.855 118.555 115.835 ;
        RECT 118.725 114.865 118.935 116.005 ;
        RECT 120.145 114.865 120.355 116.005 ;
        RECT 116.405 114.225 117.615 114.745 ;
        RECT 117.805 114.445 118.135 114.695 ;
        RECT 113.640 114.005 114.390 114.175 ;
        RECT 113.635 113.455 113.965 113.835 ;
        RECT 114.135 113.715 114.390 114.005 ;
        RECT 114.565 113.455 114.855 114.180 ;
        RECT 115.025 113.455 117.615 114.225 ;
        RECT 117.825 113.455 118.055 114.275 ;
        RECT 118.305 114.255 118.555 114.855 ;
        RECT 120.525 114.855 120.855 115.835 ;
        RECT 121.025 114.865 121.255 116.005 ;
        RECT 121.465 114.915 124.975 116.005 ;
        RECT 125.145 114.930 125.415 115.835 ;
        RECT 125.585 115.245 125.915 116.005 ;
        RECT 126.095 115.075 126.275 115.835 ;
        RECT 118.225 113.625 118.555 114.255 ;
        RECT 118.725 113.455 118.935 114.275 ;
        RECT 120.145 113.455 120.355 114.275 ;
        RECT 120.525 114.255 120.775 114.855 ;
        RECT 120.945 114.445 121.275 114.695 ;
        RECT 121.465 114.395 123.155 114.915 ;
        RECT 120.525 113.625 120.855 114.255 ;
        RECT 121.025 113.455 121.255 114.275 ;
        RECT 123.325 114.225 124.975 114.745 ;
        RECT 121.465 113.455 124.975 114.225 ;
        RECT 125.145 114.130 125.325 114.930 ;
        RECT 125.600 114.905 126.275 115.075 ;
        RECT 126.525 114.915 127.735 116.005 ;
        RECT 125.600 114.760 125.770 114.905 ;
        RECT 125.495 114.430 125.770 114.760 ;
        RECT 125.600 114.175 125.770 114.430 ;
        RECT 125.995 114.355 126.335 114.725 ;
        RECT 126.525 114.375 127.045 114.915 ;
        RECT 127.215 114.205 127.735 114.745 ;
        RECT 125.145 113.625 125.405 114.130 ;
        RECT 125.600 114.005 126.265 114.175 ;
        RECT 125.585 113.455 125.915 113.835 ;
        RECT 126.095 113.625 126.265 114.005 ;
        RECT 126.525 113.455 127.735 114.205 ;
        RECT 29.840 113.285 127.820 113.455 ;
        RECT 19.165 66.070 30.165 66.940 ;
        RECT 19.165 54.930 20.835 66.070 ;
        RECT 21.465 65.555 26.465 65.725 ;
        RECT 21.235 55.300 21.405 65.340 ;
        RECT 26.525 55.300 26.695 65.340 ;
        RECT 27.095 54.930 27.265 66.070 ;
        RECT 27.895 65.555 28.895 65.725 ;
        RECT 27.665 55.300 27.835 65.340 ;
        RECT 28.955 55.300 29.125 65.340 ;
        RECT 29.525 54.930 30.165 66.070 ;
        RECT 19.165 52.860 30.165 54.930 ;
        RECT 19.165 49.370 21.005 52.860 ;
        RECT 22.765 52.780 30.165 52.860 ;
        RECT 21.635 52.350 22.135 52.520 ;
        RECT 21.405 50.095 21.575 52.135 ;
        RECT 22.195 50.095 22.365 52.135 ;
        RECT 21.635 49.710 22.135 49.880 ;
        RECT 22.765 49.370 25.085 52.780 ;
        RECT 25.715 52.270 26.215 52.440 ;
        RECT 19.165 48.650 25.085 49.370 ;
        RECT 19.135 48.040 23.045 48.260 ;
        RECT 19.135 45.640 20.855 48.040 ;
        RECT 21.485 47.530 21.985 47.700 ;
        RECT 21.255 46.320 21.425 47.360 ;
        RECT 22.045 46.320 22.215 47.360 ;
        RECT 21.485 45.980 21.985 46.150 ;
        RECT 22.615 45.640 23.045 48.040 ;
        RECT 24.025 46.290 25.085 48.650 ;
        RECT 25.485 47.015 25.655 52.055 ;
        RECT 26.275 47.015 26.445 52.055 ;
        RECT 25.715 46.630 26.215 46.800 ;
        RECT 26.845 46.290 27.015 52.780 ;
        RECT 27.645 52.270 28.145 52.440 ;
        RECT 27.415 47.015 27.585 52.055 ;
        RECT 28.205 47.015 28.375 52.055 ;
        RECT 27.645 46.630 28.145 46.800 ;
        RECT 28.775 46.290 30.165 52.780 ;
        RECT 30.365 66.080 41.365 66.950 ;
        RECT 30.365 54.940 32.035 66.080 ;
        RECT 32.665 65.565 37.665 65.735 ;
        RECT 32.435 55.310 32.605 65.350 ;
        RECT 37.725 55.310 37.895 65.350 ;
        RECT 38.295 54.940 38.465 66.080 ;
        RECT 39.095 65.565 40.095 65.735 ;
        RECT 38.865 55.310 39.035 65.350 ;
        RECT 40.155 55.310 40.325 65.350 ;
        RECT 40.725 54.940 41.365 66.080 ;
        RECT 30.365 52.870 41.365 54.940 ;
        RECT 30.365 49.380 32.205 52.870 ;
        RECT 33.965 52.790 41.365 52.870 ;
        RECT 32.835 52.360 33.335 52.530 ;
        RECT 32.605 50.105 32.775 52.145 ;
        RECT 33.395 50.105 33.565 52.145 ;
        RECT 32.835 49.720 33.335 49.890 ;
        RECT 33.965 49.380 36.285 52.790 ;
        RECT 36.915 52.280 37.415 52.450 ;
        RECT 30.365 48.660 36.285 49.380 ;
        RECT 24.025 45.800 30.165 46.290 ;
        RECT 30.335 48.050 34.245 48.270 ;
        RECT 19.135 45.370 23.045 45.640 ;
        RECT 30.335 45.650 32.055 48.050 ;
        RECT 32.685 47.540 33.185 47.710 ;
        RECT 32.455 46.330 32.625 47.370 ;
        RECT 33.245 46.330 33.415 47.370 ;
        RECT 32.685 45.990 33.185 46.160 ;
        RECT 33.815 45.650 34.245 48.050 ;
        RECT 35.225 46.300 36.285 48.660 ;
        RECT 36.685 47.025 36.855 52.065 ;
        RECT 37.475 47.025 37.645 52.065 ;
        RECT 36.915 46.640 37.415 46.810 ;
        RECT 38.045 46.300 38.215 52.790 ;
        RECT 38.845 52.280 39.345 52.450 ;
        RECT 38.615 47.025 38.785 52.065 ;
        RECT 39.405 47.025 39.575 52.065 ;
        RECT 38.845 46.640 39.345 46.810 ;
        RECT 39.975 46.300 41.365 52.790 ;
        RECT 41.585 66.050 52.585 66.920 ;
        RECT 41.585 54.910 43.255 66.050 ;
        RECT 43.885 65.535 48.885 65.705 ;
        RECT 43.655 55.280 43.825 65.320 ;
        RECT 48.945 55.280 49.115 65.320 ;
        RECT 49.515 54.910 49.685 66.050 ;
        RECT 50.315 65.535 51.315 65.705 ;
        RECT 50.085 55.280 50.255 65.320 ;
        RECT 51.375 55.280 51.545 65.320 ;
        RECT 51.945 54.910 52.585 66.050 ;
        RECT 41.585 52.840 52.585 54.910 ;
        RECT 41.585 49.350 43.425 52.840 ;
        RECT 45.185 52.760 52.585 52.840 ;
        RECT 44.055 52.330 44.555 52.500 ;
        RECT 43.825 50.075 43.995 52.115 ;
        RECT 44.615 50.075 44.785 52.115 ;
        RECT 44.055 49.690 44.555 49.860 ;
        RECT 45.185 49.350 47.505 52.760 ;
        RECT 48.135 52.250 48.635 52.420 ;
        RECT 41.585 48.630 47.505 49.350 ;
        RECT 35.225 45.810 41.365 46.300 ;
        RECT 41.555 48.020 45.465 48.240 ;
        RECT 30.335 45.380 34.245 45.650 ;
        RECT 41.555 45.620 43.275 48.020 ;
        RECT 43.905 47.510 44.405 47.680 ;
        RECT 43.675 46.300 43.845 47.340 ;
        RECT 44.465 46.300 44.635 47.340 ;
        RECT 43.905 45.960 44.405 46.130 ;
        RECT 45.035 45.620 45.465 48.020 ;
        RECT 46.445 46.270 47.505 48.630 ;
        RECT 47.905 46.995 48.075 52.035 ;
        RECT 48.695 46.995 48.865 52.035 ;
        RECT 48.135 46.610 48.635 46.780 ;
        RECT 49.265 46.270 49.435 52.760 ;
        RECT 50.065 52.250 50.565 52.420 ;
        RECT 49.835 46.995 50.005 52.035 ;
        RECT 50.625 46.995 50.795 52.035 ;
        RECT 50.065 46.610 50.565 46.780 ;
        RECT 51.195 46.270 52.585 52.760 ;
        RECT 52.835 66.030 63.835 66.900 ;
        RECT 52.835 54.890 54.505 66.030 ;
        RECT 55.135 65.515 60.135 65.685 ;
        RECT 54.905 55.260 55.075 65.300 ;
        RECT 60.195 55.260 60.365 65.300 ;
        RECT 60.765 54.890 60.935 66.030 ;
        RECT 61.565 65.515 62.565 65.685 ;
        RECT 61.335 55.260 61.505 65.300 ;
        RECT 62.625 55.260 62.795 65.300 ;
        RECT 63.195 54.890 63.835 66.030 ;
        RECT 52.835 52.820 63.835 54.890 ;
        RECT 52.835 49.330 54.675 52.820 ;
        RECT 56.435 52.740 63.835 52.820 ;
        RECT 55.305 52.310 55.805 52.480 ;
        RECT 55.075 50.055 55.245 52.095 ;
        RECT 55.865 50.055 56.035 52.095 ;
        RECT 55.305 49.670 55.805 49.840 ;
        RECT 56.435 49.330 58.755 52.740 ;
        RECT 59.385 52.230 59.885 52.400 ;
        RECT 52.835 48.610 58.755 49.330 ;
        RECT 46.445 45.780 52.585 46.270 ;
        RECT 52.805 48.000 56.715 48.220 ;
        RECT 41.555 45.350 45.465 45.620 ;
        RECT 52.805 45.600 54.525 48.000 ;
        RECT 55.155 47.490 55.655 47.660 ;
        RECT 54.925 46.280 55.095 47.320 ;
        RECT 55.715 46.280 55.885 47.320 ;
        RECT 55.155 45.940 55.655 46.110 ;
        RECT 56.285 45.600 56.715 48.000 ;
        RECT 57.695 46.250 58.755 48.610 ;
        RECT 59.155 46.975 59.325 52.015 ;
        RECT 59.945 46.975 60.115 52.015 ;
        RECT 59.385 46.590 59.885 46.760 ;
        RECT 60.515 46.250 60.685 52.740 ;
        RECT 61.315 52.230 61.815 52.400 ;
        RECT 61.085 46.975 61.255 52.015 ;
        RECT 61.875 46.975 62.045 52.015 ;
        RECT 61.315 46.590 61.815 46.760 ;
        RECT 62.445 46.250 63.835 52.740 ;
        RECT 64.055 66.020 75.055 66.890 ;
        RECT 64.055 54.880 65.725 66.020 ;
        RECT 66.355 65.505 71.355 65.675 ;
        RECT 66.125 55.250 66.295 65.290 ;
        RECT 71.415 55.250 71.585 65.290 ;
        RECT 71.985 54.880 72.155 66.020 ;
        RECT 72.785 65.505 73.785 65.675 ;
        RECT 72.555 55.250 72.725 65.290 ;
        RECT 73.845 55.250 74.015 65.290 ;
        RECT 74.415 54.880 75.055 66.020 ;
        RECT 64.055 52.810 75.055 54.880 ;
        RECT 64.055 49.320 65.895 52.810 ;
        RECT 67.655 52.730 75.055 52.810 ;
        RECT 66.525 52.300 67.025 52.470 ;
        RECT 66.295 50.045 66.465 52.085 ;
        RECT 67.085 50.045 67.255 52.085 ;
        RECT 66.525 49.660 67.025 49.830 ;
        RECT 67.655 49.320 69.975 52.730 ;
        RECT 70.605 52.220 71.105 52.390 ;
        RECT 64.055 48.600 69.975 49.320 ;
        RECT 57.695 45.760 63.835 46.250 ;
        RECT 64.025 47.990 67.935 48.210 ;
        RECT 52.805 45.330 56.715 45.600 ;
        RECT 64.025 45.590 65.745 47.990 ;
        RECT 66.375 47.480 66.875 47.650 ;
        RECT 66.145 46.270 66.315 47.310 ;
        RECT 66.935 46.270 67.105 47.310 ;
        RECT 66.375 45.930 66.875 46.100 ;
        RECT 67.505 45.590 67.935 47.990 ;
        RECT 68.915 46.240 69.975 48.600 ;
        RECT 70.375 46.965 70.545 52.005 ;
        RECT 71.165 46.965 71.335 52.005 ;
        RECT 70.605 46.580 71.105 46.750 ;
        RECT 71.735 46.240 71.905 52.730 ;
        RECT 72.535 52.220 73.035 52.390 ;
        RECT 72.305 46.965 72.475 52.005 ;
        RECT 73.095 46.965 73.265 52.005 ;
        RECT 72.535 46.580 73.035 46.750 ;
        RECT 73.665 46.240 75.055 52.730 ;
        RECT 75.295 66.010 86.295 66.880 ;
        RECT 75.295 54.870 76.965 66.010 ;
        RECT 77.595 65.495 82.595 65.665 ;
        RECT 77.365 55.240 77.535 65.280 ;
        RECT 82.655 55.240 82.825 65.280 ;
        RECT 83.225 54.870 83.395 66.010 ;
        RECT 84.025 65.495 85.025 65.665 ;
        RECT 83.795 55.240 83.965 65.280 ;
        RECT 85.085 55.240 85.255 65.280 ;
        RECT 85.655 54.870 86.295 66.010 ;
        RECT 75.295 52.800 86.295 54.870 ;
        RECT 75.295 49.310 77.135 52.800 ;
        RECT 78.895 52.720 86.295 52.800 ;
        RECT 77.765 52.290 78.265 52.460 ;
        RECT 77.535 50.035 77.705 52.075 ;
        RECT 78.325 50.035 78.495 52.075 ;
        RECT 77.765 49.650 78.265 49.820 ;
        RECT 78.895 49.310 81.215 52.720 ;
        RECT 81.845 52.210 82.345 52.380 ;
        RECT 75.295 48.590 81.215 49.310 ;
        RECT 68.915 45.750 75.055 46.240 ;
        RECT 75.265 47.980 79.175 48.200 ;
        RECT 64.025 45.320 67.935 45.590 ;
        RECT 75.265 45.580 76.985 47.980 ;
        RECT 77.615 47.470 78.115 47.640 ;
        RECT 77.385 46.260 77.555 47.300 ;
        RECT 78.175 46.260 78.345 47.300 ;
        RECT 77.615 45.920 78.115 46.090 ;
        RECT 78.745 45.580 79.175 47.980 ;
        RECT 80.155 46.230 81.215 48.590 ;
        RECT 81.615 46.955 81.785 51.995 ;
        RECT 82.405 46.955 82.575 51.995 ;
        RECT 81.845 46.570 82.345 46.740 ;
        RECT 82.975 46.230 83.145 52.720 ;
        RECT 83.775 52.210 84.275 52.380 ;
        RECT 83.545 46.955 83.715 51.995 ;
        RECT 84.335 46.955 84.505 51.995 ;
        RECT 83.775 46.570 84.275 46.740 ;
        RECT 84.905 46.230 86.295 52.720 ;
        RECT 86.545 66.020 97.545 66.890 ;
        RECT 131.125 66.880 140.025 66.890 ;
        RECT 86.545 54.880 88.215 66.020 ;
        RECT 88.845 65.505 93.845 65.675 ;
        RECT 88.615 55.250 88.785 65.290 ;
        RECT 93.905 55.250 94.075 65.290 ;
        RECT 94.475 54.880 94.645 66.020 ;
        RECT 95.275 65.505 96.275 65.675 ;
        RECT 95.045 55.250 95.215 65.290 ;
        RECT 96.335 55.250 96.505 65.290 ;
        RECT 96.905 54.880 97.545 66.020 ;
        RECT 86.545 52.810 97.545 54.880 ;
        RECT 86.545 49.320 88.385 52.810 ;
        RECT 90.145 52.730 97.545 52.810 ;
        RECT 89.015 52.300 89.515 52.470 ;
        RECT 88.785 50.045 88.955 52.085 ;
        RECT 89.575 50.045 89.745 52.085 ;
        RECT 89.015 49.660 89.515 49.830 ;
        RECT 90.145 49.320 92.465 52.730 ;
        RECT 93.095 52.220 93.595 52.390 ;
        RECT 86.545 48.600 92.465 49.320 ;
        RECT 80.155 45.740 86.295 46.230 ;
        RECT 86.515 47.990 90.425 48.210 ;
        RECT 75.265 45.310 79.175 45.580 ;
        RECT 86.515 45.590 88.235 47.990 ;
        RECT 88.865 47.480 89.365 47.650 ;
        RECT 88.635 46.270 88.805 47.310 ;
        RECT 89.425 46.270 89.595 47.310 ;
        RECT 88.865 45.930 89.365 46.100 ;
        RECT 89.995 45.590 90.425 47.990 ;
        RECT 91.405 46.240 92.465 48.600 ;
        RECT 92.865 46.965 93.035 52.005 ;
        RECT 93.655 46.965 93.825 52.005 ;
        RECT 93.095 46.580 93.595 46.750 ;
        RECT 94.225 46.240 94.395 52.730 ;
        RECT 95.025 52.220 95.525 52.390 ;
        RECT 94.795 46.965 94.965 52.005 ;
        RECT 95.585 46.965 95.755 52.005 ;
        RECT 95.025 46.580 95.525 46.750 ;
        RECT 96.155 46.240 97.545 52.730 ;
        RECT 97.825 66.010 108.825 66.880 ;
        RECT 97.825 54.870 99.495 66.010 ;
        RECT 100.125 65.495 105.125 65.665 ;
        RECT 99.895 55.240 100.065 65.280 ;
        RECT 105.185 55.240 105.355 65.280 ;
        RECT 105.755 54.870 105.925 66.010 ;
        RECT 106.555 65.495 107.555 65.665 ;
        RECT 106.325 55.240 106.495 65.280 ;
        RECT 107.615 55.240 107.785 65.280 ;
        RECT 108.185 54.870 108.825 66.010 ;
        RECT 97.825 52.800 108.825 54.870 ;
        RECT 97.825 49.310 99.665 52.800 ;
        RECT 101.425 52.720 108.825 52.800 ;
        RECT 100.295 52.290 100.795 52.460 ;
        RECT 100.065 50.035 100.235 52.075 ;
        RECT 100.855 50.035 101.025 52.075 ;
        RECT 100.295 49.650 100.795 49.820 ;
        RECT 101.425 49.310 103.745 52.720 ;
        RECT 104.375 52.210 104.875 52.380 ;
        RECT 97.825 48.590 103.745 49.310 ;
        RECT 91.405 45.750 97.545 46.240 ;
        RECT 97.795 47.980 101.705 48.200 ;
        RECT 86.515 45.320 90.425 45.590 ;
        RECT 97.795 45.580 99.515 47.980 ;
        RECT 100.145 47.470 100.645 47.640 ;
        RECT 99.915 46.260 100.085 47.300 ;
        RECT 100.705 46.260 100.875 47.300 ;
        RECT 100.145 45.920 100.645 46.090 ;
        RECT 101.275 45.580 101.705 47.980 ;
        RECT 102.685 46.230 103.745 48.590 ;
        RECT 104.145 46.955 104.315 51.995 ;
        RECT 104.935 46.955 105.105 51.995 ;
        RECT 104.375 46.570 104.875 46.740 ;
        RECT 105.505 46.230 105.675 52.720 ;
        RECT 106.305 52.210 106.805 52.380 ;
        RECT 106.075 46.955 106.245 51.995 ;
        RECT 106.865 46.955 107.035 51.995 ;
        RECT 106.305 46.570 106.805 46.740 ;
        RECT 107.435 46.230 108.825 52.720 ;
        RECT 109.095 66.010 120.095 66.880 ;
        RECT 109.095 54.870 110.765 66.010 ;
        RECT 111.395 65.495 116.395 65.665 ;
        RECT 111.165 55.240 111.335 65.280 ;
        RECT 116.455 55.240 116.625 65.280 ;
        RECT 117.025 54.870 117.195 66.010 ;
        RECT 117.825 65.495 118.825 65.665 ;
        RECT 117.595 55.240 117.765 65.280 ;
        RECT 118.885 55.240 119.055 65.280 ;
        RECT 119.455 54.870 120.095 66.010 ;
        RECT 109.095 52.800 120.095 54.870 ;
        RECT 109.095 49.310 110.935 52.800 ;
        RECT 112.695 52.720 120.095 52.800 ;
        RECT 111.565 52.290 112.065 52.460 ;
        RECT 111.335 50.035 111.505 52.075 ;
        RECT 112.125 50.035 112.295 52.075 ;
        RECT 111.565 49.650 112.065 49.820 ;
        RECT 112.695 49.310 115.015 52.720 ;
        RECT 115.645 52.210 116.145 52.380 ;
        RECT 109.095 48.590 115.015 49.310 ;
        RECT 102.685 45.740 108.825 46.230 ;
        RECT 109.065 47.980 112.975 48.200 ;
        RECT 97.795 45.310 101.705 45.580 ;
        RECT 109.065 45.580 110.785 47.980 ;
        RECT 111.415 47.470 111.915 47.640 ;
        RECT 111.185 46.260 111.355 47.300 ;
        RECT 111.975 46.260 112.145 47.300 ;
        RECT 111.415 45.920 111.915 46.090 ;
        RECT 112.545 45.580 112.975 47.980 ;
        RECT 113.955 46.230 115.015 48.590 ;
        RECT 115.415 46.955 115.585 51.995 ;
        RECT 116.205 46.955 116.375 51.995 ;
        RECT 115.645 46.570 116.145 46.740 ;
        RECT 116.775 46.230 116.945 52.720 ;
        RECT 117.575 52.210 118.075 52.380 ;
        RECT 117.345 46.955 117.515 51.995 ;
        RECT 118.135 46.955 118.305 51.995 ;
        RECT 117.575 46.570 118.075 46.740 ;
        RECT 118.705 46.230 120.095 52.720 ;
        RECT 120.345 66.010 140.025 66.880 ;
        RECT 120.345 54.870 122.015 66.010 ;
        RECT 122.645 65.495 127.645 65.665 ;
        RECT 122.415 55.240 122.585 65.280 ;
        RECT 127.705 55.240 127.875 65.280 ;
        RECT 128.275 54.870 128.445 66.010 ;
        RECT 130.705 65.980 140.025 66.010 ;
        RECT 129.075 65.495 130.075 65.665 ;
        RECT 128.845 55.240 129.015 65.280 ;
        RECT 130.135 55.240 130.305 65.280 ;
        RECT 130.705 54.870 132.765 65.980 ;
        RECT 133.395 65.465 138.395 65.635 ;
        RECT 133.165 55.210 133.335 65.250 ;
        RECT 138.455 55.210 138.625 65.250 ;
        RECT 120.345 54.840 132.765 54.870 ;
        RECT 139.025 54.840 140.025 65.980 ;
        RECT 120.345 54.720 140.025 54.840 ;
        RECT 120.345 53.550 140.035 54.720 ;
        RECT 120.345 52.800 131.345 53.550 ;
        RECT 120.345 49.310 122.185 52.800 ;
        RECT 123.945 52.720 131.345 52.800 ;
        RECT 122.815 52.290 123.315 52.460 ;
        RECT 122.585 50.035 122.755 52.075 ;
        RECT 123.375 50.035 123.545 52.075 ;
        RECT 122.815 49.650 123.315 49.820 ;
        RECT 123.945 49.310 126.265 52.720 ;
        RECT 126.895 52.210 127.395 52.380 ;
        RECT 120.345 48.590 126.265 49.310 ;
        RECT 113.955 45.740 120.095 46.230 ;
        RECT 120.315 47.980 124.225 48.200 ;
        RECT 109.065 45.310 112.975 45.580 ;
        RECT 120.315 45.580 122.035 47.980 ;
        RECT 122.665 47.470 123.165 47.640 ;
        RECT 122.435 46.260 122.605 47.300 ;
        RECT 123.225 46.260 123.395 47.300 ;
        RECT 122.665 45.920 123.165 46.090 ;
        RECT 123.795 45.580 124.225 47.980 ;
        RECT 125.205 46.230 126.265 48.590 ;
        RECT 126.665 46.955 126.835 51.995 ;
        RECT 127.455 46.955 127.625 51.995 ;
        RECT 126.895 46.570 127.395 46.740 ;
        RECT 128.025 46.230 128.195 52.720 ;
        RECT 128.825 52.210 129.325 52.380 ;
        RECT 128.595 46.955 128.765 51.995 ;
        RECT 129.385 46.955 129.555 51.995 ;
        RECT 128.825 46.570 129.325 46.740 ;
        RECT 129.955 46.230 131.345 52.720 ;
        RECT 125.205 45.740 131.345 46.230 ;
        RECT 120.315 45.310 124.225 45.580 ;
        RECT 25.695 39.770 29.605 40.040 ;
        RECT 18.575 39.120 24.715 39.610 ;
        RECT 18.575 32.630 19.965 39.120 ;
        RECT 20.595 38.610 21.095 38.780 ;
        RECT 20.365 33.355 20.535 38.395 ;
        RECT 21.155 33.355 21.325 38.395 ;
        RECT 20.595 32.970 21.095 33.140 ;
        RECT 21.725 32.630 21.895 39.120 ;
        RECT 22.525 38.610 23.025 38.780 ;
        RECT 22.295 33.355 22.465 38.395 ;
        RECT 23.085 33.355 23.255 38.395 ;
        RECT 23.655 36.760 24.715 39.120 ;
        RECT 25.695 37.370 26.125 39.770 ;
        RECT 26.755 39.260 27.255 39.430 ;
        RECT 26.525 38.050 26.695 39.090 ;
        RECT 27.315 38.050 27.485 39.090 ;
        RECT 26.755 37.710 27.255 37.880 ;
        RECT 27.885 37.370 29.605 39.770 ;
        RECT 36.975 39.770 40.885 40.040 ;
        RECT 25.695 37.150 29.605 37.370 ;
        RECT 29.855 39.120 35.995 39.610 ;
        RECT 23.655 36.040 29.575 36.760 ;
        RECT 22.525 32.970 23.025 33.140 ;
        RECT 23.655 32.630 25.975 36.040 ;
        RECT 26.605 35.530 27.105 35.700 ;
        RECT 26.375 33.275 26.545 35.315 ;
        RECT 27.165 33.275 27.335 35.315 ;
        RECT 26.605 32.890 27.105 33.060 ;
        RECT 18.575 32.550 25.975 32.630 ;
        RECT 27.735 32.550 29.575 36.040 ;
        RECT 18.575 30.480 29.575 32.550 ;
        RECT 18.575 19.340 19.215 30.480 ;
        RECT 19.615 20.070 19.785 30.110 ;
        RECT 20.905 20.070 21.075 30.110 ;
        RECT 19.845 19.685 20.845 19.855 ;
        RECT 21.475 19.340 21.645 30.480 ;
        RECT 22.045 20.070 22.215 30.110 ;
        RECT 27.335 20.070 27.505 30.110 ;
        RECT 22.275 19.685 27.275 19.855 ;
        RECT 27.905 19.340 29.575 30.480 ;
        RECT 18.575 18.470 29.575 19.340 ;
        RECT 29.855 32.630 31.245 39.120 ;
        RECT 31.875 38.610 32.375 38.780 ;
        RECT 31.645 33.355 31.815 38.395 ;
        RECT 32.435 33.355 32.605 38.395 ;
        RECT 31.875 32.970 32.375 33.140 ;
        RECT 33.005 32.630 33.175 39.120 ;
        RECT 33.805 38.610 34.305 38.780 ;
        RECT 33.575 33.355 33.745 38.395 ;
        RECT 34.365 33.355 34.535 38.395 ;
        RECT 34.935 36.760 35.995 39.120 ;
        RECT 36.975 37.370 37.405 39.770 ;
        RECT 38.035 39.260 38.535 39.430 ;
        RECT 37.805 38.050 37.975 39.090 ;
        RECT 38.595 38.050 38.765 39.090 ;
        RECT 38.035 37.710 38.535 37.880 ;
        RECT 39.165 37.370 40.885 39.770 ;
        RECT 48.265 39.750 52.175 40.020 ;
        RECT 36.975 37.150 40.885 37.370 ;
        RECT 41.145 39.100 47.285 39.590 ;
        RECT 34.935 36.040 40.855 36.760 ;
        RECT 33.805 32.970 34.305 33.140 ;
        RECT 34.935 32.630 37.255 36.040 ;
        RECT 37.885 35.530 38.385 35.700 ;
        RECT 37.655 33.275 37.825 35.315 ;
        RECT 38.445 33.275 38.615 35.315 ;
        RECT 37.885 32.890 38.385 33.060 ;
        RECT 29.855 32.550 37.255 32.630 ;
        RECT 39.015 32.550 40.855 36.040 ;
        RECT 29.855 30.480 40.855 32.550 ;
        RECT 29.855 19.340 30.495 30.480 ;
        RECT 30.895 20.070 31.065 30.110 ;
        RECT 32.185 20.070 32.355 30.110 ;
        RECT 31.125 19.685 32.125 19.855 ;
        RECT 32.755 19.340 32.925 30.480 ;
        RECT 33.325 20.070 33.495 30.110 ;
        RECT 38.615 20.070 38.785 30.110 ;
        RECT 33.555 19.685 38.555 19.855 ;
        RECT 39.185 19.340 40.855 30.480 ;
        RECT 29.855 18.470 40.855 19.340 ;
        RECT 41.145 32.610 42.535 39.100 ;
        RECT 43.165 38.590 43.665 38.760 ;
        RECT 42.935 33.335 43.105 38.375 ;
        RECT 43.725 33.335 43.895 38.375 ;
        RECT 43.165 32.950 43.665 33.120 ;
        RECT 44.295 32.610 44.465 39.100 ;
        RECT 45.095 38.590 45.595 38.760 ;
        RECT 44.865 33.335 45.035 38.375 ;
        RECT 45.655 33.335 45.825 38.375 ;
        RECT 46.225 36.740 47.285 39.100 ;
        RECT 48.265 37.350 48.695 39.750 ;
        RECT 49.325 39.240 49.825 39.410 ;
        RECT 49.095 38.030 49.265 39.070 ;
        RECT 49.885 38.030 50.055 39.070 ;
        RECT 49.325 37.690 49.825 37.860 ;
        RECT 50.455 37.350 52.175 39.750 ;
        RECT 59.485 39.750 63.395 40.020 ;
        RECT 48.265 37.130 52.175 37.350 ;
        RECT 52.365 39.100 58.505 39.590 ;
        RECT 46.225 36.020 52.145 36.740 ;
        RECT 45.095 32.950 45.595 33.120 ;
        RECT 46.225 32.610 48.545 36.020 ;
        RECT 49.175 35.510 49.675 35.680 ;
        RECT 48.945 33.255 49.115 35.295 ;
        RECT 49.735 33.255 49.905 35.295 ;
        RECT 49.175 32.870 49.675 33.040 ;
        RECT 41.145 32.530 48.545 32.610 ;
        RECT 50.305 32.530 52.145 36.020 ;
        RECT 41.145 30.460 52.145 32.530 ;
        RECT 41.145 19.320 41.785 30.460 ;
        RECT 42.185 20.050 42.355 30.090 ;
        RECT 43.475 20.050 43.645 30.090 ;
        RECT 42.415 19.665 43.415 19.835 ;
        RECT 44.045 19.320 44.215 30.460 ;
        RECT 44.615 20.050 44.785 30.090 ;
        RECT 49.905 20.050 50.075 30.090 ;
        RECT 44.845 19.665 49.845 19.835 ;
        RECT 50.475 19.320 52.145 30.460 ;
        RECT 41.145 18.450 52.145 19.320 ;
        RECT 52.365 32.610 53.755 39.100 ;
        RECT 54.385 38.590 54.885 38.760 ;
        RECT 54.155 33.335 54.325 38.375 ;
        RECT 54.945 33.335 55.115 38.375 ;
        RECT 54.385 32.950 54.885 33.120 ;
        RECT 55.515 32.610 55.685 39.100 ;
        RECT 56.315 38.590 56.815 38.760 ;
        RECT 56.085 33.335 56.255 38.375 ;
        RECT 56.875 33.335 57.045 38.375 ;
        RECT 57.445 36.740 58.505 39.100 ;
        RECT 59.485 37.350 59.915 39.750 ;
        RECT 60.545 39.240 61.045 39.410 ;
        RECT 60.315 38.030 60.485 39.070 ;
        RECT 61.105 38.030 61.275 39.070 ;
        RECT 60.545 37.690 61.045 37.860 ;
        RECT 61.675 37.350 63.395 39.750 ;
        RECT 70.685 39.750 74.595 40.020 ;
        RECT 59.485 37.130 63.395 37.350 ;
        RECT 63.565 39.100 69.705 39.590 ;
        RECT 57.445 36.020 63.365 36.740 ;
        RECT 56.315 32.950 56.815 33.120 ;
        RECT 57.445 32.610 59.765 36.020 ;
        RECT 60.395 35.510 60.895 35.680 ;
        RECT 60.165 33.255 60.335 35.295 ;
        RECT 60.955 33.255 61.125 35.295 ;
        RECT 60.395 32.870 60.895 33.040 ;
        RECT 52.365 32.530 59.765 32.610 ;
        RECT 61.525 32.530 63.365 36.020 ;
        RECT 52.365 30.460 63.365 32.530 ;
        RECT 52.365 19.320 53.005 30.460 ;
        RECT 53.405 20.050 53.575 30.090 ;
        RECT 54.695 20.050 54.865 30.090 ;
        RECT 53.635 19.665 54.635 19.835 ;
        RECT 55.265 19.320 55.435 30.460 ;
        RECT 55.835 20.050 56.005 30.090 ;
        RECT 61.125 20.050 61.295 30.090 ;
        RECT 56.065 19.665 61.065 19.835 ;
        RECT 61.695 19.320 63.365 30.460 ;
        RECT 52.365 18.450 63.365 19.320 ;
        RECT 63.565 32.610 64.955 39.100 ;
        RECT 65.585 38.590 66.085 38.760 ;
        RECT 65.355 33.335 65.525 38.375 ;
        RECT 66.145 33.335 66.315 38.375 ;
        RECT 65.585 32.950 66.085 33.120 ;
        RECT 66.715 32.610 66.885 39.100 ;
        RECT 67.515 38.590 68.015 38.760 ;
        RECT 67.285 33.335 67.455 38.375 ;
        RECT 68.075 33.335 68.245 38.375 ;
        RECT 68.645 36.740 69.705 39.100 ;
        RECT 70.685 37.350 71.115 39.750 ;
        RECT 71.745 39.240 72.245 39.410 ;
        RECT 71.515 38.030 71.685 39.070 ;
        RECT 72.305 38.030 72.475 39.070 ;
        RECT 71.745 37.690 72.245 37.860 ;
        RECT 72.875 37.350 74.595 39.750 ;
        RECT 81.975 39.740 85.885 40.010 ;
        RECT 70.685 37.130 74.595 37.350 ;
        RECT 74.855 39.090 80.995 39.580 ;
        RECT 68.645 36.020 74.565 36.740 ;
        RECT 67.515 32.950 68.015 33.120 ;
        RECT 68.645 32.610 70.965 36.020 ;
        RECT 71.595 35.510 72.095 35.680 ;
        RECT 71.365 33.255 71.535 35.295 ;
        RECT 72.155 33.255 72.325 35.295 ;
        RECT 71.595 32.870 72.095 33.040 ;
        RECT 63.565 32.530 70.965 32.610 ;
        RECT 72.725 32.530 74.565 36.020 ;
        RECT 63.565 30.460 74.565 32.530 ;
        RECT 63.565 19.320 64.205 30.460 ;
        RECT 64.605 20.050 64.775 30.090 ;
        RECT 65.895 20.050 66.065 30.090 ;
        RECT 64.835 19.665 65.835 19.835 ;
        RECT 66.465 19.320 66.635 30.460 ;
        RECT 67.035 20.050 67.205 30.090 ;
        RECT 72.325 20.050 72.495 30.090 ;
        RECT 67.265 19.665 72.265 19.835 ;
        RECT 72.895 19.320 74.565 30.460 ;
        RECT 63.565 18.450 74.565 19.320 ;
        RECT 74.855 32.600 76.245 39.090 ;
        RECT 76.875 38.580 77.375 38.750 ;
        RECT 76.645 33.325 76.815 38.365 ;
        RECT 77.435 33.325 77.605 38.365 ;
        RECT 76.875 32.940 77.375 33.110 ;
        RECT 78.005 32.600 78.175 39.090 ;
        RECT 78.805 38.580 79.305 38.750 ;
        RECT 78.575 33.325 78.745 38.365 ;
        RECT 79.365 33.325 79.535 38.365 ;
        RECT 79.935 36.730 80.995 39.090 ;
        RECT 81.975 37.340 82.405 39.740 ;
        RECT 83.035 39.230 83.535 39.400 ;
        RECT 82.805 38.020 82.975 39.060 ;
        RECT 83.595 38.020 83.765 39.060 ;
        RECT 83.035 37.680 83.535 37.850 ;
        RECT 84.165 37.340 85.885 39.740 ;
        RECT 93.215 39.760 97.125 40.030 ;
        RECT 81.975 37.120 85.885 37.340 ;
        RECT 86.095 39.110 92.235 39.600 ;
        RECT 79.935 36.010 85.855 36.730 ;
        RECT 78.805 32.940 79.305 33.110 ;
        RECT 79.935 32.600 82.255 36.010 ;
        RECT 82.885 35.500 83.385 35.670 ;
        RECT 82.655 33.245 82.825 35.285 ;
        RECT 83.445 33.245 83.615 35.285 ;
        RECT 82.885 32.860 83.385 33.030 ;
        RECT 74.855 32.520 82.255 32.600 ;
        RECT 84.015 32.520 85.855 36.010 ;
        RECT 74.855 30.450 85.855 32.520 ;
        RECT 74.855 19.310 75.495 30.450 ;
        RECT 75.895 20.040 76.065 30.080 ;
        RECT 77.185 20.040 77.355 30.080 ;
        RECT 76.125 19.655 77.125 19.825 ;
        RECT 77.755 19.310 77.925 30.450 ;
        RECT 78.325 20.040 78.495 30.080 ;
        RECT 83.615 20.040 83.785 30.080 ;
        RECT 78.555 19.655 83.555 19.825 ;
        RECT 84.185 19.310 85.855 30.450 ;
        RECT 74.855 18.440 85.855 19.310 ;
        RECT 86.095 32.620 87.485 39.110 ;
        RECT 88.115 38.600 88.615 38.770 ;
        RECT 87.885 33.345 88.055 38.385 ;
        RECT 88.675 33.345 88.845 38.385 ;
        RECT 88.115 32.960 88.615 33.130 ;
        RECT 89.245 32.620 89.415 39.110 ;
        RECT 90.045 38.600 90.545 38.770 ;
        RECT 89.815 33.345 89.985 38.385 ;
        RECT 90.605 33.345 90.775 38.385 ;
        RECT 91.175 36.750 92.235 39.110 ;
        RECT 93.215 37.360 93.645 39.760 ;
        RECT 94.275 39.250 94.775 39.420 ;
        RECT 94.045 38.040 94.215 39.080 ;
        RECT 94.835 38.040 95.005 39.080 ;
        RECT 94.275 37.700 94.775 37.870 ;
        RECT 95.405 37.360 97.125 39.760 ;
        RECT 104.425 39.780 108.335 40.050 ;
        RECT 93.215 37.140 97.125 37.360 ;
        RECT 97.305 39.130 103.445 39.620 ;
        RECT 91.175 36.030 97.095 36.750 ;
        RECT 90.045 32.960 90.545 33.130 ;
        RECT 91.175 32.620 93.495 36.030 ;
        RECT 94.125 35.520 94.625 35.690 ;
        RECT 93.895 33.265 94.065 35.305 ;
        RECT 94.685 33.265 94.855 35.305 ;
        RECT 94.125 32.880 94.625 33.050 ;
        RECT 86.095 32.540 93.495 32.620 ;
        RECT 95.255 32.540 97.095 36.030 ;
        RECT 86.095 30.470 97.095 32.540 ;
        RECT 86.095 19.330 86.735 30.470 ;
        RECT 87.135 20.060 87.305 30.100 ;
        RECT 88.425 20.060 88.595 30.100 ;
        RECT 87.365 19.675 88.365 19.845 ;
        RECT 88.995 19.330 89.165 30.470 ;
        RECT 89.565 20.060 89.735 30.100 ;
        RECT 94.855 20.060 95.025 30.100 ;
        RECT 89.795 19.675 94.795 19.845 ;
        RECT 95.425 19.330 97.095 30.470 ;
        RECT 86.095 18.460 97.095 19.330 ;
        RECT 97.305 32.640 98.695 39.130 ;
        RECT 99.325 38.620 99.825 38.790 ;
        RECT 99.095 33.365 99.265 38.405 ;
        RECT 99.885 33.365 100.055 38.405 ;
        RECT 99.325 32.980 99.825 33.150 ;
        RECT 100.455 32.640 100.625 39.130 ;
        RECT 101.255 38.620 101.755 38.790 ;
        RECT 101.025 33.365 101.195 38.405 ;
        RECT 101.815 33.365 101.985 38.405 ;
        RECT 102.385 36.770 103.445 39.130 ;
        RECT 104.425 37.380 104.855 39.780 ;
        RECT 105.485 39.270 105.985 39.440 ;
        RECT 105.255 38.060 105.425 39.100 ;
        RECT 106.045 38.060 106.215 39.100 ;
        RECT 105.485 37.720 105.985 37.890 ;
        RECT 106.615 37.380 108.335 39.780 ;
        RECT 115.625 39.820 119.535 40.090 ;
        RECT 104.425 37.160 108.335 37.380 ;
        RECT 108.505 39.170 114.645 39.660 ;
        RECT 102.385 36.050 108.305 36.770 ;
        RECT 101.255 32.980 101.755 33.150 ;
        RECT 102.385 32.640 104.705 36.050 ;
        RECT 105.335 35.540 105.835 35.710 ;
        RECT 105.105 33.285 105.275 35.325 ;
        RECT 105.895 33.285 106.065 35.325 ;
        RECT 105.335 32.900 105.835 33.070 ;
        RECT 97.305 32.560 104.705 32.640 ;
        RECT 106.465 32.560 108.305 36.050 ;
        RECT 97.305 30.490 108.305 32.560 ;
        RECT 97.305 19.350 97.945 30.490 ;
        RECT 98.345 20.080 98.515 30.120 ;
        RECT 99.635 20.080 99.805 30.120 ;
        RECT 98.575 19.695 99.575 19.865 ;
        RECT 100.205 19.350 100.375 30.490 ;
        RECT 100.775 20.080 100.945 30.120 ;
        RECT 106.065 20.080 106.235 30.120 ;
        RECT 101.005 19.695 106.005 19.865 ;
        RECT 106.635 19.350 108.305 30.490 ;
        RECT 97.305 18.480 108.305 19.350 ;
        RECT 108.505 32.680 109.895 39.170 ;
        RECT 110.525 38.660 111.025 38.830 ;
        RECT 110.295 33.405 110.465 38.445 ;
        RECT 111.085 33.405 111.255 38.445 ;
        RECT 110.525 33.020 111.025 33.190 ;
        RECT 111.655 32.680 111.825 39.170 ;
        RECT 112.455 38.660 112.955 38.830 ;
        RECT 112.225 33.405 112.395 38.445 ;
        RECT 113.015 33.405 113.185 38.445 ;
        RECT 113.585 36.810 114.645 39.170 ;
        RECT 115.625 37.420 116.055 39.820 ;
        RECT 116.685 39.310 117.185 39.480 ;
        RECT 116.455 38.100 116.625 39.140 ;
        RECT 117.245 38.100 117.415 39.140 ;
        RECT 116.685 37.760 117.185 37.930 ;
        RECT 117.815 37.420 119.535 39.820 ;
        RECT 126.835 39.840 130.745 40.110 ;
        RECT 115.625 37.200 119.535 37.420 ;
        RECT 119.715 39.190 125.855 39.680 ;
        RECT 113.585 36.090 119.505 36.810 ;
        RECT 112.455 33.020 112.955 33.190 ;
        RECT 113.585 32.680 115.905 36.090 ;
        RECT 116.535 35.580 117.035 35.750 ;
        RECT 116.305 33.325 116.475 35.365 ;
        RECT 117.095 33.325 117.265 35.365 ;
        RECT 116.535 32.940 117.035 33.110 ;
        RECT 108.505 32.600 115.905 32.680 ;
        RECT 117.665 32.600 119.505 36.090 ;
        RECT 108.505 30.530 119.505 32.600 ;
        RECT 108.505 19.390 109.145 30.530 ;
        RECT 109.545 20.120 109.715 30.160 ;
        RECT 110.835 20.120 111.005 30.160 ;
        RECT 109.775 19.735 110.775 19.905 ;
        RECT 111.405 19.390 111.575 30.530 ;
        RECT 111.975 20.120 112.145 30.160 ;
        RECT 117.265 20.120 117.435 30.160 ;
        RECT 112.205 19.735 117.205 19.905 ;
        RECT 117.835 19.390 119.505 30.530 ;
        RECT 108.505 18.520 119.505 19.390 ;
        RECT 119.715 32.700 121.105 39.190 ;
        RECT 121.735 38.680 122.235 38.850 ;
        RECT 121.505 33.425 121.675 38.465 ;
        RECT 122.295 33.425 122.465 38.465 ;
        RECT 121.735 33.040 122.235 33.210 ;
        RECT 122.865 32.700 123.035 39.190 ;
        RECT 123.665 38.680 124.165 38.850 ;
        RECT 123.435 33.425 123.605 38.465 ;
        RECT 124.225 33.425 124.395 38.465 ;
        RECT 124.795 36.830 125.855 39.190 ;
        RECT 126.835 37.440 127.265 39.840 ;
        RECT 127.895 39.330 128.395 39.500 ;
        RECT 127.665 38.120 127.835 39.160 ;
        RECT 128.455 38.120 128.625 39.160 ;
        RECT 127.895 37.780 128.395 37.950 ;
        RECT 129.025 37.440 130.745 39.840 ;
        RECT 126.835 37.220 130.745 37.440 ;
        RECT 124.795 36.110 130.715 36.830 ;
        RECT 123.665 33.040 124.165 33.210 ;
        RECT 124.795 32.700 127.115 36.110 ;
        RECT 127.745 35.600 128.245 35.770 ;
        RECT 127.515 33.345 127.685 35.385 ;
        RECT 128.305 33.345 128.475 35.385 ;
        RECT 127.745 32.960 128.245 33.130 ;
        RECT 119.715 32.620 127.115 32.700 ;
        RECT 128.875 32.620 130.715 36.110 ;
        RECT 119.715 31.140 130.715 32.620 ;
        RECT 119.715 30.550 139.465 31.140 ;
        RECT 119.715 19.410 120.355 30.550 ;
        RECT 120.755 20.140 120.925 30.180 ;
        RECT 122.045 20.140 122.215 30.180 ;
        RECT 120.985 19.755 121.985 19.925 ;
        RECT 122.615 19.410 122.785 30.550 ;
        RECT 129.045 30.520 139.465 30.550 ;
        RECT 123.185 20.140 123.355 30.180 ;
        RECT 128.475 20.140 128.645 30.180 ;
        RECT 123.415 19.755 128.415 19.925 ;
        RECT 129.045 19.410 132.075 30.520 ;
        RECT 132.475 20.110 132.645 30.150 ;
        RECT 137.765 20.110 137.935 30.150 ;
        RECT 132.705 19.725 137.705 19.895 ;
        RECT 119.715 19.380 132.075 19.410 ;
        RECT 138.335 19.380 139.465 30.520 ;
        RECT 119.715 18.540 139.465 19.380 ;
        RECT 131.925 18.520 139.465 18.540 ;
      LAYER met1 ;
        RECT 135.340 223.880 136.790 225.180 ;
        RECT 29.840 211.050 127.820 211.530 ;
        RECT 29.840 208.330 127.820 208.810 ;
        RECT 68.550 208.130 68.870 208.190 ;
        RECT 80.065 208.130 80.355 208.175 ;
        RECT 83.730 208.130 84.050 208.190 ;
        RECT 68.550 207.990 79.820 208.130 ;
        RECT 68.550 207.930 68.870 207.990 ;
        RECT 69.125 207.790 69.415 207.835 ;
        RECT 72.245 207.790 72.535 207.835 ;
        RECT 74.135 207.790 74.425 207.835 ;
        RECT 69.125 207.650 74.425 207.790 ;
        RECT 79.680 207.790 79.820 207.990 ;
        RECT 80.065 207.990 84.050 208.130 ;
        RECT 80.065 207.945 80.355 207.990 ;
        RECT 83.730 207.930 84.050 207.990 ;
        RECT 82.810 207.790 83.130 207.850 ;
        RECT 84.305 207.790 84.595 207.835 ;
        RECT 87.425 207.790 87.715 207.835 ;
        RECT 89.315 207.790 89.605 207.835 ;
        RECT 79.680 207.650 83.960 207.790 ;
        RECT 69.125 207.605 69.415 207.650 ;
        RECT 72.245 207.605 72.535 207.650 ;
        RECT 74.135 207.605 74.425 207.650 ;
        RECT 82.810 207.590 83.130 207.650 ;
        RECT 66.265 207.450 66.555 207.495 ;
        RECT 71.310 207.450 71.630 207.510 ;
        RECT 66.265 207.310 71.630 207.450 ;
        RECT 66.265 207.265 66.555 207.310 ;
        RECT 71.310 207.250 71.630 207.310 ;
        RECT 73.625 207.450 73.915 207.495 ;
        RECT 80.050 207.450 80.370 207.510 ;
        RECT 73.625 207.310 80.370 207.450 ;
        RECT 73.625 207.265 73.915 207.310 ;
        RECT 80.050 207.250 80.370 207.310 ;
        RECT 81.430 207.250 81.750 207.510 ;
        RECT 83.820 207.450 83.960 207.650 ;
        RECT 84.305 207.650 89.605 207.790 ;
        RECT 84.305 207.605 84.595 207.650 ;
        RECT 87.425 207.605 87.715 207.650 ;
        RECT 89.315 207.605 89.605 207.650 ;
        RECT 88.330 207.450 88.650 207.510 ;
        RECT 83.820 207.310 92.700 207.450 ;
        RECT 88.330 207.250 88.650 207.310 ;
        RECT 68.090 207.130 68.410 207.170 ;
        RECT 68.045 206.910 68.410 207.130 ;
        RECT 69.125 207.110 69.415 207.155 ;
        RECT 72.705 207.110 72.995 207.155 ;
        RECT 74.540 207.110 74.830 207.155 ;
        RECT 69.125 206.970 74.830 207.110 ;
        RECT 69.125 206.925 69.415 206.970 ;
        RECT 72.705 206.925 72.995 206.970 ;
        RECT 74.540 206.925 74.830 206.970 ;
        RECT 75.005 207.110 75.295 207.155 ;
        RECT 75.450 207.110 75.770 207.170 ;
        RECT 75.005 206.970 75.770 207.110 ;
        RECT 75.005 206.925 75.295 206.970 ;
        RECT 75.450 206.910 75.770 206.970 ;
        RECT 76.385 206.925 76.675 207.155 ;
        RECT 76.830 207.110 77.150 207.170 ;
        RECT 78.225 207.110 78.515 207.155 ;
        RECT 76.830 206.970 78.515 207.110 ;
        RECT 68.045 206.815 68.335 206.910 ;
        RECT 67.745 206.770 68.335 206.815 ;
        RECT 70.985 206.770 71.635 206.815 ;
        RECT 67.745 206.630 71.635 206.770 ;
        RECT 76.460 206.770 76.600 206.925 ;
        RECT 76.830 206.910 77.150 206.970 ;
        RECT 78.225 206.925 78.515 206.970 ;
        RECT 79.130 207.110 79.450 207.170 ;
        RECT 79.605 207.110 79.895 207.155 ;
        RECT 79.130 206.970 79.895 207.110 ;
        RECT 79.130 206.910 79.450 206.970 ;
        RECT 79.605 206.925 79.895 206.970 ;
        RECT 82.350 206.770 82.670 206.830 ;
        RECT 83.225 206.815 83.515 207.130 ;
        RECT 84.305 207.110 84.595 207.155 ;
        RECT 87.885 207.110 88.175 207.155 ;
        RECT 89.720 207.110 90.010 207.155 ;
        RECT 84.305 206.970 90.010 207.110 ;
        RECT 84.305 206.925 84.595 206.970 ;
        RECT 87.885 206.925 88.175 206.970 ;
        RECT 89.720 206.925 90.010 206.970 ;
        RECT 90.170 206.910 90.490 207.170 ;
        RECT 92.560 207.155 92.700 207.310 ;
        RECT 92.485 207.110 92.775 207.155 ;
        RECT 94.310 207.110 94.630 207.170 ;
        RECT 92.485 206.970 94.630 207.110 ;
        RECT 92.485 206.925 92.775 206.970 ;
        RECT 94.310 206.910 94.630 206.970 ;
        RECT 76.460 206.630 82.670 206.770 ;
        RECT 67.745 206.585 68.035 206.630 ;
        RECT 70.985 206.585 71.635 206.630 ;
        RECT 82.350 206.570 82.670 206.630 ;
        RECT 82.925 206.770 83.515 206.815 ;
        RECT 86.165 206.770 86.815 206.815 ;
        RECT 82.925 206.630 87.180 206.770 ;
        RECT 82.925 206.585 83.215 206.630 ;
        RECT 86.165 206.585 86.815 206.630 ;
        RECT 76.370 206.430 76.690 206.490 ;
        RECT 77.305 206.430 77.595 206.475 ;
        RECT 76.370 206.290 77.595 206.430 ;
        RECT 76.370 206.230 76.690 206.290 ;
        RECT 77.305 206.245 77.595 206.290 ;
        RECT 80.985 206.430 81.275 206.475 ;
        RECT 84.190 206.430 84.510 206.490 ;
        RECT 80.985 206.290 84.510 206.430 ;
        RECT 87.040 206.430 87.180 206.630 ;
        RECT 88.790 206.570 89.110 206.830 ;
        RECT 89.250 206.770 89.570 206.830 ;
        RECT 92.025 206.770 92.315 206.815 ;
        RECT 89.250 206.630 92.315 206.770 ;
        RECT 89.250 206.570 89.570 206.630 ;
        RECT 92.025 206.585 92.315 206.630 ;
        RECT 89.710 206.430 90.030 206.490 ;
        RECT 87.040 206.290 90.030 206.430 ;
        RECT 80.985 206.245 81.275 206.290 ;
        RECT 84.190 206.230 84.510 206.290 ;
        RECT 89.710 206.230 90.030 206.290 ;
        RECT 29.840 205.610 127.820 206.090 ;
        RECT 67.645 205.410 67.935 205.455 ;
        RECT 68.090 205.410 68.410 205.470 ;
        RECT 67.645 205.270 68.410 205.410 ;
        RECT 67.645 205.225 67.935 205.270 ;
        RECT 68.090 205.210 68.410 205.270 ;
        RECT 76.370 205.410 76.690 205.470 ;
        RECT 79.145 205.410 79.435 205.455 ;
        RECT 80.050 205.410 80.370 205.470 ;
        RECT 76.370 205.270 77.520 205.410 ;
        RECT 76.370 205.210 76.690 205.270 ;
        RECT 68.550 205.070 68.870 205.130 ;
        RECT 77.380 205.115 77.520 205.270 ;
        RECT 79.145 205.270 80.370 205.410 ;
        RECT 79.145 205.225 79.435 205.270 ;
        RECT 80.050 205.210 80.370 205.270 ;
        RECT 82.350 205.210 82.670 205.470 ;
        RECT 88.345 205.410 88.635 205.455 ;
        RECT 88.790 205.410 89.110 205.470 ;
        RECT 88.345 205.270 89.110 205.410 ;
        RECT 88.345 205.225 88.635 205.270 ;
        RECT 88.790 205.210 89.110 205.270 ;
        RECT 89.710 205.210 90.030 205.470 ;
        RECT 68.180 204.930 68.870 205.070 ;
        RECT 68.180 204.775 68.320 204.930 ;
        RECT 68.550 204.870 68.870 204.930 ;
        RECT 71.425 205.070 71.715 205.115 ;
        RECT 74.665 205.070 75.315 205.115 ;
        RECT 71.425 204.930 75.315 205.070 ;
        RECT 71.425 204.885 72.015 204.930 ;
        RECT 74.665 204.885 75.315 204.930 ;
        RECT 77.305 204.885 77.595 205.115 ;
        RECT 83.125 205.070 83.415 205.115 ;
        RECT 79.220 204.930 83.415 205.070 ;
        RECT 68.105 204.545 68.395 204.775 ;
        RECT 69.010 204.730 69.330 204.790 ;
        RECT 71.725 204.730 72.015 204.885 ;
        RECT 69.010 204.590 72.015 204.730 ;
        RECT 69.010 204.530 69.330 204.590 ;
        RECT 71.725 204.570 72.015 204.590 ;
        RECT 72.805 204.730 73.095 204.775 ;
        RECT 76.385 204.730 76.675 204.775 ;
        RECT 78.220 204.730 78.510 204.775 ;
        RECT 72.805 204.590 78.510 204.730 ;
        RECT 72.805 204.545 73.095 204.590 ;
        RECT 76.385 204.545 76.675 204.590 ;
        RECT 78.220 204.545 78.510 204.590 ;
        RECT 68.565 204.390 68.855 204.435 ;
        RECT 72.230 204.390 72.550 204.450 ;
        RECT 68.565 204.250 72.550 204.390 ;
        RECT 68.565 204.205 68.855 204.250 ;
        RECT 72.230 204.190 72.550 204.250 ;
        RECT 75.450 204.390 75.770 204.450 ;
        RECT 78.685 204.390 78.975 204.435 ;
        RECT 75.450 204.250 78.975 204.390 ;
        RECT 75.450 204.190 75.770 204.250 ;
        RECT 78.685 204.205 78.975 204.250 ;
        RECT 72.805 204.050 73.095 204.095 ;
        RECT 75.925 204.050 76.215 204.095 ;
        RECT 77.815 204.050 78.105 204.095 ;
        RECT 72.805 203.910 78.105 204.050 ;
        RECT 72.805 203.865 73.095 203.910 ;
        RECT 75.925 203.865 76.215 203.910 ;
        RECT 77.815 203.865 78.105 203.910 ;
        RECT 76.370 203.710 76.690 203.770 ;
        RECT 79.220 203.710 79.360 204.930 ;
        RECT 83.125 204.885 83.415 204.930 ;
        RECT 84.190 204.870 84.510 205.130 ;
        RECT 91.105 205.070 91.395 205.115 ;
        RECT 86.120 204.930 91.395 205.070 ;
        RECT 80.970 204.530 81.290 204.790 ;
        RECT 86.120 204.450 86.260 204.930 ;
        RECT 91.105 204.885 91.395 204.930 ;
        RECT 86.505 204.545 86.795 204.775 ;
        RECT 88.330 204.730 88.650 204.790 ;
        RECT 90.185 204.730 90.475 204.775 ;
        RECT 88.330 204.590 90.475 204.730 ;
        RECT 80.050 204.390 80.370 204.450 ;
        RECT 80.525 204.390 80.815 204.435 ;
        RECT 80.050 204.250 80.815 204.390 ;
        RECT 80.050 204.190 80.370 204.250 ;
        RECT 80.525 204.205 80.815 204.250 ;
        RECT 76.370 203.570 79.360 203.710 ;
        RECT 80.600 203.710 80.740 204.205 ;
        RECT 86.030 204.190 86.350 204.450 ;
        RECT 84.650 204.050 84.970 204.110 ;
        RECT 86.580 204.050 86.720 204.545 ;
        RECT 88.330 204.530 88.650 204.590 ;
        RECT 90.185 204.545 90.475 204.590 ;
        RECT 90.630 204.530 90.950 204.790 ;
        RECT 91.550 204.730 91.870 204.790 ;
        RECT 92.945 204.730 93.235 204.775 ;
        RECT 91.550 204.590 93.235 204.730 ;
        RECT 91.550 204.530 91.870 204.590 ;
        RECT 92.945 204.545 93.235 204.590 ;
        RECT 95.245 204.545 95.535 204.775 ;
        RECT 87.410 204.390 87.730 204.450 ;
        RECT 95.320 204.390 95.460 204.545 ;
        RECT 87.410 204.250 95.460 204.390 ;
        RECT 87.410 204.190 87.730 204.250 ;
        RECT 94.325 204.050 94.615 204.095 ;
        RECT 84.650 203.910 86.720 204.050 ;
        RECT 87.040 203.910 94.615 204.050 ;
        RECT 84.650 203.850 84.970 203.910 ;
        RECT 87.040 203.770 87.180 203.910 ;
        RECT 94.325 203.865 94.615 203.910 ;
        RECT 83.285 203.710 83.575 203.755 ;
        RECT 80.600 203.570 83.575 203.710 ;
        RECT 76.370 203.510 76.690 203.570 ;
        RECT 83.285 203.525 83.575 203.570 ;
        RECT 86.950 203.510 87.270 203.770 ;
        RECT 93.405 203.710 93.695 203.755 ;
        RECT 96.150 203.710 96.470 203.770 ;
        RECT 93.405 203.570 96.470 203.710 ;
        RECT 93.405 203.525 93.695 203.570 ;
        RECT 96.150 203.510 96.470 203.570 ;
        RECT 29.840 202.890 127.820 203.370 ;
        RECT 69.010 202.490 69.330 202.750 ;
        RECT 71.310 202.690 71.630 202.750 ;
        RECT 76.845 202.690 77.135 202.735 ;
        RECT 71.310 202.550 77.135 202.690 ;
        RECT 71.310 202.490 71.630 202.550 ;
        RECT 76.845 202.505 77.135 202.550 ;
        RECT 79.130 202.490 79.450 202.750 ;
        RECT 90.170 202.690 90.490 202.750 ;
        RECT 110.870 202.690 111.190 202.750 ;
        RECT 88.420 202.550 97.760 202.690 ;
        RECT 73.165 202.350 73.455 202.395 ;
        RECT 80.970 202.350 81.290 202.410 ;
        RECT 73.165 202.210 81.290 202.350 ;
        RECT 73.165 202.165 73.455 202.210 ;
        RECT 80.970 202.150 81.290 202.210 ;
        RECT 82.465 202.350 82.755 202.395 ;
        RECT 85.585 202.350 85.875 202.395 ;
        RECT 87.475 202.350 87.765 202.395 ;
        RECT 82.465 202.210 87.765 202.350 ;
        RECT 82.465 202.165 82.755 202.210 ;
        RECT 85.585 202.165 85.875 202.210 ;
        RECT 87.475 202.165 87.765 202.210 ;
        RECT 79.130 202.010 79.450 202.070 ;
        RECT 76.460 201.870 79.450 202.010 ;
        RECT 68.550 201.470 68.870 201.730 ;
        RECT 70.405 201.670 70.695 201.715 ;
        RECT 71.310 201.670 71.630 201.730 ;
        RECT 76.460 201.715 76.600 201.870 ;
        RECT 79.130 201.810 79.450 201.870 ;
        RECT 86.950 201.810 87.270 202.070 ;
        RECT 88.420 202.055 88.560 202.550 ;
        RECT 90.170 202.490 90.490 202.550 ;
        RECT 91.665 202.350 91.955 202.395 ;
        RECT 94.785 202.350 95.075 202.395 ;
        RECT 96.675 202.350 96.965 202.395 ;
        RECT 91.665 202.210 96.965 202.350 ;
        RECT 91.665 202.165 91.955 202.210 ;
        RECT 94.785 202.165 95.075 202.210 ;
        RECT 96.675 202.165 96.965 202.210 ;
        RECT 88.345 201.825 88.635 202.055 ;
        RECT 96.150 201.810 96.470 202.070 ;
        RECT 70.405 201.530 71.630 201.670 ;
        RECT 70.405 201.485 70.695 201.530 ;
        RECT 71.310 201.470 71.630 201.530 ;
        RECT 76.385 201.485 76.675 201.715 ;
        RECT 78.225 201.670 78.515 201.715 ;
        RECT 79.590 201.670 79.910 201.730 ;
        RECT 97.620 201.715 97.760 202.550 ;
        RECT 110.870 202.550 119.380 202.690 ;
        RECT 110.870 202.490 111.190 202.550 ;
        RECT 109.965 202.350 110.255 202.395 ;
        RECT 112.250 202.350 112.570 202.410 ;
        RECT 109.965 202.210 112.570 202.350 ;
        RECT 109.965 202.165 110.255 202.210 ;
        RECT 112.250 202.150 112.570 202.210 ;
        RECT 113.285 202.350 113.575 202.395 ;
        RECT 116.405 202.350 116.695 202.395 ;
        RECT 118.295 202.350 118.585 202.395 ;
        RECT 113.285 202.210 118.585 202.350 ;
        RECT 113.285 202.165 113.575 202.210 ;
        RECT 116.405 202.165 116.695 202.210 ;
        RECT 118.295 202.165 118.585 202.210 ;
        RECT 107.205 202.010 107.495 202.055 ;
        RECT 110.410 202.010 110.730 202.070 ;
        RECT 107.205 201.870 110.730 202.010 ;
        RECT 107.205 201.825 107.495 201.870 ;
        RECT 110.410 201.810 110.730 201.870 ;
        RECT 114.090 202.010 114.410 202.070 ;
        RECT 117.785 202.010 118.075 202.055 ;
        RECT 114.090 201.870 118.075 202.010 ;
        RECT 114.090 201.810 114.410 201.870 ;
        RECT 117.785 201.825 118.075 201.870 ;
        RECT 78.225 201.530 79.910 201.670 ;
        RECT 78.225 201.485 78.515 201.530 ;
        RECT 73.610 201.330 73.930 201.390 ;
        RECT 78.300 201.330 78.440 201.485 ;
        RECT 79.590 201.470 79.910 201.530 ;
        RECT 81.385 201.375 81.675 201.690 ;
        RECT 82.465 201.670 82.755 201.715 ;
        RECT 86.045 201.670 86.335 201.715 ;
        RECT 87.880 201.670 88.170 201.715 ;
        RECT 82.465 201.530 88.170 201.670 ;
        RECT 82.465 201.485 82.755 201.530 ;
        RECT 86.045 201.485 86.335 201.530 ;
        RECT 87.880 201.485 88.170 201.530 ;
        RECT 73.610 201.190 78.440 201.330 ;
        RECT 81.085 201.330 81.675 201.375 ;
        RECT 84.325 201.330 84.975 201.375 ;
        RECT 89.250 201.330 89.570 201.390 ;
        RECT 90.585 201.375 90.875 201.690 ;
        RECT 91.665 201.670 91.955 201.715 ;
        RECT 95.245 201.670 95.535 201.715 ;
        RECT 97.080 201.670 97.370 201.715 ;
        RECT 91.665 201.530 97.370 201.670 ;
        RECT 91.665 201.485 91.955 201.530 ;
        RECT 95.245 201.485 95.535 201.530 ;
        RECT 97.080 201.485 97.370 201.530 ;
        RECT 97.545 201.670 97.835 201.715 ;
        RECT 110.870 201.670 111.190 201.730 ;
        RECT 119.240 201.715 119.380 202.550 ;
        RECT 97.545 201.530 111.190 201.670 ;
        RECT 97.545 201.485 97.835 201.530 ;
        RECT 110.870 201.470 111.190 201.530 ;
        RECT 93.850 201.375 94.170 201.390 ;
        RECT 112.205 201.375 112.495 201.690 ;
        RECT 113.285 201.670 113.575 201.715 ;
        RECT 116.865 201.670 117.155 201.715 ;
        RECT 118.700 201.670 118.990 201.715 ;
        RECT 113.285 201.530 118.990 201.670 ;
        RECT 113.285 201.485 113.575 201.530 ;
        RECT 116.865 201.485 117.155 201.530 ;
        RECT 118.700 201.485 118.990 201.530 ;
        RECT 119.165 201.670 119.455 201.715 ;
        RECT 119.165 201.530 119.840 201.670 ;
        RECT 119.165 201.485 119.455 201.530 ;
        RECT 119.700 201.390 119.840 201.530 ;
        RECT 115.470 201.375 115.790 201.390 ;
        RECT 81.085 201.190 89.570 201.330 ;
        RECT 73.610 201.130 73.930 201.190 ;
        RECT 81.085 201.145 81.375 201.190 ;
        RECT 84.325 201.145 84.975 201.190 ;
        RECT 89.250 201.130 89.570 201.190 ;
        RECT 90.285 201.330 90.875 201.375 ;
        RECT 93.525 201.330 94.175 201.375 ;
        RECT 90.285 201.190 94.175 201.330 ;
        RECT 90.285 201.145 90.575 201.190 ;
        RECT 93.525 201.145 94.175 201.190 ;
        RECT 111.905 201.330 112.495 201.375 ;
        RECT 115.145 201.330 115.795 201.375 ;
        RECT 111.905 201.190 115.795 201.330 ;
        RECT 111.905 201.145 112.195 201.190 ;
        RECT 115.145 201.145 115.795 201.190 ;
        RECT 93.850 201.130 94.170 201.145 ;
        RECT 115.470 201.130 115.790 201.145 ;
        RECT 119.610 201.130 119.930 201.390 ;
        RECT 79.605 200.990 79.895 201.035 ;
        RECT 82.350 200.990 82.670 201.050 ;
        RECT 79.605 200.850 82.670 200.990 ;
        RECT 79.605 200.805 79.895 200.850 ;
        RECT 82.350 200.790 82.670 200.850 ;
        RECT 85.570 200.990 85.890 201.050 ;
        RECT 88.805 200.990 89.095 201.035 ;
        RECT 85.570 200.850 89.095 200.990 ;
        RECT 85.570 200.790 85.890 200.850 ;
        RECT 88.805 200.805 89.095 200.850 ;
        RECT 29.840 200.170 127.820 200.650 ;
        RECT 75.465 199.970 75.755 200.015 ;
        RECT 76.370 199.970 76.690 200.030 ;
        RECT 75.465 199.830 76.690 199.970 ;
        RECT 75.465 199.785 75.755 199.830 ;
        RECT 76.370 199.770 76.690 199.830 ;
        RECT 79.130 199.770 79.450 200.030 ;
        RECT 80.050 199.770 80.370 200.030 ;
        RECT 81.430 199.970 81.750 200.030 ;
        RECT 82.365 199.970 82.655 200.015 ;
        RECT 81.430 199.830 82.655 199.970 ;
        RECT 81.430 199.770 81.750 199.830 ;
        RECT 82.365 199.785 82.655 199.830 ;
        RECT 93.850 199.770 94.170 200.030 ;
        RECT 109.490 199.970 109.810 200.030 ;
        RECT 99.460 199.830 109.810 199.970 ;
        RECT 75.910 199.630 76.230 199.690 ;
        RECT 81.520 199.630 81.660 199.770 ;
        RECT 73.240 199.490 77.520 199.630 ;
        RECT 65.805 199.290 66.095 199.335 ;
        RECT 66.710 199.290 67.030 199.350 ;
        RECT 65.805 199.150 67.030 199.290 ;
        RECT 65.805 199.105 66.095 199.150 ;
        RECT 66.710 199.090 67.030 199.150 ;
        RECT 72.230 199.290 72.550 199.350 ;
        RECT 73.240 199.335 73.380 199.490 ;
        RECT 75.910 199.430 76.230 199.490 ;
        RECT 73.165 199.290 73.455 199.335 ;
        RECT 72.230 199.150 73.455 199.290 ;
        RECT 72.230 199.090 72.550 199.150 ;
        RECT 73.165 199.105 73.455 199.150 ;
        RECT 73.610 199.290 73.930 199.350 ;
        RECT 76.370 199.290 76.690 199.350 ;
        RECT 73.610 199.150 76.690 199.290 ;
        RECT 73.610 199.090 73.930 199.150 ;
        RECT 76.370 199.090 76.690 199.150 ;
        RECT 46.470 198.950 46.790 199.010 ;
        RECT 52.465 198.950 52.755 198.995 ;
        RECT 46.470 198.810 52.755 198.950 ;
        RECT 46.470 198.750 46.790 198.810 ;
        RECT 52.465 198.765 52.755 198.810 ;
        RECT 53.370 198.950 53.690 199.010 ;
        RECT 56.145 198.950 56.435 198.995 ;
        RECT 53.370 198.810 56.435 198.950 ;
        RECT 53.370 198.750 53.690 198.810 ;
        RECT 56.145 198.765 56.435 198.810 ;
        RECT 74.085 198.765 74.375 198.995 ;
        RECT 74.545 198.950 74.835 198.995 ;
        RECT 77.380 198.950 77.520 199.490 ;
        RECT 77.840 199.490 81.660 199.630 ;
        RECT 81.905 199.630 82.195 199.675 ;
        RECT 90.185 199.630 90.475 199.675 ;
        RECT 90.630 199.630 90.950 199.690 ;
        RECT 81.905 199.490 85.800 199.630 ;
        RECT 77.840 199.335 77.980 199.490 ;
        RECT 81.905 199.445 82.195 199.490 ;
        RECT 85.660 199.350 85.800 199.490 ;
        RECT 90.185 199.490 90.950 199.630 ;
        RECT 90.185 199.445 90.475 199.490 ;
        RECT 90.630 199.430 90.950 199.490 ;
        RECT 91.090 199.430 91.410 199.690 ;
        RECT 99.460 199.630 99.600 199.830 ;
        RECT 109.490 199.770 109.810 199.830 ;
        RECT 115.470 199.770 115.790 200.030 ;
        RECT 94.400 199.490 99.600 199.630 ;
        RECT 94.400 199.350 94.540 199.490 ;
        RECT 77.765 199.105 78.055 199.335 ;
        RECT 78.225 199.105 78.515 199.335 ;
        RECT 78.300 198.950 78.440 199.105 ;
        RECT 78.670 199.090 78.990 199.350 ;
        RECT 79.590 199.290 79.910 199.350 ;
        RECT 80.065 199.290 80.355 199.335 ;
        RECT 83.745 199.290 84.035 199.335 ;
        RECT 79.590 199.150 80.355 199.290 ;
        RECT 79.590 199.090 79.910 199.150 ;
        RECT 80.065 199.105 80.355 199.150 ;
        RECT 80.600 199.150 84.035 199.290 ;
        RECT 80.600 198.950 80.740 199.150 ;
        RECT 83.745 199.105 84.035 199.150 ;
        RECT 85.570 199.090 85.890 199.350 ;
        RECT 88.345 199.290 88.635 199.335 ;
        RECT 92.025 199.290 92.315 199.335 ;
        RECT 88.345 199.150 92.315 199.290 ;
        RECT 88.345 199.105 88.635 199.150 ;
        RECT 92.025 199.105 92.315 199.150 ;
        RECT 94.310 199.090 94.630 199.350 ;
        RECT 99.460 199.335 99.600 199.490 ;
        RECT 99.845 199.630 100.135 199.675 ;
        RECT 102.245 199.630 102.535 199.675 ;
        RECT 105.485 199.630 106.135 199.675 ;
        RECT 99.845 199.490 106.135 199.630 ;
        RECT 109.580 199.630 109.720 199.770 ;
        RECT 109.580 199.490 116.160 199.630 ;
        RECT 99.845 199.445 100.135 199.490 ;
        RECT 102.245 199.445 102.835 199.490 ;
        RECT 105.485 199.445 106.135 199.490 ;
        RECT 96.165 199.105 96.455 199.335 ;
        RECT 99.385 199.105 99.675 199.335 ;
        RECT 102.545 199.130 102.835 199.445 ;
        RECT 103.625 199.290 103.915 199.335 ;
        RECT 107.205 199.290 107.495 199.335 ;
        RECT 109.040 199.290 109.330 199.335 ;
        RECT 103.625 199.150 109.330 199.290 ;
        RECT 103.625 199.105 103.915 199.150 ;
        RECT 107.205 199.105 107.495 199.150 ;
        RECT 109.040 199.105 109.330 199.150 ;
        RECT 109.505 199.290 109.795 199.335 ;
        RECT 110.870 199.290 111.190 199.350 ;
        RECT 109.505 199.150 111.190 199.290 ;
        RECT 109.505 199.105 109.795 199.150 ;
        RECT 74.545 198.810 77.060 198.950 ;
        RECT 77.380 198.810 80.740 198.950 ;
        RECT 81.320 198.950 81.610 198.995 ;
        RECT 82.350 198.950 82.670 199.010 ;
        RECT 81.320 198.810 82.670 198.950 ;
        RECT 74.545 198.765 74.835 198.810 ;
        RECT 55.670 198.070 55.990 198.330 ;
        RECT 59.350 198.070 59.670 198.330 ;
        RECT 65.790 198.270 66.110 198.330 ;
        RECT 66.265 198.270 66.555 198.315 ;
        RECT 65.790 198.130 66.555 198.270 ;
        RECT 74.160 198.270 74.300 198.765 ;
        RECT 76.920 198.655 77.060 198.810 ;
        RECT 81.320 198.765 81.610 198.810 ;
        RECT 82.350 198.750 82.670 198.810 ;
        RECT 86.950 198.950 87.270 199.010 ;
        RECT 96.240 198.950 96.380 199.105 ;
        RECT 110.870 199.090 111.190 199.150 ;
        RECT 112.250 199.090 112.570 199.350 ;
        RECT 116.020 199.335 116.160 199.490 ;
        RECT 115.945 199.290 116.235 199.335 ;
        RECT 116.865 199.290 117.155 199.335 ;
        RECT 115.945 199.150 117.155 199.290 ;
        RECT 115.945 199.105 116.235 199.150 ;
        RECT 116.865 199.105 117.155 199.150 ;
        RECT 119.165 199.105 119.455 199.335 ;
        RECT 86.950 198.810 96.380 198.950 ;
        RECT 86.950 198.750 87.270 198.810 ;
        RECT 108.110 198.750 108.430 199.010 ;
        RECT 109.950 198.950 110.270 199.010 ;
        RECT 111.345 198.950 111.635 198.995 ;
        RECT 109.950 198.810 111.635 198.950 ;
        RECT 109.950 198.750 110.270 198.810 ;
        RECT 111.345 198.765 111.635 198.810 ;
        RECT 111.790 198.750 112.110 199.010 ;
        RECT 119.240 198.950 119.380 199.105 ;
        RECT 114.180 198.810 119.380 198.950 ;
        RECT 76.845 198.610 77.135 198.655 ;
        RECT 78.670 198.610 78.990 198.670 ;
        RECT 76.845 198.470 78.990 198.610 ;
        RECT 76.845 198.425 77.135 198.470 ;
        RECT 78.670 198.410 78.990 198.470 ;
        RECT 79.130 198.610 79.450 198.670 ;
        RECT 83.730 198.610 84.050 198.670 ;
        RECT 91.090 198.610 91.410 198.670 ;
        RECT 114.180 198.655 114.320 198.810 ;
        RECT 92.945 198.610 93.235 198.655 ;
        RECT 79.130 198.470 93.235 198.610 ;
        RECT 79.130 198.410 79.450 198.470 ;
        RECT 83.730 198.410 84.050 198.470 ;
        RECT 91.090 198.410 91.410 198.470 ;
        RECT 92.945 198.425 93.235 198.470 ;
        RECT 103.625 198.610 103.915 198.655 ;
        RECT 106.745 198.610 107.035 198.655 ;
        RECT 108.635 198.610 108.925 198.655 ;
        RECT 103.625 198.470 108.925 198.610 ;
        RECT 103.625 198.425 103.915 198.470 ;
        RECT 106.745 198.425 107.035 198.470 ;
        RECT 108.635 198.425 108.925 198.470 ;
        RECT 114.105 198.425 114.395 198.655 ;
        RECT 79.220 198.270 79.360 198.410 ;
        RECT 74.160 198.130 79.360 198.270 ;
        RECT 65.790 198.070 66.110 198.130 ;
        RECT 66.265 198.085 66.555 198.130 ;
        RECT 80.510 198.070 80.830 198.330 ;
        RECT 86.490 198.270 86.810 198.330 ;
        RECT 89.265 198.270 89.555 198.315 ;
        RECT 86.490 198.130 89.555 198.270 ;
        RECT 86.490 198.070 86.810 198.130 ;
        RECT 89.265 198.085 89.555 198.130 ;
        RECT 97.085 198.270 97.375 198.315 ;
        RECT 97.990 198.270 98.310 198.330 ;
        RECT 97.085 198.130 98.310 198.270 ;
        RECT 97.085 198.085 97.375 198.130 ;
        RECT 97.990 198.070 98.310 198.130 ;
        RECT 100.750 198.070 101.070 198.330 ;
        RECT 117.325 198.270 117.615 198.315 ;
        RECT 117.770 198.270 118.090 198.330 ;
        RECT 117.325 198.130 118.090 198.270 ;
        RECT 117.325 198.085 117.615 198.130 ;
        RECT 117.770 198.070 118.090 198.130 ;
        RECT 120.085 198.270 120.375 198.315 ;
        RECT 121.450 198.270 121.770 198.330 ;
        RECT 120.085 198.130 121.770 198.270 ;
        RECT 120.085 198.085 120.375 198.130 ;
        RECT 121.450 198.070 121.770 198.130 ;
        RECT 29.840 197.450 127.820 197.930 ;
        RECT 84.190 197.250 84.510 197.310 ;
        RECT 84.190 197.110 85.340 197.250 ;
        RECT 84.190 197.050 84.510 197.110 ;
        RECT 66.710 196.910 67.030 196.970 ;
        RECT 58.520 196.770 67.030 196.910 ;
        RECT 55.210 196.570 55.530 196.630 ;
        RECT 58.520 196.570 58.660 196.770 ;
        RECT 66.710 196.710 67.030 196.770 ;
        RECT 67.645 196.725 67.935 196.955 ;
        RECT 78.670 196.910 78.990 196.970 ;
        RECT 81.890 196.910 82.210 196.970 ;
        RECT 84.650 196.910 84.970 196.970 ;
        RECT 78.670 196.770 84.970 196.910 ;
        RECT 85.200 196.910 85.340 197.110 ;
        RECT 86.490 197.050 86.810 197.310 ;
        RECT 87.410 197.050 87.730 197.310 ;
        RECT 105.810 197.250 106.130 197.310 ;
        RECT 100.840 197.110 106.130 197.250 ;
        RECT 87.870 196.910 88.190 196.970 ;
        RECT 89.265 196.910 89.555 196.955 ;
        RECT 90.630 196.910 90.950 196.970 ;
        RECT 85.200 196.770 86.720 196.910 ;
        RECT 53.460 196.430 58.660 196.570 ;
        RECT 49.705 196.230 49.995 196.275 ;
        RECT 50.150 196.230 50.470 196.290 ;
        RECT 49.705 196.090 50.470 196.230 ;
        RECT 49.705 196.045 49.995 196.090 ;
        RECT 50.150 196.030 50.470 196.090 ;
        RECT 51.990 196.030 52.310 196.290 ;
        RECT 53.460 196.275 53.600 196.430 ;
        RECT 55.210 196.370 55.530 196.430 ;
        RECT 53.385 196.045 53.675 196.275 ;
        RECT 54.305 196.230 54.595 196.275 ;
        RECT 56.590 196.230 56.910 196.290 ;
        RECT 54.305 196.090 56.910 196.230 ;
        RECT 54.305 196.045 54.595 196.090 ;
        RECT 56.590 196.030 56.910 196.090 ;
        RECT 57.065 196.230 57.355 196.275 ;
        RECT 57.970 196.230 58.290 196.290 ;
        RECT 58.520 196.275 58.660 196.430 ;
        RECT 60.730 196.570 61.050 196.630 ;
        RECT 64.425 196.570 64.715 196.615 ;
        RECT 60.730 196.430 64.715 196.570 ;
        RECT 60.730 196.370 61.050 196.430 ;
        RECT 64.425 196.385 64.715 196.430 ;
        RECT 57.065 196.090 58.290 196.230 ;
        RECT 57.065 196.045 57.355 196.090 ;
        RECT 57.970 196.030 58.290 196.090 ;
        RECT 58.445 196.045 58.735 196.275 ;
        RECT 58.905 196.230 59.195 196.275 ;
        RECT 60.285 196.230 60.575 196.275 ;
        RECT 58.905 196.090 60.575 196.230 ;
        RECT 58.905 196.045 59.195 196.090 ;
        RECT 60.285 196.045 60.575 196.090 ;
        RECT 63.505 196.230 63.795 196.275 ;
        RECT 63.950 196.230 64.270 196.290 ;
        RECT 63.505 196.090 64.270 196.230 ;
        RECT 67.720 196.230 67.860 196.725 ;
        RECT 78.670 196.710 78.990 196.770 ;
        RECT 81.890 196.710 82.210 196.770 ;
        RECT 84.650 196.710 84.970 196.770 ;
        RECT 85.570 196.370 85.890 196.630 ;
        RECT 68.105 196.230 68.395 196.275 ;
        RECT 67.720 196.090 68.395 196.230 ;
        RECT 63.505 196.045 63.795 196.090 ;
        RECT 63.950 196.030 64.270 196.090 ;
        RECT 68.105 196.045 68.395 196.090 ;
        RECT 81.905 196.230 82.195 196.275 ;
        RECT 85.660 196.230 85.800 196.370 ;
        RECT 81.905 196.090 85.800 196.230 ;
        RECT 81.905 196.045 82.195 196.090 ;
        RECT 59.350 195.890 59.670 195.950 ;
        RECT 65.805 195.890 66.095 195.935 ;
        RECT 59.350 195.750 66.095 195.890 ;
        RECT 59.350 195.690 59.670 195.750 ;
        RECT 65.805 195.705 66.095 195.750 ;
        RECT 80.985 195.890 81.275 195.935 ;
        RECT 83.270 195.890 83.590 195.950 ;
        RECT 80.985 195.750 83.590 195.890 ;
        RECT 80.985 195.705 81.275 195.750 ;
        RECT 83.270 195.690 83.590 195.750 ;
        RECT 84.190 195.890 84.510 195.950 ;
        RECT 84.665 195.890 84.955 195.935 ;
        RECT 84.190 195.750 84.955 195.890 ;
        RECT 84.190 195.690 84.510 195.750 ;
        RECT 84.665 195.705 84.955 195.750 ;
        RECT 85.585 195.890 85.875 195.935 ;
        RECT 86.030 195.890 86.350 195.950 ;
        RECT 85.585 195.750 86.350 195.890 ;
        RECT 86.580 195.935 86.720 196.770 ;
        RECT 87.870 196.770 90.950 196.910 ;
        RECT 87.870 196.710 88.190 196.770 ;
        RECT 89.265 196.725 89.555 196.770 ;
        RECT 90.630 196.710 90.950 196.770 ;
        RECT 91.090 196.570 91.410 196.630 ;
        RECT 98.005 196.570 98.295 196.615 ;
        RECT 100.840 196.570 100.980 197.110 ;
        RECT 105.810 197.050 106.130 197.110 ;
        RECT 106.745 197.250 107.035 197.295 ;
        RECT 108.110 197.250 108.430 197.310 ;
        RECT 106.745 197.110 108.430 197.250 ;
        RECT 106.745 197.065 107.035 197.110 ;
        RECT 108.110 197.050 108.430 197.110 ;
        RECT 119.610 197.250 119.930 197.310 ;
        RECT 119.610 197.110 123.060 197.250 ;
        RECT 119.610 197.050 119.930 197.110 ;
        RECT 101.225 196.725 101.515 196.955 ;
        RECT 91.090 196.430 100.980 196.570 ;
        RECT 91.090 196.370 91.410 196.430 ;
        RECT 98.005 196.385 98.295 196.430 ;
        RECT 92.485 196.230 92.775 196.275 ;
        RECT 93.390 196.230 93.710 196.290 ;
        RECT 92.485 196.090 93.710 196.230 ;
        RECT 92.485 196.045 92.775 196.090 ;
        RECT 93.390 196.030 93.710 196.090 ;
        RECT 94.325 196.230 94.615 196.275 ;
        RECT 100.750 196.230 101.070 196.290 ;
        RECT 94.325 196.090 101.070 196.230 ;
        RECT 101.300 196.230 101.440 196.725 ;
        RECT 105.900 196.570 106.040 197.050 ;
        RECT 116.965 196.910 117.255 196.955 ;
        RECT 120.085 196.910 120.375 196.955 ;
        RECT 121.975 196.910 122.265 196.955 ;
        RECT 116.965 196.770 122.265 196.910 ;
        RECT 116.965 196.725 117.255 196.770 ;
        RECT 120.085 196.725 120.375 196.770 ;
        RECT 121.975 196.725 122.265 196.770 ;
        RECT 109.950 196.570 110.270 196.630 ;
        RECT 110.425 196.570 110.715 196.615 ;
        RECT 105.900 196.430 110.715 196.570 ;
        RECT 109.950 196.370 110.270 196.430 ;
        RECT 110.425 196.385 110.715 196.430 ;
        RECT 111.345 196.570 111.635 196.615 ;
        RECT 112.250 196.570 112.570 196.630 ;
        RECT 111.345 196.430 112.570 196.570 ;
        RECT 111.345 196.385 111.635 196.430 ;
        RECT 105.825 196.230 106.115 196.275 ;
        RECT 101.300 196.090 106.115 196.230 ;
        RECT 94.325 196.045 94.615 196.090 ;
        RECT 100.750 196.030 101.070 196.090 ;
        RECT 105.825 196.045 106.115 196.090 ;
        RECT 108.585 196.230 108.875 196.275 ;
        RECT 109.030 196.230 109.350 196.290 ;
        RECT 108.585 196.090 109.350 196.230 ;
        RECT 110.500 196.230 110.640 196.385 ;
        RECT 112.250 196.370 112.570 196.430 ;
        RECT 121.450 196.370 121.770 196.630 ;
        RECT 122.920 196.615 123.060 197.110 ;
        RECT 122.845 196.570 123.135 196.615 ;
        RECT 124.670 196.570 124.990 196.630 ;
        RECT 122.845 196.430 124.990 196.570 ;
        RECT 122.845 196.385 123.135 196.430 ;
        RECT 124.670 196.370 124.990 196.430 ;
        RECT 110.500 196.090 112.480 196.230 ;
        RECT 108.585 196.045 108.875 196.090 ;
        RECT 109.030 196.030 109.350 196.090 ;
        RECT 112.340 195.950 112.480 196.090 ;
        RECT 86.580 195.750 86.875 195.935 ;
        RECT 85.585 195.705 85.875 195.750 ;
        RECT 86.030 195.690 86.350 195.750 ;
        RECT 86.585 195.705 86.875 195.750 ;
        RECT 88.345 195.705 88.635 195.935 ;
        RECT 91.550 195.890 91.870 195.950 ;
        RECT 97.085 195.890 97.375 195.935 ;
        RECT 98.925 195.890 99.215 195.935 ;
        RECT 111.805 195.890 112.095 195.935 ;
        RECT 91.550 195.750 93.620 195.890 ;
        RECT 46.010 195.550 46.330 195.610 ;
        RECT 48.785 195.550 49.075 195.595 ;
        RECT 46.010 195.410 49.075 195.550 ;
        RECT 46.010 195.350 46.330 195.410 ;
        RECT 48.785 195.365 49.075 195.410 ;
        RECT 49.230 195.550 49.550 195.610 ;
        RECT 51.085 195.550 51.375 195.595 ;
        RECT 49.230 195.410 51.375 195.550 ;
        RECT 49.230 195.350 49.550 195.410 ;
        RECT 51.085 195.365 51.375 195.410 ;
        RECT 52.910 195.350 53.230 195.610 ;
        RECT 56.130 195.550 56.450 195.610 ;
        RECT 57.985 195.550 58.275 195.595 ;
        RECT 56.130 195.410 58.275 195.550 ;
        RECT 56.130 195.350 56.450 195.410 ;
        RECT 57.985 195.365 58.275 195.410 ;
        RECT 59.825 195.550 60.115 195.595 ;
        RECT 61.190 195.550 61.510 195.610 ;
        RECT 59.825 195.410 61.510 195.550 ;
        RECT 59.825 195.365 60.115 195.410 ;
        RECT 61.190 195.350 61.510 195.410 ;
        RECT 65.330 195.350 65.650 195.610 ;
        RECT 69.025 195.550 69.315 195.595 ;
        RECT 70.850 195.550 71.170 195.610 ;
        RECT 69.025 195.410 71.170 195.550 ;
        RECT 69.025 195.365 69.315 195.410 ;
        RECT 70.850 195.350 71.170 195.410 ;
        RECT 82.350 195.550 82.670 195.610 ;
        RECT 88.420 195.550 88.560 195.705 ;
        RECT 91.550 195.690 91.870 195.750 ;
        RECT 82.350 195.410 88.560 195.550 ;
        RECT 82.350 195.350 82.670 195.410 ;
        RECT 92.930 195.350 93.250 195.610 ;
        RECT 93.480 195.550 93.620 195.750 ;
        RECT 97.085 195.750 112.095 195.890 ;
        RECT 97.085 195.705 97.375 195.750 ;
        RECT 98.925 195.705 99.215 195.750 ;
        RECT 111.805 195.705 112.095 195.750 ;
        RECT 112.250 195.690 112.570 195.950 ;
        RECT 115.885 195.935 116.175 196.250 ;
        RECT 116.965 196.230 117.255 196.275 ;
        RECT 120.545 196.230 120.835 196.275 ;
        RECT 122.380 196.230 122.670 196.275 ;
        RECT 116.965 196.090 122.670 196.230 ;
        RECT 116.965 196.045 117.255 196.090 ;
        RECT 120.545 196.045 120.835 196.090 ;
        RECT 122.380 196.045 122.670 196.090 ;
        RECT 115.585 195.890 116.175 195.935 ;
        RECT 117.770 195.890 118.090 195.950 ;
        RECT 118.825 195.890 119.475 195.935 ;
        RECT 115.585 195.750 119.475 195.890 ;
        RECT 115.585 195.705 115.875 195.750 ;
        RECT 117.770 195.690 118.090 195.750 ;
        RECT 118.825 195.705 119.475 195.750 ;
        RECT 99.385 195.550 99.675 195.595 ;
        RECT 93.480 195.410 99.675 195.550 ;
        RECT 99.385 195.365 99.675 195.410 ;
        RECT 109.505 195.550 109.795 195.595 ;
        RECT 109.950 195.550 110.270 195.610 ;
        RECT 109.505 195.410 110.270 195.550 ;
        RECT 109.505 195.365 109.795 195.410 ;
        RECT 109.950 195.350 110.270 195.410 ;
        RECT 113.170 195.550 113.490 195.610 ;
        RECT 113.645 195.550 113.935 195.595 ;
        RECT 113.170 195.410 113.935 195.550 ;
        RECT 113.170 195.350 113.490 195.410 ;
        RECT 113.645 195.365 113.935 195.410 ;
        RECT 114.105 195.550 114.395 195.595 ;
        RECT 115.010 195.550 115.330 195.610 ;
        RECT 114.105 195.410 115.330 195.550 ;
        RECT 114.105 195.365 114.395 195.410 ;
        RECT 115.010 195.350 115.330 195.410 ;
        RECT 29.840 194.730 127.820 195.210 ;
        RECT 75.910 194.530 76.230 194.590 ;
        RECT 77.750 194.530 78.070 194.590 ;
        RECT 84.190 194.530 84.510 194.590 ;
        RECT 93.390 194.530 93.710 194.590 ;
        RECT 97.530 194.530 97.850 194.590 ;
        RECT 75.910 194.390 80.280 194.530 ;
        RECT 75.910 194.330 76.230 194.390 ;
        RECT 77.750 194.330 78.070 194.390 ;
        RECT 46.010 193.990 46.330 194.250 ;
        RECT 48.305 194.190 48.955 194.235 ;
        RECT 51.905 194.190 52.195 194.235 ;
        RECT 52.910 194.190 53.230 194.250 ;
        RECT 48.305 194.050 53.230 194.190 ;
        RECT 48.305 194.005 48.955 194.050 ;
        RECT 51.605 194.005 52.195 194.050 ;
        RECT 35.430 193.850 35.750 193.910 ;
        RECT 43.265 193.850 43.555 193.895 ;
        RECT 35.430 193.710 43.555 193.850 ;
        RECT 35.430 193.650 35.750 193.710 ;
        RECT 43.265 193.665 43.555 193.710 ;
        RECT 45.110 193.850 45.400 193.895 ;
        RECT 46.945 193.850 47.235 193.895 ;
        RECT 50.525 193.850 50.815 193.895 ;
        RECT 45.110 193.710 50.815 193.850 ;
        RECT 45.110 193.665 45.400 193.710 ;
        RECT 46.945 193.665 47.235 193.710 ;
        RECT 50.525 193.665 50.815 193.710 ;
        RECT 51.605 193.690 51.895 194.005 ;
        RECT 52.910 193.990 53.230 194.050 ;
        RECT 55.325 194.190 55.615 194.235 ;
        RECT 56.130 194.190 56.450 194.250 ;
        RECT 58.565 194.190 59.215 194.235 ;
        RECT 55.325 194.050 59.215 194.190 ;
        RECT 55.325 194.005 55.915 194.050 ;
        RECT 55.625 193.690 55.915 194.005 ;
        RECT 56.130 193.990 56.450 194.050 ;
        RECT 58.565 194.005 59.215 194.050 ;
        RECT 61.190 193.990 61.510 194.250 ;
        RECT 64.985 194.190 65.275 194.235 ;
        RECT 65.790 194.190 66.110 194.250 ;
        RECT 68.225 194.190 68.875 194.235 ;
        RECT 64.985 194.050 68.875 194.190 ;
        RECT 64.985 194.005 65.575 194.050 ;
        RECT 56.705 193.850 56.995 193.895 ;
        RECT 60.285 193.850 60.575 193.895 ;
        RECT 62.120 193.850 62.410 193.895 ;
        RECT 56.705 193.710 62.410 193.850 ;
        RECT 56.705 193.665 56.995 193.710 ;
        RECT 60.285 193.665 60.575 193.710 ;
        RECT 62.120 193.665 62.410 193.710 ;
        RECT 65.285 193.690 65.575 194.005 ;
        RECT 65.790 193.990 66.110 194.050 ;
        RECT 68.225 194.005 68.875 194.050 ;
        RECT 70.850 193.990 71.170 194.250 ;
        RECT 71.310 194.190 71.630 194.250 ;
        RECT 80.140 194.190 80.280 194.390 ;
        RECT 82.900 194.390 84.510 194.530 ;
        RECT 82.900 194.190 83.040 194.390 ;
        RECT 84.190 194.330 84.510 194.390 ;
        RECT 92.560 194.390 104.660 194.530 ;
        RECT 87.870 194.190 88.190 194.250 ;
        RECT 71.310 194.050 79.820 194.190 ;
        RECT 71.310 193.990 71.630 194.050 ;
        RECT 66.365 193.850 66.655 193.895 ;
        RECT 69.945 193.850 70.235 193.895 ;
        RECT 71.780 193.850 72.070 193.895 ;
        RECT 66.365 193.710 72.070 193.850 ;
        RECT 66.365 193.665 66.655 193.710 ;
        RECT 69.945 193.665 70.235 193.710 ;
        RECT 71.780 193.665 72.070 193.710 ;
        RECT 73.150 193.850 73.470 193.910 ;
        RECT 73.625 193.850 73.915 193.895 ;
        RECT 76.845 193.850 77.135 193.895 ;
        RECT 73.150 193.710 73.915 193.850 ;
        RECT 73.150 193.650 73.470 193.710 ;
        RECT 73.625 193.665 73.915 193.710 ;
        RECT 76.000 193.710 77.135 193.850 ;
        RECT 44.645 193.510 44.935 193.555 ;
        RECT 49.690 193.510 50.010 193.570 ;
        RECT 44.645 193.370 50.010 193.510 ;
        RECT 44.645 193.325 44.935 193.370 ;
        RECT 49.690 193.310 50.010 193.370 ;
        RECT 61.190 193.510 61.510 193.570 ;
        RECT 62.585 193.510 62.875 193.555 ;
        RECT 72.245 193.510 72.535 193.555 ;
        RECT 75.450 193.510 75.770 193.570 ;
        RECT 61.190 193.370 75.770 193.510 ;
        RECT 61.190 193.310 61.510 193.370 ;
        RECT 62.585 193.325 62.875 193.370 ;
        RECT 72.245 193.325 72.535 193.370 ;
        RECT 75.450 193.310 75.770 193.370 ;
        RECT 45.515 193.170 45.805 193.215 ;
        RECT 47.405 193.170 47.695 193.215 ;
        RECT 50.525 193.170 50.815 193.215 ;
        RECT 53.845 193.170 54.135 193.215 ;
        RECT 45.515 193.030 50.815 193.170 ;
        RECT 45.515 192.985 45.805 193.030 ;
        RECT 47.405 192.985 47.695 193.030 ;
        RECT 50.525 192.985 50.815 193.030 ;
        RECT 53.000 193.030 54.135 193.170 ;
        RECT 43.710 192.630 44.030 192.890 ;
        RECT 46.010 192.830 46.330 192.890 ;
        RECT 53.000 192.830 53.140 193.030 ;
        RECT 53.845 192.985 54.135 193.030 ;
        RECT 56.705 193.170 56.995 193.215 ;
        RECT 59.825 193.170 60.115 193.215 ;
        RECT 61.715 193.170 62.005 193.215 ;
        RECT 56.705 193.030 62.005 193.170 ;
        RECT 56.705 192.985 56.995 193.030 ;
        RECT 59.825 192.985 60.115 193.030 ;
        RECT 61.715 192.985 62.005 193.030 ;
        RECT 66.365 193.170 66.655 193.215 ;
        RECT 69.485 193.170 69.775 193.215 ;
        RECT 71.375 193.170 71.665 193.215 ;
        RECT 66.365 193.030 71.665 193.170 ;
        RECT 66.365 192.985 66.655 193.030 ;
        RECT 69.485 192.985 69.775 193.030 ;
        RECT 71.375 192.985 71.665 193.030 ;
        RECT 74.545 193.170 74.835 193.215 ;
        RECT 74.990 193.170 75.310 193.230 ;
        RECT 74.545 193.030 75.310 193.170 ;
        RECT 76.000 193.170 76.140 193.710 ;
        RECT 76.845 193.665 77.135 193.710 ;
        RECT 77.290 193.650 77.610 193.910 ;
        RECT 77.750 193.650 78.070 193.910 ;
        RECT 79.680 193.895 79.820 194.050 ;
        RECT 80.140 194.050 83.040 194.190 ;
        RECT 80.140 193.895 80.280 194.050 ;
        RECT 79.605 193.665 79.895 193.895 ;
        RECT 80.065 193.665 80.355 193.895 ;
        RECT 80.525 193.850 80.815 193.895 ;
        RECT 81.430 193.850 81.750 193.910 ;
        RECT 82.900 193.895 83.040 194.050 ;
        RECT 83.820 194.050 88.190 194.190 ;
        RECT 83.820 193.895 83.960 194.050 ;
        RECT 87.870 193.990 88.190 194.050 ;
        RECT 80.525 193.710 81.750 193.850 ;
        RECT 80.525 193.665 80.815 193.710 ;
        RECT 81.430 193.650 81.750 193.710 ;
        RECT 82.810 193.665 83.100 193.895 ;
        RECT 83.745 193.665 84.035 193.895 ;
        RECT 76.385 193.510 76.675 193.555 ;
        RECT 80.985 193.510 81.275 193.555 ;
        RECT 81.890 193.510 82.210 193.570 ;
        RECT 83.285 193.510 83.575 193.555 ;
        RECT 76.385 193.370 83.575 193.510 ;
        RECT 76.385 193.325 76.675 193.370 ;
        RECT 80.140 193.230 80.280 193.370 ;
        RECT 80.985 193.325 81.275 193.370 ;
        RECT 81.890 193.310 82.210 193.370 ;
        RECT 83.285 193.325 83.575 193.370 ;
        RECT 79.130 193.170 79.450 193.230 ;
        RECT 76.000 193.030 79.450 193.170 ;
        RECT 74.545 192.985 74.835 193.030 ;
        RECT 46.010 192.690 53.140 192.830 ;
        RECT 46.010 192.630 46.330 192.690 ;
        RECT 53.370 192.630 53.690 192.890 ;
        RECT 53.920 192.830 54.060 192.985 ;
        RECT 74.990 192.970 75.310 193.030 ;
        RECT 79.130 192.970 79.450 193.030 ;
        RECT 80.050 192.970 80.370 193.230 ;
        RECT 81.430 193.170 81.750 193.230 ;
        RECT 83.820 193.170 83.960 193.665 ;
        RECT 84.190 193.650 84.510 193.910 ;
        RECT 89.265 193.850 89.555 193.895 ;
        RECT 92.560 193.850 92.700 194.390 ;
        RECT 93.390 194.330 93.710 194.390 ;
        RECT 97.530 194.330 97.850 194.390 ;
        RECT 92.930 194.235 93.250 194.250 ;
        RECT 92.880 194.190 93.250 194.235 ;
        RECT 96.140 194.190 96.430 194.235 ;
        RECT 92.880 194.050 96.430 194.190 ;
        RECT 92.880 194.005 93.250 194.050 ;
        RECT 96.140 194.005 96.430 194.050 ;
        RECT 97.060 194.190 97.350 194.235 ;
        RECT 98.920 194.190 99.210 194.235 ;
        RECT 97.060 194.050 99.210 194.190 ;
        RECT 97.060 194.005 97.350 194.050 ;
        RECT 98.920 194.005 99.210 194.050 ;
        RECT 92.930 193.990 93.250 194.005 ;
        RECT 89.265 193.710 92.700 193.850 ;
        RECT 94.740 193.850 95.030 193.895 ;
        RECT 97.060 193.850 97.275 194.005 ;
        RECT 94.740 193.710 97.275 193.850 ;
        RECT 89.265 193.665 89.555 193.710 ;
        RECT 94.740 193.665 95.030 193.710 ;
        RECT 97.990 193.650 98.310 193.910 ;
        RECT 104.520 193.895 104.660 194.390 ;
        RECT 109.030 194.330 109.350 194.590 ;
        RECT 114.090 194.330 114.410 194.590 ;
        RECT 111.790 194.190 112.110 194.250 ;
        RECT 115.025 194.190 115.315 194.235 ;
        RECT 111.790 194.050 115.315 194.190 ;
        RECT 111.790 193.990 112.110 194.050 ;
        RECT 115.025 194.005 115.315 194.050 ;
        RECT 104.445 193.665 104.735 193.895 ;
        RECT 106.270 193.650 106.590 193.910 ;
        RECT 113.170 193.650 113.490 193.910 ;
        RECT 98.450 193.510 98.770 193.570 ;
        RECT 99.845 193.510 100.135 193.555 ;
        RECT 110.870 193.510 111.190 193.570 ;
        RECT 98.450 193.370 111.190 193.510 ;
        RECT 98.450 193.310 98.770 193.370 ;
        RECT 99.845 193.325 100.135 193.370 ;
        RECT 110.870 193.310 111.190 193.370 ;
        RECT 112.710 193.310 113.030 193.570 ;
        RECT 115.010 193.510 115.330 193.570 ;
        RECT 117.785 193.510 118.075 193.555 ;
        RECT 115.010 193.370 118.075 193.510 ;
        RECT 115.010 193.310 115.330 193.370 ;
        RECT 117.785 193.325 118.075 193.370 ;
        RECT 81.430 193.030 83.960 193.170 ;
        RECT 85.570 193.170 85.890 193.230 ;
        RECT 90.875 193.170 91.165 193.215 ;
        RECT 91.550 193.170 91.870 193.230 ;
        RECT 85.570 193.030 91.870 193.170 ;
        RECT 81.430 192.970 81.750 193.030 ;
        RECT 85.570 192.970 85.890 193.030 ;
        RECT 90.875 192.985 91.165 193.030 ;
        RECT 91.550 192.970 91.870 193.030 ;
        RECT 94.740 193.170 95.030 193.215 ;
        RECT 97.520 193.170 97.810 193.215 ;
        RECT 99.380 193.170 99.670 193.215 ;
        RECT 94.740 193.030 99.670 193.170 ;
        RECT 94.740 192.985 95.030 193.030 ;
        RECT 97.520 192.985 97.810 193.030 ;
        RECT 99.380 192.985 99.670 193.030 ;
        RECT 58.890 192.830 59.210 192.890 ;
        RECT 53.920 192.690 59.210 192.830 ;
        RECT 58.890 192.630 59.210 192.690 ;
        RECT 60.270 192.830 60.590 192.890 ;
        RECT 63.505 192.830 63.795 192.875 ;
        RECT 71.770 192.830 72.090 192.890 ;
        RECT 60.270 192.690 72.090 192.830 ;
        RECT 60.270 192.630 60.590 192.690 ;
        RECT 63.505 192.645 63.795 192.690 ;
        RECT 71.770 192.630 72.090 192.690 ;
        RECT 73.610 192.830 73.930 192.890 ;
        RECT 75.465 192.830 75.755 192.875 ;
        RECT 73.610 192.690 75.755 192.830 ;
        RECT 73.610 192.630 73.930 192.690 ;
        RECT 75.465 192.645 75.755 192.690 ;
        RECT 78.670 192.630 78.990 192.890 ;
        RECT 81.890 192.630 82.210 192.890 ;
        RECT 89.710 192.630 90.030 192.890 ;
        RECT 104.890 192.630 105.210 192.890 ;
        RECT 109.490 192.630 109.810 192.890 ;
        RECT 29.840 192.010 127.820 192.490 ;
        RECT 50.150 191.810 50.470 191.870 ;
        RECT 50.625 191.810 50.915 191.855 ;
        RECT 50.150 191.670 50.915 191.810 ;
        RECT 50.150 191.610 50.470 191.670 ;
        RECT 50.625 191.625 50.915 191.670 ;
        RECT 56.590 191.610 56.910 191.870 ;
        RECT 58.890 191.810 59.210 191.870 ;
        RECT 63.950 191.810 64.270 191.870 ;
        RECT 64.425 191.810 64.715 191.855 ;
        RECT 58.890 191.670 62.340 191.810 ;
        RECT 58.890 191.610 59.210 191.670 ;
        RECT 44.600 191.470 44.890 191.515 ;
        RECT 47.380 191.470 47.670 191.515 ;
        RECT 49.240 191.470 49.530 191.515 ;
        RECT 59.350 191.470 59.670 191.530 ;
        RECT 44.600 191.330 49.530 191.470 ;
        RECT 44.600 191.285 44.890 191.330 ;
        RECT 47.380 191.285 47.670 191.330 ;
        RECT 49.240 191.285 49.530 191.330 ;
        RECT 53.000 191.330 59.670 191.470 ;
        RECT 53.000 191.175 53.140 191.330 ;
        RECT 59.350 191.270 59.670 191.330 ;
        RECT 52.925 190.945 53.215 191.175 ;
        RECT 53.845 191.130 54.135 191.175 ;
        RECT 54.290 191.130 54.610 191.190 ;
        RECT 53.845 190.990 54.610 191.130 ;
        RECT 53.845 190.945 54.135 190.990 ;
        RECT 54.290 190.930 54.610 190.990 ;
        RECT 54.750 191.130 55.070 191.190 ;
        RECT 58.905 191.130 59.195 191.175 ;
        RECT 59.825 191.130 60.115 191.175 ;
        RECT 60.730 191.130 61.050 191.190 ;
        RECT 62.200 191.175 62.340 191.670 ;
        RECT 63.950 191.670 64.715 191.810 ;
        RECT 63.950 191.610 64.270 191.670 ;
        RECT 64.425 191.625 64.715 191.670 ;
        RECT 86.950 191.610 87.270 191.870 ;
        RECT 67.745 191.470 68.035 191.515 ;
        RECT 70.865 191.470 71.155 191.515 ;
        RECT 72.755 191.470 73.045 191.515 ;
        RECT 67.745 191.330 73.045 191.470 ;
        RECT 67.745 191.285 68.035 191.330 ;
        RECT 70.865 191.285 71.155 191.330 ;
        RECT 72.755 191.285 73.045 191.330 ;
        RECT 77.765 191.470 78.055 191.515 ;
        RECT 79.130 191.470 79.450 191.530 ;
        RECT 77.765 191.330 79.450 191.470 ;
        RECT 77.765 191.285 78.055 191.330 ;
        RECT 79.130 191.270 79.450 191.330 ;
        RECT 91.520 191.470 91.810 191.515 ;
        RECT 94.300 191.470 94.590 191.515 ;
        RECT 96.160 191.470 96.450 191.515 ;
        RECT 91.520 191.330 96.450 191.470 ;
        RECT 91.520 191.285 91.810 191.330 ;
        RECT 94.300 191.285 94.590 191.330 ;
        RECT 96.160 191.285 96.450 191.330 ;
        RECT 98.450 191.270 98.770 191.530 ;
        RECT 105.465 191.470 105.755 191.515 ;
        RECT 108.585 191.470 108.875 191.515 ;
        RECT 110.475 191.470 110.765 191.515 ;
        RECT 105.465 191.330 110.765 191.470 ;
        RECT 105.465 191.285 105.755 191.330 ;
        RECT 108.585 191.285 108.875 191.330 ;
        RECT 110.475 191.285 110.765 191.330 ;
        RECT 119.725 191.470 120.015 191.515 ;
        RECT 122.845 191.470 123.135 191.515 ;
        RECT 124.735 191.470 125.025 191.515 ;
        RECT 119.725 191.330 125.025 191.470 ;
        RECT 119.725 191.285 120.015 191.330 ;
        RECT 122.845 191.285 123.135 191.330 ;
        RECT 124.735 191.285 125.025 191.330 ;
        RECT 61.205 191.130 61.495 191.175 ;
        RECT 54.750 190.990 59.195 191.130 ;
        RECT 54.750 190.930 55.070 190.990 ;
        RECT 58.905 190.945 59.195 190.990 ;
        RECT 59.440 190.990 61.495 191.130 ;
        RECT 59.440 190.850 59.580 190.990 ;
        RECT 59.825 190.945 60.115 190.990 ;
        RECT 60.730 190.930 61.050 190.990 ;
        RECT 61.205 190.945 61.495 190.990 ;
        RECT 62.125 190.945 62.415 191.175 ;
        RECT 64.885 191.130 65.175 191.175 ;
        RECT 69.470 191.130 69.790 191.190 ;
        RECT 64.885 190.990 69.790 191.130 ;
        RECT 64.885 190.945 65.175 190.990 ;
        RECT 69.470 190.930 69.790 190.990 ;
        RECT 73.625 191.130 73.915 191.175 ;
        RECT 75.450 191.130 75.770 191.190 ;
        RECT 73.625 190.990 75.770 191.130 ;
        RECT 73.625 190.945 73.915 190.990 ;
        RECT 75.450 190.930 75.770 190.990 ;
        RECT 80.050 190.930 80.370 191.190 ;
        RECT 84.205 191.130 84.495 191.175 ;
        RECT 87.410 191.130 87.730 191.190 ;
        RECT 91.090 191.130 91.410 191.190 ;
        RECT 84.205 190.990 91.410 191.130 ;
        RECT 84.205 190.945 84.495 190.990 ;
        RECT 87.410 190.930 87.730 190.990 ;
        RECT 91.090 190.930 91.410 190.990 ;
        RECT 96.625 191.130 96.915 191.175 ;
        RECT 98.540 191.130 98.680 191.270 ;
        RECT 96.625 190.990 98.680 191.130 ;
        RECT 96.625 190.945 96.915 190.990 ;
        RECT 109.950 190.930 110.270 191.190 ;
        RECT 111.330 190.930 111.650 191.190 ;
        RECT 112.250 191.130 112.570 191.190 ;
        RECT 113.185 191.130 113.475 191.175 ;
        RECT 112.250 190.990 113.475 191.130 ;
        RECT 112.250 190.930 112.570 190.990 ;
        RECT 113.185 190.945 113.475 190.990 ;
        RECT 37.270 190.590 37.590 190.850 ;
        RECT 44.600 190.790 44.890 190.835 ;
        RECT 47.865 190.790 48.155 190.835 ;
        RECT 49.230 190.790 49.550 190.850 ;
        RECT 44.600 190.650 47.135 190.790 ;
        RECT 44.600 190.605 44.890 190.650 ;
        RECT 38.190 190.450 38.510 190.510 ;
        RECT 40.735 190.450 41.025 190.495 ;
        RECT 38.190 190.310 41.025 190.450 ;
        RECT 38.190 190.250 38.510 190.310 ;
        RECT 40.735 190.265 41.025 190.310 ;
        RECT 42.740 190.450 43.030 190.495 ;
        RECT 43.710 190.450 44.030 190.510 ;
        RECT 46.920 190.495 47.135 190.650 ;
        RECT 47.865 190.650 49.550 190.790 ;
        RECT 47.865 190.605 48.155 190.650 ;
        RECT 49.230 190.590 49.550 190.650 ;
        RECT 49.690 190.590 50.010 190.850 ;
        RECT 55.210 190.590 55.530 190.850 ;
        RECT 55.670 190.790 55.990 190.850 ;
        RECT 58.445 190.790 58.735 190.835 ;
        RECT 55.670 190.650 58.735 190.790 ;
        RECT 55.670 190.590 55.990 190.650 ;
        RECT 58.445 190.605 58.735 190.650 ;
        RECT 59.350 190.590 59.670 190.850 ;
        RECT 66.665 190.495 66.955 190.810 ;
        RECT 67.745 190.790 68.035 190.835 ;
        RECT 71.325 190.790 71.615 190.835 ;
        RECT 73.160 190.790 73.450 190.835 ;
        RECT 67.745 190.650 73.450 190.790 ;
        RECT 67.745 190.605 68.035 190.650 ;
        RECT 71.325 190.605 71.615 190.650 ;
        RECT 73.160 190.605 73.450 190.650 ;
        RECT 74.085 190.605 74.375 190.835 ;
        RECT 77.290 190.790 77.610 190.850 ;
        RECT 80.525 190.790 80.815 190.835 ;
        RECT 81.430 190.790 81.750 190.850 ;
        RECT 77.290 190.650 81.750 190.790 ;
        RECT 46.000 190.450 46.290 190.495 ;
        RECT 42.740 190.310 46.290 190.450 ;
        RECT 42.740 190.265 43.030 190.310 ;
        RECT 43.710 190.250 44.030 190.310 ;
        RECT 46.000 190.265 46.290 190.310 ;
        RECT 46.920 190.450 47.210 190.495 ;
        RECT 48.780 190.450 49.070 190.495 ;
        RECT 66.365 190.450 66.955 190.495 ;
        RECT 69.605 190.450 70.255 190.495 ;
        RECT 72.245 190.450 72.535 190.495 ;
        RECT 46.920 190.310 49.070 190.450 ;
        RECT 46.920 190.265 47.210 190.310 ;
        RECT 48.780 190.265 49.070 190.310 ;
        RECT 55.760 190.310 70.255 190.450 ;
        RECT 40.045 190.110 40.335 190.155 ;
        RECT 45.550 190.110 45.870 190.170 ;
        RECT 40.045 189.970 45.870 190.110 ;
        RECT 40.045 189.925 40.335 189.970 ;
        RECT 45.550 189.910 45.870 189.970 ;
        RECT 50.150 190.110 50.470 190.170 ;
        RECT 55.760 190.155 55.900 190.310 ;
        RECT 66.365 190.265 66.655 190.310 ;
        RECT 69.605 190.265 70.255 190.310 ;
        RECT 71.170 190.310 72.535 190.450 ;
        RECT 52.465 190.110 52.755 190.155 ;
        RECT 50.150 189.970 52.755 190.110 ;
        RECT 50.150 189.910 50.470 189.970 ;
        RECT 52.465 189.925 52.755 189.970 ;
        RECT 55.685 189.925 55.975 190.155 ;
        RECT 57.050 190.110 57.370 190.170 ;
        RECT 62.585 190.110 62.875 190.155 ;
        RECT 57.050 189.970 62.875 190.110 ;
        RECT 57.050 189.910 57.370 189.970 ;
        RECT 62.585 189.925 62.875 189.970 ;
        RECT 64.870 190.110 65.190 190.170 ;
        RECT 71.170 190.110 71.310 190.310 ;
        RECT 72.245 190.265 72.535 190.310 ;
        RECT 73.610 190.450 73.930 190.510 ;
        RECT 74.160 190.450 74.300 190.605 ;
        RECT 77.290 190.590 77.610 190.650 ;
        RECT 80.525 190.605 80.815 190.650 ;
        RECT 81.430 190.590 81.750 190.650 ;
        RECT 84.665 190.790 84.955 190.835 ;
        RECT 85.570 190.790 85.890 190.850 ;
        RECT 84.665 190.650 85.890 190.790 ;
        RECT 84.665 190.605 84.955 190.650 ;
        RECT 85.570 190.590 85.890 190.650 ;
        RECT 91.520 190.790 91.810 190.835 ;
        RECT 94.785 190.790 95.075 190.835 ;
        RECT 91.520 190.650 94.055 190.790 ;
        RECT 91.520 190.605 91.810 190.650 ;
        RECT 73.610 190.310 74.300 190.450 ;
        RECT 77.750 190.450 78.070 190.510 ;
        RECT 79.590 190.450 79.910 190.510 ;
        RECT 89.710 190.495 90.030 190.510 ;
        RECT 93.840 190.495 94.055 190.650 ;
        RECT 94.785 190.650 97.300 190.790 ;
        RECT 94.785 190.605 95.075 190.650 ;
        RECT 77.750 190.310 79.910 190.450 ;
        RECT 73.610 190.250 73.930 190.310 ;
        RECT 77.750 190.250 78.070 190.310 ;
        RECT 79.590 190.250 79.910 190.310 ;
        RECT 89.660 190.450 90.030 190.495 ;
        RECT 92.920 190.450 93.210 190.495 ;
        RECT 89.660 190.310 93.210 190.450 ;
        RECT 89.660 190.265 90.030 190.310 ;
        RECT 92.920 190.265 93.210 190.310 ;
        RECT 93.840 190.450 94.130 190.495 ;
        RECT 95.700 190.450 95.990 190.495 ;
        RECT 93.840 190.310 95.990 190.450 ;
        RECT 93.840 190.265 94.130 190.310 ;
        RECT 95.700 190.265 95.990 190.310 ;
        RECT 89.710 190.250 90.030 190.265 ;
        RECT 64.870 189.970 71.310 190.110 ;
        RECT 74.530 190.110 74.850 190.170 ;
        RECT 75.005 190.110 75.295 190.155 ;
        RECT 74.530 189.970 75.295 190.110 ;
        RECT 64.870 189.910 65.190 189.970 ;
        RECT 74.530 189.910 74.850 189.970 ;
        RECT 75.005 189.925 75.295 189.970 ;
        RECT 80.970 190.110 81.290 190.170 ;
        RECT 81.445 190.110 81.735 190.155 ;
        RECT 80.970 189.970 81.735 190.110 ;
        RECT 80.970 189.910 81.290 189.970 ;
        RECT 81.445 189.925 81.735 189.970 ;
        RECT 84.650 190.110 84.970 190.170 ;
        RECT 97.160 190.155 97.300 190.650 ;
        RECT 97.990 190.590 98.310 190.850 ;
        RECT 98.465 190.605 98.755 190.835 ;
        RECT 97.530 190.450 97.850 190.510 ;
        RECT 98.540 190.450 98.680 190.605 ;
        RECT 104.385 190.495 104.675 190.810 ;
        RECT 105.465 190.790 105.755 190.835 ;
        RECT 109.045 190.790 109.335 190.835 ;
        RECT 110.880 190.790 111.170 190.835 ;
        RECT 105.465 190.650 111.170 190.790 ;
        RECT 105.465 190.605 105.755 190.650 ;
        RECT 109.045 190.605 109.335 190.650 ;
        RECT 110.880 190.605 111.170 190.650 ;
        RECT 111.790 190.790 112.110 190.850 ;
        RECT 114.565 190.790 114.855 190.835 ;
        RECT 111.790 190.650 114.855 190.790 ;
        RECT 111.790 190.590 112.110 190.650 ;
        RECT 114.565 190.605 114.855 190.650 ;
        RECT 97.530 190.310 98.680 190.450 ;
        RECT 104.085 190.450 104.675 190.495 ;
        RECT 104.890 190.450 105.210 190.510 ;
        RECT 107.325 190.450 107.975 190.495 ;
        RECT 104.085 190.310 107.975 190.450 ;
        RECT 97.530 190.250 97.850 190.310 ;
        RECT 104.085 190.265 104.375 190.310 ;
        RECT 104.890 190.250 105.210 190.310 ;
        RECT 107.325 190.265 107.975 190.310 ;
        RECT 112.250 190.450 112.570 190.510 ;
        RECT 118.645 190.495 118.935 190.810 ;
        RECT 119.725 190.790 120.015 190.835 ;
        RECT 123.305 190.790 123.595 190.835 ;
        RECT 125.140 190.790 125.430 190.835 ;
        RECT 119.725 190.650 125.430 190.790 ;
        RECT 119.725 190.605 120.015 190.650 ;
        RECT 123.305 190.605 123.595 190.650 ;
        RECT 125.140 190.605 125.430 190.650 ;
        RECT 125.605 190.605 125.895 190.835 ;
        RECT 118.345 190.450 118.935 190.495 ;
        RECT 121.585 190.450 122.235 190.495 ;
        RECT 112.250 190.310 122.235 190.450 ;
        RECT 112.250 190.250 112.570 190.310 ;
        RECT 118.345 190.265 118.635 190.310 ;
        RECT 121.585 190.265 122.235 190.310 ;
        RECT 124.210 190.250 124.530 190.510 ;
        RECT 124.670 190.450 124.990 190.510 ;
        RECT 125.680 190.450 125.820 190.605 ;
        RECT 124.670 190.310 125.820 190.450 ;
        RECT 124.670 190.250 124.990 190.310 ;
        RECT 85.125 190.110 85.415 190.155 ;
        RECT 87.655 190.110 87.945 190.155 ;
        RECT 84.650 189.970 87.945 190.110 ;
        RECT 84.650 189.910 84.970 189.970 ;
        RECT 85.125 189.925 85.415 189.970 ;
        RECT 87.655 189.925 87.945 189.970 ;
        RECT 97.085 189.925 97.375 190.155 ;
        RECT 98.910 189.910 99.230 190.170 ;
        RECT 102.605 190.110 102.895 190.155 ;
        RECT 111.330 190.110 111.650 190.170 ;
        RECT 102.605 189.970 111.650 190.110 ;
        RECT 102.605 189.925 102.895 189.970 ;
        RECT 111.330 189.910 111.650 189.970 ;
        RECT 114.105 190.110 114.395 190.155 ;
        RECT 115.930 190.110 116.250 190.170 ;
        RECT 114.105 189.970 116.250 190.110 ;
        RECT 114.105 189.925 114.395 189.970 ;
        RECT 115.930 189.910 116.250 189.970 ;
        RECT 116.390 189.910 116.710 190.170 ;
        RECT 116.865 190.110 117.155 190.155 ;
        RECT 117.310 190.110 117.630 190.170 ;
        RECT 116.865 189.970 117.630 190.110 ;
        RECT 116.865 189.925 117.155 189.970 ;
        RECT 117.310 189.910 117.630 189.970 ;
        RECT 29.840 189.290 127.820 189.770 ;
        RECT 38.190 189.090 38.510 189.150 ;
        RECT 48.325 189.090 48.615 189.135 ;
        RECT 50.150 189.090 50.470 189.150 ;
        RECT 38.190 188.950 50.470 189.090 ;
        RECT 38.190 188.890 38.510 188.950 ;
        RECT 48.325 188.905 48.615 188.950 ;
        RECT 50.150 188.890 50.470 188.950 ;
        RECT 50.625 189.090 50.915 189.135 ;
        RECT 51.990 189.090 52.310 189.150 ;
        RECT 50.625 188.950 52.310 189.090 ;
        RECT 50.625 188.905 50.915 188.950 ;
        RECT 51.990 188.890 52.310 188.950 ;
        RECT 64.870 188.890 65.190 189.150 ;
        RECT 65.330 189.090 65.650 189.150 ;
        RECT 69.025 189.090 69.315 189.135 ;
        RECT 65.330 188.950 69.315 189.090 ;
        RECT 65.330 188.890 65.650 188.950 ;
        RECT 69.025 188.905 69.315 188.950 ;
        RECT 79.130 189.090 79.450 189.150 ;
        RECT 79.130 188.950 80.280 189.090 ;
        RECT 79.130 188.890 79.450 188.950 ;
        RECT 34.985 188.750 35.275 188.795 ;
        RECT 39.225 188.750 39.515 188.795 ;
        RECT 42.465 188.750 43.115 188.795 ;
        RECT 34.985 188.610 43.115 188.750 ;
        RECT 34.985 188.565 35.275 188.610 ;
        RECT 39.225 188.565 39.815 188.610 ;
        RECT 42.465 188.565 43.115 188.610 ;
        RECT 45.550 188.750 45.870 188.810 ;
        RECT 48.785 188.750 49.075 188.795 ;
        RECT 45.550 188.610 49.075 188.750 ;
        RECT 34.525 188.410 34.815 188.455 ;
        RECT 35.430 188.410 35.750 188.470 ;
        RECT 35.905 188.410 36.195 188.455 ;
        RECT 34.525 188.270 36.195 188.410 ;
        RECT 34.525 188.225 34.815 188.270 ;
        RECT 35.430 188.210 35.750 188.270 ;
        RECT 35.905 188.225 36.195 188.270 ;
        RECT 39.525 188.250 39.815 188.565 ;
        RECT 45.550 188.550 45.870 188.610 ;
        RECT 48.785 188.565 49.075 188.610 ;
        RECT 49.230 188.750 49.550 188.810 ;
        RECT 53.945 188.750 54.235 188.795 ;
        RECT 57.185 188.750 57.835 188.795 ;
        RECT 49.230 188.610 57.835 188.750 ;
        RECT 49.230 188.550 49.550 188.610 ;
        RECT 53.945 188.565 54.535 188.610 ;
        RECT 57.185 188.565 57.835 188.610 ;
        RECT 62.125 188.750 62.415 188.795 ;
        RECT 73.150 188.750 73.470 188.810 ;
        RECT 62.125 188.610 73.470 188.750 ;
        RECT 80.140 188.750 80.280 188.950 ;
        RECT 81.430 188.890 81.750 189.150 ;
        RECT 82.350 189.090 82.670 189.150 ;
        RECT 84.650 189.090 84.970 189.150 ;
        RECT 86.045 189.090 86.335 189.135 ;
        RECT 82.350 188.950 86.335 189.090 ;
        RECT 82.350 188.890 82.670 188.950 ;
        RECT 84.650 188.890 84.970 188.950 ;
        RECT 86.045 188.905 86.335 188.950 ;
        RECT 88.345 189.090 88.635 189.135 ;
        RECT 97.990 189.090 98.310 189.150 ;
        RECT 88.345 188.950 98.310 189.090 ;
        RECT 88.345 188.905 88.635 188.950 ;
        RECT 97.990 188.890 98.310 188.950 ;
        RECT 106.270 189.090 106.590 189.150 ;
        RECT 108.585 189.090 108.875 189.135 ;
        RECT 106.270 188.950 108.875 189.090 ;
        RECT 106.270 188.890 106.590 188.950 ;
        RECT 108.585 188.905 108.875 188.950 ;
        RECT 109.490 189.090 109.810 189.150 ;
        RECT 110.425 189.090 110.715 189.135 ;
        RECT 109.490 188.950 110.715 189.090 ;
        RECT 109.490 188.890 109.810 188.950 ;
        RECT 110.425 188.905 110.715 188.950 ;
        RECT 110.885 189.090 111.175 189.135 ;
        RECT 111.330 189.090 111.650 189.150 ;
        RECT 110.885 188.950 111.650 189.090 ;
        RECT 110.885 188.905 111.175 188.950 ;
        RECT 111.330 188.890 111.650 188.950 ;
        RECT 112.710 189.090 113.030 189.150 ;
        RECT 115.025 189.090 115.315 189.135 ;
        RECT 112.710 188.950 115.315 189.090 ;
        RECT 112.710 188.890 113.030 188.950 ;
        RECT 115.025 188.905 115.315 188.950 ;
        RECT 81.520 188.750 81.660 188.890 ;
        RECT 80.140 188.610 80.740 188.750 ;
        RECT 62.125 188.565 62.415 188.610 ;
        RECT 40.605 188.410 40.895 188.455 ;
        RECT 44.185 188.410 44.475 188.455 ;
        RECT 46.020 188.410 46.310 188.455 ;
        RECT 40.605 188.270 46.310 188.410 ;
        RECT 40.605 188.225 40.895 188.270 ;
        RECT 44.185 188.225 44.475 188.270 ;
        RECT 46.020 188.225 46.310 188.270 ;
        RECT 46.470 188.410 46.790 188.470 ;
        RECT 49.690 188.410 50.010 188.470 ;
        RECT 46.470 188.270 50.010 188.410 ;
        RECT 46.470 188.210 46.790 188.270 ;
        RECT 49.690 188.210 50.010 188.270 ;
        RECT 50.150 188.410 50.470 188.470 ;
        RECT 51.085 188.410 51.375 188.455 ;
        RECT 50.150 188.270 51.375 188.410 ;
        RECT 50.150 188.210 50.470 188.270 ;
        RECT 51.085 188.225 51.375 188.270 ;
        RECT 54.245 188.250 54.535 188.565 ;
        RECT 73.150 188.550 73.470 188.610 ;
        RECT 55.325 188.410 55.615 188.455 ;
        RECT 58.905 188.410 59.195 188.455 ;
        RECT 60.740 188.410 61.030 188.455 ;
        RECT 55.325 188.270 61.030 188.410 ;
        RECT 55.325 188.225 55.615 188.270 ;
        RECT 58.905 188.225 59.195 188.270 ;
        RECT 60.740 188.225 61.030 188.270 ;
        RECT 61.190 188.210 61.510 188.470 ;
        RECT 62.585 188.225 62.875 188.455 ;
        RECT 63.965 188.410 64.255 188.455 ;
        RECT 67.630 188.410 67.950 188.470 ;
        RECT 63.965 188.270 67.950 188.410 ;
        RECT 63.965 188.225 64.255 188.270 ;
        RECT 36.365 188.070 36.655 188.115 ;
        RECT 36.810 188.070 37.130 188.130 ;
        RECT 36.365 187.930 37.130 188.070 ;
        RECT 36.365 187.885 36.655 187.930 ;
        RECT 36.810 187.870 37.130 187.930 ;
        RECT 37.270 188.070 37.590 188.130 ;
        RECT 37.745 188.070 38.035 188.115 ;
        RECT 45.090 188.070 45.410 188.130 ;
        RECT 37.270 187.930 45.410 188.070 ;
        RECT 37.270 187.870 37.590 187.930 ;
        RECT 37.745 187.885 38.035 187.930 ;
        RECT 45.090 187.870 45.410 187.930 ;
        RECT 47.390 187.870 47.710 188.130 ;
        RECT 59.350 188.070 59.670 188.130 ;
        RECT 54.380 187.930 59.670 188.070 ;
        RECT 54.380 187.790 54.520 187.930 ;
        RECT 59.350 187.870 59.670 187.930 ;
        RECT 59.810 187.870 60.130 188.130 ;
        RECT 62.660 188.070 62.800 188.225 ;
        RECT 67.630 188.210 67.950 188.270 ;
        RECT 68.090 188.210 68.410 188.470 ;
        RECT 71.310 188.410 71.630 188.470 ;
        RECT 69.100 188.270 71.630 188.410 ;
        RECT 69.100 188.070 69.240 188.270 ;
        RECT 71.310 188.210 71.630 188.270 ;
        RECT 71.770 188.210 72.090 188.470 ;
        RECT 75.005 188.410 75.295 188.455 ;
        RECT 75.450 188.410 75.770 188.470 ;
        RECT 75.005 188.270 75.770 188.410 ;
        RECT 75.005 188.225 75.295 188.270 ;
        RECT 75.450 188.210 75.770 188.270 ;
        RECT 77.750 188.210 78.070 188.470 ;
        RECT 79.590 188.210 79.910 188.470 ;
        RECT 80.050 188.210 80.370 188.470 ;
        RECT 80.600 188.455 80.740 188.610 ;
        RECT 81.060 188.610 81.660 188.750 ;
        RECT 82.810 188.750 83.130 188.810 ;
        RECT 83.285 188.750 83.575 188.795 ;
        RECT 82.810 188.610 83.575 188.750 ;
        RECT 81.060 188.455 81.200 188.610 ;
        RECT 82.810 188.550 83.130 188.610 ;
        RECT 83.285 188.565 83.575 188.610 ;
        RECT 86.490 188.550 86.810 188.810 ;
        RECT 98.450 188.550 98.770 188.810 ;
        RECT 98.910 188.750 99.230 188.810 ;
        RECT 100.865 188.750 101.155 188.795 ;
        RECT 104.105 188.750 104.755 188.795 ;
        RECT 98.910 188.610 104.755 188.750 ;
        RECT 98.910 188.550 99.230 188.610 ;
        RECT 100.865 188.565 101.455 188.610 ;
        RECT 104.105 188.565 104.755 188.610 ;
        RECT 109.030 188.750 109.350 188.810 ;
        RECT 109.950 188.750 110.270 188.810 ;
        RECT 113.185 188.750 113.475 188.795 ;
        RECT 116.505 188.750 116.795 188.795 ;
        RECT 119.745 188.750 120.395 188.795 ;
        RECT 109.030 188.610 112.940 188.750 ;
        RECT 80.525 188.225 80.815 188.455 ;
        RECT 80.985 188.225 81.275 188.455 ;
        RECT 81.430 188.410 81.750 188.470 ;
        RECT 81.905 188.410 82.195 188.455 ;
        RECT 81.430 188.270 82.195 188.410 ;
        RECT 81.430 188.210 81.750 188.270 ;
        RECT 81.905 188.225 82.195 188.270 ;
        RECT 85.110 188.410 85.430 188.470 ;
        RECT 90.185 188.410 90.475 188.455 ;
        RECT 85.110 188.270 90.475 188.410 ;
        RECT 85.110 188.210 85.430 188.270 ;
        RECT 90.185 188.225 90.475 188.270 ;
        RECT 101.165 188.250 101.455 188.565 ;
        RECT 109.030 188.550 109.350 188.610 ;
        RECT 109.950 188.550 110.270 188.610 ;
        RECT 102.245 188.410 102.535 188.455 ;
        RECT 105.825 188.410 106.115 188.455 ;
        RECT 107.660 188.410 107.950 188.455 ;
        RECT 102.245 188.270 107.950 188.410 ;
        RECT 102.245 188.225 102.535 188.270 ;
        RECT 105.825 188.225 106.115 188.270 ;
        RECT 107.660 188.225 107.950 188.270 ;
        RECT 108.125 188.410 108.415 188.455 ;
        RECT 110.870 188.410 111.190 188.470 ;
        RECT 112.800 188.455 112.940 188.610 ;
        RECT 113.185 188.610 120.395 188.750 ;
        RECT 113.185 188.565 113.475 188.610 ;
        RECT 116.505 188.565 117.095 188.610 ;
        RECT 119.745 188.565 120.395 188.610 ;
        RECT 108.125 188.270 111.190 188.410 ;
        RECT 108.125 188.225 108.415 188.270 ;
        RECT 110.870 188.210 111.190 188.270 ;
        RECT 112.725 188.225 113.015 188.455 ;
        RECT 116.805 188.250 117.095 188.565 ;
        RECT 117.885 188.410 118.175 188.455 ;
        RECT 121.465 188.410 121.755 188.455 ;
        RECT 123.300 188.410 123.590 188.455 ;
        RECT 117.885 188.270 123.590 188.410 ;
        RECT 117.885 188.225 118.175 188.270 ;
        RECT 121.465 188.225 121.755 188.270 ;
        RECT 123.300 188.225 123.590 188.270 ;
        RECT 62.660 187.930 69.240 188.070 ;
        RECT 78.685 188.070 78.975 188.115 ;
        RECT 85.585 188.070 85.875 188.115 ;
        RECT 87.410 188.070 87.730 188.130 ;
        RECT 78.685 187.930 79.820 188.070 ;
        RECT 78.685 187.885 78.975 187.930 ;
        RECT 79.680 187.790 79.820 187.930 ;
        RECT 80.140 187.930 87.730 188.070 ;
        RECT 40.605 187.730 40.895 187.775 ;
        RECT 43.725 187.730 44.015 187.775 ;
        RECT 45.615 187.730 45.905 187.775 ;
        RECT 40.605 187.590 45.905 187.730 ;
        RECT 40.605 187.545 40.895 187.590 ;
        RECT 43.725 187.545 44.015 187.590 ;
        RECT 45.615 187.545 45.905 187.590 ;
        RECT 51.990 187.530 52.310 187.790 ;
        RECT 52.450 187.530 52.770 187.790 ;
        RECT 54.290 187.530 54.610 187.790 ;
        RECT 55.325 187.730 55.615 187.775 ;
        RECT 58.445 187.730 58.735 187.775 ;
        RECT 60.335 187.730 60.625 187.775 ;
        RECT 55.325 187.590 60.625 187.730 ;
        RECT 55.325 187.545 55.615 187.590 ;
        RECT 58.445 187.545 58.735 187.590 ;
        RECT 60.335 187.545 60.625 187.590 ;
        RECT 79.590 187.530 79.910 187.790 ;
        RECT 39.570 187.390 39.890 187.450 ;
        RECT 45.170 187.390 45.460 187.435 ;
        RECT 39.570 187.250 45.460 187.390 ;
        RECT 39.570 187.190 39.890 187.250 ;
        RECT 45.170 187.205 45.460 187.250 ;
        RECT 49.690 187.390 50.010 187.450 ;
        RECT 61.190 187.390 61.510 187.450 ;
        RECT 49.690 187.250 61.510 187.390 ;
        RECT 49.690 187.190 50.010 187.250 ;
        RECT 61.190 187.190 61.510 187.250 ;
        RECT 65.330 187.190 65.650 187.450 ;
        RECT 77.305 187.390 77.595 187.435 ;
        RECT 80.140 187.390 80.280 187.930 ;
        RECT 85.585 187.885 85.875 187.930 ;
        RECT 87.410 187.870 87.730 187.930 ;
        RECT 106.270 188.070 106.590 188.130 ;
        RECT 111.345 188.070 111.635 188.115 ;
        RECT 111.790 188.070 112.110 188.130 ;
        RECT 106.270 187.930 112.110 188.070 ;
        RECT 106.270 187.870 106.590 187.930 ;
        RECT 111.345 187.885 111.635 187.930 ;
        RECT 111.790 187.870 112.110 187.930 ;
        RECT 123.765 188.070 124.055 188.115 ;
        RECT 124.670 188.070 124.990 188.130 ;
        RECT 123.765 187.930 124.990 188.070 ;
        RECT 123.765 187.885 124.055 187.930 ;
        RECT 124.670 187.870 124.990 187.930 ;
        RECT 102.245 187.730 102.535 187.775 ;
        RECT 105.365 187.730 105.655 187.775 ;
        RECT 107.255 187.730 107.545 187.775 ;
        RECT 102.245 187.590 107.545 187.730 ;
        RECT 102.245 187.545 102.535 187.590 ;
        RECT 105.365 187.545 105.655 187.590 ;
        RECT 107.255 187.545 107.545 187.590 ;
        RECT 117.885 187.730 118.175 187.775 ;
        RECT 121.005 187.730 121.295 187.775 ;
        RECT 122.895 187.730 123.185 187.775 ;
        RECT 117.885 187.590 123.185 187.730 ;
        RECT 117.885 187.545 118.175 187.590 ;
        RECT 121.005 187.545 121.295 187.590 ;
        RECT 122.895 187.545 123.185 187.590 ;
        RECT 77.305 187.250 80.280 187.390 ;
        RECT 99.385 187.390 99.675 187.435 ;
        RECT 99.830 187.390 100.150 187.450 ;
        RECT 99.385 187.250 100.150 187.390 ;
        RECT 77.305 187.205 77.595 187.250 ;
        RECT 99.385 187.205 99.675 187.250 ;
        RECT 99.830 187.190 100.150 187.250 ;
        RECT 101.210 187.390 101.530 187.450 ;
        RECT 106.810 187.390 107.100 187.435 ;
        RECT 101.210 187.250 107.100 187.390 ;
        RECT 101.210 187.190 101.530 187.250 ;
        RECT 106.810 187.205 107.100 187.250 ;
        RECT 121.450 187.390 121.770 187.450 ;
        RECT 122.450 187.390 122.740 187.435 ;
        RECT 121.450 187.250 122.740 187.390 ;
        RECT 121.450 187.190 121.770 187.250 ;
        RECT 122.450 187.205 122.740 187.250 ;
        RECT 29.840 186.570 127.820 187.050 ;
        RECT 34.985 186.370 35.275 186.415 ;
        RECT 40.030 186.370 40.350 186.430 ;
        RECT 34.985 186.230 40.350 186.370 ;
        RECT 34.985 186.185 35.275 186.230 ;
        RECT 31.765 185.690 32.055 185.735 ;
        RECT 35.060 185.690 35.200 186.185 ;
        RECT 40.030 186.170 40.350 186.230 ;
        RECT 49.230 186.170 49.550 186.430 ;
        RECT 54.765 186.370 55.055 186.415 ;
        RECT 57.050 186.370 57.370 186.430 ;
        RECT 54.765 186.230 57.370 186.370 ;
        RECT 54.765 186.185 55.055 186.230 ;
        RECT 57.050 186.170 57.370 186.230 ;
        RECT 61.190 186.170 61.510 186.430 ;
        RECT 67.630 186.370 67.950 186.430 ;
        RECT 80.050 186.370 80.370 186.430 ;
        RECT 86.030 186.370 86.350 186.430 ;
        RECT 89.265 186.370 89.555 186.415 ;
        RECT 67.630 186.230 71.310 186.370 ;
        RECT 67.630 186.170 67.950 186.230 ;
        RECT 37.845 186.030 38.135 186.075 ;
        RECT 40.965 186.030 41.255 186.075 ;
        RECT 42.855 186.030 43.145 186.075 ;
        RECT 46.470 186.030 46.790 186.090 ;
        RECT 69.470 186.030 69.790 186.090 ;
        RECT 37.845 185.890 43.145 186.030 ;
        RECT 37.845 185.845 38.135 185.890 ;
        RECT 40.965 185.845 41.255 185.890 ;
        RECT 42.855 185.845 43.145 185.890 ;
        RECT 43.800 185.890 46.790 186.030 ;
        RECT 31.765 185.550 35.200 185.690 ;
        RECT 41.870 185.690 42.190 185.750 ;
        RECT 43.800 185.735 43.940 185.890 ;
        RECT 46.470 185.830 46.790 185.890 ;
        RECT 56.220 185.890 69.790 186.030 ;
        RECT 71.170 186.030 71.310 186.230 ;
        RECT 80.050 186.230 85.800 186.370 ;
        RECT 80.050 186.170 80.370 186.230 ;
        RECT 72.245 186.030 72.535 186.075 ;
        RECT 71.170 185.890 72.535 186.030 ;
        RECT 42.345 185.690 42.635 185.735 ;
        RECT 41.870 185.550 42.635 185.690 ;
        RECT 31.765 185.505 32.055 185.550 ;
        RECT 41.870 185.490 42.190 185.550 ;
        RECT 42.345 185.505 42.635 185.550 ;
        RECT 43.725 185.505 44.015 185.735 ;
        RECT 45.090 185.690 45.410 185.750 ;
        RECT 47.390 185.690 47.710 185.750 ;
        RECT 52.005 185.690 52.295 185.735 ;
        RECT 56.220 185.690 56.360 185.890 ;
        RECT 69.470 185.830 69.790 185.890 ;
        RECT 72.245 185.845 72.535 185.890 ;
        RECT 74.990 186.030 75.310 186.090 ;
        RECT 85.660 186.030 85.800 186.230 ;
        RECT 86.030 186.230 89.555 186.370 ;
        RECT 86.030 186.170 86.350 186.230 ;
        RECT 89.265 186.185 89.555 186.230 ;
        RECT 91.640 186.230 100.980 186.370 ;
        RECT 91.640 186.030 91.780 186.230 ;
        RECT 74.990 185.890 84.880 186.030 ;
        RECT 85.660 185.890 91.780 186.030 ;
        RECT 92.125 186.030 92.415 186.075 ;
        RECT 95.245 186.030 95.535 186.075 ;
        RECT 97.135 186.030 97.425 186.075 ;
        RECT 100.840 186.030 100.980 186.230 ;
        RECT 101.210 186.170 101.530 186.430 ;
        RECT 121.450 186.370 121.770 186.430 ;
        RECT 122.845 186.370 123.135 186.415 ;
        RECT 121.450 186.230 123.135 186.370 ;
        RECT 121.450 186.170 121.770 186.230 ;
        RECT 122.845 186.185 123.135 186.230 ;
        RECT 124.210 186.170 124.530 186.430 ;
        RECT 105.810 186.030 106.130 186.090 ;
        RECT 92.125 185.890 97.425 186.030 ;
        RECT 74.990 185.830 75.310 185.890 ;
        RECT 45.090 185.550 51.760 185.690 ;
        RECT 45.090 185.490 45.410 185.550 ;
        RECT 47.390 185.490 47.710 185.550 ;
        RECT 36.810 185.370 37.130 185.410 ;
        RECT 36.765 185.150 37.130 185.370 ;
        RECT 37.845 185.350 38.135 185.395 ;
        RECT 41.425 185.350 41.715 185.395 ;
        RECT 43.260 185.350 43.550 185.395 ;
        RECT 37.845 185.210 43.550 185.350 ;
        RECT 37.845 185.165 38.135 185.210 ;
        RECT 41.425 185.165 41.715 185.210 ;
        RECT 43.260 185.165 43.550 185.210 ;
        RECT 45.180 185.210 48.540 185.350 ;
        RECT 36.765 185.055 37.055 185.150 ;
        RECT 36.465 185.010 37.055 185.055 ;
        RECT 39.705 185.010 40.355 185.055 ;
        RECT 36.465 184.870 40.355 185.010 ;
        RECT 36.465 184.825 36.755 184.870 ;
        RECT 39.705 184.825 40.355 184.870 ;
        RECT 42.790 185.010 43.110 185.070 ;
        RECT 45.180 185.010 45.320 185.210 ;
        RECT 42.790 184.870 45.320 185.010 ;
        RECT 42.790 184.810 43.110 184.870 ;
        RECT 45.550 184.810 45.870 185.070 ;
        RECT 48.400 185.010 48.540 185.210 ;
        RECT 48.770 185.150 49.090 185.410 ;
        RECT 51.620 185.350 51.760 185.550 ;
        RECT 52.005 185.550 56.360 185.690 ;
        RECT 52.005 185.505 52.295 185.550 ;
        RECT 54.290 185.350 54.610 185.410 ;
        RECT 51.620 185.210 54.610 185.350 ;
        RECT 54.290 185.150 54.610 185.210 ;
        RECT 55.210 185.150 55.530 185.410 ;
        RECT 56.220 185.395 56.360 185.550 ;
        RECT 63.950 185.690 64.270 185.750 ;
        RECT 68.565 185.690 68.855 185.735 ;
        RECT 76.845 185.690 77.135 185.735 ;
        RECT 63.950 185.550 77.135 185.690 ;
        RECT 63.950 185.490 64.270 185.550 ;
        RECT 68.565 185.505 68.855 185.550 ;
        RECT 76.845 185.505 77.135 185.550 ;
        RECT 81.890 185.490 82.210 185.750 ;
        RECT 56.145 185.165 56.435 185.395 ;
        RECT 56.590 185.150 56.910 185.410 ;
        RECT 57.065 185.350 57.355 185.395 ;
        RECT 61.190 185.350 61.510 185.410 ;
        RECT 57.065 185.210 61.510 185.350 ;
        RECT 57.065 185.165 57.355 185.210 ;
        RECT 61.190 185.150 61.510 185.210 ;
        RECT 65.330 185.350 65.650 185.410 ;
        RECT 69.945 185.350 70.235 185.395 ;
        RECT 75.005 185.350 75.295 185.395 ;
        RECT 65.330 185.210 70.235 185.350 ;
        RECT 65.330 185.150 65.650 185.210 ;
        RECT 69.945 185.165 70.235 185.210 ;
        RECT 71.860 185.210 75.295 185.350 ;
        RECT 52.450 185.010 52.770 185.070 ;
        RECT 54.750 185.010 55.070 185.070 ;
        RECT 48.400 184.870 55.070 185.010 ;
        RECT 52.450 184.810 52.770 184.870 ;
        RECT 54.750 184.810 55.070 184.870 ;
        RECT 64.410 185.010 64.730 185.070 ;
        RECT 67.630 185.010 67.950 185.070 ;
        RECT 64.410 184.870 67.950 185.010 ;
        RECT 64.410 184.810 64.730 184.870 ;
        RECT 67.630 184.810 67.950 184.870 ;
        RECT 69.470 184.810 69.790 185.070 ;
        RECT 34.525 184.670 34.815 184.715 ;
        RECT 42.330 184.670 42.650 184.730 ;
        RECT 46.025 184.670 46.315 184.715 ;
        RECT 34.525 184.530 46.315 184.670 ;
        RECT 34.525 184.485 34.815 184.530 ;
        RECT 42.330 184.470 42.650 184.530 ;
        RECT 46.025 184.485 46.315 184.530 ;
        RECT 46.470 184.670 46.790 184.730 ;
        RECT 47.865 184.670 48.155 184.715 ;
        RECT 46.470 184.530 48.155 184.670 ;
        RECT 46.470 184.470 46.790 184.530 ;
        RECT 47.865 184.485 48.155 184.530 ;
        RECT 58.430 184.470 58.750 184.730 ;
        RECT 71.860 184.715 72.000 185.210 ;
        RECT 75.005 185.165 75.295 185.210 ;
        RECT 79.145 185.350 79.435 185.395 ;
        RECT 80.050 185.350 80.370 185.410 ;
        RECT 81.980 185.350 82.120 185.490 ;
        RECT 84.740 185.410 84.880 185.890 ;
        RECT 92.125 185.845 92.415 185.890 ;
        RECT 95.245 185.845 95.535 185.890 ;
        RECT 97.135 185.845 97.425 185.890 ;
        RECT 97.620 185.890 100.060 186.030 ;
        RECT 100.840 185.890 106.130 186.030 ;
        RECT 86.045 185.505 86.335 185.735 ;
        RECT 97.620 185.690 97.760 185.890 ;
        RECT 99.920 185.750 100.060 185.890 ;
        RECT 105.810 185.830 106.130 185.890 ;
        RECT 106.270 186.030 106.590 186.090 ;
        RECT 111.330 186.030 111.650 186.090 ;
        RECT 106.270 185.890 111.650 186.030 ;
        RECT 106.270 185.830 106.590 185.890 ;
        RECT 90.720 185.550 97.760 185.690 ;
        RECT 98.005 185.690 98.295 185.735 ;
        RECT 98.450 185.690 98.770 185.750 ;
        RECT 98.005 185.550 98.770 185.690 ;
        RECT 79.145 185.210 82.120 185.350 ;
        RECT 79.145 185.165 79.435 185.210 ;
        RECT 80.050 185.150 80.370 185.210 ;
        RECT 82.810 185.150 83.130 185.410 ;
        RECT 83.285 185.165 83.575 185.395 ;
        RECT 83.745 185.165 84.035 185.395 ;
        RECT 76.370 185.010 76.690 185.070 ;
        RECT 77.750 185.010 78.070 185.070 ;
        RECT 78.225 185.010 78.515 185.055 ;
        RECT 76.370 184.870 78.515 185.010 ;
        RECT 76.370 184.810 76.690 184.870 ;
        RECT 77.750 184.810 78.070 184.870 ;
        RECT 78.225 184.825 78.515 184.870 ;
        RECT 71.785 184.485 72.075 184.715 ;
        RECT 81.430 184.470 81.750 184.730 ;
        RECT 83.360 184.670 83.500 185.165 ;
        RECT 83.820 185.010 83.960 185.165 ;
        RECT 84.650 185.150 84.970 185.410 ;
        RECT 86.120 185.350 86.260 185.505 ;
        RECT 87.410 185.350 87.730 185.410 ;
        RECT 90.720 185.350 90.860 185.550 ;
        RECT 98.005 185.505 98.295 185.550 ;
        RECT 98.450 185.490 98.770 185.550 ;
        RECT 99.830 185.690 100.150 185.750 ;
        RECT 104.445 185.690 104.735 185.735 ;
        RECT 99.830 185.550 104.735 185.690 ;
        RECT 99.830 185.490 100.150 185.550 ;
        RECT 104.445 185.505 104.735 185.550 ;
        RECT 105.350 185.490 105.670 185.750 ;
        RECT 109.580 185.735 109.720 185.890 ;
        RECT 111.330 185.830 111.650 185.890 ;
        RECT 111.790 186.030 112.110 186.090 ;
        RECT 116.390 186.030 116.710 186.090 ;
        RECT 111.790 185.890 114.780 186.030 ;
        RECT 111.790 185.830 112.110 185.890 ;
        RECT 114.640 185.735 114.780 185.890 ;
        RECT 116.390 185.890 123.520 186.030 ;
        RECT 116.390 185.830 116.710 185.890 ;
        RECT 109.505 185.505 109.795 185.735 ;
        RECT 114.565 185.505 114.855 185.735 ;
        RECT 117.310 185.690 117.630 185.750 ;
        RECT 121.005 185.690 121.295 185.735 ;
        RECT 117.310 185.550 121.295 185.690 ;
        RECT 117.310 185.490 117.630 185.550 ;
        RECT 121.005 185.505 121.295 185.550 ;
        RECT 86.120 185.210 87.730 185.350 ;
        RECT 87.410 185.150 87.730 185.210 ;
        RECT 88.420 185.210 90.860 185.350 ;
        RECT 83.820 184.870 87.180 185.010 ;
        RECT 84.190 184.670 84.510 184.730 ;
        RECT 83.360 184.530 84.510 184.670 ;
        RECT 84.190 184.470 84.510 184.530 ;
        RECT 86.490 184.470 86.810 184.730 ;
        RECT 87.040 184.715 87.180 184.870 ;
        RECT 86.965 184.670 87.255 184.715 ;
        RECT 88.420 184.670 88.560 185.210 ;
        RECT 89.250 185.010 89.570 185.070 ;
        RECT 91.045 185.055 91.335 185.370 ;
        RECT 92.125 185.350 92.415 185.395 ;
        RECT 95.705 185.350 95.995 185.395 ;
        RECT 97.540 185.350 97.830 185.395 ;
        RECT 92.125 185.210 97.830 185.350 ;
        RECT 92.125 185.165 92.415 185.210 ;
        RECT 95.705 185.165 95.995 185.210 ;
        RECT 97.540 185.165 97.830 185.210 ;
        RECT 99.385 185.165 99.675 185.395 ;
        RECT 90.745 185.010 91.335 185.055 ;
        RECT 93.985 185.010 94.635 185.055 ;
        RECT 89.250 184.870 94.635 185.010 ;
        RECT 89.250 184.810 89.570 184.870 ;
        RECT 90.745 184.825 91.035 184.870 ;
        RECT 93.985 184.825 94.635 184.870 ;
        RECT 96.625 184.825 96.915 185.055 ;
        RECT 97.070 185.010 97.390 185.070 ;
        RECT 99.460 185.010 99.600 185.165 ;
        RECT 100.290 185.150 100.610 185.410 ;
        RECT 103.985 185.350 104.275 185.395 ;
        RECT 106.285 185.350 106.575 185.395 ;
        RECT 103.985 185.210 106.575 185.350 ;
        RECT 103.985 185.165 104.275 185.210 ;
        RECT 106.285 185.165 106.575 185.210 ;
        RECT 109.030 185.350 109.350 185.410 ;
        RECT 111.345 185.350 111.635 185.395 ;
        RECT 109.030 185.210 111.635 185.350 ;
        RECT 109.030 185.150 109.350 185.210 ;
        RECT 111.345 185.165 111.635 185.210 ;
        RECT 111.805 185.165 112.095 185.395 ;
        RECT 112.265 185.350 112.555 185.395 ;
        RECT 112.710 185.350 113.030 185.410 ;
        RECT 112.265 185.210 113.030 185.350 ;
        RECT 112.265 185.165 112.555 185.210 ;
        RECT 97.070 184.870 99.600 185.010 ;
        RECT 109.490 185.010 109.810 185.070 ;
        RECT 111.880 185.010 112.020 185.165 ;
        RECT 112.710 185.150 113.030 185.210 ;
        RECT 113.170 185.150 113.490 185.410 ;
        RECT 115.930 185.350 116.250 185.410 ;
        RECT 118.245 185.350 118.535 185.395 ;
        RECT 115.930 185.210 118.535 185.350 ;
        RECT 115.930 185.150 116.250 185.210 ;
        RECT 118.245 185.165 118.535 185.210 ;
        RECT 121.910 185.150 122.230 185.410 ;
        RECT 123.380 185.395 123.520 185.890 ;
        RECT 123.305 185.165 123.595 185.395 ;
        RECT 109.490 184.870 112.020 185.010 ;
        RECT 112.800 185.010 112.940 185.150 ;
        RECT 115.485 185.010 115.775 185.055 ;
        RECT 112.800 184.870 115.775 185.010 ;
        RECT 86.965 184.530 88.560 184.670 ;
        RECT 88.805 184.670 89.095 184.715 ;
        RECT 90.170 184.670 90.490 184.730 ;
        RECT 88.805 184.530 90.490 184.670 ;
        RECT 96.700 184.670 96.840 184.825 ;
        RECT 97.070 184.810 97.390 184.870 ;
        RECT 109.490 184.810 109.810 184.870 ;
        RECT 115.485 184.825 115.775 184.870 ;
        RECT 98.465 184.670 98.755 184.715 ;
        RECT 96.700 184.530 98.755 184.670 ;
        RECT 86.965 184.485 87.255 184.530 ;
        RECT 88.805 184.485 89.095 184.530 ;
        RECT 90.170 184.470 90.490 184.530 ;
        RECT 98.465 184.485 98.755 184.530 ;
        RECT 102.130 184.470 102.450 184.730 ;
        RECT 109.965 184.670 110.255 184.715 ;
        RECT 111.790 184.670 112.110 184.730 ;
        RECT 109.965 184.530 112.110 184.670 ;
        RECT 109.965 184.485 110.255 184.530 ;
        RECT 111.790 184.470 112.110 184.530 ;
        RECT 117.785 184.670 118.075 184.715 ;
        RECT 118.690 184.670 119.010 184.730 ;
        RECT 117.785 184.530 119.010 184.670 ;
        RECT 117.785 184.485 118.075 184.530 ;
        RECT 118.690 184.470 119.010 184.530 ;
        RECT 29.840 183.850 127.820 184.330 ;
        RECT 39.570 183.450 39.890 183.710 ;
        RECT 42.330 183.450 42.650 183.710 ;
        RECT 44.630 183.650 44.950 183.710 ;
        RECT 53.385 183.650 53.675 183.695 ;
        RECT 44.630 183.510 53.675 183.650 ;
        RECT 44.630 183.450 44.950 183.510 ;
        RECT 53.385 183.465 53.675 183.510 ;
        RECT 54.750 183.650 55.070 183.710 ;
        RECT 55.225 183.650 55.515 183.695 ;
        RECT 54.750 183.510 55.515 183.650 ;
        RECT 54.750 183.450 55.070 183.510 ;
        RECT 55.225 183.465 55.515 183.510 ;
        RECT 58.445 183.650 58.735 183.695 ;
        RECT 59.810 183.650 60.130 183.710 ;
        RECT 58.445 183.510 60.130 183.650 ;
        RECT 58.445 183.465 58.735 183.510 ;
        RECT 59.810 183.450 60.130 183.510 ;
        RECT 65.330 183.450 65.650 183.710 ;
        RECT 65.790 183.450 66.110 183.710 ;
        RECT 68.090 183.450 68.410 183.710 ;
        RECT 72.230 183.650 72.550 183.710 ;
        RECT 74.530 183.650 74.850 183.710 ;
        RECT 84.650 183.650 84.970 183.710 ;
        RECT 87.885 183.650 88.175 183.695 ;
        RECT 89.250 183.650 89.570 183.710 ;
        RECT 72.230 183.510 82.120 183.650 ;
        RECT 72.230 183.450 72.550 183.510 ;
        RECT 74.530 183.450 74.850 183.510 ;
        RECT 32.685 183.310 32.975 183.355 ;
        RECT 45.665 183.310 45.955 183.355 ;
        RECT 48.905 183.310 49.555 183.355 ;
        RECT 32.685 183.170 49.555 183.310 ;
        RECT 32.685 183.125 32.975 183.170 ;
        RECT 45.665 183.125 46.255 183.170 ;
        RECT 48.905 183.125 49.555 183.170 ;
        RECT 51.545 183.310 51.835 183.355 ;
        RECT 51.990 183.310 52.310 183.370 ;
        RECT 63.950 183.310 64.270 183.370 ;
        RECT 69.585 183.310 69.875 183.355 ;
        RECT 70.390 183.310 70.710 183.370 ;
        RECT 72.825 183.310 73.475 183.355 ;
        RECT 51.545 183.170 52.310 183.310 ;
        RECT 51.545 183.125 51.835 183.170 ;
        RECT 33.145 182.970 33.435 183.015 ;
        RECT 35.430 182.970 35.750 183.030 ;
        RECT 33.145 182.830 35.750 182.970 ;
        RECT 33.145 182.785 33.435 182.830 ;
        RECT 35.430 182.770 35.750 182.830 ;
        RECT 38.650 182.770 38.970 183.030 ;
        RECT 41.885 182.970 42.175 183.015 ;
        RECT 41.885 182.830 44.860 182.970 ;
        RECT 41.885 182.785 42.175 182.830 ;
        RECT 34.065 182.445 34.355 182.675 ;
        RECT 36.825 182.630 37.115 182.675 ;
        RECT 41.960 182.630 42.100 182.785 ;
        RECT 36.825 182.490 42.100 182.630 ;
        RECT 43.265 182.630 43.555 182.675 ;
        RECT 43.710 182.630 44.030 182.690 ;
        RECT 43.265 182.490 44.030 182.630 ;
        RECT 36.825 182.445 37.115 182.490 ;
        RECT 43.265 182.445 43.555 182.490 ;
        RECT 34.140 182.290 34.280 182.445 ;
        RECT 43.710 182.430 44.030 182.490 ;
        RECT 36.350 182.290 36.670 182.350 ;
        RECT 44.185 182.290 44.475 182.335 ;
        RECT 34.140 182.150 44.475 182.290 ;
        RECT 36.350 182.090 36.670 182.150 ;
        RECT 44.185 182.105 44.475 182.150 ;
        RECT 37.270 181.950 37.590 182.010 ;
        RECT 40.045 181.950 40.335 181.995 ;
        RECT 37.270 181.810 40.335 181.950 ;
        RECT 37.270 181.750 37.590 181.810 ;
        RECT 40.045 181.765 40.335 181.810 ;
        RECT 41.410 181.950 41.730 182.010 ;
        RECT 42.790 181.950 43.110 182.010 ;
        RECT 41.410 181.810 43.110 181.950 ;
        RECT 44.720 181.950 44.860 182.830 ;
        RECT 45.965 182.810 46.255 183.125 ;
        RECT 51.990 183.110 52.310 183.170 ;
        RECT 56.680 183.170 64.640 183.310 ;
        RECT 47.045 182.970 47.335 183.015 ;
        RECT 50.625 182.970 50.915 183.015 ;
        RECT 52.460 182.970 52.750 183.015 ;
        RECT 47.045 182.830 52.750 182.970 ;
        RECT 47.045 182.785 47.335 182.830 ;
        RECT 50.625 182.785 50.915 182.830 ;
        RECT 52.460 182.785 52.750 182.830 ;
        RECT 54.290 182.970 54.610 183.030 ;
        RECT 56.680 182.970 56.820 183.170 ;
        RECT 63.950 183.110 64.270 183.170 ;
        RECT 54.290 182.830 56.820 182.970 ;
        RECT 54.290 182.770 54.610 182.830 ;
        RECT 49.690 182.630 50.010 182.690 ;
        RECT 56.680 182.675 56.820 182.830 ;
        RECT 57.525 182.970 57.815 183.015 ;
        RECT 57.970 182.970 58.290 183.030 ;
        RECT 57.525 182.830 58.290 182.970 ;
        RECT 57.525 182.785 57.815 182.830 ;
        RECT 57.970 182.770 58.290 182.830 ;
        RECT 59.365 182.785 59.655 183.015 ;
        RECT 52.925 182.630 53.215 182.675 ;
        RECT 49.690 182.490 53.215 182.630 ;
        RECT 49.690 182.430 50.010 182.490 ;
        RECT 52.925 182.445 53.215 182.490 ;
        RECT 55.685 182.445 55.975 182.675 ;
        RECT 56.605 182.445 56.895 182.675 ;
        RECT 57.050 182.630 57.370 182.690 ;
        RECT 59.440 182.630 59.580 182.785 ;
        RECT 60.270 182.770 60.590 183.030 ;
        RECT 60.745 182.785 61.035 183.015 ;
        RECT 57.050 182.490 59.580 182.630 ;
        RECT 47.045 182.290 47.335 182.335 ;
        RECT 50.165 182.290 50.455 182.335 ;
        RECT 52.055 182.290 52.345 182.335 ;
        RECT 47.045 182.150 52.345 182.290 ;
        RECT 47.045 182.105 47.335 182.150 ;
        RECT 50.165 182.105 50.455 182.150 ;
        RECT 52.055 182.105 52.345 182.150 ;
        RECT 55.760 181.950 55.900 182.445 ;
        RECT 57.050 182.430 57.370 182.490 ;
        RECT 56.130 182.290 56.450 182.350 ;
        RECT 60.820 182.290 60.960 182.785 ;
        RECT 61.190 182.770 61.510 183.030 ;
        RECT 64.500 182.675 64.640 183.170 ;
        RECT 69.585 183.170 73.475 183.310 ;
        RECT 69.585 183.125 70.175 183.170 ;
        RECT 69.885 182.810 70.175 183.125 ;
        RECT 70.390 183.110 70.710 183.170 ;
        RECT 72.825 183.125 73.475 183.170 ;
        RECT 74.990 183.310 75.310 183.370 ;
        RECT 75.465 183.310 75.755 183.355 ;
        RECT 77.750 183.310 78.070 183.370 ;
        RECT 80.050 183.310 80.370 183.370 ;
        RECT 74.990 183.170 75.755 183.310 ;
        RECT 74.990 183.110 75.310 183.170 ;
        RECT 75.465 183.125 75.755 183.170 ;
        RECT 77.380 183.170 80.370 183.310 ;
        RECT 77.380 183.015 77.520 183.170 ;
        RECT 77.750 183.110 78.070 183.170 ;
        RECT 80.050 183.110 80.370 183.170 ;
        RECT 81.980 183.310 82.120 183.510 ;
        RECT 84.650 183.510 86.720 183.650 ;
        RECT 84.650 183.450 84.970 183.510 ;
        RECT 84.190 183.310 84.510 183.370 ;
        RECT 81.980 183.170 85.800 183.310 ;
        RECT 70.965 182.970 71.255 183.015 ;
        RECT 74.545 182.970 74.835 183.015 ;
        RECT 76.380 182.970 76.670 183.015 ;
        RECT 70.965 182.830 76.670 182.970 ;
        RECT 70.965 182.785 71.255 182.830 ;
        RECT 74.545 182.785 74.835 182.830 ;
        RECT 76.380 182.785 76.670 182.830 ;
        RECT 77.305 182.785 77.595 183.015 ;
        RECT 78.210 182.970 78.530 183.030 ;
        RECT 81.980 183.015 82.120 183.170 ;
        RECT 84.190 183.110 84.510 183.170 ;
        RECT 79.145 182.970 79.435 183.015 ;
        RECT 81.445 182.970 81.735 183.015 ;
        RECT 78.210 182.830 79.435 182.970 ;
        RECT 78.210 182.770 78.530 182.830 ;
        RECT 79.145 182.785 79.435 182.830 ;
        RECT 79.680 182.830 81.735 182.970 ;
        RECT 64.425 182.445 64.715 182.675 ;
        RECT 75.450 182.630 75.770 182.690 ;
        RECT 76.845 182.630 77.135 182.675 ;
        RECT 75.450 182.490 77.135 182.630 ;
        RECT 75.450 182.430 75.770 182.490 ;
        RECT 76.845 182.445 77.135 182.490 ;
        RECT 78.685 182.445 78.975 182.675 ;
        RECT 69.010 182.290 69.330 182.350 ;
        RECT 56.130 182.150 69.330 182.290 ;
        RECT 56.130 182.090 56.450 182.150 ;
        RECT 69.010 182.090 69.330 182.150 ;
        RECT 70.965 182.290 71.255 182.335 ;
        RECT 74.085 182.290 74.375 182.335 ;
        RECT 75.975 182.290 76.265 182.335 ;
        RECT 70.965 182.150 76.265 182.290 ;
        RECT 70.965 182.105 71.255 182.150 ;
        RECT 74.085 182.105 74.375 182.150 ;
        RECT 75.975 182.105 76.265 182.150 ;
        RECT 77.290 182.290 77.610 182.350 ;
        RECT 78.225 182.290 78.515 182.335 ;
        RECT 77.290 182.150 78.515 182.290 ;
        RECT 78.760 182.290 78.900 182.445 ;
        RECT 79.130 182.290 79.450 182.350 ;
        RECT 78.760 182.150 79.450 182.290 ;
        RECT 77.290 182.090 77.610 182.150 ;
        RECT 78.225 182.105 78.515 182.150 ;
        RECT 79.130 182.090 79.450 182.150 ;
        RECT 44.720 181.810 55.900 181.950 ;
        RECT 59.350 181.950 59.670 182.010 ;
        RECT 62.585 181.950 62.875 181.995 ;
        RECT 59.350 181.810 62.875 181.950 ;
        RECT 41.410 181.750 41.730 181.810 ;
        RECT 42.790 181.750 43.110 181.810 ;
        RECT 59.350 181.750 59.670 181.810 ;
        RECT 62.585 181.765 62.875 181.810 ;
        RECT 67.645 181.950 67.935 181.995 ;
        RECT 69.930 181.950 70.250 182.010 ;
        RECT 67.645 181.810 70.250 181.950 ;
        RECT 67.645 181.765 67.935 181.810 ;
        RECT 69.930 181.750 70.250 181.810 ;
        RECT 73.610 181.950 73.930 182.010 ;
        RECT 77.765 181.950 78.055 181.995 ;
        RECT 73.610 181.810 78.055 181.950 ;
        RECT 73.610 181.750 73.930 181.810 ;
        RECT 77.765 181.765 78.055 181.810 ;
        RECT 78.670 181.950 78.990 182.010 ;
        RECT 79.680 181.950 79.820 182.830 ;
        RECT 81.445 182.785 81.735 182.830 ;
        RECT 81.905 182.785 82.195 183.015 ;
        RECT 81.520 182.630 81.660 182.785 ;
        RECT 82.350 182.770 82.670 183.030 ;
        RECT 83.285 182.970 83.575 183.015 ;
        RECT 84.650 182.970 84.970 183.030 ;
        RECT 85.660 183.015 85.800 183.170 ;
        RECT 83.285 182.830 84.970 182.970 ;
        RECT 83.285 182.785 83.575 182.830 ;
        RECT 84.650 182.770 84.970 182.830 ;
        RECT 85.125 182.785 85.415 183.015 ;
        RECT 85.585 182.785 85.875 183.015 ;
        RECT 82.810 182.630 83.130 182.690 ;
        RECT 85.200 182.630 85.340 182.785 ;
        RECT 86.030 182.770 86.350 183.030 ;
        RECT 86.580 182.970 86.720 183.510 ;
        RECT 87.885 183.510 89.570 183.650 ;
        RECT 87.885 183.465 88.175 183.510 ;
        RECT 89.250 183.450 89.570 183.510 ;
        RECT 100.290 183.450 100.610 183.710 ;
        RECT 105.810 183.650 106.130 183.710 ;
        RECT 109.030 183.650 109.350 183.710 ;
        RECT 105.810 183.510 109.350 183.650 ;
        RECT 105.810 183.450 106.130 183.510 ;
        RECT 109.030 183.450 109.350 183.510 ;
        RECT 109.950 183.650 110.270 183.710 ;
        RECT 109.950 183.510 112.020 183.650 ;
        RECT 109.950 183.450 110.270 183.510 ;
        RECT 100.750 183.310 101.070 183.370 ;
        RECT 100.750 183.170 110.180 183.310 ;
        RECT 100.750 183.110 101.070 183.170 ;
        RECT 86.965 182.970 87.255 183.015 ;
        RECT 86.580 182.830 87.255 182.970 ;
        RECT 86.965 182.785 87.255 182.830 ;
        RECT 87.410 182.770 87.730 183.030 ;
        RECT 98.450 182.970 98.770 183.030 ;
        RECT 98.925 182.970 99.215 183.015 ;
        RECT 98.450 182.830 99.215 182.970 ;
        RECT 98.450 182.770 98.770 182.830 ;
        RECT 98.925 182.785 99.215 182.830 ;
        RECT 102.130 182.970 102.450 183.030 ;
        RECT 103.065 182.970 103.355 183.015 ;
        RECT 102.130 182.830 103.355 182.970 ;
        RECT 102.130 182.770 102.450 182.830 ;
        RECT 103.065 182.785 103.355 182.830 ;
        RECT 105.350 182.770 105.670 183.030 ;
        RECT 105.810 182.770 106.130 183.030 ;
        RECT 106.270 182.770 106.590 183.030 ;
        RECT 106.730 182.970 107.050 183.030 ;
        RECT 107.205 182.970 107.495 183.015 ;
        RECT 106.730 182.830 107.495 182.970 ;
        RECT 106.730 182.770 107.050 182.830 ;
        RECT 107.205 182.785 107.495 182.830 ;
        RECT 109.030 182.770 109.350 183.030 ;
        RECT 109.490 182.770 109.810 183.030 ;
        RECT 110.040 183.015 110.180 183.170 ;
        RECT 109.965 182.785 110.255 183.015 ;
        RECT 110.885 182.970 111.175 183.015 ;
        RECT 111.330 182.970 111.650 183.030 ;
        RECT 111.880 183.015 112.020 183.510 ;
        RECT 112.250 183.450 112.570 183.710 ;
        RECT 113.170 183.650 113.490 183.710 ;
        RECT 113.170 183.510 118.460 183.650 ;
        RECT 113.170 183.450 113.490 183.510 ;
        RECT 112.340 183.170 117.080 183.310 ;
        RECT 110.885 182.830 111.650 182.970 ;
        RECT 110.885 182.785 111.175 182.830 ;
        RECT 111.330 182.770 111.650 182.830 ;
        RECT 111.805 182.785 112.095 183.015 ;
        RECT 81.520 182.490 85.340 182.630 ;
        RECT 105.900 182.630 106.040 182.770 ;
        RECT 109.580 182.630 109.720 182.770 ;
        RECT 112.340 182.630 112.480 183.170 ;
        RECT 113.185 182.970 113.475 183.015 ;
        RECT 115.930 182.970 116.250 183.030 ;
        RECT 116.940 183.015 117.080 183.170 ;
        RECT 113.185 182.830 116.250 182.970 ;
        RECT 113.185 182.785 113.475 182.830 ;
        RECT 115.930 182.770 116.250 182.830 ;
        RECT 116.405 182.785 116.695 183.015 ;
        RECT 116.865 182.785 117.155 183.015 ;
        RECT 105.900 182.490 112.480 182.630 ;
        RECT 82.810 182.430 83.130 182.490 ;
        RECT 109.030 182.290 109.350 182.350 ;
        RECT 116.480 182.290 116.620 182.785 ;
        RECT 117.310 182.770 117.630 183.030 ;
        RECT 118.320 183.015 118.460 183.510 ;
        RECT 121.910 183.450 122.230 183.710 ;
        RECT 118.245 182.785 118.535 183.015 ;
        RECT 118.690 182.770 119.010 183.030 ;
        RECT 119.150 182.970 119.470 183.030 ;
        RECT 122.385 182.970 122.675 183.015 ;
        RECT 119.150 182.830 122.675 182.970 ;
        RECT 119.150 182.770 119.470 182.830 ;
        RECT 122.385 182.785 122.675 182.830 ;
        RECT 109.030 182.150 116.620 182.290 ;
        RECT 109.030 182.090 109.350 182.150 ;
        RECT 78.670 181.810 79.820 181.950 ;
        RECT 78.670 181.750 78.990 181.810 ;
        RECT 80.050 181.750 80.370 182.010 ;
        RECT 83.730 181.750 84.050 182.010 ;
        RECT 103.050 181.950 103.370 182.010 ;
        RECT 103.985 181.950 104.275 181.995 ;
        RECT 103.050 181.810 104.275 181.950 ;
        RECT 103.050 181.750 103.370 181.810 ;
        RECT 103.985 181.765 104.275 181.810 ;
        RECT 107.665 181.950 107.955 181.995 ;
        RECT 110.870 181.950 111.190 182.010 ;
        RECT 107.665 181.810 111.190 181.950 ;
        RECT 107.665 181.765 107.955 181.810 ;
        RECT 110.870 181.750 111.190 181.810 ;
        RECT 113.630 181.750 113.950 182.010 ;
        RECT 114.550 181.950 114.870 182.010 ;
        RECT 115.025 181.950 115.315 181.995 ;
        RECT 114.550 181.810 115.315 181.950 ;
        RECT 114.550 181.750 114.870 181.810 ;
        RECT 115.025 181.765 115.315 181.810 ;
        RECT 123.305 181.950 123.595 181.995 ;
        RECT 124.210 181.950 124.530 182.010 ;
        RECT 123.305 181.810 124.530 181.950 ;
        RECT 123.305 181.765 123.595 181.810 ;
        RECT 124.210 181.750 124.530 181.810 ;
        RECT 29.840 181.130 127.820 181.610 ;
        RECT 35.430 180.930 35.750 180.990 ;
        RECT 40.950 180.930 41.270 180.990 ;
        RECT 55.210 180.930 55.530 180.990 ;
        RECT 57.050 180.930 57.370 180.990 ;
        RECT 35.430 180.790 41.270 180.930 ;
        RECT 35.430 180.730 35.750 180.790 ;
        RECT 40.950 180.730 41.270 180.790 ;
        RECT 45.640 180.790 57.370 180.930 ;
        RECT 31.765 180.590 32.055 180.635 ;
        RECT 44.170 180.590 44.490 180.650 ;
        RECT 45.640 180.590 45.780 180.790 ;
        RECT 55.210 180.730 55.530 180.790 ;
        RECT 57.050 180.730 57.370 180.790 ;
        RECT 69.010 180.930 69.330 180.990 ;
        RECT 72.230 180.930 72.550 180.990 ;
        RECT 69.010 180.790 72.550 180.930 ;
        RECT 69.010 180.730 69.330 180.790 ;
        RECT 72.230 180.730 72.550 180.790 ;
        RECT 74.530 180.730 74.850 180.990 ;
        RECT 87.410 180.930 87.730 180.990 ;
        RECT 98.450 180.930 98.770 180.990 ;
        RECT 81.980 180.790 87.730 180.930 ;
        RECT 31.765 180.450 44.490 180.590 ;
        RECT 31.765 180.405 32.055 180.450 ;
        RECT 44.170 180.390 44.490 180.450 ;
        RECT 45.180 180.450 45.780 180.590 ;
        RECT 46.025 180.590 46.315 180.635 ;
        RECT 48.310 180.590 48.630 180.650 ;
        RECT 46.025 180.450 48.630 180.590 ;
        RECT 42.790 180.250 43.110 180.310 ;
        RECT 33.680 180.110 43.110 180.250 ;
        RECT 33.680 179.955 33.820 180.110 ;
        RECT 33.145 179.725 33.435 179.955 ;
        RECT 33.605 179.725 33.895 179.955 ;
        RECT 34.065 179.725 34.355 179.955 ;
        RECT 34.985 179.910 35.275 179.955 ;
        RECT 35.445 179.910 35.735 179.955 ;
        RECT 35.890 179.910 36.210 179.970 ;
        RECT 34.985 179.770 36.210 179.910 ;
        RECT 34.985 179.725 35.275 179.770 ;
        RECT 35.445 179.725 35.735 179.770 ;
        RECT 33.220 179.570 33.360 179.725 ;
        RECT 34.140 179.570 34.280 179.725 ;
        RECT 35.890 179.710 36.210 179.770 ;
        RECT 36.350 179.710 36.670 179.970 ;
        RECT 36.900 179.955 37.040 180.110 ;
        RECT 36.825 179.725 37.115 179.955 ;
        RECT 37.285 179.910 37.575 179.955 ;
        RECT 37.730 179.910 38.050 179.970 ;
        RECT 40.490 179.910 40.810 179.970 ;
        RECT 41.040 179.955 41.180 180.110 ;
        RECT 42.790 180.050 43.110 180.110 ;
        RECT 43.250 180.050 43.570 180.310 ;
        RECT 37.285 179.770 40.810 179.910 ;
        RECT 37.285 179.725 37.575 179.770 ;
        RECT 37.730 179.710 38.050 179.770 ;
        RECT 40.490 179.710 40.810 179.770 ;
        RECT 40.965 179.725 41.255 179.955 ;
        RECT 41.410 179.710 41.730 179.970 ;
        RECT 42.345 179.910 42.635 179.955 ;
        RECT 45.180 179.910 45.320 180.450 ;
        RECT 46.025 180.405 46.315 180.450 ;
        RECT 48.310 180.390 48.630 180.450 ;
        RECT 49.690 180.390 50.010 180.650 ;
        RECT 56.130 180.590 56.450 180.650 ;
        RECT 61.190 180.590 61.510 180.650 ;
        RECT 71.785 180.590 72.075 180.635 ;
        RECT 74.990 180.590 75.310 180.650 ;
        RECT 52.540 180.450 56.450 180.590 ;
        RECT 45.550 180.250 45.870 180.310 ;
        RECT 52.540 180.250 52.680 180.450 ;
        RECT 56.130 180.390 56.450 180.450 ;
        RECT 57.140 180.450 71.540 180.590 ;
        RECT 45.550 180.110 49.000 180.250 ;
        RECT 45.550 180.050 45.870 180.110 ;
        RECT 46.485 179.910 46.775 179.955 ;
        RECT 42.345 179.770 46.775 179.910 ;
        RECT 42.345 179.725 42.635 179.770 ;
        RECT 46.485 179.725 46.775 179.770 ;
        RECT 47.405 179.725 47.695 179.955 ;
        RECT 47.865 179.725 48.155 179.955 ;
        RECT 48.325 179.725 48.615 179.955 ;
        RECT 48.860 179.910 49.000 180.110 ;
        RECT 50.240 180.110 51.760 180.250 ;
        RECT 50.240 179.910 50.380 180.110 ;
        RECT 48.860 179.770 50.380 179.910 ;
        RECT 50.625 179.910 50.915 179.955 ;
        RECT 51.070 179.910 51.390 179.970 ;
        RECT 51.620 179.955 51.760 180.110 ;
        RECT 52.080 180.110 52.680 180.250 ;
        RECT 53.370 180.250 53.690 180.310 ;
        RECT 53.370 180.110 56.820 180.250 ;
        RECT 52.080 179.970 52.220 180.110 ;
        RECT 53.370 180.050 53.690 180.110 ;
        RECT 50.625 179.770 51.390 179.910 ;
        RECT 50.625 179.725 50.915 179.770 ;
        RECT 38.190 179.570 38.510 179.630 ;
        RECT 33.220 179.430 33.820 179.570 ;
        RECT 34.140 179.430 38.510 179.570 ;
        RECT 33.680 179.230 33.820 179.430 ;
        RECT 38.190 179.370 38.510 179.430 ;
        RECT 38.665 179.570 38.955 179.615 ;
        RECT 46.010 179.570 46.330 179.630 ;
        RECT 47.480 179.570 47.620 179.725 ;
        RECT 38.665 179.430 42.560 179.570 ;
        RECT 38.665 179.385 38.955 179.430 ;
        RECT 42.420 179.290 42.560 179.430 ;
        RECT 46.010 179.430 47.620 179.570 ;
        RECT 46.010 179.370 46.330 179.430 ;
        RECT 37.730 179.230 38.050 179.290 ;
        RECT 33.680 179.090 38.050 179.230 ;
        RECT 37.730 179.030 38.050 179.090 ;
        RECT 39.125 179.230 39.415 179.275 ;
        RECT 41.410 179.230 41.730 179.290 ;
        RECT 39.125 179.090 41.730 179.230 ;
        RECT 39.125 179.045 39.415 179.090 ;
        RECT 41.410 179.030 41.730 179.090 ;
        RECT 42.330 179.030 42.650 179.290 ;
        RECT 47.940 179.230 48.080 179.725 ;
        RECT 48.400 179.570 48.540 179.725 ;
        RECT 51.070 179.710 51.390 179.770 ;
        RECT 51.545 179.725 51.835 179.955 ;
        RECT 51.990 179.710 52.310 179.970 ;
        RECT 52.465 179.910 52.755 179.955 ;
        RECT 55.685 179.910 55.975 179.955 ;
        RECT 52.465 179.770 55.975 179.910 ;
        RECT 52.465 179.725 52.755 179.770 ;
        RECT 55.685 179.725 55.975 179.770 ;
        RECT 52.540 179.570 52.680 179.725 ;
        RECT 48.400 179.430 52.680 179.570 ;
        RECT 55.760 179.570 55.900 179.725 ;
        RECT 56.130 179.710 56.450 179.970 ;
        RECT 56.680 179.955 56.820 180.110 ;
        RECT 56.605 179.725 56.895 179.955 ;
        RECT 57.140 179.570 57.280 180.450 ;
        RECT 61.190 180.390 61.510 180.450 ;
        RECT 60.730 180.250 61.050 180.310 ;
        RECT 61.665 180.250 61.955 180.295 ;
        RECT 60.730 180.110 61.955 180.250 ;
        RECT 60.730 180.050 61.050 180.110 ;
        RECT 61.665 180.065 61.955 180.110 ;
        RECT 57.510 179.710 57.830 179.970 ;
        RECT 61.205 179.910 61.495 179.955 ;
        RECT 63.950 179.910 64.270 179.970 ;
        RECT 61.205 179.770 64.270 179.910 ;
        RECT 67.720 179.910 67.860 180.450 ;
        RECT 68.090 180.250 68.410 180.310 ;
        RECT 69.930 180.250 70.250 180.310 ;
        RECT 71.400 180.250 71.540 180.450 ;
        RECT 71.785 180.450 75.310 180.590 ;
        RECT 71.785 180.405 72.075 180.450 ;
        RECT 74.990 180.390 75.310 180.450 ;
        RECT 76.845 180.590 77.135 180.635 ;
        RECT 78.670 180.590 78.990 180.650 ;
        RECT 76.845 180.450 78.990 180.590 ;
        RECT 76.845 180.405 77.135 180.450 ;
        RECT 76.920 180.250 77.060 180.405 ;
        RECT 78.670 180.390 78.990 180.450 ;
        RECT 78.210 180.250 78.530 180.310 ;
        RECT 68.090 180.110 69.700 180.250 ;
        RECT 68.090 180.050 68.410 180.110 ;
        RECT 68.565 179.910 68.855 179.955 ;
        RECT 67.720 179.770 68.855 179.910 ;
        RECT 61.205 179.725 61.495 179.770 ;
        RECT 63.950 179.710 64.270 179.770 ;
        RECT 68.565 179.725 68.855 179.770 ;
        RECT 69.010 179.710 69.330 179.970 ;
        RECT 69.560 179.955 69.700 180.110 ;
        RECT 69.930 180.110 71.080 180.250 ;
        RECT 71.400 180.110 77.060 180.250 ;
        RECT 77.380 180.110 78.530 180.250 ;
        RECT 69.930 180.050 70.250 180.110 ;
        RECT 70.940 179.955 71.080 180.110 ;
        RECT 69.485 179.725 69.775 179.955 ;
        RECT 70.405 179.725 70.695 179.955 ;
        RECT 70.865 179.725 71.155 179.955 ;
        RECT 55.760 179.430 57.280 179.570 ;
        RECT 57.600 179.570 57.740 179.710 ;
        RECT 70.480 179.570 70.620 179.725 ;
        RECT 73.610 179.710 73.930 179.970 ;
        RECT 74.070 179.910 74.390 179.970 ;
        RECT 75.465 179.910 75.755 179.955 ;
        RECT 76.370 179.910 76.690 179.970 ;
        RECT 77.380 179.910 77.520 180.110 ;
        RECT 78.210 180.050 78.530 180.110 ;
        RECT 80.985 180.250 81.275 180.295 ;
        RECT 81.980 180.250 82.120 180.790 ;
        RECT 87.410 180.730 87.730 180.790 ;
        RECT 95.320 180.790 98.770 180.930 ;
        RECT 84.650 180.590 84.970 180.650 ;
        RECT 80.985 180.110 82.120 180.250 ;
        RECT 82.440 180.450 84.970 180.590 ;
        RECT 80.985 180.065 81.275 180.110 ;
        RECT 74.070 179.770 77.520 179.910 ;
        RECT 74.070 179.710 74.390 179.770 ;
        RECT 75.465 179.725 75.755 179.770 ;
        RECT 76.370 179.710 76.690 179.770 ;
        RECT 77.750 179.710 78.070 179.970 ;
        RECT 79.605 179.910 79.895 179.955 ;
        RECT 81.890 179.910 82.210 179.970 ;
        RECT 82.440 179.955 82.580 180.450 ;
        RECT 84.650 180.390 84.970 180.450 ;
        RECT 90.140 180.590 90.430 180.635 ;
        RECT 92.920 180.590 93.210 180.635 ;
        RECT 94.780 180.590 95.070 180.635 ;
        RECT 90.140 180.450 95.070 180.590 ;
        RECT 90.140 180.405 90.430 180.450 ;
        RECT 92.920 180.405 93.210 180.450 ;
        RECT 94.780 180.405 95.070 180.450 ;
        RECT 82.810 180.250 83.130 180.310 ;
        RECT 87.410 180.250 87.730 180.310 ;
        RECT 93.405 180.250 93.695 180.295 ;
        RECT 94.310 180.250 94.630 180.310 ;
        RECT 95.320 180.295 95.460 180.790 ;
        RECT 98.450 180.730 98.770 180.790 ;
        RECT 106.730 180.930 107.050 180.990 ;
        RECT 111.330 180.930 111.650 180.990 ;
        RECT 112.710 180.930 113.030 180.990 ;
        RECT 106.730 180.790 113.030 180.930 ;
        RECT 106.730 180.730 107.050 180.790 ;
        RECT 111.330 180.730 111.650 180.790 ;
        RECT 112.710 180.730 113.030 180.790 ;
        RECT 97.530 180.390 97.850 180.650 ;
        RECT 115.010 180.590 115.330 180.650 ;
        RECT 106.820 180.450 115.330 180.590 ;
        RECT 82.810 180.110 84.420 180.250 ;
        RECT 82.810 180.050 83.130 180.110 ;
        RECT 79.605 179.770 82.210 179.910 ;
        RECT 79.605 179.725 79.895 179.770 ;
        RECT 81.890 179.710 82.210 179.770 ;
        RECT 82.365 179.725 82.655 179.955 ;
        RECT 83.285 179.725 83.575 179.955 ;
        RECT 82.440 179.570 82.580 179.725 ;
        RECT 57.600 179.430 82.580 179.570 ;
        RECT 83.360 179.570 83.500 179.725 ;
        RECT 83.730 179.710 84.050 179.970 ;
        RECT 84.280 179.955 84.420 180.110 ;
        RECT 87.410 180.110 93.160 180.250 ;
        RECT 87.410 180.050 87.730 180.110 ;
        RECT 84.205 179.725 84.495 179.955 ;
        RECT 90.140 179.910 90.430 179.955 ;
        RECT 93.020 179.910 93.160 180.110 ;
        RECT 93.405 180.110 94.630 180.250 ;
        RECT 93.405 180.065 93.695 180.110 ;
        RECT 94.310 180.050 94.630 180.110 ;
        RECT 95.245 180.065 95.535 180.295 ;
        RECT 97.620 180.250 97.760 180.390 ;
        RECT 104.430 180.250 104.750 180.310 ;
        RECT 95.780 180.110 104.750 180.250 ;
        RECT 95.780 179.955 95.920 180.110 ;
        RECT 104.430 180.050 104.750 180.110 ;
        RECT 95.705 179.910 95.995 179.955 ;
        RECT 90.140 179.770 92.675 179.910 ;
        RECT 93.020 179.770 95.995 179.910 ;
        RECT 90.140 179.725 90.430 179.770 ;
        RECT 84.650 179.570 84.970 179.630 ;
        RECT 88.280 179.570 88.570 179.615 ;
        RECT 89.710 179.570 90.030 179.630 ;
        RECT 92.460 179.615 92.675 179.770 ;
        RECT 95.705 179.725 95.995 179.770 ;
        RECT 97.530 179.910 97.850 179.970 ;
        RECT 98.005 179.910 98.295 179.955 ;
        RECT 97.530 179.770 98.295 179.910 ;
        RECT 97.530 179.710 97.850 179.770 ;
        RECT 98.005 179.725 98.295 179.770 ;
        RECT 102.130 179.710 102.450 179.970 ;
        RECT 105.825 179.910 106.115 179.955 ;
        RECT 106.270 179.910 106.590 179.970 ;
        RECT 106.820 179.955 106.960 180.450 ;
        RECT 115.010 180.390 115.330 180.450 ;
        RECT 116.865 180.590 117.155 180.635 ;
        RECT 118.690 180.590 119.010 180.650 ;
        RECT 116.865 180.450 119.010 180.590 ;
        RECT 116.865 180.405 117.155 180.450 ;
        RECT 118.690 180.390 119.010 180.450 ;
        RECT 119.725 180.590 120.015 180.635 ;
        RECT 122.845 180.590 123.135 180.635 ;
        RECT 124.735 180.590 125.025 180.635 ;
        RECT 119.725 180.450 125.025 180.590 ;
        RECT 119.725 180.405 120.015 180.450 ;
        RECT 122.845 180.405 123.135 180.450 ;
        RECT 124.735 180.405 125.025 180.450 ;
        RECT 110.410 180.250 110.730 180.310 ;
        RECT 113.645 180.250 113.935 180.295 ;
        RECT 116.390 180.250 116.710 180.310 ;
        RECT 110.410 180.110 112.020 180.250 ;
        RECT 110.410 180.050 110.730 180.110 ;
        RECT 105.825 179.770 106.590 179.910 ;
        RECT 105.825 179.725 106.115 179.770 ;
        RECT 106.270 179.710 106.590 179.770 ;
        RECT 106.745 179.725 107.035 179.955 ;
        RECT 107.205 179.725 107.495 179.955 ;
        RECT 107.665 179.910 107.955 179.955 ;
        RECT 109.030 179.910 109.350 179.970 ;
        RECT 111.880 179.955 112.020 180.110 ;
        RECT 113.645 180.110 116.710 180.250 ;
        RECT 113.645 180.065 113.935 180.110 ;
        RECT 116.390 180.050 116.710 180.110 ;
        RECT 124.210 180.050 124.530 180.310 ;
        RECT 110.885 179.910 111.175 179.955 ;
        RECT 107.665 179.770 111.175 179.910 ;
        RECT 107.665 179.725 107.955 179.770 ;
        RECT 91.540 179.570 91.830 179.615 ;
        RECT 83.360 179.430 84.970 179.570 ;
        RECT 84.650 179.370 84.970 179.430 ;
        RECT 85.200 179.430 88.100 179.570 ;
        RECT 51.990 179.230 52.310 179.290 ;
        RECT 47.940 179.090 52.310 179.230 ;
        RECT 51.990 179.030 52.310 179.090 ;
        RECT 53.370 179.230 53.690 179.290 ;
        RECT 53.845 179.230 54.135 179.275 ;
        RECT 53.370 179.090 54.135 179.230 ;
        RECT 53.370 179.030 53.690 179.090 ;
        RECT 53.845 179.045 54.135 179.090 ;
        RECT 54.290 179.030 54.610 179.290 ;
        RECT 57.985 179.230 58.275 179.275 ;
        RECT 60.270 179.230 60.590 179.290 ;
        RECT 57.985 179.090 60.590 179.230 ;
        RECT 57.985 179.045 58.275 179.090 ;
        RECT 60.270 179.030 60.590 179.090 ;
        RECT 64.870 179.030 65.190 179.290 ;
        RECT 66.250 179.230 66.570 179.290 ;
        RECT 67.185 179.230 67.475 179.275 ;
        RECT 66.250 179.090 67.475 179.230 ;
        RECT 66.250 179.030 66.570 179.090 ;
        RECT 67.185 179.045 67.475 179.090 ;
        RECT 67.630 179.230 67.950 179.290 ;
        RECT 72.705 179.230 72.995 179.275 ;
        RECT 85.200 179.230 85.340 179.430 ;
        RECT 67.630 179.090 85.340 179.230 ;
        RECT 67.630 179.030 67.950 179.090 ;
        RECT 72.705 179.045 72.995 179.090 ;
        RECT 85.570 179.030 85.890 179.290 ;
        RECT 86.275 179.230 86.565 179.275 ;
        RECT 86.950 179.230 87.270 179.290 ;
        RECT 86.275 179.090 87.270 179.230 ;
        RECT 87.960 179.230 88.100 179.430 ;
        RECT 88.280 179.430 91.830 179.570 ;
        RECT 88.280 179.385 88.570 179.430 ;
        RECT 89.710 179.370 90.030 179.430 ;
        RECT 91.540 179.385 91.830 179.430 ;
        RECT 92.460 179.570 92.750 179.615 ;
        RECT 94.320 179.570 94.610 179.615 ;
        RECT 107.280 179.570 107.420 179.725 ;
        RECT 109.030 179.710 109.350 179.770 ;
        RECT 110.885 179.725 111.175 179.770 ;
        RECT 111.345 179.725 111.635 179.955 ;
        RECT 111.805 179.725 112.095 179.955 ;
        RECT 111.420 179.570 111.560 179.725 ;
        RECT 112.710 179.710 113.030 179.970 ;
        RECT 92.460 179.430 94.610 179.570 ;
        RECT 92.460 179.385 92.750 179.430 ;
        RECT 94.320 179.385 94.610 179.430 ;
        RECT 95.780 179.430 111.560 179.570 ;
        RECT 113.630 179.570 113.950 179.630 ;
        RECT 118.645 179.615 118.935 179.930 ;
        RECT 119.725 179.910 120.015 179.955 ;
        RECT 123.305 179.910 123.595 179.955 ;
        RECT 125.140 179.910 125.430 179.955 ;
        RECT 119.725 179.770 125.430 179.910 ;
        RECT 119.725 179.725 120.015 179.770 ;
        RECT 123.305 179.725 123.595 179.770 ;
        RECT 125.140 179.725 125.430 179.770 ;
        RECT 125.605 179.910 125.895 179.955 ;
        RECT 126.050 179.910 126.370 179.970 ;
        RECT 125.605 179.770 126.370 179.910 ;
        RECT 125.605 179.725 125.895 179.770 ;
        RECT 126.050 179.710 126.370 179.770 ;
        RECT 118.345 179.570 118.935 179.615 ;
        RECT 121.585 179.570 122.235 179.615 ;
        RECT 113.630 179.430 122.235 179.570 ;
        RECT 95.780 179.230 95.920 179.430 ;
        RECT 105.900 179.290 106.040 179.430 ;
        RECT 113.630 179.370 113.950 179.430 ;
        RECT 118.345 179.385 118.635 179.430 ;
        RECT 121.585 179.385 122.235 179.430 ;
        RECT 87.960 179.090 95.920 179.230 ;
        RECT 86.275 179.045 86.565 179.090 ;
        RECT 86.950 179.030 87.270 179.090 ;
        RECT 96.150 179.030 96.470 179.290 ;
        RECT 101.210 179.030 101.530 179.290 ;
        RECT 103.065 179.230 103.355 179.275 ;
        RECT 103.970 179.230 104.290 179.290 ;
        RECT 103.065 179.090 104.290 179.230 ;
        RECT 103.065 179.045 103.355 179.090 ;
        RECT 103.970 179.030 104.290 179.090 ;
        RECT 105.810 179.030 106.130 179.290 ;
        RECT 109.030 179.030 109.350 179.290 ;
        RECT 109.505 179.230 109.795 179.275 ;
        RECT 109.950 179.230 110.270 179.290 ;
        RECT 109.505 179.090 110.270 179.230 ;
        RECT 109.505 179.045 109.795 179.090 ;
        RECT 109.950 179.030 110.270 179.090 ;
        RECT 116.405 179.230 116.695 179.275 ;
        RECT 117.310 179.230 117.630 179.290 ;
        RECT 116.405 179.090 117.630 179.230 ;
        RECT 116.405 179.045 116.695 179.090 ;
        RECT 117.310 179.030 117.630 179.090 ;
        RECT 29.840 178.410 127.820 178.890 ;
        RECT 36.365 178.210 36.655 178.255 ;
        RECT 42.790 178.210 43.110 178.270 ;
        RECT 48.770 178.210 49.090 178.270 ;
        RECT 67.630 178.210 67.950 178.270 ;
        RECT 36.365 178.070 41.180 178.210 ;
        RECT 36.365 178.025 36.655 178.070 ;
        RECT 37.270 177.870 37.590 177.930 ;
        RECT 34.600 177.730 37.590 177.870 ;
        RECT 34.600 177.575 34.740 177.730 ;
        RECT 37.270 177.670 37.590 177.730 ;
        RECT 39.110 177.670 39.430 177.930 ;
        RECT 41.040 177.870 41.180 178.070 ;
        RECT 42.790 178.070 67.950 178.210 ;
        RECT 42.790 178.010 43.110 178.070 ;
        RECT 48.770 178.010 49.090 178.070 ;
        RECT 67.630 178.010 67.950 178.070 ;
        RECT 70.390 178.210 70.710 178.270 ;
        RECT 71.325 178.210 71.615 178.255 ;
        RECT 70.390 178.070 71.615 178.210 ;
        RECT 70.390 178.010 70.710 178.070 ;
        RECT 71.325 178.025 71.615 178.070 ;
        RECT 75.450 178.010 75.770 178.270 ;
        RECT 76.370 178.210 76.690 178.270 ;
        RECT 84.665 178.210 84.955 178.255 ;
        RECT 86.490 178.210 86.810 178.270 ;
        RECT 76.370 178.070 82.580 178.210 ;
        RECT 76.370 178.010 76.690 178.070 ;
        RECT 41.405 177.870 42.055 177.915 ;
        RECT 45.005 177.870 45.295 177.915 ;
        RECT 50.610 177.870 50.930 177.930 ;
        RECT 41.040 177.730 45.295 177.870 ;
        RECT 41.405 177.685 42.055 177.730 ;
        RECT 44.705 177.685 45.295 177.730 ;
        RECT 48.300 177.730 50.930 177.870 ;
        RECT 34.525 177.345 34.815 177.575 ;
        RECT 35.430 177.530 35.750 177.590 ;
        RECT 35.905 177.530 36.195 177.575 ;
        RECT 35.430 177.390 36.195 177.530 ;
        RECT 35.430 177.330 35.750 177.390 ;
        RECT 35.905 177.345 36.195 177.390 ;
        RECT 38.210 177.530 38.500 177.575 ;
        RECT 40.045 177.530 40.335 177.575 ;
        RECT 43.625 177.530 43.915 177.575 ;
        RECT 38.210 177.390 43.915 177.530 ;
        RECT 38.210 177.345 38.500 177.390 ;
        RECT 40.045 177.345 40.335 177.390 ;
        RECT 43.625 177.345 43.915 177.390 ;
        RECT 44.705 177.370 44.995 177.685 ;
        RECT 48.300 177.575 48.440 177.730 ;
        RECT 50.610 177.670 50.930 177.730 ;
        RECT 51.990 177.670 52.310 177.930 ;
        RECT 52.450 177.870 52.770 177.930 ;
        RECT 54.285 177.870 54.935 177.915 ;
        RECT 57.885 177.870 58.175 177.915 ;
        RECT 52.450 177.730 58.175 177.870 ;
        RECT 52.450 177.670 52.770 177.730 ;
        RECT 54.285 177.685 54.935 177.730 ;
        RECT 57.585 177.685 58.175 177.730 ;
        RECT 68.550 177.870 68.870 177.930 ;
        RECT 68.550 177.730 77.060 177.870 ;
        RECT 48.300 177.380 48.615 177.575 ;
        RECT 48.325 177.345 48.615 177.380 ;
        RECT 48.770 177.330 49.090 177.590 ;
        RECT 49.230 177.330 49.550 177.590 ;
        RECT 50.150 177.330 50.470 177.590 ;
        RECT 51.090 177.530 51.380 177.575 ;
        RECT 52.925 177.530 53.215 177.575 ;
        RECT 56.505 177.530 56.795 177.575 ;
        RECT 51.090 177.390 56.795 177.530 ;
        RECT 51.090 177.345 51.380 177.390 ;
        RECT 52.925 177.345 53.215 177.390 ;
        RECT 56.505 177.345 56.795 177.390 ;
        RECT 57.585 177.370 57.875 177.685 ;
        RECT 68.550 177.670 68.870 177.730 ;
        RECT 60.270 177.330 60.590 177.590 ;
        RECT 66.710 177.530 67.030 177.590 ;
        RECT 71.785 177.530 72.075 177.575 ;
        RECT 74.990 177.530 75.310 177.590 ;
        RECT 66.710 177.390 75.310 177.530 ;
        RECT 66.710 177.330 67.030 177.390 ;
        RECT 71.785 177.345 72.075 177.390 ;
        RECT 74.990 177.330 75.310 177.390 ;
        RECT 76.370 177.330 76.690 177.590 ;
        RECT 76.920 177.530 77.060 177.730 ;
        RECT 77.290 177.670 77.610 177.930 ;
        RECT 79.145 177.870 79.435 177.915 ;
        RECT 81.890 177.870 82.210 177.930 ;
        RECT 79.145 177.730 82.210 177.870 ;
        RECT 79.145 177.685 79.435 177.730 ;
        RECT 79.220 177.530 79.360 177.685 ;
        RECT 81.890 177.670 82.210 177.730 ;
        RECT 76.920 177.390 79.360 177.530 ;
        RECT 79.590 177.330 79.910 177.590 ;
        RECT 80.065 177.530 80.355 177.575 ;
        RECT 80.510 177.530 80.830 177.590 ;
        RECT 80.065 177.390 80.830 177.530 ;
        RECT 80.065 177.345 80.355 177.390 ;
        RECT 80.510 177.330 80.830 177.390 ;
        RECT 81.445 177.530 81.735 177.575 ;
        RECT 82.440 177.530 82.580 178.070 ;
        RECT 84.665 178.070 86.810 178.210 ;
        RECT 84.665 178.025 84.955 178.070 ;
        RECT 86.490 178.010 86.810 178.070 ;
        RECT 89.710 178.010 90.030 178.270 ;
        RECT 94.310 178.010 94.630 178.270 ;
        RECT 100.750 178.210 101.070 178.270 ;
        RECT 112.265 178.210 112.555 178.255 ;
        RECT 100.750 178.070 112.555 178.210 ;
        RECT 100.750 178.010 101.070 178.070 ;
        RECT 112.265 178.025 112.555 178.070 ;
        RECT 114.105 178.210 114.395 178.255 ;
        RECT 119.150 178.210 119.470 178.270 ;
        RECT 114.105 178.070 119.470 178.210 ;
        RECT 114.105 178.025 114.395 178.070 ;
        RECT 119.150 178.010 119.470 178.070 ;
        RECT 95.690 177.870 96.010 177.930 ;
        RECT 89.340 177.730 96.010 177.870 ;
        RECT 81.445 177.390 82.580 177.530 ;
        RECT 86.030 177.530 86.350 177.590 ;
        RECT 89.340 177.575 89.480 177.730 ;
        RECT 95.690 177.670 96.010 177.730 ;
        RECT 96.150 177.870 96.470 177.930 ;
        RECT 98.105 177.870 98.395 177.915 ;
        RECT 101.345 177.870 101.995 177.915 ;
        RECT 96.150 177.730 101.995 177.870 ;
        RECT 96.150 177.670 96.470 177.730 ;
        RECT 98.105 177.685 98.695 177.730 ;
        RECT 101.345 177.685 101.995 177.730 ;
        RECT 87.425 177.530 87.715 177.575 ;
        RECT 86.030 177.390 87.715 177.530 ;
        RECT 81.445 177.345 81.735 177.390 ;
        RECT 86.030 177.330 86.350 177.390 ;
        RECT 87.425 177.345 87.715 177.390 ;
        RECT 89.265 177.345 89.555 177.575 ;
        RECT 90.170 177.530 90.490 177.590 ;
        RECT 90.645 177.530 90.935 177.575 ;
        RECT 90.170 177.390 90.935 177.530 ;
        RECT 90.170 177.330 90.490 177.390 ;
        RECT 90.645 177.345 90.935 177.390 ;
        RECT 95.245 177.345 95.535 177.575 ;
        RECT 97.070 177.530 97.390 177.590 ;
        RECT 95.780 177.390 97.390 177.530 ;
        RECT 37.745 177.190 38.035 177.235 ;
        RECT 39.570 177.190 39.890 177.250 ;
        RECT 50.625 177.190 50.915 177.235 ;
        RECT 59.365 177.190 59.655 177.235 ;
        RECT 63.965 177.190 64.255 177.235 ;
        RECT 67.630 177.190 67.950 177.250 ;
        RECT 37.745 177.050 57.740 177.190 ;
        RECT 37.745 177.005 38.035 177.050 ;
        RECT 39.570 176.990 39.890 177.050 ;
        RECT 50.625 177.005 50.915 177.050 ;
        RECT 57.600 176.910 57.740 177.050 ;
        RECT 59.365 177.050 67.950 177.190 ;
        RECT 59.365 177.005 59.655 177.050 ;
        RECT 63.965 177.005 64.255 177.050 ;
        RECT 67.630 176.990 67.950 177.050 ;
        RECT 79.130 177.190 79.450 177.250 ;
        RECT 80.985 177.190 81.275 177.235 ;
        RECT 82.810 177.190 83.130 177.250 ;
        RECT 79.130 177.050 83.130 177.190 ;
        RECT 79.130 176.990 79.450 177.050 ;
        RECT 80.985 177.005 81.275 177.050 ;
        RECT 82.810 176.990 83.130 177.050 ;
        RECT 88.330 177.190 88.650 177.250 ;
        RECT 95.320 177.190 95.460 177.345 ;
        RECT 88.330 177.050 95.460 177.190 ;
        RECT 88.330 176.990 88.650 177.050 ;
        RECT 38.615 176.850 38.905 176.895 ;
        RECT 40.505 176.850 40.795 176.895 ;
        RECT 43.625 176.850 43.915 176.895 ;
        RECT 38.615 176.710 43.915 176.850 ;
        RECT 38.615 176.665 38.905 176.710 ;
        RECT 40.505 176.665 40.795 176.710 ;
        RECT 43.625 176.665 43.915 176.710 ;
        RECT 46.010 176.850 46.330 176.910 ;
        RECT 46.945 176.850 47.235 176.895 ;
        RECT 46.010 176.710 47.235 176.850 ;
        RECT 46.010 176.650 46.330 176.710 ;
        RECT 46.945 176.665 47.235 176.710 ;
        RECT 51.495 176.850 51.785 176.895 ;
        RECT 53.385 176.850 53.675 176.895 ;
        RECT 56.505 176.850 56.795 176.895 ;
        RECT 51.495 176.710 56.795 176.850 ;
        RECT 51.495 176.665 51.785 176.710 ;
        RECT 53.385 176.665 53.675 176.710 ;
        RECT 56.505 176.665 56.795 176.710 ;
        RECT 57.510 176.650 57.830 176.910 ;
        RECT 74.530 176.850 74.850 176.910 ;
        RECT 93.865 176.850 94.155 176.895 ;
        RECT 95.780 176.850 95.920 177.390 ;
        RECT 97.070 177.330 97.390 177.390 ;
        RECT 98.405 177.370 98.695 177.685 ;
        RECT 103.970 177.670 104.290 177.930 ;
        RECT 104.430 177.870 104.750 177.930 ;
        RECT 115.485 177.870 115.775 177.915 ;
        RECT 117.885 177.870 118.175 177.915 ;
        RECT 121.125 177.870 121.775 177.915 ;
        RECT 104.430 177.730 106.040 177.870 ;
        RECT 104.430 177.670 104.750 177.730 ;
        RECT 105.900 177.575 106.040 177.730 ;
        RECT 115.485 177.730 121.775 177.870 ;
        RECT 115.485 177.685 115.775 177.730 ;
        RECT 117.885 177.685 118.475 177.730 ;
        RECT 121.125 177.685 121.775 177.730 ;
        RECT 123.765 177.870 124.055 177.915 ;
        RECT 124.210 177.870 124.530 177.930 ;
        RECT 123.765 177.730 124.530 177.870 ;
        RECT 123.765 177.685 124.055 177.730 ;
        RECT 99.485 177.530 99.775 177.575 ;
        RECT 103.065 177.530 103.355 177.575 ;
        RECT 104.900 177.530 105.190 177.575 ;
        RECT 99.485 177.390 105.190 177.530 ;
        RECT 99.485 177.345 99.775 177.390 ;
        RECT 103.065 177.345 103.355 177.390 ;
        RECT 104.900 177.345 105.190 177.390 ;
        RECT 105.825 177.530 106.115 177.575 ;
        RECT 115.025 177.530 115.315 177.575 ;
        RECT 115.930 177.530 116.250 177.590 ;
        RECT 105.825 177.390 116.250 177.530 ;
        RECT 105.825 177.345 106.115 177.390 ;
        RECT 115.025 177.345 115.315 177.390 ;
        RECT 115.930 177.330 116.250 177.390 ;
        RECT 118.185 177.370 118.475 177.685 ;
        RECT 124.210 177.670 124.530 177.730 ;
        RECT 119.265 177.530 119.555 177.575 ;
        RECT 122.845 177.530 123.135 177.575 ;
        RECT 124.680 177.530 124.970 177.575 ;
        RECT 119.265 177.390 124.970 177.530 ;
        RECT 119.265 177.345 119.555 177.390 ;
        RECT 122.845 177.345 123.135 177.390 ;
        RECT 124.680 177.345 124.970 177.390 ;
        RECT 58.060 176.710 93.620 176.850 ;
        RECT 35.445 176.510 35.735 176.555 ;
        RECT 41.870 176.510 42.190 176.570 ;
        RECT 35.445 176.370 42.190 176.510 ;
        RECT 35.445 176.325 35.735 176.370 ;
        RECT 41.870 176.310 42.190 176.370 ;
        RECT 45.090 176.510 45.410 176.570 ;
        RECT 46.485 176.510 46.775 176.555 ;
        RECT 45.090 176.370 46.775 176.510 ;
        RECT 45.090 176.310 45.410 176.370 ;
        RECT 46.485 176.325 46.775 176.370 ;
        RECT 50.150 176.510 50.470 176.570 ;
        RECT 52.910 176.510 53.230 176.570 ;
        RECT 58.060 176.510 58.200 176.710 ;
        RECT 74.530 176.650 74.850 176.710 ;
        RECT 50.150 176.370 58.200 176.510 ;
        RECT 50.150 176.310 50.470 176.370 ;
        RECT 52.910 176.310 53.230 176.370 ;
        RECT 61.190 176.310 61.510 176.570 ;
        RECT 66.725 176.510 67.015 176.555 ;
        RECT 68.090 176.510 68.410 176.570 ;
        RECT 66.725 176.370 68.410 176.510 ;
        RECT 66.725 176.325 67.015 176.370 ;
        RECT 68.090 176.310 68.410 176.370 ;
        RECT 76.370 176.510 76.690 176.570 ;
        RECT 80.525 176.510 80.815 176.555 ;
        RECT 76.370 176.370 80.815 176.510 ;
        RECT 93.480 176.510 93.620 176.710 ;
        RECT 93.865 176.710 95.920 176.850 ;
        RECT 96.240 177.050 105.120 177.190 ;
        RECT 93.865 176.665 94.155 176.710 ;
        RECT 96.240 176.510 96.380 177.050 ;
        RECT 99.485 176.850 99.775 176.895 ;
        RECT 102.605 176.850 102.895 176.895 ;
        RECT 104.495 176.850 104.785 176.895 ;
        RECT 99.485 176.710 104.785 176.850 ;
        RECT 104.980 176.850 105.120 177.050 ;
        RECT 105.350 176.990 105.670 177.250 ;
        RECT 106.270 176.990 106.590 177.250 ;
        RECT 111.330 176.990 111.650 177.250 ;
        RECT 111.805 177.190 112.095 177.235 ;
        RECT 117.770 177.190 118.090 177.250 ;
        RECT 111.805 177.050 118.090 177.190 ;
        RECT 111.805 177.005 112.095 177.050 ;
        RECT 117.770 176.990 118.090 177.050 ;
        RECT 125.145 177.190 125.435 177.235 ;
        RECT 126.050 177.190 126.370 177.250 ;
        RECT 125.145 177.050 126.370 177.190 ;
        RECT 125.145 177.005 125.435 177.050 ;
        RECT 126.050 176.990 126.370 177.050 ;
        RECT 106.360 176.850 106.500 176.990 ;
        RECT 104.980 176.710 106.500 176.850 ;
        RECT 119.265 176.850 119.555 176.895 ;
        RECT 122.385 176.850 122.675 176.895 ;
        RECT 124.275 176.850 124.565 176.895 ;
        RECT 119.265 176.710 124.565 176.850 ;
        RECT 99.485 176.665 99.775 176.710 ;
        RECT 102.605 176.665 102.895 176.710 ;
        RECT 104.495 176.665 104.785 176.710 ;
        RECT 119.265 176.665 119.555 176.710 ;
        RECT 122.385 176.665 122.675 176.710 ;
        RECT 124.275 176.665 124.565 176.710 ;
        RECT 93.480 176.370 96.380 176.510 ;
        RECT 96.625 176.510 96.915 176.555 ;
        RECT 97.530 176.510 97.850 176.570 ;
        RECT 96.625 176.370 97.850 176.510 ;
        RECT 76.370 176.310 76.690 176.370 ;
        RECT 80.525 176.325 80.815 176.370 ;
        RECT 96.625 176.325 96.915 176.370 ;
        RECT 97.530 176.310 97.850 176.370 ;
        RECT 106.270 176.310 106.590 176.570 ;
        RECT 116.390 176.310 116.710 176.570 ;
        RECT 29.840 175.690 127.820 176.170 ;
        RECT 38.650 175.490 38.970 175.550 ;
        RECT 45.105 175.490 45.395 175.535 ;
        RECT 38.650 175.350 45.395 175.490 ;
        RECT 38.650 175.290 38.970 175.350 ;
        RECT 45.105 175.305 45.395 175.350 ;
        RECT 49.245 175.490 49.535 175.535 ;
        RECT 52.450 175.490 52.770 175.550 ;
        RECT 49.245 175.350 52.770 175.490 ;
        RECT 49.245 175.305 49.535 175.350 ;
        RECT 52.450 175.290 52.770 175.350 ;
        RECT 57.510 175.490 57.830 175.550 ;
        RECT 63.045 175.490 63.335 175.535 ;
        RECT 63.950 175.490 64.270 175.550 ;
        RECT 57.510 175.350 62.800 175.490 ;
        RECT 57.510 175.290 57.830 175.350 ;
        RECT 35.400 175.150 35.690 175.195 ;
        RECT 38.180 175.150 38.470 175.195 ;
        RECT 40.040 175.150 40.330 175.195 ;
        RECT 35.400 175.010 40.330 175.150 ;
        RECT 35.400 174.965 35.690 175.010 ;
        RECT 38.180 174.965 38.470 175.010 ;
        RECT 40.040 174.965 40.330 175.010 ;
        RECT 56.705 175.150 56.995 175.195 ;
        RECT 59.825 175.150 60.115 175.195 ;
        RECT 61.715 175.150 62.005 175.195 ;
        RECT 56.705 175.010 62.005 175.150 ;
        RECT 56.705 174.965 56.995 175.010 ;
        RECT 59.825 174.965 60.115 175.010 ;
        RECT 61.715 174.965 62.005 175.010 ;
        RECT 35.890 174.810 36.210 174.870 ;
        RECT 39.570 174.810 39.890 174.870 ;
        RECT 40.505 174.810 40.795 174.855 ;
        RECT 35.890 174.670 39.340 174.810 ;
        RECT 35.890 174.610 36.210 174.670 ;
        RECT 35.400 174.470 35.690 174.515 ;
        RECT 35.400 174.330 37.935 174.470 ;
        RECT 35.400 174.285 35.690 174.330 ;
        RECT 33.540 174.130 33.830 174.175 ;
        RECT 35.890 174.130 36.210 174.190 ;
        RECT 37.720 174.175 37.935 174.330 ;
        RECT 38.650 174.270 38.970 174.530 ;
        RECT 39.200 174.470 39.340 174.670 ;
        RECT 39.570 174.670 40.795 174.810 ;
        RECT 39.570 174.610 39.890 174.670 ;
        RECT 40.505 174.625 40.795 174.670 ;
        RECT 40.950 174.810 41.270 174.870 ;
        RECT 46.470 174.810 46.790 174.870 ;
        RECT 47.865 174.810 48.155 174.855 ;
        RECT 57.970 174.810 58.290 174.870 ;
        RECT 40.950 174.670 46.240 174.810 ;
        RECT 40.950 174.610 41.270 174.670 ;
        RECT 44.645 174.470 44.935 174.515 ;
        RECT 45.090 174.470 45.410 174.530 ;
        RECT 39.200 174.330 40.260 174.470 ;
        RECT 36.800 174.130 37.090 174.175 ;
        RECT 33.540 173.990 37.090 174.130 ;
        RECT 33.540 173.945 33.830 173.990 ;
        RECT 35.890 173.930 36.210 173.990 ;
        RECT 36.800 173.945 37.090 173.990 ;
        RECT 37.720 174.130 38.010 174.175 ;
        RECT 39.580 174.130 39.870 174.175 ;
        RECT 37.720 173.990 39.870 174.130 ;
        RECT 40.120 174.130 40.260 174.330 ;
        RECT 44.645 174.330 45.410 174.470 ;
        RECT 46.100 174.470 46.240 174.670 ;
        RECT 46.470 174.670 48.155 174.810 ;
        RECT 46.470 174.610 46.790 174.670 ;
        RECT 47.865 174.625 48.155 174.670 ;
        RECT 52.540 174.670 58.290 174.810 ;
        RECT 52.540 174.515 52.680 174.670 ;
        RECT 57.970 174.610 58.290 174.670 ;
        RECT 61.190 174.610 61.510 174.870 ;
        RECT 62.660 174.855 62.800 175.350 ;
        RECT 63.045 175.350 64.270 175.490 ;
        RECT 63.045 175.305 63.335 175.350 ;
        RECT 63.950 175.290 64.270 175.350 ;
        RECT 86.030 175.490 86.350 175.550 ;
        RECT 86.950 175.490 87.270 175.550 ;
        RECT 100.765 175.490 101.055 175.535 ;
        RECT 102.130 175.490 102.450 175.550 ;
        RECT 86.030 175.350 94.540 175.490 ;
        RECT 86.030 175.290 86.350 175.350 ;
        RECT 86.950 175.290 87.270 175.350 ;
        RECT 75.450 175.150 75.770 175.210 ;
        RECT 89.220 175.150 89.510 175.195 ;
        RECT 92.000 175.150 92.290 175.195 ;
        RECT 93.860 175.150 94.150 175.195 ;
        RECT 75.450 175.010 89.020 175.150 ;
        RECT 75.450 174.950 75.770 175.010 ;
        RECT 62.585 174.625 62.875 174.855 ;
        RECT 63.490 174.810 63.810 174.870 ;
        RECT 66.265 174.810 66.555 174.855 ;
        RECT 69.930 174.810 70.250 174.870 ;
        RECT 74.085 174.810 74.375 174.855 ;
        RECT 63.490 174.670 66.020 174.810 ;
        RECT 63.490 174.610 63.810 174.670 ;
        RECT 48.785 174.470 49.075 174.515 ;
        RECT 52.465 174.470 52.755 174.515 ;
        RECT 46.100 174.330 52.755 174.470 ;
        RECT 44.645 174.285 44.935 174.330 ;
        RECT 45.090 174.270 45.410 174.330 ;
        RECT 48.785 174.285 49.075 174.330 ;
        RECT 52.465 174.285 52.755 174.330 ;
        RECT 50.150 174.130 50.470 174.190 ;
        RECT 55.625 174.175 55.915 174.490 ;
        RECT 56.705 174.470 56.995 174.515 ;
        RECT 60.285 174.470 60.575 174.515 ;
        RECT 62.120 174.470 62.410 174.515 ;
        RECT 56.705 174.330 62.410 174.470 ;
        RECT 56.705 174.285 56.995 174.330 ;
        RECT 60.285 174.285 60.575 174.330 ;
        RECT 62.120 174.285 62.410 174.330 ;
        RECT 64.870 174.270 65.190 174.530 ;
        RECT 65.345 174.285 65.635 174.515 ;
        RECT 65.880 174.470 66.020 174.670 ;
        RECT 66.265 174.670 70.250 174.810 ;
        RECT 66.265 174.625 66.555 174.670 ;
        RECT 69.930 174.610 70.250 174.670 ;
        RECT 70.940 174.670 74.375 174.810 ;
        RECT 70.940 174.515 71.080 174.670 ;
        RECT 74.085 174.625 74.375 174.670 ;
        RECT 74.990 174.810 75.310 174.870 ;
        RECT 77.765 174.810 78.055 174.855 ;
        RECT 74.990 174.670 78.055 174.810 ;
        RECT 88.880 174.810 89.020 175.010 ;
        RECT 89.220 175.010 94.150 175.150 ;
        RECT 89.220 174.965 89.510 175.010 ;
        RECT 92.000 174.965 92.290 175.010 ;
        RECT 93.860 174.965 94.150 175.010 ;
        RECT 90.170 174.810 90.490 174.870 ;
        RECT 88.880 174.670 90.490 174.810 ;
        RECT 74.990 174.610 75.310 174.670 ;
        RECT 77.765 174.625 78.055 174.670 ;
        RECT 90.170 174.610 90.490 174.670 ;
        RECT 91.090 174.810 91.410 174.870 ;
        RECT 92.485 174.810 92.775 174.855 ;
        RECT 91.090 174.670 92.775 174.810 ;
        RECT 94.400 174.810 94.540 175.350 ;
        RECT 100.765 175.350 102.450 175.490 ;
        RECT 100.765 175.305 101.055 175.350 ;
        RECT 102.130 175.290 102.450 175.350 ;
        RECT 96.165 175.150 96.455 175.195 ;
        RECT 101.670 175.150 101.990 175.210 ;
        RECT 96.165 175.010 101.990 175.150 ;
        RECT 96.165 174.965 96.455 175.010 ;
        RECT 101.670 174.950 101.990 175.010 ;
        RECT 109.145 175.150 109.435 175.195 ;
        RECT 112.265 175.150 112.555 175.195 ;
        RECT 114.155 175.150 114.445 175.195 ;
        RECT 109.145 175.010 114.445 175.150 ;
        RECT 109.145 174.965 109.435 175.010 ;
        RECT 112.265 174.965 112.555 175.010 ;
        RECT 114.155 174.965 114.445 175.010 ;
        RECT 118.690 175.150 119.010 175.210 ;
        RECT 118.690 175.010 123.060 175.150 ;
        RECT 118.690 174.950 119.010 175.010 ;
        RECT 94.400 174.670 96.380 174.810 ;
        RECT 91.090 174.610 91.410 174.670 ;
        RECT 92.485 174.625 92.775 174.670 ;
        RECT 70.865 174.470 71.155 174.515 ;
        RECT 65.880 174.330 71.155 174.470 ;
        RECT 70.865 174.285 71.155 174.330 ;
        RECT 71.325 174.285 71.615 174.515 ;
        RECT 75.465 174.470 75.755 174.515 ;
        RECT 75.910 174.470 76.230 174.530 ;
        RECT 77.290 174.470 77.610 174.530 ;
        RECT 79.130 174.470 79.450 174.530 ;
        RECT 75.465 174.330 79.450 174.470 ;
        RECT 75.465 174.285 75.755 174.330 ;
        RECT 40.120 173.990 50.470 174.130 ;
        RECT 37.720 173.945 38.010 173.990 ;
        RECT 39.580 173.945 39.870 173.990 ;
        RECT 50.150 173.930 50.470 173.990 ;
        RECT 52.925 174.130 53.215 174.175 ;
        RECT 55.325 174.130 55.915 174.175 ;
        RECT 58.565 174.130 59.215 174.175 ;
        RECT 65.420 174.130 65.560 174.285 ;
        RECT 52.925 173.990 59.215 174.130 ;
        RECT 52.925 173.945 53.215 173.990 ;
        RECT 55.325 173.945 55.615 173.990 ;
        RECT 58.565 173.945 59.215 173.990 ;
        RECT 60.360 173.990 65.560 174.130 ;
        RECT 60.360 173.850 60.500 173.990 ;
        RECT 70.390 173.930 70.710 174.190 ;
        RECT 31.535 173.790 31.825 173.835 ;
        RECT 40.030 173.790 40.350 173.850 ;
        RECT 31.535 173.650 40.350 173.790 ;
        RECT 31.535 173.605 31.825 173.650 ;
        RECT 40.030 173.590 40.350 173.650 ;
        RECT 41.425 173.790 41.715 173.835 ;
        RECT 41.870 173.790 42.190 173.850 ;
        RECT 41.425 173.650 42.190 173.790 ;
        RECT 41.425 173.605 41.715 173.650 ;
        RECT 41.870 173.590 42.190 173.650 ;
        RECT 53.845 173.790 54.135 173.835 ;
        RECT 60.270 173.790 60.590 173.850 ;
        RECT 53.845 173.650 60.590 173.790 ;
        RECT 53.845 173.605 54.135 173.650 ;
        RECT 60.270 173.590 60.590 173.650 ;
        RECT 65.330 173.790 65.650 173.850 ;
        RECT 71.400 173.790 71.540 174.285 ;
        RECT 75.910 174.270 76.230 174.330 ;
        RECT 77.290 174.270 77.610 174.330 ;
        RECT 79.130 174.270 79.450 174.330 ;
        RECT 82.825 174.470 83.115 174.515 ;
        RECT 85.110 174.470 85.430 174.530 ;
        RECT 82.825 174.330 85.430 174.470 ;
        RECT 82.825 174.285 83.115 174.330 ;
        RECT 85.110 174.270 85.430 174.330 ;
        RECT 89.220 174.470 89.510 174.515 ;
        RECT 89.220 174.330 91.755 174.470 ;
        RECT 89.220 174.285 89.510 174.330 ;
        RECT 76.370 174.130 76.690 174.190 ;
        RECT 80.985 174.130 81.275 174.175 ;
        RECT 76.370 173.990 81.275 174.130 ;
        RECT 76.370 173.930 76.690 173.990 ;
        RECT 80.985 173.945 81.275 173.990 ;
        RECT 83.730 174.130 84.050 174.190 ;
        RECT 91.540 174.175 91.755 174.330 ;
        RECT 94.325 174.285 94.615 174.515 ;
        RECT 87.360 174.130 87.650 174.175 ;
        RECT 90.620 174.130 90.910 174.175 ;
        RECT 83.730 173.990 90.910 174.130 ;
        RECT 83.730 173.930 84.050 173.990 ;
        RECT 87.360 173.945 87.650 173.990 ;
        RECT 90.620 173.945 90.910 173.990 ;
        RECT 91.540 174.130 91.830 174.175 ;
        RECT 93.400 174.130 93.690 174.175 ;
        RECT 91.540 173.990 93.690 174.130 ;
        RECT 94.400 174.130 94.540 174.285 ;
        RECT 95.690 174.270 96.010 174.530 ;
        RECT 96.240 174.470 96.380 174.670 ;
        RECT 97.990 174.610 98.310 174.870 ;
        RECT 98.465 174.810 98.755 174.855 ;
        RECT 101.210 174.810 101.530 174.870 ;
        RECT 98.465 174.670 101.530 174.810 ;
        RECT 98.465 174.625 98.755 174.670 ;
        RECT 101.210 174.610 101.530 174.670 ;
        RECT 105.810 174.810 106.130 174.870 ;
        RECT 106.285 174.810 106.575 174.855 ;
        RECT 105.810 174.670 106.575 174.810 ;
        RECT 105.810 174.610 106.130 174.670 ;
        RECT 106.285 174.625 106.575 174.670 ;
        RECT 111.330 174.810 111.650 174.870 ;
        RECT 116.405 174.810 116.695 174.855 ;
        RECT 111.330 174.670 116.695 174.810 ;
        RECT 111.330 174.610 111.650 174.670 ;
        RECT 116.405 174.625 116.695 174.670 ;
        RECT 117.310 174.610 117.630 174.870 ;
        RECT 122.920 174.855 123.060 175.010 ;
        RECT 122.845 174.625 123.135 174.855 ;
        RECT 123.750 174.610 124.070 174.870 ;
        RECT 135.635 174.550 136.775 223.880 ;
        RECT 138.130 223.810 139.580 225.110 ;
        RECT 143.180 223.840 144.630 225.140 ;
        RECT 98.925 174.470 99.215 174.515 ;
        RECT 96.240 174.330 99.215 174.470 ;
        RECT 98.925 174.285 99.215 174.330 ;
        RECT 104.905 174.470 105.195 174.515 ;
        RECT 105.350 174.470 105.670 174.530 ;
        RECT 115.010 174.515 115.330 174.530 ;
        RECT 104.905 174.330 105.670 174.470 ;
        RECT 104.905 174.285 105.195 174.330 ;
        RECT 105.350 174.270 105.670 174.330 ;
        RECT 99.370 174.130 99.690 174.190 ;
        RECT 104.430 174.130 104.750 174.190 ;
        RECT 94.400 173.990 99.690 174.130 ;
        RECT 91.540 173.945 91.830 173.990 ;
        RECT 93.400 173.945 93.690 173.990 ;
        RECT 99.370 173.930 99.690 173.990 ;
        RECT 99.920 173.990 104.750 174.130 ;
        RECT 65.330 173.650 71.540 173.790 ;
        RECT 65.330 173.590 65.650 173.650 ;
        RECT 72.230 173.590 72.550 173.850 ;
        RECT 85.355 173.790 85.645 173.835 ;
        RECT 86.490 173.790 86.810 173.850 ;
        RECT 85.355 173.650 86.810 173.790 ;
        RECT 85.355 173.605 85.645 173.650 ;
        RECT 86.490 173.590 86.810 173.650 ;
        RECT 90.170 173.790 90.490 173.850 ;
        RECT 99.920 173.790 100.060 173.990 ;
        RECT 104.430 173.930 104.750 173.990 ;
        RECT 106.270 174.130 106.590 174.190 ;
        RECT 108.065 174.175 108.355 174.490 ;
        RECT 109.145 174.470 109.435 174.515 ;
        RECT 112.725 174.470 113.015 174.515 ;
        RECT 114.560 174.470 114.850 174.515 ;
        RECT 109.145 174.330 114.850 174.470 ;
        RECT 109.145 174.285 109.435 174.330 ;
        RECT 112.725 174.285 113.015 174.330 ;
        RECT 114.560 174.285 114.850 174.330 ;
        RECT 114.990 174.470 115.330 174.515 ;
        RECT 117.770 174.470 118.090 174.530 ;
        RECT 120.085 174.470 120.375 174.515 ;
        RECT 114.990 174.330 117.540 174.470 ;
        RECT 114.990 174.285 115.330 174.330 ;
        RECT 115.010 174.270 115.330 174.285 ;
        RECT 107.765 174.130 108.355 174.175 ;
        RECT 111.005 174.130 111.655 174.175 ;
        RECT 106.270 173.990 111.655 174.130 ;
        RECT 106.270 173.930 106.590 173.990 ;
        RECT 107.765 173.945 108.055 173.990 ;
        RECT 111.005 173.945 111.655 173.990 ;
        RECT 112.250 174.130 112.570 174.190 ;
        RECT 113.645 174.130 113.935 174.175 ;
        RECT 112.250 173.990 113.935 174.130 ;
        RECT 117.400 174.130 117.540 174.330 ;
        RECT 117.770 174.330 120.375 174.470 ;
        RECT 117.770 174.270 118.090 174.330 ;
        RECT 120.085 174.285 120.375 174.330 ;
        RECT 124.685 174.470 124.975 174.515 ;
        RECT 130.650 174.470 130.970 174.530 ;
        RECT 124.685 174.330 130.970 174.470 ;
        RECT 124.685 174.285 124.975 174.330 ;
        RECT 130.650 174.270 130.970 174.330 ;
        RECT 126.050 174.130 126.370 174.190 ;
        RECT 117.400 173.990 126.370 174.130 ;
        RECT 112.250 173.930 112.570 173.990 ;
        RECT 113.645 173.945 113.935 173.990 ;
        RECT 126.050 173.930 126.370 173.990 ;
        RECT 90.170 173.650 100.060 173.790 ;
        RECT 119.625 173.790 119.915 173.835 ;
        RECT 122.830 173.790 123.150 173.850 ;
        RECT 119.625 173.650 123.150 173.790 ;
        RECT 90.170 173.590 90.490 173.650 ;
        RECT 119.625 173.605 119.915 173.650 ;
        RECT 122.830 173.590 123.150 173.650 ;
        RECT 29.840 172.970 127.820 173.450 ;
        RECT 135.580 173.430 136.830 174.550 ;
        RECT 135.635 173.420 136.775 173.430 ;
        RECT 35.445 172.770 35.735 172.815 ;
        RECT 35.890 172.770 36.210 172.830 ;
        RECT 35.445 172.630 36.210 172.770 ;
        RECT 35.445 172.585 35.735 172.630 ;
        RECT 35.890 172.570 36.210 172.630 ;
        RECT 38.650 172.570 38.970 172.830 ;
        RECT 39.110 172.770 39.430 172.830 ;
        RECT 40.045 172.770 40.335 172.815 ;
        RECT 39.110 172.630 40.335 172.770 ;
        RECT 39.110 172.570 39.430 172.630 ;
        RECT 40.045 172.585 40.335 172.630 ;
        RECT 41.425 172.585 41.715 172.815 ;
        RECT 56.145 172.770 56.435 172.815 ;
        RECT 57.510 172.770 57.830 172.830 ;
        RECT 56.145 172.630 57.830 172.770 ;
        RECT 56.145 172.585 56.435 172.630 ;
        RECT 35.430 172.090 35.750 172.150 ;
        RECT 35.905 172.090 36.195 172.135 ;
        RECT 35.430 171.950 36.195 172.090 ;
        RECT 35.430 171.890 35.750 171.950 ;
        RECT 35.905 171.905 36.195 171.950 ;
        RECT 39.585 172.090 39.875 172.135 ;
        RECT 40.490 172.090 40.810 172.150 ;
        RECT 39.585 171.950 40.810 172.090 ;
        RECT 39.585 171.905 39.875 171.950 ;
        RECT 40.490 171.890 40.810 171.950 ;
        RECT 40.965 172.090 41.255 172.135 ;
        RECT 41.500 172.090 41.640 172.585 ;
        RECT 57.510 172.570 57.830 172.630 ;
        RECT 57.970 172.770 58.290 172.830 ;
        RECT 62.570 172.770 62.890 172.830 ;
        RECT 68.090 172.770 68.410 172.830 ;
        RECT 57.970 172.630 62.890 172.770 ;
        RECT 57.970 172.570 58.290 172.630 ;
        RECT 62.570 172.570 62.890 172.630 ;
        RECT 63.120 172.630 68.410 172.770 ;
        RECT 41.870 172.430 42.190 172.490 ;
        RECT 43.725 172.430 44.015 172.475 ;
        RECT 51.545 172.430 51.835 172.475 ;
        RECT 41.870 172.290 51.835 172.430 ;
        RECT 41.870 172.230 42.190 172.290 ;
        RECT 43.725 172.245 44.015 172.290 ;
        RECT 51.545 172.245 51.835 172.290 ;
        RECT 52.005 172.430 52.295 172.475 ;
        RECT 63.120 172.430 63.260 172.630 ;
        RECT 68.090 172.570 68.410 172.630 ;
        RECT 83.730 172.570 84.050 172.830 ;
        RECT 86.030 172.570 86.350 172.830 ;
        RECT 88.330 172.570 88.650 172.830 ;
        RECT 97.545 172.770 97.835 172.815 ;
        RECT 99.370 172.770 99.690 172.830 ;
        RECT 102.590 172.770 102.910 172.830 ;
        RECT 105.350 172.770 105.670 172.830 ;
        RECT 117.310 172.770 117.630 172.830 ;
        RECT 117.785 172.770 118.075 172.815 ;
        RECT 97.545 172.630 108.800 172.770 ;
        RECT 97.545 172.585 97.835 172.630 ;
        RECT 99.370 172.570 99.690 172.630 ;
        RECT 102.590 172.570 102.910 172.630 ;
        RECT 105.350 172.570 105.670 172.630 ;
        RECT 52.005 172.290 63.260 172.430 ;
        RECT 63.965 172.430 64.255 172.475 ;
        RECT 66.365 172.430 66.655 172.475 ;
        RECT 69.605 172.430 70.255 172.475 ;
        RECT 63.965 172.290 70.255 172.430 ;
        RECT 52.005 172.245 52.295 172.290 ;
        RECT 63.965 172.245 64.255 172.290 ;
        RECT 66.365 172.245 66.955 172.290 ;
        RECT 69.605 172.245 70.255 172.290 ;
        RECT 43.250 172.090 43.570 172.150 ;
        RECT 40.965 171.950 41.640 172.090 ;
        RECT 41.960 171.950 43.570 172.090 ;
        RECT 40.965 171.905 41.255 171.950 ;
        RECT 40.030 171.750 40.350 171.810 ;
        RECT 41.960 171.750 42.100 171.950 ;
        RECT 43.250 171.890 43.570 171.950 ;
        RECT 46.485 172.090 46.775 172.135 ;
        RECT 60.270 172.090 60.590 172.150 ;
        RECT 46.485 171.950 60.590 172.090 ;
        RECT 46.485 171.905 46.775 171.950 ;
        RECT 60.270 171.890 60.590 171.950 ;
        RECT 61.190 172.090 61.510 172.150 ;
        RECT 62.585 172.090 62.875 172.135 ;
        RECT 61.190 171.950 62.875 172.090 ;
        RECT 61.190 171.890 61.510 171.950 ;
        RECT 62.585 171.905 62.875 171.950 ;
        RECT 40.030 171.610 42.100 171.750 ;
        RECT 44.185 171.750 44.475 171.795 ;
        RECT 52.465 171.750 52.755 171.795 ;
        RECT 57.050 171.750 57.370 171.810 ;
        RECT 44.185 171.610 57.370 171.750 ;
        RECT 62.660 171.750 62.800 171.905 ;
        RECT 63.490 171.890 63.810 172.150 ;
        RECT 66.665 171.930 66.955 172.245 ;
        RECT 72.230 172.230 72.550 172.490 ;
        RECT 76.370 172.430 76.690 172.490 ;
        RECT 76.845 172.430 77.135 172.475 ;
        RECT 76.370 172.290 77.135 172.430 ;
        RECT 76.370 172.230 76.690 172.290 ;
        RECT 76.845 172.245 77.135 172.290 ;
        RECT 90.170 172.230 90.490 172.490 ;
        RECT 101.670 172.475 101.990 172.490 ;
        RECT 101.620 172.430 101.990 172.475 ;
        RECT 104.880 172.430 105.170 172.475 ;
        RECT 101.620 172.290 105.170 172.430 ;
        RECT 101.620 172.245 101.990 172.290 ;
        RECT 104.880 172.245 105.170 172.290 ;
        RECT 105.800 172.430 106.090 172.475 ;
        RECT 107.660 172.430 107.950 172.475 ;
        RECT 105.800 172.290 107.950 172.430 ;
        RECT 105.800 172.245 106.090 172.290 ;
        RECT 107.660 172.245 107.950 172.290 ;
        RECT 108.660 172.430 108.800 172.630 ;
        RECT 117.310 172.630 118.075 172.770 ;
        RECT 117.310 172.570 117.630 172.630 ;
        RECT 117.785 172.585 118.075 172.630 ;
        RECT 123.765 172.770 124.055 172.815 ;
        RECT 124.210 172.770 124.530 172.830 ;
        RECT 123.765 172.630 124.530 172.770 ;
        RECT 123.765 172.585 124.055 172.630 ;
        RECT 124.210 172.570 124.530 172.630 ;
        RECT 115.010 172.430 115.330 172.490 ;
        RECT 108.660 172.290 115.330 172.430 ;
        RECT 101.670 172.230 101.990 172.245 ;
        RECT 67.745 172.090 68.035 172.135 ;
        RECT 71.325 172.090 71.615 172.135 ;
        RECT 73.160 172.090 73.450 172.135 ;
        RECT 67.745 171.950 73.450 172.090 ;
        RECT 67.745 171.905 68.035 171.950 ;
        RECT 71.325 171.905 71.615 171.950 ;
        RECT 73.160 171.905 73.450 171.950 ;
        RECT 79.605 172.090 79.895 172.135 ;
        RECT 80.510 172.090 80.830 172.150 ;
        RECT 79.605 171.950 80.830 172.090 ;
        RECT 79.605 171.905 79.895 171.950 ;
        RECT 80.510 171.890 80.830 171.950 ;
        RECT 84.205 172.090 84.495 172.135 ;
        RECT 86.490 172.090 86.810 172.150 ;
        RECT 87.410 172.090 87.730 172.150 ;
        RECT 84.205 171.950 86.260 172.090 ;
        RECT 84.205 171.905 84.495 171.950 ;
        RECT 63.950 171.750 64.270 171.810 ;
        RECT 73.625 171.750 73.915 171.795 ;
        RECT 75.450 171.750 75.770 171.810 ;
        RECT 62.660 171.610 64.270 171.750 ;
        RECT 40.030 171.550 40.350 171.610 ;
        RECT 44.185 171.565 44.475 171.610 ;
        RECT 52.465 171.565 52.755 171.610 ;
        RECT 42.790 171.410 43.110 171.470 ;
        RECT 44.260 171.410 44.400 171.565 ;
        RECT 57.050 171.550 57.370 171.610 ;
        RECT 63.950 171.550 64.270 171.610 ;
        RECT 64.500 171.610 75.770 171.750 ;
        RECT 42.790 171.270 44.400 171.410 ;
        RECT 57.510 171.410 57.830 171.470 ;
        RECT 64.500 171.410 64.640 171.610 ;
        RECT 73.625 171.565 73.915 171.610 ;
        RECT 75.450 171.550 75.770 171.610 ;
        RECT 85.110 171.550 85.430 171.810 ;
        RECT 86.120 171.750 86.260 171.950 ;
        RECT 86.490 171.950 87.730 172.090 ;
        RECT 86.490 171.890 86.810 171.950 ;
        RECT 87.410 171.890 87.730 171.950 ;
        RECT 103.480 172.090 103.770 172.135 ;
        RECT 105.800 172.090 106.015 172.245 ;
        RECT 108.660 172.135 108.800 172.290 ;
        RECT 115.010 172.230 115.330 172.290 ;
        RECT 115.930 172.430 116.250 172.490 ;
        RECT 115.930 172.290 120.300 172.430 ;
        RECT 115.930 172.230 116.250 172.290 ;
        RECT 103.480 171.950 106.015 172.090 ;
        RECT 103.480 171.905 103.770 171.950 ;
        RECT 108.585 171.905 108.875 172.135 ;
        RECT 109.490 172.090 109.810 172.150 ;
        RECT 120.160 172.135 120.300 172.290 ;
        RECT 109.965 172.090 110.255 172.135 ;
        RECT 109.490 171.950 110.255 172.090 ;
        RECT 109.490 171.890 109.810 171.950 ;
        RECT 109.965 171.905 110.255 171.950 ;
        RECT 120.085 171.905 120.375 172.135 ;
        RECT 121.465 171.905 121.755 172.135 ;
        RECT 95.690 171.750 96.010 171.810 ;
        RECT 86.120 171.610 96.010 171.750 ;
        RECT 95.690 171.550 96.010 171.610 ;
        RECT 106.745 171.750 107.035 171.795 ;
        RECT 106.745 171.610 109.260 171.750 ;
        RECT 106.745 171.565 107.035 171.610 ;
        RECT 109.120 171.455 109.260 171.610 ;
        RECT 113.630 171.550 113.950 171.810 ;
        RECT 116.405 171.565 116.695 171.795 ;
        RECT 57.510 171.270 64.640 171.410 ;
        RECT 67.745 171.410 68.035 171.455 ;
        RECT 70.865 171.410 71.155 171.455 ;
        RECT 72.755 171.410 73.045 171.455 ;
        RECT 67.745 171.270 73.045 171.410 ;
        RECT 42.790 171.210 43.110 171.270 ;
        RECT 57.510 171.210 57.830 171.270 ;
        RECT 67.745 171.225 68.035 171.270 ;
        RECT 70.865 171.225 71.155 171.270 ;
        RECT 72.755 171.225 73.045 171.270 ;
        RECT 103.480 171.410 103.770 171.455 ;
        RECT 106.260 171.410 106.550 171.455 ;
        RECT 108.120 171.410 108.410 171.455 ;
        RECT 103.480 171.270 108.410 171.410 ;
        RECT 103.480 171.225 103.770 171.270 ;
        RECT 106.260 171.225 106.550 171.270 ;
        RECT 108.120 171.225 108.410 171.270 ;
        RECT 109.045 171.225 109.335 171.455 ;
        RECT 111.330 171.410 111.650 171.470 ;
        RECT 116.480 171.410 116.620 171.565 ;
        RECT 117.310 171.550 117.630 171.810 ;
        RECT 121.540 171.750 121.680 171.905 ;
        RECT 122.830 171.890 123.150 172.150 ;
        RECT 133.500 172.050 136.690 172.190 ;
        RECT 129.260 171.930 136.690 172.050 ;
        RECT 138.330 171.930 139.470 223.810 ;
        RECT 119.700 171.610 121.680 171.750 ;
        RECT 119.700 171.455 119.840 171.610 ;
        RECT 111.330 171.270 116.620 171.410 ;
        RECT 111.330 171.210 111.650 171.270 ;
        RECT 119.625 171.225 119.915 171.455 ;
        RECT 49.230 170.870 49.550 171.130 ;
        RECT 49.690 170.870 50.010 171.130 ;
        RECT 60.730 171.070 61.050 171.130 ;
        RECT 64.870 171.070 65.190 171.130 ;
        RECT 60.730 170.930 65.190 171.070 ;
        RECT 60.730 170.870 61.050 170.930 ;
        RECT 64.870 170.870 65.190 170.930 ;
        RECT 69.930 171.070 70.250 171.130 ;
        RECT 75.465 171.070 75.755 171.115 ;
        RECT 69.930 170.930 75.755 171.070 ;
        RECT 69.930 170.870 70.250 170.930 ;
        RECT 75.465 170.885 75.755 170.930 ;
        RECT 76.370 171.070 76.690 171.130 ;
        RECT 78.685 171.070 78.975 171.115 ;
        RECT 76.370 170.930 78.975 171.070 ;
        RECT 76.370 170.870 76.690 170.930 ;
        RECT 78.685 170.885 78.975 170.930 ;
        RECT 98.910 171.070 99.230 171.130 ;
        RECT 99.615 171.070 99.905 171.115 ;
        RECT 98.910 170.930 99.905 171.070 ;
        RECT 98.910 170.870 99.230 170.930 ;
        RECT 99.615 170.885 99.905 170.930 ;
        RECT 110.410 170.870 110.730 171.130 ;
        RECT 120.530 170.870 120.850 171.130 ;
        RECT 122.385 171.070 122.675 171.115 ;
        RECT 124.210 171.070 124.530 171.130 ;
        RECT 122.385 170.930 124.530 171.070 ;
        RECT 122.385 170.885 122.675 170.930 ;
        RECT 124.210 170.870 124.530 170.930 ;
        RECT 129.260 170.790 139.470 171.930 ;
        RECT 29.840 170.250 127.820 170.730 ;
        RECT 133.500 170.600 136.690 170.790 ;
        RECT 40.490 170.050 40.810 170.110 ;
        RECT 40.965 170.050 41.255 170.095 ;
        RECT 40.490 169.910 41.255 170.050 ;
        RECT 40.490 169.850 40.810 169.910 ;
        RECT 40.965 169.865 41.255 169.910 ;
        RECT 51.990 169.850 52.310 170.110 ;
        RECT 59.365 170.050 59.655 170.095 ;
        RECT 65.330 170.050 65.650 170.110 ;
        RECT 59.365 169.910 65.650 170.050 ;
        RECT 59.365 169.865 59.655 169.910 ;
        RECT 65.330 169.850 65.650 169.910 ;
        RECT 91.090 170.050 91.410 170.110 ;
        RECT 91.565 170.050 91.855 170.095 ;
        RECT 91.090 169.910 91.855 170.050 ;
        RECT 91.090 169.850 91.410 169.910 ;
        RECT 91.565 169.865 91.855 169.910 ;
        RECT 107.205 170.050 107.495 170.095 ;
        RECT 109.490 170.050 109.810 170.110 ;
        RECT 107.205 169.910 109.810 170.050 ;
        RECT 107.205 169.865 107.495 169.910 ;
        RECT 109.490 169.850 109.810 169.910 ;
        RECT 109.965 170.050 110.255 170.095 ;
        RECT 112.250 170.050 112.570 170.110 ;
        RECT 109.965 169.910 112.570 170.050 ;
        RECT 109.965 169.865 110.255 169.910 ;
        RECT 112.250 169.850 112.570 169.910 ;
        RECT 113.630 170.050 113.950 170.110 ;
        RECT 114.105 170.050 114.395 170.095 ;
        RECT 113.630 169.910 114.395 170.050 ;
        RECT 113.630 169.850 113.950 169.910 ;
        RECT 114.105 169.865 114.395 169.910 ;
        RECT 35.400 169.710 35.690 169.755 ;
        RECT 38.180 169.710 38.470 169.755 ;
        RECT 40.040 169.710 40.330 169.755 ;
        RECT 60.730 169.710 61.050 169.770 ;
        RECT 35.400 169.570 40.330 169.710 ;
        RECT 35.400 169.525 35.690 169.570 ;
        RECT 38.180 169.525 38.470 169.570 ;
        RECT 40.040 169.525 40.330 169.570 ;
        RECT 53.690 169.570 61.050 169.710 ;
        RECT 39.570 169.370 39.890 169.430 ;
        RECT 40.505 169.370 40.795 169.415 ;
        RECT 39.570 169.230 40.795 169.370 ;
        RECT 39.570 169.170 39.890 169.230 ;
        RECT 40.505 169.185 40.795 169.230 ;
        RECT 43.250 169.170 43.570 169.430 ;
        RECT 43.725 169.185 44.015 169.415 ;
        RECT 53.690 169.370 53.830 169.570 ;
        RECT 60.730 169.510 61.050 169.570 ;
        RECT 69.585 169.710 69.875 169.755 ;
        RECT 72.705 169.710 72.995 169.755 ;
        RECT 74.595 169.710 74.885 169.755 ;
        RECT 69.585 169.570 74.885 169.710 ;
        RECT 69.585 169.525 69.875 169.570 ;
        RECT 72.705 169.525 72.995 169.570 ;
        RECT 74.595 169.525 74.885 169.570 ;
        RECT 85.110 169.710 85.430 169.770 ;
        RECT 104.890 169.710 105.210 169.770 ;
        RECT 105.810 169.710 106.130 169.770 ;
        RECT 119.725 169.710 120.015 169.755 ;
        RECT 122.845 169.710 123.135 169.755 ;
        RECT 124.735 169.710 125.025 169.755 ;
        RECT 85.110 169.570 87.180 169.710 ;
        RECT 85.110 169.510 85.430 169.570 ;
        RECT 87.040 169.430 87.180 169.570 ;
        RECT 93.940 169.570 112.020 169.710 ;
        RECT 46.560 169.230 52.450 169.370 ;
        RECT 35.400 169.030 35.690 169.075 ;
        RECT 35.400 168.890 37.935 169.030 ;
        RECT 35.400 168.845 35.690 168.890 ;
        RECT 33.540 168.690 33.830 168.735 ;
        RECT 34.970 168.690 35.290 168.750 ;
        RECT 37.720 168.735 37.935 168.890 ;
        RECT 38.650 168.830 38.970 169.090 ;
        RECT 39.110 169.030 39.430 169.090 ;
        RECT 42.790 169.030 43.110 169.090 ;
        RECT 43.800 169.030 43.940 169.185 ;
        RECT 46.560 169.075 46.700 169.230 ;
        RECT 39.110 168.890 43.940 169.030 ;
        RECT 39.110 168.830 39.430 168.890 ;
        RECT 42.790 168.830 43.110 168.890 ;
        RECT 46.485 168.845 46.775 169.075 ;
        RECT 47.405 168.845 47.695 169.075 ;
        RECT 36.800 168.690 37.090 168.735 ;
        RECT 33.540 168.550 37.090 168.690 ;
        RECT 33.540 168.505 33.830 168.550 ;
        RECT 34.970 168.490 35.290 168.550 ;
        RECT 36.800 168.505 37.090 168.550 ;
        RECT 37.720 168.690 38.010 168.735 ;
        RECT 39.580 168.690 39.870 168.735 ;
        RECT 37.720 168.550 39.870 168.690 ;
        RECT 37.720 168.505 38.010 168.550 ;
        RECT 39.580 168.505 39.870 168.550 ;
        RECT 45.090 168.690 45.410 168.750 ;
        RECT 47.480 168.690 47.620 168.845 ;
        RECT 47.850 168.830 48.170 169.090 ;
        RECT 48.325 168.845 48.615 169.075 ;
        RECT 49.690 169.030 50.010 169.090 ;
        RECT 52.310 169.075 52.450 169.230 ;
        RECT 53.460 169.230 53.830 169.370 ;
        RECT 56.605 169.370 56.895 169.415 ;
        RECT 57.970 169.370 58.290 169.430 ;
        RECT 56.605 169.230 58.290 169.370 ;
        RECT 51.085 169.030 51.375 169.075 ;
        RECT 49.690 168.890 51.375 169.030 ;
        RECT 52.310 169.030 52.695 169.075 ;
        RECT 52.910 169.030 53.230 169.090 ;
        RECT 53.460 169.075 53.600 169.230 ;
        RECT 56.605 169.185 56.895 169.230 ;
        RECT 57.970 169.170 58.290 169.230 ;
        RECT 75.450 169.170 75.770 169.430 ;
        RECT 86.030 169.370 86.350 169.430 ;
        RECT 84.740 169.230 86.350 169.370 ;
        RECT 52.310 168.890 53.230 169.030 ;
        RECT 45.090 168.550 47.620 168.690 ;
        RECT 48.400 168.690 48.540 168.845 ;
        RECT 49.690 168.830 50.010 168.890 ;
        RECT 51.085 168.845 51.375 168.890 ;
        RECT 52.405 168.845 52.695 168.890 ;
        RECT 52.910 168.830 53.230 168.890 ;
        RECT 53.385 168.845 53.675 169.075 ;
        RECT 53.830 168.830 54.150 169.090 ;
        RECT 54.305 168.845 54.595 169.075 ;
        RECT 57.510 169.030 57.830 169.090 ;
        RECT 59.810 169.030 60.130 169.090 ;
        RECT 60.285 169.030 60.575 169.075 ;
        RECT 57.510 168.890 60.575 169.030 ;
        RECT 54.380 168.690 54.520 168.845 ;
        RECT 57.510 168.830 57.830 168.890 ;
        RECT 59.810 168.830 60.130 168.890 ;
        RECT 60.285 168.845 60.575 168.890 ;
        RECT 68.505 168.735 68.795 169.050 ;
        RECT 69.585 169.030 69.875 169.075 ;
        RECT 73.165 169.030 73.455 169.075 ;
        RECT 75.000 169.030 75.290 169.075 ;
        RECT 69.585 168.890 75.290 169.030 ;
        RECT 69.585 168.845 69.875 168.890 ;
        RECT 73.165 168.845 73.455 168.890 ;
        RECT 75.000 168.845 75.290 168.890 ;
        RECT 78.685 169.030 78.975 169.075 ;
        RECT 79.590 169.030 79.910 169.090 ;
        RECT 78.685 168.890 79.910 169.030 ;
        RECT 78.685 168.845 78.975 168.890 ;
        RECT 79.590 168.830 79.910 168.890 ;
        RECT 80.510 168.830 80.830 169.090 ;
        RECT 82.350 169.030 82.670 169.090 ;
        RECT 83.745 169.030 84.035 169.075 ;
        RECT 82.350 168.890 84.035 169.030 ;
        RECT 82.350 168.830 82.670 168.890 ;
        RECT 83.745 168.845 84.035 168.890 ;
        RECT 84.190 168.830 84.510 169.090 ;
        RECT 84.740 169.075 84.880 169.230 ;
        RECT 86.030 169.170 86.350 169.230 ;
        RECT 86.950 169.370 87.270 169.430 ;
        RECT 93.940 169.415 94.080 169.570 ;
        RECT 104.890 169.510 105.210 169.570 ;
        RECT 105.810 169.510 106.130 169.570 ;
        RECT 86.950 169.230 93.620 169.370 ;
        RECT 86.950 169.170 87.270 169.230 ;
        RECT 84.665 168.845 84.955 169.075 ;
        RECT 85.585 169.030 85.875 169.075 ;
        RECT 86.490 169.030 86.810 169.090 ;
        RECT 90.645 169.030 90.935 169.075 ;
        RECT 85.585 168.890 86.810 169.030 ;
        RECT 85.585 168.845 85.875 168.890 ;
        RECT 86.490 168.830 86.810 168.890 ;
        RECT 89.800 168.890 90.935 169.030 ;
        RECT 93.480 169.030 93.620 169.230 ;
        RECT 93.865 169.185 94.155 169.415 ;
        RECT 97.545 169.370 97.835 169.415 ;
        RECT 97.990 169.370 98.310 169.430 ;
        RECT 103.985 169.370 104.275 169.415 ;
        RECT 110.885 169.370 111.175 169.415 ;
        RECT 111.330 169.370 111.650 169.430 ;
        RECT 111.880 169.415 112.020 169.570 ;
        RECT 119.725 169.570 125.025 169.710 ;
        RECT 119.725 169.525 120.015 169.570 ;
        RECT 122.845 169.525 123.135 169.570 ;
        RECT 124.735 169.525 125.025 169.570 ;
        RECT 97.545 169.230 111.650 169.370 ;
        RECT 97.545 169.185 97.835 169.230 ;
        RECT 97.620 169.030 97.760 169.185 ;
        RECT 97.990 169.170 98.310 169.230 ;
        RECT 103.985 169.185 104.275 169.230 ;
        RECT 110.885 169.185 111.175 169.230 ;
        RECT 111.330 169.170 111.650 169.230 ;
        RECT 111.805 169.185 112.095 169.415 ;
        RECT 124.210 169.170 124.530 169.430 ;
        RECT 93.480 168.890 97.760 169.030 ;
        RECT 98.910 169.030 99.230 169.090 ;
        RECT 104.905 169.030 105.195 169.075 ;
        RECT 98.910 168.890 105.195 169.030 ;
        RECT 48.400 168.550 54.520 168.690 ;
        RECT 68.205 168.690 68.795 168.735 ;
        RECT 70.390 168.690 70.710 168.750 ;
        RECT 71.445 168.690 72.095 168.735 ;
        RECT 68.205 168.550 72.095 168.690 ;
        RECT 45.090 168.490 45.410 168.550 ;
        RECT 53.920 168.410 54.060 168.550 ;
        RECT 68.205 168.505 68.495 168.550 ;
        RECT 70.390 168.490 70.710 168.550 ;
        RECT 71.445 168.505 72.095 168.550 ;
        RECT 73.610 168.690 73.930 168.750 ;
        RECT 74.085 168.690 74.375 168.735 ;
        RECT 73.610 168.550 74.375 168.690 ;
        RECT 73.610 168.490 73.930 168.550 ;
        RECT 74.085 168.505 74.375 168.550 ;
        RECT 87.410 168.490 87.730 168.750 ;
        RECT 31.535 168.350 31.825 168.395 ;
        RECT 37.270 168.350 37.590 168.410 ;
        RECT 42.790 168.350 43.110 168.410 ;
        RECT 31.535 168.210 43.110 168.350 ;
        RECT 31.535 168.165 31.825 168.210 ;
        RECT 37.270 168.150 37.590 168.210 ;
        RECT 42.790 168.150 43.110 168.210 ;
        RECT 43.710 168.350 44.030 168.410 ;
        RECT 49.705 168.350 49.995 168.395 ;
        RECT 43.710 168.210 49.995 168.350 ;
        RECT 43.710 168.150 44.030 168.210 ;
        RECT 49.705 168.165 49.995 168.210 ;
        RECT 53.830 168.150 54.150 168.410 ;
        RECT 55.670 168.150 55.990 168.410 ;
        RECT 66.710 168.150 67.030 168.410 ;
        RECT 69.010 168.350 69.330 168.410 ;
        RECT 77.765 168.350 78.055 168.395 ;
        RECT 79.130 168.350 79.450 168.410 ;
        RECT 69.010 168.210 79.450 168.350 ;
        RECT 69.010 168.150 69.330 168.210 ;
        RECT 77.765 168.165 78.055 168.210 ;
        RECT 79.130 168.150 79.450 168.210 ;
        RECT 79.605 168.350 79.895 168.395 ;
        RECT 80.050 168.350 80.370 168.410 ;
        RECT 79.605 168.210 80.370 168.350 ;
        RECT 79.605 168.165 79.895 168.210 ;
        RECT 80.050 168.150 80.370 168.210 ;
        RECT 82.365 168.350 82.655 168.395 ;
        RECT 83.730 168.350 84.050 168.410 ;
        RECT 82.365 168.210 84.050 168.350 ;
        RECT 82.365 168.165 82.655 168.210 ;
        RECT 83.730 168.150 84.050 168.210 ;
        RECT 86.030 168.350 86.350 168.410 ;
        RECT 89.800 168.395 89.940 168.890 ;
        RECT 90.645 168.845 90.935 168.890 ;
        RECT 98.910 168.830 99.230 168.890 ;
        RECT 104.905 168.845 105.195 168.890 ;
        RECT 109.045 169.030 109.335 169.075 ;
        RECT 110.410 169.030 110.730 169.090 ;
        RECT 109.045 168.890 110.730 169.030 ;
        RECT 109.045 168.845 109.335 168.890 ;
        RECT 110.410 168.830 110.730 168.890 ;
        RECT 112.265 169.030 112.555 169.075 ;
        RECT 117.310 169.030 117.630 169.090 ;
        RECT 112.265 168.890 117.630 169.030 ;
        RECT 112.265 168.845 112.555 168.890 ;
        RECT 117.310 168.830 117.630 168.890 ;
        RECT 118.645 168.735 118.935 169.050 ;
        RECT 119.725 169.030 120.015 169.075 ;
        RECT 123.305 169.030 123.595 169.075 ;
        RECT 125.140 169.030 125.430 169.075 ;
        RECT 119.725 168.890 125.430 169.030 ;
        RECT 119.725 168.845 120.015 168.890 ;
        RECT 123.305 168.845 123.595 168.890 ;
        RECT 125.140 168.845 125.430 168.890 ;
        RECT 125.605 169.030 125.895 169.075 ;
        RECT 126.050 169.030 126.370 169.090 ;
        RECT 125.605 168.890 126.370 169.030 ;
        RECT 125.605 168.845 125.895 168.890 ;
        RECT 126.050 168.830 126.370 168.890 ;
        RECT 96.625 168.690 96.915 168.735 ;
        RECT 105.365 168.690 105.655 168.735 ;
        RECT 96.625 168.550 105.655 168.690 ;
        RECT 96.625 168.505 96.915 168.550 ;
        RECT 105.365 168.505 105.655 168.550 ;
        RECT 118.345 168.690 118.935 168.735 ;
        RECT 120.530 168.690 120.850 168.750 ;
        RECT 121.585 168.690 122.235 168.735 ;
        RECT 118.345 168.550 122.235 168.690 ;
        RECT 118.345 168.505 118.635 168.550 ;
        RECT 120.530 168.490 120.850 168.550 ;
        RECT 121.585 168.505 122.235 168.550 ;
        RECT 87.885 168.350 88.175 168.395 ;
        RECT 86.030 168.210 88.175 168.350 ;
        RECT 86.030 168.150 86.350 168.210 ;
        RECT 87.885 168.165 88.175 168.210 ;
        RECT 89.725 168.165 90.015 168.395 ;
        RECT 96.150 168.350 96.470 168.410 ;
        RECT 98.465 168.350 98.755 168.395 ;
        RECT 96.150 168.210 98.755 168.350 ;
        RECT 96.150 168.150 96.470 168.210 ;
        RECT 98.465 168.165 98.755 168.210 ;
        RECT 98.910 168.150 99.230 168.410 ;
        RECT 100.765 168.350 101.055 168.395 ;
        RECT 103.970 168.350 104.290 168.410 ;
        RECT 100.765 168.210 104.290 168.350 ;
        RECT 100.765 168.165 101.055 168.210 ;
        RECT 103.970 168.150 104.290 168.210 ;
        RECT 115.470 168.350 115.790 168.410 ;
        RECT 116.865 168.350 117.155 168.395 ;
        RECT 115.470 168.210 117.155 168.350 ;
        RECT 115.470 168.150 115.790 168.210 ;
        RECT 116.865 168.165 117.155 168.210 ;
        RECT 29.840 167.530 127.820 168.010 ;
        RECT 34.970 167.130 35.290 167.390 ;
        RECT 38.650 167.130 38.970 167.390 ;
        RECT 51.070 167.130 51.390 167.390 ;
        RECT 64.870 167.330 65.190 167.390 ;
        RECT 67.645 167.330 67.935 167.375 ;
        RECT 64.870 167.190 67.935 167.330 ;
        RECT 64.870 167.130 65.190 167.190 ;
        RECT 67.645 167.145 67.935 167.190 ;
        RECT 86.030 167.130 86.350 167.390 ;
        RECT 88.345 167.330 88.635 167.375 ;
        RECT 109.950 167.330 110.270 167.390 ;
        RECT 113.170 167.330 113.490 167.390 ;
        RECT 88.345 167.190 91.780 167.330 ;
        RECT 88.345 167.145 88.635 167.190 ;
        RECT 39.110 166.990 39.430 167.050 ;
        RECT 49.230 166.990 49.550 167.050 ;
        RECT 57.525 166.990 57.815 167.035 ;
        RECT 39.110 166.850 47.160 166.990 ;
        RECT 39.110 166.790 39.430 166.850 ;
        RECT 35.430 166.450 35.750 166.710 ;
        RECT 37.730 166.450 38.050 166.710 ;
        RECT 42.805 166.465 43.095 166.695 ;
        RECT 43.250 166.650 43.570 166.710 ;
        RECT 43.725 166.650 44.015 166.695 ;
        RECT 43.250 166.510 44.015 166.650 ;
        RECT 42.880 166.310 43.020 166.465 ;
        RECT 43.250 166.450 43.570 166.510 ;
        RECT 43.725 166.465 44.015 166.510 ;
        RECT 44.170 166.450 44.490 166.710 ;
        RECT 44.645 166.650 44.935 166.695 ;
        RECT 45.090 166.650 45.410 166.710 ;
        RECT 44.645 166.510 45.410 166.650 ;
        RECT 44.645 166.465 44.935 166.510 ;
        RECT 45.090 166.450 45.410 166.510 ;
        RECT 46.470 166.310 46.790 166.370 ;
        RECT 47.020 166.355 47.160 166.850 ;
        RECT 49.230 166.850 57.815 166.990 ;
        RECT 49.230 166.790 49.550 166.850 ;
        RECT 57.525 166.805 57.815 166.850 ;
        RECT 68.090 166.990 68.410 167.050 ;
        RECT 71.325 166.990 71.615 167.035 ;
        RECT 68.090 166.850 71.615 166.990 ;
        RECT 68.090 166.790 68.410 166.850 ;
        RECT 71.325 166.805 71.615 166.850 ;
        RECT 79.130 166.990 79.450 167.050 ;
        RECT 87.410 166.990 87.730 167.050 ;
        RECT 79.130 166.850 82.580 166.990 ;
        RECT 79.130 166.790 79.450 166.850 ;
        RECT 82.440 166.710 82.580 166.850 ;
        RECT 83.360 166.850 87.730 166.990 ;
        RECT 48.310 166.450 48.630 166.710 ;
        RECT 50.610 166.450 50.930 166.710 ;
        RECT 51.990 166.450 52.310 166.710 ;
        RECT 52.925 166.650 53.215 166.695 ;
        RECT 52.540 166.510 53.215 166.650 ;
        RECT 42.880 166.170 46.790 166.310 ;
        RECT 46.470 166.110 46.790 166.170 ;
        RECT 46.945 166.125 47.235 166.355 ;
        RECT 47.865 166.310 48.155 166.355 ;
        RECT 49.230 166.310 49.550 166.370 ;
        RECT 47.865 166.170 49.550 166.310 ;
        RECT 47.865 166.125 48.155 166.170 ;
        RECT 49.230 166.110 49.550 166.170 ;
        RECT 42.790 165.970 43.110 166.030 ;
        RECT 52.540 165.970 52.680 166.510 ;
        RECT 52.925 166.465 53.215 166.510 ;
        RECT 53.385 166.465 53.675 166.695 ;
        RECT 53.460 166.310 53.600 166.465 ;
        RECT 53.830 166.450 54.150 166.710 ;
        RECT 57.985 166.650 58.275 166.695 ;
        RECT 56.680 166.510 58.275 166.650 ;
        RECT 54.750 166.310 55.070 166.370 ;
        RECT 53.460 166.170 55.070 166.310 ;
        RECT 54.750 166.110 55.070 166.170 ;
        RECT 42.790 165.830 52.680 165.970 ;
        RECT 56.680 165.970 56.820 166.510 ;
        RECT 57.985 166.465 58.275 166.510 ;
        RECT 67.170 166.650 67.490 166.710 ;
        RECT 70.865 166.650 71.155 166.695 ;
        RECT 67.170 166.510 71.155 166.650 ;
        RECT 67.170 166.450 67.490 166.510 ;
        RECT 70.865 166.465 71.155 166.510 ;
        RECT 75.910 166.650 76.230 166.710 ;
        RECT 76.385 166.650 76.675 166.695 ;
        RECT 75.910 166.510 76.675 166.650 ;
        RECT 75.910 166.450 76.230 166.510 ;
        RECT 76.385 166.465 76.675 166.510 ;
        RECT 78.685 166.650 78.975 166.695 ;
        RECT 79.590 166.650 79.910 166.710 ;
        RECT 78.685 166.510 79.910 166.650 ;
        RECT 78.685 166.465 78.975 166.510 ;
        RECT 79.590 166.450 79.910 166.510 ;
        RECT 82.350 166.450 82.670 166.710 ;
        RECT 83.360 166.695 83.500 166.850 ;
        RECT 87.410 166.790 87.730 166.850 ;
        RECT 82.825 166.465 83.115 166.695 ;
        RECT 83.285 166.465 83.575 166.695 ;
        RECT 84.205 166.465 84.495 166.695 ;
        RECT 85.110 166.650 85.430 166.710 ;
        RECT 91.640 166.695 91.780 167.190 ;
        RECT 108.200 167.190 110.270 167.330 ;
        RECT 95.640 166.990 95.930 167.035 ;
        RECT 97.070 166.990 97.390 167.050 ;
        RECT 98.900 166.990 99.190 167.035 ;
        RECT 95.640 166.850 99.190 166.990 ;
        RECT 95.640 166.805 95.930 166.850 ;
        RECT 97.070 166.790 97.390 166.850 ;
        RECT 98.900 166.805 99.190 166.850 ;
        RECT 99.820 166.990 100.110 167.035 ;
        RECT 101.680 166.990 101.970 167.035 ;
        RECT 99.820 166.850 101.970 166.990 ;
        RECT 99.820 166.805 100.110 166.850 ;
        RECT 101.680 166.805 101.970 166.850 ;
        RECT 86.505 166.650 86.795 166.695 ;
        RECT 85.110 166.510 90.860 166.650 ;
        RECT 57.050 166.310 57.370 166.370 ;
        RECT 58.445 166.310 58.735 166.355 ;
        RECT 68.105 166.310 68.395 166.355 ;
        RECT 69.930 166.310 70.250 166.370 ;
        RECT 57.050 166.170 70.250 166.310 ;
        RECT 57.050 166.110 57.370 166.170 ;
        RECT 58.445 166.125 58.735 166.170 ;
        RECT 68.105 166.125 68.395 166.170 ;
        RECT 69.930 166.110 70.250 166.170 ;
        RECT 72.230 166.310 72.550 166.370 ;
        RECT 75.005 166.310 75.295 166.355 ;
        RECT 72.230 166.170 75.295 166.310 ;
        RECT 72.230 166.110 72.550 166.170 ;
        RECT 75.005 166.125 75.295 166.170 ;
        RECT 76.830 166.310 77.150 166.370 ;
        RECT 82.900 166.310 83.040 166.465 ;
        RECT 76.830 166.170 83.040 166.310 ;
        RECT 76.830 166.110 77.150 166.170 ;
        RECT 57.510 165.970 57.830 166.030 ;
        RECT 56.680 165.830 57.830 165.970 ;
        RECT 42.790 165.770 43.110 165.830 ;
        RECT 57.510 165.770 57.830 165.830 ;
        RECT 57.970 165.970 58.290 166.030 ;
        RECT 65.345 165.970 65.635 166.015 ;
        RECT 77.765 165.970 78.055 166.015 ;
        RECT 81.890 165.970 82.210 166.030 ;
        RECT 57.970 165.830 65.635 165.970 ;
        RECT 57.970 165.770 58.290 165.830 ;
        RECT 65.345 165.785 65.635 165.830 ;
        RECT 65.880 165.830 82.210 165.970 ;
        RECT 45.550 165.630 45.870 165.690 ;
        RECT 46.025 165.630 46.315 165.675 ;
        RECT 45.550 165.490 46.315 165.630 ;
        RECT 45.550 165.430 45.870 165.490 ;
        RECT 46.025 165.445 46.315 165.490 ;
        RECT 50.150 165.430 50.470 165.690 ;
        RECT 54.750 165.630 55.070 165.690 ;
        RECT 55.225 165.630 55.515 165.675 ;
        RECT 54.750 165.490 55.515 165.630 ;
        RECT 54.750 165.430 55.070 165.490 ;
        RECT 55.225 165.445 55.515 165.490 ;
        RECT 55.670 165.430 55.990 165.690 ;
        RECT 56.130 165.630 56.450 165.690 ;
        RECT 65.880 165.630 66.020 165.830 ;
        RECT 77.765 165.785 78.055 165.830 ;
        RECT 81.890 165.770 82.210 165.830 ;
        RECT 56.130 165.490 66.020 165.630 ;
        RECT 72.690 165.630 73.010 165.690 ;
        RECT 73.165 165.630 73.455 165.675 ;
        RECT 72.690 165.490 73.455 165.630 ;
        RECT 56.130 165.430 56.450 165.490 ;
        RECT 72.690 165.430 73.010 165.490 ;
        RECT 73.165 165.445 73.455 165.490 ;
        RECT 80.970 165.430 81.290 165.690 ;
        RECT 82.900 165.630 83.040 166.170 ;
        RECT 84.280 165.970 84.420 166.465 ;
        RECT 85.110 166.450 85.430 166.510 ;
        RECT 86.505 166.465 86.795 166.510 ;
        RECT 85.585 166.310 85.875 166.355 ;
        RECT 86.950 166.310 87.270 166.370 ;
        RECT 85.585 166.170 87.270 166.310 ;
        RECT 85.585 166.125 85.875 166.170 ;
        RECT 86.950 166.110 87.270 166.170 ;
        RECT 86.490 165.970 86.810 166.030 ;
        RECT 84.280 165.830 86.810 165.970 ;
        RECT 90.720 165.970 90.860 166.510 ;
        RECT 91.105 166.465 91.395 166.695 ;
        RECT 91.565 166.465 91.855 166.695 ;
        RECT 97.500 166.650 97.790 166.695 ;
        RECT 99.820 166.650 100.035 166.805 ;
        RECT 97.500 166.510 100.035 166.650 ;
        RECT 97.500 166.465 97.790 166.510 ;
        RECT 91.180 166.310 91.320 166.465 ;
        RECT 102.590 166.450 102.910 166.710 ;
        RECT 103.970 166.450 104.290 166.710 ;
        RECT 107.650 166.450 107.970 166.710 ;
        RECT 108.200 166.695 108.340 167.190 ;
        RECT 109.950 167.130 110.270 167.190 ;
        RECT 111.420 167.190 113.490 167.330 ;
        RECT 108.660 166.850 110.640 166.990 ;
        RECT 108.125 166.465 108.415 166.695 ;
        RECT 95.690 166.310 96.010 166.370 ;
        RECT 96.610 166.310 96.930 166.370 ;
        RECT 91.180 166.170 96.930 166.310 ;
        RECT 95.690 166.110 96.010 166.170 ;
        RECT 96.610 166.110 96.930 166.170 ;
        RECT 100.765 166.310 101.055 166.355 ;
        RECT 100.765 166.170 103.280 166.310 ;
        RECT 100.765 166.125 101.055 166.170 ;
        RECT 93.635 165.970 93.925 166.015 ;
        RECT 96.150 165.970 96.470 166.030 ;
        RECT 103.140 166.015 103.280 166.170 ;
        RECT 90.720 165.830 96.470 165.970 ;
        RECT 86.490 165.770 86.810 165.830 ;
        RECT 93.635 165.785 93.925 165.830 ;
        RECT 96.150 165.770 96.470 165.830 ;
        RECT 97.500 165.970 97.790 166.015 ;
        RECT 100.280 165.970 100.570 166.015 ;
        RECT 102.140 165.970 102.430 166.015 ;
        RECT 97.500 165.830 102.430 165.970 ;
        RECT 97.500 165.785 97.790 165.830 ;
        RECT 100.280 165.785 100.570 165.830 ;
        RECT 102.140 165.785 102.430 165.830 ;
        RECT 103.065 165.785 103.355 166.015 ;
        RECT 108.660 165.970 108.800 166.850 ;
        RECT 109.030 166.450 109.350 166.710 ;
        RECT 110.500 166.310 110.640 166.850 ;
        RECT 110.870 166.450 111.190 166.710 ;
        RECT 111.420 166.695 111.560 167.190 ;
        RECT 113.170 167.130 113.490 167.190 ;
        RECT 117.310 167.330 117.630 167.390 ;
        RECT 118.245 167.330 118.535 167.375 ;
        RECT 117.310 167.190 118.535 167.330 ;
        RECT 117.310 167.130 117.630 167.190 ;
        RECT 118.245 167.145 118.535 167.190 ;
        RECT 111.880 166.850 115.700 166.990 ;
        RECT 111.880 166.695 112.020 166.850 ;
        RECT 115.560 166.710 115.700 166.850 ;
        RECT 111.345 166.465 111.635 166.695 ;
        RECT 111.805 166.465 112.095 166.695 ;
        RECT 112.710 166.650 113.030 166.710 ;
        RECT 114.090 166.650 114.410 166.710 ;
        RECT 112.710 166.510 114.410 166.650 ;
        RECT 112.710 166.450 113.030 166.510 ;
        RECT 114.090 166.450 114.410 166.510 ;
        RECT 115.470 166.450 115.790 166.710 ;
        RECT 121.005 166.650 121.295 166.695 ;
        RECT 123.765 166.650 124.055 166.695 ;
        RECT 124.670 166.650 124.990 166.710 ;
        RECT 121.005 166.510 124.990 166.650 ;
        RECT 121.005 166.465 121.295 166.510 ;
        RECT 123.765 166.465 124.055 166.510 ;
        RECT 124.670 166.450 124.990 166.510 ;
        RECT 115.930 166.310 116.250 166.370 ;
        RECT 119.625 166.310 119.915 166.355 ;
        RECT 110.500 166.170 114.320 166.310 ;
        RECT 113.630 165.970 113.950 166.030 ;
        RECT 103.600 165.830 108.800 165.970 ;
        RECT 109.120 165.830 113.950 165.970 ;
        RECT 114.180 165.970 114.320 166.170 ;
        RECT 115.930 166.170 119.915 166.310 ;
        RECT 115.930 166.110 116.250 166.170 ;
        RECT 119.625 166.125 119.915 166.170 ;
        RECT 122.385 166.125 122.675 166.355 ;
        RECT 122.460 165.970 122.600 166.125 ;
        RECT 114.180 165.830 122.600 165.970 ;
        RECT 84.650 165.630 84.970 165.690 ;
        RECT 82.900 165.490 84.970 165.630 ;
        RECT 84.650 165.430 84.970 165.490 ;
        RECT 90.645 165.630 90.935 165.675 ;
        RECT 91.090 165.630 91.410 165.690 ;
        RECT 90.645 165.490 91.410 165.630 ;
        RECT 90.645 165.445 90.935 165.490 ;
        RECT 91.090 165.430 91.410 165.490 ;
        RECT 92.485 165.630 92.775 165.675 ;
        RECT 92.930 165.630 93.250 165.690 ;
        RECT 92.485 165.490 93.250 165.630 ;
        RECT 92.485 165.445 92.775 165.490 ;
        RECT 92.930 165.430 93.250 165.490 ;
        RECT 94.310 165.630 94.630 165.690 ;
        RECT 103.600 165.630 103.740 165.830 ;
        RECT 94.310 165.490 103.740 165.630 ;
        RECT 105.810 165.630 106.130 165.690 ;
        RECT 109.120 165.675 109.260 165.830 ;
        RECT 113.630 165.770 113.950 165.830 ;
        RECT 106.745 165.630 107.035 165.675 ;
        RECT 105.810 165.490 107.035 165.630 ;
        RECT 94.310 165.430 94.630 165.490 ;
        RECT 105.810 165.430 106.130 165.490 ;
        RECT 106.745 165.445 107.035 165.490 ;
        RECT 109.045 165.445 109.335 165.675 ;
        RECT 109.505 165.630 109.795 165.675 ;
        RECT 111.330 165.630 111.650 165.690 ;
        RECT 109.505 165.490 111.650 165.630 ;
        RECT 109.505 165.445 109.795 165.490 ;
        RECT 111.330 165.430 111.650 165.490 ;
        RECT 135.580 165.470 136.830 166.590 ;
        RECT 29.840 164.810 127.820 165.290 ;
        RECT 35.905 164.610 36.195 164.655 ;
        RECT 37.730 164.610 38.050 164.670 ;
        RECT 35.905 164.470 38.050 164.610 ;
        RECT 35.905 164.425 36.195 164.470 ;
        RECT 37.730 164.410 38.050 164.470 ;
        RECT 48.310 164.610 48.630 164.670 ;
        RECT 50.855 164.610 51.145 164.655 ;
        RECT 57.050 164.610 57.370 164.670 ;
        RECT 48.310 164.470 57.370 164.610 ;
        RECT 48.310 164.410 48.630 164.470 ;
        RECT 50.855 164.425 51.145 164.470 ;
        RECT 57.050 164.410 57.370 164.470 ;
        RECT 63.505 164.610 63.795 164.655 ;
        RECT 67.170 164.610 67.490 164.670 ;
        RECT 63.505 164.470 67.490 164.610 ;
        RECT 63.505 164.425 63.795 164.470 ;
        RECT 67.170 164.410 67.490 164.470 ;
        RECT 73.610 164.410 73.930 164.670 ;
        RECT 75.450 164.610 75.770 164.670 ;
        RECT 79.605 164.610 79.895 164.655 ;
        RECT 81.430 164.610 81.750 164.670 ;
        RECT 75.450 164.470 81.750 164.610 ;
        RECT 75.450 164.410 75.770 164.470 ;
        RECT 79.605 164.425 79.895 164.470 ;
        RECT 81.430 164.410 81.750 164.470 ;
        RECT 81.890 164.610 82.210 164.670 ;
        RECT 81.890 164.470 89.480 164.610 ;
        RECT 81.890 164.410 82.210 164.470 ;
        RECT 37.270 164.270 37.590 164.330 ;
        RECT 33.680 164.130 37.590 164.270 ;
        RECT 33.680 163.975 33.820 164.130 ;
        RECT 37.270 164.070 37.590 164.130 ;
        RECT 44.600 164.270 44.890 164.315 ;
        RECT 47.380 164.270 47.670 164.315 ;
        RECT 49.240 164.270 49.530 164.315 ;
        RECT 44.600 164.130 49.530 164.270 ;
        RECT 44.600 164.085 44.890 164.130 ;
        RECT 47.380 164.085 47.670 164.130 ;
        RECT 49.240 164.085 49.530 164.130 ;
        RECT 54.720 164.270 55.010 164.315 ;
        RECT 57.500 164.270 57.790 164.315 ;
        RECT 59.360 164.270 59.650 164.315 ;
        RECT 54.720 164.130 59.650 164.270 ;
        RECT 54.720 164.085 55.010 164.130 ;
        RECT 57.500 164.085 57.790 164.130 ;
        RECT 59.360 164.085 59.650 164.130 ;
        RECT 65.330 164.270 65.650 164.330 ;
        RECT 69.010 164.270 69.330 164.330 ;
        RECT 65.330 164.130 69.330 164.270 ;
        RECT 65.330 164.070 65.650 164.130 ;
        RECT 69.010 164.070 69.330 164.130 ;
        RECT 83.270 164.070 83.590 164.330 ;
        RECT 84.650 164.270 84.970 164.330 ;
        RECT 83.820 164.130 84.970 164.270 ;
        RECT 33.145 163.745 33.435 163.975 ;
        RECT 33.605 163.745 33.895 163.975 ;
        RECT 36.825 163.930 37.115 163.975 ;
        RECT 39.110 163.930 39.430 163.990 ;
        RECT 36.825 163.790 39.430 163.930 ;
        RECT 36.825 163.745 37.115 163.790 ;
        RECT 33.220 163.590 33.360 163.745 ;
        RECT 36.900 163.590 37.040 163.745 ;
        RECT 39.110 163.730 39.430 163.790 ;
        RECT 39.570 163.930 39.890 163.990 ;
        RECT 47.865 163.930 48.155 163.975 ;
        RECT 50.610 163.930 50.930 163.990 ;
        RECT 39.570 163.790 47.620 163.930 ;
        RECT 39.570 163.730 39.890 163.790 ;
        RECT 33.220 163.450 37.040 163.590 ;
        RECT 44.600 163.590 44.890 163.635 ;
        RECT 47.480 163.590 47.620 163.790 ;
        RECT 47.865 163.790 50.930 163.930 ;
        RECT 47.865 163.745 48.155 163.790 ;
        RECT 50.610 163.730 50.930 163.790 ;
        RECT 53.830 163.930 54.150 163.990 ;
        RECT 53.830 163.790 59.580 163.930 ;
        RECT 53.830 163.730 54.150 163.790 ;
        RECT 49.705 163.590 49.995 163.635 ;
        RECT 44.600 163.450 47.135 163.590 ;
        RECT 47.480 163.450 49.995 163.590 ;
        RECT 44.600 163.405 44.890 163.450 ;
        RECT 42.790 163.295 43.110 163.310 ;
        RECT 46.920 163.295 47.135 163.450 ;
        RECT 49.705 163.405 49.995 163.450 ;
        RECT 54.720 163.590 55.010 163.635 ;
        RECT 54.720 163.450 57.255 163.590 ;
        RECT 54.720 163.405 55.010 163.450 ;
        RECT 38.205 163.250 38.495 163.295 ;
        RECT 42.740 163.250 43.110 163.295 ;
        RECT 46.000 163.250 46.290 163.295 ;
        RECT 38.205 163.110 40.950 163.250 ;
        RECT 38.205 163.065 38.495 163.110 ;
        RECT 34.050 162.910 34.370 162.970 ;
        RECT 36.350 162.910 36.670 162.970 ;
        RECT 37.745 162.910 38.035 162.955 ;
        RECT 34.050 162.770 38.035 162.910 ;
        RECT 34.050 162.710 34.370 162.770 ;
        RECT 36.350 162.710 36.670 162.770 ;
        RECT 37.745 162.725 38.035 162.770 ;
        RECT 40.030 162.710 40.350 162.970 ;
        RECT 40.810 162.955 40.950 163.110 ;
        RECT 42.740 163.110 46.290 163.250 ;
        RECT 42.740 163.065 43.110 163.110 ;
        RECT 46.000 163.065 46.290 163.110 ;
        RECT 46.920 163.250 47.210 163.295 ;
        RECT 48.780 163.250 49.070 163.295 ;
        RECT 46.920 163.110 49.070 163.250 ;
        RECT 46.920 163.065 47.210 163.110 ;
        RECT 48.780 163.065 49.070 163.110 ;
        RECT 51.070 163.250 51.390 163.310 ;
        RECT 57.040 163.295 57.255 163.450 ;
        RECT 57.970 163.390 58.290 163.650 ;
        RECT 59.440 163.590 59.580 163.790 ;
        RECT 59.810 163.730 60.130 163.990 ;
        RECT 60.745 163.930 61.035 163.975 ;
        RECT 66.710 163.930 67.030 163.990 ;
        RECT 79.590 163.930 79.910 163.990 ;
        RECT 83.360 163.930 83.500 164.070 ;
        RECT 60.745 163.790 70.160 163.930 ;
        RECT 60.745 163.745 61.035 163.790 ;
        RECT 66.710 163.730 67.030 163.790 ;
        RECT 60.270 163.590 60.590 163.650 ;
        RECT 65.330 163.590 65.650 163.650 ;
        RECT 59.440 163.450 65.650 163.590 ;
        RECT 60.270 163.390 60.590 163.450 ;
        RECT 65.330 163.390 65.650 163.450 ;
        RECT 65.805 163.405 66.095 163.635 ;
        RECT 66.265 163.405 66.555 163.635 ;
        RECT 67.170 163.590 67.490 163.650 ;
        RECT 67.170 163.450 68.780 163.590 ;
        RECT 52.860 163.250 53.150 163.295 ;
        RECT 56.120 163.250 56.410 163.295 ;
        RECT 51.070 163.110 56.410 163.250 ;
        RECT 42.790 163.050 43.110 163.065 ;
        RECT 51.070 163.050 51.390 163.110 ;
        RECT 52.860 163.065 53.150 163.110 ;
        RECT 56.120 163.065 56.410 163.110 ;
        RECT 57.040 163.250 57.330 163.295 ;
        RECT 58.900 163.250 59.190 163.295 ;
        RECT 64.870 163.250 65.190 163.310 ;
        RECT 65.880 163.250 66.020 163.405 ;
        RECT 57.040 163.110 59.190 163.250 ;
        RECT 57.040 163.065 57.330 163.110 ;
        RECT 58.900 163.065 59.190 163.110 ;
        RECT 61.280 163.110 66.020 163.250 ;
        RECT 66.340 163.250 66.480 163.405 ;
        RECT 67.170 163.390 67.490 163.450 ;
        RECT 68.090 163.250 68.410 163.310 ;
        RECT 66.340 163.110 68.410 163.250 ;
        RECT 68.640 163.250 68.780 163.450 ;
        RECT 69.010 163.390 69.330 163.650 ;
        RECT 69.470 163.390 69.790 163.650 ;
        RECT 70.020 163.635 70.160 163.790 ;
        RECT 78.300 163.790 83.500 163.930 ;
        RECT 69.945 163.405 70.235 163.635 ;
        RECT 70.865 163.405 71.155 163.635 ;
        RECT 70.940 163.250 71.080 163.405 ;
        RECT 72.690 163.390 73.010 163.650 ;
        RECT 74.070 163.590 74.390 163.650 ;
        RECT 78.300 163.635 78.440 163.790 ;
        RECT 79.590 163.730 79.910 163.790 ;
        RECT 75.465 163.590 75.755 163.635 ;
        RECT 74.070 163.450 75.755 163.590 ;
        RECT 74.070 163.390 74.390 163.450 ;
        RECT 75.465 163.405 75.755 163.450 ;
        RECT 78.225 163.405 78.515 163.635 ;
        RECT 78.685 163.590 78.975 163.635 ;
        RECT 80.510 163.590 80.830 163.650 ;
        RECT 78.685 163.450 80.830 163.590 ;
        RECT 78.685 163.405 78.975 163.450 ;
        RECT 80.510 163.390 80.830 163.450 ;
        RECT 82.350 163.590 82.670 163.650 ;
        RECT 83.820 163.635 83.960 164.130 ;
        RECT 84.650 164.070 84.970 164.130 ;
        RECT 86.030 163.975 86.350 163.990 ;
        RECT 85.815 163.930 86.350 163.975 ;
        RECT 84.280 163.790 86.350 163.930 ;
        RECT 89.340 163.930 89.480 164.470 ;
        RECT 97.070 164.410 97.390 164.670 ;
        RECT 107.650 164.610 107.970 164.670 ;
        RECT 111.345 164.610 111.635 164.655 ;
        RECT 107.650 164.470 111.635 164.610 ;
        RECT 107.650 164.410 107.970 164.470 ;
        RECT 111.345 164.425 111.635 164.470 ;
        RECT 113.170 164.610 113.490 164.670 ;
        RECT 113.170 164.470 117.080 164.610 ;
        RECT 113.170 164.410 113.490 164.470 ;
        RECT 89.680 164.270 89.970 164.315 ;
        RECT 92.460 164.270 92.750 164.315 ;
        RECT 94.320 164.270 94.610 164.315 ;
        RECT 89.680 164.130 94.610 164.270 ;
        RECT 89.680 164.085 89.970 164.130 ;
        RECT 92.460 164.085 92.750 164.130 ;
        RECT 94.320 164.085 94.610 164.130 ;
        RECT 97.530 164.270 97.850 164.330 ;
        RECT 110.870 164.270 111.190 164.330 ;
        RECT 116.390 164.270 116.710 164.330 ;
        RECT 97.530 164.130 110.180 164.270 ;
        RECT 97.530 164.070 97.850 164.130 ;
        RECT 92.945 163.930 93.235 163.975 ;
        RECT 93.850 163.930 94.170 163.990 ;
        RECT 89.340 163.790 92.700 163.930 ;
        RECT 84.280 163.635 84.420 163.790 ;
        RECT 85.815 163.745 86.350 163.790 ;
        RECT 86.030 163.730 86.350 163.745 ;
        RECT 83.285 163.590 83.575 163.635 ;
        RECT 82.350 163.450 83.575 163.590 ;
        RECT 82.350 163.390 82.670 163.450 ;
        RECT 83.285 163.405 83.575 163.450 ;
        RECT 83.745 163.405 84.035 163.635 ;
        RECT 84.205 163.405 84.495 163.635 ;
        RECT 85.125 163.405 85.415 163.635 ;
        RECT 89.680 163.590 89.970 163.635 ;
        RECT 92.560 163.590 92.700 163.790 ;
        RECT 92.945 163.790 94.170 163.930 ;
        RECT 92.945 163.745 93.235 163.790 ;
        RECT 93.850 163.730 94.170 163.790 ;
        RECT 94.785 163.930 95.075 163.975 ;
        RECT 102.590 163.930 102.910 163.990 ;
        RECT 94.785 163.790 102.910 163.930 ;
        RECT 94.785 163.745 95.075 163.790 ;
        RECT 102.590 163.730 102.910 163.790 ;
        RECT 107.650 163.930 107.970 163.990 ;
        RECT 107.650 163.790 109.720 163.930 ;
        RECT 107.650 163.730 107.970 163.790 ;
        RECT 96.610 163.590 96.930 163.650 ;
        RECT 97.530 163.590 97.850 163.650 ;
        RECT 89.680 163.450 92.215 163.590 ;
        RECT 92.560 163.450 96.380 163.590 ;
        RECT 89.680 163.405 89.970 163.450 ;
        RECT 85.200 163.250 85.340 163.405 ;
        RECT 86.030 163.250 86.350 163.310 ;
        RECT 91.090 163.295 91.410 163.310 ;
        RECT 68.640 163.110 71.080 163.250 ;
        RECT 61.280 162.970 61.420 163.110 ;
        RECT 64.870 163.050 65.190 163.110 ;
        RECT 68.090 163.050 68.410 163.110 ;
        RECT 40.735 162.910 41.025 162.955 ;
        RECT 49.230 162.910 49.550 162.970 ;
        RECT 40.735 162.770 49.550 162.910 ;
        RECT 40.735 162.725 41.025 162.770 ;
        RECT 49.230 162.710 49.550 162.770 ;
        RECT 55.210 162.910 55.530 162.970 ;
        RECT 61.190 162.910 61.510 162.970 ;
        RECT 55.210 162.770 61.510 162.910 ;
        RECT 55.210 162.710 55.530 162.770 ;
        RECT 61.190 162.710 61.510 162.770 ;
        RECT 63.950 162.710 64.270 162.970 ;
        RECT 65.330 162.910 65.650 162.970 ;
        RECT 67.645 162.910 67.935 162.955 ;
        RECT 65.330 162.770 67.935 162.910 ;
        RECT 70.940 162.910 71.080 163.110 ;
        RECT 74.620 163.110 86.350 163.250 ;
        RECT 74.620 162.955 74.760 163.110 ;
        RECT 86.030 163.050 86.350 163.110 ;
        RECT 87.820 163.250 88.110 163.295 ;
        RECT 91.080 163.250 91.410 163.295 ;
        RECT 87.820 163.110 91.410 163.250 ;
        RECT 87.820 163.065 88.110 163.110 ;
        RECT 91.080 163.065 91.410 163.110 ;
        RECT 92.000 163.295 92.215 163.450 ;
        RECT 92.000 163.250 92.290 163.295 ;
        RECT 93.860 163.250 94.150 163.295 ;
        RECT 92.000 163.110 94.150 163.250 ;
        RECT 96.240 163.250 96.380 163.450 ;
        RECT 96.610 163.450 97.850 163.590 ;
        RECT 96.610 163.390 96.930 163.450 ;
        RECT 97.530 163.390 97.850 163.450 ;
        RECT 97.990 163.390 98.310 163.650 ;
        RECT 98.910 163.390 99.230 163.650 ;
        RECT 99.370 163.390 99.690 163.650 ;
        RECT 99.845 163.405 100.135 163.635 ;
        RECT 103.510 163.590 103.830 163.650 ;
        RECT 103.985 163.590 104.275 163.635 ;
        RECT 103.510 163.450 104.275 163.590 ;
        RECT 99.920 163.250 100.060 163.405 ;
        RECT 103.510 163.390 103.830 163.450 ;
        RECT 103.985 163.405 104.275 163.450 ;
        RECT 104.890 163.390 105.210 163.650 ;
        RECT 105.350 163.590 105.670 163.650 ;
        RECT 109.580 163.635 109.720 163.790 ;
        RECT 106.055 163.590 106.345 163.635 ;
        RECT 108.945 163.600 109.235 163.635 ;
        RECT 108.200 163.590 109.260 163.600 ;
        RECT 105.350 163.450 105.865 163.590 ;
        RECT 106.055 163.460 109.260 163.590 ;
        RECT 106.055 163.450 108.340 163.460 ;
        RECT 105.350 163.390 105.670 163.450 ;
        RECT 106.055 163.405 106.345 163.450 ;
        RECT 106.820 163.250 106.960 163.450 ;
        RECT 96.240 163.110 106.960 163.250 ;
        RECT 92.000 163.065 92.290 163.110 ;
        RECT 93.860 163.065 94.150 163.110 ;
        RECT 91.090 163.050 91.410 163.065 ;
        RECT 107.190 163.050 107.510 163.310 ;
        RECT 74.545 162.910 74.835 162.955 ;
        RECT 70.940 162.770 74.835 162.910 ;
        RECT 65.330 162.710 65.650 162.770 ;
        RECT 67.645 162.725 67.935 162.770 ;
        RECT 74.545 162.725 74.835 162.770 ;
        RECT 77.305 162.910 77.595 162.955 ;
        RECT 79.130 162.910 79.450 162.970 ;
        RECT 77.305 162.770 79.450 162.910 ;
        RECT 77.305 162.725 77.595 162.770 ;
        RECT 79.130 162.710 79.450 162.770 ;
        RECT 81.430 162.910 81.750 162.970 ;
        RECT 81.905 162.910 82.195 162.955 ;
        RECT 81.430 162.770 82.195 162.910 ;
        RECT 81.430 162.710 81.750 162.770 ;
        RECT 81.905 162.725 82.195 162.770 ;
        RECT 100.290 162.910 100.610 162.970 ;
        RECT 101.225 162.910 101.515 162.955 ;
        RECT 100.290 162.770 101.515 162.910 ;
        RECT 100.290 162.710 100.610 162.770 ;
        RECT 101.225 162.725 101.515 162.770 ;
        RECT 106.730 162.910 107.050 162.970 ;
        RECT 107.665 162.910 107.955 162.955 ;
        RECT 106.730 162.770 107.955 162.910 ;
        RECT 108.200 162.910 108.340 163.450 ;
        RECT 108.945 163.450 109.260 163.460 ;
        RECT 108.945 163.405 109.235 163.450 ;
        RECT 109.490 163.405 109.780 163.635 ;
        RECT 110.040 163.620 110.180 164.130 ;
        RECT 110.870 164.130 112.940 164.270 ;
        RECT 110.870 164.070 111.190 164.130 ;
        RECT 112.250 163.930 112.570 163.990 ;
        RECT 111.420 163.790 112.570 163.930 ;
        RECT 109.965 163.390 110.255 163.620 ;
        RECT 110.855 163.600 111.145 163.635 ;
        RECT 111.420 163.600 111.560 163.790 ;
        RECT 112.250 163.730 112.570 163.790 ;
        RECT 112.800 163.650 112.940 164.130 ;
        RECT 115.995 164.130 116.710 164.270 ;
        RECT 114.090 163.930 114.410 163.990 ;
        RECT 114.090 163.790 114.780 163.930 ;
        RECT 114.090 163.730 114.410 163.790 ;
        RECT 110.855 163.460 111.560 163.600 ;
        RECT 112.710 163.590 113.030 163.650 ;
        RECT 110.855 163.405 111.145 163.460 ;
        RECT 111.880 163.450 113.030 163.590 ;
        RECT 111.880 162.910 112.020 163.450 ;
        RECT 112.710 163.390 113.030 163.450 ;
        RECT 113.170 163.390 113.490 163.650 ;
        RECT 114.640 163.635 114.780 163.790 ;
        RECT 115.995 163.635 116.135 164.130 ;
        RECT 116.390 164.070 116.710 164.130 ;
        RECT 116.940 163.930 117.080 164.470 ;
        RECT 116.480 163.790 117.080 163.930 ;
        RECT 116.480 163.635 116.620 163.790 ;
        RECT 113.645 163.590 113.935 163.635 ;
        RECT 114.565 163.590 114.855 163.635 ;
        RECT 115.025 163.590 115.315 163.635 ;
        RECT 113.645 163.450 114.320 163.590 ;
        RECT 113.645 163.405 113.935 163.450 ;
        RECT 114.180 163.250 114.320 163.450 ;
        RECT 114.565 163.450 115.315 163.590 ;
        RECT 114.565 163.405 114.855 163.450 ;
        RECT 115.025 163.405 115.315 163.450 ;
        RECT 115.945 163.405 116.235 163.635 ;
        RECT 116.405 163.405 116.695 163.635 ;
        RECT 116.850 163.390 117.170 163.650 ;
        RECT 118.690 163.250 119.010 163.310 ;
        RECT 114.180 163.110 119.010 163.250 ;
        RECT 118.690 163.050 119.010 163.110 ;
        RECT 108.200 162.770 112.020 162.910 ;
        RECT 112.250 162.910 112.570 162.970 ;
        RECT 118.245 162.910 118.535 162.955 ;
        RECT 112.250 162.770 118.535 162.910 ;
        RECT 106.730 162.710 107.050 162.770 ;
        RECT 107.665 162.725 107.955 162.770 ;
        RECT 112.250 162.710 112.570 162.770 ;
        RECT 118.245 162.725 118.535 162.770 ;
        RECT 29.840 162.090 127.820 162.570 ;
        RECT 42.345 161.890 42.635 161.935 ;
        RECT 42.790 161.890 43.110 161.950 ;
        RECT 42.345 161.750 43.110 161.890 ;
        RECT 42.345 161.705 42.635 161.750 ;
        RECT 42.790 161.690 43.110 161.750 ;
        RECT 50.610 161.690 50.930 161.950 ;
        RECT 55.225 161.890 55.515 161.935 ;
        RECT 57.050 161.890 57.370 161.950 ;
        RECT 55.225 161.750 57.370 161.890 ;
        RECT 55.225 161.705 55.515 161.750 ;
        RECT 57.050 161.690 57.370 161.750 ;
        RECT 79.130 161.890 79.450 161.950 ;
        RECT 96.150 161.890 96.470 161.950 ;
        RECT 79.130 161.750 96.470 161.890 ;
        RECT 79.130 161.690 79.450 161.750 ;
        RECT 96.150 161.690 96.470 161.750 ;
        RECT 107.205 161.890 107.495 161.935 ;
        RECT 109.030 161.890 109.350 161.950 ;
        RECT 120.070 161.890 120.390 161.950 ;
        RECT 107.205 161.750 109.350 161.890 ;
        RECT 107.205 161.705 107.495 161.750 ;
        RECT 109.030 161.690 109.350 161.750 ;
        RECT 109.580 161.750 120.390 161.890 ;
        RECT 36.350 161.550 36.670 161.610 ;
        RECT 49.230 161.550 49.550 161.610 ;
        RECT 56.130 161.550 56.450 161.610 ;
        RECT 67.170 161.550 67.490 161.610 ;
        RECT 36.350 161.410 42.560 161.550 ;
        RECT 36.350 161.350 36.670 161.410 ;
        RECT 35.430 161.210 35.750 161.270 ;
        RECT 36.825 161.210 37.115 161.255 ;
        RECT 35.430 161.070 37.115 161.210 ;
        RECT 35.430 161.010 35.750 161.070 ;
        RECT 36.825 161.025 37.115 161.070 ;
        RECT 40.030 161.210 40.350 161.270 ;
        RECT 41.425 161.210 41.715 161.255 ;
        RECT 40.030 161.070 41.715 161.210 ;
        RECT 36.900 160.870 37.040 161.025 ;
        RECT 40.030 161.010 40.350 161.070 ;
        RECT 41.425 161.025 41.715 161.070 ;
        RECT 41.870 161.010 42.190 161.270 ;
        RECT 41.960 160.870 42.100 161.010 ;
        RECT 36.900 160.730 42.100 160.870 ;
        RECT 42.420 160.870 42.560 161.410 ;
        RECT 43.800 161.410 47.160 161.550 ;
        RECT 43.295 161.210 43.585 161.255 ;
        RECT 43.800 161.210 43.940 161.410 ;
        RECT 47.020 161.270 47.160 161.410 ;
        RECT 47.940 161.410 49.550 161.550 ;
        RECT 43.295 161.070 43.940 161.210 ;
        RECT 43.295 161.025 43.585 161.070 ;
        RECT 44.185 161.025 44.475 161.255 ;
        RECT 44.645 161.025 44.935 161.255 ;
        RECT 44.260 160.870 44.400 161.025 ;
        RECT 42.420 160.730 44.400 160.870 ;
        RECT 44.170 160.530 44.490 160.590 ;
        RECT 44.720 160.530 44.860 161.025 ;
        RECT 45.090 161.010 45.410 161.270 ;
        RECT 46.930 161.010 47.250 161.270 ;
        RECT 47.940 161.255 48.080 161.410 ;
        RECT 49.230 161.350 49.550 161.410 ;
        RECT 49.780 161.410 57.050 161.550 ;
        RECT 47.865 161.025 48.155 161.255 ;
        RECT 48.310 161.010 48.630 161.270 ;
        RECT 48.785 161.210 49.075 161.255 ;
        RECT 49.780 161.210 49.920 161.410 ;
        RECT 56.130 161.350 56.450 161.410 ;
        RECT 48.785 161.070 49.920 161.210 ;
        RECT 50.150 161.210 50.470 161.270 ;
        RECT 51.545 161.210 51.835 161.255 ;
        RECT 50.150 161.070 51.835 161.210 ;
        RECT 48.785 161.025 49.075 161.070 ;
        RECT 45.180 160.870 45.320 161.010 ;
        RECT 48.860 160.870 49.000 161.025 ;
        RECT 50.150 161.010 50.470 161.070 ;
        RECT 51.545 161.025 51.835 161.070 ;
        RECT 54.305 161.210 54.595 161.255 ;
        RECT 55.670 161.210 55.990 161.270 ;
        RECT 54.305 161.070 55.990 161.210 ;
        RECT 56.910 161.255 57.050 161.410 ;
        RECT 59.900 161.410 67.490 161.550 ;
        RECT 56.910 161.230 57.255 161.255 ;
        RECT 56.910 161.090 57.280 161.230 ;
        RECT 54.305 161.025 54.595 161.070 ;
        RECT 55.670 161.010 55.990 161.070 ;
        RECT 56.965 161.070 57.280 161.090 ;
        RECT 56.965 161.025 57.255 161.070 ;
        RECT 57.510 161.010 57.830 161.270 ;
        RECT 57.970 161.040 58.290 161.300 ;
        RECT 59.900 161.270 60.040 161.410 ;
        RECT 58.905 161.210 59.195 161.255 ;
        RECT 59.810 161.210 60.130 161.270 ;
        RECT 58.905 161.070 60.130 161.210 ;
        RECT 58.905 161.025 59.195 161.070 ;
        RECT 59.810 161.010 60.130 161.070 ;
        RECT 60.270 161.210 60.590 161.270 ;
        RECT 60.745 161.210 61.035 161.255 ;
        RECT 60.270 161.070 61.035 161.210 ;
        RECT 60.270 161.010 60.590 161.070 ;
        RECT 60.745 161.025 61.035 161.070 ;
        RECT 61.190 161.010 61.510 161.270 ;
        RECT 61.650 161.010 61.970 161.270 ;
        RECT 62.660 161.255 62.800 161.410 ;
        RECT 67.170 161.350 67.490 161.410 ;
        RECT 73.150 161.350 73.470 161.610 ;
        RECT 98.105 161.550 98.395 161.595 ;
        RECT 101.345 161.550 101.995 161.595 ;
        RECT 98.105 161.410 101.995 161.550 ;
        RECT 98.105 161.365 98.695 161.410 ;
        RECT 101.345 161.365 101.995 161.410 ;
        RECT 102.590 161.550 102.910 161.610 ;
        RECT 105.810 161.550 106.130 161.610 ;
        RECT 109.580 161.550 109.720 161.750 ;
        RECT 120.070 161.690 120.390 161.750 ;
        RECT 116.405 161.550 116.695 161.595 ;
        RECT 118.805 161.550 119.095 161.595 ;
        RECT 122.045 161.550 122.695 161.595 ;
        RECT 102.590 161.410 105.580 161.550 ;
        RECT 98.405 161.270 98.695 161.365 ;
        RECT 102.590 161.350 102.910 161.410 ;
        RECT 62.585 161.025 62.875 161.255 ;
        RECT 63.950 161.210 64.270 161.270 ;
        RECT 67.630 161.210 67.950 161.270 ;
        RECT 63.950 161.070 67.950 161.210 ;
        RECT 63.950 161.010 64.270 161.070 ;
        RECT 67.630 161.010 67.950 161.070 ;
        RECT 68.105 161.210 68.395 161.255 ;
        RECT 69.010 161.210 69.330 161.270 ;
        RECT 68.105 161.070 69.330 161.210 ;
        RECT 68.105 161.025 68.395 161.070 ;
        RECT 69.010 161.010 69.330 161.070 ;
        RECT 72.705 161.210 72.995 161.255 ;
        RECT 74.070 161.210 74.390 161.270 ;
        RECT 72.705 161.070 74.390 161.210 ;
        RECT 72.705 161.025 72.995 161.070 ;
        RECT 74.070 161.010 74.390 161.070 ;
        RECT 81.890 161.010 82.210 161.270 ;
        RECT 82.350 161.210 82.670 161.270 ;
        RECT 84.205 161.210 84.495 161.255 ;
        RECT 82.350 161.070 84.495 161.210 ;
        RECT 82.350 161.010 82.670 161.070 ;
        RECT 84.205 161.025 84.495 161.070 ;
        RECT 84.650 161.010 84.970 161.270 ;
        RECT 85.110 161.010 85.430 161.270 ;
        RECT 86.030 161.010 86.350 161.270 ;
        RECT 92.945 161.210 93.235 161.255 ;
        RECT 94.310 161.210 94.630 161.270 ;
        RECT 92.945 161.070 94.630 161.210 ;
        RECT 92.945 161.025 93.235 161.070 ;
        RECT 94.310 161.010 94.630 161.070 ;
        RECT 98.405 161.050 98.770 161.270 ;
        RECT 105.440 161.255 105.580 161.410 ;
        RECT 105.810 161.410 109.720 161.550 ;
        RECT 110.040 161.410 111.560 161.550 ;
        RECT 105.810 161.350 106.130 161.410 ;
        RECT 98.450 161.010 98.770 161.050 ;
        RECT 99.485 161.210 99.775 161.255 ;
        RECT 103.065 161.210 103.355 161.255 ;
        RECT 104.900 161.210 105.190 161.255 ;
        RECT 99.485 161.070 105.190 161.210 ;
        RECT 99.485 161.025 99.775 161.070 ;
        RECT 103.065 161.025 103.355 161.070 ;
        RECT 104.900 161.025 105.190 161.070 ;
        RECT 105.365 161.025 105.655 161.255 ;
        RECT 108.570 161.010 108.890 161.270 ;
        RECT 109.045 161.025 109.335 161.255 ;
        RECT 109.505 161.210 109.795 161.255 ;
        RECT 110.040 161.210 110.180 161.410 ;
        RECT 109.505 161.070 110.180 161.210 ;
        RECT 109.505 161.025 109.795 161.070 ;
        RECT 110.425 161.025 110.715 161.255 ;
        RECT 79.130 160.870 79.450 160.930 ;
        RECT 97.990 160.870 98.310 160.930 ;
        RECT 103.510 160.870 103.830 160.930 ;
        RECT 45.180 160.730 49.000 160.870 ;
        RECT 60.820 160.730 79.450 160.870 ;
        RECT 60.820 160.590 60.960 160.730 ;
        RECT 79.130 160.670 79.450 160.730 ;
        RECT 79.680 160.730 103.830 160.870 ;
        RECT 48.310 160.530 48.630 160.590 ;
        RECT 44.170 160.390 48.630 160.530 ;
        RECT 44.170 160.330 44.490 160.390 ;
        RECT 48.310 160.330 48.630 160.390 ;
        RECT 48.860 160.390 60.040 160.530 ;
        RECT 35.890 160.190 36.210 160.250 ;
        RECT 36.365 160.190 36.655 160.235 ;
        RECT 35.890 160.050 36.655 160.190 ;
        RECT 35.890 159.990 36.210 160.050 ;
        RECT 36.365 160.005 36.655 160.050 ;
        RECT 39.570 160.190 39.890 160.250 ;
        RECT 40.505 160.190 40.795 160.235 ;
        RECT 39.570 160.050 40.795 160.190 ;
        RECT 39.570 159.990 39.890 160.050 ;
        RECT 40.505 160.005 40.795 160.050 ;
        RECT 46.470 159.990 46.790 160.250 ;
        RECT 46.930 160.190 47.250 160.250 ;
        RECT 48.860 160.190 49.000 160.390 ;
        RECT 46.930 160.050 49.000 160.190 ;
        RECT 46.930 159.990 47.250 160.050 ;
        RECT 50.150 159.990 50.470 160.250 ;
        RECT 55.685 160.190 55.975 160.235 ;
        RECT 57.050 160.190 57.370 160.250 ;
        RECT 55.685 160.050 57.370 160.190 ;
        RECT 55.685 160.005 55.975 160.050 ;
        RECT 57.050 159.990 57.370 160.050 ;
        RECT 58.890 160.190 59.210 160.250 ;
        RECT 59.365 160.190 59.655 160.235 ;
        RECT 58.890 160.050 59.655 160.190 ;
        RECT 59.900 160.190 60.040 160.390 ;
        RECT 60.730 160.330 61.050 160.590 ;
        RECT 65.790 160.530 66.110 160.590 ;
        RECT 71.785 160.530 72.075 160.575 ;
        RECT 79.680 160.530 79.820 160.730 ;
        RECT 97.990 160.670 98.310 160.730 ;
        RECT 103.510 160.670 103.830 160.730 ;
        RECT 103.970 160.670 104.290 160.930 ;
        RECT 108.110 160.870 108.430 160.930 ;
        RECT 109.120 160.870 109.260 161.025 ;
        RECT 108.110 160.730 109.260 160.870 ;
        RECT 108.110 160.670 108.430 160.730 ;
        RECT 65.790 160.390 79.820 160.530 ;
        RECT 84.190 160.530 84.510 160.590 ;
        RECT 98.910 160.530 99.230 160.590 ;
        RECT 84.190 160.390 99.230 160.530 ;
        RECT 65.790 160.330 66.110 160.390 ;
        RECT 71.785 160.345 72.075 160.390 ;
        RECT 84.190 160.330 84.510 160.390 ;
        RECT 98.910 160.330 99.230 160.390 ;
        RECT 99.485 160.530 99.775 160.575 ;
        RECT 102.605 160.530 102.895 160.575 ;
        RECT 104.495 160.530 104.785 160.575 ;
        RECT 99.485 160.390 104.785 160.530 ;
        RECT 99.485 160.345 99.775 160.390 ;
        RECT 102.605 160.345 102.895 160.390 ;
        RECT 104.495 160.345 104.785 160.390 ;
        RECT 105.810 160.530 106.130 160.590 ;
        RECT 110.500 160.530 110.640 161.025 ;
        RECT 111.420 160.915 111.560 161.410 ;
        RECT 116.405 161.410 122.695 161.550 ;
        RECT 116.405 161.365 116.695 161.410 ;
        RECT 118.805 161.365 119.395 161.410 ;
        RECT 122.045 161.365 122.695 161.410 ;
        RECT 115.930 161.010 116.250 161.270 ;
        RECT 119.105 161.050 119.395 161.365 ;
        RECT 120.185 161.210 120.475 161.255 ;
        RECT 123.765 161.210 124.055 161.255 ;
        RECT 125.600 161.210 125.890 161.255 ;
        RECT 120.185 161.070 125.890 161.210 ;
        RECT 120.185 161.025 120.475 161.070 ;
        RECT 123.765 161.025 124.055 161.070 ;
        RECT 125.600 161.025 125.890 161.070 ;
        RECT 126.050 161.010 126.370 161.270 ;
        RECT 111.345 160.870 111.635 160.915 ;
        RECT 117.325 160.870 117.615 160.915 ;
        RECT 111.345 160.730 117.615 160.870 ;
        RECT 111.345 160.685 111.635 160.730 ;
        RECT 117.325 160.685 117.615 160.730 ;
        RECT 124.670 160.670 124.990 160.930 ;
        RECT 112.710 160.530 113.030 160.590 ;
        RECT 105.810 160.390 113.030 160.530 ;
        RECT 105.810 160.330 106.130 160.390 ;
        RECT 112.710 160.330 113.030 160.390 ;
        RECT 120.185 160.530 120.475 160.575 ;
        RECT 123.305 160.530 123.595 160.575 ;
        RECT 125.195 160.530 125.485 160.575 ;
        RECT 120.185 160.390 125.485 160.530 ;
        RECT 120.185 160.345 120.475 160.390 ;
        RECT 123.305 160.345 123.595 160.390 ;
        RECT 125.195 160.345 125.485 160.390 ;
        RECT 65.880 160.190 66.020 160.330 ;
        RECT 59.900 160.050 66.020 160.190 ;
        RECT 67.185 160.190 67.475 160.235 ;
        RECT 67.630 160.190 67.950 160.250 ;
        RECT 67.185 160.050 67.950 160.190 ;
        RECT 58.890 159.990 59.210 160.050 ;
        RECT 59.365 160.005 59.655 160.050 ;
        RECT 67.185 160.005 67.475 160.050 ;
        RECT 67.630 159.990 67.950 160.050 ;
        RECT 69.025 160.190 69.315 160.235 ;
        RECT 70.390 160.190 70.710 160.250 ;
        RECT 69.025 160.050 70.710 160.190 ;
        RECT 69.025 160.005 69.315 160.050 ;
        RECT 70.390 159.990 70.710 160.050 ;
        RECT 82.350 160.190 82.670 160.250 ;
        RECT 82.825 160.190 83.115 160.235 ;
        RECT 82.350 160.050 83.115 160.190 ;
        RECT 82.350 159.990 82.670 160.050 ;
        RECT 82.825 160.005 83.115 160.050 ;
        RECT 92.485 160.190 92.775 160.235 ;
        RECT 93.850 160.190 94.170 160.250 ;
        RECT 92.485 160.050 94.170 160.190 ;
        RECT 92.485 160.005 92.775 160.050 ;
        RECT 93.850 159.990 94.170 160.050 ;
        RECT 96.610 159.990 96.930 160.250 ;
        RECT 99.000 160.190 99.140 160.330 ;
        RECT 108.110 160.190 108.430 160.250 ;
        RECT 109.490 160.190 109.810 160.250 ;
        RECT 99.000 160.050 109.810 160.190 ;
        RECT 108.110 159.990 108.430 160.050 ;
        RECT 109.490 159.990 109.810 160.050 ;
        RECT 114.105 160.190 114.395 160.235 ;
        RECT 115.470 160.190 115.790 160.250 ;
        RECT 114.105 160.050 115.790 160.190 ;
        RECT 114.105 160.005 114.395 160.050 ;
        RECT 115.470 159.990 115.790 160.050 ;
        RECT 29.840 159.370 127.820 159.850 ;
        RECT 32.455 159.170 32.745 159.215 ;
        RECT 34.050 159.170 34.370 159.230 ;
        RECT 32.455 159.030 34.370 159.170 ;
        RECT 32.455 158.985 32.745 159.030 ;
        RECT 34.050 158.970 34.370 159.030 ;
        RECT 53.830 158.970 54.150 159.230 ;
        RECT 79.145 159.170 79.435 159.215 ;
        RECT 79.590 159.170 79.910 159.230 ;
        RECT 79.145 159.030 79.910 159.170 ;
        RECT 79.145 158.985 79.435 159.030 ;
        RECT 79.590 158.970 79.910 159.030 ;
        RECT 84.665 159.170 84.955 159.215 ;
        RECT 86.490 159.170 86.810 159.230 ;
        RECT 84.665 159.030 86.810 159.170 ;
        RECT 84.665 158.985 84.955 159.030 ;
        RECT 86.490 158.970 86.810 159.030 ;
        RECT 98.450 159.170 98.770 159.230 ;
        RECT 99.845 159.170 100.135 159.215 ;
        RECT 98.450 159.030 100.135 159.170 ;
        RECT 98.450 158.970 98.770 159.030 ;
        RECT 99.845 158.985 100.135 159.030 ;
        RECT 105.350 159.170 105.670 159.230 ;
        RECT 106.745 159.170 107.035 159.215 ;
        RECT 105.350 159.030 107.035 159.170 ;
        RECT 105.350 158.970 105.670 159.030 ;
        RECT 106.745 158.985 107.035 159.030 ;
        RECT 124.670 158.970 124.990 159.230 ;
        RECT 36.320 158.830 36.610 158.875 ;
        RECT 39.100 158.830 39.390 158.875 ;
        RECT 40.960 158.830 41.250 158.875 ;
        RECT 59.365 158.830 59.655 158.875 ;
        RECT 64.870 158.830 65.190 158.890 ;
        RECT 36.320 158.690 41.250 158.830 ;
        RECT 36.320 158.645 36.610 158.690 ;
        RECT 39.100 158.645 39.390 158.690 ;
        RECT 40.960 158.645 41.250 158.690 ;
        RECT 53.920 158.690 65.190 158.830 ;
        RECT 39.570 158.290 39.890 158.550 ;
        RECT 36.320 158.150 36.610 158.195 ;
        RECT 41.425 158.150 41.715 158.195 ;
        RECT 42.790 158.150 43.110 158.210 ;
        RECT 53.920 158.195 54.060 158.690 ;
        RECT 59.365 158.645 59.655 158.690 ;
        RECT 64.870 158.630 65.190 158.690 ;
        RECT 67.140 158.830 67.430 158.875 ;
        RECT 69.920 158.830 70.210 158.875 ;
        RECT 71.780 158.830 72.070 158.875 ;
        RECT 67.140 158.690 72.070 158.830 ;
        RECT 67.140 158.645 67.430 158.690 ;
        RECT 69.920 158.645 70.210 158.690 ;
        RECT 71.780 158.645 72.070 158.690 ;
        RECT 74.530 158.830 74.850 158.890 ;
        RECT 76.370 158.830 76.690 158.890 ;
        RECT 91.980 158.830 92.270 158.875 ;
        RECT 94.760 158.830 95.050 158.875 ;
        RECT 96.620 158.830 96.910 158.875 ;
        RECT 74.530 158.690 82.120 158.830 ;
        RECT 74.530 158.630 74.850 158.690 ;
        RECT 76.370 158.630 76.690 158.690 ;
        RECT 54.750 158.290 55.070 158.550 ;
        RECT 70.390 158.290 70.710 158.550 ;
        RECT 80.510 158.490 80.830 158.550 ;
        RECT 81.980 158.535 82.120 158.690 ;
        RECT 91.980 158.690 96.910 158.830 ;
        RECT 91.980 158.645 92.270 158.690 ;
        RECT 94.760 158.645 95.050 158.690 ;
        RECT 96.620 158.645 96.910 158.690 ;
        RECT 105.825 158.830 106.115 158.875 ;
        RECT 120.530 158.830 120.850 158.890 ;
        RECT 105.825 158.690 120.850 158.830 ;
        RECT 105.825 158.645 106.115 158.690 ;
        RECT 120.530 158.630 120.850 158.690 ;
        RECT 121.005 158.645 121.295 158.875 ;
        RECT 78.300 158.350 80.830 158.490 ;
        RECT 36.320 158.010 38.855 158.150 ;
        RECT 36.320 157.965 36.610 158.010 ;
        RECT 34.460 157.810 34.750 157.855 ;
        RECT 35.890 157.810 36.210 157.870 ;
        RECT 38.640 157.855 38.855 158.010 ;
        RECT 41.425 158.010 43.110 158.150 ;
        RECT 41.425 157.965 41.715 158.010 ;
        RECT 42.790 157.950 43.110 158.010 ;
        RECT 53.845 157.965 54.135 158.195 ;
        RECT 55.670 158.150 55.990 158.210 ;
        RECT 60.730 158.150 61.050 158.210 ;
        RECT 55.670 158.010 61.050 158.150 ;
        RECT 55.670 157.950 55.990 158.010 ;
        RECT 60.730 157.950 61.050 158.010 ;
        RECT 61.205 157.965 61.495 158.195 ;
        RECT 37.720 157.810 38.010 157.855 ;
        RECT 34.460 157.670 38.010 157.810 ;
        RECT 34.460 157.625 34.750 157.670 ;
        RECT 35.890 157.610 36.210 157.670 ;
        RECT 37.720 157.625 38.010 157.670 ;
        RECT 38.640 157.810 38.930 157.855 ;
        RECT 40.500 157.810 40.790 157.855 ;
        RECT 38.640 157.670 40.790 157.810 ;
        RECT 38.640 157.625 38.930 157.670 ;
        RECT 40.500 157.625 40.790 157.670 ;
        RECT 53.370 157.810 53.690 157.870 ;
        RECT 55.225 157.810 55.515 157.855 ;
        RECT 53.370 157.670 55.515 157.810 ;
        RECT 53.370 157.610 53.690 157.670 ;
        RECT 55.225 157.625 55.515 157.670 ;
        RECT 44.630 157.470 44.950 157.530 ;
        RECT 52.925 157.470 53.215 157.515 ;
        RECT 44.630 157.330 53.215 157.470 ;
        RECT 44.630 157.270 44.950 157.330 ;
        RECT 52.925 157.285 53.215 157.330 ;
        RECT 54.750 157.470 55.070 157.530 ;
        RECT 61.280 157.470 61.420 157.965 ;
        RECT 61.650 157.950 61.970 158.210 ;
        RECT 62.585 158.150 62.875 158.195 ;
        RECT 65.790 158.150 66.110 158.210 ;
        RECT 62.585 158.010 66.110 158.150 ;
        RECT 62.585 157.965 62.875 158.010 ;
        RECT 65.790 157.950 66.110 158.010 ;
        RECT 67.140 158.150 67.430 158.195 ;
        RECT 72.245 158.150 72.535 158.195 ;
        RECT 73.610 158.150 73.930 158.210 ;
        RECT 78.300 158.195 78.440 158.350 ;
        RECT 80.510 158.290 80.830 158.350 ;
        RECT 81.905 158.305 82.195 158.535 ;
        RECT 84.665 158.490 84.955 158.535 ;
        RECT 85.570 158.490 85.890 158.550 ;
        RECT 84.665 158.350 85.890 158.490 ;
        RECT 84.665 158.305 84.955 158.350 ;
        RECT 85.570 158.290 85.890 158.350 ;
        RECT 107.650 158.290 107.970 158.550 ;
        RECT 109.490 158.490 109.810 158.550 ;
        RECT 116.405 158.490 116.695 158.535 ;
        RECT 117.770 158.490 118.090 158.550 ;
        RECT 109.490 158.350 110.640 158.490 ;
        RECT 109.490 158.290 109.810 158.350 ;
        RECT 67.140 158.010 69.675 158.150 ;
        RECT 67.140 157.965 67.430 158.010 ;
        RECT 61.740 157.810 61.880 157.950 ;
        RECT 63.275 157.810 63.565 157.855 ;
        RECT 61.740 157.670 63.565 157.810 ;
        RECT 63.275 157.625 63.565 157.670 ;
        RECT 65.280 157.810 65.570 157.855 ;
        RECT 67.630 157.810 67.950 157.870 ;
        RECT 69.460 157.855 69.675 158.010 ;
        RECT 72.245 158.010 73.930 158.150 ;
        RECT 72.245 157.965 72.535 158.010 ;
        RECT 73.610 157.950 73.930 158.010 ;
        RECT 77.765 157.965 78.055 158.195 ;
        RECT 78.225 157.965 78.515 158.195 ;
        RECT 80.050 158.150 80.370 158.210 ;
        RECT 81.445 158.150 81.735 158.195 ;
        RECT 83.270 158.150 83.590 158.210 ;
        RECT 78.760 158.010 80.565 158.150 ;
        RECT 81.445 158.010 83.590 158.150 ;
        RECT 68.540 157.810 68.830 157.855 ;
        RECT 65.280 157.670 68.830 157.810 ;
        RECT 65.280 157.625 65.570 157.670 ;
        RECT 67.630 157.610 67.950 157.670 ;
        RECT 68.540 157.625 68.830 157.670 ;
        RECT 69.460 157.810 69.750 157.855 ;
        RECT 71.320 157.810 71.610 157.855 ;
        RECT 69.460 157.670 71.610 157.810 ;
        RECT 77.840 157.810 77.980 157.965 ;
        RECT 78.760 157.810 78.900 158.010 ;
        RECT 80.050 157.950 80.370 158.010 ;
        RECT 81.445 157.965 81.735 158.010 ;
        RECT 77.840 157.670 78.900 157.810 ;
        RECT 80.510 157.810 80.830 157.870 ;
        RECT 81.520 157.810 81.660 157.965 ;
        RECT 83.270 157.950 83.590 158.010 ;
        RECT 83.730 157.950 84.050 158.210 ;
        RECT 91.980 158.150 92.270 158.195 ;
        RECT 91.980 158.010 94.515 158.150 ;
        RECT 91.980 157.965 92.270 158.010 ;
        RECT 80.510 157.670 81.660 157.810 ;
        RECT 69.460 157.625 69.750 157.670 ;
        RECT 71.320 157.625 71.610 157.670 ;
        RECT 80.510 157.610 80.830 157.670 ;
        RECT 85.110 157.610 85.430 157.870 ;
        RECT 93.390 157.855 93.710 157.870 ;
        RECT 90.120 157.810 90.410 157.855 ;
        RECT 93.380 157.810 93.710 157.855 ;
        RECT 90.120 157.670 93.710 157.810 ;
        RECT 90.120 157.625 90.410 157.670 ;
        RECT 93.380 157.625 93.710 157.670 ;
        RECT 94.300 157.855 94.515 158.010 ;
        RECT 95.230 157.950 95.550 158.210 ;
        RECT 95.690 158.150 96.010 158.210 ;
        RECT 97.085 158.150 97.375 158.195 ;
        RECT 95.690 158.010 97.375 158.150 ;
        RECT 95.690 157.950 96.010 158.010 ;
        RECT 97.085 157.965 97.375 158.010 ;
        RECT 97.530 158.150 97.850 158.210 ;
        RECT 100.305 158.150 100.595 158.195 ;
        RECT 97.530 158.010 100.595 158.150 ;
        RECT 97.530 157.950 97.850 158.010 ;
        RECT 100.305 157.965 100.595 158.010 ;
        RECT 106.270 158.150 106.590 158.210 ;
        RECT 110.500 158.195 110.640 158.350 ;
        RECT 116.405 158.350 118.090 158.490 ;
        RECT 116.405 158.305 116.695 158.350 ;
        RECT 117.770 158.290 118.090 158.350 ;
        RECT 106.745 158.150 107.035 158.195 ;
        RECT 106.270 158.010 107.035 158.150 ;
        RECT 106.270 157.950 106.590 158.010 ;
        RECT 106.745 157.965 107.035 158.010 ;
        RECT 109.965 157.965 110.255 158.195 ;
        RECT 110.425 157.965 110.715 158.195 ;
        RECT 110.885 157.965 111.175 158.195 ;
        RECT 111.805 158.150 112.095 158.195 ;
        RECT 112.250 158.150 112.570 158.210 ;
        RECT 115.025 158.150 115.315 158.195 ;
        RECT 111.805 158.010 112.570 158.150 ;
        RECT 111.805 157.965 112.095 158.010 ;
        RECT 94.300 157.810 94.590 157.855 ;
        RECT 96.160 157.810 96.450 157.855 ;
        RECT 94.300 157.670 96.450 157.810 ;
        RECT 94.300 157.625 94.590 157.670 ;
        RECT 96.160 157.625 96.450 157.670 ;
        RECT 108.125 157.810 108.415 157.855 ;
        RECT 108.585 157.810 108.875 157.855 ;
        RECT 108.125 157.670 108.875 157.810 ;
        RECT 108.125 157.625 108.415 157.670 ;
        RECT 108.585 157.625 108.875 157.670 ;
        RECT 109.030 157.810 109.350 157.870 ;
        RECT 110.040 157.810 110.180 157.965 ;
        RECT 109.030 157.670 110.180 157.810 ;
        RECT 110.960 157.810 111.100 157.965 ;
        RECT 112.250 157.950 112.570 158.010 ;
        RECT 112.800 158.010 115.315 158.150 ;
        RECT 112.800 157.810 112.940 158.010 ;
        RECT 115.025 157.965 115.315 158.010 ;
        RECT 115.470 158.150 115.790 158.210 ;
        RECT 119.165 158.150 119.455 158.195 ;
        RECT 115.470 158.010 119.455 158.150 ;
        RECT 121.080 158.150 121.220 158.645 ;
        RECT 122.385 158.150 122.675 158.195 ;
        RECT 121.080 158.010 122.675 158.150 ;
        RECT 115.470 157.950 115.790 158.010 ;
        RECT 119.165 157.965 119.455 158.010 ;
        RECT 122.385 157.965 122.675 158.010 ;
        RECT 123.765 157.965 124.055 158.195 ;
        RECT 110.960 157.670 112.940 157.810 ;
        RECT 114.090 157.810 114.410 157.870 ;
        RECT 123.840 157.810 123.980 157.965 ;
        RECT 114.090 157.670 123.980 157.810 ;
        RECT 93.390 157.610 93.710 157.625 ;
        RECT 109.030 157.610 109.350 157.670 ;
        RECT 75.450 157.470 75.770 157.530 ;
        RECT 54.750 157.330 75.770 157.470 ;
        RECT 54.750 157.270 55.070 157.330 ;
        RECT 75.450 157.270 75.770 157.330 ;
        RECT 75.910 157.470 76.230 157.530 ;
        RECT 76.845 157.470 77.135 157.515 ;
        RECT 75.910 157.330 77.135 157.470 ;
        RECT 75.910 157.270 76.230 157.330 ;
        RECT 76.845 157.285 77.135 157.330 ;
        RECT 79.130 157.470 79.450 157.530 ;
        RECT 81.905 157.470 82.195 157.515 ;
        RECT 79.130 157.330 82.195 157.470 ;
        RECT 79.130 157.270 79.450 157.330 ;
        RECT 81.905 157.285 82.195 157.330 ;
        RECT 82.825 157.470 83.115 157.515 ;
        RECT 85.570 157.470 85.890 157.530 ;
        RECT 82.825 157.330 85.890 157.470 ;
        RECT 82.825 157.285 83.115 157.330 ;
        RECT 85.570 157.270 85.890 157.330 ;
        RECT 87.870 157.515 88.190 157.530 ;
        RECT 87.870 157.285 88.405 157.515 ;
        RECT 96.610 157.470 96.930 157.530 ;
        RECT 110.960 157.470 111.100 157.670 ;
        RECT 114.090 157.610 114.410 157.670 ;
        RECT 96.610 157.330 111.100 157.470 ;
        RECT 87.870 157.270 88.190 157.285 ;
        RECT 96.610 157.270 96.930 157.330 ;
        RECT 113.170 157.270 113.490 157.530 ;
        RECT 118.690 157.270 119.010 157.530 ;
        RECT 123.305 157.470 123.595 157.515 ;
        RECT 124.210 157.470 124.530 157.530 ;
        RECT 123.305 157.330 124.530 157.470 ;
        RECT 123.305 157.285 123.595 157.330 ;
        RECT 124.210 157.270 124.530 157.330 ;
        RECT 29.840 156.650 127.820 157.130 ;
        RECT 52.235 156.450 52.525 156.495 ;
        RECT 61.650 156.450 61.970 156.510 ;
        RECT 64.885 156.450 65.175 156.495 ;
        RECT 50.700 156.310 60.960 156.450 ;
        RECT 47.865 156.110 48.155 156.155 ;
        RECT 48.325 156.110 48.615 156.155 ;
        RECT 47.865 155.970 48.615 156.110 ;
        RECT 47.865 155.925 48.155 155.970 ;
        RECT 48.325 155.925 48.615 155.970 ;
        RECT 49.320 155.970 50.380 156.110 ;
        RECT 31.290 155.770 31.610 155.830 ;
        RECT 34.065 155.770 34.355 155.815 ;
        RECT 31.290 155.630 34.355 155.770 ;
        RECT 31.290 155.570 31.610 155.630 ;
        RECT 34.065 155.585 34.355 155.630 ;
        RECT 36.810 155.770 37.130 155.830 ;
        RECT 37.745 155.770 38.035 155.815 ;
        RECT 36.810 155.630 38.035 155.770 ;
        RECT 36.810 155.570 37.130 155.630 ;
        RECT 37.745 155.585 38.035 155.630 ;
        RECT 46.470 155.570 46.790 155.830 ;
        RECT 46.010 155.430 46.330 155.490 ;
        RECT 46.945 155.430 47.235 155.475 ;
        RECT 46.010 155.290 47.235 155.430 ;
        RECT 46.010 155.230 46.330 155.290 ;
        RECT 46.945 155.245 47.235 155.290 ;
        RECT 49.320 155.090 49.460 155.970 ;
        RECT 50.240 155.815 50.380 155.970 ;
        RECT 50.700 155.815 50.840 156.310 ;
        RECT 52.235 156.265 52.525 156.310 ;
        RECT 60.820 156.170 60.960 156.310 ;
        RECT 61.650 156.310 65.175 156.450 ;
        RECT 61.650 156.250 61.970 156.310 ;
        RECT 64.885 156.265 65.175 156.310 ;
        RECT 67.185 156.450 67.475 156.495 ;
        RECT 69.010 156.450 69.330 156.510 ;
        RECT 82.810 156.450 83.130 156.510 ;
        RECT 67.185 156.310 69.330 156.450 ;
        RECT 67.185 156.265 67.475 156.310 ;
        RECT 69.010 156.250 69.330 156.310 ;
        RECT 81.980 156.310 83.130 156.450 ;
        RECT 53.370 156.110 53.690 156.170 ;
        RECT 54.240 156.110 54.530 156.155 ;
        RECT 57.500 156.110 57.790 156.155 ;
        RECT 53.370 155.970 57.790 156.110 ;
        RECT 53.370 155.910 53.690 155.970 ;
        RECT 54.240 155.925 54.530 155.970 ;
        RECT 57.500 155.925 57.790 155.970 ;
        RECT 58.420 156.110 58.710 156.155 ;
        RECT 60.280 156.110 60.570 156.155 ;
        RECT 58.420 155.970 60.570 156.110 ;
        RECT 58.420 155.925 58.710 155.970 ;
        RECT 60.280 155.925 60.570 155.970 ;
        RECT 60.730 156.110 61.050 156.170 ;
        RECT 65.345 156.110 65.635 156.155 ;
        RECT 60.730 155.970 65.635 156.110 ;
        RECT 49.705 155.585 49.995 155.815 ;
        RECT 50.165 155.585 50.455 155.815 ;
        RECT 50.625 155.585 50.915 155.815 ;
        RECT 49.780 155.430 49.920 155.585 ;
        RECT 51.530 155.570 51.850 155.830 ;
        RECT 56.100 155.770 56.390 155.815 ;
        RECT 58.420 155.770 58.635 155.925 ;
        RECT 60.730 155.910 61.050 155.970 ;
        RECT 65.345 155.925 65.635 155.970 ;
        RECT 66.710 156.110 67.030 156.170 ;
        RECT 70.405 156.110 70.695 156.155 ;
        RECT 66.710 155.970 70.695 156.110 ;
        RECT 66.710 155.910 67.030 155.970 ;
        RECT 70.405 155.925 70.695 155.970 ;
        RECT 76.845 156.110 77.135 156.155 ;
        RECT 78.685 156.110 78.975 156.155 ;
        RECT 79.130 156.110 79.450 156.170 ;
        RECT 76.845 155.970 79.450 156.110 ;
        RECT 76.845 155.925 77.135 155.970 ;
        RECT 78.685 155.925 78.975 155.970 ;
        RECT 79.130 155.910 79.450 155.970 ;
        RECT 79.590 156.110 79.910 156.170 ;
        RECT 79.590 155.970 81.660 156.110 ;
        RECT 79.590 155.910 79.910 155.970 ;
        RECT 62.585 155.770 62.875 155.815 ;
        RECT 63.490 155.770 63.810 155.830 ;
        RECT 56.100 155.630 58.635 155.770 ;
        RECT 58.980 155.630 63.810 155.770 ;
        RECT 56.100 155.585 56.390 155.630 ;
        RECT 55.670 155.430 55.990 155.490 ;
        RECT 49.780 155.290 55.990 155.430 ;
        RECT 55.670 155.230 55.990 155.290 ;
        RECT 56.590 155.430 56.910 155.490 ;
        RECT 58.980 155.430 59.120 155.630 ;
        RECT 62.585 155.585 62.875 155.630 ;
        RECT 63.490 155.570 63.810 155.630 ;
        RECT 69.930 155.570 70.250 155.830 ;
        RECT 70.850 155.770 71.170 155.830 ;
        RECT 72.230 155.770 72.550 155.830 ;
        RECT 73.625 155.770 73.915 155.815 ;
        RECT 70.850 155.630 73.915 155.770 ;
        RECT 70.850 155.570 71.170 155.630 ;
        RECT 72.230 155.570 72.550 155.630 ;
        RECT 73.625 155.585 73.915 155.630 ;
        RECT 80.985 155.585 81.275 155.815 ;
        RECT 56.590 155.290 59.120 155.430 ;
        RECT 56.590 155.230 56.910 155.290 ;
        RECT 59.350 155.230 59.670 155.490 ;
        RECT 61.190 155.230 61.510 155.490 ;
        RECT 64.425 155.430 64.715 155.475 ;
        RECT 65.790 155.430 66.110 155.490 ;
        RECT 69.025 155.430 69.315 155.475 ;
        RECT 75.465 155.430 75.755 155.475 ;
        RECT 64.425 155.290 75.755 155.430 ;
        RECT 64.425 155.245 64.715 155.290 ;
        RECT 65.790 155.230 66.110 155.290 ;
        RECT 69.025 155.245 69.315 155.290 ;
        RECT 75.465 155.245 75.755 155.290 ;
        RECT 75.910 155.430 76.230 155.490 ;
        RECT 79.130 155.430 79.450 155.490 ;
        RECT 81.060 155.430 81.200 155.585 ;
        RECT 75.910 155.290 77.980 155.430 ;
        RECT 75.910 155.230 76.230 155.290 ;
        RECT 54.750 155.090 55.070 155.150 ;
        RECT 49.320 154.950 55.070 155.090 ;
        RECT 54.750 154.890 55.070 154.950 ;
        RECT 56.100 155.090 56.390 155.135 ;
        RECT 58.880 155.090 59.170 155.135 ;
        RECT 60.740 155.090 61.030 155.135 ;
        RECT 56.100 154.950 61.030 155.090 ;
        RECT 56.100 154.905 56.390 154.950 ;
        RECT 58.880 154.905 59.170 154.950 ;
        RECT 60.740 154.905 61.030 154.950 ;
        RECT 72.245 155.090 72.535 155.135 ;
        RECT 77.290 155.090 77.610 155.150 ;
        RECT 72.245 154.950 77.610 155.090 ;
        RECT 77.840 155.090 77.980 155.290 ;
        RECT 79.130 155.290 81.200 155.430 ;
        RECT 81.520 155.430 81.660 155.970 ;
        RECT 81.980 155.815 82.120 156.310 ;
        RECT 82.810 156.250 83.130 156.310 ;
        RECT 83.730 156.250 84.050 156.510 ;
        RECT 84.205 156.450 84.495 156.495 ;
        RECT 85.110 156.450 85.430 156.510 ;
        RECT 84.205 156.310 85.430 156.450 ;
        RECT 84.205 156.265 84.495 156.310 ;
        RECT 85.110 156.250 85.430 156.310 ;
        RECT 93.405 156.450 93.695 156.495 ;
        RECT 95.230 156.450 95.550 156.510 ;
        RECT 93.405 156.310 95.550 156.450 ;
        RECT 93.405 156.265 93.695 156.310 ;
        RECT 95.230 156.250 95.550 156.310 ;
        RECT 97.085 156.450 97.375 156.495 ;
        RECT 98.925 156.450 99.215 156.495 ;
        RECT 97.085 156.310 99.215 156.450 ;
        RECT 97.085 156.265 97.375 156.310 ;
        RECT 98.925 156.265 99.215 156.310 ;
        RECT 101.225 156.265 101.515 156.495 ;
        RECT 102.605 156.450 102.895 156.495 ;
        RECT 103.970 156.450 104.290 156.510 ;
        RECT 102.605 156.310 104.290 156.450 ;
        RECT 102.605 156.265 102.895 156.310 ;
        RECT 83.820 156.110 83.960 156.250 ;
        RECT 86.045 156.110 86.335 156.155 ;
        RECT 87.870 156.110 88.190 156.170 ;
        RECT 99.385 156.110 99.675 156.155 ;
        RECT 83.820 155.970 99.675 156.110 ;
        RECT 86.045 155.925 86.335 155.970 ;
        RECT 87.870 155.910 88.190 155.970 ;
        RECT 99.385 155.925 99.675 155.970 ;
        RECT 81.905 155.585 82.195 155.815 ;
        RECT 82.365 155.585 82.655 155.815 ;
        RECT 82.825 155.770 83.115 155.815 ;
        RECT 83.730 155.770 84.050 155.830 ;
        RECT 82.825 155.630 84.050 155.770 ;
        RECT 82.825 155.585 83.115 155.630 ;
        RECT 82.440 155.430 82.580 155.585 ;
        RECT 83.730 155.570 84.050 155.630 ;
        RECT 85.110 155.770 85.430 155.830 ;
        RECT 86.505 155.770 86.795 155.815 ;
        RECT 85.110 155.630 86.795 155.770 ;
        RECT 85.110 155.570 85.430 155.630 ;
        RECT 86.505 155.585 86.795 155.630 ;
        RECT 91.565 155.770 91.855 155.815 ;
        RECT 92.010 155.770 92.330 155.830 ;
        RECT 91.565 155.630 92.330 155.770 ;
        RECT 91.565 155.585 91.855 155.630 ;
        RECT 92.010 155.570 92.330 155.630 ;
        RECT 92.485 155.585 92.775 155.815 ;
        RECT 94.325 155.770 94.615 155.815 ;
        RECT 96.610 155.770 96.930 155.830 ;
        RECT 94.325 155.630 96.930 155.770 ;
        RECT 101.300 155.770 101.440 156.265 ;
        RECT 103.970 156.250 104.290 156.310 ;
        RECT 114.090 156.250 114.410 156.510 ;
        RECT 111.790 156.110 112.110 156.170 ;
        RECT 109.580 155.970 112.110 156.110 ;
        RECT 101.685 155.770 101.975 155.815 ;
        RECT 101.300 155.630 101.975 155.770 ;
        RECT 94.325 155.585 94.615 155.630 ;
        RECT 83.270 155.430 83.590 155.490 ;
        RECT 85.585 155.430 85.875 155.475 ;
        RECT 86.950 155.430 87.270 155.490 ;
        RECT 92.560 155.430 92.700 155.585 ;
        RECT 96.610 155.570 96.930 155.630 ;
        RECT 101.685 155.585 101.975 155.630 ;
        RECT 107.650 155.770 107.970 155.830 ;
        RECT 109.580 155.815 109.720 155.970 ;
        RECT 111.790 155.910 112.110 155.970 ;
        RECT 115.945 156.110 116.235 156.155 ;
        RECT 119.100 156.110 119.390 156.155 ;
        RECT 122.360 156.110 122.650 156.155 ;
        RECT 115.945 155.970 122.650 156.110 ;
        RECT 115.945 155.925 116.235 155.970 ;
        RECT 119.100 155.925 119.390 155.970 ;
        RECT 122.360 155.925 122.650 155.970 ;
        RECT 123.280 156.110 123.570 156.155 ;
        RECT 125.140 156.110 125.430 156.155 ;
        RECT 123.280 155.970 125.430 156.110 ;
        RECT 123.280 155.925 123.570 155.970 ;
        RECT 125.140 155.925 125.430 155.970 ;
        RECT 108.125 155.770 108.415 155.815 ;
        RECT 107.650 155.630 108.415 155.770 ;
        RECT 107.650 155.570 107.970 155.630 ;
        RECT 108.125 155.585 108.415 155.630 ;
        RECT 109.505 155.585 109.795 155.815 ;
        RECT 111.345 155.770 111.635 155.815 ;
        RECT 113.170 155.770 113.490 155.830 ;
        RECT 111.345 155.630 113.490 155.770 ;
        RECT 111.345 155.585 111.635 155.630 ;
        RECT 113.170 155.570 113.490 155.630 ;
        RECT 115.485 155.585 115.775 155.815 ;
        RECT 120.960 155.770 121.250 155.815 ;
        RECT 123.280 155.770 123.495 155.925 ;
        RECT 120.960 155.630 123.495 155.770 ;
        RECT 120.960 155.585 121.250 155.630 ;
        RECT 98.005 155.430 98.295 155.475 ;
        RECT 103.510 155.430 103.830 155.490 ;
        RECT 81.520 155.290 83.590 155.430 ;
        RECT 79.130 155.230 79.450 155.290 ;
        RECT 83.270 155.230 83.590 155.290 ;
        RECT 84.740 155.290 87.270 155.430 ;
        RECT 83.730 155.090 84.050 155.150 ;
        RECT 77.840 154.950 84.050 155.090 ;
        RECT 72.245 154.905 72.535 154.950 ;
        RECT 77.290 154.890 77.610 154.950 ;
        RECT 83.730 154.890 84.050 154.950 ;
        RECT 34.510 154.550 34.830 154.810 ;
        RECT 38.650 154.550 38.970 154.810 ;
        RECT 41.870 154.750 42.190 154.810 ;
        RECT 45.565 154.750 45.855 154.795 ;
        RECT 41.870 154.610 45.855 154.750 ;
        RECT 41.870 154.550 42.190 154.610 ;
        RECT 45.565 154.565 45.855 154.610 ;
        RECT 47.865 154.750 48.155 154.795 ;
        RECT 49.690 154.750 50.010 154.810 ;
        RECT 47.865 154.610 50.010 154.750 ;
        RECT 47.865 154.565 48.155 154.610 ;
        RECT 49.690 154.550 50.010 154.610 ;
        RECT 60.270 154.750 60.590 154.810 ;
        RECT 62.125 154.750 62.415 154.795 ;
        RECT 60.270 154.610 62.415 154.750 ;
        RECT 60.270 154.550 60.590 154.610 ;
        RECT 62.125 154.565 62.415 154.610 ;
        RECT 70.850 154.750 71.170 154.810 ;
        RECT 73.165 154.750 73.455 154.795 ;
        RECT 70.850 154.610 73.455 154.750 ;
        RECT 70.850 154.550 71.170 154.610 ;
        RECT 73.165 154.565 73.455 154.610 ;
        RECT 80.065 154.750 80.355 154.795 ;
        RECT 84.740 154.750 84.880 155.290 ;
        RECT 85.585 155.245 85.875 155.290 ;
        RECT 86.950 155.230 87.270 155.290 ;
        RECT 88.420 155.290 92.700 155.430 ;
        RECT 97.160 155.290 103.830 155.430 ;
        RECT 88.420 155.135 88.560 155.290 ;
        RECT 88.345 154.905 88.635 155.135 ;
        RECT 97.160 155.090 97.300 155.290 ;
        RECT 98.005 155.245 98.295 155.290 ;
        RECT 103.510 155.230 103.830 155.290 ;
        RECT 109.045 155.430 109.335 155.475 ;
        RECT 109.950 155.430 110.270 155.490 ;
        RECT 109.045 155.290 110.270 155.430 ;
        RECT 109.045 155.245 109.335 155.290 ;
        RECT 109.950 155.230 110.270 155.290 ;
        RECT 90.260 154.950 97.300 155.090 ;
        RECT 97.530 155.090 97.850 155.150 ;
        RECT 115.560 155.090 115.700 155.585 ;
        RECT 124.210 155.570 124.530 155.830 ;
        RECT 126.050 155.230 126.370 155.490 ;
        RECT 116.390 155.090 116.710 155.150 ;
        RECT 97.530 154.950 116.710 155.090 ;
        RECT 80.065 154.610 84.880 154.750 ;
        RECT 86.950 154.750 87.270 154.810 ;
        RECT 90.260 154.750 90.400 154.950 ;
        RECT 97.530 154.890 97.850 154.950 ;
        RECT 116.390 154.890 116.710 154.950 ;
        RECT 117.095 155.090 117.385 155.135 ;
        RECT 118.690 155.090 119.010 155.150 ;
        RECT 117.095 154.950 119.010 155.090 ;
        RECT 117.095 154.905 117.385 154.950 ;
        RECT 118.690 154.890 119.010 154.950 ;
        RECT 120.960 155.090 121.250 155.135 ;
        RECT 123.740 155.090 124.030 155.135 ;
        RECT 125.600 155.090 125.890 155.135 ;
        RECT 120.960 154.950 125.890 155.090 ;
        RECT 120.960 154.905 121.250 154.950 ;
        RECT 123.740 154.905 124.030 154.950 ;
        RECT 125.600 154.905 125.890 154.950 ;
        RECT 86.950 154.610 90.400 154.750 ;
        RECT 90.630 154.750 90.950 154.810 ;
        RECT 91.105 154.750 91.395 154.795 ;
        RECT 90.630 154.610 91.395 154.750 ;
        RECT 80.065 154.565 80.355 154.610 ;
        RECT 86.950 154.550 87.270 154.610 ;
        RECT 90.630 154.550 90.950 154.610 ;
        RECT 91.105 154.565 91.395 154.610 ;
        RECT 106.270 154.750 106.590 154.810 ;
        RECT 108.125 154.750 108.415 154.795 ;
        RECT 106.270 154.610 108.415 154.750 ;
        RECT 106.270 154.550 106.590 154.610 ;
        RECT 108.125 154.565 108.415 154.610 ;
        RECT 110.425 154.750 110.715 154.795 ;
        RECT 111.790 154.750 112.110 154.810 ;
        RECT 110.425 154.610 112.110 154.750 ;
        RECT 110.425 154.565 110.715 154.610 ;
        RECT 111.790 154.550 112.110 154.610 ;
        RECT 29.840 153.930 127.820 154.410 ;
        RECT 43.250 153.730 43.570 153.790 ;
        RECT 44.645 153.730 44.935 153.775 ;
        RECT 43.250 153.590 44.935 153.730 ;
        RECT 43.250 153.530 43.570 153.590 ;
        RECT 44.645 153.545 44.935 153.590 ;
        RECT 46.470 153.530 46.790 153.790 ;
        RECT 48.785 153.730 49.075 153.775 ;
        RECT 49.230 153.730 49.550 153.790 ;
        RECT 48.785 153.590 49.550 153.730 ;
        RECT 48.785 153.545 49.075 153.590 ;
        RECT 49.230 153.530 49.550 153.590 ;
        RECT 49.705 153.730 49.995 153.775 ;
        RECT 50.610 153.730 50.930 153.790 ;
        RECT 49.705 153.590 50.930 153.730 ;
        RECT 49.705 153.545 49.995 153.590 ;
        RECT 50.610 153.530 50.930 153.590 ;
        RECT 51.530 153.730 51.850 153.790 ;
        RECT 56.835 153.730 57.125 153.775 ;
        RECT 58.430 153.730 58.750 153.790 ;
        RECT 66.710 153.730 67.030 153.790 ;
        RECT 51.530 153.590 56.360 153.730 ;
        RECT 51.530 153.530 51.850 153.590 ;
        RECT 35.400 153.390 35.690 153.435 ;
        RECT 38.180 153.390 38.470 153.435 ;
        RECT 40.040 153.390 40.330 153.435 ;
        RECT 52.465 153.390 52.755 153.435 ;
        RECT 53.830 153.390 54.150 153.450 ;
        RECT 35.400 153.250 40.330 153.390 ;
        RECT 35.400 153.205 35.690 153.250 ;
        RECT 38.180 153.205 38.470 153.250 ;
        RECT 40.040 153.205 40.330 153.250 ;
        RECT 41.960 153.250 46.700 153.390 ;
        RECT 38.650 152.850 38.970 153.110 ;
        RECT 41.960 153.050 42.100 153.250 ;
        RECT 40.120 152.910 42.100 153.050 ;
        RECT 42.330 153.050 42.650 153.110 ;
        RECT 45.090 153.050 45.410 153.110 ;
        RECT 46.025 153.050 46.315 153.095 ;
        RECT 42.330 152.910 43.940 153.050 ;
        RECT 35.400 152.710 35.690 152.755 ;
        RECT 35.400 152.570 37.935 152.710 ;
        RECT 35.400 152.525 35.690 152.570 ;
        RECT 33.540 152.370 33.830 152.415 ;
        RECT 34.510 152.370 34.830 152.430 ;
        RECT 37.720 152.415 37.935 152.570 ;
        RECT 36.800 152.370 37.090 152.415 ;
        RECT 33.540 152.230 37.090 152.370 ;
        RECT 33.540 152.185 33.830 152.230 ;
        RECT 34.510 152.170 34.830 152.230 ;
        RECT 36.800 152.185 37.090 152.230 ;
        RECT 37.720 152.370 38.010 152.415 ;
        RECT 39.580 152.370 39.870 152.415 ;
        RECT 37.720 152.230 39.870 152.370 ;
        RECT 37.720 152.185 38.010 152.230 ;
        RECT 39.580 152.185 39.870 152.230 ;
        RECT 31.535 152.030 31.825 152.075 ;
        RECT 34.970 152.030 35.290 152.090 ;
        RECT 40.120 152.030 40.260 152.910 ;
        RECT 42.330 152.850 42.650 152.910 ;
        RECT 40.505 152.710 40.795 152.755 ;
        RECT 42.790 152.710 43.110 152.770 ;
        RECT 40.505 152.570 43.110 152.710 ;
        RECT 40.505 152.525 40.795 152.570 ;
        RECT 42.790 152.510 43.110 152.570 ;
        RECT 43.265 152.525 43.555 152.755 ;
        RECT 42.330 152.370 42.650 152.430 ;
        RECT 43.340 152.370 43.480 152.525 ;
        RECT 42.330 152.230 43.480 152.370 ;
        RECT 43.800 152.370 43.940 152.910 ;
        RECT 45.090 152.910 46.315 153.050 ;
        RECT 46.560 153.050 46.700 153.250 ;
        RECT 52.465 153.250 54.150 153.390 ;
        RECT 52.465 153.205 52.755 153.250 ;
        RECT 53.830 153.190 54.150 153.250 ;
        RECT 50.625 153.050 50.915 153.095 ;
        RECT 46.560 152.910 50.915 153.050 ;
        RECT 45.090 152.850 45.410 152.910 ;
        RECT 46.025 152.865 46.315 152.910 ;
        RECT 50.625 152.865 50.915 152.910 ;
        RECT 52.925 153.050 53.215 153.095 ;
        RECT 55.670 153.050 55.990 153.110 ;
        RECT 52.925 152.910 53.600 153.050 ;
        RECT 52.925 152.865 53.215 152.910 ;
        RECT 45.550 152.510 45.870 152.770 ;
        RECT 48.325 152.710 48.615 152.755 ;
        RECT 46.100 152.570 48.615 152.710 ;
        RECT 46.100 152.370 46.240 152.570 ;
        RECT 48.325 152.525 48.615 152.570 ;
        RECT 48.785 152.710 49.075 152.755 ;
        RECT 50.150 152.710 50.470 152.770 ;
        RECT 48.785 152.570 50.470 152.710 ;
        RECT 48.785 152.525 49.075 152.570 ;
        RECT 50.150 152.510 50.470 152.570 ;
        RECT 51.070 152.710 51.390 152.770 ;
        RECT 51.545 152.710 51.835 152.755 ;
        RECT 51.070 152.570 51.835 152.710 ;
        RECT 51.070 152.510 51.390 152.570 ;
        RECT 51.545 152.525 51.835 152.570 ;
        RECT 43.800 152.230 46.240 152.370 ;
        RECT 42.330 152.170 42.650 152.230 ;
        RECT 46.945 152.185 47.235 152.415 ;
        RECT 47.405 152.370 47.695 152.415 ;
        RECT 52.910 152.370 53.230 152.430 ;
        RECT 47.405 152.230 53.230 152.370 ;
        RECT 47.405 152.185 47.695 152.230 ;
        RECT 31.535 151.890 40.260 152.030 ;
        RECT 44.185 152.030 44.475 152.075 ;
        RECT 45.090 152.030 45.410 152.090 ;
        RECT 44.185 151.890 45.410 152.030 ;
        RECT 47.020 152.030 47.160 152.185 ;
        RECT 52.910 152.170 53.230 152.230 ;
        RECT 53.460 152.030 53.600 152.910 ;
        RECT 54.380 152.910 55.990 153.050 ;
        RECT 54.380 152.755 54.520 152.910 ;
        RECT 55.670 152.850 55.990 152.910 ;
        RECT 56.220 152.770 56.360 153.590 ;
        RECT 56.835 153.590 67.030 153.730 ;
        RECT 56.835 153.545 57.125 153.590 ;
        RECT 54.305 152.525 54.595 152.755 ;
        RECT 54.750 152.510 55.070 152.770 ;
        RECT 55.225 152.525 55.515 152.755 ;
        RECT 55.300 152.370 55.440 152.525 ;
        RECT 56.130 152.510 56.450 152.770 ;
        RECT 56.910 152.370 57.050 153.545 ;
        RECT 58.430 153.530 58.750 153.590 ;
        RECT 66.710 153.530 67.030 153.590 ;
        RECT 80.050 153.530 80.370 153.790 ;
        RECT 107.650 153.530 107.970 153.790 ;
        RECT 115.470 153.730 115.790 153.790 ;
        RECT 117.770 153.730 118.090 153.790 ;
        RECT 109.120 153.590 118.460 153.730 ;
        RECT 60.700 153.390 60.990 153.435 ;
        RECT 63.480 153.390 63.770 153.435 ;
        RECT 65.340 153.390 65.630 153.435 ;
        RECT 60.700 153.250 65.630 153.390 ;
        RECT 60.700 153.205 60.990 153.250 ;
        RECT 63.480 153.205 63.770 153.250 ;
        RECT 65.340 153.205 65.630 153.250 ;
        RECT 69.585 153.390 69.875 153.435 ;
        RECT 72.705 153.390 72.995 153.435 ;
        RECT 74.595 153.390 74.885 153.435 ;
        RECT 69.585 153.250 74.885 153.390 ;
        RECT 69.585 153.205 69.875 153.250 ;
        RECT 72.705 153.205 72.995 153.250 ;
        RECT 74.595 153.205 74.885 153.250 ;
        RECT 76.385 153.205 76.675 153.435 ;
        RECT 78.685 153.390 78.975 153.435 ;
        RECT 79.130 153.390 79.450 153.450 ;
        RECT 83.270 153.390 83.590 153.450 ;
        RECT 78.685 153.250 83.590 153.390 ;
        RECT 78.685 153.205 78.975 153.250 ;
        RECT 61.190 153.050 61.510 153.110 ;
        RECT 61.190 152.910 63.720 153.050 ;
        RECT 61.190 152.850 61.510 152.910 ;
        RECT 60.700 152.710 60.990 152.755 ;
        RECT 63.580 152.710 63.720 152.910 ;
        RECT 63.950 152.850 64.270 153.110 ;
        RECT 73.610 153.050 73.930 153.110 ;
        RECT 65.880 152.910 73.930 153.050 ;
        RECT 65.880 152.755 66.020 152.910 ;
        RECT 73.610 152.850 73.930 152.910 ;
        RECT 74.085 153.050 74.375 153.095 ;
        RECT 76.460 153.050 76.600 153.205 ;
        RECT 79.130 153.190 79.450 153.250 ;
        RECT 83.270 153.190 83.590 153.250 ;
        RECT 90.140 153.390 90.430 153.435 ;
        RECT 92.920 153.390 93.210 153.435 ;
        RECT 94.780 153.390 95.070 153.435 ;
        RECT 90.140 153.250 95.070 153.390 ;
        RECT 90.140 153.205 90.430 153.250 ;
        RECT 92.920 153.205 93.210 153.250 ;
        RECT 94.780 153.205 95.070 153.250 ;
        RECT 103.510 153.390 103.830 153.450 ;
        RECT 109.120 153.390 109.260 153.590 ;
        RECT 115.470 153.530 115.790 153.590 ;
        RECT 117.770 153.530 118.090 153.590 ;
        RECT 112.710 153.390 113.030 153.450 ;
        RECT 103.510 153.250 109.260 153.390 ;
        RECT 109.580 153.250 113.030 153.390 ;
        RECT 103.510 153.190 103.830 153.250 ;
        RECT 74.085 152.910 76.600 153.050 ;
        RECT 74.085 152.865 74.375 152.910 ;
        RECT 80.510 152.850 80.830 153.110 ;
        RECT 82.810 153.050 83.130 153.110 ;
        RECT 86.275 153.050 86.565 153.095 ;
        RECT 82.810 152.910 84.420 153.050 ;
        RECT 82.810 152.850 83.130 152.910 ;
        RECT 65.805 152.710 66.095 152.755 ;
        RECT 60.700 152.570 63.235 152.710 ;
        RECT 63.580 152.570 66.095 152.710 ;
        RECT 60.700 152.525 60.990 152.570 ;
        RECT 55.300 152.230 57.050 152.370 ;
        RECT 58.840 152.370 59.130 152.415 ;
        RECT 60.270 152.370 60.590 152.430 ;
        RECT 63.020 152.415 63.235 152.570 ;
        RECT 65.805 152.525 66.095 152.570 ;
        RECT 68.505 152.415 68.795 152.730 ;
        RECT 69.585 152.710 69.875 152.755 ;
        RECT 73.165 152.710 73.455 152.755 ;
        RECT 75.000 152.710 75.290 152.755 ;
        RECT 69.585 152.570 75.290 152.710 ;
        RECT 69.585 152.525 69.875 152.570 ;
        RECT 73.165 152.525 73.455 152.570 ;
        RECT 75.000 152.525 75.290 152.570 ;
        RECT 75.465 152.710 75.755 152.755 ;
        RECT 75.910 152.710 76.230 152.770 ;
        RECT 75.465 152.570 76.230 152.710 ;
        RECT 75.465 152.525 75.755 152.570 ;
        RECT 62.100 152.370 62.390 152.415 ;
        RECT 58.840 152.230 62.390 152.370 ;
        RECT 58.840 152.185 59.130 152.230 ;
        RECT 60.270 152.170 60.590 152.230 ;
        RECT 62.100 152.185 62.390 152.230 ;
        RECT 63.020 152.370 63.310 152.415 ;
        RECT 64.880 152.370 65.170 152.415 ;
        RECT 63.020 152.230 65.170 152.370 ;
        RECT 63.020 152.185 63.310 152.230 ;
        RECT 64.880 152.185 65.170 152.230 ;
        RECT 68.205 152.370 68.795 152.415 ;
        RECT 70.850 152.370 71.170 152.430 ;
        RECT 71.445 152.370 72.095 152.415 ;
        RECT 68.205 152.230 72.095 152.370 ;
        RECT 68.205 152.185 68.495 152.230 ;
        RECT 70.850 152.170 71.170 152.230 ;
        RECT 71.445 152.185 72.095 152.230 ;
        RECT 73.610 152.370 73.930 152.430 ;
        RECT 75.540 152.370 75.680 152.525 ;
        RECT 75.910 152.510 76.230 152.570 ;
        RECT 77.290 152.510 77.610 152.770 ;
        RECT 77.765 152.525 78.055 152.755 ;
        RECT 73.610 152.230 75.680 152.370 ;
        RECT 76.370 152.370 76.690 152.430 ;
        RECT 77.840 152.370 77.980 152.525 ;
        RECT 80.970 152.510 81.290 152.770 ;
        RECT 83.730 152.510 84.050 152.770 ;
        RECT 84.280 152.755 84.420 152.910 ;
        RECT 85.200 152.910 86.565 153.050 ;
        RECT 85.200 152.770 85.340 152.910 ;
        RECT 86.275 152.865 86.565 152.910 ;
        RECT 98.910 153.050 99.230 153.110 ;
        RECT 109.580 153.050 109.720 153.250 ;
        RECT 112.710 153.190 113.030 153.250 ;
        RECT 118.320 153.095 118.460 153.590 ;
        RECT 98.910 152.910 109.720 153.050 ;
        RECT 98.910 152.850 99.230 152.910 ;
        RECT 84.205 152.525 84.495 152.755 ;
        RECT 84.665 152.710 84.955 152.755 ;
        RECT 85.110 152.710 85.430 152.770 ;
        RECT 84.665 152.570 85.430 152.710 ;
        RECT 84.665 152.525 84.955 152.570 ;
        RECT 85.110 152.510 85.430 152.570 ;
        RECT 85.585 152.525 85.875 152.755 ;
        RECT 90.140 152.710 90.430 152.755 ;
        RECT 90.140 152.570 92.675 152.710 ;
        RECT 90.140 152.525 90.430 152.570 ;
        RECT 76.370 152.230 77.980 152.370 ;
        RECT 79.605 152.370 79.895 152.415 ;
        RECT 82.365 152.370 82.655 152.415 ;
        RECT 79.605 152.230 82.655 152.370 ;
        RECT 73.610 152.170 73.930 152.230 ;
        RECT 76.370 152.170 76.690 152.230 ;
        RECT 79.605 152.185 79.895 152.230 ;
        RECT 82.365 152.185 82.655 152.230 ;
        RECT 83.270 152.370 83.590 152.430 ;
        RECT 85.660 152.370 85.800 152.525 ;
        RECT 83.270 152.230 85.800 152.370 ;
        RECT 88.280 152.370 88.570 152.415 ;
        RECT 90.630 152.370 90.950 152.430 ;
        RECT 92.460 152.415 92.675 152.570 ;
        RECT 93.390 152.510 93.710 152.770 ;
        RECT 95.245 152.710 95.535 152.755 ;
        RECT 95.690 152.710 96.010 152.770 ;
        RECT 95.245 152.570 96.010 152.710 ;
        RECT 95.245 152.525 95.535 152.570 ;
        RECT 95.690 152.510 96.010 152.570 ;
        RECT 99.370 152.510 99.690 152.770 ;
        RECT 99.920 152.755 100.060 152.910 ;
        RECT 109.580 152.770 109.720 152.910 ;
        RECT 110.040 152.910 118.000 153.050 ;
        RECT 99.845 152.525 100.135 152.755 ;
        RECT 100.305 152.525 100.595 152.755 ;
        RECT 101.225 152.710 101.515 152.755 ;
        RECT 105.810 152.710 106.130 152.770 ;
        RECT 101.225 152.570 106.130 152.710 ;
        RECT 101.225 152.525 101.515 152.570 ;
        RECT 91.540 152.370 91.830 152.415 ;
        RECT 88.280 152.230 91.830 152.370 ;
        RECT 83.270 152.170 83.590 152.230 ;
        RECT 88.280 152.185 88.570 152.230 ;
        RECT 90.630 152.170 90.950 152.230 ;
        RECT 91.540 152.185 91.830 152.230 ;
        RECT 92.460 152.370 92.750 152.415 ;
        RECT 94.320 152.370 94.610 152.415 ;
        RECT 92.460 152.230 94.610 152.370 ;
        RECT 92.460 152.185 92.750 152.230 ;
        RECT 94.320 152.185 94.610 152.230 ;
        RECT 98.450 152.370 98.770 152.430 ;
        RECT 100.380 152.370 100.520 152.525 ;
        RECT 105.810 152.510 106.130 152.570 ;
        RECT 109.030 152.510 109.350 152.770 ;
        RECT 109.490 152.510 109.810 152.770 ;
        RECT 110.040 152.755 110.180 152.910 ;
        RECT 109.965 152.525 110.255 152.755 ;
        RECT 110.885 152.710 111.175 152.755 ;
        RECT 111.345 152.710 111.635 152.755 ;
        RECT 110.885 152.570 111.635 152.710 ;
        RECT 110.885 152.525 111.175 152.570 ;
        RECT 111.345 152.525 111.635 152.570 ;
        RECT 112.265 152.525 112.555 152.755 ;
        RECT 98.450 152.230 100.520 152.370 ;
        RECT 105.900 152.370 106.040 152.510 ;
        RECT 110.410 152.370 110.730 152.430 ;
        RECT 110.960 152.370 111.100 152.525 ;
        RECT 105.900 152.230 111.100 152.370 ;
        RECT 112.340 152.370 112.480 152.525 ;
        RECT 112.710 152.510 113.030 152.770 ;
        RECT 113.170 152.510 113.490 152.770 ;
        RECT 117.860 152.710 118.000 152.910 ;
        RECT 118.245 152.865 118.535 153.095 ;
        RECT 118.690 152.710 119.010 152.770 ;
        RECT 119.165 152.710 119.455 152.755 ;
        RECT 117.860 152.570 119.455 152.710 ;
        RECT 118.690 152.510 119.010 152.570 ;
        RECT 119.165 152.525 119.455 152.570 ;
        RECT 112.340 152.230 115.240 152.370 ;
        RECT 98.450 152.170 98.770 152.230 ;
        RECT 110.410 152.170 110.730 152.230 ;
        RECT 47.020 151.890 53.600 152.030 ;
        RECT 66.725 152.030 67.015 152.075 ;
        RECT 67.170 152.030 67.490 152.090 ;
        RECT 66.725 151.890 67.490 152.030 ;
        RECT 31.535 151.845 31.825 151.890 ;
        RECT 34.970 151.830 35.290 151.890 ;
        RECT 44.185 151.845 44.475 151.890 ;
        RECT 45.090 151.830 45.410 151.890 ;
        RECT 66.725 151.845 67.015 151.890 ;
        RECT 67.170 151.830 67.490 151.890 ;
        RECT 81.905 152.030 82.195 152.075 ;
        RECT 84.650 152.030 84.970 152.090 ;
        RECT 81.905 151.890 84.970 152.030 ;
        RECT 81.905 151.845 82.195 151.890 ;
        RECT 84.650 151.830 84.970 151.890 ;
        RECT 97.990 151.830 98.310 152.090 ;
        RECT 99.370 152.030 99.690 152.090 ;
        RECT 109.030 152.030 109.350 152.090 ;
        RECT 113.170 152.030 113.490 152.090 ;
        RECT 99.370 151.890 113.490 152.030 ;
        RECT 99.370 151.830 99.690 151.890 ;
        RECT 109.030 151.830 109.350 151.890 ;
        RECT 113.170 151.830 113.490 151.890 ;
        RECT 114.550 151.830 114.870 152.090 ;
        RECT 115.100 152.030 115.240 152.230 ;
        RECT 116.850 152.030 117.170 152.090 ;
        RECT 118.705 152.030 118.995 152.075 ;
        RECT 115.100 151.890 118.995 152.030 ;
        RECT 116.850 151.830 117.170 151.890 ;
        RECT 118.705 151.845 118.995 151.890 ;
        RECT 121.005 152.030 121.295 152.075 ;
        RECT 121.450 152.030 121.770 152.090 ;
        RECT 121.005 151.890 121.770 152.030 ;
        RECT 121.005 151.845 121.295 151.890 ;
        RECT 121.450 151.830 121.770 151.890 ;
        RECT 29.840 151.210 127.820 151.690 ;
        RECT 34.970 150.810 35.290 151.070 ;
        RECT 36.810 150.810 37.130 151.070 ;
        RECT 47.405 151.010 47.695 151.055 ;
        RECT 49.230 151.010 49.550 151.070 ;
        RECT 47.405 150.870 49.550 151.010 ;
        RECT 47.405 150.825 47.695 150.870 ;
        RECT 49.230 150.810 49.550 150.870 ;
        RECT 49.690 150.810 50.010 151.070 ;
        RECT 52.910 150.810 53.230 151.070 ;
        RECT 53.830 151.010 54.150 151.070 ;
        RECT 55.210 151.010 55.530 151.070 ;
        RECT 59.365 151.010 59.655 151.055 ;
        RECT 53.830 150.870 59.655 151.010 ;
        RECT 53.830 150.810 54.150 150.870 ;
        RECT 55.210 150.810 55.530 150.870 ;
        RECT 59.365 150.825 59.655 150.870 ;
        RECT 61.205 150.825 61.495 151.055 ;
        RECT 70.850 151.010 71.170 151.070 ;
        RECT 79.130 151.010 79.450 151.070 ;
        RECT 68.180 150.870 79.450 151.010 ;
        RECT 32.225 150.670 32.515 150.715 ;
        RECT 39.980 150.670 40.270 150.715 ;
        RECT 43.240 150.670 43.530 150.715 ;
        RECT 32.225 150.530 43.530 150.670 ;
        RECT 32.225 150.485 32.515 150.530 ;
        RECT 39.980 150.485 40.270 150.530 ;
        RECT 43.240 150.485 43.530 150.530 ;
        RECT 44.160 150.670 44.450 150.715 ;
        RECT 46.020 150.670 46.310 150.715 ;
        RECT 55.670 150.670 55.990 150.730 ;
        RECT 44.160 150.530 46.310 150.670 ;
        RECT 44.160 150.485 44.450 150.530 ;
        RECT 46.020 150.485 46.310 150.530 ;
        RECT 48.400 150.530 50.840 150.670 ;
        RECT 31.290 150.330 31.610 150.390 ;
        RECT 32.685 150.330 32.975 150.375 ;
        RECT 31.290 150.190 32.975 150.330 ;
        RECT 31.290 150.130 31.610 150.190 ;
        RECT 32.685 150.145 32.975 150.190 ;
        RECT 41.840 150.330 42.130 150.375 ;
        RECT 44.160 150.330 44.375 150.485 ;
        RECT 41.840 150.190 44.375 150.330 ;
        RECT 41.840 150.145 42.130 150.190 ;
        RECT 45.090 150.130 45.410 150.390 ;
        RECT 48.400 150.375 48.540 150.530 ;
        RECT 50.700 150.390 50.840 150.530 ;
        RECT 54.380 150.530 55.990 150.670 ;
        RECT 48.325 150.145 48.615 150.375 ;
        RECT 48.770 150.130 49.090 150.390 ;
        RECT 50.610 150.130 50.930 150.390 ;
        RECT 51.070 150.130 51.390 150.390 ;
        RECT 54.380 150.375 54.520 150.530 ;
        RECT 55.670 150.470 55.990 150.530 ;
        RECT 58.905 150.670 59.195 150.715 ;
        RECT 60.730 150.670 61.050 150.730 ;
        RECT 58.905 150.530 61.050 150.670 ;
        RECT 58.905 150.485 59.195 150.530 ;
        RECT 60.730 150.470 61.050 150.530 ;
        RECT 54.305 150.145 54.595 150.375 ;
        RECT 54.750 150.130 55.070 150.390 ;
        RECT 55.210 150.130 55.530 150.390 ;
        RECT 56.130 150.130 56.450 150.390 ;
        RECT 61.280 150.330 61.420 150.825 ;
        RECT 62.585 150.330 62.875 150.375 ;
        RECT 61.280 150.190 62.875 150.330 ;
        RECT 62.585 150.145 62.875 150.190 ;
        RECT 66.265 150.145 66.555 150.375 ;
        RECT 66.725 150.145 67.015 150.375 ;
        RECT 34.050 149.790 34.370 150.050 ;
        RECT 34.525 149.805 34.815 150.035 ;
        RECT 42.790 149.990 43.110 150.050 ;
        RECT 46.945 149.990 47.235 150.035 ;
        RECT 58.445 149.990 58.735 150.035 ;
        RECT 65.790 149.990 66.110 150.050 ;
        RECT 42.790 149.850 56.360 149.990 ;
        RECT 34.600 149.310 34.740 149.805 ;
        RECT 42.790 149.790 43.110 149.850 ;
        RECT 46.945 149.805 47.235 149.850 ;
        RECT 56.220 149.710 56.360 149.850 ;
        RECT 58.445 149.850 66.110 149.990 ;
        RECT 58.445 149.805 58.735 149.850 ;
        RECT 65.790 149.790 66.110 149.850 ;
        RECT 41.840 149.650 42.130 149.695 ;
        RECT 44.620 149.650 44.910 149.695 ;
        RECT 46.480 149.650 46.770 149.695 ;
        RECT 41.840 149.510 46.770 149.650 ;
        RECT 41.840 149.465 42.130 149.510 ;
        RECT 44.620 149.465 44.910 149.510 ;
        RECT 46.480 149.465 46.770 149.510 ;
        RECT 56.130 149.450 56.450 149.710 ;
        RECT 59.350 149.650 59.670 149.710 ;
        RECT 61.665 149.650 61.955 149.695 ;
        RECT 59.350 149.510 61.955 149.650 ;
        RECT 66.340 149.650 66.480 150.145 ;
        RECT 66.800 149.990 66.940 150.145 ;
        RECT 67.170 150.130 67.490 150.390 ;
        RECT 68.180 150.375 68.320 150.870 ;
        RECT 70.850 150.810 71.170 150.870 ;
        RECT 79.130 150.810 79.450 150.870 ;
        RECT 79.605 150.825 79.895 151.055 ;
        RECT 85.110 151.010 85.430 151.070 ;
        RECT 86.045 151.010 86.335 151.055 ;
        RECT 85.110 150.870 86.335 151.010 ;
        RECT 69.025 150.670 69.315 150.715 ;
        RECT 72.180 150.670 72.470 150.715 ;
        RECT 75.440 150.670 75.730 150.715 ;
        RECT 69.025 150.530 75.730 150.670 ;
        RECT 69.025 150.485 69.315 150.530 ;
        RECT 72.180 150.485 72.470 150.530 ;
        RECT 75.440 150.485 75.730 150.530 ;
        RECT 76.360 150.670 76.650 150.715 ;
        RECT 78.220 150.670 78.510 150.715 ;
        RECT 76.360 150.530 78.510 150.670 ;
        RECT 76.360 150.485 76.650 150.530 ;
        RECT 78.220 150.485 78.510 150.530 ;
        RECT 68.105 150.145 68.395 150.375 ;
        RECT 68.565 150.330 68.855 150.375 ;
        RECT 70.390 150.330 70.710 150.390 ;
        RECT 68.565 150.190 70.710 150.330 ;
        RECT 68.565 150.145 68.855 150.190 ;
        RECT 70.390 150.130 70.710 150.190 ;
        RECT 74.040 150.330 74.330 150.375 ;
        RECT 76.360 150.330 76.575 150.485 ;
        RECT 74.040 150.190 76.575 150.330 ;
        RECT 77.305 150.330 77.595 150.375 ;
        RECT 79.680 150.330 79.820 150.825 ;
        RECT 85.110 150.810 85.430 150.870 ;
        RECT 86.045 150.825 86.335 150.870 ;
        RECT 88.345 150.825 88.635 151.055 ;
        RECT 92.485 151.010 92.775 151.055 ;
        RECT 93.390 151.010 93.710 151.070 ;
        RECT 92.485 150.870 93.710 151.010 ;
        RECT 92.485 150.825 92.775 150.870 ;
        RECT 77.305 150.190 79.820 150.330 ;
        RECT 74.040 150.145 74.330 150.190 ;
        RECT 77.305 150.145 77.595 150.190 ;
        RECT 80.510 150.130 80.830 150.390 ;
        RECT 86.030 150.330 86.350 150.390 ;
        RECT 86.505 150.330 86.795 150.375 ;
        RECT 86.030 150.190 86.795 150.330 ;
        RECT 88.420 150.330 88.560 150.825 ;
        RECT 93.390 150.810 93.710 150.870 ;
        RECT 108.110 151.010 108.430 151.070 ;
        RECT 112.250 151.010 112.570 151.070 ;
        RECT 108.110 150.870 112.570 151.010 ;
        RECT 108.110 150.810 108.430 150.870 ;
        RECT 112.250 150.810 112.570 150.870 ;
        RECT 99.370 150.715 99.690 150.730 ;
        RECT 99.320 150.670 99.690 150.715 ;
        RECT 102.580 150.670 102.870 150.715 ;
        RECT 99.320 150.530 102.870 150.670 ;
        RECT 99.320 150.485 99.690 150.530 ;
        RECT 102.580 150.485 102.870 150.530 ;
        RECT 103.500 150.670 103.790 150.715 ;
        RECT 105.360 150.670 105.650 150.715 ;
        RECT 112.710 150.670 113.030 150.730 ;
        RECT 103.500 150.530 105.650 150.670 ;
        RECT 103.500 150.485 103.790 150.530 ;
        RECT 105.360 150.485 105.650 150.530 ;
        RECT 110.500 150.530 113.030 150.670 ;
        RECT 99.370 150.470 99.690 150.485 ;
        RECT 91.565 150.330 91.855 150.375 ;
        RECT 88.420 150.190 91.855 150.330 ;
        RECT 86.030 150.130 86.350 150.190 ;
        RECT 86.505 150.145 86.795 150.190 ;
        RECT 91.565 150.145 91.855 150.190 ;
        RECT 101.180 150.330 101.470 150.375 ;
        RECT 103.500 150.330 103.715 150.485 ;
        RECT 101.180 150.190 103.715 150.330 ;
        RECT 101.180 150.145 101.470 150.190 ;
        RECT 104.430 150.130 104.750 150.390 ;
        RECT 109.030 150.330 109.350 150.390 ;
        RECT 110.500 150.375 110.640 150.530 ;
        RECT 112.710 150.470 113.030 150.530 ;
        RECT 113.645 150.670 113.935 150.715 ;
        RECT 119.100 150.670 119.390 150.715 ;
        RECT 122.360 150.670 122.650 150.715 ;
        RECT 113.645 150.530 122.650 150.670 ;
        RECT 113.645 150.485 113.935 150.530 ;
        RECT 119.100 150.485 119.390 150.530 ;
        RECT 122.360 150.485 122.650 150.530 ;
        RECT 123.280 150.670 123.570 150.715 ;
        RECT 125.140 150.670 125.430 150.715 ;
        RECT 123.280 150.530 125.430 150.670 ;
        RECT 123.280 150.485 123.570 150.530 ;
        RECT 125.140 150.485 125.430 150.530 ;
        RECT 109.505 150.330 109.795 150.375 ;
        RECT 109.030 150.190 109.795 150.330 ;
        RECT 109.030 150.130 109.350 150.190 ;
        RECT 109.505 150.145 109.795 150.190 ;
        RECT 109.965 150.145 110.255 150.375 ;
        RECT 110.425 150.145 110.715 150.375 ;
        RECT 111.345 150.145 111.635 150.375 ;
        RECT 113.185 150.330 113.475 150.375 ;
        RECT 115.485 150.330 115.775 150.375 ;
        RECT 116.390 150.330 116.710 150.390 ;
        RECT 113.185 150.190 116.710 150.330 ;
        RECT 113.185 150.145 113.475 150.190 ;
        RECT 115.485 150.145 115.775 150.190 ;
        RECT 67.630 149.990 67.950 150.050 ;
        RECT 66.800 149.850 67.950 149.990 ;
        RECT 67.630 149.790 67.950 149.850 ;
        RECT 75.910 149.990 76.230 150.050 ;
        RECT 79.145 149.990 79.435 150.035 ;
        RECT 75.910 149.850 79.435 149.990 ;
        RECT 75.910 149.790 76.230 149.850 ;
        RECT 79.145 149.805 79.435 149.850 ;
        RECT 85.585 149.990 85.875 150.035 ;
        RECT 86.950 149.990 87.270 150.050 ;
        RECT 85.585 149.850 87.270 149.990 ;
        RECT 85.585 149.805 85.875 149.850 ;
        RECT 86.950 149.790 87.270 149.850 ;
        RECT 102.130 149.990 102.450 150.050 ;
        RECT 106.285 149.990 106.575 150.035 ;
        RECT 102.130 149.850 108.800 149.990 ;
        RECT 102.130 149.790 102.450 149.850 ;
        RECT 106.285 149.805 106.575 149.850 ;
        RECT 68.090 149.650 68.410 149.710 ;
        RECT 66.340 149.510 68.410 149.650 ;
        RECT 59.350 149.450 59.670 149.510 ;
        RECT 61.665 149.465 61.955 149.510 ;
        RECT 68.090 149.450 68.410 149.510 ;
        RECT 74.040 149.650 74.330 149.695 ;
        RECT 76.820 149.650 77.110 149.695 ;
        RECT 78.680 149.650 78.970 149.695 ;
        RECT 74.040 149.510 78.970 149.650 ;
        RECT 74.040 149.465 74.330 149.510 ;
        RECT 76.820 149.465 77.110 149.510 ;
        RECT 78.680 149.465 78.970 149.510 ;
        RECT 101.180 149.650 101.470 149.695 ;
        RECT 103.960 149.650 104.250 149.695 ;
        RECT 105.820 149.650 106.110 149.695 ;
        RECT 101.180 149.510 106.110 149.650 ;
        RECT 101.180 149.465 101.470 149.510 ;
        RECT 103.960 149.465 104.250 149.510 ;
        RECT 105.820 149.465 106.110 149.510 ;
        RECT 37.975 149.310 38.265 149.355 ;
        RECT 51.070 149.310 51.390 149.370 ;
        RECT 34.600 149.170 51.390 149.310 ;
        RECT 37.975 149.125 38.265 149.170 ;
        RECT 51.070 149.110 51.390 149.170 ;
        RECT 55.670 149.310 55.990 149.370 ;
        RECT 64.885 149.310 65.175 149.355 ;
        RECT 55.670 149.170 65.175 149.310 ;
        RECT 55.670 149.110 55.990 149.170 ;
        RECT 64.885 149.125 65.175 149.170 ;
        RECT 70.175 149.310 70.465 149.355 ;
        RECT 73.610 149.310 73.930 149.370 ;
        RECT 70.175 149.170 73.930 149.310 ;
        RECT 70.175 149.125 70.465 149.170 ;
        RECT 73.610 149.110 73.930 149.170 ;
        RECT 97.315 149.310 97.605 149.355 ;
        RECT 98.450 149.310 98.770 149.370 ;
        RECT 97.315 149.170 98.770 149.310 ;
        RECT 97.315 149.125 97.605 149.170 ;
        RECT 98.450 149.110 98.770 149.170 ;
        RECT 107.190 149.310 107.510 149.370 ;
        RECT 108.125 149.310 108.415 149.355 ;
        RECT 107.190 149.170 108.415 149.310 ;
        RECT 108.660 149.310 108.800 149.850 ;
        RECT 109.490 149.650 109.810 149.710 ;
        RECT 110.040 149.650 110.180 150.145 ;
        RECT 111.420 149.990 111.560 150.145 ;
        RECT 116.390 150.130 116.710 150.190 ;
        RECT 116.850 150.375 117.170 150.390 ;
        RECT 116.850 150.145 117.385 150.375 ;
        RECT 120.960 150.330 121.250 150.375 ;
        RECT 123.280 150.330 123.495 150.485 ;
        RECT 120.960 150.190 123.495 150.330 ;
        RECT 120.960 150.145 121.250 150.190 ;
        RECT 116.850 150.130 117.170 150.145 ;
        RECT 124.210 150.130 124.530 150.390 ;
        RECT 126.050 150.130 126.370 150.390 ;
        RECT 126.140 149.990 126.280 150.130 ;
        RECT 110.500 149.850 111.560 149.990 ;
        RECT 119.470 149.850 126.280 149.990 ;
        RECT 110.500 149.710 110.640 149.850 ;
        RECT 109.490 149.510 110.180 149.650 ;
        RECT 109.490 149.450 109.810 149.510 ;
        RECT 110.410 149.450 110.730 149.710 ;
        RECT 119.470 149.650 119.610 149.850 ;
        RECT 112.800 149.510 119.610 149.650 ;
        RECT 120.960 149.650 121.250 149.695 ;
        RECT 123.740 149.650 124.030 149.695 ;
        RECT 125.600 149.650 125.890 149.695 ;
        RECT 120.960 149.510 125.890 149.650 ;
        RECT 112.800 149.310 112.940 149.510 ;
        RECT 120.960 149.465 121.250 149.510 ;
        RECT 123.740 149.465 124.030 149.510 ;
        RECT 125.600 149.465 125.890 149.510 ;
        RECT 108.660 149.170 112.940 149.310 ;
        RECT 107.190 149.110 107.510 149.170 ;
        RECT 108.125 149.125 108.415 149.170 ;
        RECT 115.930 149.110 116.250 149.370 ;
        RECT 29.840 148.490 127.820 148.970 ;
        RECT 42.330 148.290 42.650 148.350 ;
        RECT 42.805 148.290 43.095 148.335 ;
        RECT 42.330 148.150 43.095 148.290 ;
        RECT 42.330 148.090 42.650 148.150 ;
        RECT 42.805 148.105 43.095 148.150 ;
        RECT 46.470 148.290 46.790 148.350 ;
        RECT 46.945 148.290 47.235 148.335 ;
        RECT 46.470 148.150 47.235 148.290 ;
        RECT 46.470 148.090 46.790 148.150 ;
        RECT 46.945 148.105 47.235 148.150 ;
        RECT 51.545 148.290 51.835 148.335 ;
        RECT 53.370 148.290 53.690 148.350 ;
        RECT 51.545 148.150 53.690 148.290 ;
        RECT 51.545 148.105 51.835 148.150 ;
        RECT 53.370 148.090 53.690 148.150 ;
        RECT 54.750 148.090 55.070 148.350 ;
        RECT 68.105 148.290 68.395 148.335 ;
        RECT 69.930 148.290 70.250 148.350 ;
        RECT 68.105 148.150 70.250 148.290 ;
        RECT 68.105 148.105 68.395 148.150 ;
        RECT 69.930 148.090 70.250 148.150 ;
        RECT 74.545 148.290 74.835 148.335 ;
        RECT 80.510 148.290 80.830 148.350 ;
        RECT 74.545 148.150 80.830 148.290 ;
        RECT 74.545 148.105 74.835 148.150 ;
        RECT 80.510 148.090 80.830 148.150 ;
        RECT 98.005 148.290 98.295 148.335 ;
        RECT 99.370 148.290 99.690 148.350 ;
        RECT 98.005 148.150 99.690 148.290 ;
        RECT 98.005 148.105 98.295 148.150 ;
        RECT 99.370 148.090 99.690 148.150 ;
        RECT 99.830 148.090 100.150 148.350 ;
        RECT 108.585 148.290 108.875 148.335 ;
        RECT 109.030 148.290 109.350 148.350 ;
        RECT 108.585 148.150 109.350 148.290 ;
        RECT 108.585 148.105 108.875 148.150 ;
        RECT 109.030 148.090 109.350 148.150 ;
        RECT 112.250 148.090 112.570 148.350 ;
        RECT 124.210 148.090 124.530 148.350 ;
        RECT 35.400 147.950 35.690 147.995 ;
        RECT 38.180 147.950 38.470 147.995 ;
        RECT 40.040 147.950 40.330 147.995 ;
        RECT 35.400 147.810 40.330 147.950 ;
        RECT 35.400 147.765 35.690 147.810 ;
        RECT 38.180 147.765 38.470 147.810 ;
        RECT 40.040 147.765 40.330 147.810 ;
        RECT 43.710 147.950 44.030 148.010 ;
        RECT 52.465 147.950 52.755 147.995 ;
        RECT 74.070 147.950 74.390 148.010 ;
        RECT 43.710 147.810 49.460 147.950 ;
        RECT 43.710 147.750 44.030 147.810 ;
        RECT 40.505 147.610 40.795 147.655 ;
        RECT 42.790 147.610 43.110 147.670 ;
        RECT 40.505 147.470 43.110 147.610 ;
        RECT 40.505 147.425 40.795 147.470 ;
        RECT 42.790 147.410 43.110 147.470 ;
        RECT 45.550 147.410 45.870 147.670 ;
        RECT 48.785 147.610 49.075 147.655 ;
        RECT 46.560 147.470 49.075 147.610 ;
        RECT 49.320 147.610 49.460 147.810 ;
        RECT 52.465 147.810 74.390 147.950 ;
        RECT 52.465 147.765 52.755 147.810 ;
        RECT 74.070 147.750 74.390 147.810 ;
        RECT 90.600 147.950 90.890 147.995 ;
        RECT 93.380 147.950 93.670 147.995 ;
        RECT 95.240 147.950 95.530 147.995 ;
        RECT 102.130 147.950 102.450 148.010 ;
        RECT 90.600 147.810 95.530 147.950 ;
        RECT 90.600 147.765 90.890 147.810 ;
        RECT 93.380 147.765 93.670 147.810 ;
        RECT 95.240 147.765 95.530 147.810 ;
        RECT 99.460 147.810 102.450 147.950 ;
        RECT 49.320 147.470 53.600 147.610 ;
        RECT 35.400 147.270 35.690 147.315 ;
        RECT 35.400 147.130 37.935 147.270 ;
        RECT 35.400 147.085 35.690 147.130 ;
        RECT 32.210 146.930 32.530 146.990 ;
        RECT 37.720 146.975 37.935 147.130 ;
        RECT 38.650 147.070 38.970 147.330 ;
        RECT 46.560 147.270 46.700 147.470 ;
        RECT 48.785 147.425 49.075 147.470 ;
        RECT 40.120 147.130 46.700 147.270 ;
        RECT 47.865 147.270 48.155 147.315 ;
        RECT 50.610 147.270 50.930 147.330 ;
        RECT 53.460 147.315 53.600 147.470 ;
        RECT 54.290 147.410 54.610 147.670 ;
        RECT 58.430 147.410 58.750 147.670 ;
        RECT 65.345 147.610 65.635 147.655 ;
        RECT 67.170 147.610 67.490 147.670 ;
        RECT 65.345 147.470 67.490 147.610 ;
        RECT 65.345 147.425 65.635 147.470 ;
        RECT 67.170 147.410 67.490 147.470 ;
        RECT 71.770 147.410 72.090 147.670 ;
        RECT 89.710 147.610 90.030 147.670 ;
        RECT 93.865 147.610 94.155 147.655 ;
        RECT 89.710 147.470 94.155 147.610 ;
        RECT 89.710 147.410 90.030 147.470 ;
        RECT 93.865 147.425 94.155 147.470 ;
        RECT 95.690 147.610 96.010 147.670 ;
        RECT 99.460 147.610 99.600 147.810 ;
        RECT 102.130 147.750 102.450 147.810 ;
        RECT 117.740 147.950 118.030 147.995 ;
        RECT 120.520 147.950 120.810 147.995 ;
        RECT 122.380 147.950 122.670 147.995 ;
        RECT 117.740 147.810 122.670 147.950 ;
        RECT 117.740 147.765 118.030 147.810 ;
        RECT 120.520 147.765 120.810 147.810 ;
        RECT 122.380 147.765 122.670 147.810 ;
        RECT 95.690 147.470 99.600 147.610 ;
        RECT 99.845 147.610 100.135 147.655 ;
        RECT 103.050 147.610 103.370 147.670 ;
        RECT 99.845 147.470 103.370 147.610 ;
        RECT 95.690 147.410 96.010 147.470 ;
        RECT 99.845 147.425 100.135 147.470 ;
        RECT 103.050 147.410 103.370 147.470 ;
        RECT 103.510 147.410 103.830 147.670 ;
        RECT 108.110 147.410 108.430 147.670 ;
        RECT 111.805 147.610 112.095 147.655 ;
        RECT 114.090 147.610 114.410 147.670 ;
        RECT 111.805 147.470 114.410 147.610 ;
        RECT 111.805 147.425 112.095 147.470 ;
        RECT 114.090 147.410 114.410 147.470 ;
        RECT 122.845 147.610 123.135 147.655 ;
        RECT 126.050 147.610 126.370 147.670 ;
        RECT 122.845 147.470 126.370 147.610 ;
        RECT 122.845 147.425 123.135 147.470 ;
        RECT 126.050 147.410 126.370 147.470 ;
        RECT 47.865 147.130 51.760 147.270 ;
        RECT 33.540 146.930 33.830 146.975 ;
        RECT 36.800 146.930 37.090 146.975 ;
        RECT 32.210 146.790 37.090 146.930 ;
        RECT 32.210 146.730 32.530 146.790 ;
        RECT 33.540 146.745 33.830 146.790 ;
        RECT 36.800 146.745 37.090 146.790 ;
        RECT 37.720 146.930 38.010 146.975 ;
        RECT 39.580 146.930 39.870 146.975 ;
        RECT 37.720 146.790 39.870 146.930 ;
        RECT 37.720 146.745 38.010 146.790 ;
        RECT 39.580 146.745 39.870 146.790 ;
        RECT 31.535 146.590 31.825 146.635 ;
        RECT 34.970 146.590 35.290 146.650 ;
        RECT 40.120 146.590 40.260 147.130 ;
        RECT 47.865 147.085 48.155 147.130 ;
        RECT 50.610 147.070 50.930 147.130 ;
        RECT 44.645 146.930 44.935 146.975 ;
        RECT 51.070 146.930 51.390 146.990 ;
        RECT 44.645 146.790 51.390 146.930 ;
        RECT 44.645 146.745 44.935 146.790 ;
        RECT 51.070 146.730 51.390 146.790 ;
        RECT 31.535 146.450 40.260 146.590 ;
        RECT 45.105 146.590 45.395 146.635 ;
        RECT 48.770 146.590 49.090 146.650 ;
        RECT 49.690 146.590 50.010 146.650 ;
        RECT 45.105 146.450 50.010 146.590 ;
        RECT 51.620 146.590 51.760 147.130 ;
        RECT 52.005 147.085 52.295 147.315 ;
        RECT 53.385 147.085 53.675 147.315 ;
        RECT 54.765 147.270 55.055 147.315 ;
        RECT 55.670 147.270 55.990 147.330 ;
        RECT 54.765 147.130 55.990 147.270 ;
        RECT 54.765 147.085 55.055 147.130 ;
        RECT 52.080 146.930 52.220 147.085 ;
        RECT 55.670 147.070 55.990 147.130 ;
        RECT 56.130 147.270 56.450 147.330 ;
        RECT 61.190 147.270 61.510 147.330 ;
        RECT 56.130 147.130 61.510 147.270 ;
        RECT 56.130 147.070 56.450 147.130 ;
        RECT 61.190 147.070 61.510 147.130 ;
        RECT 69.930 147.270 70.250 147.330 ;
        RECT 72.705 147.270 72.995 147.315 ;
        RECT 69.930 147.130 72.995 147.270 ;
        RECT 69.930 147.070 70.250 147.130 ;
        RECT 72.705 147.085 72.995 147.130 ;
        RECT 90.600 147.270 90.890 147.315 ;
        RECT 94.310 147.270 94.630 147.330 ;
        RECT 97.545 147.270 97.835 147.315 ;
        RECT 90.600 147.130 93.135 147.270 ;
        RECT 90.600 147.085 90.890 147.130 ;
        RECT 56.590 146.930 56.910 146.990 ;
        RECT 76.370 146.930 76.690 146.990 ;
        RECT 52.080 146.790 56.910 146.930 ;
        RECT 56.590 146.730 56.910 146.790 ;
        RECT 61.280 146.790 76.690 146.930 ;
        RECT 61.280 146.590 61.420 146.790 ;
        RECT 76.370 146.730 76.690 146.790 ;
        RECT 88.740 146.930 89.030 146.975 ;
        RECT 91.090 146.930 91.410 146.990 ;
        RECT 92.920 146.975 93.135 147.130 ;
        RECT 94.310 147.130 97.835 147.270 ;
        RECT 94.310 147.070 94.630 147.130 ;
        RECT 97.545 147.085 97.835 147.130 ;
        RECT 97.990 147.270 98.310 147.330 ;
        RECT 98.925 147.270 99.215 147.315 ;
        RECT 97.990 147.130 99.215 147.270 ;
        RECT 97.990 147.070 98.310 147.130 ;
        RECT 98.925 147.085 99.215 147.130 ;
        RECT 100.290 147.070 100.610 147.330 ;
        RECT 107.190 147.070 107.510 147.330 ;
        RECT 108.585 147.270 108.875 147.315 ;
        RECT 110.410 147.270 110.730 147.330 ;
        RECT 108.585 147.130 110.730 147.270 ;
        RECT 108.585 147.085 108.875 147.130 ;
        RECT 110.410 147.070 110.730 147.130 ;
        RECT 110.885 147.270 111.175 147.315 ;
        RECT 111.330 147.270 111.650 147.330 ;
        RECT 110.885 147.130 111.650 147.270 ;
        RECT 110.885 147.085 111.175 147.130 ;
        RECT 111.330 147.070 111.650 147.130 ;
        RECT 112.265 147.270 112.555 147.315 ;
        RECT 114.550 147.270 114.870 147.330 ;
        RECT 112.265 147.130 114.870 147.270 ;
        RECT 112.265 147.085 112.555 147.130 ;
        RECT 114.550 147.070 114.870 147.130 ;
        RECT 117.740 147.270 118.030 147.315 ;
        RECT 120.530 147.270 120.850 147.330 ;
        RECT 121.005 147.270 121.295 147.315 ;
        RECT 117.740 147.130 120.275 147.270 ;
        RECT 117.740 147.085 118.030 147.130 ;
        RECT 92.000 146.930 92.290 146.975 ;
        RECT 88.740 146.790 92.290 146.930 ;
        RECT 88.740 146.745 89.030 146.790 ;
        RECT 91.090 146.730 91.410 146.790 ;
        RECT 92.000 146.745 92.290 146.790 ;
        RECT 92.920 146.930 93.210 146.975 ;
        RECT 94.780 146.930 95.070 146.975 ;
        RECT 92.920 146.790 95.070 146.930 ;
        RECT 92.920 146.745 93.210 146.790 ;
        RECT 94.780 146.745 95.070 146.790 ;
        RECT 98.450 146.930 98.770 146.990 ;
        RECT 115.930 146.975 116.250 146.990 ;
        RECT 120.060 146.975 120.275 147.130 ;
        RECT 120.530 147.130 121.295 147.270 ;
        RECT 120.530 147.070 120.850 147.130 ;
        RECT 121.005 147.085 121.295 147.130 ;
        RECT 121.450 147.270 121.770 147.330 ;
        RECT 123.305 147.270 123.595 147.315 ;
        RECT 121.450 147.130 123.595 147.270 ;
        RECT 121.450 147.070 121.770 147.130 ;
        RECT 123.305 147.085 123.595 147.130 ;
        RECT 104.445 146.930 104.735 146.975 ;
        RECT 98.450 146.790 104.735 146.930 ;
        RECT 98.450 146.730 98.770 146.790 ;
        RECT 104.445 146.745 104.735 146.790 ;
        RECT 104.905 146.930 105.195 146.975 ;
        RECT 115.880 146.930 116.250 146.975 ;
        RECT 119.140 146.930 119.430 146.975 ;
        RECT 104.905 146.790 112.940 146.930 ;
        RECT 104.905 146.745 105.195 146.790 ;
        RECT 112.800 146.650 112.940 146.790 ;
        RECT 115.880 146.790 119.430 146.930 ;
        RECT 115.880 146.745 116.250 146.790 ;
        RECT 119.140 146.745 119.430 146.790 ;
        RECT 120.060 146.930 120.350 146.975 ;
        RECT 121.920 146.930 122.210 146.975 ;
        RECT 120.060 146.790 122.210 146.930 ;
        RECT 120.060 146.745 120.350 146.790 ;
        RECT 121.920 146.745 122.210 146.790 ;
        RECT 115.930 146.730 116.250 146.745 ;
        RECT 51.620 146.450 61.420 146.590 ;
        RECT 61.665 146.590 61.955 146.635 ;
        RECT 67.170 146.590 67.490 146.650 ;
        RECT 61.665 146.450 67.490 146.590 ;
        RECT 31.535 146.405 31.825 146.450 ;
        RECT 34.970 146.390 35.290 146.450 ;
        RECT 45.105 146.405 45.395 146.450 ;
        RECT 48.770 146.390 49.090 146.450 ;
        RECT 49.690 146.390 50.010 146.450 ;
        RECT 61.665 146.405 61.955 146.450 ;
        RECT 67.170 146.390 67.490 146.450 ;
        RECT 72.245 146.590 72.535 146.635 ;
        RECT 73.610 146.590 73.930 146.650 ;
        RECT 72.245 146.450 73.930 146.590 ;
        RECT 72.245 146.405 72.535 146.450 ;
        RECT 73.610 146.390 73.930 146.450 ;
        RECT 86.030 146.590 86.350 146.650 ;
        RECT 86.735 146.590 87.025 146.635 ;
        RECT 86.030 146.450 87.025 146.590 ;
        RECT 86.030 146.390 86.350 146.450 ;
        RECT 86.735 146.405 87.025 146.450 ;
        RECT 101.225 146.590 101.515 146.635 ;
        RECT 103.050 146.590 103.370 146.650 ;
        RECT 101.225 146.450 103.370 146.590 ;
        RECT 101.225 146.405 101.515 146.450 ;
        RECT 103.050 146.390 103.370 146.450 ;
        RECT 105.810 146.590 106.130 146.650 ;
        RECT 106.745 146.590 107.035 146.635 ;
        RECT 105.810 146.450 107.035 146.590 ;
        RECT 105.810 146.390 106.130 146.450 ;
        RECT 106.745 146.405 107.035 146.450 ;
        RECT 109.490 146.390 109.810 146.650 ;
        RECT 109.965 146.590 110.255 146.635 ;
        RECT 110.410 146.590 110.730 146.650 ;
        RECT 109.965 146.450 110.730 146.590 ;
        RECT 109.965 146.405 110.255 146.450 ;
        RECT 110.410 146.390 110.730 146.450 ;
        RECT 112.710 146.590 113.030 146.650 ;
        RECT 113.875 146.590 114.165 146.635 ;
        RECT 116.390 146.590 116.710 146.650 ;
        RECT 112.710 146.450 116.710 146.590 ;
        RECT 112.710 146.390 113.030 146.450 ;
        RECT 113.875 146.405 114.165 146.450 ;
        RECT 116.390 146.390 116.710 146.450 ;
        RECT 29.840 145.770 127.820 146.250 ;
        RECT 32.210 145.370 32.530 145.630 ;
        RECT 34.510 145.370 34.830 145.630 ;
        RECT 34.970 145.370 35.290 145.630 ;
        RECT 36.825 145.385 37.115 145.615 ;
        RECT 31.290 144.890 31.610 144.950 ;
        RECT 32.685 144.890 32.975 144.935 ;
        RECT 36.900 144.890 37.040 145.385 ;
        RECT 38.650 145.370 38.970 145.630 ;
        RECT 63.950 145.370 64.270 145.630 ;
        RECT 83.730 145.570 84.050 145.630 ;
        RECT 68.640 145.430 84.050 145.570 ;
        RECT 62.570 145.030 62.890 145.290 ;
        RECT 65.790 145.030 66.110 145.290 ;
        RECT 37.745 144.890 38.035 144.935 ;
        RECT 31.290 144.750 33.820 144.890 ;
        RECT 36.900 144.750 38.035 144.890 ;
        RECT 62.660 144.890 62.800 145.030 ;
        RECT 63.950 144.890 64.270 144.950 ;
        RECT 62.660 144.750 64.270 144.890 ;
        RECT 31.290 144.690 31.610 144.750 ;
        RECT 32.685 144.705 32.975 144.750 ;
        RECT 33.680 144.210 33.820 144.750 ;
        RECT 37.745 144.705 38.035 144.750 ;
        RECT 63.950 144.690 64.270 144.750 ;
        RECT 64.870 144.690 65.190 144.950 ;
        RECT 65.345 144.705 65.635 144.935 ;
        RECT 66.725 144.890 67.015 144.935 ;
        RECT 67.170 144.890 67.490 144.950 ;
        RECT 66.725 144.750 67.490 144.890 ;
        RECT 66.725 144.705 67.015 144.750 ;
        RECT 34.050 144.550 34.370 144.610 ;
        RECT 45.550 144.550 45.870 144.610 ;
        RECT 34.050 144.410 45.870 144.550 ;
        RECT 34.050 144.350 34.370 144.410 ;
        RECT 45.550 144.350 45.870 144.410 ;
        RECT 37.270 144.210 37.590 144.270 ;
        RECT 33.680 144.070 37.590 144.210 ;
        RECT 65.420 144.210 65.560 144.705 ;
        RECT 67.170 144.690 67.490 144.750 ;
        RECT 68.090 144.890 68.410 144.950 ;
        RECT 68.640 144.935 68.780 145.430 ;
        RECT 76.370 145.030 76.690 145.290 ;
        RECT 77.305 145.230 77.595 145.275 ;
        RECT 78.670 145.230 78.990 145.290 ;
        RECT 77.305 145.090 78.990 145.230 ;
        RECT 77.305 145.045 77.595 145.090 ;
        RECT 78.670 145.030 78.990 145.090 ;
        RECT 80.525 145.230 80.815 145.275 ;
        RECT 80.985 145.230 81.275 145.275 ;
        RECT 80.525 145.090 81.275 145.230 ;
        RECT 80.525 145.045 80.815 145.090 ;
        RECT 80.985 145.045 81.275 145.090 ;
        RECT 68.565 144.890 68.855 144.935 ;
        RECT 68.090 144.750 68.855 144.890 ;
        RECT 68.090 144.690 68.410 144.750 ;
        RECT 68.565 144.705 68.855 144.750 ;
        RECT 69.025 144.705 69.315 144.935 ;
        RECT 69.485 144.705 69.775 144.935 ;
        RECT 69.930 144.890 70.250 144.950 ;
        RECT 70.405 144.890 70.695 144.935 ;
        RECT 70.850 144.890 71.170 144.950 ;
        RECT 69.930 144.750 71.170 144.890 ;
        RECT 67.630 144.550 67.950 144.610 ;
        RECT 69.100 144.550 69.240 144.705 ;
        RECT 67.630 144.410 69.240 144.550 ;
        RECT 69.560 144.550 69.700 144.705 ;
        RECT 69.930 144.690 70.250 144.750 ;
        RECT 70.405 144.705 70.695 144.750 ;
        RECT 70.850 144.690 71.170 144.750 ;
        RECT 74.990 144.690 75.310 144.950 ;
        RECT 79.145 144.890 79.435 144.935 ;
        RECT 81.430 144.890 81.750 144.950 ;
        RECT 79.145 144.750 81.750 144.890 ;
        RECT 81.980 144.890 82.120 145.430 ;
        RECT 83.730 145.370 84.050 145.430 ;
        RECT 91.105 145.570 91.395 145.615 ;
        RECT 98.450 145.570 98.770 145.630 ;
        RECT 91.105 145.430 98.770 145.570 ;
        RECT 91.105 145.385 91.395 145.430 ;
        RECT 98.450 145.370 98.770 145.430 ;
        RECT 104.430 145.570 104.750 145.630 ;
        RECT 104.905 145.570 105.195 145.615 ;
        RECT 104.430 145.430 105.195 145.570 ;
        RECT 104.430 145.370 104.750 145.430 ;
        RECT 104.905 145.385 105.195 145.430 ;
        RECT 116.390 145.370 116.710 145.630 ;
        RECT 116.850 145.370 117.170 145.630 ;
        RECT 120.530 145.370 120.850 145.630 ;
        RECT 86.030 145.230 86.350 145.290 ;
        RECT 83.360 145.090 86.350 145.230 ;
        RECT 82.365 144.890 82.655 144.935 ;
        RECT 81.980 144.750 82.655 144.890 ;
        RECT 79.145 144.705 79.435 144.750 ;
        RECT 81.430 144.690 81.750 144.750 ;
        RECT 82.365 144.705 82.655 144.750 ;
        RECT 73.610 144.550 73.930 144.610 ;
        RECT 69.560 144.410 73.930 144.550 ;
        RECT 67.630 144.350 67.950 144.410 ;
        RECT 73.610 144.350 73.930 144.410 ;
        RECT 80.065 144.550 80.355 144.595 ;
        RECT 81.890 144.550 82.210 144.610 ;
        RECT 80.065 144.410 82.210 144.550 ;
        RECT 80.065 144.365 80.355 144.410 ;
        RECT 81.890 144.350 82.210 144.410 ;
        RECT 79.590 144.210 79.910 144.270 ;
        RECT 81.430 144.210 81.750 144.270 ;
        RECT 65.420 144.070 81.750 144.210 ;
        RECT 82.440 144.210 82.580 144.705 ;
        RECT 82.810 144.690 83.130 144.950 ;
        RECT 83.360 144.935 83.500 145.090 ;
        RECT 86.030 145.030 86.350 145.090 ;
        RECT 102.130 145.030 102.450 145.290 ;
        RECT 83.285 144.705 83.575 144.935 ;
        RECT 84.190 144.690 84.510 144.950 ;
        RECT 86.505 144.890 86.795 144.935 ;
        RECT 93.405 144.890 93.695 144.935 ;
        RECT 93.850 144.890 94.170 144.950 ;
        RECT 86.505 144.750 90.860 144.890 ;
        RECT 86.505 144.705 86.795 144.750 ;
        RECT 82.900 144.550 83.040 144.690 ;
        RECT 90.720 144.610 90.860 144.750 ;
        RECT 93.405 144.750 94.170 144.890 ;
        RECT 93.405 144.705 93.695 144.750 ;
        RECT 93.850 144.690 94.170 144.750 ;
        RECT 105.810 144.690 106.130 144.950 ;
        RECT 119.665 144.705 119.955 144.935 ;
        RECT 85.585 144.550 85.875 144.595 ;
        RECT 86.950 144.550 87.270 144.610 ;
        RECT 89.725 144.550 90.015 144.595 ;
        RECT 82.900 144.410 85.340 144.550 ;
        RECT 83.270 144.210 83.590 144.270 ;
        RECT 82.440 144.070 83.590 144.210 ;
        RECT 85.200 144.210 85.340 144.410 ;
        RECT 85.585 144.410 90.015 144.550 ;
        RECT 85.585 144.365 85.875 144.410 ;
        RECT 86.950 144.350 87.270 144.410 ;
        RECT 89.725 144.365 90.015 144.410 ;
        RECT 90.630 144.350 90.950 144.610 ;
        RECT 115.470 144.350 115.790 144.610 ;
        RECT 119.700 144.550 119.840 144.705 ;
        RECT 118.780 144.410 119.840 144.550 ;
        RECT 86.030 144.210 86.350 144.270 ;
        RECT 118.780 144.255 118.920 144.410 ;
        RECT 85.200 144.070 86.350 144.210 ;
        RECT 37.270 144.010 37.590 144.070 ;
        RECT 79.590 144.010 79.910 144.070 ;
        RECT 81.430 144.010 81.750 144.070 ;
        RECT 83.270 144.010 83.590 144.070 ;
        RECT 86.030 144.010 86.350 144.070 ;
        RECT 118.705 144.025 118.995 144.255 ;
        RECT 56.130 143.670 56.450 143.930 ;
        RECT 66.710 143.870 67.030 143.930 ;
        RECT 67.185 143.870 67.475 143.915 ;
        RECT 66.710 143.730 67.475 143.870 ;
        RECT 66.710 143.670 67.030 143.730 ;
        RECT 67.185 143.685 67.475 143.730 ;
        RECT 75.925 143.870 76.215 143.915 ;
        RECT 76.370 143.870 76.690 143.930 ;
        RECT 75.925 143.730 76.690 143.870 ;
        RECT 75.925 143.685 76.215 143.730 ;
        RECT 76.370 143.670 76.690 143.730 ;
        RECT 78.225 143.870 78.515 143.915 ;
        RECT 79.130 143.870 79.450 143.930 ;
        RECT 78.225 143.730 79.450 143.870 ;
        RECT 78.225 143.685 78.515 143.730 ;
        RECT 79.130 143.670 79.450 143.730 ;
        RECT 80.525 143.870 80.815 143.915 ;
        RECT 82.810 143.870 83.130 143.930 ;
        RECT 80.525 143.730 83.130 143.870 ;
        RECT 80.525 143.685 80.815 143.730 ;
        RECT 82.810 143.670 83.130 143.730 ;
        RECT 88.330 143.670 88.650 143.930 ;
        RECT 92.945 143.870 93.235 143.915 ;
        RECT 94.310 143.870 94.630 143.930 ;
        RECT 92.945 143.730 94.630 143.870 ;
        RECT 92.945 143.685 93.235 143.730 ;
        RECT 94.310 143.670 94.630 143.730 ;
        RECT 29.840 143.050 127.820 143.530 ;
        RECT 41.410 142.850 41.730 142.910 ;
        RECT 54.750 142.850 55.070 142.910 ;
        RECT 55.685 142.850 55.975 142.895 ;
        RECT 41.410 142.710 54.520 142.850 ;
        RECT 41.410 142.650 41.730 142.710 ;
        RECT 36.320 142.510 36.610 142.555 ;
        RECT 39.100 142.510 39.390 142.555 ;
        RECT 40.960 142.510 41.250 142.555 ;
        RECT 36.320 142.370 41.250 142.510 ;
        RECT 36.320 142.325 36.610 142.370 ;
        RECT 39.100 142.325 39.390 142.370 ;
        RECT 40.960 142.325 41.250 142.370 ;
        RECT 42.330 142.510 42.650 142.570 ;
        RECT 46.025 142.510 46.315 142.555 ;
        RECT 42.330 142.370 46.315 142.510 ;
        RECT 42.330 142.310 42.650 142.370 ;
        RECT 46.025 142.325 46.315 142.370 ;
        RECT 32.455 142.170 32.745 142.215 ;
        RECT 35.430 142.170 35.750 142.230 ;
        RECT 32.455 142.030 35.750 142.170 ;
        RECT 32.455 141.985 32.745 142.030 ;
        RECT 35.430 141.970 35.750 142.030 ;
        RECT 37.270 142.170 37.590 142.230 ;
        RECT 41.425 142.170 41.715 142.215 ;
        RECT 42.790 142.170 43.110 142.230 ;
        RECT 37.270 142.030 40.260 142.170 ;
        RECT 37.270 141.970 37.590 142.030 ;
        RECT 36.320 141.830 36.610 141.875 ;
        RECT 36.320 141.690 38.855 141.830 ;
        RECT 36.320 141.645 36.610 141.690 ;
        RECT 32.210 141.490 32.530 141.550 ;
        RECT 38.640 141.535 38.855 141.690 ;
        RECT 39.570 141.630 39.890 141.890 ;
        RECT 40.120 141.830 40.260 142.030 ;
        RECT 41.425 142.030 43.110 142.170 ;
        RECT 41.425 141.985 41.715 142.030 ;
        RECT 42.790 141.970 43.110 142.030 ;
        RECT 45.550 142.170 45.870 142.230 ;
        RECT 48.785 142.170 49.075 142.215 ;
        RECT 53.845 142.170 54.135 142.215 ;
        RECT 45.550 142.030 49.075 142.170 ;
        RECT 45.550 141.970 45.870 142.030 ;
        RECT 48.785 141.985 49.075 142.030 ;
        RECT 53.460 142.030 54.135 142.170 ;
        RECT 54.380 142.170 54.520 142.710 ;
        RECT 54.750 142.710 55.975 142.850 ;
        RECT 54.750 142.650 55.070 142.710 ;
        RECT 55.685 142.665 55.975 142.710 ;
        RECT 57.510 142.650 57.830 142.910 ;
        RECT 63.045 142.850 63.335 142.895 ;
        RECT 60.820 142.710 63.335 142.850 ;
        RECT 56.590 142.510 56.910 142.570 ;
        RECT 60.820 142.510 60.960 142.710 ;
        RECT 63.045 142.665 63.335 142.710 ;
        RECT 65.345 142.850 65.635 142.895 ;
        RECT 69.470 142.850 69.790 142.910 ;
        RECT 65.345 142.710 69.790 142.850 ;
        RECT 65.345 142.665 65.635 142.710 ;
        RECT 69.470 142.650 69.790 142.710 ;
        RECT 74.990 142.850 75.310 142.910 ;
        RECT 75.465 142.850 75.755 142.895 ;
        RECT 74.990 142.710 75.755 142.850 ;
        RECT 74.990 142.650 75.310 142.710 ;
        RECT 75.465 142.665 75.755 142.710 ;
        RECT 83.270 142.650 83.590 142.910 ;
        RECT 83.730 142.650 84.050 142.910 ;
        RECT 89.710 142.650 90.030 142.910 ;
        RECT 90.645 142.850 90.935 142.895 ;
        RECT 91.090 142.850 91.410 142.910 ;
        RECT 90.645 142.710 91.410 142.850 ;
        RECT 90.645 142.665 90.935 142.710 ;
        RECT 91.090 142.650 91.410 142.710 ;
        RECT 94.770 142.650 95.090 142.910 ;
        RECT 108.585 142.850 108.875 142.895 ;
        RECT 109.030 142.850 109.350 142.910 ;
        RECT 108.585 142.710 109.350 142.850 ;
        RECT 108.585 142.665 108.875 142.710 ;
        RECT 109.030 142.650 109.350 142.710 ;
        RECT 112.250 142.650 112.570 142.910 ;
        RECT 112.725 142.850 113.015 142.895 ;
        RECT 113.630 142.850 113.950 142.910 ;
        RECT 112.725 142.710 113.950 142.850 ;
        RECT 112.725 142.665 113.015 142.710 ;
        RECT 113.630 142.650 113.950 142.710 ;
        RECT 56.590 142.370 60.960 142.510 ;
        RECT 65.790 142.510 66.110 142.570 ;
        RECT 83.360 142.510 83.500 142.650 ;
        RECT 94.860 142.510 95.000 142.650 ;
        RECT 65.790 142.370 72.000 142.510 ;
        RECT 83.360 142.370 85.340 142.510 ;
        RECT 56.590 142.310 56.910 142.370 ;
        RECT 65.790 142.310 66.110 142.370 ;
        RECT 71.860 142.230 72.000 142.370 ;
        RECT 57.525 142.170 57.815 142.215 ;
        RECT 54.380 142.030 57.815 142.170 ;
        RECT 44.645 141.830 44.935 141.875 ;
        RECT 53.460 141.830 53.600 142.030 ;
        RECT 53.845 141.985 54.135 142.030 ;
        RECT 57.525 141.985 57.815 142.030 ;
        RECT 59.810 142.170 60.130 142.230 ;
        RECT 63.505 142.170 63.795 142.215 ;
        RECT 66.710 142.170 67.030 142.230 ;
        RECT 70.850 142.170 71.170 142.230 ;
        RECT 59.810 142.030 63.795 142.170 ;
        RECT 59.810 141.970 60.130 142.030 ;
        RECT 63.505 141.985 63.795 142.030 ;
        RECT 64.040 142.030 67.030 142.170 ;
        RECT 54.765 141.830 55.055 141.875 ;
        RECT 40.120 141.690 44.935 141.830 ;
        RECT 44.645 141.645 44.935 141.690 ;
        RECT 45.180 141.690 53.600 141.830 ;
        RECT 53.920 141.690 55.055 141.830 ;
        RECT 34.460 141.490 34.750 141.535 ;
        RECT 37.720 141.490 38.010 141.535 ;
        RECT 32.210 141.350 38.010 141.490 ;
        RECT 32.210 141.290 32.530 141.350 ;
        RECT 34.460 141.305 34.750 141.350 ;
        RECT 37.720 141.305 38.010 141.350 ;
        RECT 38.640 141.490 38.930 141.535 ;
        RECT 40.500 141.490 40.790 141.535 ;
        RECT 45.180 141.490 45.320 141.690 ;
        RECT 38.640 141.350 40.790 141.490 ;
        RECT 38.640 141.305 38.930 141.350 ;
        RECT 40.500 141.305 40.790 141.350 ;
        RECT 41.040 141.350 45.320 141.490 ;
        RECT 48.325 141.490 48.615 141.535 ;
        RECT 50.150 141.490 50.470 141.550 ;
        RECT 48.325 141.350 50.470 141.490 ;
        RECT 35.430 141.150 35.750 141.210 ;
        RECT 41.040 141.150 41.180 141.350 ;
        RECT 48.325 141.305 48.615 141.350 ;
        RECT 50.150 141.290 50.470 141.350 ;
        RECT 53.370 141.490 53.690 141.550 ;
        RECT 53.920 141.490 54.060 141.690 ;
        RECT 54.765 141.645 55.055 141.690 ;
        RECT 57.050 141.630 57.370 141.890 ;
        RECT 63.045 141.830 63.335 141.875 ;
        RECT 64.040 141.830 64.180 142.030 ;
        RECT 66.710 141.970 67.030 142.030 ;
        RECT 68.180 142.030 71.170 142.170 ;
        RECT 58.060 141.690 62.800 141.830 ;
        RECT 53.370 141.350 54.060 141.490 ;
        RECT 54.290 141.490 54.610 141.550 ;
        RECT 58.060 141.490 58.200 141.690 ;
        RECT 54.290 141.350 58.200 141.490 ;
        RECT 53.370 141.290 53.690 141.350 ;
        RECT 54.290 141.290 54.610 141.350 ;
        RECT 58.430 141.290 58.750 141.550 ;
        RECT 62.660 141.490 62.800 141.690 ;
        RECT 63.045 141.690 64.180 141.830 ;
        RECT 63.045 141.645 63.335 141.690 ;
        RECT 64.410 141.630 64.730 141.890 ;
        RECT 67.170 141.630 67.490 141.890 ;
        RECT 67.630 141.630 67.950 141.890 ;
        RECT 68.180 141.875 68.320 142.030 ;
        RECT 70.850 141.970 71.170 142.030 ;
        RECT 71.770 142.170 72.090 142.230 ;
        RECT 72.245 142.170 72.535 142.215 ;
        RECT 71.770 142.030 72.535 142.170 ;
        RECT 71.770 141.970 72.090 142.030 ;
        RECT 72.245 141.985 72.535 142.030 ;
        RECT 78.670 141.970 78.990 142.230 ;
        RECT 80.525 142.170 80.815 142.215 ;
        RECT 81.430 142.170 81.750 142.230 ;
        RECT 80.525 142.030 81.750 142.170 ;
        RECT 80.525 141.985 80.815 142.030 ;
        RECT 81.430 141.970 81.750 142.030 ;
        RECT 83.270 141.970 83.590 142.230 ;
        RECT 84.190 142.170 84.510 142.230 ;
        RECT 84.190 142.030 84.880 142.170 ;
        RECT 84.190 141.970 84.510 142.030 ;
        RECT 68.105 141.645 68.395 141.875 ;
        RECT 69.025 141.830 69.315 141.875 ;
        RECT 69.930 141.830 70.250 141.890 ;
        RECT 69.025 141.690 70.250 141.830 ;
        RECT 69.025 141.645 69.315 141.690 ;
        RECT 69.930 141.630 70.250 141.690 ;
        RECT 70.390 141.630 70.710 141.890 ;
        RECT 73.610 141.630 73.930 141.890 ;
        RECT 77.765 141.830 78.055 141.875 ;
        RECT 78.760 141.830 78.900 141.970 ;
        RECT 79.605 141.830 79.895 141.875 ;
        RECT 77.765 141.690 79.895 141.830 ;
        RECT 77.765 141.645 78.055 141.690 ;
        RECT 79.605 141.645 79.895 141.690 ;
        RECT 82.350 141.630 82.670 141.890 ;
        RECT 78.685 141.490 78.975 141.535 ;
        RECT 80.510 141.490 80.830 141.550 ;
        RECT 62.660 141.350 80.830 141.490 ;
        RECT 78.685 141.305 78.975 141.350 ;
        RECT 80.510 141.290 80.830 141.350 ;
        RECT 83.745 141.490 84.035 141.535 ;
        RECT 84.205 141.490 84.495 141.535 ;
        RECT 83.745 141.350 84.495 141.490 ;
        RECT 84.740 141.490 84.880 142.030 ;
        RECT 85.200 141.830 85.340 142.370 ;
        RECT 94.400 142.370 95.000 142.510 ;
        RECT 95.660 142.510 95.950 142.555 ;
        RECT 98.440 142.510 98.730 142.555 ;
        RECT 100.300 142.510 100.590 142.555 ;
        RECT 95.660 142.370 100.590 142.510 ;
        RECT 90.630 142.170 90.950 142.230 ;
        RECT 91.795 142.170 92.085 142.215 ;
        RECT 86.580 142.030 92.085 142.170 ;
        RECT 85.585 141.830 85.875 141.875 ;
        RECT 85.200 141.690 85.875 141.830 ;
        RECT 85.585 141.645 85.875 141.690 ;
        RECT 86.030 141.630 86.350 141.890 ;
        RECT 86.580 141.875 86.720 142.030 ;
        RECT 90.630 141.970 90.950 142.030 ;
        RECT 91.795 141.985 92.085 142.030 ;
        RECT 86.505 141.645 86.795 141.875 ;
        RECT 87.425 141.645 87.715 141.875 ;
        RECT 88.330 141.830 88.650 141.890 ;
        RECT 88.805 141.830 89.095 141.875 ;
        RECT 88.330 141.690 89.095 141.830 ;
        RECT 87.500 141.490 87.640 141.645 ;
        RECT 88.330 141.630 88.650 141.690 ;
        RECT 88.805 141.645 89.095 141.690 ;
        RECT 91.105 141.830 91.395 141.875 ;
        RECT 94.400 141.830 94.540 142.370 ;
        RECT 95.660 142.325 95.950 142.370 ;
        RECT 98.440 142.325 98.730 142.370 ;
        RECT 100.300 142.325 100.590 142.370 ;
        RECT 94.770 142.170 95.090 142.230 ;
        RECT 98.925 142.170 99.215 142.215 ;
        RECT 94.770 142.030 99.215 142.170 ;
        RECT 94.770 141.970 95.090 142.030 ;
        RECT 98.925 141.985 99.215 142.030 ;
        RECT 100.765 142.170 101.055 142.215 ;
        RECT 102.130 142.170 102.450 142.230 ;
        RECT 100.765 142.030 102.450 142.170 ;
        RECT 100.765 141.985 101.055 142.030 ;
        RECT 102.130 141.970 102.450 142.030 ;
        RECT 113.170 142.170 113.490 142.230 ;
        RECT 115.485 142.170 115.775 142.215 ;
        RECT 113.170 142.030 115.775 142.170 ;
        RECT 113.170 141.970 113.490 142.030 ;
        RECT 115.485 141.985 115.775 142.030 ;
        RECT 91.105 141.690 94.540 141.830 ;
        RECT 95.660 141.830 95.950 141.875 ;
        RECT 106.270 141.830 106.590 141.890 ;
        RECT 106.745 141.830 107.035 141.875 ;
        RECT 95.660 141.690 98.195 141.830 ;
        RECT 91.105 141.645 91.395 141.690 ;
        RECT 95.660 141.645 95.950 141.690 ;
        RECT 84.740 141.350 87.640 141.490 ;
        RECT 93.800 141.490 94.090 141.535 ;
        RECT 96.150 141.490 96.470 141.550 ;
        RECT 97.980 141.535 98.195 141.690 ;
        RECT 106.270 141.690 107.035 141.830 ;
        RECT 106.270 141.630 106.590 141.690 ;
        RECT 106.745 141.645 107.035 141.690 ;
        RECT 107.665 141.830 107.955 141.875 ;
        RECT 109.030 141.830 109.350 141.890 ;
        RECT 107.665 141.690 109.350 141.830 ;
        RECT 107.665 141.645 107.955 141.690 ;
        RECT 109.030 141.630 109.350 141.690 ;
        RECT 110.870 141.630 111.190 141.890 ;
        RECT 111.345 141.830 111.635 141.875 ;
        RECT 113.645 141.830 113.935 141.875 ;
        RECT 111.345 141.690 113.935 141.830 ;
        RECT 111.345 141.645 111.635 141.690 ;
        RECT 113.645 141.645 113.935 141.690 ;
        RECT 114.550 141.830 114.870 141.890 ;
        RECT 116.405 141.830 116.695 141.875 ;
        RECT 114.550 141.690 116.695 141.830 ;
        RECT 97.060 141.490 97.350 141.535 ;
        RECT 93.800 141.350 97.350 141.490 ;
        RECT 83.745 141.305 84.035 141.350 ;
        RECT 84.205 141.305 84.495 141.350 ;
        RECT 93.800 141.305 94.090 141.350 ;
        RECT 96.150 141.290 96.470 141.350 ;
        RECT 97.060 141.305 97.350 141.350 ;
        RECT 97.980 141.490 98.270 141.535 ;
        RECT 99.840 141.490 100.130 141.535 ;
        RECT 97.980 141.350 100.130 141.490 ;
        RECT 109.120 141.490 109.260 141.630 ;
        RECT 111.420 141.490 111.560 141.645 ;
        RECT 114.550 141.630 114.870 141.690 ;
        RECT 116.405 141.645 116.695 141.690 ;
        RECT 109.120 141.350 111.560 141.490 ;
        RECT 97.980 141.305 98.270 141.350 ;
        RECT 99.840 141.305 100.130 141.350 ;
        RECT 135.635 141.220 136.775 165.470 ;
        RECT 35.430 141.010 41.180 141.150 ;
        RECT 45.105 141.150 45.395 141.195 ;
        RECT 46.470 141.150 46.790 141.210 ;
        RECT 45.105 141.010 46.790 141.150 ;
        RECT 35.430 140.950 35.750 141.010 ;
        RECT 45.105 140.965 45.395 141.010 ;
        RECT 46.470 140.950 46.790 141.010 ;
        RECT 47.865 141.150 48.155 141.195 ;
        RECT 49.690 141.150 50.010 141.210 ;
        RECT 47.865 141.010 50.010 141.150 ;
        RECT 47.865 140.965 48.155 141.010 ;
        RECT 49.690 140.950 50.010 141.010 ;
        RECT 54.750 141.150 55.070 141.210 ;
        RECT 56.145 141.150 56.435 141.195 ;
        RECT 54.750 141.010 56.435 141.150 ;
        RECT 54.750 140.950 55.070 141.010 ;
        RECT 56.145 140.965 56.435 141.010 ;
        RECT 60.270 141.150 60.590 141.210 ;
        RECT 65.805 141.150 66.095 141.195 ;
        RECT 60.270 141.010 66.095 141.150 ;
        RECT 60.270 140.950 60.590 141.010 ;
        RECT 65.805 140.965 66.095 141.010 ;
        RECT 67.170 141.150 67.490 141.210 ;
        RECT 68.090 141.150 68.410 141.210 ;
        RECT 67.170 141.010 68.410 141.150 ;
        RECT 67.170 140.950 67.490 141.010 ;
        RECT 68.090 140.950 68.410 141.010 ;
        RECT 70.865 141.150 71.155 141.195 ;
        RECT 72.690 141.150 73.010 141.210 ;
        RECT 70.865 141.010 73.010 141.150 ;
        RECT 70.865 140.965 71.155 141.010 ;
        RECT 72.690 140.950 73.010 141.010 ;
        RECT 73.150 140.950 73.470 141.210 ;
        RECT 75.910 141.150 76.230 141.210 ;
        RECT 77.305 141.150 77.595 141.195 ;
        RECT 75.910 141.010 77.595 141.150 ;
        RECT 75.910 140.950 76.230 141.010 ;
        RECT 77.305 140.965 77.595 141.010 ;
        RECT 81.445 141.150 81.735 141.195 ;
        RECT 99.370 141.150 99.690 141.210 ;
        RECT 81.445 141.010 99.690 141.150 ;
        RECT 81.445 140.965 81.735 141.010 ;
        RECT 99.370 140.950 99.690 141.010 ;
        RECT 116.850 140.950 117.170 141.210 ;
        RECT 118.690 140.950 119.010 141.210 ;
        RECT 29.840 140.330 127.820 140.810 ;
        RECT 135.580 140.230 136.830 141.220 ;
        RECT 32.210 139.930 32.530 140.190 ;
        RECT 34.985 140.130 35.275 140.175 ;
        RECT 35.430 140.130 35.750 140.190 ;
        RECT 34.985 139.990 35.750 140.130 ;
        RECT 34.985 139.945 35.275 139.990 ;
        RECT 35.430 139.930 35.750 139.990 ;
        RECT 36.825 139.945 37.115 140.175 ;
        RECT 39.570 140.130 39.890 140.190 ;
        RECT 40.045 140.130 40.335 140.175 ;
        RECT 39.570 139.990 40.335 140.130 ;
        RECT 32.685 139.450 32.975 139.495 ;
        RECT 34.525 139.450 34.815 139.495 ;
        RECT 34.970 139.450 35.290 139.510 ;
        RECT 32.685 139.310 33.820 139.450 ;
        RECT 32.685 139.265 32.975 139.310 ;
        RECT 33.680 138.770 33.820 139.310 ;
        RECT 34.525 139.310 35.290 139.450 ;
        RECT 36.900 139.450 37.040 139.945 ;
        RECT 39.570 139.930 39.890 139.990 ;
        RECT 40.045 139.945 40.335 139.990 ;
        RECT 46.010 140.130 46.330 140.190 ;
        RECT 46.010 139.990 50.380 140.130 ;
        RECT 46.010 139.930 46.330 139.990 ;
        RECT 46.470 139.835 46.790 139.850 ;
        RECT 43.730 139.790 44.020 139.835 ;
        RECT 45.590 139.790 45.880 139.835 ;
        RECT 43.730 139.650 45.880 139.790 ;
        RECT 43.730 139.605 44.020 139.650 ;
        RECT 45.590 139.605 45.880 139.650 ;
        RECT 39.125 139.450 39.415 139.495 ;
        RECT 36.900 139.310 39.415 139.450 ;
        RECT 34.525 139.265 34.815 139.310 ;
        RECT 34.970 139.250 35.290 139.310 ;
        RECT 39.125 139.265 39.415 139.310 ;
        RECT 41.425 139.450 41.715 139.495 ;
        RECT 42.330 139.450 42.650 139.510 ;
        RECT 41.425 139.310 42.650 139.450 ;
        RECT 41.425 139.265 41.715 139.310 ;
        RECT 42.330 139.250 42.650 139.310 ;
        RECT 42.790 139.250 43.110 139.510 ;
        RECT 45.665 139.450 45.880 139.605 ;
        RECT 46.470 139.790 46.800 139.835 ;
        RECT 49.770 139.790 50.060 139.835 ;
        RECT 46.470 139.650 50.060 139.790 ;
        RECT 50.240 139.790 50.380 139.990 ;
        RECT 55.225 139.945 55.515 140.175 ;
        RECT 55.670 140.130 55.990 140.190 ;
        RECT 56.605 140.130 56.895 140.175 ;
        RECT 55.670 139.990 56.895 140.130 ;
        RECT 51.070 139.790 51.390 139.850 ;
        RECT 52.465 139.790 52.755 139.835 ;
        RECT 50.240 139.650 52.755 139.790 ;
        RECT 46.470 139.605 46.800 139.650 ;
        RECT 49.770 139.605 50.060 139.650 ;
        RECT 46.470 139.590 46.790 139.605 ;
        RECT 51.070 139.590 51.390 139.650 ;
        RECT 52.465 139.605 52.755 139.650 ;
        RECT 54.290 139.590 54.610 139.850 ;
        RECT 47.910 139.450 48.200 139.495 ;
        RECT 45.665 139.310 48.200 139.450 ;
        RECT 47.910 139.265 48.200 139.310 ;
        RECT 48.770 139.450 49.090 139.510 ;
        RECT 55.300 139.450 55.440 139.945 ;
        RECT 55.670 139.930 55.990 139.990 ;
        RECT 56.605 139.945 56.895 139.990 ;
        RECT 58.430 140.130 58.750 140.190 ;
        RECT 59.365 140.130 59.655 140.175 ;
        RECT 65.790 140.130 66.110 140.190 ;
        RECT 58.430 139.990 59.655 140.130 ;
        RECT 58.430 139.930 58.750 139.990 ;
        RECT 59.365 139.945 59.655 139.990 ;
        RECT 62.200 139.990 66.110 140.130 ;
        RECT 59.810 139.790 60.130 139.850 ;
        RECT 57.600 139.650 59.580 139.790 ;
        RECT 48.770 139.310 55.440 139.450 ;
        RECT 55.670 139.450 55.990 139.510 ;
        RECT 57.600 139.495 57.740 139.650 ;
        RECT 59.440 139.510 59.580 139.650 ;
        RECT 59.810 139.650 61.880 139.790 ;
        RECT 59.810 139.590 60.130 139.650 ;
        RECT 56.145 139.450 56.435 139.495 ;
        RECT 55.670 139.310 56.435 139.450 ;
        RECT 48.770 139.250 49.090 139.310 ;
        RECT 55.670 139.250 55.990 139.310 ;
        RECT 56.145 139.265 56.435 139.310 ;
        RECT 57.525 139.265 57.815 139.495 ;
        RECT 57.970 139.250 58.290 139.510 ;
        RECT 58.890 139.250 59.210 139.510 ;
        RECT 59.350 139.250 59.670 139.510 ;
        RECT 61.740 139.495 61.880 139.650 ;
        RECT 60.745 139.265 61.035 139.495 ;
        RECT 61.205 139.265 61.495 139.495 ;
        RECT 61.665 139.265 61.955 139.495 ;
        RECT 34.050 138.910 34.370 139.170 ;
        RECT 44.645 139.110 44.935 139.155 ;
        RECT 42.420 138.970 44.935 139.110 ;
        RECT 37.270 138.770 37.590 138.830 ;
        RECT 42.420 138.815 42.560 138.970 ;
        RECT 44.645 138.925 44.935 138.970 ;
        RECT 49.690 139.110 50.010 139.170 ;
        RECT 51.775 139.110 52.065 139.155 ;
        RECT 49.690 138.970 52.065 139.110 ;
        RECT 49.690 138.910 50.010 138.970 ;
        RECT 51.775 138.925 52.065 138.970 ;
        RECT 33.680 138.630 37.590 138.770 ;
        RECT 37.270 138.570 37.590 138.630 ;
        RECT 42.345 138.585 42.635 138.815 ;
        RECT 43.270 138.770 43.560 138.815 ;
        RECT 45.130 138.770 45.420 138.815 ;
        RECT 47.910 138.770 48.200 138.815 ;
        RECT 43.270 138.630 48.200 138.770 ;
        RECT 43.270 138.585 43.560 138.630 ;
        RECT 45.130 138.585 45.420 138.630 ;
        RECT 47.910 138.585 48.200 138.630 ;
        RECT 58.430 138.230 58.750 138.490 ;
        RECT 60.820 138.430 60.960 139.265 ;
        RECT 61.280 139.110 61.420 139.265 ;
        RECT 62.200 139.110 62.340 139.990 ;
        RECT 65.790 139.930 66.110 139.990 ;
        RECT 66.265 140.130 66.555 140.175 ;
        RECT 69.010 140.130 69.330 140.190 ;
        RECT 66.265 139.990 69.330 140.130 ;
        RECT 66.265 139.945 66.555 139.990 ;
        RECT 69.010 139.930 69.330 139.990 ;
        RECT 75.450 140.130 75.770 140.190 ;
        RECT 75.450 139.990 81.660 140.130 ;
        RECT 75.450 139.930 75.770 139.990 ;
        RECT 72.690 139.835 73.010 139.850 ;
        RECT 63.965 139.790 64.255 139.835 ;
        RECT 66.725 139.790 67.015 139.835 ;
        RECT 72.640 139.790 73.010 139.835 ;
        RECT 75.900 139.790 76.190 139.835 ;
        RECT 63.965 139.650 67.015 139.790 ;
        RECT 63.965 139.605 64.255 139.650 ;
        RECT 66.725 139.605 67.015 139.650 ;
        RECT 67.720 139.650 70.160 139.790 ;
        RECT 62.585 139.265 62.875 139.495 ;
        RECT 61.280 138.970 62.340 139.110 ;
        RECT 62.660 138.770 62.800 139.265 ;
        RECT 65.330 139.250 65.650 139.510 ;
        RECT 64.885 139.110 65.175 139.155 ;
        RECT 66.250 139.110 66.570 139.170 ;
        RECT 64.885 138.970 66.570 139.110 ;
        RECT 64.885 138.925 65.175 138.970 ;
        RECT 66.250 138.910 66.570 138.970 ;
        RECT 67.170 138.770 67.490 138.830 ;
        RECT 67.720 138.770 67.860 139.650 ;
        RECT 70.020 139.510 70.160 139.650 ;
        RECT 72.640 139.650 76.190 139.790 ;
        RECT 72.640 139.605 73.010 139.650 ;
        RECT 75.900 139.605 76.190 139.650 ;
        RECT 76.820 139.790 77.110 139.835 ;
        RECT 78.680 139.790 78.970 139.835 ;
        RECT 76.820 139.650 78.970 139.790 ;
        RECT 76.820 139.605 77.110 139.650 ;
        RECT 78.680 139.605 78.970 139.650 ;
        RECT 72.690 139.590 73.010 139.605 ;
        RECT 68.090 139.250 68.410 139.510 ;
        RECT 68.565 139.265 68.855 139.495 ;
        RECT 69.025 139.265 69.315 139.495 ;
        RECT 68.640 139.110 68.780 139.265 ;
        RECT 62.660 138.630 67.860 138.770 ;
        RECT 68.410 138.970 68.780 139.110 ;
        RECT 67.170 138.570 67.490 138.630 ;
        RECT 63.950 138.430 64.270 138.490 ;
        RECT 60.820 138.290 64.270 138.430 ;
        RECT 63.950 138.230 64.270 138.290 ;
        RECT 65.330 138.230 65.650 138.490 ;
        RECT 65.790 138.430 66.110 138.490 ;
        RECT 67.630 138.430 67.950 138.490 ;
        RECT 68.410 138.430 68.550 138.970 ;
        RECT 65.790 138.290 68.550 138.430 ;
        RECT 69.100 138.430 69.240 139.265 ;
        RECT 69.930 139.250 70.250 139.510 ;
        RECT 74.500 139.450 74.790 139.495 ;
        RECT 76.820 139.450 77.035 139.605 ;
        RECT 80.510 139.590 80.830 139.850 ;
        RECT 81.520 139.790 81.660 139.990 ;
        RECT 93.405 139.945 93.695 140.175 ;
        RECT 93.480 139.790 93.620 139.945 ;
        RECT 94.770 139.930 95.090 140.190 ;
        RECT 95.705 140.130 95.995 140.175 ;
        RECT 96.150 140.130 96.470 140.190 ;
        RECT 95.705 139.990 96.470 140.130 ;
        RECT 95.705 139.945 95.995 139.990 ;
        RECT 96.150 139.930 96.470 139.990 ;
        RECT 105.350 140.130 105.670 140.190 ;
        RECT 108.125 140.130 108.415 140.175 ;
        RECT 135.635 140.155 136.775 140.230 ;
        RECT 105.350 139.990 108.415 140.130 ;
        RECT 105.350 139.930 105.670 139.990 ;
        RECT 108.125 139.945 108.415 139.990 ;
        RECT 96.610 139.790 96.930 139.850 ;
        RECT 106.730 139.790 107.050 139.850 ;
        RECT 110.425 139.790 110.715 139.835 ;
        RECT 81.520 139.650 92.240 139.790 ;
        RECT 93.480 139.650 96.930 139.790 ;
        RECT 74.500 139.310 77.035 139.450 ;
        RECT 77.290 139.450 77.610 139.510 ;
        RECT 77.765 139.450 78.055 139.495 ;
        RECT 77.290 139.310 78.055 139.450 ;
        RECT 74.500 139.265 74.790 139.310 ;
        RECT 77.290 139.250 77.610 139.310 ;
        RECT 77.765 139.265 78.055 139.310 ;
        RECT 86.030 139.450 86.350 139.510 ;
        RECT 87.325 139.450 87.615 139.495 ;
        RECT 86.030 139.310 87.615 139.450 ;
        RECT 86.030 139.250 86.350 139.310 ;
        RECT 87.325 139.265 87.615 139.310 ;
        RECT 75.450 139.110 75.770 139.170 ;
        RECT 79.605 139.110 79.895 139.155 ;
        RECT 75.450 138.970 79.895 139.110 ;
        RECT 75.450 138.910 75.770 138.970 ;
        RECT 79.605 138.925 79.895 138.970 ;
        RECT 86.490 138.910 86.810 139.170 ;
        RECT 88.345 139.110 88.635 139.155 ;
        RECT 90.630 139.110 90.950 139.170 ;
        RECT 88.345 138.970 90.950 139.110 ;
        RECT 92.100 139.110 92.240 139.650 ;
        RECT 96.610 139.590 96.930 139.650 ;
        RECT 98.080 139.650 105.120 139.790 ;
        RECT 92.485 139.450 92.775 139.495 ;
        RECT 93.390 139.450 93.710 139.510 ;
        RECT 92.485 139.310 93.710 139.450 ;
        RECT 92.485 139.265 92.775 139.310 ;
        RECT 93.390 139.250 93.710 139.310 ;
        RECT 93.865 139.450 94.155 139.495 ;
        RECT 94.310 139.450 94.630 139.510 ;
        RECT 93.865 139.310 94.630 139.450 ;
        RECT 93.865 139.265 94.155 139.310 ;
        RECT 94.310 139.250 94.630 139.310 ;
        RECT 95.230 139.450 95.550 139.510 ;
        RECT 98.080 139.495 98.220 139.650 ;
        RECT 96.165 139.450 96.455 139.495 ;
        RECT 98.005 139.450 98.295 139.495 ;
        RECT 95.230 139.310 96.455 139.450 ;
        RECT 95.230 139.250 95.550 139.310 ;
        RECT 96.165 139.265 96.455 139.310 ;
        RECT 96.700 139.310 98.295 139.450 ;
        RECT 96.700 139.110 96.840 139.310 ;
        RECT 98.005 139.265 98.295 139.310 ;
        RECT 101.685 139.450 101.975 139.495 ;
        RECT 102.130 139.450 102.450 139.510 ;
        RECT 104.980 139.495 105.120 139.650 ;
        RECT 106.730 139.650 110.715 139.790 ;
        RECT 106.730 139.590 107.050 139.650 ;
        RECT 110.425 139.605 110.715 139.650 ;
        RECT 115.010 139.790 115.330 139.850 ;
        RECT 119.100 139.790 119.390 139.835 ;
        RECT 122.360 139.790 122.650 139.835 ;
        RECT 115.010 139.650 122.650 139.790 ;
        RECT 115.010 139.590 115.330 139.650 ;
        RECT 119.100 139.605 119.390 139.650 ;
        RECT 122.360 139.605 122.650 139.650 ;
        RECT 123.280 139.790 123.570 139.835 ;
        RECT 125.140 139.790 125.430 139.835 ;
        RECT 123.280 139.650 125.430 139.790 ;
        RECT 123.280 139.605 123.570 139.650 ;
        RECT 125.140 139.605 125.430 139.650 ;
        RECT 101.685 139.310 102.450 139.450 ;
        RECT 101.685 139.265 101.975 139.310 ;
        RECT 102.130 139.250 102.450 139.310 ;
        RECT 104.905 139.450 105.195 139.495 ;
        RECT 107.205 139.450 107.495 139.495 ;
        RECT 108.570 139.450 108.890 139.510 ;
        RECT 104.905 139.310 108.890 139.450 ;
        RECT 104.905 139.265 105.195 139.310 ;
        RECT 107.205 139.265 107.495 139.310 ;
        RECT 108.570 139.250 108.890 139.310 ;
        RECT 109.965 139.450 110.255 139.495 ;
        RECT 110.870 139.450 111.190 139.510 ;
        RECT 109.965 139.310 111.190 139.450 ;
        RECT 109.965 139.265 110.255 139.310 ;
        RECT 110.870 139.250 111.190 139.310 ;
        RECT 120.960 139.450 121.250 139.495 ;
        RECT 123.280 139.450 123.495 139.605 ;
        RECT 120.960 139.310 123.495 139.450 ;
        RECT 120.960 139.265 121.250 139.310 ;
        RECT 129.090 139.190 134.150 139.405 ;
        RECT 143.370 139.390 144.510 223.840 ;
        RECT 137.240 139.380 144.510 139.390 ;
        RECT 136.210 139.190 144.510 139.380 ;
        RECT 92.100 138.970 96.840 139.110 ;
        RECT 88.345 138.925 88.635 138.970 ;
        RECT 90.630 138.910 90.950 138.970 ;
        RECT 97.085 138.925 97.375 139.155 ;
        RECT 98.925 139.110 99.215 139.155 ;
        RECT 99.830 139.110 100.150 139.170 ;
        RECT 98.925 138.970 100.150 139.110 ;
        RECT 98.925 138.925 99.215 138.970 ;
        RECT 74.500 138.770 74.790 138.815 ;
        RECT 77.280 138.770 77.570 138.815 ;
        RECT 79.140 138.770 79.430 138.815 ;
        RECT 74.500 138.630 79.430 138.770 ;
        RECT 97.160 138.770 97.300 138.925 ;
        RECT 99.830 138.910 100.150 138.970 ;
        RECT 103.985 138.925 104.275 139.155 ;
        RECT 97.160 138.630 99.140 138.770 ;
        RECT 74.500 138.585 74.790 138.630 ;
        RECT 77.280 138.585 77.570 138.630 ;
        RECT 79.140 138.585 79.430 138.630 ;
        RECT 99.000 138.490 99.140 138.630 ;
        RECT 70.635 138.430 70.925 138.475 ;
        RECT 73.150 138.430 73.470 138.490 ;
        RECT 69.100 138.290 73.470 138.430 ;
        RECT 65.790 138.230 66.110 138.290 ;
        RECT 67.630 138.230 67.950 138.290 ;
        RECT 70.635 138.245 70.925 138.290 ;
        RECT 73.150 138.230 73.470 138.290 ;
        RECT 81.905 138.430 82.195 138.475 ;
        RECT 83.270 138.430 83.590 138.490 ;
        RECT 81.905 138.290 83.590 138.430 ;
        RECT 81.905 138.245 82.195 138.290 ;
        RECT 83.270 138.230 83.590 138.290 ;
        RECT 98.910 138.230 99.230 138.490 ;
        RECT 104.060 138.430 104.200 138.925 ;
        RECT 105.810 138.910 106.130 139.170 ;
        RECT 106.285 139.110 106.575 139.155 ;
        RECT 109.030 139.110 109.350 139.170 ;
        RECT 106.285 138.970 109.350 139.110 ;
        RECT 106.285 138.925 106.575 138.970 ;
        RECT 109.030 138.910 109.350 138.970 ;
        RECT 109.505 139.110 109.795 139.155 ;
        RECT 113.170 139.110 113.490 139.170 ;
        RECT 109.505 138.970 113.490 139.110 ;
        RECT 109.505 138.925 109.795 138.970 ;
        RECT 113.170 138.910 113.490 138.970 ;
        RECT 124.210 138.910 124.530 139.170 ;
        RECT 126.050 138.910 126.370 139.170 ;
        RECT 116.850 138.815 117.170 138.830 ;
        RECT 116.850 138.770 117.385 138.815 ;
        RECT 111.880 138.630 117.385 138.770 ;
        RECT 111.880 138.430 112.020 138.630 ;
        RECT 116.850 138.585 117.385 138.630 ;
        RECT 120.960 138.770 121.250 138.815 ;
        RECT 123.740 138.770 124.030 138.815 ;
        RECT 125.600 138.770 125.890 138.815 ;
        RECT 120.960 138.630 125.890 138.770 ;
        RECT 120.960 138.585 121.250 138.630 ;
        RECT 123.740 138.585 124.030 138.630 ;
        RECT 125.600 138.585 125.890 138.630 ;
        RECT 116.850 138.570 117.170 138.585 ;
        RECT 104.060 138.290 112.020 138.430 ;
        RECT 112.250 138.230 112.570 138.490 ;
        RECT 112.710 138.430 113.030 138.490 ;
        RECT 126.140 138.430 126.280 138.910 ;
        RECT 112.710 138.290 126.280 138.430 ;
        RECT 129.090 138.530 144.510 139.190 ;
        RECT 112.710 138.230 113.030 138.290 ;
        RECT 129.090 138.225 134.150 138.530 ;
        RECT 136.210 138.250 144.510 138.530 ;
        RECT 136.210 138.240 138.350 138.250 ;
        RECT 29.840 137.610 127.820 138.090 ;
        RECT 40.735 137.410 41.025 137.455 ;
        RECT 50.150 137.410 50.470 137.470 ;
        RECT 40.735 137.270 50.470 137.410 ;
        RECT 40.735 137.225 41.025 137.270 ;
        RECT 50.150 137.210 50.470 137.270 ;
        RECT 54.305 137.410 54.595 137.455 ;
        RECT 55.670 137.410 55.990 137.470 ;
        RECT 54.305 137.270 55.990 137.410 ;
        RECT 54.305 137.225 54.595 137.270 ;
        RECT 55.670 137.210 55.990 137.270 ;
        RECT 56.590 137.410 56.910 137.470 ;
        RECT 57.065 137.410 57.355 137.455 ;
        RECT 56.590 137.270 57.355 137.410 ;
        RECT 56.590 137.210 56.910 137.270 ;
        RECT 57.065 137.225 57.355 137.270 ;
        RECT 80.050 137.410 80.370 137.470 ;
        RECT 80.525 137.410 80.815 137.455 ;
        RECT 80.050 137.270 80.815 137.410 ;
        RECT 80.050 137.210 80.370 137.270 ;
        RECT 80.525 137.225 80.815 137.270 ;
        RECT 82.810 137.210 83.130 137.470 ;
        RECT 83.730 137.410 84.050 137.470 ;
        RECT 85.125 137.410 85.415 137.455 ;
        RECT 83.730 137.270 85.415 137.410 ;
        RECT 83.730 137.210 84.050 137.270 ;
        RECT 85.125 137.225 85.415 137.270 ;
        RECT 95.230 137.410 95.550 137.470 ;
        RECT 109.950 137.410 110.270 137.470 ;
        RECT 95.230 137.270 114.780 137.410 ;
        RECT 95.230 137.210 95.550 137.270 ;
        RECT 44.600 137.070 44.890 137.115 ;
        RECT 47.380 137.070 47.670 137.115 ;
        RECT 49.240 137.070 49.530 137.115 ;
        RECT 44.600 136.930 49.530 137.070 ;
        RECT 44.600 136.885 44.890 136.930 ;
        RECT 47.380 136.885 47.670 136.930 ;
        RECT 49.240 136.885 49.530 136.930 ;
        RECT 53.370 137.070 53.690 137.130 ;
        RECT 75.910 137.070 76.230 137.130 ;
        RECT 53.370 136.930 76.230 137.070 ;
        RECT 53.370 136.870 53.690 136.930 ;
        RECT 47.865 136.730 48.155 136.775 ;
        RECT 48.770 136.730 49.090 136.790 ;
        RECT 47.865 136.590 49.090 136.730 ;
        RECT 47.865 136.545 48.155 136.590 ;
        RECT 48.770 136.530 49.090 136.590 ;
        RECT 50.150 136.530 50.470 136.790 ;
        RECT 51.070 136.530 51.390 136.790 ;
        RECT 51.990 136.730 52.310 136.790 ;
        RECT 55.670 136.730 55.990 136.790 ;
        RECT 51.990 136.590 55.990 136.730 ;
        RECT 51.990 136.530 52.310 136.590 ;
        RECT 55.670 136.530 55.990 136.590 ;
        RECT 37.270 136.390 37.590 136.450 ;
        RECT 39.125 136.390 39.415 136.435 ;
        RECT 37.270 136.250 39.415 136.390 ;
        RECT 37.270 136.190 37.590 136.250 ;
        RECT 39.125 136.205 39.415 136.250 ;
        RECT 44.600 136.390 44.890 136.435 ;
        RECT 44.600 136.250 47.135 136.390 ;
        RECT 44.600 136.205 44.890 136.250 ;
        RECT 46.920 136.095 47.135 136.250 ;
        RECT 49.705 136.205 49.995 136.435 ;
        RECT 50.240 136.390 50.380 136.530 ;
        RECT 52.450 136.390 52.770 136.450 ;
        RECT 50.240 136.250 52.770 136.390 ;
        RECT 39.585 136.050 39.875 136.095 ;
        RECT 42.740 136.050 43.030 136.095 ;
        RECT 46.000 136.050 46.290 136.095 ;
        RECT 39.585 135.910 46.290 136.050 ;
        RECT 39.585 135.865 39.875 135.910 ;
        RECT 42.740 135.865 43.030 135.910 ;
        RECT 46.000 135.865 46.290 135.910 ;
        RECT 46.920 136.050 47.210 136.095 ;
        RECT 48.780 136.050 49.070 136.095 ;
        RECT 46.920 135.910 49.070 136.050 ;
        RECT 49.780 136.050 49.920 136.205 ;
        RECT 52.450 136.190 52.770 136.250 ;
        RECT 52.910 136.390 53.230 136.450 ;
        RECT 56.220 136.435 56.360 136.930 ;
        RECT 75.910 136.870 76.230 136.930 ;
        RECT 83.270 137.070 83.590 137.130 ;
        RECT 83.270 136.930 97.760 137.070 ;
        RECT 83.270 136.870 83.590 136.930 ;
        RECT 69.930 136.730 70.250 136.790 ;
        RECT 70.865 136.730 71.155 136.775 ;
        RECT 71.770 136.730 72.090 136.790 ;
        RECT 69.930 136.590 72.090 136.730 ;
        RECT 69.930 136.530 70.250 136.590 ;
        RECT 70.865 136.545 71.155 136.590 ;
        RECT 71.770 136.530 72.090 136.590 ;
        RECT 55.225 136.390 55.515 136.435 ;
        RECT 52.910 136.250 55.515 136.390 ;
        RECT 52.910 136.190 53.230 136.250 ;
        RECT 55.225 136.205 55.515 136.250 ;
        RECT 56.145 136.390 56.435 136.435 ;
        RECT 57.050 136.390 57.370 136.450 ;
        RECT 56.145 136.250 57.370 136.390 ;
        RECT 56.145 136.205 56.435 136.250 ;
        RECT 57.050 136.190 57.370 136.250 ;
        RECT 64.410 136.390 64.730 136.450 ;
        RECT 66.265 136.390 66.555 136.435 ;
        RECT 64.410 136.250 66.555 136.390 ;
        RECT 64.410 136.190 64.730 136.250 ;
        RECT 66.265 136.205 66.555 136.250 ;
        RECT 72.245 136.390 72.535 136.435 ;
        RECT 73.150 136.390 73.470 136.450 ;
        RECT 72.245 136.250 73.470 136.390 ;
        RECT 76.000 136.390 76.140 136.870 ;
        RECT 97.620 136.775 97.760 136.930 ;
        RECT 81.520 136.590 85.110 136.730 ;
        RECT 81.520 136.435 81.660 136.590 ;
        RECT 81.445 136.390 81.735 136.435 ;
        RECT 76.000 136.250 81.735 136.390 ;
        RECT 72.245 136.205 72.535 136.250 ;
        RECT 73.150 136.190 73.470 136.250 ;
        RECT 81.445 136.205 81.735 136.250 ;
        RECT 81.890 136.190 82.210 136.450 ;
        RECT 83.820 136.435 83.960 136.590 ;
        RECT 83.745 136.205 84.035 136.435 ;
        RECT 84.190 136.190 84.510 136.450 ;
        RECT 84.970 136.390 85.110 136.590 ;
        RECT 97.545 136.545 97.835 136.775 ;
        RECT 86.030 136.390 86.350 136.450 ;
        RECT 84.970 136.250 86.350 136.390 ;
        RECT 86.030 136.190 86.350 136.250 ;
        RECT 86.490 136.190 86.810 136.450 ;
        RECT 87.870 136.190 88.190 136.450 ;
        RECT 102.220 136.435 102.360 137.270 ;
        RECT 109.950 137.210 110.270 137.270 ;
        RECT 107.620 137.070 107.910 137.115 ;
        RECT 110.400 137.070 110.690 137.115 ;
        RECT 112.260 137.070 112.550 137.115 ;
        RECT 107.620 136.930 112.550 137.070 ;
        RECT 107.620 136.885 107.910 136.930 ;
        RECT 110.400 136.885 110.690 136.930 ;
        RECT 112.260 136.885 112.550 136.930 ;
        RECT 113.185 136.885 113.475 137.115 ;
        RECT 105.350 136.730 105.670 136.790 ;
        RECT 112.710 136.730 113.030 136.790 ;
        RECT 105.350 136.590 113.030 136.730 ;
        RECT 105.350 136.530 105.670 136.590 ;
        RECT 112.710 136.530 113.030 136.590 ;
        RECT 98.925 136.205 99.215 136.435 ;
        RECT 102.145 136.205 102.435 136.435 ;
        RECT 107.620 136.390 107.910 136.435 ;
        RECT 110.885 136.390 111.175 136.435 ;
        RECT 113.260 136.390 113.400 136.885 ;
        RECT 114.640 136.435 114.780 137.270 ;
        RECT 115.010 137.210 115.330 137.470 ;
        RECT 120.040 137.070 120.330 137.115 ;
        RECT 122.820 137.070 123.110 137.115 ;
        RECT 124.680 137.070 124.970 137.115 ;
        RECT 120.040 136.930 124.970 137.070 ;
        RECT 120.040 136.885 120.330 136.930 ;
        RECT 122.820 136.885 123.110 136.930 ;
        RECT 124.680 136.885 124.970 136.930 ;
        RECT 107.620 136.250 110.155 136.390 ;
        RECT 107.620 136.205 107.910 136.250 ;
        RECT 50.150 136.050 50.470 136.110 ;
        RECT 57.525 136.050 57.815 136.095 ;
        RECT 49.780 135.910 57.815 136.050 ;
        RECT 86.580 136.050 86.720 136.190 ;
        RECT 99.000 136.050 99.140 136.205 ;
        RECT 109.940 136.095 110.155 136.250 ;
        RECT 110.885 136.250 113.400 136.390 ;
        RECT 110.885 136.205 111.175 136.250 ;
        RECT 114.105 136.205 114.395 136.435 ;
        RECT 114.565 136.390 114.855 136.435 ;
        RECT 119.150 136.390 119.470 136.450 ;
        RECT 114.565 136.250 119.470 136.390 ;
        RECT 114.565 136.205 114.855 136.250 ;
        RECT 86.580 135.910 99.140 136.050 ;
        RECT 102.605 136.050 102.895 136.095 ;
        RECT 105.760 136.050 106.050 136.095 ;
        RECT 109.020 136.050 109.310 136.095 ;
        RECT 102.605 135.910 109.310 136.050 ;
        RECT 46.920 135.865 47.210 135.910 ;
        RECT 48.780 135.865 49.070 135.910 ;
        RECT 50.150 135.850 50.470 135.910 ;
        RECT 57.525 135.865 57.815 135.910 ;
        RECT 102.605 135.865 102.895 135.910 ;
        RECT 105.760 135.865 106.050 135.910 ;
        RECT 109.020 135.865 109.310 135.910 ;
        RECT 109.940 136.050 110.230 136.095 ;
        RECT 111.800 136.050 112.090 136.095 ;
        RECT 109.940 135.910 112.090 136.050 ;
        RECT 109.940 135.865 110.230 135.910 ;
        RECT 111.800 135.865 112.090 135.910 ;
        RECT 112.250 136.050 112.570 136.110 ;
        RECT 114.180 136.050 114.320 136.205 ;
        RECT 119.150 136.190 119.470 136.250 ;
        RECT 120.040 136.390 120.330 136.435 ;
        RECT 122.830 136.390 123.150 136.450 ;
        RECT 123.305 136.390 123.595 136.435 ;
        RECT 120.040 136.250 122.575 136.390 ;
        RECT 120.040 136.205 120.330 136.250 ;
        RECT 112.250 135.910 114.320 136.050 ;
        RECT 118.180 136.050 118.470 136.095 ;
        RECT 119.610 136.050 119.930 136.110 ;
        RECT 122.360 136.095 122.575 136.250 ;
        RECT 122.830 136.250 123.595 136.390 ;
        RECT 122.830 136.190 123.150 136.250 ;
        RECT 123.305 136.205 123.595 136.250 ;
        RECT 125.130 136.190 125.450 136.450 ;
        RECT 121.440 136.050 121.730 136.095 ;
        RECT 118.180 135.910 121.730 136.050 ;
        RECT 112.250 135.850 112.570 135.910 ;
        RECT 118.180 135.865 118.470 135.910 ;
        RECT 119.610 135.850 119.930 135.910 ;
        RECT 121.440 135.865 121.730 135.910 ;
        RECT 122.360 136.050 122.650 136.095 ;
        RECT 124.220 136.050 124.510 136.095 ;
        RECT 122.360 135.910 124.510 136.050 ;
        RECT 122.360 135.865 122.650 135.910 ;
        RECT 124.220 135.865 124.510 135.910 ;
        RECT 34.970 135.710 35.290 135.770 ;
        RECT 52.910 135.710 53.230 135.770 ;
        RECT 34.970 135.570 53.230 135.710 ;
        RECT 34.970 135.510 35.290 135.570 ;
        RECT 52.910 135.510 53.230 135.570 ;
        RECT 70.850 135.710 71.170 135.770 ;
        RECT 71.785 135.710 72.075 135.755 ;
        RECT 70.850 135.570 72.075 135.710 ;
        RECT 70.850 135.510 71.170 135.570 ;
        RECT 71.785 135.525 72.075 135.570 ;
        RECT 74.085 135.710 74.375 135.755 ;
        RECT 74.530 135.710 74.850 135.770 ;
        RECT 74.085 135.570 74.850 135.710 ;
        RECT 74.085 135.525 74.375 135.570 ;
        RECT 74.530 135.510 74.850 135.570 ;
        RECT 95.230 135.510 95.550 135.770 ;
        RECT 98.465 135.710 98.755 135.755 ;
        RECT 98.910 135.710 99.230 135.770 ;
        RECT 98.465 135.570 99.230 135.710 ;
        RECT 98.465 135.525 98.755 135.570 ;
        RECT 98.910 135.510 99.230 135.570 ;
        RECT 100.290 135.710 100.610 135.770 ;
        RECT 100.765 135.710 101.055 135.755 ;
        RECT 100.290 135.570 101.055 135.710 ;
        RECT 100.290 135.510 100.610 135.570 ;
        RECT 100.765 135.525 101.055 135.570 ;
        RECT 103.755 135.710 104.045 135.755 ;
        RECT 106.270 135.710 106.590 135.770 ;
        RECT 103.755 135.570 106.590 135.710 ;
        RECT 103.755 135.525 104.045 135.570 ;
        RECT 106.270 135.510 106.590 135.570 ;
        RECT 110.870 135.710 111.190 135.770 ;
        RECT 116.175 135.710 116.465 135.755 ;
        RECT 116.850 135.710 117.170 135.770 ;
        RECT 110.870 135.570 117.170 135.710 ;
        RECT 110.870 135.510 111.190 135.570 ;
        RECT 116.175 135.525 116.465 135.570 ;
        RECT 116.850 135.510 117.170 135.570 ;
        RECT 29.840 134.890 127.820 135.370 ;
        RECT 34.970 134.490 35.290 134.750 ;
        RECT 35.430 134.490 35.750 134.750 ;
        RECT 43.250 134.690 43.570 134.750 ;
        RECT 46.715 134.690 47.005 134.735 ;
        RECT 51.990 134.690 52.310 134.750 ;
        RECT 43.250 134.550 45.320 134.690 ;
        RECT 43.250 134.490 43.570 134.550 ;
        RECT 41.410 134.395 41.730 134.410 ;
        RECT 38.670 134.350 38.960 134.395 ;
        RECT 40.530 134.350 40.820 134.395 ;
        RECT 38.670 134.210 40.820 134.350 ;
        RECT 38.670 134.165 38.960 134.210 ;
        RECT 40.530 134.165 40.820 134.210 ;
        RECT 39.570 133.810 39.890 134.070 ;
        RECT 40.605 134.010 40.820 134.165 ;
        RECT 41.410 134.350 41.740 134.395 ;
        RECT 44.710 134.350 45.000 134.395 ;
        RECT 41.410 134.210 45.000 134.350 ;
        RECT 41.410 134.165 41.740 134.210 ;
        RECT 44.710 134.165 45.000 134.210 ;
        RECT 41.410 134.150 41.730 134.165 ;
        RECT 42.850 134.010 43.140 134.055 ;
        RECT 40.605 133.870 43.140 134.010 ;
        RECT 45.180 134.010 45.320 134.550 ;
        RECT 46.715 134.550 52.310 134.690 ;
        RECT 46.715 134.505 47.005 134.550 ;
        RECT 51.990 134.490 52.310 134.550 ;
        RECT 52.910 134.690 53.230 134.750 ;
        RECT 56.375 134.690 56.665 134.735 ;
        RECT 52.910 134.550 56.665 134.690 ;
        RECT 52.910 134.490 53.230 134.550 ;
        RECT 56.375 134.505 56.665 134.550 ;
        RECT 58.890 134.690 59.210 134.750 ;
        RECT 63.965 134.690 64.255 134.735 ;
        RECT 68.090 134.690 68.410 134.750 ;
        RECT 58.890 134.550 64.255 134.690 ;
        RECT 58.890 134.490 59.210 134.550 ;
        RECT 63.965 134.505 64.255 134.550 ;
        RECT 64.500 134.550 68.410 134.690 ;
        RECT 48.330 134.350 48.620 134.395 ;
        RECT 50.190 134.350 50.480 134.395 ;
        RECT 48.330 134.210 50.480 134.350 ;
        RECT 48.330 134.165 48.620 134.210 ;
        RECT 50.190 134.165 50.480 134.210 ;
        RECT 51.110 134.350 51.400 134.395 ;
        RECT 54.370 134.350 54.660 134.395 ;
        RECT 51.110 134.210 54.660 134.350 ;
        RECT 51.110 134.165 51.400 134.210 ;
        RECT 49.245 134.010 49.535 134.055 ;
        RECT 45.180 133.870 49.535 134.010 ;
        RECT 50.265 134.010 50.480 134.165 ;
        RECT 52.510 134.010 52.800 134.055 ;
        RECT 50.265 133.870 52.800 134.010 ;
        RECT 42.850 133.825 43.140 133.870 ;
        RECT 49.245 133.825 49.535 133.870 ;
        RECT 52.510 133.825 52.800 133.870 ;
        RECT 34.050 133.670 34.370 133.730 ;
        RECT 35.890 133.670 36.210 133.730 ;
        RECT 34.050 133.530 36.210 133.670 ;
        RECT 34.050 133.470 34.370 133.530 ;
        RECT 35.890 133.470 36.210 133.530 ;
        RECT 37.745 133.670 38.035 133.715 ;
        RECT 44.170 133.670 44.490 133.730 ;
        RECT 47.405 133.670 47.695 133.715 ;
        RECT 50.150 133.670 50.470 133.730 ;
        RECT 37.745 133.530 50.470 133.670 ;
        RECT 37.745 133.485 38.035 133.530 ;
        RECT 44.170 133.470 44.490 133.530 ;
        RECT 47.405 133.485 47.695 133.530 ;
        RECT 50.150 133.470 50.470 133.530 ;
        RECT 38.210 133.330 38.500 133.375 ;
        RECT 40.070 133.330 40.360 133.375 ;
        RECT 42.850 133.330 43.140 133.375 ;
        RECT 38.210 133.190 43.140 133.330 ;
        RECT 38.210 133.145 38.500 133.190 ;
        RECT 40.070 133.145 40.360 133.190 ;
        RECT 42.850 133.145 43.140 133.190 ;
        RECT 47.870 133.330 48.160 133.375 ;
        RECT 49.730 133.330 50.020 133.375 ;
        RECT 52.510 133.330 52.800 133.375 ;
        RECT 47.870 133.190 52.800 133.330 ;
        RECT 47.870 133.145 48.160 133.190 ;
        RECT 49.730 133.145 50.020 133.190 ;
        RECT 52.510 133.145 52.800 133.190 ;
        RECT 33.145 132.990 33.435 133.035 ;
        RECT 34.050 132.990 34.370 133.050 ;
        RECT 33.145 132.850 34.370 132.990 ;
        RECT 33.145 132.805 33.435 132.850 ;
        RECT 34.050 132.790 34.370 132.850 ;
        RECT 35.430 132.990 35.750 133.050 ;
        RECT 53.000 132.990 53.140 134.210 ;
        RECT 54.370 134.165 54.660 134.210 ;
        RECT 60.270 134.150 60.590 134.410 ;
        RECT 57.050 134.010 57.370 134.070 ;
        RECT 58.905 134.010 59.195 134.055 ;
        RECT 57.050 133.870 59.195 134.010 ;
        RECT 57.050 133.810 57.370 133.870 ;
        RECT 58.905 133.825 59.195 133.870 ;
        RECT 61.650 133.810 61.970 134.070 ;
        RECT 63.950 134.010 64.270 134.070 ;
        RECT 64.500 134.010 64.640 134.550 ;
        RECT 68.090 134.490 68.410 134.550 ;
        RECT 81.890 134.690 82.210 134.750 ;
        RECT 85.125 134.690 85.415 134.735 ;
        RECT 90.645 134.690 90.935 134.735 ;
        RECT 81.890 134.550 90.935 134.690 ;
        RECT 81.890 134.490 82.210 134.550 ;
        RECT 85.125 134.505 85.415 134.550 ;
        RECT 90.645 134.505 90.935 134.550 ;
        RECT 92.945 134.690 93.235 134.735 ;
        RECT 93.850 134.690 94.170 134.750 ;
        RECT 92.945 134.550 94.170 134.690 ;
        RECT 92.945 134.505 93.235 134.550 ;
        RECT 93.850 134.490 94.170 134.550 ;
        RECT 96.395 134.690 96.685 134.735 ;
        RECT 98.910 134.690 99.230 134.750 ;
        RECT 107.665 134.690 107.955 134.735 ;
        RECT 96.395 134.550 107.955 134.690 ;
        RECT 96.395 134.505 96.685 134.550 ;
        RECT 98.910 134.490 99.230 134.550 ;
        RECT 107.665 134.505 107.955 134.550 ;
        RECT 116.390 134.490 116.710 134.750 ;
        RECT 116.850 134.490 117.170 134.750 ;
        RECT 119.610 134.490 119.930 134.750 ;
        RECT 121.925 134.690 122.215 134.735 ;
        RECT 122.830 134.690 123.150 134.750 ;
        RECT 121.925 134.550 123.150 134.690 ;
        RECT 121.925 134.505 122.215 134.550 ;
        RECT 122.830 134.490 123.150 134.550 ;
        RECT 123.305 134.690 123.595 134.735 ;
        RECT 124.210 134.690 124.530 134.750 ;
        RECT 123.305 134.550 124.530 134.690 ;
        RECT 123.305 134.505 123.595 134.550 ;
        RECT 124.210 134.490 124.530 134.550 ;
        RECT 135.660 134.480 136.800 134.510 ;
        RECT 64.870 134.350 65.190 134.410 ;
        RECT 70.405 134.350 70.695 134.395 ;
        RECT 64.870 134.210 70.695 134.350 ;
        RECT 64.870 134.150 65.190 134.210 ;
        RECT 65.345 134.010 65.635 134.055 ;
        RECT 63.950 133.870 65.635 134.010 ;
        RECT 63.950 133.810 64.270 133.870 ;
        RECT 65.345 133.825 65.635 133.870 ;
        RECT 65.790 133.810 66.110 134.070 ;
        RECT 66.340 134.055 66.480 134.210 ;
        RECT 70.405 134.165 70.695 134.210 ;
        RECT 74.990 134.350 75.310 134.410 ;
        RECT 101.670 134.395 101.990 134.410 ;
        RECT 98.400 134.350 98.690 134.395 ;
        RECT 101.660 134.350 101.990 134.395 ;
        RECT 74.990 134.210 80.740 134.350 ;
        RECT 74.990 134.150 75.310 134.210 ;
        RECT 66.265 133.825 66.555 134.055 ;
        RECT 67.170 133.810 67.490 134.070 ;
        RECT 67.645 134.010 67.935 134.055 ;
        RECT 67.645 133.870 70.620 134.010 ;
        RECT 67.645 133.825 67.935 133.870 ;
        RECT 70.480 133.730 70.620 133.870 ;
        RECT 70.850 133.810 71.170 134.070 ;
        RECT 74.085 133.825 74.375 134.055 ;
        RECT 74.530 134.010 74.850 134.070 ;
        RECT 80.600 134.055 80.740 134.210 ;
        RECT 81.980 134.210 87.640 134.350 ;
        RECT 81.980 134.055 82.120 134.210 ;
        RECT 75.465 134.010 75.755 134.055 ;
        RECT 74.530 133.870 75.755 134.010 ;
        RECT 53.370 133.670 53.690 133.730 ;
        RECT 57.985 133.670 58.275 133.715 ;
        RECT 53.370 133.530 58.275 133.670 ;
        RECT 53.370 133.470 53.690 133.530 ;
        RECT 57.985 133.485 58.275 133.530 ;
        RECT 60.730 133.470 61.050 133.730 ;
        RECT 68.090 133.670 68.410 133.730 ;
        RECT 69.485 133.670 69.775 133.715 ;
        RECT 69.930 133.670 70.250 133.730 ;
        RECT 68.090 133.530 70.250 133.670 ;
        RECT 68.090 133.470 68.410 133.530 ;
        RECT 69.485 133.485 69.775 133.530 ;
        RECT 69.930 133.470 70.250 133.530 ;
        RECT 70.390 133.670 70.710 133.730 ;
        RECT 74.160 133.670 74.300 133.825 ;
        RECT 74.530 133.810 74.850 133.870 ;
        RECT 75.465 133.825 75.755 133.870 ;
        RECT 80.525 134.010 80.815 134.055 ;
        RECT 81.905 134.010 82.195 134.055 ;
        RECT 80.525 133.870 82.195 134.010 ;
        RECT 80.525 133.825 80.815 133.870 ;
        RECT 81.905 133.825 82.195 133.870 ;
        RECT 83.730 134.010 84.050 134.070 ;
        RECT 87.500 134.055 87.640 134.210 ;
        RECT 98.400 134.210 101.990 134.350 ;
        RECT 98.400 134.165 98.690 134.210 ;
        RECT 101.660 134.165 101.990 134.210 ;
        RECT 101.670 134.150 101.990 134.165 ;
        RECT 102.580 134.350 102.870 134.395 ;
        RECT 104.440 134.350 104.730 134.395 ;
        RECT 102.580 134.210 104.730 134.350 ;
        RECT 102.580 134.165 102.870 134.210 ;
        RECT 104.440 134.165 104.730 134.210 ;
        RECT 106.270 134.350 106.590 134.410 ;
        RECT 108.125 134.350 108.415 134.395 ;
        RECT 106.270 134.210 108.415 134.350 ;
        RECT 84.665 134.010 84.955 134.055 ;
        RECT 83.730 133.870 84.955 134.010 ;
        RECT 83.730 133.810 84.050 133.870 ;
        RECT 84.665 133.825 84.955 133.870 ;
        RECT 87.425 134.010 87.715 134.055 ;
        RECT 88.790 134.010 89.110 134.070 ;
        RECT 87.425 133.870 89.110 134.010 ;
        RECT 87.425 133.825 87.715 133.870 ;
        RECT 88.790 133.810 89.110 133.870 ;
        RECT 90.630 134.010 90.950 134.070 ;
        RECT 91.105 134.010 91.395 134.055 ;
        RECT 90.630 133.870 91.395 134.010 ;
        RECT 90.630 133.810 90.950 133.870 ;
        RECT 91.105 133.825 91.395 133.870 ;
        RECT 95.230 133.810 95.550 134.070 ;
        RECT 100.260 134.010 100.550 134.055 ;
        RECT 102.580 134.010 102.795 134.165 ;
        RECT 106.270 134.150 106.590 134.210 ;
        RECT 108.125 134.165 108.415 134.210 ;
        RECT 118.690 134.350 119.010 134.410 ;
        RECT 118.690 134.210 122.600 134.350 ;
        RECT 118.690 134.150 119.010 134.210 ;
        RECT 100.260 133.870 102.795 134.010 ;
        RECT 103.140 133.870 105.120 134.010 ;
        RECT 100.260 133.825 100.550 133.870 ;
        RECT 70.390 133.530 74.300 133.670 ;
        RECT 83.270 133.670 83.590 133.730 ;
        RECT 84.205 133.670 84.495 133.715 ;
        RECT 89.725 133.670 90.015 133.715 ;
        RECT 103.140 133.670 103.280 133.870 ;
        RECT 83.270 133.530 103.280 133.670 ;
        RECT 70.390 133.470 70.710 133.530 ;
        RECT 83.270 133.470 83.590 133.530 ;
        RECT 84.205 133.485 84.495 133.530 ;
        RECT 89.725 133.485 90.015 133.530 ;
        RECT 103.510 133.470 103.830 133.730 ;
        RECT 104.980 133.670 105.120 133.870 ;
        RECT 105.350 133.810 105.670 134.070 ;
        RECT 119.150 133.810 119.470 134.070 ;
        RECT 122.460 134.055 122.600 134.210 ;
        RECT 121.005 133.825 121.295 134.055 ;
        RECT 122.385 133.825 122.675 134.055 ;
        RECT 106.730 133.670 107.050 133.730 ;
        RECT 108.585 133.670 108.875 133.715 ;
        RECT 113.170 133.670 113.490 133.730 ;
        RECT 115.485 133.670 115.775 133.715 ;
        RECT 121.080 133.670 121.220 133.825 ;
        RECT 104.980 133.530 115.775 133.670 ;
        RECT 106.730 133.470 107.050 133.530 ;
        RECT 108.585 133.485 108.875 133.530 ;
        RECT 113.170 133.470 113.490 133.530 ;
        RECT 115.485 133.485 115.775 133.530 ;
        RECT 119.470 133.530 121.220 133.670 ;
        RECT 87.885 133.330 88.175 133.375 ;
        RECT 93.850 133.330 94.170 133.390 ;
        RECT 87.885 133.190 94.170 133.330 ;
        RECT 87.885 133.145 88.175 133.190 ;
        RECT 93.850 133.130 94.170 133.190 ;
        RECT 100.260 133.330 100.550 133.375 ;
        RECT 103.040 133.330 103.330 133.375 ;
        RECT 104.900 133.330 105.190 133.375 ;
        RECT 100.260 133.190 105.190 133.330 ;
        RECT 100.260 133.145 100.550 133.190 ;
        RECT 103.040 133.145 103.330 133.190 ;
        RECT 104.900 133.145 105.190 133.190 ;
        RECT 118.705 133.330 118.995 133.375 ;
        RECT 119.470 133.330 119.610 133.530 ;
        RECT 135.590 133.400 136.850 134.480 ;
        RECT 118.705 133.190 119.610 133.330 ;
        RECT 118.705 133.145 118.995 133.190 ;
        RECT 35.430 132.850 53.140 132.990 ;
        RECT 59.825 132.990 60.115 133.035 ;
        RECT 60.285 132.990 60.575 133.035 ;
        RECT 59.825 132.850 60.575 132.990 ;
        RECT 35.430 132.790 35.750 132.850 ;
        RECT 59.825 132.805 60.115 132.850 ;
        RECT 60.285 132.805 60.575 132.850 ;
        RECT 61.190 132.990 61.510 133.050 ;
        RECT 62.585 132.990 62.875 133.035 ;
        RECT 61.190 132.850 62.875 132.990 ;
        RECT 61.190 132.790 61.510 132.850 ;
        RECT 62.585 132.805 62.875 132.850 ;
        RECT 68.105 132.990 68.395 133.035 ;
        RECT 68.550 132.990 68.870 133.050 ;
        RECT 68.105 132.850 68.870 132.990 ;
        RECT 68.105 132.805 68.395 132.850 ;
        RECT 68.550 132.790 68.870 132.850 ;
        RECT 72.690 132.790 73.010 133.050 ;
        RECT 73.610 132.790 73.930 133.050 ;
        RECT 74.530 132.790 74.850 133.050 ;
        RECT 80.970 132.790 81.290 133.050 ;
        RECT 82.350 132.790 82.670 133.050 ;
        RECT 86.965 132.990 87.255 133.035 ;
        RECT 91.090 132.990 91.410 133.050 ;
        RECT 86.965 132.850 91.410 132.990 ;
        RECT 86.965 132.805 87.255 132.850 ;
        RECT 91.090 132.790 91.410 132.850 ;
        RECT 104.430 132.990 104.750 133.050 ;
        RECT 105.825 132.990 106.115 133.035 ;
        RECT 104.430 132.850 106.115 132.990 ;
        RECT 104.430 132.790 104.750 132.850 ;
        RECT 105.825 132.805 106.115 132.850 ;
        RECT 29.840 132.170 127.820 132.650 ;
        RECT 34.525 131.970 34.815 132.015 ;
        RECT 43.250 131.970 43.570 132.030 ;
        RECT 34.525 131.830 43.570 131.970 ;
        RECT 34.525 131.785 34.815 131.830 ;
        RECT 43.250 131.770 43.570 131.830 ;
        RECT 46.470 131.970 46.790 132.030 ;
        RECT 48.095 131.970 48.385 132.015 ;
        RECT 53.370 131.970 53.690 132.030 ;
        RECT 46.470 131.830 53.690 131.970 ;
        RECT 46.470 131.770 46.790 131.830 ;
        RECT 48.095 131.785 48.385 131.830 ;
        RECT 53.370 131.770 53.690 131.830 ;
        RECT 57.510 131.770 57.830 132.030 ;
        RECT 66.495 131.970 66.785 132.015 ;
        RECT 70.850 131.970 71.170 132.030 ;
        RECT 83.270 131.970 83.590 132.030 ;
        RECT 86.490 131.970 86.810 132.030 ;
        RECT 92.255 131.970 92.545 132.015 ;
        RECT 66.495 131.830 71.170 131.970 ;
        RECT 66.495 131.785 66.785 131.830 ;
        RECT 70.850 131.770 71.170 131.830 ;
        RECT 77.380 131.830 83.590 131.970 ;
        RECT 32.685 131.630 32.975 131.675 ;
        RECT 35.430 131.630 35.750 131.690 ;
        RECT 32.685 131.490 35.750 131.630 ;
        RECT 32.685 131.445 32.975 131.490 ;
        RECT 35.430 131.430 35.750 131.490 ;
        RECT 39.590 131.630 39.880 131.675 ;
        RECT 41.450 131.630 41.740 131.675 ;
        RECT 44.230 131.630 44.520 131.675 ;
        RECT 39.590 131.490 44.520 131.630 ;
        RECT 39.590 131.445 39.880 131.490 ;
        RECT 41.450 131.445 41.740 131.490 ;
        RECT 44.230 131.445 44.520 131.490 ;
        RECT 50.625 131.445 50.915 131.675 ;
        RECT 52.450 131.630 52.770 131.690 ;
        RECT 70.360 131.630 70.650 131.675 ;
        RECT 73.140 131.630 73.430 131.675 ;
        RECT 75.000 131.630 75.290 131.675 ;
        RECT 52.450 131.490 55.900 131.630 ;
        RECT 35.890 131.090 36.210 131.350 ;
        RECT 36.365 131.290 36.655 131.335 ;
        RECT 46.470 131.290 46.790 131.350 ;
        RECT 36.365 131.150 46.790 131.290 ;
        RECT 36.365 131.105 36.655 131.150 ;
        RECT 46.470 131.090 46.790 131.150 ;
        RECT 33.145 130.765 33.435 130.995 ;
        RECT 33.605 130.950 33.895 130.995 ;
        RECT 34.050 130.950 34.370 131.010 ;
        RECT 33.605 130.810 34.370 130.950 ;
        RECT 33.605 130.765 33.895 130.810 ;
        RECT 33.220 130.610 33.360 130.765 ;
        RECT 34.050 130.750 34.370 130.810 ;
        RECT 39.125 130.765 39.415 130.995 ;
        RECT 37.270 130.610 37.590 130.670 ;
        RECT 33.220 130.470 37.590 130.610 ;
        RECT 37.270 130.410 37.590 130.470 ;
        RECT 36.810 130.070 37.130 130.330 ;
        RECT 38.650 130.070 38.970 130.330 ;
        RECT 39.200 130.270 39.340 130.765 ;
        RECT 40.950 130.750 41.270 131.010 ;
        RECT 44.230 130.950 44.520 130.995 ;
        RECT 41.985 130.810 44.520 130.950 ;
        RECT 41.985 130.655 42.200 130.810 ;
        RECT 44.230 130.765 44.520 130.810 ;
        RECT 48.785 130.950 49.075 130.995 ;
        RECT 50.700 130.950 50.840 131.445 ;
        RECT 52.450 131.430 52.770 131.490 ;
        RECT 52.910 131.090 53.230 131.350 ;
        RECT 55.760 131.335 55.900 131.490 ;
        RECT 70.360 131.490 75.290 131.630 ;
        RECT 70.360 131.445 70.650 131.490 ;
        RECT 73.140 131.445 73.430 131.490 ;
        RECT 75.000 131.445 75.290 131.490 ;
        RECT 53.385 131.105 53.675 131.335 ;
        RECT 55.685 131.105 55.975 131.335 ;
        RECT 58.905 131.290 59.195 131.335 ;
        RECT 62.585 131.290 62.875 131.335 ;
        RECT 68.090 131.290 68.410 131.350 ;
        RECT 58.905 131.150 68.410 131.290 ;
        RECT 58.905 131.105 59.195 131.150 ;
        RECT 62.585 131.105 62.875 131.150 ;
        RECT 48.785 130.810 50.840 130.950 ;
        RECT 51.070 130.950 51.390 131.010 ;
        RECT 53.460 130.950 53.600 131.105 ;
        RECT 68.090 131.090 68.410 131.150 ;
        RECT 73.625 131.290 73.915 131.335 ;
        RECT 74.530 131.290 74.850 131.350 ;
        RECT 73.625 131.150 74.850 131.290 ;
        RECT 73.625 131.105 73.915 131.150 ;
        RECT 74.530 131.090 74.850 131.150 ;
        RECT 75.450 131.090 75.770 131.350 ;
        RECT 77.380 131.335 77.520 131.830 ;
        RECT 83.270 131.770 83.590 131.830 ;
        RECT 84.280 131.830 92.545 131.970 ;
        RECT 84.280 131.630 84.420 131.830 ;
        RECT 86.490 131.770 86.810 131.830 ;
        RECT 92.255 131.785 92.545 131.830 ;
        RECT 101.670 131.970 101.990 132.030 ;
        RECT 102.605 131.970 102.895 132.015 ;
        RECT 101.670 131.830 102.895 131.970 ;
        RECT 101.670 131.770 101.990 131.830 ;
        RECT 102.605 131.785 102.895 131.830 ;
        RECT 103.510 131.770 103.830 132.030 ;
        RECT 77.840 131.490 84.420 131.630 ;
        RECT 84.620 131.630 84.910 131.675 ;
        RECT 87.400 131.630 87.690 131.675 ;
        RECT 89.260 131.630 89.550 131.675 ;
        RECT 84.620 131.490 89.550 131.630 ;
        RECT 77.840 131.335 77.980 131.490 ;
        RECT 84.620 131.445 84.910 131.490 ;
        RECT 87.400 131.445 87.690 131.490 ;
        RECT 89.260 131.445 89.550 131.490 ;
        RECT 96.120 131.630 96.410 131.675 ;
        RECT 98.900 131.630 99.190 131.675 ;
        RECT 100.760 131.630 101.050 131.675 ;
        RECT 96.120 131.490 101.050 131.630 ;
        RECT 96.120 131.445 96.410 131.490 ;
        RECT 98.900 131.445 99.190 131.490 ;
        RECT 100.760 131.445 101.050 131.490 ;
        RECT 109.965 131.445 110.255 131.675 ;
        RECT 116.405 131.445 116.695 131.675 ;
        RECT 77.305 131.105 77.595 131.335 ;
        RECT 77.765 131.105 78.055 131.335 ;
        RECT 80.755 131.290 81.045 131.335 ;
        RECT 83.730 131.290 84.050 131.350 ;
        RECT 95.230 131.290 95.550 131.350 ;
        RECT 78.300 131.150 84.050 131.290 ;
        RECT 51.070 130.810 53.600 130.950 ;
        RECT 56.605 130.950 56.895 130.995 ;
        RECT 57.050 130.950 57.370 131.010 ;
        RECT 78.300 130.995 78.440 131.150 ;
        RECT 80.755 131.105 81.045 131.150 ;
        RECT 83.730 131.090 84.050 131.150 ;
        RECT 89.800 131.150 95.550 131.290 ;
        RECT 56.605 130.810 57.370 130.950 ;
        RECT 48.785 130.765 49.075 130.810 ;
        RECT 51.070 130.750 51.390 130.810 ;
        RECT 56.605 130.765 56.895 130.810 ;
        RECT 57.050 130.750 57.370 130.810 ;
        RECT 70.360 130.950 70.650 130.995 ;
        RECT 70.360 130.810 72.895 130.950 ;
        RECT 70.360 130.765 70.650 130.810 ;
        RECT 40.050 130.610 40.340 130.655 ;
        RECT 41.910 130.610 42.200 130.655 ;
        RECT 40.050 130.470 42.200 130.610 ;
        RECT 40.050 130.425 40.340 130.470 ;
        RECT 41.910 130.425 42.200 130.470 ;
        RECT 42.790 130.655 43.110 130.670 ;
        RECT 42.790 130.610 43.120 130.655 ;
        RECT 46.090 130.610 46.380 130.655 ;
        RECT 42.790 130.470 46.380 130.610 ;
        RECT 42.790 130.425 43.120 130.470 ;
        RECT 46.090 130.425 46.380 130.470 ;
        RECT 50.150 130.610 50.470 130.670 ;
        RECT 52.465 130.610 52.755 130.655 ;
        RECT 63.505 130.610 63.795 130.655 ;
        RECT 50.150 130.470 52.755 130.610 ;
        RECT 42.790 130.410 43.110 130.425 ;
        RECT 50.150 130.410 50.470 130.470 ;
        RECT 52.465 130.425 52.755 130.470 ;
        RECT 59.900 130.470 63.795 130.610 ;
        RECT 59.900 130.330 60.040 130.470 ;
        RECT 63.505 130.425 63.795 130.470 ;
        RECT 63.965 130.610 64.255 130.655 ;
        RECT 64.870 130.610 65.190 130.670 ;
        RECT 68.550 130.655 68.870 130.670 ;
        RECT 72.680 130.655 72.895 130.810 ;
        RECT 78.225 130.765 78.515 130.995 ;
        RECT 84.620 130.950 84.910 130.995 ;
        RECT 87.885 130.950 88.175 130.995 ;
        RECT 88.330 130.950 88.650 131.010 ;
        RECT 84.620 130.810 87.155 130.950 ;
        RECT 84.620 130.765 84.910 130.810 ;
        RECT 63.965 130.470 65.190 130.610 ;
        RECT 63.965 130.425 64.255 130.470 ;
        RECT 64.870 130.410 65.190 130.470 ;
        RECT 68.500 130.610 68.870 130.655 ;
        RECT 71.760 130.610 72.050 130.655 ;
        RECT 68.500 130.470 72.050 130.610 ;
        RECT 68.500 130.425 68.870 130.470 ;
        RECT 71.760 130.425 72.050 130.470 ;
        RECT 72.680 130.610 72.970 130.655 ;
        RECT 74.540 130.610 74.830 130.655 ;
        RECT 72.680 130.470 74.830 130.610 ;
        RECT 72.680 130.425 72.970 130.470 ;
        RECT 74.540 130.425 74.830 130.470 ;
        RECT 80.970 130.610 81.290 130.670 ;
        RECT 86.940 130.655 87.155 130.810 ;
        RECT 87.885 130.810 88.650 130.950 ;
        RECT 87.885 130.765 88.175 130.810 ;
        RECT 88.330 130.750 88.650 130.810 ;
        RECT 89.250 130.950 89.570 131.010 ;
        RECT 89.800 130.995 89.940 131.150 ;
        RECT 95.230 131.090 95.550 131.150 ;
        RECT 98.450 131.290 98.770 131.350 ;
        RECT 101.225 131.290 101.515 131.335 ;
        RECT 105.350 131.290 105.670 131.350 ;
        RECT 98.450 131.150 100.060 131.290 ;
        RECT 98.450 131.090 98.770 131.150 ;
        RECT 89.725 130.950 90.015 130.995 ;
        RECT 89.250 130.810 90.015 130.950 ;
        RECT 89.250 130.750 89.570 130.810 ;
        RECT 89.725 130.765 90.015 130.810 ;
        RECT 91.090 130.750 91.410 131.010 ;
        RECT 96.120 130.950 96.410 130.995 ;
        RECT 96.120 130.810 98.655 130.950 ;
        RECT 96.120 130.765 96.410 130.810 ;
        RECT 82.760 130.610 83.050 130.655 ;
        RECT 86.020 130.610 86.310 130.655 ;
        RECT 80.970 130.470 86.310 130.610 ;
        RECT 68.550 130.410 68.870 130.425 ;
        RECT 80.970 130.410 81.290 130.470 ;
        RECT 82.760 130.425 83.050 130.470 ;
        RECT 86.020 130.425 86.310 130.470 ;
        RECT 86.940 130.610 87.230 130.655 ;
        RECT 88.800 130.610 89.090 130.655 ;
        RECT 86.940 130.470 89.090 130.610 ;
        RECT 86.940 130.425 87.230 130.470 ;
        RECT 88.800 130.425 89.090 130.470 ;
        RECT 94.260 130.610 94.550 130.655 ;
        RECT 95.690 130.610 96.010 130.670 ;
        RECT 98.440 130.655 98.655 130.810 ;
        RECT 99.370 130.750 99.690 131.010 ;
        RECT 99.920 130.950 100.060 131.150 ;
        RECT 101.225 131.150 105.670 131.290 ;
        RECT 101.225 131.105 101.515 131.150 ;
        RECT 105.350 131.090 105.670 131.150 ;
        RECT 106.730 131.090 107.050 131.350 ;
        RECT 102.145 130.950 102.435 130.995 ;
        RECT 99.920 130.810 102.435 130.950 ;
        RECT 102.145 130.765 102.435 130.810 ;
        RECT 104.430 130.750 104.750 131.010 ;
        RECT 108.125 130.950 108.415 130.995 ;
        RECT 109.030 130.950 109.350 131.010 ;
        RECT 108.125 130.810 109.350 130.950 ;
        RECT 110.040 130.950 110.180 131.445 ;
        RECT 113.170 131.090 113.490 131.350 ;
        RECT 116.480 131.290 116.620 131.445 ;
        RECT 116.480 131.150 118.920 131.290 ;
        RECT 118.780 130.995 118.920 131.150 ;
        RECT 110.425 130.950 110.715 130.995 ;
        RECT 110.040 130.810 110.715 130.950 ;
        RECT 108.125 130.765 108.415 130.810 ;
        RECT 109.030 130.750 109.350 130.810 ;
        RECT 110.425 130.765 110.715 130.810 ;
        RECT 117.325 130.765 117.615 130.995 ;
        RECT 118.705 130.765 118.995 130.995 ;
        RECT 97.520 130.610 97.810 130.655 ;
        RECT 94.260 130.470 97.810 130.610 ;
        RECT 94.260 130.425 94.550 130.470 ;
        RECT 95.690 130.410 96.010 130.470 ;
        RECT 97.520 130.425 97.810 130.470 ;
        RECT 98.440 130.610 98.730 130.655 ;
        RECT 100.300 130.610 100.590 130.655 ;
        RECT 98.440 130.470 100.590 130.610 ;
        RECT 109.120 130.610 109.260 130.750 ;
        RECT 114.105 130.610 114.395 130.655 ;
        RECT 109.120 130.470 114.395 130.610 ;
        RECT 117.400 130.610 117.540 130.765 ;
        RECT 119.150 130.610 119.470 130.670 ;
        RECT 117.400 130.470 119.470 130.610 ;
        RECT 98.440 130.425 98.730 130.470 ;
        RECT 100.300 130.425 100.590 130.470 ;
        RECT 114.105 130.425 114.395 130.470 ;
        RECT 119.150 130.410 119.470 130.470 ;
        RECT 44.170 130.270 44.490 130.330 ;
        RECT 39.200 130.130 44.490 130.270 ;
        RECT 44.170 130.070 44.490 130.130 ;
        RECT 49.705 130.270 49.995 130.315 ;
        RECT 51.070 130.270 51.390 130.330 ;
        RECT 49.705 130.130 51.390 130.270 ;
        RECT 49.705 130.085 49.995 130.130 ;
        RECT 51.070 130.070 51.390 130.130 ;
        RECT 54.290 130.270 54.610 130.330 ;
        RECT 59.365 130.270 59.655 130.315 ;
        RECT 54.290 130.130 59.655 130.270 ;
        RECT 54.290 130.070 54.610 130.130 ;
        RECT 59.365 130.085 59.655 130.130 ;
        RECT 59.810 130.070 60.130 130.330 ;
        RECT 61.665 130.270 61.955 130.315 ;
        RECT 64.410 130.270 64.730 130.330 ;
        RECT 61.665 130.130 64.730 130.270 ;
        RECT 61.665 130.085 61.955 130.130 ;
        RECT 64.410 130.070 64.730 130.130 ;
        RECT 65.805 130.270 66.095 130.315 ;
        RECT 66.250 130.270 66.570 130.330 ;
        RECT 65.805 130.130 66.570 130.270 ;
        RECT 65.805 130.085 66.095 130.130 ;
        RECT 66.250 130.070 66.570 130.130 ;
        RECT 80.050 130.070 80.370 130.330 ;
        RECT 90.170 130.070 90.490 130.330 ;
        RECT 90.630 130.270 90.950 130.330 ;
        RECT 107.665 130.270 107.955 130.315 ;
        RECT 90.630 130.130 107.955 130.270 ;
        RECT 90.630 130.070 90.950 130.130 ;
        RECT 107.665 130.085 107.955 130.130 ;
        RECT 111.345 130.270 111.635 130.315 ;
        RECT 112.250 130.270 112.570 130.330 ;
        RECT 111.345 130.130 112.570 130.270 ;
        RECT 111.345 130.085 111.635 130.130 ;
        RECT 112.250 130.070 112.570 130.130 ;
        RECT 114.550 130.070 114.870 130.330 ;
        RECT 117.770 130.070 118.090 130.330 ;
        RECT 119.625 130.270 119.915 130.315 ;
        RECT 122.370 130.270 122.690 130.330 ;
        RECT 119.625 130.130 122.690 130.270 ;
        RECT 119.625 130.085 119.915 130.130 ;
        RECT 122.370 130.070 122.690 130.130 ;
        RECT 29.840 129.450 127.820 129.930 ;
        RECT 39.125 129.250 39.415 129.295 ;
        RECT 39.570 129.250 39.890 129.310 ;
        RECT 39.125 129.110 39.890 129.250 ;
        RECT 39.125 129.065 39.415 129.110 ;
        RECT 39.570 129.050 39.890 129.110 ;
        RECT 40.950 129.250 41.270 129.310 ;
        RECT 41.885 129.250 42.175 129.295 ;
        RECT 40.950 129.110 42.175 129.250 ;
        RECT 40.950 129.050 41.270 129.110 ;
        RECT 41.885 129.065 42.175 129.110 ;
        RECT 53.615 129.250 53.905 129.295 ;
        RECT 54.290 129.250 54.610 129.310 ;
        RECT 53.615 129.110 54.610 129.250 ;
        RECT 53.615 129.065 53.905 129.110 ;
        RECT 54.290 129.050 54.610 129.110 ;
        RECT 56.130 129.250 56.450 129.310 ;
        RECT 64.870 129.250 65.190 129.310 ;
        RECT 68.335 129.250 68.625 129.295 ;
        RECT 56.130 129.110 62.800 129.250 ;
        RECT 56.130 129.050 56.450 129.110 ;
        RECT 35.905 128.910 36.195 128.955 ;
        RECT 41.410 128.910 41.730 128.970 ;
        RECT 35.905 128.770 41.730 128.910 ;
        RECT 35.905 128.725 36.195 128.770 ;
        RECT 41.410 128.710 41.730 128.770 ;
        RECT 42.805 128.910 43.095 128.955 ;
        RECT 45.960 128.910 46.250 128.955 ;
        RECT 49.220 128.910 49.510 128.955 ;
        RECT 42.805 128.770 49.510 128.910 ;
        RECT 42.805 128.725 43.095 128.770 ;
        RECT 45.960 128.725 46.250 128.770 ;
        RECT 49.220 128.725 49.510 128.770 ;
        RECT 50.140 128.910 50.430 128.955 ;
        RECT 52.000 128.910 52.290 128.955 ;
        RECT 50.140 128.770 52.290 128.910 ;
        RECT 50.140 128.725 50.430 128.770 ;
        RECT 52.000 128.725 52.290 128.770 ;
        RECT 55.620 128.910 55.910 128.955 ;
        RECT 56.590 128.910 56.910 128.970 ;
        RECT 58.880 128.910 59.170 128.955 ;
        RECT 55.620 128.770 59.170 128.910 ;
        RECT 55.620 128.725 55.910 128.770 ;
        RECT 35.445 128.385 35.735 128.615 ;
        RECT 38.205 128.570 38.495 128.615 ;
        RECT 38.650 128.570 38.970 128.630 ;
        RECT 38.205 128.430 38.970 128.570 ;
        RECT 38.205 128.385 38.495 128.430 ;
        RECT 35.520 128.230 35.660 128.385 ;
        RECT 38.650 128.370 38.970 128.430 ;
        RECT 39.585 128.385 39.875 128.615 ;
        RECT 37.270 128.230 37.590 128.290 ;
        RECT 39.660 128.230 39.800 128.385 ;
        RECT 40.950 128.370 41.270 128.630 ;
        RECT 42.345 128.570 42.635 128.615 ;
        RECT 47.820 128.570 48.110 128.615 ;
        RECT 50.140 128.570 50.355 128.725 ;
        RECT 56.590 128.710 56.910 128.770 ;
        RECT 58.880 128.725 59.170 128.770 ;
        RECT 59.800 128.910 60.090 128.955 ;
        RECT 61.660 128.910 61.950 128.955 ;
        RECT 59.800 128.770 61.950 128.910 ;
        RECT 59.800 128.725 60.090 128.770 ;
        RECT 61.660 128.725 61.950 128.770 ;
        RECT 42.345 128.430 43.480 128.570 ;
        RECT 42.345 128.385 42.635 128.430 ;
        RECT 35.520 128.090 39.800 128.230 ;
        RECT 37.270 128.030 37.590 128.090 ;
        RECT 39.660 127.890 39.800 128.090 ;
        RECT 40.045 128.230 40.335 128.275 ;
        RECT 42.790 128.230 43.110 128.290 ;
        RECT 40.045 128.090 43.110 128.230 ;
        RECT 40.045 128.045 40.335 128.090 ;
        RECT 42.790 128.030 43.110 128.090 ;
        RECT 43.340 128.230 43.480 128.430 ;
        RECT 47.820 128.430 50.355 128.570 ;
        RECT 47.820 128.385 48.110 128.430 ;
        RECT 51.070 128.370 51.390 128.630 ;
        RECT 57.480 128.570 57.770 128.615 ;
        RECT 59.800 128.570 60.015 128.725 ;
        RECT 62.660 128.615 62.800 129.110 ;
        RECT 64.870 129.110 68.625 129.250 ;
        RECT 64.870 129.050 65.190 129.110 ;
        RECT 68.335 129.065 68.625 129.110 ;
        RECT 79.375 129.250 79.665 129.295 ;
        RECT 81.890 129.250 82.210 129.310 ;
        RECT 79.375 129.110 82.210 129.250 ;
        RECT 79.375 129.065 79.665 129.110 ;
        RECT 81.890 129.050 82.210 129.110 ;
        RECT 89.495 129.250 89.785 129.295 ;
        RECT 90.630 129.250 90.950 129.310 ;
        RECT 89.495 129.110 90.950 129.250 ;
        RECT 89.495 129.065 89.785 129.110 ;
        RECT 90.630 129.050 90.950 129.110 ;
        RECT 99.370 129.050 99.690 129.310 ;
        RECT 105.135 129.250 105.425 129.295 ;
        RECT 109.030 129.250 109.350 129.310 ;
        RECT 105.135 129.110 109.350 129.250 ;
        RECT 105.135 129.065 105.425 129.110 ;
        RECT 109.030 129.050 109.350 129.110 ;
        RECT 114.550 129.250 114.870 129.310 ;
        RECT 115.255 129.250 115.545 129.295 ;
        RECT 114.550 129.110 115.545 129.250 ;
        RECT 114.550 129.050 114.870 129.110 ;
        RECT 115.255 129.065 115.545 129.110 ;
        RECT 73.610 128.955 73.930 128.970 ;
        RECT 70.340 128.910 70.630 128.955 ;
        RECT 73.600 128.910 73.930 128.955 ;
        RECT 70.340 128.770 73.930 128.910 ;
        RECT 70.340 128.725 70.630 128.770 ;
        RECT 73.600 128.725 73.930 128.770 ;
        RECT 73.610 128.710 73.930 128.725 ;
        RECT 74.520 128.910 74.810 128.955 ;
        RECT 76.380 128.910 76.670 128.955 ;
        RECT 74.520 128.770 76.670 128.910 ;
        RECT 74.520 128.725 74.810 128.770 ;
        RECT 76.380 128.725 76.670 128.770 ;
        RECT 81.380 128.910 81.670 128.955 ;
        RECT 82.350 128.910 82.670 128.970 ;
        RECT 84.640 128.910 84.930 128.955 ;
        RECT 81.380 128.770 84.930 128.910 ;
        RECT 81.380 128.725 81.670 128.770 ;
        RECT 57.480 128.430 60.015 128.570 ;
        RECT 57.480 128.385 57.770 128.430 ;
        RECT 62.585 128.385 62.875 128.615 ;
        RECT 64.410 128.370 64.730 128.630 ;
        RECT 65.790 128.370 66.110 128.630 ;
        RECT 66.250 128.370 66.570 128.630 ;
        RECT 72.200 128.570 72.490 128.615 ;
        RECT 74.520 128.570 74.735 128.725 ;
        RECT 82.350 128.710 82.670 128.770 ;
        RECT 84.640 128.725 84.930 128.770 ;
        RECT 85.560 128.910 85.850 128.955 ;
        RECT 87.420 128.910 87.710 128.955 ;
        RECT 85.560 128.770 87.710 128.910 ;
        RECT 85.560 128.725 85.850 128.770 ;
        RECT 87.420 128.725 87.710 128.770 ;
        RECT 91.500 128.910 91.790 128.955 ;
        RECT 93.850 128.910 94.170 128.970 ;
        RECT 94.760 128.910 95.050 128.955 ;
        RECT 91.500 128.770 95.050 128.910 ;
        RECT 91.500 128.725 91.790 128.770 ;
        RECT 72.200 128.430 74.735 128.570 ;
        RECT 75.910 128.570 76.230 128.630 ;
        RECT 77.305 128.570 77.595 128.615 ;
        RECT 75.910 128.430 77.595 128.570 ;
        RECT 72.200 128.385 72.490 128.430 ;
        RECT 75.910 128.370 76.230 128.430 ;
        RECT 77.305 128.385 77.595 128.430 ;
        RECT 83.240 128.570 83.530 128.615 ;
        RECT 85.560 128.570 85.775 128.725 ;
        RECT 93.850 128.710 94.170 128.770 ;
        RECT 94.760 128.725 95.050 128.770 ;
        RECT 95.680 128.910 95.970 128.955 ;
        RECT 97.540 128.910 97.830 128.955 ;
        RECT 95.680 128.770 97.830 128.910 ;
        RECT 95.680 128.725 95.970 128.770 ;
        RECT 97.540 128.725 97.830 128.770 ;
        RECT 107.140 128.910 107.430 128.955 ;
        RECT 108.570 128.910 108.890 128.970 ;
        RECT 110.400 128.910 110.690 128.955 ;
        RECT 107.140 128.770 110.690 128.910 ;
        RECT 107.140 128.725 107.430 128.770 ;
        RECT 83.240 128.430 85.775 128.570 ;
        RECT 86.505 128.570 86.795 128.615 ;
        RECT 90.170 128.570 90.490 128.630 ;
        RECT 86.505 128.430 90.490 128.570 ;
        RECT 83.240 128.385 83.530 128.430 ;
        RECT 86.505 128.385 86.795 128.430 ;
        RECT 90.170 128.370 90.490 128.430 ;
        RECT 93.360 128.570 93.650 128.615 ;
        RECT 95.680 128.570 95.895 128.725 ;
        RECT 108.570 128.710 108.890 128.770 ;
        RECT 110.400 128.725 110.690 128.770 ;
        RECT 111.320 128.910 111.610 128.955 ;
        RECT 113.180 128.910 113.470 128.955 ;
        RECT 111.320 128.770 113.470 128.910 ;
        RECT 111.320 128.725 111.610 128.770 ;
        RECT 113.180 128.725 113.470 128.770 ;
        RECT 117.260 128.910 117.550 128.955 ;
        RECT 117.770 128.910 118.090 128.970 ;
        RECT 120.520 128.910 120.810 128.955 ;
        RECT 117.260 128.770 120.810 128.910 ;
        RECT 117.260 128.725 117.550 128.770 ;
        RECT 93.360 128.430 95.895 128.570 ;
        RECT 93.360 128.385 93.650 128.430 ;
        RECT 96.610 128.370 96.930 128.630 ;
        RECT 100.290 128.370 100.610 128.630 ;
        RECT 109.000 128.570 109.290 128.615 ;
        RECT 111.320 128.570 111.535 128.725 ;
        RECT 117.770 128.710 118.090 128.770 ;
        RECT 120.520 128.725 120.810 128.770 ;
        RECT 121.440 128.910 121.730 128.955 ;
        RECT 123.300 128.910 123.590 128.955 ;
        RECT 121.440 128.770 123.590 128.910 ;
        RECT 121.440 128.725 121.730 128.770 ;
        RECT 123.300 128.725 123.590 128.770 ;
        RECT 109.000 128.430 111.535 128.570 ;
        RECT 109.000 128.385 109.290 128.430 ;
        RECT 112.250 128.370 112.570 128.630 ;
        RECT 119.120 128.570 119.410 128.615 ;
        RECT 121.440 128.570 121.655 128.725 ;
        RECT 119.120 128.430 121.655 128.570 ;
        RECT 119.120 128.385 119.410 128.430 ;
        RECT 122.370 128.370 122.690 128.630 ;
        RECT 124.225 128.570 124.515 128.615 ;
        RECT 125.130 128.570 125.450 128.630 ;
        RECT 124.225 128.430 125.450 128.570 ;
        RECT 124.225 128.385 124.515 128.430 ;
        RECT 45.550 128.230 45.870 128.290 ;
        RECT 43.340 128.090 45.870 128.230 ;
        RECT 43.340 127.890 43.480 128.090 ;
        RECT 45.550 128.030 45.870 128.090 ;
        RECT 49.690 128.230 50.010 128.290 ;
        RECT 52.925 128.230 53.215 128.275 ;
        RECT 57.050 128.230 57.370 128.290 ;
        RECT 49.690 128.090 57.370 128.230 ;
        RECT 49.690 128.030 50.010 128.090 ;
        RECT 52.925 128.045 53.215 128.090 ;
        RECT 57.050 128.030 57.370 128.090 ;
        RECT 60.745 128.230 61.035 128.275 ;
        RECT 74.530 128.230 74.850 128.290 ;
        RECT 75.465 128.230 75.755 128.275 ;
        RECT 60.745 128.090 63.720 128.230 ;
        RECT 60.745 128.045 61.035 128.090 ;
        RECT 63.580 127.935 63.720 128.090 ;
        RECT 74.530 128.090 75.755 128.230 ;
        RECT 74.530 128.030 74.850 128.090 ;
        RECT 75.465 128.045 75.755 128.090 ;
        RECT 88.345 128.230 88.635 128.275 ;
        RECT 89.250 128.230 89.570 128.290 ;
        RECT 88.345 128.090 89.570 128.230 ;
        RECT 88.345 128.045 88.635 128.090 ;
        RECT 89.250 128.030 89.570 128.090 ;
        RECT 95.230 128.230 95.550 128.290 ;
        RECT 98.465 128.230 98.755 128.275 ;
        RECT 95.230 128.090 98.755 128.230 ;
        RECT 95.230 128.030 95.550 128.090 ;
        RECT 98.465 128.045 98.755 128.090 ;
        RECT 114.105 128.230 114.395 128.275 ;
        RECT 124.300 128.230 124.440 128.385 ;
        RECT 125.130 128.370 125.450 128.430 ;
        RECT 114.105 128.090 124.440 128.230 ;
        RECT 114.105 128.045 114.395 128.090 ;
        RECT 39.660 127.750 43.480 127.890 ;
        RECT 47.820 127.890 48.110 127.935 ;
        RECT 50.600 127.890 50.890 127.935 ;
        RECT 52.460 127.890 52.750 127.935 ;
        RECT 47.820 127.750 52.750 127.890 ;
        RECT 47.820 127.705 48.110 127.750 ;
        RECT 50.600 127.705 50.890 127.750 ;
        RECT 52.460 127.705 52.750 127.750 ;
        RECT 57.480 127.890 57.770 127.935 ;
        RECT 60.260 127.890 60.550 127.935 ;
        RECT 62.120 127.890 62.410 127.935 ;
        RECT 57.480 127.750 62.410 127.890 ;
        RECT 57.480 127.705 57.770 127.750 ;
        RECT 60.260 127.705 60.550 127.750 ;
        RECT 62.120 127.705 62.410 127.750 ;
        RECT 63.505 127.705 63.795 127.935 ;
        RECT 72.200 127.890 72.490 127.935 ;
        RECT 74.980 127.890 75.270 127.935 ;
        RECT 76.840 127.890 77.130 127.935 ;
        RECT 72.200 127.750 77.130 127.890 ;
        RECT 72.200 127.705 72.490 127.750 ;
        RECT 74.980 127.705 75.270 127.750 ;
        RECT 76.840 127.705 77.130 127.750 ;
        RECT 83.240 127.890 83.530 127.935 ;
        RECT 86.020 127.890 86.310 127.935 ;
        RECT 87.880 127.890 88.170 127.935 ;
        RECT 83.240 127.750 88.170 127.890 ;
        RECT 83.240 127.705 83.530 127.750 ;
        RECT 86.020 127.705 86.310 127.750 ;
        RECT 87.880 127.705 88.170 127.750 ;
        RECT 93.360 127.890 93.650 127.935 ;
        RECT 96.140 127.890 96.430 127.935 ;
        RECT 98.000 127.890 98.290 127.935 ;
        RECT 93.360 127.750 98.290 127.890 ;
        RECT 93.360 127.705 93.650 127.750 ;
        RECT 96.140 127.705 96.430 127.750 ;
        RECT 98.000 127.705 98.290 127.750 ;
        RECT 109.000 127.890 109.290 127.935 ;
        RECT 111.780 127.890 112.070 127.935 ;
        RECT 113.640 127.890 113.930 127.935 ;
        RECT 109.000 127.750 113.930 127.890 ;
        RECT 109.000 127.705 109.290 127.750 ;
        RECT 111.780 127.705 112.070 127.750 ;
        RECT 113.640 127.705 113.930 127.750 ;
        RECT 119.120 127.890 119.410 127.935 ;
        RECT 121.900 127.890 122.190 127.935 ;
        RECT 123.760 127.890 124.050 127.935 ;
        RECT 119.120 127.750 124.050 127.890 ;
        RECT 119.120 127.705 119.410 127.750 ;
        RECT 121.900 127.705 122.190 127.750 ;
        RECT 123.760 127.705 124.050 127.750 ;
        RECT 43.955 127.550 44.245 127.595 ;
        RECT 50.150 127.550 50.470 127.610 ;
        RECT 43.955 127.410 50.470 127.550 ;
        RECT 43.955 127.365 44.245 127.410 ;
        RECT 50.150 127.350 50.470 127.410 ;
        RECT 63.950 127.550 64.270 127.610 ;
        RECT 65.345 127.550 65.635 127.595 ;
        RECT 63.950 127.410 65.635 127.550 ;
        RECT 63.950 127.350 64.270 127.410 ;
        RECT 65.345 127.365 65.635 127.410 ;
        RECT 66.250 127.550 66.570 127.610 ;
        RECT 67.185 127.550 67.475 127.595 ;
        RECT 66.250 127.410 67.475 127.550 ;
        RECT 66.250 127.350 66.570 127.410 ;
        RECT 67.185 127.365 67.475 127.410 ;
        RECT 29.840 126.730 127.820 127.210 ;
        RECT 36.810 126.530 37.130 126.590 ;
        RECT 55.670 126.530 55.990 126.590 ;
        RECT 36.810 126.390 55.990 126.530 ;
        RECT 36.810 126.330 37.130 126.390 ;
        RECT 55.670 126.330 55.990 126.390 ;
        RECT 59.135 126.530 59.425 126.575 ;
        RECT 59.810 126.530 60.130 126.590 ;
        RECT 59.135 126.390 60.130 126.530 ;
        RECT 59.135 126.345 59.425 126.390 ;
        RECT 59.810 126.330 60.130 126.390 ;
        RECT 74.530 126.330 74.850 126.590 ;
        RECT 88.330 126.330 88.650 126.590 ;
        RECT 38.305 126.190 38.595 126.235 ;
        RECT 41.425 126.190 41.715 126.235 ;
        RECT 43.315 126.190 43.605 126.235 ;
        RECT 50.150 126.190 50.470 126.250 ;
        RECT 63.000 126.190 63.290 126.235 ;
        RECT 65.780 126.190 66.070 126.235 ;
        RECT 67.640 126.190 67.930 126.235 ;
        RECT 38.305 126.050 43.605 126.190 ;
        RECT 38.305 126.005 38.595 126.050 ;
        RECT 41.425 126.005 41.715 126.050 ;
        RECT 43.315 126.005 43.605 126.050 ;
        RECT 47.480 126.050 54.520 126.190 ;
        RECT 42.790 125.650 43.110 125.910 ;
        RECT 47.480 125.895 47.620 126.050 ;
        RECT 50.150 125.990 50.470 126.050 ;
        RECT 47.405 125.665 47.695 125.895 ;
        RECT 48.325 125.850 48.615 125.895 ;
        RECT 50.610 125.850 50.930 125.910 ;
        RECT 54.380 125.895 54.520 126.050 ;
        RECT 63.000 126.050 67.930 126.190 ;
        RECT 63.000 126.005 63.290 126.050 ;
        RECT 65.780 126.005 66.070 126.050 ;
        RECT 67.640 126.005 67.930 126.050 ;
        RECT 122.845 126.005 123.135 126.235 ;
        RECT 48.325 125.710 50.930 125.850 ;
        RECT 48.325 125.665 48.615 125.710 ;
        RECT 50.610 125.650 50.930 125.710 ;
        RECT 54.305 125.665 54.595 125.895 ;
        RECT 55.670 125.850 55.990 125.910 ;
        RECT 56.605 125.850 56.895 125.895 ;
        RECT 55.670 125.710 56.895 125.850 ;
        RECT 55.670 125.650 55.990 125.710 ;
        RECT 56.605 125.665 56.895 125.710 ;
        RECT 57.050 125.850 57.370 125.910 ;
        RECT 57.050 125.710 66.020 125.850 ;
        RECT 57.050 125.650 57.370 125.710 ;
        RECT 34.065 125.170 34.355 125.215 ;
        RECT 35.890 125.170 36.210 125.230 ;
        RECT 37.225 125.215 37.515 125.530 ;
        RECT 38.305 125.510 38.595 125.555 ;
        RECT 41.885 125.510 42.175 125.555 ;
        RECT 43.720 125.510 44.010 125.555 ;
        RECT 38.305 125.370 44.010 125.510 ;
        RECT 38.305 125.325 38.595 125.370 ;
        RECT 41.885 125.325 42.175 125.370 ;
        RECT 43.720 125.325 44.010 125.370 ;
        RECT 44.170 125.310 44.490 125.570 ;
        RECT 46.470 125.510 46.790 125.570 ;
        RECT 46.945 125.510 47.235 125.555 ;
        RECT 46.470 125.370 47.235 125.510 ;
        RECT 46.470 125.310 46.790 125.370 ;
        RECT 46.945 125.325 47.235 125.370 ;
        RECT 53.370 125.310 53.690 125.570 ;
        RECT 55.225 125.510 55.515 125.555 ;
        RECT 57.510 125.510 57.830 125.570 ;
        RECT 55.225 125.370 57.830 125.510 ;
        RECT 55.225 125.325 55.515 125.370 ;
        RECT 57.510 125.310 57.830 125.370 ;
        RECT 58.430 125.310 58.750 125.570 ;
        RECT 63.000 125.510 63.290 125.555 ;
        RECT 65.880 125.510 66.020 125.710 ;
        RECT 66.250 125.650 66.570 125.910 ;
        RECT 75.450 125.850 75.770 125.910 ;
        RECT 71.170 125.710 75.770 125.850 ;
        RECT 68.105 125.510 68.395 125.555 ;
        RECT 68.550 125.510 68.870 125.570 ;
        RECT 71.170 125.510 71.310 125.710 ;
        RECT 75.450 125.650 75.770 125.710 ;
        RECT 88.790 125.850 89.110 125.910 ;
        RECT 98.450 125.850 98.770 125.910 ;
        RECT 88.790 125.710 98.770 125.850 ;
        RECT 88.790 125.650 89.110 125.710 ;
        RECT 63.000 125.370 65.535 125.510 ;
        RECT 65.880 125.370 71.310 125.510 ;
        RECT 72.690 125.510 73.010 125.570 ;
        RECT 73.625 125.510 73.915 125.555 ;
        RECT 72.690 125.370 73.915 125.510 ;
        RECT 63.000 125.325 63.290 125.370 ;
        RECT 34.065 125.030 36.210 125.170 ;
        RECT 34.065 124.985 34.355 125.030 ;
        RECT 35.890 124.970 36.210 125.030 ;
        RECT 36.925 125.170 37.515 125.215 ;
        RECT 37.730 125.170 38.050 125.230 ;
        RECT 40.165 125.170 40.815 125.215 ;
        RECT 36.925 125.030 40.815 125.170 ;
        RECT 44.260 125.170 44.400 125.310 ;
        RECT 49.690 125.170 50.010 125.230 ;
        RECT 44.260 125.030 50.010 125.170 ;
        RECT 36.925 124.985 37.215 125.030 ;
        RECT 37.730 124.970 38.050 125.030 ;
        RECT 40.165 124.985 40.815 125.030 ;
        RECT 49.690 124.970 50.010 125.030 ;
        RECT 52.005 124.985 52.295 125.215 ;
        RECT 61.140 125.170 61.430 125.215 ;
        RECT 63.490 125.170 63.810 125.230 ;
        RECT 65.320 125.215 65.535 125.370 ;
        RECT 68.105 125.325 68.395 125.370 ;
        RECT 68.550 125.310 68.870 125.370 ;
        RECT 72.690 125.310 73.010 125.370 ;
        RECT 73.625 125.325 73.915 125.370 ;
        RECT 80.050 125.510 80.370 125.570 ;
        RECT 87.425 125.510 87.715 125.555 ;
        RECT 80.050 125.370 87.715 125.510 ;
        RECT 80.050 125.310 80.370 125.370 ;
        RECT 87.425 125.325 87.715 125.370 ;
        RECT 95.690 125.510 96.010 125.570 ;
        RECT 96.700 125.555 96.840 125.710 ;
        RECT 98.450 125.650 98.770 125.710 ;
        RECT 96.165 125.510 96.455 125.555 ;
        RECT 95.690 125.370 96.455 125.510 ;
        RECT 95.690 125.310 96.010 125.370 ;
        RECT 96.165 125.325 96.455 125.370 ;
        RECT 96.625 125.325 96.915 125.555 ;
        RECT 108.570 125.510 108.890 125.570 ;
        RECT 109.045 125.510 109.335 125.555 ;
        RECT 108.570 125.370 109.335 125.510 ;
        RECT 108.570 125.310 108.890 125.370 ;
        RECT 109.045 125.325 109.335 125.370 ;
        RECT 109.505 125.510 109.795 125.555 ;
        RECT 109.950 125.510 110.270 125.570 ;
        RECT 109.505 125.370 110.270 125.510 ;
        RECT 109.505 125.325 109.795 125.370 ;
        RECT 109.950 125.310 110.270 125.370 ;
        RECT 119.610 125.510 119.930 125.570 ;
        RECT 120.085 125.510 120.375 125.555 ;
        RECT 119.610 125.370 120.375 125.510 ;
        RECT 119.610 125.310 119.930 125.370 ;
        RECT 120.085 125.325 120.375 125.370 ;
        RECT 120.530 125.510 120.850 125.570 ;
        RECT 121.465 125.510 121.755 125.555 ;
        RECT 120.530 125.370 121.755 125.510 ;
        RECT 120.530 125.310 120.850 125.370 ;
        RECT 121.465 125.325 121.755 125.370 ;
        RECT 64.400 125.170 64.690 125.215 ;
        RECT 61.140 125.030 64.690 125.170 ;
        RECT 61.140 124.985 61.430 125.030 ;
        RECT 40.950 124.830 41.270 124.890 ;
        RECT 45.105 124.830 45.395 124.875 ;
        RECT 40.950 124.690 45.395 124.830 ;
        RECT 40.950 124.630 41.270 124.690 ;
        RECT 45.105 124.645 45.395 124.690 ;
        RECT 45.550 124.830 45.870 124.890 ;
        RECT 52.080 124.830 52.220 124.985 ;
        RECT 63.490 124.970 63.810 125.030 ;
        RECT 64.400 124.985 64.690 125.030 ;
        RECT 65.320 125.170 65.610 125.215 ;
        RECT 67.180 125.170 67.470 125.215 ;
        RECT 65.320 125.030 67.470 125.170 ;
        RECT 65.320 124.985 65.610 125.030 ;
        RECT 67.180 124.985 67.470 125.030 ;
        RECT 117.310 125.170 117.630 125.230 ;
        RECT 122.920 125.170 123.060 126.005 ;
        RECT 123.290 125.510 123.610 125.570 ;
        RECT 123.765 125.510 124.055 125.555 ;
        RECT 123.290 125.370 124.055 125.510 ;
        RECT 123.290 125.310 123.610 125.370 ;
        RECT 123.765 125.325 124.055 125.370 ;
        RECT 117.310 125.030 123.060 125.170 ;
        RECT 117.310 124.970 117.630 125.030 ;
        RECT 45.550 124.690 52.220 124.830 ;
        RECT 56.145 124.830 56.435 124.875 ;
        RECT 64.870 124.830 65.190 124.890 ;
        RECT 56.145 124.690 65.190 124.830 ;
        RECT 45.550 124.630 45.870 124.690 ;
        RECT 56.145 124.645 56.435 124.690 ;
        RECT 64.870 124.630 65.190 124.690 ;
        RECT 120.530 124.630 120.850 124.890 ;
        RECT 122.385 124.830 122.675 124.875 ;
        RECT 124.670 124.830 124.990 124.890 ;
        RECT 122.385 124.690 124.990 124.830 ;
        RECT 122.385 124.645 122.675 124.690 ;
        RECT 124.670 124.630 124.990 124.690 ;
        RECT 29.840 124.010 127.820 124.490 ;
        RECT 42.790 123.810 43.110 123.870 ;
        RECT 48.325 123.810 48.615 123.855 ;
        RECT 42.790 123.670 48.615 123.810 ;
        RECT 42.790 123.610 43.110 123.670 ;
        RECT 48.325 123.625 48.615 123.670 ;
        RECT 56.590 123.810 56.910 123.870 ;
        RECT 57.985 123.810 58.275 123.855 ;
        RECT 56.590 123.670 58.275 123.810 ;
        RECT 56.590 123.610 56.910 123.670 ;
        RECT 57.985 123.625 58.275 123.670 ;
        RECT 81.430 123.810 81.750 123.870 ;
        RECT 84.665 123.810 84.955 123.855 ;
        RECT 81.430 123.670 84.955 123.810 ;
        RECT 81.430 123.610 81.750 123.670 ;
        RECT 84.665 123.625 84.955 123.670 ;
        RECT 36.350 123.470 36.670 123.530 ;
        RECT 40.605 123.470 40.895 123.515 ;
        RECT 43.845 123.470 44.495 123.515 ;
        RECT 36.350 123.330 44.495 123.470 ;
        RECT 36.350 123.270 36.670 123.330 ;
        RECT 40.605 123.285 41.195 123.330 ;
        RECT 43.845 123.285 44.495 123.330 ;
        RECT 45.090 123.470 45.410 123.530 ;
        RECT 79.130 123.470 79.450 123.530 ;
        RECT 45.090 123.330 49.460 123.470 ;
        RECT 40.905 122.970 41.195 123.285 ;
        RECT 45.090 123.270 45.410 123.330 ;
        RECT 49.320 123.175 49.460 123.330 ;
        RECT 79.130 123.330 95.000 123.470 ;
        RECT 79.130 123.270 79.450 123.330 ;
        RECT 41.985 123.130 42.275 123.175 ;
        RECT 45.565 123.130 45.855 123.175 ;
        RECT 47.400 123.130 47.690 123.175 ;
        RECT 41.985 122.990 47.690 123.130 ;
        RECT 41.985 122.945 42.275 122.990 ;
        RECT 45.565 122.945 45.855 122.990 ;
        RECT 47.400 122.945 47.690 122.990 ;
        RECT 49.245 122.945 49.535 123.175 ;
        RECT 53.370 123.130 53.690 123.190 ;
        RECT 58.445 123.130 58.735 123.175 ;
        RECT 53.370 122.990 58.735 123.130 ;
        RECT 53.370 122.930 53.690 122.990 ;
        RECT 58.445 122.945 58.735 122.990 ;
        RECT 61.190 123.130 61.510 123.190 ;
        RECT 64.425 123.130 64.715 123.175 ;
        RECT 61.190 122.990 64.715 123.130 ;
        RECT 30.830 122.790 31.150 122.850 ;
        RECT 37.745 122.790 38.035 122.835 ;
        RECT 30.830 122.650 38.035 122.790 ;
        RECT 30.830 122.590 31.150 122.650 ;
        RECT 37.745 122.605 38.035 122.650 ;
        RECT 38.650 122.790 38.970 122.850 ;
        RECT 46.485 122.790 46.775 122.835 ;
        RECT 38.650 122.650 46.775 122.790 ;
        RECT 38.650 122.590 38.970 122.650 ;
        RECT 46.485 122.605 46.775 122.650 ;
        RECT 47.865 122.790 48.155 122.835 ;
        RECT 49.690 122.790 50.010 122.850 ;
        RECT 47.865 122.650 50.010 122.790 ;
        RECT 58.520 122.790 58.660 122.945 ;
        RECT 61.190 122.930 61.510 122.990 ;
        RECT 64.425 122.945 64.715 122.990 ;
        RECT 65.790 123.130 66.110 123.190 ;
        RECT 70.810 123.130 71.100 123.175 ;
        RECT 65.790 122.990 71.100 123.130 ;
        RECT 65.790 122.930 66.110 122.990 ;
        RECT 70.810 122.945 71.100 122.990 ;
        RECT 65.880 122.790 66.020 122.930 ;
        RECT 58.520 122.650 66.020 122.790 ;
        RECT 70.940 122.790 71.080 122.945 ;
        RECT 72.230 122.930 72.550 123.190 ;
        RECT 85.110 122.930 85.430 123.190 ;
        RECT 86.045 122.945 86.335 123.175 ;
        RECT 87.425 123.130 87.715 123.175 ;
        RECT 91.090 123.130 91.410 123.190 ;
        RECT 94.860 123.175 95.000 123.330 ;
        RECT 117.310 123.270 117.630 123.530 ;
        RECT 119.605 123.470 120.255 123.515 ;
        RECT 120.530 123.470 120.850 123.530 ;
        RECT 123.205 123.470 123.495 123.515 ;
        RECT 119.605 123.330 123.495 123.470 ;
        RECT 119.605 123.285 120.255 123.330 ;
        RECT 120.530 123.270 120.850 123.330 ;
        RECT 122.905 123.285 123.495 123.330 ;
        RECT 94.325 123.130 94.615 123.175 ;
        RECT 87.425 122.990 94.615 123.130 ;
        RECT 87.425 122.945 87.715 122.990 ;
        RECT 86.120 122.790 86.260 122.945 ;
        RECT 91.090 122.930 91.410 122.990 ;
        RECT 94.325 122.945 94.615 122.990 ;
        RECT 94.785 122.945 95.075 123.175 ;
        RECT 98.910 122.930 99.230 123.190 ;
        RECT 103.050 122.930 103.370 123.190 ;
        RECT 108.585 123.130 108.875 123.175 ;
        RECT 109.490 123.130 109.810 123.190 ;
        RECT 108.585 122.990 109.810 123.130 ;
        RECT 108.585 122.945 108.875 122.990 ;
        RECT 109.490 122.930 109.810 122.990 ;
        RECT 111.790 123.130 112.110 123.190 ;
        RECT 112.265 123.130 112.555 123.175 ;
        RECT 111.790 122.990 112.555 123.130 ;
        RECT 111.790 122.930 112.110 122.990 ;
        RECT 112.265 122.945 112.555 122.990 ;
        RECT 116.410 123.130 116.700 123.175 ;
        RECT 118.245 123.130 118.535 123.175 ;
        RECT 121.825 123.130 122.115 123.175 ;
        RECT 116.410 122.990 122.115 123.130 ;
        RECT 116.410 122.945 116.700 122.990 ;
        RECT 118.245 122.945 118.535 122.990 ;
        RECT 121.825 122.945 122.115 122.990 ;
        RECT 122.905 122.970 123.195 123.285 ;
        RECT 70.940 122.650 86.260 122.790 ;
        RECT 113.170 122.790 113.490 122.850 ;
        RECT 115.945 122.790 116.235 122.835 ;
        RECT 125.130 122.790 125.450 122.850 ;
        RECT 113.170 122.650 125.450 122.790 ;
        RECT 47.865 122.605 48.155 122.650 ;
        RECT 49.690 122.590 50.010 122.650 ;
        RECT 113.170 122.590 113.490 122.650 ;
        RECT 115.945 122.605 116.235 122.650 ;
        RECT 125.130 122.590 125.450 122.650 ;
        RECT 126.065 122.790 126.355 122.835 ;
        RECT 126.970 122.790 127.290 122.850 ;
        RECT 126.065 122.650 127.290 122.790 ;
        RECT 126.065 122.605 126.355 122.650 ;
        RECT 126.970 122.590 127.290 122.650 ;
        RECT 41.985 122.450 42.275 122.495 ;
        RECT 45.105 122.450 45.395 122.495 ;
        RECT 46.995 122.450 47.285 122.495 ;
        RECT 41.985 122.310 47.285 122.450 ;
        RECT 41.985 122.265 42.275 122.310 ;
        RECT 45.105 122.265 45.395 122.310 ;
        RECT 46.995 122.265 47.285 122.310 ;
        RECT 116.815 122.450 117.105 122.495 ;
        RECT 118.705 122.450 118.995 122.495 ;
        RECT 121.825 122.450 122.115 122.495 ;
        RECT 116.815 122.310 122.115 122.450 ;
        RECT 116.815 122.265 117.105 122.310 ;
        RECT 118.705 122.265 118.995 122.310 ;
        RECT 121.825 122.265 122.115 122.310 ;
        RECT 65.330 121.910 65.650 122.170 ;
        RECT 93.865 122.110 94.155 122.155 ;
        RECT 94.770 122.110 95.090 122.170 ;
        RECT 93.865 121.970 95.090 122.110 ;
        RECT 93.865 121.925 94.155 121.970 ;
        RECT 94.770 121.910 95.090 121.970 ;
        RECT 95.705 122.110 95.995 122.155 ;
        RECT 97.990 122.110 98.310 122.170 ;
        RECT 95.705 121.970 98.310 122.110 ;
        RECT 95.705 121.925 95.995 121.970 ;
        RECT 97.990 121.910 98.310 121.970 ;
        RECT 99.830 121.910 100.150 122.170 ;
        RECT 103.970 121.910 104.290 122.170 ;
        RECT 109.490 121.910 109.810 122.170 ;
        RECT 113.185 122.110 113.475 122.155 ;
        RECT 117.310 122.110 117.630 122.170 ;
        RECT 113.185 121.970 117.630 122.110 ;
        RECT 113.185 121.925 113.475 121.970 ;
        RECT 117.310 121.910 117.630 121.970 ;
        RECT 29.840 121.290 127.820 121.770 ;
        RECT 37.745 121.090 38.035 121.135 ;
        RECT 38.650 121.090 38.970 121.150 ;
        RECT 37.745 120.950 38.970 121.090 ;
        RECT 37.745 120.905 38.035 120.950 ;
        RECT 38.650 120.890 38.970 120.950 ;
        RECT 44.630 121.090 44.950 121.150 ;
        RECT 55.685 121.090 55.975 121.135 ;
        RECT 44.630 120.950 55.975 121.090 ;
        RECT 44.630 120.890 44.950 120.950 ;
        RECT 55.685 120.905 55.975 120.950 ;
        RECT 42.330 120.750 42.650 120.810 ;
        RECT 36.900 120.610 42.650 120.750 ;
        RECT 36.900 120.115 37.040 120.610 ;
        RECT 42.330 120.550 42.650 120.610 ;
        RECT 43.825 120.750 44.115 120.795 ;
        RECT 46.945 120.750 47.235 120.795 ;
        RECT 48.835 120.750 49.125 120.795 ;
        RECT 50.625 120.750 50.915 120.795 ;
        RECT 43.825 120.610 49.125 120.750 ;
        RECT 43.825 120.565 44.115 120.610 ;
        RECT 46.945 120.565 47.235 120.610 ;
        RECT 48.835 120.565 49.125 120.610 ;
        RECT 49.320 120.610 50.915 120.750 ;
        RECT 39.585 120.410 39.875 120.455 ;
        RECT 46.010 120.410 46.330 120.470 ;
        RECT 39.585 120.270 46.330 120.410 ;
        RECT 39.585 120.225 39.875 120.270 ;
        RECT 46.010 120.210 46.330 120.270 ;
        RECT 48.325 120.410 48.615 120.455 ;
        RECT 49.320 120.410 49.460 120.610 ;
        RECT 50.625 120.565 50.915 120.610 ;
        RECT 62.685 120.750 62.975 120.795 ;
        RECT 65.805 120.750 66.095 120.795 ;
        RECT 67.695 120.750 67.985 120.795 ;
        RECT 62.685 120.610 67.985 120.750 ;
        RECT 62.685 120.565 62.975 120.610 ;
        RECT 65.805 120.565 66.095 120.610 ;
        RECT 67.695 120.565 67.985 120.610 ;
        RECT 83.385 120.750 83.675 120.795 ;
        RECT 86.505 120.750 86.795 120.795 ;
        RECT 88.395 120.750 88.685 120.795 ;
        RECT 83.385 120.610 88.685 120.750 ;
        RECT 83.385 120.565 83.675 120.610 ;
        RECT 86.505 120.565 86.795 120.610 ;
        RECT 88.395 120.565 88.685 120.610 ;
        RECT 95.345 120.750 95.635 120.795 ;
        RECT 98.465 120.750 98.755 120.795 ;
        RECT 100.355 120.750 100.645 120.795 ;
        RECT 95.345 120.610 100.645 120.750 ;
        RECT 95.345 120.565 95.635 120.610 ;
        RECT 98.465 120.565 98.755 120.610 ;
        RECT 100.355 120.565 100.645 120.610 ;
        RECT 107.305 120.750 107.595 120.795 ;
        RECT 110.425 120.750 110.715 120.795 ;
        RECT 112.315 120.750 112.605 120.795 ;
        RECT 107.305 120.610 112.605 120.750 ;
        RECT 107.305 120.565 107.595 120.610 ;
        RECT 110.425 120.565 110.715 120.610 ;
        RECT 112.315 120.565 112.605 120.610 ;
        RECT 120.185 120.750 120.475 120.795 ;
        RECT 123.305 120.750 123.595 120.795 ;
        RECT 125.195 120.750 125.485 120.795 ;
        RECT 120.185 120.610 125.485 120.750 ;
        RECT 120.185 120.565 120.475 120.610 ;
        RECT 123.305 120.565 123.595 120.610 ;
        RECT 125.195 120.565 125.485 120.610 ;
        RECT 48.325 120.270 49.460 120.410 ;
        RECT 48.325 120.225 48.615 120.270 ;
        RECT 49.690 120.210 50.010 120.470 ;
        RECT 50.150 120.410 50.470 120.470 ;
        RECT 53.385 120.410 53.675 120.455 ;
        RECT 50.150 120.270 53.675 120.410 ;
        RECT 50.150 120.210 50.470 120.270 ;
        RECT 53.385 120.225 53.675 120.270 ;
        RECT 55.210 120.410 55.530 120.470 ;
        RECT 58.445 120.410 58.735 120.455 ;
        RECT 61.190 120.410 61.510 120.470 ;
        RECT 55.210 120.270 57.280 120.410 ;
        RECT 55.210 120.210 55.530 120.270 ;
        RECT 36.825 119.885 37.115 120.115 ;
        RECT 38.205 120.070 38.495 120.115 ;
        RECT 41.870 120.070 42.190 120.130 ;
        RECT 38.205 119.930 42.190 120.070 ;
        RECT 38.205 119.885 38.495 119.930 ;
        RECT 41.870 119.870 42.190 119.930 ;
        RECT 40.950 119.730 41.270 119.790 ;
        RECT 42.745 119.775 43.035 120.090 ;
        RECT 43.825 120.070 44.115 120.115 ;
        RECT 47.405 120.070 47.695 120.115 ;
        RECT 49.240 120.070 49.530 120.115 ;
        RECT 51.545 120.070 51.835 120.115 ;
        RECT 43.825 119.930 49.530 120.070 ;
        RECT 43.825 119.885 44.115 119.930 ;
        RECT 47.405 119.885 47.695 119.930 ;
        RECT 49.240 119.885 49.530 119.930 ;
        RECT 50.240 119.930 51.835 120.070 ;
        RECT 42.445 119.730 43.035 119.775 ;
        RECT 45.685 119.730 46.335 119.775 ;
        RECT 40.950 119.590 46.335 119.730 ;
        RECT 40.950 119.530 41.270 119.590 ;
        RECT 42.445 119.545 42.735 119.590 ;
        RECT 45.685 119.545 46.335 119.590 ;
        RECT 39.125 119.390 39.415 119.435 ;
        RECT 41.870 119.390 42.190 119.450 ;
        RECT 39.125 119.250 42.190 119.390 ;
        RECT 39.125 119.205 39.415 119.250 ;
        RECT 41.870 119.190 42.190 119.250 ;
        RECT 49.230 119.390 49.550 119.450 ;
        RECT 50.240 119.390 50.380 119.930 ;
        RECT 51.545 119.885 51.835 119.930 ;
        RECT 53.830 119.870 54.150 120.130 ;
        RECT 54.750 120.070 55.070 120.130 ;
        RECT 57.140 120.115 57.280 120.270 ;
        RECT 58.445 120.270 61.510 120.410 ;
        RECT 58.445 120.225 58.735 120.270 ;
        RECT 61.190 120.210 61.510 120.270 ;
        RECT 65.330 120.410 65.650 120.470 ;
        RECT 67.185 120.410 67.475 120.455 ;
        RECT 65.330 120.270 67.475 120.410 ;
        RECT 65.330 120.210 65.650 120.270 ;
        RECT 67.185 120.225 67.475 120.270 ;
        RECT 69.470 120.410 69.790 120.470 ;
        RECT 84.650 120.410 84.970 120.470 ;
        RECT 91.105 120.410 91.395 120.455 ;
        RECT 96.610 120.410 96.930 120.470 ;
        RECT 69.470 120.270 73.840 120.410 ;
        RECT 69.470 120.210 69.790 120.270 ;
        RECT 56.605 120.070 56.895 120.115 ;
        RECT 54.750 119.930 56.895 120.070 ;
        RECT 54.750 119.870 55.070 119.930 ;
        RECT 56.605 119.885 56.895 119.930 ;
        RECT 57.065 119.885 57.355 120.115 ;
        RECT 61.605 119.775 61.895 120.090 ;
        RECT 62.685 120.070 62.975 120.115 ;
        RECT 66.265 120.070 66.555 120.115 ;
        RECT 68.100 120.070 68.390 120.115 ;
        RECT 62.685 119.930 68.390 120.070 ;
        RECT 62.685 119.885 62.975 119.930 ;
        RECT 66.265 119.885 66.555 119.930 ;
        RECT 68.100 119.885 68.390 119.930 ;
        RECT 68.550 119.870 68.870 120.130 ;
        RECT 69.010 119.870 69.330 120.130 ;
        RECT 70.865 120.070 71.155 120.115 ;
        RECT 72.230 120.070 72.550 120.130 ;
        RECT 73.700 120.115 73.840 120.270 ;
        RECT 84.650 120.270 89.940 120.410 ;
        RECT 84.650 120.210 84.970 120.270 ;
        RECT 69.560 119.930 72.550 120.070 ;
        RECT 61.305 119.730 61.895 119.775 ;
        RECT 63.950 119.730 64.270 119.790 ;
        RECT 64.545 119.730 65.195 119.775 ;
        RECT 61.305 119.590 65.195 119.730 ;
        RECT 61.305 119.545 61.595 119.590 ;
        RECT 63.950 119.530 64.270 119.590 ;
        RECT 64.545 119.545 65.195 119.590 ;
        RECT 49.230 119.250 50.380 119.390 ;
        RECT 57.985 119.390 58.275 119.435 ;
        RECT 59.810 119.390 60.130 119.450 ;
        RECT 57.985 119.250 60.130 119.390 ;
        RECT 49.230 119.190 49.550 119.250 ;
        RECT 57.985 119.205 58.275 119.250 ;
        RECT 59.810 119.190 60.130 119.250 ;
        RECT 66.250 119.390 66.570 119.450 ;
        RECT 69.560 119.390 69.700 119.930 ;
        RECT 70.865 119.885 71.155 119.930 ;
        RECT 72.230 119.870 72.550 119.930 ;
        RECT 73.625 119.885 73.915 120.115 ;
        RECT 74.070 120.070 74.390 120.130 ;
        RECT 77.765 120.070 78.055 120.115 ;
        RECT 74.070 119.930 78.055 120.070 ;
        RECT 74.070 119.870 74.390 119.930 ;
        RECT 77.765 119.885 78.055 119.930 ;
        RECT 70.390 119.730 70.710 119.790 ;
        RECT 72.705 119.730 72.995 119.775 ;
        RECT 70.390 119.590 72.995 119.730 ;
        RECT 70.390 119.530 70.710 119.590 ;
        RECT 72.705 119.545 72.995 119.590 ;
        RECT 79.145 119.730 79.435 119.775 ;
        RECT 81.430 119.730 81.750 119.790 ;
        RECT 82.305 119.775 82.595 120.090 ;
        RECT 83.385 120.070 83.675 120.115 ;
        RECT 86.965 120.070 87.255 120.115 ;
        RECT 88.800 120.070 89.090 120.115 ;
        RECT 83.385 119.930 89.090 120.070 ;
        RECT 83.385 119.885 83.675 119.930 ;
        RECT 86.965 119.885 87.255 119.930 ;
        RECT 88.800 119.885 89.090 119.930 ;
        RECT 89.250 119.870 89.570 120.130 ;
        RECT 89.800 120.115 89.940 120.270 ;
        RECT 91.105 120.270 96.930 120.410 ;
        RECT 91.105 120.225 91.395 120.270 ;
        RECT 96.610 120.210 96.930 120.270 ;
        RECT 99.830 120.210 100.150 120.470 ;
        RECT 103.065 120.410 103.355 120.455 ;
        RECT 105.810 120.410 106.130 120.470 ;
        RECT 103.065 120.270 106.130 120.410 ;
        RECT 103.065 120.225 103.355 120.270 ;
        RECT 105.810 120.210 106.130 120.270 ;
        RECT 109.490 120.410 109.810 120.470 ;
        RECT 111.805 120.410 112.095 120.455 ;
        RECT 109.490 120.270 112.095 120.410 ;
        RECT 109.490 120.210 109.810 120.270 ;
        RECT 111.805 120.225 112.095 120.270 ;
        RECT 115.945 120.410 116.235 120.455 ;
        RECT 121.450 120.410 121.770 120.470 ;
        RECT 115.945 120.270 121.770 120.410 ;
        RECT 115.945 120.225 116.235 120.270 ;
        RECT 121.450 120.210 121.770 120.270 ;
        RECT 124.670 120.210 124.990 120.470 ;
        RECT 89.725 119.885 90.015 120.115 ;
        RECT 79.145 119.590 81.750 119.730 ;
        RECT 79.145 119.545 79.435 119.590 ;
        RECT 81.430 119.530 81.750 119.590 ;
        RECT 82.005 119.730 82.595 119.775 ;
        RECT 84.650 119.730 84.970 119.790 ;
        RECT 85.245 119.730 85.895 119.775 ;
        RECT 82.005 119.590 85.895 119.730 ;
        RECT 82.005 119.545 82.295 119.590 ;
        RECT 84.650 119.530 84.970 119.590 ;
        RECT 85.245 119.545 85.895 119.590 ;
        RECT 86.490 119.730 86.810 119.790 ;
        RECT 94.265 119.775 94.555 120.090 ;
        RECT 95.345 120.070 95.635 120.115 ;
        RECT 98.925 120.070 99.215 120.115 ;
        RECT 100.760 120.070 101.050 120.115 ;
        RECT 95.345 119.930 101.050 120.070 ;
        RECT 95.345 119.885 95.635 119.930 ;
        RECT 98.925 119.885 99.215 119.930 ;
        RECT 100.760 119.885 101.050 119.930 ;
        RECT 101.210 119.870 101.530 120.130 ;
        RECT 97.530 119.775 97.850 119.790 ;
        RECT 106.225 119.775 106.515 120.090 ;
        RECT 107.305 120.070 107.595 120.115 ;
        RECT 110.885 120.070 111.175 120.115 ;
        RECT 112.720 120.070 113.010 120.115 ;
        RECT 107.305 119.930 113.010 120.070 ;
        RECT 107.305 119.885 107.595 119.930 ;
        RECT 110.885 119.885 111.175 119.930 ;
        RECT 112.720 119.885 113.010 119.930 ;
        RECT 113.170 119.870 113.490 120.130 ;
        RECT 114.565 119.885 114.855 120.115 ;
        RECT 119.150 120.090 119.470 120.130 ;
        RECT 109.490 119.775 109.810 119.790 ;
        RECT 87.885 119.730 88.175 119.775 ;
        RECT 86.490 119.590 88.175 119.730 ;
        RECT 86.490 119.530 86.810 119.590 ;
        RECT 87.885 119.545 88.175 119.590 ;
        RECT 93.965 119.730 94.555 119.775 ;
        RECT 97.205 119.730 97.855 119.775 ;
        RECT 93.965 119.590 97.855 119.730 ;
        RECT 93.965 119.545 94.255 119.590 ;
        RECT 97.205 119.545 97.855 119.590 ;
        RECT 105.925 119.730 106.515 119.775 ;
        RECT 109.165 119.730 109.815 119.775 ;
        RECT 105.925 119.590 109.815 119.730 ;
        RECT 105.925 119.545 106.215 119.590 ;
        RECT 109.165 119.545 109.815 119.590 ;
        RECT 110.410 119.730 110.730 119.790 ;
        RECT 114.640 119.730 114.780 119.885 ;
        RECT 119.105 119.870 119.470 120.090 ;
        RECT 120.185 120.070 120.475 120.115 ;
        RECT 123.765 120.070 124.055 120.115 ;
        RECT 125.600 120.070 125.890 120.115 ;
        RECT 120.185 119.930 125.890 120.070 ;
        RECT 120.185 119.885 120.475 119.930 ;
        RECT 123.765 119.885 124.055 119.930 ;
        RECT 125.600 119.885 125.890 119.930 ;
        RECT 126.065 119.885 126.355 120.115 ;
        RECT 119.105 119.775 119.395 119.870 ;
        RECT 110.410 119.590 114.780 119.730 ;
        RECT 118.805 119.730 119.395 119.775 ;
        RECT 122.045 119.730 122.695 119.775 ;
        RECT 118.805 119.590 122.695 119.730 ;
        RECT 97.530 119.530 97.850 119.545 ;
        RECT 109.490 119.530 109.810 119.545 ;
        RECT 110.410 119.530 110.730 119.590 ;
        RECT 118.805 119.545 119.095 119.590 ;
        RECT 122.045 119.545 122.695 119.590 ;
        RECT 125.130 119.730 125.450 119.790 ;
        RECT 126.140 119.730 126.280 119.885 ;
        RECT 125.130 119.590 126.280 119.730 ;
        RECT 125.130 119.530 125.450 119.590 ;
        RECT 66.250 119.250 69.700 119.390 ;
        RECT 69.945 119.390 70.235 119.435 ;
        RECT 70.850 119.390 71.170 119.450 ;
        RECT 69.945 119.250 71.170 119.390 ;
        RECT 66.250 119.190 66.570 119.250 ;
        RECT 69.945 119.205 70.235 119.250 ;
        RECT 70.850 119.190 71.170 119.250 ;
        RECT 71.325 119.390 71.615 119.435 ;
        RECT 73.610 119.390 73.930 119.450 ;
        RECT 71.325 119.250 73.930 119.390 ;
        RECT 71.325 119.205 71.615 119.250 ;
        RECT 73.610 119.190 73.930 119.250 ;
        RECT 74.070 119.390 74.390 119.450 ;
        RECT 74.545 119.390 74.835 119.435 ;
        RECT 74.070 119.250 74.835 119.390 ;
        RECT 74.070 119.190 74.390 119.250 ;
        RECT 74.545 119.205 74.835 119.250 ;
        RECT 78.685 119.390 78.975 119.435 ;
        RECT 82.810 119.390 83.130 119.450 ;
        RECT 78.685 119.250 83.130 119.390 ;
        RECT 78.685 119.205 78.975 119.250 ;
        RECT 82.810 119.190 83.130 119.250 ;
        RECT 90.630 119.190 90.950 119.450 ;
        RECT 112.710 119.390 113.030 119.450 ;
        RECT 113.645 119.390 113.935 119.435 ;
        RECT 112.710 119.250 113.935 119.390 ;
        RECT 112.710 119.190 113.030 119.250 ;
        RECT 113.645 119.205 113.935 119.250 ;
        RECT 29.840 118.570 127.820 119.050 ;
        RECT 35.905 118.370 36.195 118.415 ;
        RECT 36.350 118.370 36.670 118.430 ;
        RECT 35.905 118.230 36.670 118.370 ;
        RECT 35.905 118.185 36.195 118.230 ;
        RECT 36.350 118.170 36.670 118.230 ;
        RECT 37.730 118.370 38.050 118.430 ;
        RECT 38.205 118.370 38.495 118.415 ;
        RECT 37.730 118.230 38.495 118.370 ;
        RECT 37.730 118.170 38.050 118.230 ;
        RECT 38.205 118.185 38.495 118.230 ;
        RECT 40.950 118.170 41.270 118.430 ;
        RECT 53.830 118.370 54.150 118.430 ;
        RECT 41.960 118.230 54.150 118.370 ;
        RECT 36.365 117.690 36.655 117.735 ;
        RECT 37.745 117.690 38.035 117.735 ;
        RECT 39.125 117.690 39.415 117.735 ;
        RECT 40.505 117.690 40.795 117.735 ;
        RECT 41.960 117.690 42.100 118.230 ;
        RECT 53.830 118.170 54.150 118.230 ;
        RECT 86.045 118.370 86.335 118.415 ;
        RECT 86.490 118.370 86.810 118.430 ;
        RECT 86.045 118.230 86.810 118.370 ;
        RECT 86.045 118.185 86.335 118.230 ;
        RECT 86.490 118.170 86.810 118.230 ;
        RECT 90.630 118.370 90.950 118.430 ;
        RECT 103.970 118.370 104.290 118.430 ;
        RECT 109.490 118.370 109.810 118.430 ;
        RECT 110.885 118.370 111.175 118.415 ;
        RECT 119.610 118.370 119.930 118.430 ;
        RECT 90.630 118.230 98.220 118.370 ;
        RECT 90.630 118.170 90.950 118.230 ;
        RECT 43.265 118.030 43.555 118.075 ;
        RECT 44.630 118.030 44.950 118.090 ;
        RECT 43.265 117.890 44.950 118.030 ;
        RECT 43.265 117.845 43.555 117.890 ;
        RECT 44.630 117.830 44.950 117.890 ;
        RECT 45.545 118.030 46.195 118.075 ;
        RECT 49.145 118.030 49.435 118.075 ;
        RECT 50.150 118.030 50.470 118.090 ;
        RECT 45.545 117.890 50.470 118.030 ;
        RECT 45.545 117.845 46.195 117.890 ;
        RECT 48.845 117.845 49.435 117.890 ;
        RECT 36.365 117.550 42.100 117.690 ;
        RECT 42.350 117.690 42.640 117.735 ;
        RECT 44.185 117.690 44.475 117.735 ;
        RECT 47.765 117.690 48.055 117.735 ;
        RECT 42.350 117.550 48.055 117.690 ;
        RECT 36.365 117.505 36.655 117.550 ;
        RECT 37.745 117.505 38.035 117.550 ;
        RECT 39.125 117.505 39.415 117.550 ;
        RECT 40.505 117.505 40.795 117.550 ;
        RECT 42.350 117.505 42.640 117.550 ;
        RECT 44.185 117.505 44.475 117.550 ;
        RECT 47.765 117.505 48.055 117.550 ;
        RECT 48.845 117.530 49.135 117.845 ;
        RECT 50.150 117.830 50.470 117.890 ;
        RECT 55.325 118.030 55.615 118.075 ;
        RECT 57.970 118.030 58.290 118.090 ;
        RECT 58.565 118.030 59.215 118.075 ;
        RECT 55.325 117.890 59.215 118.030 ;
        RECT 55.325 117.845 55.915 117.890 ;
        RECT 55.625 117.530 55.915 117.845 ;
        RECT 57.970 117.830 58.290 117.890 ;
        RECT 58.565 117.845 59.215 117.890 ;
        RECT 59.810 118.030 60.130 118.090 ;
        RECT 61.205 118.030 61.495 118.075 ;
        RECT 59.810 117.890 61.495 118.030 ;
        RECT 59.810 117.830 60.130 117.890 ;
        RECT 61.205 117.845 61.495 117.890 ;
        RECT 64.410 118.030 64.730 118.090 ;
        RECT 66.365 118.030 66.655 118.075 ;
        RECT 69.605 118.030 70.255 118.075 ;
        RECT 64.410 117.890 70.255 118.030 ;
        RECT 64.410 117.830 64.730 117.890 ;
        RECT 66.365 117.845 66.955 117.890 ;
        RECT 69.605 117.845 70.255 117.890 ;
        RECT 70.850 118.030 71.170 118.090 ;
        RECT 72.245 118.030 72.535 118.075 ;
        RECT 70.850 117.890 72.535 118.030 ;
        RECT 56.705 117.690 56.995 117.735 ;
        RECT 60.285 117.690 60.575 117.735 ;
        RECT 62.120 117.690 62.410 117.735 ;
        RECT 56.705 117.550 62.410 117.690 ;
        RECT 56.705 117.505 56.995 117.550 ;
        RECT 60.285 117.505 60.575 117.550 ;
        RECT 62.120 117.505 62.410 117.550 ;
        RECT 63.505 117.690 63.795 117.735 ;
        RECT 65.790 117.690 66.110 117.750 ;
        RECT 63.505 117.550 66.110 117.690 ;
        RECT 63.505 117.505 63.795 117.550 ;
        RECT 65.790 117.490 66.110 117.550 ;
        RECT 66.665 117.530 66.955 117.845 ;
        RECT 70.850 117.830 71.170 117.890 ;
        RECT 72.245 117.845 72.535 117.890 ;
        RECT 73.610 118.030 73.930 118.090 ;
        RECT 76.945 118.030 77.235 118.075 ;
        RECT 80.185 118.030 80.835 118.075 ;
        RECT 73.610 117.890 80.835 118.030 ;
        RECT 73.610 117.830 73.930 117.890 ;
        RECT 76.945 117.845 77.535 117.890 ;
        RECT 80.185 117.845 80.835 117.890 ;
        RECT 67.745 117.690 68.035 117.735 ;
        RECT 71.325 117.690 71.615 117.735 ;
        RECT 73.160 117.690 73.450 117.735 ;
        RECT 67.745 117.550 73.450 117.690 ;
        RECT 67.745 117.505 68.035 117.550 ;
        RECT 71.325 117.505 71.615 117.550 ;
        RECT 73.160 117.505 73.450 117.550 ;
        RECT 74.085 117.690 74.375 117.735 ;
        RECT 76.370 117.690 76.690 117.750 ;
        RECT 74.085 117.550 76.690 117.690 ;
        RECT 74.085 117.505 74.375 117.550 ;
        RECT 76.370 117.490 76.690 117.550 ;
        RECT 77.245 117.530 77.535 117.845 ;
        RECT 82.810 117.830 83.130 118.090 ;
        RECT 84.650 118.030 84.970 118.090 ;
        RECT 86.965 118.030 87.255 118.075 ;
        RECT 84.650 117.890 87.255 118.030 ;
        RECT 84.650 117.830 84.970 117.890 ;
        RECT 86.965 117.845 87.255 117.890 ;
        RECT 88.330 118.030 88.650 118.090 ;
        RECT 98.080 118.075 98.220 118.230 ;
        RECT 103.970 118.230 108.800 118.370 ;
        RECT 103.970 118.170 104.290 118.230 ;
        RECT 108.660 118.075 108.800 118.230 ;
        RECT 109.490 118.230 111.175 118.370 ;
        RECT 109.490 118.170 109.810 118.230 ;
        RECT 110.885 118.185 111.175 118.230 ;
        RECT 112.800 118.230 119.930 118.370 ;
        RECT 89.265 118.030 89.555 118.075 ;
        RECT 88.330 117.890 89.555 118.030 ;
        RECT 88.330 117.830 88.650 117.890 ;
        RECT 89.265 117.845 89.555 117.890 ;
        RECT 92.125 118.030 92.415 118.075 ;
        RECT 95.365 118.030 96.015 118.075 ;
        RECT 92.125 117.890 96.015 118.030 ;
        RECT 92.125 117.845 92.715 117.890 ;
        RECT 95.365 117.845 96.015 117.890 ;
        RECT 98.005 117.845 98.295 118.075 ;
        RECT 102.705 118.030 102.995 118.075 ;
        RECT 105.945 118.030 106.595 118.075 ;
        RECT 102.705 117.890 106.595 118.030 ;
        RECT 102.705 117.845 103.295 117.890 ;
        RECT 105.945 117.845 106.595 117.890 ;
        RECT 108.585 117.845 108.875 118.075 ;
        RECT 78.325 117.690 78.615 117.735 ;
        RECT 81.905 117.690 82.195 117.735 ;
        RECT 83.740 117.690 84.030 117.735 ;
        RECT 78.325 117.550 84.030 117.690 ;
        RECT 78.325 117.505 78.615 117.550 ;
        RECT 81.905 117.505 82.195 117.550 ;
        RECT 83.740 117.505 84.030 117.550 ;
        RECT 85.125 117.690 85.415 117.735 ;
        RECT 85.570 117.690 85.890 117.750 ;
        RECT 85.125 117.550 85.890 117.690 ;
        RECT 85.125 117.505 85.415 117.550 ;
        RECT 85.570 117.490 85.890 117.550 ;
        RECT 87.410 117.490 87.730 117.750 ;
        RECT 87.870 117.690 88.190 117.750 ;
        RECT 92.425 117.690 92.715 117.845 ;
        RECT 103.005 117.750 103.295 117.845 ;
        RECT 87.870 117.550 92.715 117.690 ;
        RECT 87.870 117.490 88.190 117.550 ;
        RECT 92.425 117.530 92.715 117.550 ;
        RECT 93.505 117.690 93.795 117.735 ;
        RECT 97.085 117.690 97.375 117.735 ;
        RECT 98.920 117.690 99.210 117.735 ;
        RECT 93.505 117.550 99.210 117.690 ;
        RECT 93.505 117.505 93.795 117.550 ;
        RECT 97.085 117.505 97.375 117.550 ;
        RECT 98.920 117.505 99.210 117.550 ;
        RECT 99.845 117.690 100.135 117.735 ;
        RECT 101.670 117.690 101.990 117.750 ;
        RECT 99.845 117.550 101.990 117.690 ;
        RECT 99.845 117.505 100.135 117.550 ;
        RECT 101.670 117.490 101.990 117.550 ;
        RECT 103.005 117.530 103.370 117.750 ;
        RECT 103.050 117.490 103.370 117.530 ;
        RECT 104.085 117.690 104.375 117.735 ;
        RECT 107.665 117.690 107.955 117.735 ;
        RECT 109.500 117.690 109.790 117.735 ;
        RECT 104.085 117.550 109.790 117.690 ;
        RECT 104.085 117.505 104.375 117.550 ;
        RECT 107.665 117.505 107.955 117.550 ;
        RECT 109.500 117.505 109.790 117.550 ;
        RECT 110.410 117.690 110.730 117.750 ;
        RECT 112.800 117.735 112.940 118.230 ;
        RECT 119.610 118.170 119.930 118.230 ;
        RECT 117.885 118.030 118.175 118.075 ;
        RECT 121.125 118.030 121.775 118.075 ;
        RECT 117.885 117.890 121.775 118.030 ;
        RECT 117.885 117.845 118.475 117.890 ;
        RECT 121.125 117.845 121.775 117.890 ;
        RECT 118.185 117.750 118.475 117.845 ;
        RECT 111.345 117.690 111.635 117.735 ;
        RECT 112.725 117.690 113.015 117.735 ;
        RECT 110.410 117.550 113.015 117.690 ;
        RECT 110.410 117.490 110.730 117.550 ;
        RECT 111.345 117.505 111.635 117.550 ;
        RECT 112.725 117.505 113.015 117.550 ;
        RECT 118.185 117.530 118.550 117.750 ;
        RECT 118.230 117.490 118.550 117.530 ;
        RECT 119.265 117.690 119.555 117.735 ;
        RECT 122.845 117.690 123.135 117.735 ;
        RECT 124.680 117.690 124.970 117.735 ;
        RECT 119.265 117.550 124.970 117.690 ;
        RECT 119.265 117.505 119.555 117.550 ;
        RECT 122.845 117.505 123.135 117.550 ;
        RECT 124.680 117.505 124.970 117.550 ;
        RECT 125.130 117.490 125.450 117.750 ;
        RECT 41.885 117.350 42.175 117.395 ;
        RECT 49.690 117.350 50.010 117.410 ;
        RECT 41.885 117.210 50.010 117.350 ;
        RECT 41.885 117.165 42.175 117.210 ;
        RECT 49.690 117.150 50.010 117.210 ;
        RECT 51.070 117.350 51.390 117.410 ;
        RECT 52.005 117.350 52.295 117.395 ;
        RECT 51.070 117.210 52.295 117.350 ;
        RECT 51.070 117.150 51.390 117.210 ;
        RECT 52.005 117.165 52.295 117.210 ;
        RECT 52.465 117.350 52.755 117.395 ;
        RECT 56.130 117.350 56.450 117.410 ;
        RECT 52.465 117.210 56.450 117.350 ;
        RECT 52.465 117.165 52.755 117.210 ;
        RECT 56.130 117.150 56.450 117.210 ;
        RECT 62.585 117.350 62.875 117.395 ;
        RECT 68.550 117.350 68.870 117.410 ;
        RECT 73.625 117.350 73.915 117.395 ;
        RECT 75.450 117.350 75.770 117.410 ;
        RECT 62.585 117.210 75.770 117.350 ;
        RECT 62.585 117.165 62.875 117.210 ;
        RECT 68.550 117.150 68.870 117.210 ;
        RECT 73.625 117.165 73.915 117.210 ;
        RECT 75.450 117.150 75.770 117.210 ;
        RECT 84.205 117.350 84.495 117.395 ;
        RECT 89.250 117.350 89.570 117.410 ;
        RECT 99.370 117.350 99.690 117.410 ;
        RECT 101.210 117.350 101.530 117.410 ;
        RECT 109.965 117.350 110.255 117.395 ;
        RECT 113.170 117.350 113.490 117.410 ;
        RECT 84.205 117.210 113.490 117.350 ;
        RECT 84.205 117.165 84.495 117.210 ;
        RECT 89.250 117.150 89.570 117.210 ;
        RECT 99.370 117.150 99.690 117.210 ;
        RECT 101.210 117.150 101.530 117.210 ;
        RECT 109.965 117.165 110.255 117.210 ;
        RECT 113.170 117.150 113.490 117.210 ;
        RECT 115.025 117.350 115.315 117.395 ;
        RECT 116.850 117.350 117.170 117.410 ;
        RECT 115.025 117.210 117.170 117.350 ;
        RECT 115.025 117.165 115.315 117.210 ;
        RECT 116.850 117.150 117.170 117.210 ;
        RECT 117.310 117.350 117.630 117.410 ;
        RECT 123.765 117.350 124.055 117.395 ;
        RECT 117.310 117.210 124.055 117.350 ;
        RECT 117.310 117.150 117.630 117.210 ;
        RECT 123.765 117.165 124.055 117.210 ;
        RECT 42.755 117.010 43.045 117.055 ;
        RECT 44.645 117.010 44.935 117.055 ;
        RECT 47.765 117.010 48.055 117.055 ;
        RECT 42.755 116.870 48.055 117.010 ;
        RECT 42.755 116.825 43.045 116.870 ;
        RECT 44.645 116.825 44.935 116.870 ;
        RECT 47.765 116.825 48.055 116.870 ;
        RECT 56.705 117.010 56.995 117.055 ;
        RECT 59.825 117.010 60.115 117.055 ;
        RECT 61.715 117.010 62.005 117.055 ;
        RECT 56.705 116.870 62.005 117.010 ;
        RECT 56.705 116.825 56.995 116.870 ;
        RECT 59.825 116.825 60.115 116.870 ;
        RECT 61.715 116.825 62.005 116.870 ;
        RECT 67.745 117.010 68.035 117.055 ;
        RECT 70.865 117.010 71.155 117.055 ;
        RECT 72.755 117.010 73.045 117.055 ;
        RECT 67.745 116.870 73.045 117.010 ;
        RECT 67.745 116.825 68.035 116.870 ;
        RECT 70.865 116.825 71.155 116.870 ;
        RECT 72.755 116.825 73.045 116.870 ;
        RECT 78.325 117.010 78.615 117.055 ;
        RECT 81.445 117.010 81.735 117.055 ;
        RECT 83.335 117.010 83.625 117.055 ;
        RECT 78.325 116.870 83.625 117.010 ;
        RECT 78.325 116.825 78.615 116.870 ;
        RECT 81.445 116.825 81.735 116.870 ;
        RECT 83.335 116.825 83.625 116.870 ;
        RECT 93.505 117.010 93.795 117.055 ;
        RECT 96.625 117.010 96.915 117.055 ;
        RECT 98.515 117.010 98.805 117.055 ;
        RECT 93.505 116.870 98.805 117.010 ;
        RECT 93.505 116.825 93.795 116.870 ;
        RECT 96.625 116.825 96.915 116.870 ;
        RECT 98.515 116.825 98.805 116.870 ;
        RECT 104.085 117.010 104.375 117.055 ;
        RECT 107.205 117.010 107.495 117.055 ;
        RECT 109.095 117.010 109.385 117.055 ;
        RECT 104.085 116.870 109.385 117.010 ;
        RECT 104.085 116.825 104.375 116.870 ;
        RECT 107.205 116.825 107.495 116.870 ;
        RECT 109.095 116.825 109.385 116.870 ;
        RECT 119.265 117.010 119.555 117.055 ;
        RECT 122.385 117.010 122.675 117.055 ;
        RECT 124.275 117.010 124.565 117.055 ;
        RECT 119.265 116.870 124.565 117.010 ;
        RECT 119.265 116.825 119.555 116.870 ;
        RECT 122.385 116.825 122.675 116.870 ;
        RECT 124.275 116.825 124.565 116.870 ;
        RECT 39.570 116.470 39.890 116.730 ;
        RECT 85.110 116.670 85.430 116.730 ;
        RECT 103.510 116.670 103.830 116.730 ;
        RECT 85.110 116.530 103.830 116.670 ;
        RECT 85.110 116.470 85.430 116.530 ;
        RECT 103.510 116.470 103.830 116.530 ;
        RECT 112.250 116.470 112.570 116.730 ;
        RECT 29.840 115.850 127.820 116.330 ;
        RECT 57.970 115.450 58.290 115.710 ;
        RECT 62.125 115.650 62.415 115.695 ;
        RECT 63.950 115.650 64.270 115.710 ;
        RECT 62.125 115.510 64.270 115.650 ;
        RECT 62.125 115.465 62.415 115.510 ;
        RECT 63.950 115.450 64.270 115.510 ;
        RECT 64.410 115.450 64.730 115.710 ;
        RECT 87.870 115.450 88.190 115.710 ;
        RECT 97.530 115.650 97.850 115.710 ;
        RECT 100.305 115.650 100.595 115.695 ;
        RECT 97.530 115.510 100.595 115.650 ;
        RECT 97.530 115.450 97.850 115.510 ;
        RECT 100.305 115.465 100.595 115.510 ;
        RECT 103.050 115.450 103.370 115.710 ;
        RECT 103.510 115.650 103.830 115.710 ;
        RECT 103.510 115.510 113.860 115.650 ;
        RECT 103.510 115.450 103.830 115.510 ;
        RECT 42.445 115.310 42.735 115.355 ;
        RECT 45.565 115.310 45.855 115.355 ;
        RECT 47.455 115.310 47.745 115.355 ;
        RECT 42.445 115.170 47.745 115.310 ;
        RECT 42.445 115.125 42.735 115.170 ;
        RECT 45.565 115.125 45.855 115.170 ;
        RECT 47.455 115.125 47.745 115.170 ;
        RECT 69.585 115.310 69.875 115.355 ;
        RECT 72.705 115.310 72.995 115.355 ;
        RECT 74.595 115.310 74.885 115.355 ;
        RECT 69.585 115.170 74.885 115.310 ;
        RECT 69.585 115.125 69.875 115.170 ;
        RECT 72.705 115.125 72.995 115.170 ;
        RECT 74.595 115.125 74.885 115.170 ;
        RECT 93.505 115.310 93.795 115.355 ;
        RECT 96.625 115.310 96.915 115.355 ;
        RECT 98.515 115.310 98.805 115.355 ;
        RECT 93.505 115.170 98.805 115.310 ;
        RECT 93.505 115.125 93.795 115.170 ;
        RECT 96.625 115.125 96.915 115.170 ;
        RECT 98.515 115.125 98.805 115.170 ;
        RECT 108.225 115.310 108.515 115.355 ;
        RECT 111.345 115.310 111.635 115.355 ;
        RECT 113.235 115.310 113.525 115.355 ;
        RECT 108.225 115.170 113.525 115.310 ;
        RECT 113.720 115.310 113.860 115.510 ;
        RECT 118.230 115.450 118.550 115.710 ;
        RECT 119.150 115.650 119.470 115.710 ;
        RECT 120.545 115.650 120.835 115.695 ;
        RECT 119.150 115.510 120.835 115.650 ;
        RECT 119.150 115.450 119.470 115.510 ;
        RECT 120.545 115.465 120.835 115.510 ;
        RECT 125.145 115.465 125.435 115.695 ;
        RECT 125.220 115.310 125.360 115.465 ;
        RECT 113.720 115.170 125.360 115.310 ;
        RECT 108.225 115.125 108.515 115.170 ;
        RECT 111.345 115.125 111.635 115.170 ;
        RECT 113.235 115.125 113.525 115.170 ;
        RECT 38.205 114.970 38.495 115.015 ;
        RECT 40.950 114.970 41.270 115.030 ;
        RECT 38.205 114.830 41.270 114.970 ;
        RECT 38.205 114.785 38.495 114.830 ;
        RECT 40.950 114.770 41.270 114.830 ;
        RECT 41.870 114.970 42.190 115.030 ;
        RECT 46.945 114.970 47.235 115.015 ;
        RECT 41.870 114.830 47.235 114.970 ;
        RECT 41.870 114.770 42.190 114.830 ;
        RECT 46.945 114.785 47.235 114.830 ;
        RECT 48.325 114.970 48.615 115.015 ;
        RECT 49.690 114.970 50.010 115.030 ;
        RECT 48.325 114.830 50.010 114.970 ;
        RECT 48.325 114.785 48.615 114.830 ;
        RECT 49.690 114.770 50.010 114.830 ;
        RECT 65.345 114.970 65.635 115.015 ;
        RECT 71.310 114.970 71.630 115.030 ;
        RECT 65.345 114.830 71.630 114.970 ;
        RECT 65.345 114.785 65.635 114.830 ;
        RECT 71.310 114.770 71.630 114.830 ;
        RECT 74.070 114.770 74.390 115.030 ;
        RECT 75.450 114.770 75.770 115.030 ;
        RECT 97.990 114.770 98.310 115.030 ;
        RECT 99.370 114.770 99.690 115.030 ;
        RECT 110.410 114.970 110.730 115.030 ;
        RECT 102.680 114.830 110.730 114.970 ;
        RECT 39.570 114.290 39.890 114.350 ;
        RECT 41.365 114.335 41.655 114.650 ;
        RECT 42.445 114.630 42.735 114.675 ;
        RECT 46.025 114.630 46.315 114.675 ;
        RECT 47.860 114.630 48.150 114.675 ;
        RECT 42.445 114.490 48.150 114.630 ;
        RECT 42.445 114.445 42.735 114.490 ;
        RECT 46.025 114.445 46.315 114.490 ;
        RECT 47.860 114.445 48.150 114.490 ;
        RECT 53.830 114.630 54.150 114.690 ;
        RECT 58.445 114.630 58.735 114.675 ;
        RECT 61.665 114.630 61.955 114.675 ;
        RECT 63.965 114.630 64.255 114.675 ;
        RECT 66.250 114.630 66.570 114.690 ;
        RECT 53.830 114.490 66.570 114.630 ;
        RECT 53.830 114.430 54.150 114.490 ;
        RECT 58.445 114.445 58.735 114.490 ;
        RECT 61.665 114.445 61.955 114.490 ;
        RECT 63.965 114.445 64.255 114.490 ;
        RECT 66.250 114.430 66.570 114.490 ;
        RECT 68.505 114.335 68.795 114.650 ;
        RECT 69.585 114.630 69.875 114.675 ;
        RECT 73.165 114.630 73.455 114.675 ;
        RECT 75.000 114.630 75.290 114.675 ;
        RECT 69.585 114.490 75.290 114.630 ;
        RECT 69.585 114.445 69.875 114.490 ;
        RECT 73.165 114.445 73.455 114.490 ;
        RECT 75.000 114.445 75.290 114.490 ;
        RECT 87.410 114.630 87.730 114.690 ;
        RECT 91.090 114.630 91.410 114.690 ;
        RECT 102.680 114.675 102.820 114.830 ;
        RECT 110.410 114.770 110.730 114.830 ;
        RECT 112.710 114.770 113.030 115.030 ;
        RECT 114.105 114.970 114.395 115.015 ;
        RECT 125.130 114.970 125.450 115.030 ;
        RECT 114.105 114.830 125.450 114.970 ;
        RECT 114.105 114.785 114.395 114.830 ;
        RECT 125.130 114.770 125.450 114.830 ;
        RECT 87.410 114.490 91.410 114.630 ;
        RECT 87.410 114.430 87.730 114.490 ;
        RECT 91.090 114.430 91.410 114.490 ;
        RECT 41.065 114.290 41.655 114.335 ;
        RECT 44.305 114.290 44.955 114.335 ;
        RECT 39.570 114.150 44.955 114.290 ;
        RECT 39.570 114.090 39.890 114.150 ;
        RECT 41.065 114.105 41.355 114.150 ;
        RECT 44.305 114.105 44.955 114.150 ;
        RECT 68.205 114.290 68.795 114.335 ;
        RECT 70.390 114.290 70.710 114.350 ;
        RECT 71.445 114.290 72.095 114.335 ;
        RECT 68.205 114.150 72.095 114.290 ;
        RECT 68.205 114.105 68.495 114.150 ;
        RECT 70.390 114.090 70.710 114.150 ;
        RECT 71.445 114.105 72.095 114.150 ;
        RECT 89.265 114.290 89.555 114.335 ;
        RECT 91.550 114.290 91.870 114.350 ;
        RECT 92.425 114.335 92.715 114.650 ;
        RECT 93.505 114.630 93.795 114.675 ;
        RECT 97.085 114.630 97.375 114.675 ;
        RECT 98.920 114.630 99.210 114.675 ;
        RECT 93.505 114.490 99.210 114.630 ;
        RECT 93.505 114.445 93.795 114.490 ;
        RECT 97.085 114.445 97.375 114.490 ;
        RECT 98.920 114.445 99.210 114.490 ;
        RECT 100.765 114.630 101.055 114.675 ;
        RECT 102.605 114.630 102.895 114.675 ;
        RECT 100.765 114.490 102.895 114.630 ;
        RECT 100.765 114.445 101.055 114.490 ;
        RECT 102.605 114.445 102.895 114.490 ;
        RECT 89.265 114.150 91.870 114.290 ;
        RECT 89.265 114.105 89.555 114.150 ;
        RECT 91.550 114.090 91.870 114.150 ;
        RECT 92.125 114.290 92.715 114.335 ;
        RECT 94.770 114.290 95.090 114.350 ;
        RECT 95.365 114.290 96.015 114.335 ;
        RECT 92.125 114.150 96.015 114.290 ;
        RECT 92.125 114.105 92.415 114.150 ;
        RECT 94.770 114.090 95.090 114.150 ;
        RECT 95.365 114.105 96.015 114.150 ;
        RECT 91.090 113.950 91.410 114.010 ;
        RECT 100.840 113.950 100.980 114.445 ;
        RECT 107.145 114.335 107.435 114.650 ;
        RECT 108.225 114.630 108.515 114.675 ;
        RECT 111.805 114.630 112.095 114.675 ;
        RECT 113.640 114.630 113.930 114.675 ;
        RECT 108.225 114.490 113.930 114.630 ;
        RECT 108.225 114.445 108.515 114.490 ;
        RECT 111.805 114.445 112.095 114.490 ;
        RECT 113.640 114.445 113.930 114.490 ;
        RECT 117.785 114.630 118.075 114.675 ;
        RECT 119.610 114.630 119.930 114.690 ;
        RECT 121.005 114.630 121.295 114.675 ;
        RECT 117.785 114.490 121.295 114.630 ;
        RECT 117.785 114.445 118.075 114.490 ;
        RECT 119.610 114.430 119.930 114.490 ;
        RECT 121.005 114.445 121.295 114.490 ;
        RECT 126.065 114.630 126.355 114.675 ;
        RECT 130.190 114.630 130.510 114.690 ;
        RECT 126.065 114.490 130.510 114.630 ;
        RECT 126.065 114.445 126.355 114.490 ;
        RECT 130.190 114.430 130.510 114.490 ;
        RECT 103.985 114.105 104.275 114.335 ;
        RECT 106.845 114.290 107.435 114.335 ;
        RECT 110.085 114.290 110.735 114.335 ;
        RECT 112.250 114.290 112.570 114.350 ;
        RECT 106.845 114.150 112.570 114.290 ;
        RECT 106.845 114.105 107.135 114.150 ;
        RECT 110.085 114.105 110.735 114.150 ;
        RECT 91.090 113.810 100.980 113.950 ;
        RECT 104.060 113.950 104.200 114.105 ;
        RECT 112.250 114.090 112.570 114.150 ;
        RECT 111.790 113.950 112.110 114.010 ;
        RECT 104.060 113.810 112.110 113.950 ;
        RECT 91.090 113.750 91.410 113.810 ;
        RECT 111.790 113.750 112.110 113.810 ;
        RECT 29.840 113.130 127.820 113.610 ;
        RECT 135.660 106.690 136.800 133.400 ;
        RECT 133.100 106.600 136.850 106.690 ;
        RECT 129.700 105.630 136.850 106.600 ;
        RECT 133.100 105.500 136.850 105.630 ;
        RECT 133.330 76.630 136.060 77.830 ;
        RECT 137.920 77.810 143.450 77.960 ;
        RECT 21.115 74.380 23.065 74.390 ;
        RECT 19.415 73.240 23.065 74.380 ;
        RECT 19.415 73.230 21.125 73.240 ;
        RECT 28.135 73.230 30.305 74.410 ;
        RECT 32.315 74.390 34.265 74.400 ;
        RECT 30.615 73.250 34.265 74.390 ;
        RECT 30.615 73.240 32.325 73.250 ;
        RECT 39.425 73.200 41.595 74.380 ;
        RECT 43.535 74.360 45.485 74.370 ;
        RECT 41.835 73.220 45.485 74.360 ;
        RECT 54.785 74.340 56.735 74.350 ;
        RECT 41.835 73.210 43.545 73.220 ;
        RECT 3.910 73.080 6.100 73.190 ;
        RECT 50.005 73.140 52.175 74.320 ;
        RECT 53.085 73.200 56.735 74.340 ;
        RECT 53.085 73.190 54.795 73.200 ;
        RECT 61.425 73.170 63.595 74.350 ;
        RECT 66.005 74.330 67.955 74.340 ;
        RECT 64.305 73.190 67.955 74.330 ;
        RECT 64.305 73.180 66.015 73.190 ;
        RECT 72.535 73.180 74.705 74.360 ;
        RECT 77.245 74.320 79.195 74.330 ;
        RECT 75.545 73.180 79.195 74.320 ;
        RECT 75.545 73.170 77.255 73.180 ;
        RECT 83.805 73.170 85.975 74.350 ;
        RECT 88.495 74.330 90.445 74.340 ;
        RECT 86.795 73.190 90.445 74.330 ;
        RECT 99.775 74.320 101.725 74.330 ;
        RECT 86.795 73.180 88.505 73.190 ;
        RECT 94.995 73.110 97.165 74.290 ;
        RECT 98.075 73.180 101.725 74.320 ;
        RECT 98.075 73.170 99.785 73.180 ;
        RECT 106.405 73.160 108.575 74.340 ;
        RECT 111.045 74.320 112.995 74.330 ;
        RECT 109.345 73.180 112.995 74.320 ;
        RECT 109.345 73.170 111.055 73.180 ;
        RECT 117.605 73.160 119.775 74.340 ;
        RECT 122.295 74.320 124.245 74.330 ;
        RECT 120.595 73.180 124.245 74.320 ;
        RECT 129.455 73.240 131.625 74.420 ;
        RECT 120.595 73.170 122.305 73.180 ;
        RECT 3.910 72.820 12.240 73.080 ;
        RECT 29.635 72.840 43.235 72.850 ;
        RECT 18.435 72.820 43.235 72.840 ;
        RECT 3.910 72.800 54.455 72.820 ;
        RECT 3.910 72.790 65.705 72.800 ;
        RECT 133.960 72.790 135.640 76.630 ;
        RECT 137.190 76.610 143.450 77.810 ;
        RECT 137.920 75.460 143.450 76.610 ;
        RECT 3.910 72.780 76.925 72.790 ;
        RECT 85.815 72.780 99.415 72.790 ;
        RECT 132.085 72.780 140.600 72.790 ;
        RECT 3.910 71.700 140.600 72.780 ;
        RECT 3.910 71.690 32.035 71.700 ;
        RECT 3.910 71.670 19.135 71.690 ;
        RECT 40.855 71.670 140.600 71.700 ;
        RECT 3.910 71.500 12.240 71.670 ;
        RECT 52.105 71.650 140.600 71.670 ;
        RECT 63.325 71.640 140.600 71.650 ;
        RECT 74.565 71.630 88.165 71.640 ;
        RECT 97.095 71.630 133.215 71.640 ;
        RECT 3.910 71.370 6.100 71.500 ;
        RECT 10.800 71.180 11.950 71.500 ;
        RECT 10.800 69.480 11.915 71.180 ;
        RECT 29.635 71.170 43.285 71.180 ;
        RECT 15.510 71.155 17.040 71.160 ;
        RECT 18.435 71.155 43.285 71.170 ;
        RECT 12.285 71.150 43.285 71.155 ;
        RECT 12.285 71.130 54.505 71.150 ;
        RECT 141.810 71.140 143.230 75.460 ;
        RECT 12.285 71.120 65.755 71.130 ;
        RECT 12.285 71.110 76.975 71.120 ;
        RECT 85.815 71.110 99.465 71.120 ;
        RECT 140.220 71.110 143.240 71.140 ;
        RECT 12.285 70.030 143.240 71.110 ;
        RECT 12.285 70.020 32.085 70.030 ;
        RECT 12.285 70.005 19.375 70.020 ;
        RECT 10.800 13.800 11.950 69.480 ;
        RECT 12.320 15.450 13.470 70.005 ;
        RECT 15.510 68.660 17.040 70.005 ;
        RECT 40.855 70.000 143.240 70.030 ;
        RECT 52.105 69.980 143.240 70.000 ;
        RECT 63.325 69.970 143.240 69.980 ;
        RECT 74.565 69.960 88.215 69.970 ;
        RECT 97.095 69.960 143.240 69.970 ;
        RECT 140.220 69.910 143.240 69.960 ;
        RECT 29.645 69.670 43.315 69.680 ;
        RECT 18.445 69.650 43.315 69.670 ;
        RECT 18.445 69.630 54.535 69.650 ;
        RECT 18.445 69.620 65.785 69.630 ;
        RECT 139.590 69.620 150.610 69.640 ;
        RECT 18.445 69.610 77.005 69.620 ;
        RECT 85.825 69.610 99.495 69.620 ;
        RECT 132.155 69.610 150.610 69.620 ;
        RECT 18.445 69.570 150.610 69.610 ;
        RECT 18.445 68.530 150.740 69.570 ;
        RECT 18.445 68.520 32.115 68.530 ;
        RECT 40.865 68.500 150.740 68.530 ;
        RECT 52.115 68.490 143.320 68.500 ;
        RECT 52.115 68.480 140.670 68.490 ;
        RECT 63.335 68.470 140.670 68.480 ;
        RECT 74.575 68.460 88.245 68.470 ;
        RECT 97.105 68.460 133.295 68.470 ;
        RECT 141.080 68.450 142.300 68.490 ;
        RECT 149.360 68.470 150.740 68.500 ;
        RECT 29.655 68.100 43.325 68.110 ;
        RECT 13.950 68.080 43.325 68.100 ;
        RECT 13.950 68.060 54.545 68.080 ;
        RECT 13.950 68.050 65.795 68.060 ;
        RECT 13.950 68.040 77.015 68.050 ;
        RECT 85.835 68.040 99.505 68.050 ;
        RECT 139.530 68.040 143.320 68.060 ;
        RECT 13.950 66.960 152.870 68.040 ;
        RECT 13.950 66.950 32.125 66.960 ;
        RECT 13.950 18.530 15.100 66.950 ;
        RECT 40.875 66.930 152.870 66.960 ;
        RECT 52.125 66.910 152.870 66.930 ;
        RECT 63.345 66.900 152.870 66.910 ;
        RECT 74.585 66.890 88.255 66.900 ;
        RECT 97.115 66.890 143.320 66.900 ;
        RECT 141.030 66.770 142.490 66.890 ;
        RECT 21.405 65.510 26.555 65.790 ;
        RECT 27.815 65.490 28.965 65.800 ;
        RECT 32.605 65.520 37.755 65.800 ;
        RECT 39.015 65.500 40.165 65.810 ;
        RECT 43.825 65.490 48.975 65.770 ;
        RECT 50.235 65.470 51.385 65.780 ;
        RECT 149.460 65.760 150.600 65.780 ;
        RECT 55.075 65.470 60.225 65.750 ;
        RECT 61.485 65.450 62.635 65.760 ;
        RECT 66.295 65.460 71.445 65.740 ;
        RECT 72.705 65.440 73.855 65.750 ;
        RECT 77.535 65.450 82.685 65.730 ;
        RECT 83.945 65.430 85.095 65.740 ;
        RECT 88.785 65.460 93.935 65.740 ;
        RECT 95.195 65.440 96.345 65.750 ;
        RECT 100.065 65.450 105.215 65.730 ;
        RECT 106.475 65.430 107.625 65.740 ;
        RECT 111.335 65.450 116.485 65.730 ;
        RECT 117.745 65.430 118.895 65.740 ;
        RECT 122.585 65.450 127.735 65.730 ;
        RECT 128.995 65.430 130.145 65.740 ;
        RECT 133.315 65.430 138.455 65.690 ;
        RECT 21.205 65.140 21.435 65.320 ;
        RECT 26.495 65.190 26.725 65.320 ;
        RECT 21.125 55.220 21.485 65.140 ;
        RECT 26.435 55.240 26.805 65.190 ;
        RECT 27.635 65.150 27.865 65.320 ;
        RECT 27.565 55.200 27.935 65.150 ;
        RECT 28.925 65.140 29.155 65.320 ;
        RECT 32.405 65.150 32.635 65.330 ;
        RECT 37.695 65.200 37.925 65.330 ;
        RECT 28.835 55.250 29.255 65.140 ;
        RECT 32.325 55.230 32.685 65.150 ;
        RECT 37.635 55.250 38.005 65.200 ;
        RECT 38.835 65.160 39.065 65.330 ;
        RECT 38.765 55.210 39.135 65.160 ;
        RECT 40.125 65.150 40.355 65.330 ;
        RECT 40.035 55.260 40.455 65.150 ;
        RECT 43.625 65.120 43.855 65.300 ;
        RECT 48.915 65.170 49.145 65.300 ;
        RECT 43.545 55.200 43.905 65.120 ;
        RECT 48.855 55.220 49.225 65.170 ;
        RECT 50.055 65.130 50.285 65.300 ;
        RECT 49.985 55.180 50.355 65.130 ;
        RECT 51.345 65.120 51.575 65.300 ;
        RECT 51.255 55.230 51.675 65.120 ;
        RECT 54.875 65.100 55.105 65.280 ;
        RECT 60.165 65.150 60.395 65.280 ;
        RECT 54.795 55.180 55.155 65.100 ;
        RECT 60.105 55.200 60.475 65.150 ;
        RECT 61.305 65.110 61.535 65.280 ;
        RECT 61.235 55.160 61.605 65.110 ;
        RECT 62.595 65.100 62.825 65.280 ;
        RECT 62.505 55.210 62.925 65.100 ;
        RECT 66.095 65.090 66.325 65.270 ;
        RECT 71.385 65.140 71.615 65.270 ;
        RECT 66.015 55.170 66.375 65.090 ;
        RECT 71.325 55.190 71.695 65.140 ;
        RECT 72.525 65.100 72.755 65.270 ;
        RECT 72.455 55.150 72.825 65.100 ;
        RECT 73.815 65.090 74.045 65.270 ;
        RECT 73.725 55.200 74.145 65.090 ;
        RECT 77.335 65.080 77.565 65.260 ;
        RECT 82.625 65.130 82.855 65.260 ;
        RECT 77.255 55.160 77.615 65.080 ;
        RECT 82.565 55.180 82.935 65.130 ;
        RECT 83.765 65.090 83.995 65.260 ;
        RECT 83.695 55.140 84.065 65.090 ;
        RECT 85.055 65.080 85.285 65.260 ;
        RECT 88.585 65.090 88.815 65.270 ;
        RECT 93.875 65.140 94.105 65.270 ;
        RECT 84.965 55.190 85.385 65.080 ;
        RECT 88.505 55.170 88.865 65.090 ;
        RECT 93.815 55.190 94.185 65.140 ;
        RECT 95.015 65.100 95.245 65.270 ;
        RECT 94.945 55.150 95.315 65.100 ;
        RECT 96.305 65.090 96.535 65.270 ;
        RECT 96.215 55.200 96.635 65.090 ;
        RECT 99.865 65.080 100.095 65.260 ;
        RECT 105.155 65.130 105.385 65.260 ;
        RECT 99.785 55.160 100.145 65.080 ;
        RECT 105.095 55.180 105.465 65.130 ;
        RECT 106.295 65.090 106.525 65.260 ;
        RECT 106.225 55.140 106.595 65.090 ;
        RECT 107.585 65.080 107.815 65.260 ;
        RECT 111.135 65.080 111.365 65.260 ;
        RECT 116.425 65.130 116.655 65.260 ;
        RECT 107.495 55.190 107.915 65.080 ;
        RECT 111.055 55.160 111.415 65.080 ;
        RECT 116.365 55.180 116.735 65.130 ;
        RECT 117.565 65.090 117.795 65.260 ;
        RECT 117.495 55.140 117.865 65.090 ;
        RECT 118.855 65.080 119.085 65.260 ;
        RECT 122.385 65.080 122.615 65.260 ;
        RECT 127.675 65.130 127.905 65.260 ;
        RECT 118.765 55.190 119.185 65.080 ;
        RECT 122.305 55.160 122.665 65.080 ;
        RECT 127.615 55.180 127.985 65.130 ;
        RECT 128.815 65.090 129.045 65.260 ;
        RECT 128.745 55.140 129.115 65.090 ;
        RECT 130.105 65.080 130.335 65.260 ;
        RECT 133.135 65.130 133.365 65.230 ;
        RECT 130.015 55.190 130.435 65.080 ;
        RECT 133.005 55.240 133.405 65.130 ;
        RECT 138.425 65.100 138.655 65.230 ;
        RECT 133.135 55.230 133.365 55.240 ;
        RECT 138.345 55.130 138.725 65.100 ;
        RECT 149.340 64.660 150.720 65.760 ;
        RECT 20.815 54.230 25.555 54.530 ;
        RECT 32.015 54.240 36.755 54.540 ;
        RECT 43.235 54.210 47.975 54.510 ;
        RECT 54.485 54.190 59.225 54.490 ;
        RECT 65.705 54.180 70.445 54.480 ;
        RECT 76.945 54.170 81.685 54.470 ;
        RECT 88.195 54.180 92.935 54.480 ;
        RECT 99.475 54.170 104.215 54.470 ;
        RECT 110.745 54.170 115.485 54.470 ;
        RECT 121.995 54.170 126.735 54.470 ;
        RECT 21.655 52.320 22.115 52.550 ;
        RECT 25.625 52.280 26.255 52.560 ;
        RECT 25.735 52.240 26.195 52.280 ;
        RECT 27.665 52.240 28.125 52.470 ;
        RECT 32.855 52.330 33.315 52.560 ;
        RECT 36.825 52.290 37.455 52.570 ;
        RECT 36.935 52.250 37.395 52.290 ;
        RECT 38.865 52.250 39.325 52.480 ;
        RECT 44.075 52.300 44.535 52.530 ;
        RECT 48.045 52.260 48.675 52.540 ;
        RECT 48.155 52.220 48.615 52.260 ;
        RECT 50.085 52.220 50.545 52.450 ;
        RECT 55.325 52.280 55.785 52.510 ;
        RECT 59.295 52.240 59.925 52.520 ;
        RECT 59.405 52.200 59.865 52.240 ;
        RECT 61.335 52.200 61.795 52.430 ;
        RECT 66.545 52.270 67.005 52.500 ;
        RECT 70.515 52.230 71.145 52.510 ;
        RECT 70.625 52.190 71.085 52.230 ;
        RECT 72.555 52.190 73.015 52.420 ;
        RECT 77.785 52.260 78.245 52.490 ;
        RECT 81.755 52.220 82.385 52.500 ;
        RECT 81.865 52.180 82.325 52.220 ;
        RECT 83.795 52.180 84.255 52.410 ;
        RECT 89.035 52.270 89.495 52.500 ;
        RECT 93.005 52.230 93.635 52.510 ;
        RECT 93.115 52.190 93.575 52.230 ;
        RECT 95.045 52.190 95.505 52.420 ;
        RECT 100.315 52.260 100.775 52.490 ;
        RECT 104.285 52.220 104.915 52.500 ;
        RECT 104.395 52.180 104.855 52.220 ;
        RECT 106.325 52.180 106.785 52.410 ;
        RECT 111.585 52.260 112.045 52.490 ;
        RECT 115.555 52.220 116.185 52.500 ;
        RECT 115.665 52.180 116.125 52.220 ;
        RECT 117.595 52.180 118.055 52.410 ;
        RECT 122.835 52.260 123.295 52.490 ;
        RECT 126.805 52.220 127.435 52.500 ;
        RECT 126.915 52.180 127.375 52.220 ;
        RECT 128.845 52.180 129.305 52.410 ;
        RECT 21.375 52.010 21.605 52.115 ;
        RECT 21.245 50.290 21.615 52.010 ;
        RECT 22.165 51.890 22.395 52.115 ;
        RECT 25.455 51.980 25.685 52.035 ;
        RECT 21.375 50.115 21.605 50.290 ;
        RECT 22.155 50.210 22.525 51.890 ;
        RECT 22.165 50.115 22.395 50.210 ;
        RECT 21.525 49.670 22.245 49.930 ;
        RECT 19.295 46.650 20.065 47.720 ;
        RECT 21.385 47.490 22.105 47.750 ;
        RECT 21.225 47.200 21.455 47.340 ;
        RECT 21.085 46.430 21.475 47.200 ;
        RECT 22.015 47.190 22.245 47.340 ;
        RECT 22.005 46.450 22.375 47.190 ;
        RECT 25.305 47.010 25.735 51.980 ;
        RECT 26.245 51.970 26.475 52.035 ;
        RECT 27.385 51.970 27.615 52.035 ;
        RECT 26.185 46.970 26.585 51.970 ;
        RECT 27.265 46.970 27.665 51.970 ;
        RECT 28.175 51.940 28.405 52.035 ;
        RECT 32.575 52.020 32.805 52.125 ;
        RECT 28.115 46.970 28.545 51.940 ;
        RECT 32.445 50.300 32.815 52.020 ;
        RECT 33.365 51.900 33.595 52.125 ;
        RECT 36.655 51.990 36.885 52.045 ;
        RECT 32.575 50.125 32.805 50.300 ;
        RECT 33.355 50.220 33.725 51.900 ;
        RECT 33.365 50.125 33.595 50.220 ;
        RECT 32.725 49.680 33.445 49.940 ;
        RECT 25.735 46.600 26.195 46.830 ;
        RECT 27.665 46.710 28.125 46.830 ;
        RECT 27.515 46.600 28.125 46.710 ;
        RECT 30.495 46.660 31.265 47.730 ;
        RECT 32.585 47.500 33.305 47.760 ;
        RECT 32.425 47.210 32.655 47.350 ;
        RECT 21.225 46.340 21.455 46.430 ;
        RECT 22.015 46.340 22.245 46.450 ;
        RECT 27.515 46.430 28.095 46.600 ;
        RECT 32.285 46.440 32.675 47.210 ;
        RECT 33.215 47.200 33.445 47.350 ;
        RECT 33.205 46.460 33.575 47.200 ;
        RECT 36.505 47.020 36.935 51.990 ;
        RECT 37.445 51.980 37.675 52.045 ;
        RECT 38.585 51.980 38.815 52.045 ;
        RECT 37.385 46.980 37.785 51.980 ;
        RECT 38.465 46.980 38.865 51.980 ;
        RECT 39.375 51.950 39.605 52.045 ;
        RECT 43.795 51.990 44.025 52.095 ;
        RECT 39.315 46.980 39.745 51.950 ;
        RECT 43.665 50.270 44.035 51.990 ;
        RECT 44.585 51.870 44.815 52.095 ;
        RECT 47.875 51.960 48.105 52.015 ;
        RECT 43.795 50.095 44.025 50.270 ;
        RECT 44.575 50.190 44.945 51.870 ;
        RECT 44.585 50.095 44.815 50.190 ;
        RECT 43.945 49.650 44.665 49.910 ;
        RECT 36.935 46.610 37.395 46.840 ;
        RECT 38.865 46.720 39.325 46.840 ;
        RECT 38.715 46.610 39.325 46.720 ;
        RECT 41.715 46.630 42.485 47.700 ;
        RECT 43.805 47.470 44.525 47.730 ;
        RECT 43.645 47.180 43.875 47.320 ;
        RECT 32.425 46.350 32.655 46.440 ;
        RECT 33.215 46.350 33.445 46.460 ;
        RECT 38.715 46.440 39.295 46.610 ;
        RECT 43.505 46.410 43.895 47.180 ;
        RECT 44.435 47.170 44.665 47.320 ;
        RECT 44.425 46.430 44.795 47.170 ;
        RECT 47.725 46.990 48.155 51.960 ;
        RECT 48.665 51.950 48.895 52.015 ;
        RECT 49.805 51.950 50.035 52.015 ;
        RECT 48.605 46.950 49.005 51.950 ;
        RECT 49.685 46.950 50.085 51.950 ;
        RECT 50.595 51.920 50.825 52.015 ;
        RECT 55.045 51.970 55.275 52.075 ;
        RECT 50.535 46.950 50.965 51.920 ;
        RECT 54.915 50.250 55.285 51.970 ;
        RECT 55.835 51.850 56.065 52.075 ;
        RECT 59.125 51.940 59.355 51.995 ;
        RECT 55.045 50.075 55.275 50.250 ;
        RECT 55.825 50.170 56.195 51.850 ;
        RECT 55.835 50.075 56.065 50.170 ;
        RECT 55.195 49.630 55.915 49.890 ;
        RECT 48.155 46.580 48.615 46.810 ;
        RECT 50.085 46.690 50.545 46.810 ;
        RECT 49.935 46.580 50.545 46.690 ;
        RECT 52.965 46.610 53.735 47.680 ;
        RECT 55.055 47.450 55.775 47.710 ;
        RECT 54.895 47.160 55.125 47.300 ;
        RECT 43.645 46.320 43.875 46.410 ;
        RECT 44.435 46.320 44.665 46.430 ;
        RECT 49.935 46.410 50.515 46.580 ;
        RECT 54.755 46.390 55.145 47.160 ;
        RECT 55.685 47.150 55.915 47.300 ;
        RECT 55.675 46.410 56.045 47.150 ;
        RECT 58.975 46.970 59.405 51.940 ;
        RECT 59.915 51.930 60.145 51.995 ;
        RECT 61.055 51.930 61.285 51.995 ;
        RECT 59.855 46.930 60.255 51.930 ;
        RECT 60.935 46.930 61.335 51.930 ;
        RECT 61.845 51.900 62.075 51.995 ;
        RECT 66.265 51.960 66.495 52.065 ;
        RECT 61.785 46.930 62.215 51.900 ;
        RECT 66.135 50.240 66.505 51.960 ;
        RECT 67.055 51.840 67.285 52.065 ;
        RECT 70.345 51.930 70.575 51.985 ;
        RECT 66.265 50.065 66.495 50.240 ;
        RECT 67.045 50.160 67.415 51.840 ;
        RECT 67.055 50.065 67.285 50.160 ;
        RECT 66.415 49.620 67.135 49.880 ;
        RECT 59.405 46.560 59.865 46.790 ;
        RECT 61.335 46.670 61.795 46.790 ;
        RECT 61.185 46.560 61.795 46.670 ;
        RECT 64.185 46.600 64.955 47.670 ;
        RECT 66.275 47.440 66.995 47.700 ;
        RECT 66.115 47.150 66.345 47.290 ;
        RECT 54.895 46.300 55.125 46.390 ;
        RECT 55.685 46.300 55.915 46.410 ;
        RECT 61.185 46.390 61.765 46.560 ;
        RECT 65.975 46.380 66.365 47.150 ;
        RECT 66.905 47.140 67.135 47.290 ;
        RECT 66.895 46.400 67.265 47.140 ;
        RECT 70.195 46.960 70.625 51.930 ;
        RECT 71.135 51.920 71.365 51.985 ;
        RECT 72.275 51.920 72.505 51.985 ;
        RECT 71.075 46.920 71.475 51.920 ;
        RECT 72.155 46.920 72.555 51.920 ;
        RECT 73.065 51.890 73.295 51.985 ;
        RECT 77.505 51.950 77.735 52.055 ;
        RECT 73.005 46.920 73.435 51.890 ;
        RECT 77.375 50.230 77.745 51.950 ;
        RECT 78.295 51.830 78.525 52.055 ;
        RECT 81.585 51.920 81.815 51.975 ;
        RECT 77.505 50.055 77.735 50.230 ;
        RECT 78.285 50.150 78.655 51.830 ;
        RECT 78.295 50.055 78.525 50.150 ;
        RECT 77.655 49.610 78.375 49.870 ;
        RECT 70.625 46.550 71.085 46.780 ;
        RECT 72.555 46.660 73.015 46.780 ;
        RECT 72.405 46.550 73.015 46.660 ;
        RECT 75.425 46.590 76.195 47.660 ;
        RECT 77.515 47.430 78.235 47.690 ;
        RECT 77.355 47.140 77.585 47.280 ;
        RECT 66.115 46.290 66.345 46.380 ;
        RECT 66.905 46.290 67.135 46.400 ;
        RECT 72.405 46.380 72.985 46.550 ;
        RECT 77.215 46.370 77.605 47.140 ;
        RECT 78.145 47.130 78.375 47.280 ;
        RECT 78.135 46.390 78.505 47.130 ;
        RECT 81.435 46.950 81.865 51.920 ;
        RECT 82.375 51.910 82.605 51.975 ;
        RECT 83.515 51.910 83.745 51.975 ;
        RECT 82.315 46.910 82.715 51.910 ;
        RECT 83.395 46.910 83.795 51.910 ;
        RECT 84.305 51.880 84.535 51.975 ;
        RECT 88.755 51.960 88.985 52.065 ;
        RECT 84.245 46.910 84.675 51.880 ;
        RECT 88.625 50.240 88.995 51.960 ;
        RECT 89.545 51.840 89.775 52.065 ;
        RECT 92.835 51.930 93.065 51.985 ;
        RECT 88.755 50.065 88.985 50.240 ;
        RECT 89.535 50.160 89.905 51.840 ;
        RECT 89.545 50.065 89.775 50.160 ;
        RECT 88.905 49.620 89.625 49.880 ;
        RECT 81.865 46.540 82.325 46.770 ;
        RECT 83.795 46.650 84.255 46.770 ;
        RECT 83.645 46.540 84.255 46.650 ;
        RECT 86.675 46.600 87.445 47.670 ;
        RECT 88.765 47.440 89.485 47.700 ;
        RECT 88.605 47.150 88.835 47.290 ;
        RECT 77.355 46.280 77.585 46.370 ;
        RECT 78.145 46.280 78.375 46.390 ;
        RECT 83.645 46.370 84.225 46.540 ;
        RECT 88.465 46.380 88.855 47.150 ;
        RECT 89.395 47.140 89.625 47.290 ;
        RECT 89.385 46.400 89.755 47.140 ;
        RECT 92.685 46.960 93.115 51.930 ;
        RECT 93.625 51.920 93.855 51.985 ;
        RECT 94.765 51.920 94.995 51.985 ;
        RECT 93.565 46.920 93.965 51.920 ;
        RECT 94.645 46.920 95.045 51.920 ;
        RECT 95.555 51.890 95.785 51.985 ;
        RECT 100.035 51.950 100.265 52.055 ;
        RECT 95.495 46.920 95.925 51.890 ;
        RECT 99.905 50.230 100.275 51.950 ;
        RECT 100.825 51.830 101.055 52.055 ;
        RECT 104.115 51.920 104.345 51.975 ;
        RECT 100.035 50.055 100.265 50.230 ;
        RECT 100.815 50.150 101.185 51.830 ;
        RECT 100.825 50.055 101.055 50.150 ;
        RECT 100.185 49.610 100.905 49.870 ;
        RECT 93.115 46.550 93.575 46.780 ;
        RECT 95.045 46.660 95.505 46.780 ;
        RECT 94.895 46.550 95.505 46.660 ;
        RECT 97.955 46.590 98.725 47.660 ;
        RECT 100.045 47.430 100.765 47.690 ;
        RECT 99.885 47.140 100.115 47.280 ;
        RECT 88.605 46.290 88.835 46.380 ;
        RECT 89.395 46.290 89.625 46.400 ;
        RECT 94.895 46.380 95.475 46.550 ;
        RECT 99.745 46.370 100.135 47.140 ;
        RECT 100.675 47.130 100.905 47.280 ;
        RECT 100.665 46.390 101.035 47.130 ;
        RECT 103.965 46.950 104.395 51.920 ;
        RECT 104.905 51.910 105.135 51.975 ;
        RECT 106.045 51.910 106.275 51.975 ;
        RECT 104.845 46.910 105.245 51.910 ;
        RECT 105.925 46.910 106.325 51.910 ;
        RECT 106.835 51.880 107.065 51.975 ;
        RECT 111.305 51.950 111.535 52.055 ;
        RECT 106.775 46.910 107.205 51.880 ;
        RECT 111.175 50.230 111.545 51.950 ;
        RECT 112.095 51.830 112.325 52.055 ;
        RECT 115.385 51.920 115.615 51.975 ;
        RECT 111.305 50.055 111.535 50.230 ;
        RECT 112.085 50.150 112.455 51.830 ;
        RECT 112.095 50.055 112.325 50.150 ;
        RECT 111.455 49.610 112.175 49.870 ;
        RECT 104.395 46.540 104.855 46.770 ;
        RECT 106.325 46.650 106.785 46.770 ;
        RECT 106.175 46.540 106.785 46.650 ;
        RECT 109.225 46.590 109.995 47.660 ;
        RECT 111.315 47.430 112.035 47.690 ;
        RECT 111.155 47.140 111.385 47.280 ;
        RECT 99.885 46.280 100.115 46.370 ;
        RECT 100.675 46.280 100.905 46.390 ;
        RECT 106.175 46.370 106.755 46.540 ;
        RECT 111.015 46.370 111.405 47.140 ;
        RECT 111.945 47.130 112.175 47.280 ;
        RECT 111.935 46.390 112.305 47.130 ;
        RECT 115.235 46.950 115.665 51.920 ;
        RECT 116.175 51.910 116.405 51.975 ;
        RECT 117.315 51.910 117.545 51.975 ;
        RECT 116.115 46.910 116.515 51.910 ;
        RECT 117.195 46.910 117.595 51.910 ;
        RECT 118.105 51.880 118.335 51.975 ;
        RECT 122.555 51.950 122.785 52.055 ;
        RECT 118.045 46.910 118.475 51.880 ;
        RECT 122.425 50.230 122.795 51.950 ;
        RECT 123.345 51.830 123.575 52.055 ;
        RECT 126.635 51.920 126.865 51.975 ;
        RECT 122.555 50.055 122.785 50.230 ;
        RECT 123.335 50.150 123.705 51.830 ;
        RECT 123.345 50.055 123.575 50.150 ;
        RECT 122.705 49.610 123.425 49.870 ;
        RECT 115.665 46.540 116.125 46.770 ;
        RECT 117.595 46.650 118.055 46.770 ;
        RECT 117.445 46.540 118.055 46.650 ;
        RECT 120.475 46.590 121.245 47.660 ;
        RECT 122.565 47.430 123.285 47.690 ;
        RECT 122.405 47.140 122.635 47.280 ;
        RECT 111.155 46.280 111.385 46.370 ;
        RECT 111.945 46.280 112.175 46.390 ;
        RECT 117.445 46.370 118.025 46.540 ;
        RECT 122.265 46.370 122.655 47.140 ;
        RECT 123.195 47.130 123.425 47.280 ;
        RECT 123.185 46.390 123.555 47.130 ;
        RECT 126.485 46.950 126.915 51.920 ;
        RECT 127.425 51.910 127.655 51.975 ;
        RECT 128.565 51.910 128.795 51.975 ;
        RECT 127.365 46.910 127.765 51.910 ;
        RECT 128.445 46.910 128.845 51.910 ;
        RECT 129.355 51.880 129.585 51.975 ;
        RECT 129.295 46.910 129.725 51.880 ;
        RECT 126.915 46.540 127.375 46.770 ;
        RECT 128.845 46.650 129.305 46.770 ;
        RECT 128.695 46.540 129.305 46.650 ;
        RECT 122.405 46.280 122.635 46.370 ;
        RECT 123.195 46.280 123.425 46.390 ;
        RECT 128.695 46.370 129.275 46.540 ;
        RECT 21.505 45.950 21.965 46.180 ;
        RECT 32.705 45.960 33.165 46.190 ;
        RECT 43.925 45.930 44.385 46.160 ;
        RECT 55.175 45.910 55.635 46.140 ;
        RECT 66.395 45.900 66.855 46.130 ;
        RECT 77.635 45.890 78.095 46.120 ;
        RECT 88.885 45.900 89.345 46.130 ;
        RECT 100.165 45.890 100.625 46.120 ;
        RECT 111.435 45.890 111.895 46.120 ;
        RECT 122.685 45.890 123.145 46.120 ;
        RECT 29.055 45.020 41.225 45.030 ;
        RECT 17.855 45.005 41.225 45.020 ;
        RECT 15.900 45.000 41.225 45.005 ;
        RECT 15.900 44.980 52.445 45.000 ;
        RECT 15.900 44.970 63.695 44.980 ;
        RECT 15.900 44.960 74.915 44.970 ;
        RECT 85.235 44.960 97.405 44.970 ;
        RECT 15.900 43.880 131.205 44.960 ;
        RECT 15.900 43.870 30.025 43.880 ;
        RECT 15.900 43.855 18.690 43.870 ;
        RECT 15.900 41.620 17.050 43.855 ;
        RECT 40.275 43.850 131.205 43.880 ;
        RECT 51.525 43.830 131.205 43.850 ;
        RECT 62.745 43.820 131.205 43.830 ;
        RECT 73.985 43.810 86.155 43.820 ;
        RECT 96.515 43.810 131.205 43.820 ;
        RECT 29.015 43.330 41.185 43.340 ;
        RECT 17.815 43.310 41.185 43.330 ;
        RECT 142.830 43.320 144.150 43.340 ;
        RECT 17.815 43.290 52.405 43.310 ;
        RECT 140.750 43.300 144.150 43.320 ;
        RECT 17.815 43.280 63.655 43.290 ;
        RECT 119.895 43.280 144.150 43.300 ;
        RECT 17.815 43.270 74.875 43.280 ;
        RECT 85.195 43.270 97.365 43.280 ;
        RECT 108.685 43.270 144.150 43.280 ;
        RECT 17.815 42.180 144.150 43.270 ;
        RECT 18.755 42.150 144.150 42.180 ;
        RECT 18.755 42.120 131.165 42.150 ;
        RECT 18.755 42.090 109.655 42.120 ;
        RECT 18.755 42.080 98.445 42.090 ;
        RECT 41.325 42.070 98.445 42.080 ;
        RECT 142.830 42.070 144.150 42.150 ;
        RECT 41.325 42.060 87.205 42.070 ;
        RECT 75.035 42.050 87.205 42.060 ;
        RECT 15.900 41.540 19.685 41.620 ;
        RECT 142.070 41.610 146.210 41.640 ;
        RECT 119.855 41.590 146.210 41.610 ;
        RECT 108.645 41.550 146.210 41.590 ;
        RECT 15.900 41.520 42.165 41.540 ;
        RECT 97.445 41.530 146.210 41.550 ;
        RECT 15.900 41.510 75.875 41.520 ;
        RECT 86.235 41.510 146.210 41.530 ;
        RECT 15.900 40.500 146.210 41.510 ;
        RECT 15.900 40.480 142.320 40.500 ;
        RECT 15.900 40.470 140.920 40.480 ;
        RECT 18.715 40.460 140.920 40.470 ;
        RECT 142.070 40.460 142.250 40.480 ;
        RECT 18.715 40.440 120.815 40.460 ;
        RECT 18.715 40.400 109.615 40.440 ;
        RECT 18.715 40.390 98.405 40.400 ;
        RECT 41.285 40.380 98.405 40.390 ;
        RECT 41.285 40.370 87.165 40.380 ;
        RECT 74.995 40.360 87.165 40.370 ;
        RECT 26.775 39.230 27.235 39.460 ;
        RECT 38.055 39.230 38.515 39.460 ;
        RECT 49.345 39.210 49.805 39.440 ;
        RECT 60.565 39.210 61.025 39.440 ;
        RECT 71.765 39.210 72.225 39.440 ;
        RECT 83.055 39.200 83.515 39.430 ;
        RECT 94.295 39.220 94.755 39.450 ;
        RECT 105.505 39.240 105.965 39.470 ;
        RECT 116.705 39.280 117.165 39.510 ;
        RECT 127.915 39.300 128.375 39.530 ;
        RECT 20.645 38.810 21.225 38.980 ;
        RECT 26.495 38.960 26.725 39.070 ;
        RECT 27.285 38.980 27.515 39.070 ;
        RECT 20.615 38.700 21.225 38.810 ;
        RECT 20.615 38.580 21.075 38.700 ;
        RECT 22.545 38.580 23.005 38.810 ;
        RECT 20.195 33.470 20.625 38.440 ;
        RECT 20.335 33.375 20.565 33.470 ;
        RECT 21.075 33.440 21.475 38.440 ;
        RECT 22.155 33.440 22.555 38.440 ;
        RECT 21.125 33.375 21.355 33.440 ;
        RECT 22.265 33.375 22.495 33.440 ;
        RECT 23.005 33.430 23.435 38.400 ;
        RECT 26.365 38.220 26.735 38.960 ;
        RECT 26.495 38.070 26.725 38.220 ;
        RECT 27.265 38.210 27.655 38.980 ;
        RECT 31.925 38.810 32.505 38.980 ;
        RECT 37.775 38.960 38.005 39.070 ;
        RECT 38.565 38.980 38.795 39.070 ;
        RECT 27.285 38.070 27.515 38.210 ;
        RECT 26.635 37.660 27.355 37.920 ;
        RECT 28.675 37.690 29.445 38.760 ;
        RECT 31.895 38.700 32.505 38.810 ;
        RECT 31.895 38.580 32.355 38.700 ;
        RECT 33.825 38.580 34.285 38.810 ;
        RECT 26.495 35.480 27.215 35.740 ;
        RECT 26.345 35.200 26.575 35.295 ;
        RECT 26.215 33.520 26.585 35.200 ;
        RECT 27.135 35.120 27.365 35.295 ;
        RECT 23.055 33.375 23.285 33.430 ;
        RECT 26.345 33.295 26.575 33.520 ;
        RECT 27.125 33.400 27.495 35.120 ;
        RECT 31.475 33.470 31.905 38.440 ;
        RECT 27.135 33.295 27.365 33.400 ;
        RECT 31.615 33.375 31.845 33.470 ;
        RECT 32.355 33.440 32.755 38.440 ;
        RECT 33.435 33.440 33.835 38.440 ;
        RECT 32.405 33.375 32.635 33.440 ;
        RECT 33.545 33.375 33.775 33.440 ;
        RECT 34.285 33.430 34.715 38.400 ;
        RECT 37.645 38.220 38.015 38.960 ;
        RECT 37.775 38.070 38.005 38.220 ;
        RECT 38.545 38.210 38.935 38.980 ;
        RECT 43.215 38.790 43.795 38.960 ;
        RECT 49.065 38.940 49.295 39.050 ;
        RECT 49.855 38.960 50.085 39.050 ;
        RECT 38.565 38.070 38.795 38.210 ;
        RECT 37.915 37.660 38.635 37.920 ;
        RECT 39.955 37.690 40.725 38.760 ;
        RECT 43.185 38.680 43.795 38.790 ;
        RECT 43.185 38.560 43.645 38.680 ;
        RECT 45.115 38.560 45.575 38.790 ;
        RECT 37.775 35.480 38.495 35.740 ;
        RECT 37.625 35.200 37.855 35.295 ;
        RECT 37.495 33.520 37.865 35.200 ;
        RECT 38.415 35.120 38.645 35.295 ;
        RECT 34.335 33.375 34.565 33.430 ;
        RECT 37.625 33.295 37.855 33.520 ;
        RECT 38.405 33.400 38.775 35.120 ;
        RECT 42.765 33.450 43.195 38.420 ;
        RECT 38.415 33.295 38.645 33.400 ;
        RECT 42.905 33.355 43.135 33.450 ;
        RECT 43.645 33.420 44.045 38.420 ;
        RECT 44.725 33.420 45.125 38.420 ;
        RECT 43.695 33.355 43.925 33.420 ;
        RECT 44.835 33.355 45.065 33.420 ;
        RECT 45.575 33.410 46.005 38.380 ;
        RECT 48.935 38.200 49.305 38.940 ;
        RECT 49.065 38.050 49.295 38.200 ;
        RECT 49.835 38.190 50.225 38.960 ;
        RECT 54.435 38.790 55.015 38.960 ;
        RECT 60.285 38.940 60.515 39.050 ;
        RECT 61.075 38.960 61.305 39.050 ;
        RECT 49.855 38.050 50.085 38.190 ;
        RECT 49.205 37.640 49.925 37.900 ;
        RECT 51.245 37.670 52.015 38.740 ;
        RECT 54.405 38.680 55.015 38.790 ;
        RECT 54.405 38.560 54.865 38.680 ;
        RECT 56.335 38.560 56.795 38.790 ;
        RECT 49.065 35.460 49.785 35.720 ;
        RECT 48.915 35.180 49.145 35.275 ;
        RECT 48.785 33.500 49.155 35.180 ;
        RECT 49.705 35.100 49.935 35.275 ;
        RECT 45.625 33.355 45.855 33.410 ;
        RECT 48.915 33.275 49.145 33.500 ;
        RECT 49.695 33.380 50.065 35.100 ;
        RECT 53.985 33.450 54.415 38.420 ;
        RECT 49.705 33.275 49.935 33.380 ;
        RECT 54.125 33.355 54.355 33.450 ;
        RECT 54.865 33.420 55.265 38.420 ;
        RECT 55.945 33.420 56.345 38.420 ;
        RECT 54.915 33.355 55.145 33.420 ;
        RECT 56.055 33.355 56.285 33.420 ;
        RECT 56.795 33.410 57.225 38.380 ;
        RECT 60.155 38.200 60.525 38.940 ;
        RECT 60.285 38.050 60.515 38.200 ;
        RECT 61.055 38.190 61.445 38.960 ;
        RECT 65.635 38.790 66.215 38.960 ;
        RECT 71.485 38.940 71.715 39.050 ;
        RECT 72.275 38.960 72.505 39.050 ;
        RECT 61.075 38.050 61.305 38.190 ;
        RECT 60.425 37.640 61.145 37.900 ;
        RECT 62.465 37.670 63.235 38.740 ;
        RECT 65.605 38.680 66.215 38.790 ;
        RECT 65.605 38.560 66.065 38.680 ;
        RECT 67.535 38.560 67.995 38.790 ;
        RECT 60.285 35.460 61.005 35.720 ;
        RECT 60.135 35.180 60.365 35.275 ;
        RECT 60.005 33.500 60.375 35.180 ;
        RECT 60.925 35.100 61.155 35.275 ;
        RECT 56.845 33.355 57.075 33.410 ;
        RECT 60.135 33.275 60.365 33.500 ;
        RECT 60.915 33.380 61.285 35.100 ;
        RECT 65.185 33.450 65.615 38.420 ;
        RECT 60.925 33.275 61.155 33.380 ;
        RECT 65.325 33.355 65.555 33.450 ;
        RECT 66.065 33.420 66.465 38.420 ;
        RECT 67.145 33.420 67.545 38.420 ;
        RECT 66.115 33.355 66.345 33.420 ;
        RECT 67.255 33.355 67.485 33.420 ;
        RECT 67.995 33.410 68.425 38.380 ;
        RECT 71.355 38.200 71.725 38.940 ;
        RECT 71.485 38.050 71.715 38.200 ;
        RECT 72.255 38.190 72.645 38.960 ;
        RECT 76.925 38.780 77.505 38.950 ;
        RECT 82.775 38.930 83.005 39.040 ;
        RECT 83.565 38.950 83.795 39.040 ;
        RECT 72.275 38.050 72.505 38.190 ;
        RECT 71.625 37.640 72.345 37.900 ;
        RECT 73.665 37.670 74.435 38.740 ;
        RECT 76.895 38.670 77.505 38.780 ;
        RECT 76.895 38.550 77.355 38.670 ;
        RECT 78.825 38.550 79.285 38.780 ;
        RECT 71.485 35.460 72.205 35.720 ;
        RECT 71.335 35.180 71.565 35.275 ;
        RECT 71.205 33.500 71.575 35.180 ;
        RECT 72.125 35.100 72.355 35.275 ;
        RECT 68.045 33.355 68.275 33.410 ;
        RECT 71.335 33.275 71.565 33.500 ;
        RECT 72.115 33.380 72.485 35.100 ;
        RECT 76.475 33.440 76.905 38.410 ;
        RECT 72.125 33.275 72.355 33.380 ;
        RECT 76.615 33.345 76.845 33.440 ;
        RECT 77.355 33.410 77.755 38.410 ;
        RECT 78.435 33.410 78.835 38.410 ;
        RECT 77.405 33.345 77.635 33.410 ;
        RECT 78.545 33.345 78.775 33.410 ;
        RECT 79.285 33.400 79.715 38.370 ;
        RECT 82.645 38.190 83.015 38.930 ;
        RECT 82.775 38.040 83.005 38.190 ;
        RECT 83.545 38.180 83.935 38.950 ;
        RECT 88.165 38.800 88.745 38.970 ;
        RECT 94.015 38.950 94.245 39.060 ;
        RECT 94.805 38.970 95.035 39.060 ;
        RECT 83.565 38.040 83.795 38.180 ;
        RECT 82.915 37.630 83.635 37.890 ;
        RECT 84.955 37.660 85.725 38.730 ;
        RECT 88.135 38.690 88.745 38.800 ;
        RECT 88.135 38.570 88.595 38.690 ;
        RECT 90.065 38.570 90.525 38.800 ;
        RECT 82.775 35.450 83.495 35.710 ;
        RECT 82.625 35.170 82.855 35.265 ;
        RECT 82.495 33.490 82.865 35.170 ;
        RECT 83.415 35.090 83.645 35.265 ;
        RECT 79.335 33.345 79.565 33.400 ;
        RECT 82.625 33.265 82.855 33.490 ;
        RECT 83.405 33.370 83.775 35.090 ;
        RECT 87.715 33.460 88.145 38.430 ;
        RECT 83.415 33.265 83.645 33.370 ;
        RECT 87.855 33.365 88.085 33.460 ;
        RECT 88.595 33.430 88.995 38.430 ;
        RECT 89.675 33.430 90.075 38.430 ;
        RECT 88.645 33.365 88.875 33.430 ;
        RECT 89.785 33.365 90.015 33.430 ;
        RECT 90.525 33.420 90.955 38.390 ;
        RECT 93.885 38.210 94.255 38.950 ;
        RECT 94.015 38.060 94.245 38.210 ;
        RECT 94.785 38.200 95.175 38.970 ;
        RECT 99.375 38.820 99.955 38.990 ;
        RECT 105.225 38.970 105.455 39.080 ;
        RECT 106.015 38.990 106.245 39.080 ;
        RECT 94.805 38.060 95.035 38.200 ;
        RECT 94.155 37.650 94.875 37.910 ;
        RECT 96.195 37.680 96.965 38.750 ;
        RECT 99.345 38.710 99.955 38.820 ;
        RECT 99.345 38.590 99.805 38.710 ;
        RECT 101.275 38.590 101.735 38.820 ;
        RECT 94.015 35.470 94.735 35.730 ;
        RECT 93.865 35.190 94.095 35.285 ;
        RECT 93.735 33.510 94.105 35.190 ;
        RECT 94.655 35.110 94.885 35.285 ;
        RECT 90.575 33.365 90.805 33.420 ;
        RECT 93.865 33.285 94.095 33.510 ;
        RECT 94.645 33.390 95.015 35.110 ;
        RECT 98.925 33.480 99.355 38.450 ;
        RECT 94.655 33.285 94.885 33.390 ;
        RECT 99.065 33.385 99.295 33.480 ;
        RECT 99.805 33.450 100.205 38.450 ;
        RECT 100.885 33.450 101.285 38.450 ;
        RECT 99.855 33.385 100.085 33.450 ;
        RECT 100.995 33.385 101.225 33.450 ;
        RECT 101.735 33.440 102.165 38.410 ;
        RECT 105.095 38.230 105.465 38.970 ;
        RECT 105.225 38.080 105.455 38.230 ;
        RECT 105.995 38.220 106.385 38.990 ;
        RECT 110.575 38.860 111.155 39.030 ;
        RECT 116.425 39.010 116.655 39.120 ;
        RECT 117.215 39.030 117.445 39.120 ;
        RECT 106.015 38.080 106.245 38.220 ;
        RECT 105.365 37.670 106.085 37.930 ;
        RECT 107.405 37.700 108.175 38.770 ;
        RECT 110.545 38.750 111.155 38.860 ;
        RECT 110.545 38.630 111.005 38.750 ;
        RECT 112.475 38.630 112.935 38.860 ;
        RECT 105.225 35.490 105.945 35.750 ;
        RECT 105.075 35.210 105.305 35.305 ;
        RECT 104.945 33.530 105.315 35.210 ;
        RECT 105.865 35.130 106.095 35.305 ;
        RECT 101.785 33.385 102.015 33.440 ;
        RECT 105.075 33.305 105.305 33.530 ;
        RECT 105.855 33.410 106.225 35.130 ;
        RECT 110.125 33.520 110.555 38.490 ;
        RECT 110.265 33.425 110.495 33.520 ;
        RECT 111.005 33.490 111.405 38.490 ;
        RECT 112.085 33.490 112.485 38.490 ;
        RECT 111.055 33.425 111.285 33.490 ;
        RECT 112.195 33.425 112.425 33.490 ;
        RECT 112.935 33.480 113.365 38.450 ;
        RECT 116.295 38.270 116.665 39.010 ;
        RECT 116.425 38.120 116.655 38.270 ;
        RECT 117.195 38.260 117.585 39.030 ;
        RECT 121.785 38.880 122.365 39.050 ;
        RECT 127.635 39.030 127.865 39.140 ;
        RECT 128.425 39.050 128.655 39.140 ;
        RECT 117.215 38.120 117.445 38.260 ;
        RECT 116.565 37.710 117.285 37.970 ;
        RECT 118.605 37.740 119.375 38.810 ;
        RECT 121.755 38.770 122.365 38.880 ;
        RECT 121.755 38.650 122.215 38.770 ;
        RECT 123.685 38.650 124.145 38.880 ;
        RECT 116.425 35.530 117.145 35.790 ;
        RECT 116.275 35.250 116.505 35.345 ;
        RECT 116.145 33.570 116.515 35.250 ;
        RECT 117.065 35.170 117.295 35.345 ;
        RECT 112.985 33.425 113.215 33.480 ;
        RECT 105.865 33.305 106.095 33.410 ;
        RECT 116.275 33.345 116.505 33.570 ;
        RECT 117.055 33.450 117.425 35.170 ;
        RECT 121.335 33.540 121.765 38.510 ;
        RECT 117.065 33.345 117.295 33.450 ;
        RECT 121.475 33.445 121.705 33.540 ;
        RECT 122.215 33.510 122.615 38.510 ;
        RECT 123.295 33.510 123.695 38.510 ;
        RECT 122.265 33.445 122.495 33.510 ;
        RECT 123.405 33.445 123.635 33.510 ;
        RECT 124.145 33.500 124.575 38.470 ;
        RECT 127.505 38.290 127.875 39.030 ;
        RECT 127.635 38.140 127.865 38.290 ;
        RECT 128.405 38.280 128.795 39.050 ;
        RECT 128.425 38.140 128.655 38.280 ;
        RECT 127.775 37.730 128.495 37.990 ;
        RECT 129.815 37.760 130.585 38.830 ;
        RECT 142.850 37.630 144.170 38.900 ;
        RECT 127.635 35.550 128.355 35.810 ;
        RECT 127.485 35.270 127.715 35.365 ;
        RECT 127.355 33.590 127.725 35.270 ;
        RECT 128.275 35.190 128.505 35.365 ;
        RECT 124.195 33.445 124.425 33.500 ;
        RECT 127.485 33.365 127.715 33.590 ;
        RECT 128.265 33.470 128.635 35.190 ;
        RECT 128.275 33.365 128.505 33.470 ;
        RECT 20.615 32.940 21.075 33.170 ;
        RECT 22.545 33.130 23.005 33.170 ;
        RECT 22.485 32.850 23.115 33.130 ;
        RECT 26.625 32.860 27.085 33.090 ;
        RECT 31.895 32.940 32.355 33.170 ;
        RECT 33.825 33.130 34.285 33.170 ;
        RECT 33.765 32.850 34.395 33.130 ;
        RECT 37.905 32.860 38.365 33.090 ;
        RECT 43.185 32.920 43.645 33.150 ;
        RECT 45.115 33.110 45.575 33.150 ;
        RECT 45.055 32.830 45.685 33.110 ;
        RECT 49.195 32.840 49.655 33.070 ;
        RECT 54.405 32.920 54.865 33.150 ;
        RECT 56.335 33.110 56.795 33.150 ;
        RECT 56.275 32.830 56.905 33.110 ;
        RECT 60.415 32.840 60.875 33.070 ;
        RECT 65.605 32.920 66.065 33.150 ;
        RECT 67.535 33.110 67.995 33.150 ;
        RECT 67.475 32.830 68.105 33.110 ;
        RECT 71.615 32.840 72.075 33.070 ;
        RECT 76.895 32.910 77.355 33.140 ;
        RECT 78.825 33.100 79.285 33.140 ;
        RECT 78.765 32.820 79.395 33.100 ;
        RECT 82.905 32.830 83.365 33.060 ;
        RECT 88.135 32.930 88.595 33.160 ;
        RECT 90.065 33.120 90.525 33.160 ;
        RECT 90.005 32.840 90.635 33.120 ;
        RECT 94.145 32.850 94.605 33.080 ;
        RECT 99.345 32.950 99.805 33.180 ;
        RECT 101.275 33.140 101.735 33.180 ;
        RECT 101.215 32.860 101.845 33.140 ;
        RECT 105.355 32.870 105.815 33.100 ;
        RECT 110.545 32.990 111.005 33.220 ;
        RECT 112.475 33.180 112.935 33.220 ;
        RECT 112.415 32.900 113.045 33.180 ;
        RECT 116.555 32.910 117.015 33.140 ;
        RECT 121.755 33.010 122.215 33.240 ;
        RECT 123.685 33.200 124.145 33.240 ;
        RECT 123.625 32.920 124.255 33.200 ;
        RECT 127.765 32.930 128.225 33.160 ;
        RECT 23.185 30.880 27.925 31.180 ;
        RECT 34.465 30.880 39.205 31.180 ;
        RECT 45.755 30.860 50.495 31.160 ;
        RECT 56.975 30.860 61.715 31.160 ;
        RECT 68.175 30.860 72.915 31.160 ;
        RECT 79.465 30.850 84.205 31.150 ;
        RECT 90.705 30.870 95.445 31.170 ;
        RECT 101.915 30.890 106.655 31.190 ;
        RECT 113.115 30.930 117.855 31.230 ;
        RECT 124.325 30.950 129.065 31.250 ;
        RECT 19.485 20.270 19.905 30.160 ;
        RECT 19.585 20.090 19.815 20.270 ;
        RECT 20.805 20.260 21.175 30.210 ;
        RECT 20.875 20.090 21.105 20.260 ;
        RECT 21.935 20.220 22.305 30.170 ;
        RECT 27.255 20.270 27.615 30.190 ;
        RECT 30.765 20.270 31.185 30.160 ;
        RECT 22.015 20.090 22.245 20.220 ;
        RECT 27.305 20.090 27.535 20.270 ;
        RECT 30.865 20.090 31.095 20.270 ;
        RECT 32.085 20.260 32.455 30.210 ;
        RECT 32.155 20.090 32.385 20.260 ;
        RECT 33.215 20.220 33.585 30.170 ;
        RECT 38.535 20.270 38.895 30.190 ;
        RECT 33.295 20.090 33.525 20.220 ;
        RECT 38.585 20.090 38.815 20.270 ;
        RECT 42.055 20.250 42.475 30.140 ;
        RECT 42.155 20.070 42.385 20.250 ;
        RECT 43.375 20.240 43.745 30.190 ;
        RECT 43.445 20.070 43.675 20.240 ;
        RECT 44.505 20.200 44.875 30.150 ;
        RECT 49.825 20.250 50.185 30.170 ;
        RECT 53.275 20.250 53.695 30.140 ;
        RECT 44.585 20.070 44.815 20.200 ;
        RECT 49.875 20.070 50.105 20.250 ;
        RECT 53.375 20.070 53.605 20.250 ;
        RECT 54.595 20.240 54.965 30.190 ;
        RECT 54.665 20.070 54.895 20.240 ;
        RECT 55.725 20.200 56.095 30.150 ;
        RECT 61.045 20.250 61.405 30.170 ;
        RECT 64.475 20.250 64.895 30.140 ;
        RECT 55.805 20.070 56.035 20.200 ;
        RECT 61.095 20.070 61.325 20.250 ;
        RECT 64.575 20.070 64.805 20.250 ;
        RECT 65.795 20.240 66.165 30.190 ;
        RECT 65.865 20.070 66.095 20.240 ;
        RECT 66.925 20.200 67.295 30.150 ;
        RECT 72.245 20.250 72.605 30.170 ;
        RECT 67.005 20.070 67.235 20.200 ;
        RECT 72.295 20.070 72.525 20.250 ;
        RECT 75.765 20.240 76.185 30.130 ;
        RECT 75.865 20.060 76.095 20.240 ;
        RECT 77.085 20.230 77.455 30.180 ;
        RECT 77.155 20.060 77.385 20.230 ;
        RECT 78.215 20.190 78.585 30.140 ;
        RECT 83.535 20.240 83.895 30.160 ;
        RECT 87.005 20.260 87.425 30.150 ;
        RECT 78.295 20.060 78.525 20.190 ;
        RECT 83.585 20.060 83.815 20.240 ;
        RECT 87.105 20.080 87.335 20.260 ;
        RECT 88.325 20.250 88.695 30.200 ;
        RECT 88.395 20.080 88.625 20.250 ;
        RECT 89.455 20.210 89.825 30.160 ;
        RECT 94.775 20.260 95.135 30.180 ;
        RECT 98.215 20.280 98.635 30.170 ;
        RECT 89.535 20.080 89.765 20.210 ;
        RECT 94.825 20.080 95.055 20.260 ;
        RECT 98.315 20.100 98.545 20.280 ;
        RECT 99.535 20.270 99.905 30.220 ;
        RECT 99.605 20.100 99.835 20.270 ;
        RECT 100.665 20.230 101.035 30.180 ;
        RECT 105.985 20.280 106.345 30.200 ;
        RECT 109.415 20.320 109.835 30.210 ;
        RECT 100.745 20.100 100.975 20.230 ;
        RECT 106.035 20.100 106.265 20.280 ;
        RECT 109.515 20.140 109.745 20.320 ;
        RECT 110.735 20.310 111.105 30.260 ;
        RECT 110.805 20.140 111.035 20.310 ;
        RECT 111.865 20.270 112.235 30.220 ;
        RECT 117.185 20.320 117.545 30.240 ;
        RECT 120.625 20.340 121.045 30.230 ;
        RECT 111.945 20.140 112.175 20.270 ;
        RECT 117.235 20.140 117.465 20.320 ;
        RECT 120.725 20.160 120.955 20.340 ;
        RECT 121.945 20.330 122.315 30.280 ;
        RECT 122.015 20.160 122.245 20.330 ;
        RECT 123.075 20.290 123.445 30.240 ;
        RECT 128.395 20.340 128.755 30.260 ;
        RECT 123.155 20.160 123.385 20.290 ;
        RECT 128.445 20.160 128.675 20.340 ;
        RECT 132.345 20.170 132.755 30.180 ;
        RECT 137.735 30.120 137.965 30.130 ;
        RECT 132.445 20.130 132.675 20.170 ;
        RECT 137.665 20.080 138.055 30.120 ;
        RECT 19.775 19.610 20.925 19.920 ;
        RECT 22.185 19.620 27.335 19.900 ;
        RECT 31.055 19.610 32.205 19.920 ;
        RECT 33.465 19.620 38.615 19.900 ;
        RECT 42.345 19.590 43.495 19.900 ;
        RECT 44.755 19.600 49.905 19.880 ;
        RECT 53.565 19.590 54.715 19.900 ;
        RECT 55.975 19.600 61.125 19.880 ;
        RECT 64.765 19.590 65.915 19.900 ;
        RECT 67.175 19.600 72.325 19.880 ;
        RECT 76.055 19.580 77.205 19.890 ;
        RECT 78.465 19.590 83.615 19.870 ;
        RECT 87.295 19.600 88.445 19.910 ;
        RECT 89.705 19.610 94.855 19.890 ;
        RECT 98.505 19.620 99.655 19.930 ;
        RECT 100.915 19.630 106.065 19.910 ;
        RECT 109.705 19.660 110.855 19.970 ;
        RECT 112.115 19.670 117.265 19.950 ;
        RECT 120.915 19.680 122.065 19.990 ;
        RECT 123.325 19.690 128.475 19.970 ;
        RECT 132.635 19.640 138.025 19.930 ;
        RECT 142.940 19.110 144.080 37.630 ;
        RECT 13.940 18.460 17.635 18.530 ;
        RECT 117.755 18.510 131.425 18.530 ;
        RECT 106.545 18.470 131.425 18.510 ;
        RECT 13.940 18.440 41.565 18.460 ;
        RECT 95.345 18.450 131.425 18.470 ;
        RECT 13.940 18.430 75.275 18.440 ;
        RECT 84.135 18.430 131.425 18.450 ;
        RECT 13.940 17.380 131.425 18.430 ;
        RECT 142.890 17.990 144.140 19.110 ;
        RECT 145.070 18.880 146.210 40.500 ;
        RECT 145.030 17.960 146.250 18.880 ;
        RECT 13.950 17.370 15.100 17.380 ;
        RECT 16.615 17.360 120.215 17.380 ;
        RECT 16.615 17.320 109.015 17.360 ;
        RECT 16.615 17.310 97.805 17.320 ;
        RECT 39.185 17.300 97.805 17.310 ;
        RECT 39.185 17.290 86.565 17.300 ;
        RECT 72.895 17.280 86.565 17.290 ;
        RECT 117.765 16.950 140.620 16.960 ;
        RECT 142.040 16.950 148.010 16.980 ;
        RECT 117.765 16.940 148.010 16.950 ;
        RECT 106.555 16.900 148.010 16.940 ;
        RECT 16.625 16.870 41.575 16.890 ;
        RECT 95.355 16.880 148.010 16.900 ;
        RECT 16.625 16.860 75.285 16.870 ;
        RECT 84.145 16.860 148.010 16.880 ;
        RECT 16.625 15.840 148.010 16.860 ;
        RECT 16.625 15.820 142.660 15.840 ;
        RECT 16.625 15.810 140.620 15.820 ;
        RECT 142.040 15.810 142.660 15.820 ;
        RECT 16.625 15.790 120.225 15.810 ;
        RECT 16.625 15.750 109.025 15.790 ;
        RECT 16.625 15.740 97.815 15.750 ;
        RECT 39.195 15.730 97.815 15.740 ;
        RECT 39.195 15.720 86.575 15.730 ;
        RECT 72.905 15.710 86.575 15.720 ;
        RECT 131.215 15.460 132.585 15.470 ;
        RECT 12.290 15.390 17.625 15.450 ;
        RECT 117.795 15.440 132.785 15.460 ;
        RECT 106.585 15.400 132.785 15.440 ;
        RECT 12.290 15.370 41.585 15.390 ;
        RECT 95.385 15.380 132.785 15.400 ;
        RECT 12.290 15.360 75.295 15.370 ;
        RECT 84.175 15.360 132.785 15.380 ;
        RECT 12.290 14.320 132.785 15.360 ;
        RECT 142.905 15.040 144.045 15.050 ;
        RECT 12.290 14.310 131.445 14.320 ;
        RECT 12.290 14.300 120.235 14.310 ;
        RECT 12.320 14.280 13.470 14.300 ;
        RECT 16.655 14.290 120.235 14.300 ;
        RECT 16.655 14.250 109.035 14.290 ;
        RECT 16.655 14.240 97.825 14.250 ;
        RECT 39.225 14.230 97.825 14.240 ;
        RECT 39.225 14.220 86.585 14.230 ;
        RECT 72.935 14.210 86.585 14.220 ;
        RECT 142.850 13.920 144.100 15.040 ;
        RECT 145.020 14.870 146.160 14.980 ;
        RECT 144.980 13.950 146.200 14.870 ;
        RECT 16.965 13.800 17.435 13.810 ;
        RECT 10.800 13.780 17.435 13.800 ;
        RECT 10.800 13.720 17.555 13.780 ;
        RECT 117.845 13.770 131.445 13.790 ;
        RECT 106.635 13.730 131.445 13.770 ;
        RECT 10.800 13.700 41.585 13.720 ;
        RECT 95.435 13.710 131.445 13.730 ;
        RECT 10.800 13.690 75.295 13.700 ;
        RECT 84.225 13.690 131.445 13.710 ;
        RECT 10.800 12.650 131.445 13.690 ;
        RECT 16.705 12.640 131.445 12.650 ;
        RECT 16.705 12.620 120.235 12.640 ;
        RECT 16.705 12.580 109.035 12.620 ;
        RECT 16.705 12.570 97.825 12.580 ;
        RECT 39.275 12.560 97.825 12.570 ;
        RECT 39.275 12.550 86.585 12.560 ;
        RECT 72.985 12.540 86.585 12.550 ;
        RECT 128.755 12.240 130.465 12.250 ;
        RECT 117.545 12.220 119.255 12.230 ;
        RECT 106.345 12.180 108.055 12.190 ;
        RECT 27.615 12.170 29.325 12.180 ;
        RECT 38.895 12.170 40.605 12.180 ;
        RECT 25.675 11.030 29.325 12.170 ;
        RECT 36.955 11.030 40.605 12.170 ;
        RECT 95.135 12.160 96.845 12.170 ;
        RECT 50.185 12.150 51.895 12.160 ;
        RECT 61.405 12.150 63.115 12.160 ;
        RECT 72.605 12.150 74.315 12.160 ;
        RECT 25.675 11.020 27.625 11.030 ;
        RECT 36.955 11.020 38.905 11.030 ;
        RECT 48.245 11.010 51.895 12.150 ;
        RECT 59.465 11.010 63.115 12.150 ;
        RECT 70.665 11.010 74.315 12.150 ;
        RECT 83.895 12.140 85.605 12.150 ;
        RECT 48.245 11.000 50.195 11.010 ;
        RECT 59.465 11.000 61.415 11.010 ;
        RECT 70.665 11.000 72.615 11.010 ;
        RECT 81.955 11.000 85.605 12.140 ;
        RECT 93.195 11.020 96.845 12.160 ;
        RECT 104.405 11.040 108.055 12.180 ;
        RECT 115.605 11.080 119.255 12.220 ;
        RECT 126.815 11.100 130.465 12.240 ;
        RECT 126.815 11.090 128.765 11.100 ;
        RECT 115.605 11.070 117.555 11.080 ;
        RECT 104.405 11.030 106.355 11.040 ;
        RECT 93.195 11.010 95.145 11.020 ;
        RECT 81.955 10.990 83.905 11.000 ;
        RECT 142.905 8.580 144.045 13.920 ;
        RECT 74.420 7.440 144.045 8.580 ;
        RECT 74.420 1.410 75.560 7.440 ;
        RECT 145.020 6.630 146.160 13.950 ;
        RECT 93.650 5.490 146.160 6.630 ;
        RECT 93.650 1.480 94.790 5.490 ;
        RECT 146.870 4.560 148.010 15.840 ;
        RECT 113.130 3.420 148.010 4.560 ;
        RECT 113.130 1.610 114.270 3.420 ;
        RECT 149.460 2.770 150.600 64.660 ;
        RECT 131.940 1.880 150.600 2.770 ;
        RECT 131.800 1.630 150.600 1.880 ;
        RECT 74.290 0.160 75.680 1.410 ;
        RECT 93.500 0.230 94.890 1.480 ;
        RECT 112.900 0.360 114.290 1.610 ;
        RECT 131.800 1.380 133.490 1.630 ;
        RECT 151.730 1.420 152.870 66.900 ;
        RECT 131.800 0.430 133.540 1.380 ;
        RECT 113.130 0.330 114.270 0.360 ;
        RECT 151.600 0.300 152.970 1.420 ;
        RECT 93.650 0.150 94.790 0.230 ;
      LAYER met2 ;
        RECT 135.390 223.830 136.740 225.230 ;
        RECT 138.180 223.760 139.530 225.160 ;
        RECT 143.230 223.790 144.580 225.190 ;
        RECT 46.880 211.105 48.760 211.475 ;
        RECT 76.880 211.105 78.760 211.475 ;
        RECT 106.880 211.105 108.760 211.475 ;
        RECT 31.880 208.385 33.760 208.755 ;
        RECT 61.880 208.385 63.760 208.755 ;
        RECT 91.880 208.385 93.760 208.755 ;
        RECT 121.880 208.385 123.760 208.755 ;
        RECT 68.580 207.900 68.840 208.220 ;
        RECT 83.760 208.130 84.020 208.220 ;
        RECT 83.760 207.990 84.880 208.130 ;
        RECT 83.760 207.900 84.020 207.990 ;
        RECT 68.120 206.880 68.380 207.200 ;
        RECT 46.880 205.665 48.760 206.035 ;
        RECT 68.180 205.500 68.320 206.880 ;
        RECT 68.120 205.180 68.380 205.500 ;
        RECT 68.640 205.160 68.780 207.900 ;
        RECT 82.840 207.560 83.100 207.880 ;
        RECT 71.340 207.220 71.600 207.540 ;
        RECT 80.080 207.220 80.340 207.540 ;
        RECT 81.460 207.220 81.720 207.540 ;
        RECT 68.580 204.840 68.840 205.160 ;
        RECT 31.880 202.945 33.760 203.315 ;
        RECT 61.880 202.945 63.760 203.315 ;
        RECT 68.640 201.760 68.780 204.840 ;
        RECT 69.040 204.500 69.300 204.820 ;
        RECT 69.100 202.780 69.240 204.500 ;
        RECT 71.400 202.780 71.540 207.220 ;
        RECT 75.480 206.880 75.740 207.200 ;
        RECT 76.860 207.110 77.120 207.200 ;
        RECT 76.000 206.970 77.120 207.110 ;
        RECT 75.540 204.480 75.680 206.880 ;
        RECT 72.260 204.160 72.520 204.480 ;
        RECT 75.480 204.160 75.740 204.480 ;
        RECT 69.040 202.460 69.300 202.780 ;
        RECT 71.340 202.460 71.600 202.780 ;
        RECT 71.400 201.760 71.540 202.460 ;
        RECT 68.580 201.440 68.840 201.760 ;
        RECT 71.340 201.440 71.600 201.760 ;
        RECT 46.880 200.225 48.760 200.595 ;
        RECT 66.740 199.060 67.000 199.380 ;
        RECT 46.500 198.720 46.760 199.040 ;
        RECT 53.400 198.720 53.660 199.040 ;
        RECT 31.880 197.505 33.760 197.875 ;
        RECT 46.040 195.320 46.300 195.640 ;
        RECT 46.100 194.280 46.240 195.320 ;
        RECT 46.040 193.960 46.300 194.280 ;
        RECT 35.460 193.620 35.720 193.940 ;
        RECT 31.880 192.065 33.760 192.435 ;
        RECT 35.520 188.500 35.660 193.620 ;
        RECT 43.740 192.600 44.000 192.920 ;
        RECT 46.040 192.830 46.300 192.920 ;
        RECT 46.560 192.830 46.700 198.720 ;
        RECT 50.180 196.000 50.440 196.320 ;
        RECT 52.020 196.000 52.280 196.320 ;
        RECT 49.260 195.320 49.520 195.640 ;
        RECT 46.880 194.785 48.760 195.155 ;
        RECT 46.040 192.690 46.700 192.830 ;
        RECT 46.040 192.600 46.300 192.690 ;
        RECT 37.300 190.560 37.560 190.880 ;
        RECT 35.460 188.180 35.720 188.500 ;
        RECT 31.880 186.625 33.760 186.995 ;
        RECT 35.520 183.060 35.660 188.180 ;
        RECT 37.360 188.160 37.500 190.560 ;
        RECT 43.800 190.540 43.940 192.600 ;
        RECT 38.220 190.220 38.480 190.540 ;
        RECT 43.740 190.220 44.000 190.540 ;
        RECT 38.280 189.180 38.420 190.220 ;
        RECT 45.580 189.880 45.840 190.200 ;
        RECT 38.220 188.860 38.480 189.180 ;
        RECT 36.840 187.840 37.100 188.160 ;
        RECT 37.300 187.840 37.560 188.160 ;
        RECT 36.900 185.440 37.040 187.840 ;
        RECT 36.840 185.120 37.100 185.440 ;
        RECT 35.460 182.740 35.720 183.060 ;
        RECT 31.880 181.185 33.760 181.555 ;
        RECT 35.520 181.020 35.660 182.740 ;
        RECT 36.380 182.060 36.640 182.380 ;
        RECT 35.460 180.700 35.720 181.020 ;
        RECT 35.520 177.620 35.660 180.700 ;
        RECT 36.440 180.000 36.580 182.060 ;
        RECT 37.300 181.720 37.560 182.040 ;
        RECT 35.920 179.680 36.180 180.000 ;
        RECT 36.380 179.680 36.640 180.000 ;
        RECT 35.460 177.300 35.720 177.620 ;
        RECT 31.880 175.745 33.760 176.115 ;
        RECT 35.980 174.900 36.120 179.680 ;
        RECT 37.360 177.960 37.500 181.720 ;
        RECT 37.760 179.680 38.020 180.000 ;
        RECT 37.820 179.320 37.960 179.680 ;
        RECT 38.280 179.660 38.420 188.860 ;
        RECT 45.640 188.840 45.780 189.880 ;
        RECT 45.580 188.520 45.840 188.840 ;
        RECT 45.120 187.900 45.380 188.160 ;
        RECT 45.120 187.840 45.780 187.900 ;
        RECT 45.180 187.760 45.780 187.840 ;
        RECT 39.600 187.160 39.860 187.480 ;
        RECT 39.660 183.740 39.800 187.160 ;
        RECT 40.060 186.140 40.320 186.460 ;
        RECT 39.600 183.420 39.860 183.740 ;
        RECT 38.680 182.740 38.940 183.060 ;
        RECT 38.220 179.340 38.480 179.660 ;
        RECT 37.760 179.000 38.020 179.320 ;
        RECT 37.300 177.640 37.560 177.960 ;
        RECT 38.740 175.580 38.880 182.740 ;
        RECT 40.120 180.535 40.260 186.140 ;
        RECT 40.510 185.605 40.790 185.975 ;
        RECT 40.050 180.165 40.330 180.535 ;
        RECT 40.580 180.000 40.720 185.605 ;
        RECT 41.900 185.460 42.160 185.780 ;
        RECT 45.120 185.460 45.380 185.780 ;
        RECT 40.970 184.925 41.250 185.295 ;
        RECT 41.040 181.020 41.180 184.925 ;
        RECT 41.440 181.720 41.700 182.040 ;
        RECT 40.980 180.700 41.240 181.020 ;
        RECT 40.520 179.680 40.780 180.000 ;
        RECT 39.140 177.640 39.400 177.960 ;
        RECT 38.680 175.260 38.940 175.580 ;
        RECT 35.920 174.580 36.180 174.900 ;
        RECT 38.680 174.240 38.940 174.560 ;
        RECT 35.920 173.900 36.180 174.220 ;
        RECT 35.980 172.860 36.120 173.900 ;
        RECT 38.740 172.860 38.880 174.240 ;
        RECT 39.200 172.860 39.340 177.640 ;
        RECT 39.600 176.960 39.860 177.280 ;
        RECT 39.660 174.900 39.800 176.960 ;
        RECT 41.040 174.900 41.180 180.700 ;
        RECT 41.500 180.000 41.640 181.720 ;
        RECT 41.440 179.680 41.700 180.000 ;
        RECT 41.440 179.000 41.700 179.320 ;
        RECT 39.600 174.580 39.860 174.900 ;
        RECT 40.980 174.580 41.240 174.900 ;
        RECT 35.920 172.540 36.180 172.860 ;
        RECT 38.680 172.540 38.940 172.860 ;
        RECT 39.140 172.540 39.400 172.860 ;
        RECT 35.460 171.860 35.720 172.180 ;
        RECT 31.880 170.305 33.760 170.675 ;
        RECT 35.000 168.460 35.260 168.780 ;
        RECT 35.060 167.420 35.200 168.460 ;
        RECT 35.000 167.100 35.260 167.420 ;
        RECT 35.520 166.740 35.660 171.860 ;
        RECT 39.660 169.460 39.800 174.580 ;
        RECT 40.060 173.560 40.320 173.880 ;
        RECT 40.120 171.840 40.260 173.560 ;
        RECT 40.520 171.860 40.780 172.180 ;
        RECT 40.060 171.520 40.320 171.840 ;
        RECT 40.580 170.140 40.720 171.860 ;
        RECT 40.520 169.820 40.780 170.140 ;
        RECT 39.600 169.140 39.860 169.460 ;
        RECT 38.680 168.800 38.940 169.120 ;
        RECT 39.140 168.800 39.400 169.120 ;
        RECT 37.300 168.120 37.560 168.440 ;
        RECT 35.460 166.420 35.720 166.740 ;
        RECT 31.880 164.865 33.760 165.235 ;
        RECT 34.080 162.680 34.340 163.000 ;
        RECT 31.880 159.425 33.760 159.795 ;
        RECT 34.140 159.260 34.280 162.680 ;
        RECT 35.520 161.300 35.660 166.420 ;
        RECT 37.360 164.360 37.500 168.120 ;
        RECT 38.740 167.420 38.880 168.800 ;
        RECT 38.680 167.100 38.940 167.420 ;
        RECT 39.200 167.080 39.340 168.800 ;
        RECT 39.140 166.760 39.400 167.080 ;
        RECT 37.760 166.420 38.020 166.740 ;
        RECT 37.820 164.700 37.960 166.420 ;
        RECT 37.760 164.380 38.020 164.700 ;
        RECT 37.300 164.040 37.560 164.360 ;
        RECT 39.200 164.020 39.340 166.760 ;
        RECT 39.660 164.020 39.800 169.140 ;
        RECT 39.140 163.700 39.400 164.020 ;
        RECT 39.600 163.700 39.860 164.020 ;
        RECT 36.380 162.680 36.640 163.000 ;
        RECT 40.060 162.680 40.320 163.000 ;
        RECT 36.440 161.640 36.580 162.680 ;
        RECT 36.380 161.320 36.640 161.640 ;
        RECT 40.120 161.300 40.260 162.680 ;
        RECT 35.460 160.980 35.720 161.300 ;
        RECT 40.060 160.980 40.320 161.300 ;
        RECT 35.920 159.960 36.180 160.280 ;
        RECT 39.600 159.960 39.860 160.280 ;
        RECT 34.080 158.940 34.340 159.260 ;
        RECT 35.980 157.900 36.120 159.960 ;
        RECT 39.660 158.580 39.800 159.960 ;
        RECT 39.600 158.260 39.860 158.580 ;
        RECT 35.920 157.580 36.180 157.900 ;
        RECT 31.320 155.540 31.580 155.860 ;
        RECT 36.840 155.540 37.100 155.860 ;
        RECT 31.380 150.420 31.520 155.540 ;
        RECT 34.540 154.520 34.800 154.840 ;
        RECT 31.880 153.985 33.760 154.355 ;
        RECT 34.600 152.460 34.740 154.520 ;
        RECT 34.540 152.140 34.800 152.460 ;
        RECT 35.000 151.800 35.260 152.120 ;
        RECT 35.060 151.100 35.200 151.800 ;
        RECT 36.900 151.100 37.040 155.540 ;
        RECT 38.680 154.520 38.940 154.840 ;
        RECT 38.740 153.140 38.880 154.520 ;
        RECT 38.680 152.820 38.940 153.140 ;
        RECT 35.000 150.780 35.260 151.100 ;
        RECT 36.840 150.780 37.100 151.100 ;
        RECT 35.060 150.500 35.200 150.780 ;
        RECT 31.320 150.100 31.580 150.420 ;
        RECT 34.600 150.360 35.200 150.500 ;
        RECT 31.380 144.980 31.520 150.100 ;
        RECT 34.080 149.760 34.340 150.080 ;
        RECT 31.880 148.545 33.760 148.915 ;
        RECT 32.240 146.700 32.500 147.020 ;
        RECT 32.300 145.660 32.440 146.700 ;
        RECT 32.240 145.340 32.500 145.660 ;
        RECT 31.320 144.660 31.580 144.980 ;
        RECT 34.140 144.640 34.280 149.760 ;
        RECT 34.600 145.660 34.740 150.360 ;
        RECT 38.680 147.040 38.940 147.360 ;
        RECT 35.000 146.360 35.260 146.680 ;
        RECT 35.060 145.660 35.200 146.360 ;
        RECT 38.740 145.660 38.880 147.040 ;
        RECT 34.540 145.340 34.800 145.660 ;
        RECT 35.000 145.340 35.260 145.660 ;
        RECT 38.680 145.340 38.940 145.660 ;
        RECT 34.080 144.320 34.340 144.640 ;
        RECT 31.880 143.105 33.760 143.475 ;
        RECT 32.240 141.260 32.500 141.580 ;
        RECT 32.300 140.220 32.440 141.260 ;
        RECT 32.240 139.900 32.500 140.220 ;
        RECT 34.140 139.200 34.280 144.320 ;
        RECT 35.060 139.540 35.200 145.340 ;
        RECT 37.300 143.980 37.560 144.300 ;
        RECT 37.360 142.260 37.500 143.980 ;
        RECT 41.500 142.940 41.640 179.000 ;
        RECT 41.960 176.600 42.100 185.460 ;
        RECT 42.820 184.780 43.080 185.100 ;
        RECT 42.360 184.440 42.620 184.760 ;
        RECT 42.420 183.740 42.560 184.440 ;
        RECT 42.360 183.420 42.620 183.740 ;
        RECT 42.880 182.040 43.020 184.780 ;
        RECT 43.340 183.740 44.860 183.820 ;
        RECT 43.340 183.680 44.920 183.740 ;
        RECT 42.820 181.720 43.080 182.040 ;
        RECT 43.340 180.340 43.480 183.680 ;
        RECT 44.660 183.420 44.920 183.680 ;
        RECT 45.180 183.140 45.320 185.460 ;
        RECT 45.640 185.100 45.780 187.760 ;
        RECT 45.580 184.780 45.840 185.100 ;
        RECT 43.800 183.000 45.320 183.140 ;
        RECT 43.800 182.720 43.940 183.000 ;
        RECT 43.740 182.400 44.000 182.720 ;
        RECT 44.200 180.360 44.460 180.680 ;
        RECT 42.820 180.020 43.080 180.340 ;
        RECT 43.280 180.020 43.540 180.340 ;
        RECT 42.360 179.000 42.620 179.320 ;
        RECT 41.900 176.280 42.160 176.600 ;
        RECT 41.900 173.560 42.160 173.880 ;
        RECT 41.960 172.520 42.100 173.560 ;
        RECT 41.900 172.200 42.160 172.520 ;
        RECT 41.890 165.885 42.170 166.255 ;
        RECT 41.960 161.300 42.100 165.885 ;
        RECT 41.900 160.980 42.160 161.300 ;
        RECT 41.900 154.520 42.160 154.840 ;
        RECT 41.440 142.620 41.700 142.940 ;
        RECT 35.460 141.940 35.720 142.260 ;
        RECT 37.300 141.940 37.560 142.260 ;
        RECT 35.520 141.240 35.660 141.940 ;
        RECT 35.460 140.920 35.720 141.240 ;
        RECT 35.520 140.220 35.660 140.920 ;
        RECT 35.460 139.900 35.720 140.220 ;
        RECT 35.000 139.220 35.260 139.540 ;
        RECT 34.080 138.880 34.340 139.200 ;
        RECT 31.880 137.665 33.760 138.035 ;
        RECT 34.140 133.760 34.280 138.880 ;
        RECT 35.000 135.480 35.260 135.800 ;
        RECT 35.060 134.780 35.200 135.480 ;
        RECT 35.520 134.780 35.660 139.900 ;
        RECT 37.360 138.860 37.500 141.940 ;
        RECT 39.600 141.600 39.860 141.920 ;
        RECT 39.660 140.220 39.800 141.600 ;
        RECT 39.600 139.900 39.860 140.220 ;
        RECT 37.300 138.540 37.560 138.860 ;
        RECT 37.360 136.480 37.500 138.540 ;
        RECT 37.300 136.160 37.560 136.480 ;
        RECT 35.000 134.460 35.260 134.780 ;
        RECT 35.460 134.460 35.720 134.780 ;
        RECT 34.080 133.440 34.340 133.760 ;
        RECT 35.920 133.440 36.180 133.760 ;
        RECT 34.080 132.760 34.340 133.080 ;
        RECT 35.460 132.760 35.720 133.080 ;
        RECT 31.880 132.225 33.760 132.595 ;
        RECT 34.140 131.040 34.280 132.760 ;
        RECT 35.520 131.720 35.660 132.760 ;
        RECT 35.460 131.400 35.720 131.720 ;
        RECT 35.980 131.380 36.120 133.440 ;
        RECT 35.920 131.060 36.180 131.380 ;
        RECT 34.080 130.720 34.340 131.040 ;
        RECT 37.360 130.700 37.500 136.160 ;
        RECT 41.440 134.120 41.700 134.440 ;
        RECT 39.600 133.780 39.860 134.100 ;
        RECT 37.300 130.380 37.560 130.700 ;
        RECT 36.840 130.040 37.100 130.360 ;
        RECT 31.880 126.785 33.760 127.155 ;
        RECT 36.900 126.620 37.040 130.040 ;
        RECT 37.360 128.320 37.500 130.380 ;
        RECT 38.680 130.040 38.940 130.360 ;
        RECT 38.740 128.660 38.880 130.040 ;
        RECT 39.660 129.340 39.800 133.780 ;
        RECT 40.980 130.720 41.240 131.040 ;
        RECT 41.040 129.340 41.180 130.720 ;
        RECT 39.600 129.020 39.860 129.340 ;
        RECT 40.980 129.020 41.240 129.340 ;
        RECT 41.500 129.000 41.640 134.120 ;
        RECT 41.440 128.680 41.700 129.000 ;
        RECT 38.680 128.340 38.940 128.660 ;
        RECT 40.980 128.340 41.240 128.660 ;
        RECT 37.300 128.000 37.560 128.320 ;
        RECT 36.840 126.300 37.100 126.620 ;
        RECT 35.920 124.940 36.180 125.260 ;
        RECT 37.760 124.940 38.020 125.260 ;
        RECT 30.860 122.560 31.120 122.880 ;
        RECT 30.920 104.340 31.060 122.560 ;
        RECT 31.880 121.345 33.760 121.715 ;
        RECT 31.880 115.905 33.760 116.275 ;
        RECT 35.980 104.340 36.120 124.940 ;
        RECT 36.380 123.240 36.640 123.560 ;
        RECT 36.440 118.460 36.580 123.240 ;
        RECT 37.820 118.460 37.960 124.940 ;
        RECT 41.040 124.920 41.180 128.340 ;
        RECT 40.980 124.600 41.240 124.920 ;
        RECT 38.680 122.560 38.940 122.880 ;
        RECT 38.740 121.180 38.880 122.560 ;
        RECT 38.680 120.860 38.940 121.180 ;
        RECT 41.960 120.160 42.100 154.520 ;
        RECT 42.420 153.140 42.560 179.000 ;
        RECT 42.880 178.300 43.020 180.020 ;
        RECT 42.820 177.980 43.080 178.300 ;
        RECT 43.280 171.860 43.540 172.180 ;
        RECT 42.820 171.180 43.080 171.500 ;
        RECT 42.880 169.120 43.020 171.180 ;
        RECT 43.340 169.460 43.480 171.860 ;
        RECT 43.280 169.140 43.540 169.460 ;
        RECT 42.820 168.800 43.080 169.120 ;
        RECT 42.820 168.120 43.080 168.440 ;
        RECT 42.880 166.060 43.020 168.120 ;
        RECT 43.340 166.740 43.480 169.140 ;
        RECT 44.260 168.860 44.400 180.360 ;
        RECT 45.640 180.340 45.780 184.780 ;
        RECT 45.580 180.020 45.840 180.340 ;
        RECT 46.100 179.660 46.240 192.600 ;
        RECT 49.320 190.880 49.460 195.320 ;
        RECT 49.720 193.280 49.980 193.600 ;
        RECT 49.780 190.880 49.920 193.280 ;
        RECT 50.240 191.900 50.380 196.000 ;
        RECT 50.180 191.580 50.440 191.900 ;
        RECT 49.260 190.560 49.520 190.880 ;
        RECT 49.720 190.560 49.980 190.880 ;
        RECT 46.880 189.345 48.760 189.715 ;
        RECT 49.260 188.520 49.520 188.840 ;
        RECT 46.500 188.180 46.760 188.500 ;
        RECT 46.560 186.120 46.700 188.180 ;
        RECT 47.420 187.840 47.680 188.160 ;
        RECT 46.500 185.800 46.760 186.120 ;
        RECT 47.480 185.780 47.620 187.840 ;
        RECT 49.320 186.460 49.460 188.520 ;
        RECT 49.780 188.500 49.920 190.560 ;
        RECT 50.180 189.880 50.440 190.200 ;
        RECT 50.240 189.180 50.380 189.880 ;
        RECT 52.080 189.180 52.220 196.000 ;
        RECT 52.940 195.320 53.200 195.640 ;
        RECT 53.000 194.280 53.140 195.320 ;
        RECT 52.940 193.960 53.200 194.280 ;
        RECT 53.460 192.920 53.600 198.720 ;
        RECT 55.700 198.040 55.960 198.360 ;
        RECT 59.380 198.040 59.640 198.360 ;
        RECT 65.820 198.040 66.080 198.360 ;
        RECT 55.240 196.340 55.500 196.660 ;
        RECT 53.400 192.600 53.660 192.920 ;
        RECT 50.180 188.860 50.440 189.180 ;
        RECT 52.020 188.860 52.280 189.180 ;
        RECT 49.720 188.180 49.980 188.500 ;
        RECT 50.180 188.180 50.440 188.500 ;
        RECT 49.780 187.480 49.920 188.180 ;
        RECT 49.720 187.160 49.980 187.480 ;
        RECT 49.260 186.140 49.520 186.460 ;
        RECT 47.420 185.460 47.680 185.780 ;
        RECT 48.800 185.295 49.060 185.440 ;
        RECT 48.790 184.925 49.070 185.295 ;
        RECT 46.500 184.440 46.760 184.760 ;
        RECT 46.040 179.340 46.300 179.660 ;
        RECT 46.040 176.620 46.300 176.940 ;
        RECT 45.120 176.280 45.380 176.600 ;
        RECT 45.180 174.560 45.320 176.280 ;
        RECT 45.120 174.240 45.380 174.560 ;
        RECT 44.260 168.720 44.860 168.860 ;
        RECT 45.180 168.780 45.320 174.240 ;
        RECT 43.740 168.120 44.000 168.440 ;
        RECT 43.280 166.420 43.540 166.740 ;
        RECT 42.820 165.740 43.080 166.060 ;
        RECT 42.820 163.020 43.080 163.340 ;
        RECT 42.880 161.980 43.020 163.020 ;
        RECT 42.820 161.660 43.080 161.980 ;
        RECT 42.820 157.920 43.080 158.240 ;
        RECT 42.360 152.820 42.620 153.140 ;
        RECT 42.880 152.800 43.020 157.920 ;
        RECT 43.280 153.500 43.540 153.820 ;
        RECT 42.820 152.480 43.080 152.800 ;
        RECT 42.360 152.140 42.620 152.460 ;
        RECT 42.420 148.380 42.560 152.140 ;
        RECT 42.880 150.080 43.020 152.480 ;
        RECT 42.820 149.760 43.080 150.080 ;
        RECT 42.360 148.060 42.620 148.380 ;
        RECT 42.880 147.700 43.020 149.760 ;
        RECT 42.820 147.380 43.080 147.700 ;
        RECT 42.360 142.280 42.620 142.600 ;
        RECT 42.420 139.540 42.560 142.280 ;
        RECT 42.880 142.260 43.020 147.380 ;
        RECT 42.820 141.940 43.080 142.260 ;
        RECT 42.880 139.540 43.020 141.940 ;
        RECT 42.360 139.220 42.620 139.540 ;
        RECT 42.820 139.220 43.080 139.540 ;
        RECT 43.340 138.940 43.480 153.500 ;
        RECT 43.800 148.040 43.940 168.120 ;
        RECT 44.200 166.420 44.460 166.740 ;
        RECT 44.260 160.620 44.400 166.420 ;
        RECT 44.200 160.300 44.460 160.620 ;
        RECT 44.720 160.140 44.860 168.720 ;
        RECT 45.120 168.460 45.380 168.780 ;
        RECT 45.120 166.420 45.380 166.740 ;
        RECT 45.180 161.300 45.320 166.420 ;
        RECT 45.580 165.400 45.840 165.720 ;
        RECT 45.120 160.980 45.380 161.300 ;
        RECT 44.720 160.000 45.320 160.140 ;
        RECT 44.660 157.240 44.920 157.560 ;
        RECT 44.720 149.820 44.860 157.240 ;
        RECT 45.180 153.140 45.320 160.000 ;
        RECT 45.120 152.820 45.380 153.140 ;
        RECT 45.640 152.800 45.780 165.400 ;
        RECT 46.100 155.520 46.240 176.620 ;
        RECT 46.560 174.900 46.700 184.440 ;
        RECT 46.880 183.905 48.760 184.275 ;
        RECT 49.780 182.720 49.920 187.160 ;
        RECT 49.720 182.400 49.980 182.720 ;
        RECT 50.240 181.950 50.380 188.180 ;
        RECT 52.020 187.500 52.280 187.820 ;
        RECT 52.480 187.500 52.740 187.820 ;
        RECT 50.630 185.605 50.910 185.975 ;
        RECT 48.400 181.810 50.380 181.950 ;
        RECT 48.400 180.680 48.540 181.810 ;
        RECT 48.340 180.360 48.600 180.680 ;
        RECT 49.250 180.165 49.530 180.535 ;
        RECT 49.720 180.360 49.980 180.680 ;
        RECT 46.880 178.465 48.760 178.835 ;
        RECT 48.800 177.980 49.060 178.300 ;
        RECT 48.860 177.620 49.000 177.980 ;
        RECT 49.320 177.620 49.460 180.165 ;
        RECT 49.780 179.855 49.920 180.360 ;
        RECT 49.710 179.485 49.990 179.855 ;
        RECT 50.700 177.960 50.840 185.605 ;
        RECT 52.080 183.400 52.220 187.500 ;
        RECT 52.540 185.100 52.680 187.500 ;
        RECT 52.480 184.780 52.740 185.100 ;
        RECT 52.020 183.080 52.280 183.400 ;
        RECT 51.090 180.165 51.370 180.535 ;
        RECT 53.460 180.340 53.600 192.600 ;
        RECT 54.320 190.900 54.580 191.220 ;
        RECT 54.780 190.900 55.040 191.220 ;
        RECT 54.380 187.820 54.520 190.900 ;
        RECT 54.320 187.500 54.580 187.820 ;
        RECT 54.380 185.440 54.520 187.500 ;
        RECT 54.320 185.120 54.580 185.440 ;
        RECT 54.380 183.060 54.520 185.120 ;
        RECT 54.840 185.100 54.980 190.900 ;
        RECT 55.300 190.880 55.440 196.340 ;
        RECT 55.760 190.880 55.900 198.040 ;
        RECT 56.620 196.000 56.880 196.320 ;
        RECT 58.000 196.000 58.260 196.320 ;
        RECT 56.160 195.320 56.420 195.640 ;
        RECT 56.220 194.280 56.360 195.320 ;
        RECT 56.160 193.960 56.420 194.280 ;
        RECT 56.680 191.900 56.820 196.000 ;
        RECT 56.620 191.580 56.880 191.900 ;
        RECT 55.240 190.560 55.500 190.880 ;
        RECT 55.700 190.560 55.960 190.880 ;
        RECT 57.080 189.880 57.340 190.200 ;
        RECT 57.140 186.460 57.280 189.880 ;
        RECT 57.080 186.140 57.340 186.460 ;
        RECT 55.240 185.120 55.500 185.440 ;
        RECT 56.620 185.120 56.880 185.440 ;
        RECT 54.780 184.780 55.040 185.100 ;
        RECT 54.840 183.740 54.980 184.780 ;
        RECT 54.780 183.420 55.040 183.740 ;
        RECT 54.320 182.740 54.580 183.060 ;
        RECT 55.300 181.020 55.440 185.120 ;
        RECT 56.680 182.460 56.820 185.120 ;
        RECT 58.060 183.060 58.200 196.000 ;
        RECT 59.440 195.980 59.580 198.040 ;
        RECT 61.880 197.505 63.760 197.875 ;
        RECT 60.760 196.340 61.020 196.660 ;
        RECT 59.380 195.660 59.640 195.980 ;
        RECT 58.920 192.600 59.180 192.920 ;
        RECT 58.980 191.900 59.120 192.600 ;
        RECT 58.920 191.580 59.180 191.900 ;
        RECT 59.440 191.560 59.580 195.660 ;
        RECT 60.300 192.600 60.560 192.920 ;
        RECT 59.380 191.240 59.640 191.560 ;
        RECT 59.380 190.560 59.640 190.880 ;
        RECT 59.440 188.160 59.580 190.560 ;
        RECT 59.380 187.840 59.640 188.160 ;
        RECT 59.840 187.840 60.100 188.160 ;
        RECT 58.460 184.440 58.720 184.760 ;
        RECT 58.000 182.740 58.260 183.060 ;
        RECT 56.220 182.380 56.820 182.460 ;
        RECT 57.080 182.400 57.340 182.720 ;
        RECT 56.160 182.320 56.820 182.380 ;
        RECT 56.160 182.060 56.420 182.320 ;
        RECT 55.240 180.700 55.500 181.020 ;
        RECT 56.220 180.680 56.360 182.060 ;
        RECT 57.140 181.020 57.280 182.400 ;
        RECT 57.080 180.700 57.340 181.020 ;
        RECT 56.160 180.360 56.420 180.680 ;
        RECT 57.140 180.420 57.280 180.700 ;
        RECT 51.160 180.000 51.300 180.165 ;
        RECT 53.400 180.020 53.660 180.340 ;
        RECT 56.220 180.000 56.360 180.360 ;
        RECT 57.140 180.280 57.740 180.420 ;
        RECT 57.600 180.000 57.740 180.280 ;
        RECT 51.100 179.680 51.360 180.000 ;
        RECT 52.020 179.680 52.280 180.000 ;
        RECT 56.160 179.680 56.420 180.000 ;
        RECT 57.540 179.680 57.800 180.000 ;
        RECT 50.640 177.640 50.900 177.960 ;
        RECT 48.800 177.300 49.060 177.620 ;
        RECT 49.260 177.300 49.520 177.620 ;
        RECT 50.180 177.300 50.440 177.620 ;
        RECT 50.240 176.600 50.380 177.300 ;
        RECT 50.180 176.280 50.440 176.600 ;
        RECT 46.500 174.580 46.760 174.900 ;
        RECT 50.240 174.220 50.380 176.280 ;
        RECT 50.180 173.900 50.440 174.220 ;
        RECT 46.880 173.025 48.760 173.395 ;
        RECT 51.160 172.940 51.300 179.680 ;
        RECT 52.080 179.320 52.220 179.680 ;
        RECT 52.020 179.000 52.280 179.320 ;
        RECT 53.400 179.000 53.660 179.320 ;
        RECT 54.320 179.000 54.580 179.320 ;
        RECT 52.020 177.640 52.280 177.960 ;
        RECT 52.480 177.640 52.740 177.960 ;
        RECT 51.160 172.800 51.760 172.940 ;
        RECT 49.260 170.840 49.520 171.160 ;
        RECT 49.720 170.840 49.980 171.160 ;
        RECT 47.880 168.975 48.140 169.120 ;
        RECT 47.870 168.605 48.150 168.975 ;
        RECT 46.880 167.585 48.760 167.955 ;
        RECT 49.320 167.080 49.460 170.840 ;
        RECT 49.780 169.120 49.920 170.840 ;
        RECT 49.720 168.800 49.980 169.120 ;
        RECT 51.100 167.100 51.360 167.420 ;
        RECT 49.260 166.760 49.520 167.080 ;
        RECT 48.340 166.420 48.600 166.740 ;
        RECT 50.640 166.420 50.900 166.740 ;
        RECT 46.500 166.080 46.760 166.400 ;
        RECT 46.560 161.890 46.700 166.080 ;
        RECT 48.400 164.700 48.540 166.420 ;
        RECT 49.260 166.080 49.520 166.400 ;
        RECT 50.700 166.255 50.840 166.420 ;
        RECT 48.340 164.380 48.600 164.700 ;
        RECT 49.320 163.000 49.460 166.080 ;
        RECT 50.630 165.885 50.910 166.255 ;
        RECT 50.180 165.400 50.440 165.720 ;
        RECT 49.260 162.680 49.520 163.000 ;
        RECT 46.880 162.145 48.760 162.515 ;
        RECT 46.560 161.750 47.160 161.890 ;
        RECT 47.020 161.300 47.160 161.750 ;
        RECT 49.320 161.640 49.460 162.680 ;
        RECT 46.960 160.980 47.220 161.300 ;
        RECT 48.330 161.125 48.610 161.495 ;
        RECT 49.260 161.320 49.520 161.640 ;
        RECT 50.240 161.300 50.380 165.400 ;
        RECT 50.640 163.700 50.900 164.020 ;
        RECT 50.700 161.980 50.840 163.700 ;
        RECT 51.160 163.340 51.300 167.100 ;
        RECT 51.100 163.020 51.360 163.340 ;
        RECT 50.640 161.660 50.900 161.980 ;
        RECT 48.340 160.980 48.600 161.125 ;
        RECT 50.180 160.980 50.440 161.300 ;
        RECT 47.020 160.280 47.160 160.980 ;
        RECT 48.400 160.620 48.540 160.980 ;
        RECT 48.340 160.300 48.600 160.620 ;
        RECT 46.500 159.960 46.760 160.280 ;
        RECT 46.960 159.960 47.220 160.280 ;
        RECT 50.180 159.960 50.440 160.280 ;
        RECT 46.560 155.860 46.700 159.960 ;
        RECT 46.880 156.705 48.760 157.075 ;
        RECT 46.500 155.540 46.760 155.860 ;
        RECT 46.040 155.200 46.300 155.520 ;
        RECT 49.720 154.520 49.980 154.840 ;
        RECT 46.500 153.500 46.760 153.820 ;
        RECT 49.260 153.500 49.520 153.820 ;
        RECT 45.580 152.480 45.840 152.800 ;
        RECT 45.120 151.800 45.380 152.120 ;
        RECT 45.180 150.420 45.320 151.800 ;
        RECT 45.120 150.100 45.380 150.420 ;
        RECT 44.720 149.680 45.320 149.820 ;
        RECT 43.740 147.720 44.000 148.040 ;
        RECT 42.420 138.800 43.480 138.940 ;
        RECT 42.420 120.840 42.560 138.800 ;
        RECT 43.280 134.460 43.540 134.780 ;
        RECT 43.340 132.060 43.480 134.460 ;
        RECT 44.200 133.440 44.460 133.760 ;
        RECT 43.280 131.740 43.540 132.060 ;
        RECT 42.820 130.380 43.080 130.700 ;
        RECT 42.880 128.320 43.020 130.380 ;
        RECT 44.260 130.360 44.400 133.440 ;
        RECT 44.200 130.040 44.460 130.360 ;
        RECT 42.820 128.000 43.080 128.320 ;
        RECT 42.820 125.620 43.080 125.940 ;
        RECT 42.880 123.900 43.020 125.620 ;
        RECT 44.260 125.600 44.400 130.040 ;
        RECT 44.200 125.280 44.460 125.600 ;
        RECT 42.820 123.580 43.080 123.900 ;
        RECT 45.180 123.560 45.320 149.680 ;
        RECT 46.560 148.380 46.700 153.500 ;
        RECT 46.880 151.265 48.760 151.635 ;
        RECT 49.320 151.100 49.460 153.500 ;
        RECT 49.780 151.100 49.920 154.520 ;
        RECT 50.240 152.800 50.380 159.960 ;
        RECT 51.620 155.860 51.760 172.800 ;
        RECT 52.080 170.140 52.220 177.640 ;
        RECT 52.540 175.580 52.680 177.640 ;
        RECT 52.940 176.280 53.200 176.600 ;
        RECT 52.480 175.260 52.740 175.580 ;
        RECT 52.020 169.820 52.280 170.140 ;
        RECT 53.000 169.540 53.140 176.280 ;
        RECT 52.080 169.400 53.140 169.540 ;
        RECT 52.080 166.740 52.220 169.400 ;
        RECT 52.940 168.800 53.200 169.120 ;
        RECT 52.020 166.420 52.280 166.740 ;
        RECT 53.000 162.855 53.140 168.800 ;
        RECT 52.930 162.485 53.210 162.855 ;
        RECT 53.460 157.900 53.600 179.000 ;
        RECT 53.860 168.975 54.120 169.120 ;
        RECT 53.850 168.605 54.130 168.975 ;
        RECT 53.860 168.120 54.120 168.440 ;
        RECT 53.920 166.740 54.060 168.120 ;
        RECT 53.860 166.420 54.120 166.740 ;
        RECT 53.920 164.020 54.060 166.420 ;
        RECT 53.860 163.700 54.120 164.020 ;
        RECT 53.860 158.940 54.120 159.260 ;
        RECT 53.400 157.580 53.660 157.900 ;
        RECT 53.400 155.880 53.660 156.200 ;
        RECT 51.560 155.540 51.820 155.860 ;
        RECT 51.620 153.820 51.760 155.540 ;
        RECT 50.640 153.500 50.900 153.820 ;
        RECT 51.560 153.500 51.820 153.820 ;
        RECT 50.180 152.480 50.440 152.800 ;
        RECT 50.700 151.860 50.840 153.500 ;
        RECT 51.100 152.480 51.360 152.800 ;
        RECT 50.240 151.720 50.840 151.860 ;
        RECT 49.260 150.780 49.520 151.100 ;
        RECT 49.720 150.780 49.980 151.100 ;
        RECT 50.240 150.500 50.380 151.720 ;
        RECT 51.160 151.180 51.300 152.480 ;
        RECT 52.940 152.140 53.200 152.460 ;
        RECT 48.800 150.100 49.060 150.420 ;
        RECT 49.320 150.360 50.380 150.500 ;
        RECT 50.700 151.040 51.300 151.180 ;
        RECT 53.000 151.100 53.140 152.140 ;
        RECT 50.700 150.420 50.840 151.040 ;
        RECT 52.940 150.780 53.200 151.100 ;
        RECT 46.500 148.060 46.760 148.380 ;
        RECT 45.580 147.380 45.840 147.700 ;
        RECT 45.640 144.640 45.780 147.380 ;
        RECT 48.860 146.680 49.000 150.100 ;
        RECT 48.800 146.360 49.060 146.680 ;
        RECT 46.880 145.825 48.760 146.195 ;
        RECT 45.580 144.320 45.840 144.640 ;
        RECT 45.640 142.260 45.780 144.320 ;
        RECT 45.580 142.170 45.840 142.260 ;
        RECT 45.580 142.030 46.240 142.170 ;
        RECT 45.580 141.940 45.840 142.030 ;
        RECT 46.100 140.220 46.240 142.030 ;
        RECT 46.500 140.920 46.760 141.240 ;
        RECT 46.040 139.900 46.300 140.220 ;
        RECT 46.560 139.880 46.700 140.920 ;
        RECT 46.880 140.385 48.760 140.755 ;
        RECT 46.500 139.560 46.760 139.880 ;
        RECT 48.800 139.220 49.060 139.540 ;
        RECT 48.860 136.820 49.000 139.220 ;
        RECT 48.800 136.500 49.060 136.820 ;
        RECT 46.880 134.945 48.760 135.315 ;
        RECT 46.500 131.740 46.760 132.060 ;
        RECT 46.560 131.380 46.700 131.740 ;
        RECT 46.500 131.060 46.760 131.380 ;
        RECT 45.580 128.000 45.840 128.320 ;
        RECT 45.640 124.920 45.780 128.000 ;
        RECT 46.560 125.600 46.700 131.060 ;
        RECT 46.880 129.505 48.760 129.875 ;
        RECT 46.500 125.280 46.760 125.600 ;
        RECT 45.580 124.600 45.840 124.920 ;
        RECT 46.880 124.065 48.760 124.435 ;
        RECT 45.120 123.240 45.380 123.560 ;
        RECT 44.660 120.860 44.920 121.180 ;
        RECT 42.360 120.520 42.620 120.840 ;
        RECT 41.900 119.840 42.160 120.160 ;
        RECT 40.980 119.500 41.240 119.820 ;
        RECT 41.040 118.460 41.180 119.500 ;
        RECT 41.900 119.160 42.160 119.480 ;
        RECT 36.380 118.140 36.640 118.460 ;
        RECT 37.760 118.140 38.020 118.460 ;
        RECT 40.980 118.140 41.240 118.460 ;
        RECT 39.600 116.440 39.860 116.760 ;
        RECT 39.660 114.380 39.800 116.440 ;
        RECT 41.960 115.060 42.100 119.160 ;
        RECT 44.720 118.120 44.860 120.860 ;
        RECT 46.040 120.180 46.300 120.500 ;
        RECT 44.660 117.800 44.920 118.120 ;
        RECT 40.980 114.740 41.240 115.060 ;
        RECT 41.900 114.740 42.160 115.060 ;
        RECT 39.600 114.060 39.860 114.380 ;
        RECT 41.040 104.340 41.180 114.740 ;
        RECT 46.100 104.340 46.240 120.180 ;
        RECT 49.320 119.480 49.460 150.360 ;
        RECT 50.640 150.100 50.900 150.420 ;
        RECT 51.100 150.100 51.360 150.420 ;
        RECT 50.700 147.360 50.840 150.100 ;
        RECT 51.160 149.400 51.300 150.100 ;
        RECT 51.100 149.080 51.360 149.400 ;
        RECT 50.640 147.040 50.900 147.360 ;
        RECT 51.160 147.020 51.300 149.080 ;
        RECT 53.460 148.380 53.600 155.880 ;
        RECT 53.920 153.480 54.060 158.940 ;
        RECT 53.860 153.160 54.120 153.480 ;
        RECT 53.860 150.780 54.120 151.100 ;
        RECT 53.400 148.060 53.660 148.380 ;
        RECT 51.100 146.700 51.360 147.020 ;
        RECT 49.720 146.360 49.980 146.680 ;
        RECT 49.780 141.240 49.920 146.360 ;
        RECT 50.180 141.260 50.440 141.580 ;
        RECT 53.400 141.260 53.660 141.580 ;
        RECT 49.720 140.920 49.980 141.240 ;
        RECT 49.780 139.200 49.920 140.920 ;
        RECT 49.720 138.880 49.980 139.200 ;
        RECT 50.240 137.500 50.380 141.260 ;
        RECT 51.100 139.560 51.360 139.880 ;
        RECT 50.180 137.180 50.440 137.500 ;
        RECT 50.240 136.820 50.380 137.180 ;
        RECT 51.160 136.820 51.300 139.560 ;
        RECT 53.460 137.160 53.600 141.260 ;
        RECT 53.920 138.940 54.060 150.780 ;
        RECT 54.380 147.700 54.520 179.000 ;
        RECT 57.540 176.620 57.800 176.940 ;
        RECT 57.600 175.580 57.740 176.620 ;
        RECT 57.540 175.260 57.800 175.580 ;
        RECT 57.600 172.860 57.740 175.260 ;
        RECT 58.000 174.580 58.260 174.900 ;
        RECT 58.060 172.860 58.200 174.580 ;
        RECT 57.540 172.540 57.800 172.860 ;
        RECT 58.000 172.540 58.260 172.860 ;
        RECT 57.080 171.520 57.340 171.840 ;
        RECT 54.770 168.605 55.050 168.975 ;
        RECT 54.840 166.400 54.980 168.605 ;
        RECT 55.700 168.295 55.960 168.440 ;
        RECT 55.690 167.925 55.970 168.295 ;
        RECT 57.140 166.400 57.280 171.520 ;
        RECT 57.600 171.500 57.740 172.540 ;
        RECT 57.540 171.180 57.800 171.500 ;
        RECT 57.600 169.120 57.740 171.180 ;
        RECT 58.000 169.140 58.260 169.460 ;
        RECT 57.540 168.800 57.800 169.120 ;
        RECT 54.780 166.310 55.040 166.400 ;
        RECT 54.780 166.170 55.440 166.310 ;
        RECT 54.780 166.080 55.040 166.170 ;
        RECT 54.780 165.400 55.040 165.720 ;
        RECT 54.840 158.580 54.980 165.400 ;
        RECT 55.300 163.000 55.440 166.170 ;
        RECT 57.080 166.080 57.340 166.400 ;
        RECT 58.060 166.060 58.200 169.140 ;
        RECT 57.540 165.740 57.800 166.060 ;
        RECT 58.000 165.740 58.260 166.060 ;
        RECT 55.700 165.400 55.960 165.720 ;
        RECT 56.160 165.400 56.420 165.720 ;
        RECT 55.240 162.680 55.500 163.000 ;
        RECT 55.760 161.300 55.900 165.400 ;
        RECT 56.220 161.640 56.360 165.400 ;
        RECT 57.080 164.610 57.340 164.700 ;
        RECT 57.600 164.610 57.740 165.740 ;
        RECT 57.080 164.470 57.740 164.610 ;
        RECT 57.080 164.380 57.340 164.470 ;
        RECT 57.070 163.165 57.350 163.535 ;
        RECT 57.140 161.980 57.280 163.165 ;
        RECT 57.600 162.910 57.740 164.470 ;
        RECT 58.000 163.535 58.260 163.680 ;
        RECT 57.990 163.165 58.270 163.535 ;
        RECT 57.600 162.770 58.200 162.910 ;
        RECT 57.080 161.660 57.340 161.980 ;
        RECT 56.160 161.320 56.420 161.640 ;
        RECT 55.700 160.980 55.960 161.300 ;
        RECT 57.530 161.125 57.810 161.495 ;
        RECT 58.060 161.330 58.200 162.770 ;
        RECT 58.520 162.175 58.660 184.440 ;
        RECT 59.900 183.740 60.040 187.840 ;
        RECT 59.840 183.420 60.100 183.740 ;
        RECT 60.360 183.060 60.500 192.600 ;
        RECT 60.820 191.220 60.960 196.340 ;
        RECT 63.980 196.000 64.240 196.320 ;
        RECT 61.220 195.320 61.480 195.640 ;
        RECT 61.280 194.280 61.420 195.320 ;
        RECT 61.220 193.960 61.480 194.280 ;
        RECT 61.220 193.280 61.480 193.600 ;
        RECT 60.760 190.900 61.020 191.220 ;
        RECT 61.280 188.500 61.420 193.280 ;
        RECT 61.880 192.065 63.760 192.435 ;
        RECT 64.040 191.900 64.180 196.000 ;
        RECT 65.360 195.320 65.620 195.640 ;
        RECT 63.980 191.580 64.240 191.900 ;
        RECT 64.900 189.880 65.160 190.200 ;
        RECT 64.960 189.180 65.100 189.880 ;
        RECT 65.420 189.180 65.560 195.320 ;
        RECT 65.880 194.280 66.020 198.040 ;
        RECT 66.800 197.000 66.940 199.060 ;
        RECT 66.740 196.680 67.000 197.000 ;
        RECT 65.820 193.960 66.080 194.280 ;
        RECT 64.900 188.860 65.160 189.180 ;
        RECT 65.360 188.860 65.620 189.180 ;
        RECT 65.420 188.580 65.560 188.860 ;
        RECT 61.220 188.180 61.480 188.500 ;
        RECT 65.420 188.440 66.020 188.580 ;
        RECT 61.280 187.480 61.420 188.180 ;
        RECT 61.220 187.160 61.480 187.480 ;
        RECT 65.360 187.160 65.620 187.480 ;
        RECT 61.280 186.460 61.420 187.160 ;
        RECT 61.880 186.625 63.760 186.995 ;
        RECT 61.220 186.140 61.480 186.460 ;
        RECT 63.980 185.460 64.240 185.780 ;
        RECT 61.220 185.120 61.480 185.440 ;
        RECT 61.280 183.060 61.420 185.120 ;
        RECT 64.040 183.400 64.180 185.460 ;
        RECT 65.420 185.440 65.560 187.160 ;
        RECT 65.360 185.120 65.620 185.440 ;
        RECT 64.440 184.780 64.700 185.100 ;
        RECT 63.980 183.080 64.240 183.400 ;
        RECT 60.300 182.740 60.560 183.060 ;
        RECT 61.220 182.740 61.480 183.060 ;
        RECT 59.380 181.720 59.640 182.040 ;
        RECT 58.910 179.485 59.190 179.855 ;
        RECT 58.450 161.805 58.730 162.175 ;
        RECT 57.540 160.980 57.800 161.125 ;
        RECT 58.000 161.010 58.260 161.330 ;
        RECT 58.980 160.700 59.120 179.485 ;
        RECT 58.520 160.560 59.120 160.700 ;
        RECT 58.520 160.530 58.660 160.560 ;
        RECT 58.165 160.390 58.660 160.530 ;
        RECT 57.080 159.960 57.340 160.280 ;
        RECT 54.780 158.260 55.040 158.580 ;
        RECT 55.700 157.920 55.960 158.240 ;
        RECT 54.780 157.240 55.040 157.560 ;
        RECT 54.840 155.180 54.980 157.240 ;
        RECT 55.760 155.520 55.900 157.920 ;
        RECT 55.700 155.200 55.960 155.520 ;
        RECT 56.620 155.200 56.880 155.520 ;
        RECT 54.780 154.860 55.040 155.180 ;
        RECT 54.840 152.800 54.980 154.860 ;
        RECT 55.760 153.140 55.900 155.200 ;
        RECT 55.700 152.820 55.960 153.140 ;
        RECT 54.780 152.480 55.040 152.800 ;
        RECT 54.840 150.420 54.980 152.480 ;
        RECT 55.240 150.780 55.500 151.100 ;
        RECT 55.300 150.420 55.440 150.780 ;
        RECT 55.760 150.760 55.900 152.820 ;
        RECT 56.160 152.480 56.420 152.800 ;
        RECT 55.700 150.440 55.960 150.760 ;
        RECT 56.220 150.420 56.360 152.480 ;
        RECT 54.780 150.100 55.040 150.420 ;
        RECT 55.240 150.100 55.500 150.420 ;
        RECT 56.160 150.100 56.420 150.420 ;
        RECT 56.160 149.420 56.420 149.740 ;
        RECT 55.700 149.080 55.960 149.400 ;
        RECT 54.780 148.060 55.040 148.380 ;
        RECT 54.320 147.380 54.580 147.700 ;
        RECT 54.840 142.940 54.980 148.060 ;
        RECT 55.760 147.360 55.900 149.080 ;
        RECT 56.220 147.360 56.360 149.420 ;
        RECT 55.700 147.040 55.960 147.360 ;
        RECT 56.160 147.040 56.420 147.360 ;
        RECT 56.220 143.960 56.360 147.040 ;
        RECT 56.680 147.020 56.820 155.200 ;
        RECT 56.620 146.700 56.880 147.020 ;
        RECT 56.680 146.535 56.820 146.700 ;
        RECT 56.610 146.165 56.890 146.535 ;
        RECT 56.160 143.640 56.420 143.960 ;
        RECT 54.780 142.620 55.040 142.940 ;
        RECT 54.320 141.260 54.580 141.580 ;
        RECT 54.380 139.880 54.520 141.260 ;
        RECT 54.780 140.920 55.040 141.240 ;
        RECT 54.320 139.560 54.580 139.880 ;
        RECT 53.920 138.800 54.520 138.940 ;
        RECT 53.400 136.840 53.660 137.160 ;
        RECT 50.180 136.500 50.440 136.820 ;
        RECT 51.100 136.500 51.360 136.820 ;
        RECT 52.020 136.500 52.280 136.820 ;
        RECT 50.180 135.820 50.440 136.140 ;
        RECT 50.240 133.760 50.380 135.820 ;
        RECT 50.180 133.440 50.440 133.760 ;
        RECT 51.160 131.040 51.300 136.500 ;
        RECT 52.080 134.780 52.220 136.500 ;
        RECT 52.480 136.160 52.740 136.480 ;
        RECT 52.940 136.160 53.200 136.480 ;
        RECT 52.020 134.460 52.280 134.780 ;
        RECT 52.540 131.720 52.680 136.160 ;
        RECT 53.000 135.800 53.140 136.160 ;
        RECT 52.940 135.480 53.200 135.800 ;
        RECT 53.000 134.780 53.140 135.480 ;
        RECT 52.940 134.460 53.200 134.780 ;
        RECT 52.480 131.400 52.740 131.720 ;
        RECT 53.000 131.380 53.140 134.460 ;
        RECT 53.400 133.440 53.660 133.760 ;
        RECT 53.460 132.060 53.600 133.440 ;
        RECT 53.400 131.740 53.660 132.060 ;
        RECT 52.940 131.060 53.200 131.380 ;
        RECT 51.100 130.950 51.360 131.040 ;
        RECT 50.700 130.810 51.360 130.950 ;
        RECT 50.180 130.380 50.440 130.700 ;
        RECT 49.720 128.000 49.980 128.320 ;
        RECT 49.780 125.260 49.920 128.000 ;
        RECT 50.240 127.640 50.380 130.380 ;
        RECT 50.180 127.320 50.440 127.640 ;
        RECT 50.240 126.280 50.380 127.320 ;
        RECT 50.180 125.960 50.440 126.280 ;
        RECT 50.700 125.940 50.840 130.810 ;
        RECT 51.100 130.720 51.360 130.810 ;
        RECT 54.380 130.360 54.520 138.800 ;
        RECT 51.100 130.040 51.360 130.360 ;
        RECT 54.320 130.040 54.580 130.360 ;
        RECT 51.160 128.660 51.300 130.040 ;
        RECT 54.380 129.340 54.520 130.040 ;
        RECT 54.320 129.020 54.580 129.340 ;
        RECT 51.100 128.340 51.360 128.660 ;
        RECT 50.640 125.620 50.900 125.940 ;
        RECT 53.400 125.455 53.660 125.600 ;
        RECT 49.720 124.940 49.980 125.260 ;
        RECT 53.390 125.085 53.670 125.455 ;
        RECT 49.780 122.880 49.920 124.940 ;
        RECT 53.460 123.220 53.600 125.085 ;
        RECT 53.400 122.900 53.660 123.220 ;
        RECT 49.720 122.560 49.980 122.880 ;
        RECT 49.780 120.500 49.920 122.560 ;
        RECT 49.720 120.180 49.980 120.500 ;
        RECT 50.180 120.180 50.440 120.500 ;
        RECT 49.260 119.160 49.520 119.480 ;
        RECT 46.880 118.625 48.760 118.995 ;
        RECT 49.780 117.440 49.920 120.180 ;
        RECT 50.240 118.120 50.380 120.180 ;
        RECT 54.840 120.160 54.980 140.920 ;
        RECT 55.300 140.220 55.900 140.300 ;
        RECT 55.300 140.160 55.960 140.220 ;
        RECT 55.300 120.500 55.440 140.160 ;
        RECT 55.700 139.900 55.960 140.160 ;
        RECT 55.700 139.220 55.960 139.540 ;
        RECT 55.760 137.500 55.900 139.220 ;
        RECT 55.700 137.180 55.960 137.500 ;
        RECT 55.700 136.500 55.960 136.820 ;
        RECT 55.760 126.620 55.900 136.500 ;
        RECT 56.220 129.340 56.360 143.640 ;
        RECT 56.620 142.280 56.880 142.600 ;
        RECT 56.680 137.500 56.820 142.280 ;
        RECT 57.140 141.920 57.280 159.960 ;
        RECT 58.165 159.340 58.305 160.390 ;
        RECT 58.920 159.960 59.180 160.280 ;
        RECT 59.440 160.140 59.580 181.720 ;
        RECT 61.280 180.680 61.420 182.740 ;
        RECT 61.880 181.185 63.760 181.555 ;
        RECT 61.220 180.360 61.480 180.680 ;
        RECT 60.760 180.020 61.020 180.340 ;
        RECT 60.300 179.000 60.560 179.320 ;
        RECT 60.360 177.620 60.500 179.000 ;
        RECT 60.300 177.300 60.560 177.620 ;
        RECT 60.300 173.560 60.560 173.880 ;
        RECT 60.360 172.180 60.500 173.560 ;
        RECT 60.300 171.860 60.560 172.180 ;
        RECT 59.840 168.800 60.100 169.120 ;
        RECT 59.900 164.020 60.040 168.800 ;
        RECT 60.360 164.100 60.500 171.860 ;
        RECT 60.820 171.160 60.960 180.020 ;
        RECT 63.980 179.680 64.240 180.000 ;
        RECT 61.220 176.280 61.480 176.600 ;
        RECT 61.280 174.900 61.420 176.280 ;
        RECT 61.880 175.745 63.760 176.115 ;
        RECT 64.040 175.580 64.180 179.680 ;
        RECT 63.980 175.260 64.240 175.580 ;
        RECT 61.220 174.580 61.480 174.900 ;
        RECT 63.520 174.580 63.780 174.900 ;
        RECT 63.580 172.940 63.720 174.580 ;
        RECT 64.500 173.790 64.640 184.780 ;
        RECT 65.420 183.740 65.560 185.120 ;
        RECT 65.880 183.740 66.020 188.440 ;
        RECT 65.360 183.420 65.620 183.740 ;
        RECT 65.820 183.420 66.080 183.740 ;
        RECT 64.900 179.000 65.160 179.320 ;
        RECT 66.280 179.000 66.540 179.320 ;
        RECT 64.960 174.560 65.100 179.000 ;
        RECT 64.900 174.240 65.160 174.560 ;
        RECT 62.660 172.860 63.720 172.940 ;
        RECT 62.600 172.800 63.720 172.860 ;
        RECT 62.600 172.540 62.860 172.800 ;
        RECT 63.580 172.180 63.720 172.800 ;
        RECT 64.040 173.650 64.640 173.790 ;
        RECT 61.220 171.860 61.480 172.180 ;
        RECT 63.520 171.860 63.780 172.180 ;
        RECT 60.760 170.840 61.020 171.160 ;
        RECT 60.820 169.800 60.960 170.840 ;
        RECT 60.760 169.480 61.020 169.800 ;
        RECT 61.280 167.615 61.420 171.860 ;
        RECT 64.040 171.840 64.180 173.650 ;
        RECT 65.360 173.560 65.620 173.880 ;
        RECT 63.980 171.520 64.240 171.840 ;
        RECT 64.900 170.840 65.160 171.160 ;
        RECT 61.880 170.305 63.760 170.675 ;
        RECT 61.210 167.245 61.490 167.615 ;
        RECT 64.960 167.420 65.100 170.840 ;
        RECT 65.420 170.140 65.560 173.560 ;
        RECT 65.360 169.820 65.620 170.140 ;
        RECT 64.900 167.100 65.160 167.420 ;
        RECT 61.880 164.865 63.760 165.235 ;
        RECT 59.840 163.700 60.100 164.020 ;
        RECT 60.360 163.960 61.880 164.100 ;
        RECT 65.360 164.040 65.620 164.360 ;
        RECT 60.300 163.360 60.560 163.680 ;
        RECT 59.830 162.485 60.110 162.855 ;
        RECT 59.900 161.300 60.040 162.485 ;
        RECT 60.360 161.300 60.500 163.360 ;
        RECT 61.220 162.680 61.480 163.000 ;
        RECT 61.280 161.300 61.420 162.680 ;
        RECT 61.740 161.300 61.880 163.960 ;
        RECT 65.420 163.680 65.560 164.040 ;
        RECT 64.890 163.165 65.170 163.535 ;
        RECT 65.360 163.360 65.620 163.680 ;
        RECT 64.900 163.020 65.160 163.165 ;
        RECT 63.980 162.680 64.240 163.000 ;
        RECT 65.360 162.680 65.620 163.000 ;
        RECT 64.040 162.060 64.180 162.680 ;
        RECT 64.040 161.920 64.640 162.060 ;
        RECT 59.840 160.980 60.100 161.300 ;
        RECT 60.300 160.980 60.560 161.300 ;
        RECT 61.220 160.980 61.480 161.300 ;
        RECT 61.680 160.980 61.940 161.300 ;
        RECT 63.980 160.980 64.240 161.300 ;
        RECT 60.760 160.300 61.020 160.620 ;
        RECT 59.440 160.000 60.040 160.140 ;
        RECT 58.060 159.200 58.305 159.340 ;
        RECT 57.540 142.620 57.800 142.940 ;
        RECT 57.080 141.600 57.340 141.920 ;
        RECT 56.620 137.180 56.880 137.500 ;
        RECT 57.080 136.160 57.340 136.480 ;
        RECT 57.140 134.100 57.280 136.160 ;
        RECT 57.080 133.780 57.340 134.100 ;
        RECT 57.140 131.040 57.280 133.780 ;
        RECT 57.600 132.060 57.740 142.620 ;
        RECT 58.060 139.540 58.200 159.200 ;
        RECT 58.460 153.500 58.720 153.820 ;
        RECT 58.520 147.700 58.660 153.500 ;
        RECT 58.980 149.140 59.120 159.960 ;
        RECT 59.380 155.200 59.640 155.520 ;
        RECT 59.440 149.740 59.580 155.200 ;
        RECT 59.380 149.420 59.640 149.740 ;
        RECT 58.980 149.000 59.580 149.140 ;
        RECT 58.460 147.380 58.720 147.700 ;
        RECT 58.460 141.260 58.720 141.580 ;
        RECT 58.520 140.220 58.660 141.260 ;
        RECT 58.460 139.900 58.720 140.220 ;
        RECT 59.440 139.540 59.580 149.000 ;
        RECT 59.900 142.260 60.040 160.000 ;
        RECT 60.820 158.240 60.960 160.300 ;
        RECT 61.880 159.425 63.760 159.795 ;
        RECT 60.760 157.920 61.020 158.240 ;
        RECT 61.680 157.920 61.940 158.240 ;
        RECT 61.740 156.540 61.880 157.920 ;
        RECT 64.040 156.620 64.180 160.980 ;
        RECT 61.680 156.220 61.940 156.540 ;
        RECT 63.580 156.480 64.180 156.620 ;
        RECT 60.760 155.880 61.020 156.200 ;
        RECT 60.300 154.520 60.560 154.840 ;
        RECT 60.360 152.460 60.500 154.520 ;
        RECT 60.300 152.140 60.560 152.460 ;
        RECT 60.820 150.760 60.960 155.880 ;
        RECT 63.580 155.860 63.720 156.480 ;
        RECT 63.520 155.540 63.780 155.860 ;
        RECT 61.220 155.200 61.480 155.520 ;
        RECT 61.280 153.140 61.420 155.200 ;
        RECT 61.880 153.985 63.760 154.355 ;
        RECT 61.220 152.820 61.480 153.140 ;
        RECT 63.980 152.820 64.240 153.140 ;
        RECT 60.760 150.440 61.020 150.760 ;
        RECT 61.280 147.360 61.420 152.820 ;
        RECT 61.880 148.545 63.760 148.915 ;
        RECT 61.220 147.040 61.480 147.360 ;
        RECT 62.590 145.485 62.870 145.855 ;
        RECT 64.040 145.660 64.180 152.820 ;
        RECT 62.660 145.320 62.800 145.485 ;
        RECT 63.980 145.340 64.240 145.660 ;
        RECT 60.750 144.805 61.030 145.175 ;
        RECT 62.600 145.000 62.860 145.320 ;
        RECT 59.840 141.940 60.100 142.260 ;
        RECT 60.300 140.920 60.560 141.240 ;
        RECT 59.840 139.560 60.100 139.880 ;
        RECT 58.000 139.220 58.260 139.540 ;
        RECT 58.920 139.220 59.180 139.540 ;
        RECT 59.380 139.220 59.640 139.540 ;
        RECT 58.460 138.200 58.720 138.520 ;
        RECT 57.540 131.740 57.800 132.060 ;
        RECT 57.080 130.720 57.340 131.040 ;
        RECT 56.160 129.020 56.420 129.340 ;
        RECT 56.620 128.680 56.880 129.000 ;
        RECT 57.140 128.740 57.280 130.720 ;
        RECT 55.700 126.300 55.960 126.620 ;
        RECT 55.760 125.940 55.900 126.300 ;
        RECT 55.700 125.620 55.960 125.940 ;
        RECT 56.680 123.900 56.820 128.680 ;
        RECT 57.140 128.600 57.740 128.740 ;
        RECT 57.080 128.000 57.340 128.320 ;
        RECT 57.140 125.940 57.280 128.000 ;
        RECT 57.080 125.620 57.340 125.940 ;
        RECT 57.600 125.600 57.740 128.600 ;
        RECT 58.520 125.600 58.660 138.200 ;
        RECT 58.980 134.780 59.120 139.220 ;
        RECT 58.920 134.460 59.180 134.780 ;
        RECT 59.900 130.360 60.040 139.560 ;
        RECT 60.360 134.440 60.500 140.920 ;
        RECT 60.300 134.120 60.560 134.440 ;
        RECT 60.820 133.760 60.960 144.805 ;
        RECT 63.980 144.660 64.240 144.980 ;
        RECT 61.880 143.105 63.760 143.475 ;
        RECT 64.040 139.620 64.180 144.660 ;
        RECT 64.500 141.920 64.640 161.920 ;
        RECT 64.900 158.600 65.160 158.920 ;
        RECT 64.960 144.980 65.100 158.600 ;
        RECT 64.900 144.660 65.160 144.980 ;
        RECT 64.440 141.600 64.700 141.920 ;
        RECT 64.040 139.480 64.640 139.620 ;
        RECT 65.420 139.540 65.560 162.680 ;
        RECT 65.820 160.300 66.080 160.620 ;
        RECT 65.880 158.240 66.020 160.300 ;
        RECT 65.820 157.920 66.080 158.240 ;
        RECT 65.820 155.200 66.080 155.520 ;
        RECT 65.880 150.080 66.020 155.200 ;
        RECT 65.820 149.760 66.080 150.080 ;
        RECT 65.880 145.320 66.020 149.760 ;
        RECT 65.820 145.000 66.080 145.320 ;
        RECT 65.880 142.600 66.020 145.000 ;
        RECT 65.820 142.280 66.080 142.600 ;
        RECT 65.820 139.900 66.080 140.220 ;
        RECT 63.980 138.200 64.240 138.520 ;
        RECT 61.880 137.665 63.760 138.035 ;
        RECT 61.670 136.645 61.950 137.015 ;
        RECT 61.740 134.100 61.880 136.645 ;
        RECT 64.040 134.100 64.180 138.200 ;
        RECT 64.500 136.480 64.640 139.480 ;
        RECT 65.360 139.220 65.620 139.540 ;
        RECT 65.880 138.520 66.020 139.900 ;
        RECT 66.340 139.200 66.480 179.000 ;
        RECT 66.800 177.620 66.940 196.680 ;
        RECT 70.880 195.320 71.140 195.640 ;
        RECT 70.940 194.280 71.080 195.320 ;
        RECT 71.400 194.280 71.540 201.440 ;
        RECT 72.320 199.380 72.460 204.160 ;
        RECT 73.640 201.100 73.900 201.420 ;
        RECT 73.700 199.380 73.840 201.100 ;
        RECT 72.260 199.060 72.520 199.380 ;
        RECT 73.640 199.060 73.900 199.380 ;
        RECT 70.880 193.960 71.140 194.280 ;
        RECT 71.340 193.960 71.600 194.280 ;
        RECT 69.500 190.900 69.760 191.220 ;
        RECT 67.660 188.180 67.920 188.500 ;
        RECT 68.120 188.180 68.380 188.500 ;
        RECT 67.720 186.460 67.860 188.180 ;
        RECT 67.660 186.140 67.920 186.460 ;
        RECT 67.650 184.925 67.930 185.295 ;
        RECT 67.660 184.780 67.920 184.925 ;
        RECT 68.180 183.740 68.320 188.180 ;
        RECT 69.560 186.120 69.700 190.900 ;
        RECT 71.400 188.500 71.540 193.960 ;
        RECT 73.180 193.620 73.440 193.940 ;
        RECT 71.800 192.600 72.060 192.920 ;
        RECT 71.860 188.500 72.000 192.600 ;
        RECT 73.240 188.840 73.380 193.620 ;
        RECT 75.540 193.600 75.680 204.160 ;
        RECT 76.000 199.720 76.140 206.970 ;
        RECT 76.860 206.880 77.120 206.970 ;
        RECT 79.160 206.880 79.420 207.200 ;
        RECT 76.400 206.200 76.660 206.520 ;
        RECT 76.460 205.500 76.600 206.200 ;
        RECT 76.880 205.665 78.760 206.035 ;
        RECT 76.400 205.180 76.660 205.500 ;
        RECT 76.400 203.480 76.660 203.800 ;
        RECT 76.460 200.060 76.600 203.480 ;
        RECT 79.220 202.780 79.360 206.880 ;
        RECT 80.140 205.500 80.280 207.220 ;
        RECT 80.080 205.180 80.340 205.500 ;
        RECT 81.000 204.500 81.260 204.820 ;
        RECT 80.080 204.160 80.340 204.480 ;
        RECT 79.160 202.460 79.420 202.780 ;
        RECT 79.160 201.780 79.420 202.100 ;
        RECT 76.880 200.225 78.760 200.595 ;
        RECT 79.220 200.060 79.360 201.780 ;
        RECT 79.620 201.440 79.880 201.760 ;
        RECT 76.400 199.740 76.660 200.060 ;
        RECT 79.160 199.740 79.420 200.060 ;
        RECT 75.940 199.400 76.200 199.720 ;
        RECT 76.000 194.620 76.140 199.400 ;
        RECT 76.400 199.060 76.660 199.380 ;
        RECT 78.700 199.060 78.960 199.380 ;
        RECT 75.940 194.300 76.200 194.620 ;
        RECT 76.460 194.530 76.600 199.060 ;
        RECT 78.760 198.700 78.900 199.060 ;
        RECT 79.220 198.700 79.360 199.740 ;
        RECT 79.680 199.380 79.820 201.440 ;
        RECT 80.140 200.060 80.280 204.160 ;
        RECT 81.060 202.440 81.200 204.500 ;
        RECT 81.000 202.120 81.260 202.440 ;
        RECT 81.520 200.060 81.660 207.220 ;
        RECT 82.380 206.540 82.640 206.860 ;
        RECT 82.440 205.500 82.580 206.540 ;
        RECT 82.380 205.180 82.640 205.500 ;
        RECT 82.380 200.760 82.640 201.080 ;
        RECT 80.080 199.740 80.340 200.060 ;
        RECT 81.460 199.740 81.720 200.060 ;
        RECT 79.620 199.060 79.880 199.380 ;
        RECT 82.440 199.040 82.580 200.760 ;
        RECT 82.380 198.720 82.640 199.040 ;
        RECT 78.700 198.380 78.960 198.700 ;
        RECT 79.160 198.380 79.420 198.700 ;
        RECT 78.760 197.000 78.900 198.380 ;
        RECT 78.700 196.680 78.960 197.000 ;
        RECT 76.880 194.785 78.760 195.155 ;
        RECT 76.460 194.390 77.520 194.530 ;
        RECT 77.380 193.940 77.520 194.390 ;
        RECT 77.780 194.300 78.040 194.620 ;
        RECT 77.840 193.940 77.980 194.300 ;
        RECT 77.320 193.620 77.580 193.940 ;
        RECT 77.780 193.620 78.040 193.940 ;
        RECT 75.480 193.280 75.740 193.600 ;
        RECT 75.020 192.940 75.280 193.260 ;
        RECT 73.640 192.600 73.900 192.920 ;
        RECT 73.700 190.540 73.840 192.600 ;
        RECT 73.640 190.220 73.900 190.540 ;
        RECT 73.180 188.520 73.440 188.840 ;
        RECT 71.340 188.180 71.600 188.500 ;
        RECT 71.800 188.180 72.060 188.500 ;
        RECT 69.500 185.800 69.760 186.120 ;
        RECT 69.560 185.100 69.700 185.800 ;
        RECT 69.500 184.780 69.760 185.100 ;
        RECT 68.120 183.420 68.380 183.740 ;
        RECT 72.260 183.420 72.520 183.740 ;
        RECT 68.180 180.340 68.320 183.420 ;
        RECT 70.420 183.080 70.680 183.400 ;
        RECT 69.040 182.060 69.300 182.380 ;
        RECT 69.100 181.020 69.240 182.060 ;
        RECT 69.960 181.720 70.220 182.040 ;
        RECT 69.040 180.700 69.300 181.020 ;
        RECT 68.120 180.020 68.380 180.340 ;
        RECT 69.100 180.000 69.240 180.700 ;
        RECT 70.020 180.340 70.160 181.720 ;
        RECT 69.960 180.020 70.220 180.340 ;
        RECT 69.040 179.680 69.300 180.000 ;
        RECT 67.660 179.000 67.920 179.320 ;
        RECT 67.720 178.300 67.860 179.000 ;
        RECT 70.480 178.300 70.620 183.080 ;
        RECT 72.320 181.020 72.460 183.420 ;
        RECT 72.260 180.700 72.520 181.020 ;
        RECT 73.240 179.060 73.380 188.520 ;
        RECT 73.700 182.040 73.840 190.220 ;
        RECT 74.560 189.880 74.820 190.200 ;
        RECT 74.620 183.740 74.760 189.880 ;
        RECT 75.080 186.120 75.220 192.940 ;
        RECT 75.540 191.220 75.680 193.280 ;
        RECT 75.480 190.900 75.740 191.220 ;
        RECT 75.540 188.500 75.680 190.900 ;
        RECT 77.380 190.880 77.520 193.620 ;
        RECT 77.320 190.560 77.580 190.880 ;
        RECT 77.840 190.540 77.980 193.620 ;
        RECT 79.220 193.260 79.360 198.380 ;
        RECT 80.540 198.040 80.800 198.360 ;
        RECT 79.160 192.940 79.420 193.260 ;
        RECT 80.080 192.940 80.340 193.260 ;
        RECT 78.700 192.775 78.960 192.920 ;
        RECT 78.690 192.405 78.970 192.775 ;
        RECT 79.220 191.560 79.360 192.940 ;
        RECT 79.160 191.240 79.420 191.560 ;
        RECT 77.780 190.220 78.040 190.540 ;
        RECT 76.880 189.345 78.760 189.715 ;
        RECT 79.220 189.180 79.360 191.240 ;
        RECT 80.140 191.220 80.280 192.940 ;
        RECT 80.080 190.900 80.340 191.220 ;
        RECT 79.620 190.220 79.880 190.540 ;
        RECT 79.160 188.860 79.420 189.180 ;
        RECT 79.680 188.500 79.820 190.220 ;
        RECT 80.140 188.500 80.280 190.900 ;
        RECT 75.480 188.180 75.740 188.500 ;
        RECT 77.780 188.180 78.040 188.500 ;
        RECT 79.620 188.180 79.880 188.500 ;
        RECT 80.080 188.180 80.340 188.500 ;
        RECT 75.020 185.800 75.280 186.120 ;
        RECT 74.560 183.420 74.820 183.740 ;
        RECT 75.020 183.080 75.280 183.400 ;
        RECT 73.640 181.720 73.900 182.040 ;
        RECT 73.700 180.000 73.840 181.720 ;
        RECT 74.560 180.700 74.820 181.020 ;
        RECT 73.640 179.680 73.900 180.000 ;
        RECT 74.100 179.680 74.360 180.000 ;
        RECT 74.160 179.060 74.300 179.680 ;
        RECT 73.240 178.920 74.300 179.060 ;
        RECT 67.660 177.980 67.920 178.300 ;
        RECT 70.420 177.980 70.680 178.300 ;
        RECT 68.580 177.640 68.840 177.960 ;
        RECT 66.740 177.300 67.000 177.620 ;
        RECT 67.660 176.960 67.920 177.280 ;
        RECT 66.740 168.120 67.000 168.440 ;
        RECT 66.800 164.020 66.940 168.120 ;
        RECT 67.200 166.420 67.460 166.740 ;
        RECT 67.260 164.700 67.400 166.420 ;
        RECT 67.720 166.140 67.860 176.960 ;
        RECT 68.120 176.280 68.380 176.600 ;
        RECT 68.180 172.860 68.320 176.280 ;
        RECT 68.120 172.540 68.380 172.860 ;
        RECT 68.180 167.080 68.320 172.540 ;
        RECT 68.120 166.760 68.380 167.080 ;
        RECT 67.720 166.000 68.320 166.140 ;
        RECT 67.200 164.380 67.460 164.700 ;
        RECT 66.740 163.700 67.000 164.020 ;
        RECT 67.200 163.360 67.460 163.680 ;
        RECT 67.260 161.640 67.400 163.360 ;
        RECT 68.180 163.340 68.320 166.000 ;
        RECT 68.120 163.020 68.380 163.340 ;
        RECT 68.640 162.740 68.780 177.640 ;
        RECT 69.960 174.580 70.220 174.900 ;
        RECT 70.020 171.160 70.160 174.580 ;
        RECT 70.420 173.900 70.680 174.220 ;
        RECT 69.960 170.840 70.220 171.160 ;
        RECT 69.040 168.120 69.300 168.440 ;
        RECT 69.100 164.360 69.240 168.120 ;
        RECT 70.020 166.400 70.160 170.840 ;
        RECT 70.480 168.780 70.620 173.900 ;
        RECT 72.260 173.560 72.520 173.880 ;
        RECT 72.320 172.520 72.460 173.560 ;
        RECT 72.260 172.200 72.520 172.520 ;
        RECT 70.420 168.460 70.680 168.780 ;
        RECT 73.640 168.460 73.900 168.780 ;
        RECT 73.170 166.565 73.450 166.935 ;
        RECT 69.960 166.080 70.220 166.400 ;
        RECT 72.260 166.255 72.520 166.400 ;
        RECT 72.250 165.885 72.530 166.255 ;
        RECT 69.040 164.040 69.300 164.360 ;
        RECT 69.100 163.680 69.240 164.040 ;
        RECT 69.040 163.360 69.300 163.680 ;
        RECT 69.500 163.535 69.760 163.680 ;
        RECT 69.490 163.165 69.770 163.535 ;
        RECT 67.720 162.600 68.780 162.740 ;
        RECT 67.200 161.320 67.460 161.640 ;
        RECT 67.720 161.300 67.860 162.600 ;
        RECT 67.660 160.980 67.920 161.300 ;
        RECT 69.040 160.980 69.300 161.300 ;
        RECT 67.660 159.960 67.920 160.280 ;
        RECT 67.720 157.900 67.860 159.960 ;
        RECT 67.660 157.580 67.920 157.900 ;
        RECT 69.100 156.540 69.240 160.980 ;
        RECT 70.420 159.960 70.680 160.280 ;
        RECT 70.480 158.580 70.620 159.960 ;
        RECT 70.420 158.260 70.680 158.580 ;
        RECT 69.040 156.220 69.300 156.540 ;
        RECT 66.740 155.880 67.000 156.200 ;
        RECT 66.800 153.820 66.940 155.880 ;
        RECT 72.320 155.860 72.460 165.885 ;
        RECT 72.720 165.400 72.980 165.720 ;
        RECT 72.780 163.680 72.920 165.400 ;
        RECT 72.720 163.360 72.980 163.680 ;
        RECT 73.240 161.640 73.380 166.565 ;
        RECT 73.700 164.700 73.840 168.460 ;
        RECT 73.640 164.380 73.900 164.700 ;
        RECT 74.160 163.680 74.300 178.920 ;
        RECT 74.620 176.940 74.760 180.700 ;
        RECT 75.080 180.680 75.220 183.080 ;
        RECT 75.540 182.720 75.680 188.180 ;
        RECT 77.840 185.100 77.980 188.180 ;
        RECT 79.620 187.500 79.880 187.820 ;
        RECT 76.400 184.780 76.660 185.100 ;
        RECT 77.780 184.780 78.040 185.100 ;
        RECT 75.480 182.400 75.740 182.720 ;
        RECT 76.460 182.290 76.600 184.780 ;
        RECT 76.880 183.905 78.760 184.275 ;
        RECT 77.780 183.080 78.040 183.400 ;
        RECT 77.320 182.290 77.580 182.380 ;
        RECT 76.460 182.150 77.580 182.290 ;
        RECT 77.320 182.060 77.580 182.150 ;
        RECT 75.020 180.360 75.280 180.680 ;
        RECT 75.470 180.165 75.750 180.535 ;
        RECT 75.540 178.300 75.680 180.165 ;
        RECT 77.840 180.000 77.980 183.080 ;
        RECT 78.240 182.740 78.500 183.060 ;
        RECT 78.300 180.340 78.440 182.740 ;
        RECT 79.160 182.060 79.420 182.380 ;
        RECT 78.700 181.720 78.960 182.040 ;
        RECT 78.760 180.680 78.900 181.720 ;
        RECT 78.700 180.360 78.960 180.680 ;
        RECT 78.240 180.020 78.500 180.340 ;
        RECT 76.400 179.680 76.660 180.000 ;
        RECT 77.780 179.680 78.040 180.000 ;
        RECT 76.460 178.300 76.600 179.680 ;
        RECT 76.880 178.465 78.760 178.835 ;
        RECT 75.480 177.980 75.740 178.300 ;
        RECT 76.400 177.980 76.660 178.300 ;
        RECT 75.020 177.300 75.280 177.620 ;
        RECT 74.560 176.620 74.820 176.940 ;
        RECT 75.080 174.900 75.220 177.300 ;
        RECT 75.540 175.240 75.680 177.980 ;
        RECT 76.460 177.620 76.600 177.980 ;
        RECT 77.320 177.640 77.580 177.960 ;
        RECT 76.400 177.300 76.660 177.620 ;
        RECT 76.400 176.280 76.660 176.600 ;
        RECT 75.480 174.920 75.740 175.240 ;
        RECT 75.020 174.580 75.280 174.900 ;
        RECT 74.100 163.360 74.360 163.680 ;
        RECT 73.180 161.320 73.440 161.640 ;
        RECT 74.160 161.300 74.300 163.360 ;
        RECT 74.100 160.980 74.360 161.300 ;
        RECT 74.160 160.140 74.300 160.980 ;
        RECT 74.160 160.000 74.760 160.140 ;
        RECT 74.620 158.920 74.760 160.000 ;
        RECT 74.560 158.600 74.820 158.920 ;
        RECT 73.640 157.920 73.900 158.240 ;
        RECT 69.960 155.540 70.220 155.860 ;
        RECT 70.880 155.770 71.140 155.860 ;
        RECT 70.480 155.630 71.140 155.770 ;
        RECT 66.740 153.500 67.000 153.820 ;
        RECT 67.200 151.800 67.460 152.120 ;
        RECT 67.260 150.420 67.400 151.800 ;
        RECT 67.200 150.100 67.460 150.420 ;
        RECT 67.260 147.700 67.400 150.100 ;
        RECT 67.660 149.760 67.920 150.080 ;
        RECT 67.200 147.380 67.460 147.700 ;
        RECT 67.200 146.360 67.460 146.680 ;
        RECT 67.260 144.980 67.400 146.360 ;
        RECT 67.200 144.660 67.460 144.980 ;
        RECT 67.720 144.640 67.860 149.760 ;
        RECT 68.120 149.420 68.380 149.740 ;
        RECT 68.180 144.980 68.320 149.420 ;
        RECT 70.020 148.380 70.160 155.540 ;
        RECT 70.480 150.420 70.620 155.630 ;
        RECT 70.880 155.540 71.140 155.630 ;
        RECT 72.260 155.540 72.520 155.860 ;
        RECT 70.880 154.520 71.140 154.840 ;
        RECT 70.940 152.460 71.080 154.520 ;
        RECT 73.700 153.140 73.840 157.920 ;
        RECT 73.640 152.820 73.900 153.140 ;
        RECT 73.700 152.460 73.840 152.820 ;
        RECT 70.880 152.140 71.140 152.460 ;
        RECT 73.640 152.140 73.900 152.460 ;
        RECT 70.880 150.780 71.140 151.100 ;
        RECT 70.420 150.100 70.680 150.420 ;
        RECT 69.960 148.060 70.220 148.380 ;
        RECT 70.020 147.360 70.160 148.060 ;
        RECT 69.960 147.040 70.220 147.360 ;
        RECT 68.120 144.660 68.380 144.980 ;
        RECT 69.960 144.660 70.220 144.980 ;
        RECT 67.660 144.495 67.920 144.640 ;
        RECT 67.650 144.125 67.930 144.495 ;
        RECT 66.740 143.640 67.000 143.960 ;
        RECT 66.800 142.260 66.940 143.640 ;
        RECT 66.740 141.940 67.000 142.260 ;
        RECT 67.720 141.920 67.860 144.125 ;
        RECT 67.200 141.600 67.460 141.920 ;
        RECT 67.660 141.600 67.920 141.920 ;
        RECT 67.260 141.240 67.400 141.600 ;
        RECT 67.200 140.920 67.460 141.240 ;
        RECT 66.280 138.880 66.540 139.200 ;
        RECT 67.200 138.540 67.460 138.860 ;
        RECT 65.360 138.200 65.620 138.520 ;
        RECT 65.820 138.200 66.080 138.520 ;
        RECT 64.440 136.335 64.700 136.480 ;
        RECT 64.430 135.965 64.710 136.335 ;
        RECT 64.900 134.120 65.160 134.440 ;
        RECT 61.680 133.780 61.940 134.100 ;
        RECT 63.980 133.780 64.240 134.100 ;
        RECT 60.760 133.440 61.020 133.760 ;
        RECT 61.220 132.760 61.480 133.080 ;
        RECT 59.840 130.040 60.100 130.360 ;
        RECT 59.900 126.620 60.040 130.040 ;
        RECT 59.840 126.300 60.100 126.620 ;
        RECT 57.540 125.280 57.800 125.600 ;
        RECT 58.460 125.280 58.720 125.600 ;
        RECT 56.620 123.580 56.880 123.900 ;
        RECT 61.280 123.220 61.420 132.760 ;
        RECT 61.880 132.225 63.760 132.595 ;
        RECT 64.960 130.700 65.100 134.120 ;
        RECT 64.900 130.380 65.160 130.700 ;
        RECT 64.440 130.040 64.700 130.360 ;
        RECT 64.500 128.660 64.640 130.040 ;
        RECT 64.960 129.340 65.100 130.380 ;
        RECT 64.900 129.020 65.160 129.340 ;
        RECT 65.420 128.740 65.560 138.200 ;
        RECT 65.880 134.100 66.020 138.200 ;
        RECT 67.260 134.100 67.400 138.540 ;
        RECT 67.720 138.520 67.860 141.600 ;
        RECT 68.180 141.240 68.320 144.660 ;
        RECT 69.500 142.620 69.760 142.940 ;
        RECT 68.120 140.920 68.380 141.240 ;
        RECT 68.180 139.540 68.320 140.920 ;
        RECT 69.040 139.900 69.300 140.220 ;
        RECT 68.120 139.220 68.380 139.540 ;
        RECT 67.660 138.200 67.920 138.520 ;
        RECT 68.180 134.780 68.320 139.220 ;
        RECT 68.120 134.460 68.380 134.780 ;
        RECT 65.820 133.780 66.080 134.100 ;
        RECT 67.200 133.780 67.460 134.100 ;
        RECT 68.120 133.440 68.380 133.760 ;
        RECT 68.180 131.380 68.320 133.440 ;
        RECT 68.580 132.760 68.840 133.080 ;
        RECT 68.120 131.060 68.380 131.380 ;
        RECT 68.640 130.700 68.780 132.760 ;
        RECT 68.580 130.380 68.840 130.700 ;
        RECT 66.280 130.040 66.540 130.360 ;
        RECT 64.440 128.340 64.700 128.660 ;
        RECT 64.960 128.600 65.560 128.740 ;
        RECT 66.340 128.660 66.480 130.040 ;
        RECT 63.980 127.320 64.240 127.640 ;
        RECT 61.880 126.785 63.760 127.155 ;
        RECT 64.040 126.020 64.180 127.320 ;
        RECT 63.580 125.880 64.180 126.020 ;
        RECT 63.580 125.260 63.720 125.880 ;
        RECT 63.520 124.940 63.780 125.260 ;
        RECT 64.960 124.920 65.100 128.600 ;
        RECT 65.820 128.340 66.080 128.660 ;
        RECT 66.280 128.340 66.540 128.660 ;
        RECT 64.900 124.600 65.160 124.920 ;
        RECT 65.880 123.220 66.020 128.340 ;
        RECT 66.280 127.320 66.540 127.640 ;
        RECT 66.340 125.940 66.480 127.320 ;
        RECT 66.280 125.620 66.540 125.940 ;
        RECT 68.580 125.280 68.840 125.600 ;
        RECT 61.220 122.900 61.480 123.220 ;
        RECT 65.820 122.900 66.080 123.220 ;
        RECT 65.360 121.880 65.620 122.200 ;
        RECT 61.880 121.345 63.760 121.715 ;
        RECT 65.420 120.500 65.560 121.880 ;
        RECT 55.240 120.180 55.500 120.500 ;
        RECT 61.220 120.180 61.480 120.500 ;
        RECT 65.360 120.180 65.620 120.500 ;
        RECT 53.860 119.840 54.120 120.160 ;
        RECT 54.780 119.840 55.040 120.160 ;
        RECT 53.920 118.460 54.060 119.840 ;
        RECT 59.840 119.160 60.100 119.480 ;
        RECT 53.860 118.140 54.120 118.460 ;
        RECT 50.180 117.800 50.440 118.120 ;
        RECT 49.720 117.120 49.980 117.440 ;
        RECT 51.100 117.120 51.360 117.440 ;
        RECT 49.780 115.060 49.920 117.120 ;
        RECT 49.720 114.740 49.980 115.060 ;
        RECT 46.880 113.185 48.760 113.555 ;
        RECT 51.160 104.340 51.300 117.120 ;
        RECT 53.920 114.720 54.060 118.140 ;
        RECT 59.900 118.120 60.040 119.160 ;
        RECT 58.000 117.800 58.260 118.120 ;
        RECT 59.840 117.800 60.100 118.120 ;
        RECT 56.160 117.120 56.420 117.440 ;
        RECT 53.860 114.400 54.120 114.720 ;
        RECT 56.220 104.340 56.360 117.120 ;
        RECT 58.060 115.740 58.200 117.800 ;
        RECT 58.000 115.420 58.260 115.740 ;
        RECT 61.280 104.340 61.420 120.180 ;
        RECT 68.640 120.160 68.780 125.280 ;
        RECT 69.100 120.160 69.240 139.900 ;
        RECT 69.560 120.500 69.700 142.620 ;
        RECT 70.020 141.920 70.160 144.660 ;
        RECT 70.480 141.920 70.620 150.100 ;
        RECT 70.940 144.980 71.080 150.780 ;
        RECT 73.640 149.080 73.900 149.400 ;
        RECT 71.800 147.380 72.060 147.700 ;
        RECT 70.880 144.660 71.140 144.980 ;
        RECT 71.860 142.260 72.000 147.380 ;
        RECT 73.700 146.680 73.840 149.080 ;
        RECT 74.100 147.720 74.360 148.040 ;
        RECT 73.640 146.360 73.900 146.680 ;
        RECT 73.700 144.640 73.840 146.360 ;
        RECT 73.640 144.320 73.900 144.640 ;
        RECT 70.880 141.940 71.140 142.260 ;
        RECT 71.800 141.940 72.060 142.260 ;
        RECT 69.960 141.600 70.220 141.920 ;
        RECT 70.420 141.600 70.680 141.920 ;
        RECT 70.020 139.540 70.160 141.600 ;
        RECT 69.960 139.220 70.220 139.540 ;
        RECT 69.960 136.500 70.220 136.820 ;
        RECT 70.020 133.760 70.160 136.500 ;
        RECT 70.480 133.760 70.620 141.600 ;
        RECT 70.940 135.800 71.080 141.940 ;
        RECT 71.860 136.820 72.000 141.940 ;
        RECT 73.700 141.920 73.840 144.320 ;
        RECT 73.640 141.600 73.900 141.920 ;
        RECT 72.720 140.920 72.980 141.240 ;
        RECT 73.180 140.920 73.440 141.240 ;
        RECT 72.780 139.880 72.920 140.920 ;
        RECT 72.720 139.560 72.980 139.880 ;
        RECT 73.240 138.520 73.380 140.920 ;
        RECT 73.180 138.200 73.440 138.520 ;
        RECT 71.800 136.500 72.060 136.820 ;
        RECT 73.240 136.480 73.380 138.200 ;
        RECT 73.180 136.160 73.440 136.480 ;
        RECT 70.880 135.480 71.140 135.800 ;
        RECT 70.940 134.100 71.080 135.480 ;
        RECT 70.880 133.780 71.140 134.100 ;
        RECT 69.960 133.440 70.220 133.760 ;
        RECT 70.420 133.440 70.680 133.760 ;
        RECT 70.940 132.060 71.080 133.780 ;
        RECT 72.720 132.760 72.980 133.080 ;
        RECT 73.640 132.760 73.900 133.080 ;
        RECT 70.880 131.740 71.140 132.060 ;
        RECT 72.780 125.600 72.920 132.760 ;
        RECT 73.700 129.000 73.840 132.760 ;
        RECT 73.640 128.680 73.900 129.000 ;
        RECT 72.720 125.280 72.980 125.600 ;
        RECT 72.260 122.900 72.520 123.220 ;
        RECT 69.500 120.180 69.760 120.500 ;
        RECT 72.320 120.160 72.460 122.900 ;
        RECT 74.160 120.160 74.300 147.720 ;
        RECT 75.080 145.570 75.220 174.580 ;
        RECT 75.940 174.240 76.200 174.560 ;
        RECT 75.480 171.520 75.740 171.840 ;
        RECT 75.540 169.460 75.680 171.520 ;
        RECT 75.480 169.140 75.740 169.460 ;
        RECT 76.000 166.740 76.140 174.240 ;
        RECT 76.460 174.220 76.600 176.280 ;
        RECT 77.380 174.560 77.520 177.640 ;
        RECT 79.220 177.280 79.360 182.060 ;
        RECT 79.680 177.620 79.820 187.500 ;
        RECT 80.080 186.140 80.340 186.460 ;
        RECT 80.140 185.975 80.280 186.140 ;
        RECT 80.070 185.605 80.350 185.975 ;
        RECT 80.080 185.120 80.340 185.440 ;
        RECT 80.140 183.400 80.280 185.120 ;
        RECT 80.080 183.080 80.340 183.400 ;
        RECT 80.080 181.895 80.340 182.040 ;
        RECT 80.070 181.525 80.350 181.895 ;
        RECT 80.600 177.620 80.740 198.040 ;
        RECT 81.920 196.680 82.180 197.000 ;
        RECT 81.460 193.620 81.720 193.940 ;
        RECT 81.520 193.260 81.660 193.620 ;
        RECT 81.980 193.600 82.120 196.680 ;
        RECT 82.440 195.640 82.580 198.720 ;
        RECT 82.380 195.320 82.640 195.640 ;
        RECT 81.920 193.280 82.180 193.600 ;
        RECT 81.460 192.940 81.720 193.260 ;
        RECT 81.520 190.880 81.660 192.940 ;
        RECT 81.920 192.600 82.180 192.920 ;
        RECT 81.460 190.560 81.720 190.880 ;
        RECT 81.000 189.880 81.260 190.200 ;
        RECT 79.620 177.300 79.880 177.620 ;
        RECT 80.540 177.300 80.800 177.620 ;
        RECT 79.160 176.960 79.420 177.280 ;
        RECT 79.150 174.725 79.430 175.095 ;
        RECT 79.220 174.560 79.360 174.725 ;
        RECT 77.320 174.240 77.580 174.560 ;
        RECT 79.160 174.240 79.420 174.560 ;
        RECT 76.400 173.900 76.660 174.220 ;
        RECT 76.460 172.520 76.600 173.900 ;
        RECT 76.880 173.025 78.760 173.395 ;
        RECT 76.400 172.200 76.660 172.520 ;
        RECT 76.400 170.840 76.660 171.160 ;
        RECT 75.940 166.420 76.200 166.740 ;
        RECT 76.460 166.310 76.600 170.840 ;
        RECT 79.680 169.120 79.820 177.300 ;
        RECT 80.600 172.180 80.740 177.300 ;
        RECT 80.540 171.860 80.800 172.180 ;
        RECT 80.600 169.120 80.740 171.860 ;
        RECT 79.620 168.800 79.880 169.120 ;
        RECT 80.540 168.800 80.800 169.120 ;
        RECT 79.160 168.120 79.420 168.440 ;
        RECT 76.880 167.585 78.760 167.955 ;
        RECT 79.220 167.080 79.360 168.120 ;
        RECT 79.160 166.760 79.420 167.080 ;
        RECT 79.680 166.740 79.820 168.800 ;
        RECT 80.080 168.120 80.340 168.440 ;
        RECT 79.620 166.420 79.880 166.740 ;
        RECT 76.860 166.310 77.120 166.400 ;
        RECT 76.460 166.170 77.120 166.310 ;
        RECT 75.480 164.380 75.740 164.700 ;
        RECT 75.540 157.560 75.680 164.380 ;
        RECT 76.460 163.535 76.600 166.170 ;
        RECT 76.860 166.080 77.120 166.170 ;
        RECT 79.620 163.700 79.880 164.020 ;
        RECT 76.390 163.165 76.670 163.535 ;
        RECT 79.160 162.680 79.420 163.000 ;
        RECT 76.880 162.145 78.760 162.515 ;
        RECT 79.220 161.980 79.360 162.680 ;
        RECT 79.160 161.660 79.420 161.980 ;
        RECT 79.220 160.960 79.360 161.660 ;
        RECT 79.160 160.640 79.420 160.960 ;
        RECT 79.680 160.190 79.820 163.700 ;
        RECT 80.140 161.495 80.280 168.120 ;
        RECT 81.060 166.140 81.200 189.880 ;
        RECT 81.520 189.180 81.660 190.560 ;
        RECT 81.460 188.860 81.720 189.180 ;
        RECT 81.460 188.180 81.720 188.500 ;
        RECT 81.520 185.180 81.660 188.180 ;
        RECT 81.980 185.780 82.120 192.600 ;
        RECT 82.380 188.860 82.640 189.180 ;
        RECT 81.920 185.460 82.180 185.780 ;
        RECT 81.520 185.040 82.120 185.180 ;
        RECT 81.460 184.615 81.720 184.760 ;
        RECT 81.450 184.245 81.730 184.615 ;
        RECT 81.980 180.000 82.120 185.040 ;
        RECT 82.440 183.060 82.580 188.860 ;
        RECT 82.900 188.840 83.040 207.560 ;
        RECT 84.220 206.200 84.480 206.520 ;
        RECT 84.280 205.160 84.420 206.200 ;
        RECT 84.220 204.840 84.480 205.160 ;
        RECT 83.760 198.380 84.020 198.700 ;
        RECT 83.300 195.660 83.560 195.980 ;
        RECT 82.840 188.520 83.100 188.840 ;
        RECT 82.840 185.120 83.100 185.440 ;
        RECT 82.380 182.740 82.640 183.060 ;
        RECT 82.900 182.720 83.040 185.120 ;
        RECT 82.840 182.400 83.100 182.720 ;
        RECT 82.900 180.340 83.040 182.400 ;
        RECT 82.840 180.020 83.100 180.340 ;
        RECT 81.920 179.680 82.180 180.000 ;
        RECT 81.980 177.960 82.120 179.680 ;
        RECT 81.920 177.640 82.180 177.960 ;
        RECT 82.840 176.960 83.100 177.280 ;
        RECT 82.380 168.800 82.640 169.120 ;
        RECT 82.440 166.740 82.580 168.800 ;
        RECT 82.380 166.420 82.640 166.740 ;
        RECT 80.600 166.000 81.200 166.140 ;
        RECT 80.600 163.680 80.740 166.000 ;
        RECT 81.920 165.740 82.180 166.060 ;
        RECT 81.000 165.400 81.260 165.720 ;
        RECT 80.540 163.360 80.800 163.680 ;
        RECT 80.070 161.125 80.350 161.495 ;
        RECT 79.680 160.050 80.280 160.190 ;
        RECT 79.620 158.940 79.880 159.260 ;
        RECT 76.400 158.600 76.660 158.920 ;
        RECT 75.480 157.240 75.740 157.560 ;
        RECT 75.940 157.240 76.200 157.560 ;
        RECT 76.000 155.520 76.140 157.240 ;
        RECT 75.940 155.200 76.200 155.520 ;
        RECT 75.940 152.480 76.200 152.800 ;
        RECT 76.000 150.080 76.140 152.480 ;
        RECT 76.460 152.460 76.600 158.600 ;
        RECT 79.160 157.240 79.420 157.560 ;
        RECT 76.880 156.705 78.760 157.075 ;
        RECT 79.220 156.200 79.360 157.240 ;
        RECT 79.680 156.200 79.820 158.940 ;
        RECT 80.140 158.240 80.280 160.050 ;
        RECT 80.600 158.580 80.740 163.360 ;
        RECT 80.540 158.260 80.800 158.580 ;
        RECT 80.080 157.920 80.340 158.240 ;
        RECT 80.540 157.580 80.800 157.900 ;
        RECT 79.160 155.880 79.420 156.200 ;
        RECT 79.620 155.880 79.880 156.200 ;
        RECT 79.160 155.200 79.420 155.520 ;
        RECT 77.320 154.860 77.580 155.180 ;
        RECT 77.380 152.800 77.520 154.860 ;
        RECT 79.220 153.480 79.360 155.200 ;
        RECT 80.600 154.580 80.740 157.580 ;
        RECT 79.680 154.440 80.740 154.580 ;
        RECT 79.160 153.160 79.420 153.480 ;
        RECT 77.320 152.480 77.580 152.800 ;
        RECT 76.400 152.140 76.660 152.460 ;
        RECT 76.880 151.265 78.760 151.635 ;
        RECT 79.220 151.100 79.360 153.160 ;
        RECT 79.160 150.780 79.420 151.100 ;
        RECT 75.940 149.760 76.200 150.080 ;
        RECT 76.400 146.700 76.660 147.020 ;
        RECT 74.620 145.430 75.220 145.570 ;
        RECT 74.620 136.220 74.760 145.430 ;
        RECT 76.460 145.320 76.600 146.700 ;
        RECT 76.880 145.825 78.760 146.195 ;
        RECT 76.400 145.000 76.660 145.320 ;
        RECT 78.700 145.175 78.960 145.320 ;
        RECT 75.020 144.660 75.280 144.980 ;
        RECT 75.080 142.940 75.220 144.660 ;
        RECT 76.460 144.380 76.600 145.000 ;
        RECT 78.690 144.805 78.970 145.175 ;
        RECT 75.540 144.240 76.600 144.380 ;
        RECT 75.020 142.620 75.280 142.940 ;
        RECT 75.540 140.220 75.680 144.240 ;
        RECT 76.400 143.640 76.660 143.960 ;
        RECT 75.940 140.920 76.200 141.240 ;
        RECT 75.480 139.900 75.740 140.220 ;
        RECT 75.480 138.880 75.740 139.200 ;
        RECT 74.620 136.080 75.220 136.220 ;
        RECT 74.560 135.480 74.820 135.800 ;
        RECT 74.620 134.100 74.760 135.480 ;
        RECT 75.080 134.440 75.220 136.080 ;
        RECT 75.020 134.120 75.280 134.440 ;
        RECT 74.560 133.780 74.820 134.100 ;
        RECT 74.560 132.760 74.820 133.080 ;
        RECT 74.620 131.380 74.760 132.760 ;
        RECT 75.540 131.380 75.680 138.880 ;
        RECT 76.000 137.160 76.140 140.920 ;
        RECT 76.460 139.450 76.600 143.640 ;
        RECT 78.760 142.260 78.900 144.805 ;
        RECT 79.680 144.300 79.820 154.440 ;
        RECT 80.080 153.500 80.340 153.820 ;
        RECT 79.620 143.980 79.880 144.300 ;
        RECT 79.160 143.640 79.420 143.960 ;
        RECT 78.700 141.940 78.960 142.260 ;
        RECT 76.880 140.385 78.760 140.755 ;
        RECT 77.320 139.450 77.580 139.540 ;
        RECT 76.460 139.310 77.580 139.450 ;
        RECT 77.320 139.220 77.580 139.310 ;
        RECT 75.940 136.840 76.200 137.160 ;
        RECT 76.880 134.945 78.760 135.315 ;
        RECT 74.560 131.060 74.820 131.380 ;
        RECT 75.480 131.060 75.740 131.380 ;
        RECT 75.540 128.740 75.680 131.060 ;
        RECT 76.880 129.505 78.760 129.875 ;
        RECT 75.540 128.660 76.140 128.740 ;
        RECT 75.540 128.600 76.200 128.660 ;
        RECT 74.560 128.000 74.820 128.320 ;
        RECT 74.620 126.620 74.760 128.000 ;
        RECT 74.560 126.300 74.820 126.620 ;
        RECT 75.540 125.940 75.680 128.600 ;
        RECT 75.940 128.340 76.200 128.600 ;
        RECT 75.480 125.620 75.740 125.940 ;
        RECT 76.880 124.065 78.760 124.435 ;
        RECT 79.220 123.560 79.360 143.640 ;
        RECT 80.140 137.500 80.280 153.500 ;
        RECT 80.530 152.965 80.810 153.335 ;
        RECT 80.540 152.820 80.800 152.965 ;
        RECT 81.060 152.800 81.200 165.400 ;
        RECT 81.980 164.700 82.120 165.740 ;
        RECT 81.460 164.380 81.720 164.700 ;
        RECT 81.920 164.380 82.180 164.700 ;
        RECT 81.520 164.215 81.660 164.380 ;
        RECT 81.450 163.845 81.730 164.215 ;
        RECT 82.440 163.680 82.580 166.420 ;
        RECT 82.380 163.360 82.640 163.680 ;
        RECT 81.460 162.680 81.720 163.000 ;
        RECT 81.000 152.480 81.260 152.800 ;
        RECT 80.540 150.100 80.800 150.420 ;
        RECT 80.600 148.380 80.740 150.100 ;
        RECT 80.540 148.060 80.800 148.380 ;
        RECT 81.520 144.980 81.660 162.680 ;
        RECT 82.440 161.300 82.580 163.360 ;
        RECT 81.920 160.980 82.180 161.300 ;
        RECT 82.380 160.980 82.640 161.300 ;
        RECT 81.980 160.815 82.120 160.980 ;
        RECT 81.910 160.445 82.190 160.815 ;
        RECT 82.380 159.960 82.640 160.280 ;
        RECT 82.900 160.140 83.040 176.960 ;
        RECT 83.360 164.360 83.500 195.660 ;
        RECT 83.820 194.020 83.960 198.380 ;
        RECT 84.280 197.340 84.420 204.840 ;
        RECT 84.740 204.140 84.880 207.990 ;
        RECT 88.360 207.220 88.620 207.540 ;
        RECT 88.420 204.820 88.560 207.220 ;
        RECT 90.200 206.880 90.460 207.200 ;
        RECT 94.340 206.880 94.600 207.200 ;
        RECT 88.820 206.540 89.080 206.860 ;
        RECT 89.280 206.540 89.540 206.860 ;
        RECT 88.880 205.500 89.020 206.540 ;
        RECT 88.820 205.180 89.080 205.500 ;
        RECT 88.360 204.500 88.620 204.820 ;
        RECT 86.060 204.160 86.320 204.480 ;
        RECT 87.440 204.160 87.700 204.480 ;
        RECT 84.680 203.820 84.940 204.140 ;
        RECT 84.220 197.020 84.480 197.340 ;
        RECT 84.740 197.000 84.880 203.820 ;
        RECT 85.600 200.760 85.860 201.080 ;
        RECT 85.660 199.380 85.800 200.760 ;
        RECT 85.600 199.060 85.860 199.380 ;
        RECT 84.680 196.680 84.940 197.000 ;
        RECT 85.660 196.660 85.800 199.060 ;
        RECT 85.600 196.340 85.860 196.660 ;
        RECT 86.120 195.980 86.260 204.160 ;
        RECT 86.980 203.480 87.240 203.800 ;
        RECT 87.040 202.100 87.180 203.480 ;
        RECT 86.980 201.780 87.240 202.100 ;
        RECT 86.980 198.720 87.240 199.040 ;
        RECT 86.520 198.040 86.780 198.360 ;
        RECT 86.580 197.340 86.720 198.040 ;
        RECT 86.520 197.020 86.780 197.340 ;
        RECT 84.220 195.660 84.480 195.980 ;
        RECT 86.060 195.660 86.320 195.980 ;
        RECT 84.280 194.620 84.420 195.660 ;
        RECT 84.220 194.300 84.480 194.620 ;
        RECT 83.820 193.940 84.420 194.020 ;
        RECT 83.820 193.880 84.480 193.940 ;
        RECT 84.220 193.620 84.480 193.880 ;
        RECT 85.600 192.940 85.860 193.260 ;
        RECT 85.660 190.880 85.800 192.940 ;
        RECT 87.040 191.900 87.180 198.720 ;
        RECT 87.500 197.340 87.640 204.160 ;
        RECT 89.340 201.420 89.480 206.540 ;
        RECT 89.740 206.200 90.000 206.520 ;
        RECT 89.800 205.500 89.940 206.200 ;
        RECT 89.740 205.180 90.000 205.500 ;
        RECT 90.260 202.780 90.400 206.880 ;
        RECT 90.660 204.500 90.920 204.820 ;
        RECT 91.580 204.730 91.840 204.820 ;
        RECT 91.180 204.590 91.840 204.730 ;
        RECT 90.200 202.460 90.460 202.780 ;
        RECT 89.280 201.100 89.540 201.420 ;
        RECT 90.720 199.720 90.860 204.500 ;
        RECT 91.180 199.720 91.320 204.590 ;
        RECT 91.580 204.500 91.840 204.590 ;
        RECT 91.880 202.945 93.760 203.315 ;
        RECT 93.880 201.100 94.140 201.420 ;
        RECT 93.940 200.060 94.080 201.100 ;
        RECT 93.880 199.740 94.140 200.060 ;
        RECT 90.660 199.400 90.920 199.720 ;
        RECT 91.120 199.400 91.380 199.720 ;
        RECT 87.440 197.020 87.700 197.340 ;
        RECT 90.720 197.000 90.860 199.400 ;
        RECT 91.180 198.700 91.320 199.400 ;
        RECT 94.400 199.380 94.540 206.880 ;
        RECT 106.880 205.665 108.760 206.035 ;
        RECT 96.180 203.480 96.440 203.800 ;
        RECT 96.240 202.100 96.380 203.480 ;
        RECT 121.880 202.945 123.760 203.315 ;
        RECT 110.900 202.460 111.160 202.780 ;
        RECT 96.180 201.780 96.440 202.100 ;
        RECT 110.440 201.780 110.700 202.100 ;
        RECT 106.880 200.225 108.760 200.595 ;
        RECT 109.520 199.740 109.780 200.060 ;
        RECT 94.340 199.060 94.600 199.380 ;
        RECT 108.140 198.720 108.400 199.040 ;
        RECT 91.120 198.380 91.380 198.700 ;
        RECT 98.020 198.040 98.280 198.360 ;
        RECT 100.780 198.040 101.040 198.360 ;
        RECT 91.880 197.505 93.760 197.875 ;
        RECT 87.900 196.680 88.160 197.000 ;
        RECT 90.660 196.680 90.920 197.000 ;
        RECT 87.960 194.280 88.100 196.680 ;
        RECT 91.120 196.340 91.380 196.660 ;
        RECT 87.900 193.960 88.160 194.280 ;
        RECT 89.740 192.600 90.000 192.920 ;
        RECT 86.980 191.580 87.240 191.900 ;
        RECT 87.440 190.900 87.700 191.220 ;
        RECT 85.600 190.560 85.860 190.880 ;
        RECT 84.680 189.880 84.940 190.200 ;
        RECT 84.740 189.180 84.880 189.880 ;
        RECT 84.680 188.860 84.940 189.180 ;
        RECT 85.140 188.180 85.400 188.500 ;
        RECT 84.680 185.120 84.940 185.440 ;
        RECT 85.200 185.295 85.340 188.180 ;
        RECT 84.220 184.440 84.480 184.760 ;
        RECT 84.280 183.400 84.420 184.440 ;
        RECT 84.740 183.740 84.880 185.120 ;
        RECT 85.130 184.925 85.410 185.295 ;
        RECT 84.680 183.420 84.940 183.740 ;
        RECT 84.220 183.080 84.480 183.400 ;
        RECT 83.760 181.895 84.020 182.040 ;
        RECT 83.750 181.525 84.030 181.895 ;
        RECT 83.760 179.910 84.020 180.000 ;
        RECT 84.280 179.910 84.420 183.080 ;
        RECT 84.740 183.060 84.880 183.420 ;
        RECT 84.680 182.740 84.940 183.060 ;
        RECT 84.740 180.680 84.880 182.740 ;
        RECT 84.680 180.360 84.940 180.680 ;
        RECT 83.760 179.770 84.420 179.910 ;
        RECT 83.760 179.680 84.020 179.770 ;
        RECT 85.660 179.740 85.800 190.560 ;
        RECT 86.520 188.520 86.780 188.840 ;
        RECT 86.060 186.140 86.320 186.460 ;
        RECT 86.120 183.060 86.260 186.140 ;
        RECT 86.580 184.760 86.720 188.520 ;
        RECT 87.500 188.160 87.640 190.900 ;
        RECT 89.800 190.540 89.940 192.600 ;
        RECT 91.180 191.220 91.320 196.340 ;
        RECT 93.420 196.000 93.680 196.320 ;
        RECT 91.580 195.660 91.840 195.980 ;
        RECT 91.640 193.260 91.780 195.660 ;
        RECT 92.960 195.320 93.220 195.640 ;
        RECT 93.020 194.280 93.160 195.320 ;
        RECT 93.480 194.620 93.620 196.000 ;
        RECT 93.420 194.300 93.680 194.620 ;
        RECT 97.560 194.300 97.820 194.620 ;
        RECT 92.960 193.960 93.220 194.280 ;
        RECT 91.580 192.940 91.840 193.260 ;
        RECT 91.880 192.065 93.760 192.435 ;
        RECT 91.120 190.900 91.380 191.220 ;
        RECT 97.620 190.540 97.760 194.300 ;
        RECT 98.080 193.940 98.220 198.040 ;
        RECT 100.840 196.320 100.980 198.040 ;
        RECT 108.200 197.340 108.340 198.720 ;
        RECT 105.840 197.020 106.100 197.340 ;
        RECT 108.140 197.020 108.400 197.340 ;
        RECT 100.780 196.000 101.040 196.320 ;
        RECT 98.020 193.620 98.280 193.940 ;
        RECT 98.480 193.280 98.740 193.600 ;
        RECT 98.540 191.560 98.680 193.280 ;
        RECT 98.480 191.240 98.740 191.560 ;
        RECT 98.020 190.560 98.280 190.880 ;
        RECT 89.740 190.220 90.000 190.540 ;
        RECT 97.560 190.220 97.820 190.540 ;
        RECT 87.440 187.840 87.700 188.160 ;
        RECT 87.500 185.440 87.640 187.840 ;
        RECT 91.880 186.625 93.760 186.995 ;
        RECT 87.440 185.120 87.700 185.440 ;
        RECT 89.280 184.780 89.540 185.100 ;
        RECT 97.100 184.780 97.360 185.100 ;
        RECT 86.520 184.440 86.780 184.760 ;
        RECT 86.060 182.740 86.320 183.060 ;
        RECT 84.740 179.660 85.800 179.740 ;
        RECT 84.680 179.600 85.800 179.660 ;
        RECT 84.680 179.340 84.940 179.600 ;
        RECT 85.600 179.000 85.860 179.320 ;
        RECT 85.140 174.240 85.400 174.560 ;
        RECT 83.760 173.900 84.020 174.220 ;
        RECT 83.820 172.860 83.960 173.900 ;
        RECT 83.760 172.540 84.020 172.860 ;
        RECT 85.200 171.840 85.340 174.240 ;
        RECT 85.140 171.520 85.400 171.840 ;
        RECT 85.200 169.800 85.340 171.520 ;
        RECT 85.140 169.480 85.400 169.800 ;
        RECT 84.220 169.030 84.480 169.120 ;
        RECT 84.220 168.890 84.880 169.030 ;
        RECT 84.220 168.800 84.480 168.890 ;
        RECT 83.760 168.120 84.020 168.440 ;
        RECT 83.300 164.040 83.560 164.360 ;
        RECT 82.900 160.000 83.500 160.140 ;
        RECT 81.910 145.485 82.190 145.855 ;
        RECT 81.460 144.660 81.720 144.980 ;
        RECT 81.980 144.640 82.120 145.485 ;
        RECT 81.920 144.320 82.180 144.640 ;
        RECT 81.460 143.980 81.720 144.300 ;
        RECT 81.520 142.260 81.660 143.980 ;
        RECT 81.460 141.940 81.720 142.260 ;
        RECT 80.540 141.260 80.800 141.580 ;
        RECT 80.600 139.880 80.740 141.260 ;
        RECT 80.540 139.560 80.800 139.880 ;
        RECT 80.080 137.180 80.340 137.500 ;
        RECT 81.000 132.760 81.260 133.080 ;
        RECT 81.060 130.700 81.200 132.760 ;
        RECT 81.000 130.380 81.260 130.700 ;
        RECT 80.080 130.040 80.340 130.360 ;
        RECT 80.140 125.600 80.280 130.040 ;
        RECT 80.080 125.280 80.340 125.600 ;
        RECT 81.520 123.900 81.660 141.940 ;
        RECT 82.440 141.920 82.580 159.960 ;
        RECT 83.360 158.240 83.500 160.000 ;
        RECT 83.820 158.240 83.960 168.120 ;
        RECT 84.740 165.720 84.880 168.890 ;
        RECT 85.140 166.420 85.400 166.740 ;
        RECT 84.680 165.400 84.940 165.720 ;
        RECT 84.740 164.360 84.880 165.400 ;
        RECT 84.210 163.845 84.490 164.215 ;
        RECT 84.680 164.040 84.940 164.360 ;
        RECT 84.280 160.620 84.420 163.845 ;
        RECT 84.740 161.300 84.880 164.040 ;
        RECT 85.200 161.300 85.340 166.420 ;
        RECT 84.680 160.980 84.940 161.300 ;
        RECT 85.140 160.980 85.400 161.300 ;
        RECT 84.220 160.300 84.480 160.620 ;
        RECT 85.660 158.580 85.800 179.000 ;
        RECT 86.120 177.620 86.260 182.740 ;
        RECT 86.580 178.300 86.720 184.440 ;
        RECT 89.340 183.740 89.480 184.780 ;
        RECT 90.200 184.440 90.460 184.760 ;
        RECT 89.280 183.420 89.540 183.740 ;
        RECT 87.440 182.740 87.700 183.060 ;
        RECT 87.500 181.020 87.640 182.740 ;
        RECT 87.440 180.700 87.700 181.020 ;
        RECT 87.500 180.340 87.640 180.700 ;
        RECT 87.440 180.020 87.700 180.340 ;
        RECT 89.740 179.340 90.000 179.660 ;
        RECT 86.980 179.000 87.240 179.320 ;
        RECT 86.520 177.980 86.780 178.300 ;
        RECT 86.060 177.300 86.320 177.620 ;
        RECT 87.040 175.580 87.180 179.000 ;
        RECT 89.800 178.300 89.940 179.340 ;
        RECT 89.740 177.980 90.000 178.300 ;
        RECT 90.260 177.620 90.400 184.440 ;
        RECT 91.880 181.185 93.760 181.555 ;
        RECT 94.340 180.020 94.600 180.340 ;
        RECT 94.400 178.300 94.540 180.020 ;
        RECT 96.180 179.000 96.440 179.320 ;
        RECT 94.340 177.980 94.600 178.300 ;
        RECT 96.240 177.960 96.380 179.000 ;
        RECT 95.720 177.640 95.980 177.960 ;
        RECT 96.180 177.640 96.440 177.960 ;
        RECT 90.200 177.300 90.460 177.620 ;
        RECT 88.360 176.960 88.620 177.280 ;
        RECT 86.060 175.260 86.320 175.580 ;
        RECT 86.980 175.260 87.240 175.580 ;
        RECT 86.120 172.860 86.260 175.260 ;
        RECT 86.520 173.560 86.780 173.880 ;
        RECT 86.060 172.540 86.320 172.860 ;
        RECT 86.120 169.460 86.260 172.540 ;
        RECT 86.580 172.180 86.720 173.560 ;
        RECT 88.420 172.860 88.560 176.960 ;
        RECT 91.880 175.745 93.760 176.115 ;
        RECT 90.200 174.580 90.460 174.900 ;
        RECT 91.120 174.580 91.380 174.900 ;
        RECT 90.260 173.880 90.400 174.580 ;
        RECT 90.200 173.560 90.460 173.880 ;
        RECT 88.360 172.540 88.620 172.860 ;
        RECT 90.190 172.685 90.470 173.055 ;
        RECT 90.260 172.520 90.400 172.685 ;
        RECT 90.200 172.200 90.460 172.520 ;
        RECT 86.520 171.860 86.780 172.180 ;
        RECT 87.440 171.860 87.700 172.180 ;
        RECT 86.060 169.140 86.320 169.460 ;
        RECT 86.980 169.140 87.240 169.460 ;
        RECT 86.520 168.800 86.780 169.120 ;
        RECT 86.060 168.120 86.320 168.440 ;
        RECT 86.120 167.420 86.260 168.120 ;
        RECT 86.060 167.100 86.320 167.420 ;
        RECT 86.120 164.020 86.260 167.100 ;
        RECT 86.580 166.060 86.720 168.800 ;
        RECT 87.040 166.400 87.180 169.140 ;
        RECT 87.500 168.780 87.640 171.860 ;
        RECT 91.180 170.140 91.320 174.580 ;
        RECT 95.780 174.560 95.920 177.640 ;
        RECT 97.160 177.620 97.300 184.780 ;
        RECT 97.620 180.680 97.760 190.220 ;
        RECT 98.080 189.180 98.220 190.560 ;
        RECT 98.020 188.860 98.280 189.180 ;
        RECT 98.540 188.840 98.680 191.240 ;
        RECT 98.940 189.880 99.200 190.200 ;
        RECT 99.000 188.840 99.140 189.880 ;
        RECT 98.480 188.520 98.740 188.840 ;
        RECT 98.940 188.520 99.200 188.840 ;
        RECT 98.540 185.780 98.680 188.520 ;
        RECT 99.860 187.160 100.120 187.480 ;
        RECT 99.920 185.780 100.060 187.160 ;
        RECT 98.480 185.460 98.740 185.780 ;
        RECT 99.860 185.460 100.120 185.780 ;
        RECT 98.540 183.060 98.680 185.460 ;
        RECT 100.320 185.120 100.580 185.440 ;
        RECT 100.380 183.740 100.520 185.120 ;
        RECT 100.320 183.420 100.580 183.740 ;
        RECT 100.840 183.400 100.980 196.000 ;
        RECT 104.920 192.600 105.180 192.920 ;
        RECT 104.980 190.540 105.120 192.600 ;
        RECT 104.920 190.220 105.180 190.540 ;
        RECT 105.900 187.900 106.040 197.020 ;
        RECT 109.060 196.000 109.320 196.320 ;
        RECT 106.880 194.785 108.760 195.155 ;
        RECT 109.120 194.620 109.260 196.000 ;
        RECT 109.060 194.300 109.320 194.620 ;
        RECT 106.300 193.620 106.560 193.940 ;
        RECT 106.360 189.180 106.500 193.620 ;
        RECT 109.580 193.340 109.720 199.740 ;
        RECT 109.980 198.720 110.240 199.040 ;
        RECT 110.040 196.660 110.180 198.720 ;
        RECT 109.980 196.340 110.240 196.660 ;
        RECT 109.980 195.320 110.240 195.640 ;
        RECT 109.120 193.200 109.720 193.340 ;
        RECT 106.880 189.345 108.760 189.715 ;
        RECT 106.300 188.860 106.560 189.180 ;
        RECT 109.120 188.840 109.260 193.200 ;
        RECT 109.520 192.600 109.780 192.920 ;
        RECT 109.580 189.180 109.720 192.600 ;
        RECT 110.040 191.220 110.180 195.320 ;
        RECT 109.980 190.900 110.240 191.220 ;
        RECT 109.520 188.860 109.780 189.180 ;
        RECT 109.060 188.520 109.320 188.840 ;
        RECT 109.980 188.520 110.240 188.840 ;
        RECT 106.300 187.900 106.560 188.160 ;
        RECT 105.900 187.840 106.560 187.900 ;
        RECT 105.900 187.760 106.500 187.840 ;
        RECT 101.240 187.160 101.500 187.480 ;
        RECT 101.300 186.460 101.440 187.160 ;
        RECT 105.900 186.540 106.040 187.760 ;
        RECT 101.240 186.140 101.500 186.460 ;
        RECT 105.440 186.400 106.040 186.540 ;
        RECT 105.440 185.780 105.580 186.400 ;
        RECT 105.840 185.800 106.100 186.120 ;
        RECT 106.300 185.800 106.560 186.120 ;
        RECT 105.380 185.460 105.640 185.780 ;
        RECT 102.160 184.440 102.420 184.760 ;
        RECT 100.780 183.080 101.040 183.400 ;
        RECT 102.220 183.060 102.360 184.440 ;
        RECT 105.900 183.820 106.040 185.800 ;
        RECT 105.440 183.740 106.040 183.820 ;
        RECT 105.440 183.680 106.100 183.740 ;
        RECT 105.440 183.060 105.580 183.680 ;
        RECT 105.840 183.420 106.100 183.680 ;
        RECT 106.360 183.060 106.500 185.800 ;
        RECT 109.060 185.120 109.320 185.440 ;
        RECT 106.880 183.905 108.760 184.275 ;
        RECT 109.120 183.740 109.260 185.120 ;
        RECT 109.520 184.780 109.780 185.100 ;
        RECT 109.060 183.420 109.320 183.740 ;
        RECT 109.120 183.060 109.260 183.420 ;
        RECT 109.580 183.060 109.720 184.780 ;
        RECT 110.040 183.740 110.180 188.520 ;
        RECT 109.980 183.420 110.240 183.740 ;
        RECT 98.480 182.740 98.740 183.060 ;
        RECT 102.160 182.740 102.420 183.060 ;
        RECT 105.380 182.740 105.640 183.060 ;
        RECT 105.840 182.740 106.100 183.060 ;
        RECT 106.300 182.740 106.560 183.060 ;
        RECT 106.760 182.740 107.020 183.060 ;
        RECT 109.060 182.740 109.320 183.060 ;
        RECT 109.520 182.740 109.780 183.060 ;
        RECT 98.540 181.020 98.680 182.740 ;
        RECT 103.080 181.720 103.340 182.040 ;
        RECT 98.480 180.700 98.740 181.020 ;
        RECT 97.560 180.360 97.820 180.680 ;
        RECT 97.560 179.680 97.820 180.000 ;
        RECT 102.160 179.680 102.420 180.000 ;
        RECT 97.100 177.300 97.360 177.620 ;
        RECT 97.620 176.600 97.760 179.680 ;
        RECT 101.240 179.000 101.500 179.320 ;
        RECT 100.780 178.210 101.040 178.300 ;
        RECT 101.300 178.210 101.440 179.000 ;
        RECT 100.780 178.070 101.440 178.210 ;
        RECT 100.780 177.980 101.040 178.070 ;
        RECT 97.560 176.280 97.820 176.600 ;
        RECT 95.720 174.240 95.980 174.560 ;
        RECT 95.780 171.840 95.920 174.240 ;
        RECT 95.720 171.520 95.980 171.840 ;
        RECT 91.880 170.305 93.760 170.675 ;
        RECT 91.120 169.820 91.380 170.140 ;
        RECT 87.440 168.460 87.700 168.780 ;
        RECT 87.500 167.080 87.640 168.460 ;
        RECT 87.440 166.760 87.700 167.080 ;
        RECT 95.780 166.400 95.920 171.520 ;
        RECT 96.180 168.120 96.440 168.440 ;
        RECT 86.980 166.080 87.240 166.400 ;
        RECT 86.520 165.740 86.780 166.060 ;
        RECT 93.020 166.000 94.080 166.140 ;
        RECT 95.720 166.080 95.980 166.400 ;
        RECT 96.240 166.060 96.380 168.120 ;
        RECT 97.100 166.760 97.360 167.080 ;
        RECT 96.640 166.080 96.900 166.400 ;
        RECT 86.060 163.700 86.320 164.020 ;
        RECT 86.580 163.420 86.720 165.740 ;
        RECT 93.020 165.720 93.160 166.000 ;
        RECT 91.120 165.400 91.380 165.720 ;
        RECT 92.960 165.400 93.220 165.720 ;
        RECT 86.120 163.340 86.720 163.420 ;
        RECT 91.180 163.340 91.320 165.400 ;
        RECT 91.880 164.865 93.760 165.235 ;
        RECT 93.940 164.020 94.080 166.000 ;
        RECT 96.180 165.740 96.440 166.060 ;
        RECT 94.340 165.400 94.600 165.720 ;
        RECT 93.880 163.700 94.140 164.020 ;
        RECT 86.060 163.280 86.720 163.340 ;
        RECT 86.060 163.020 86.320 163.280 ;
        RECT 91.120 163.020 91.380 163.340 ;
        RECT 86.120 161.300 86.260 163.020 ;
        RECT 94.400 161.300 94.540 165.400 ;
        RECT 96.700 163.680 96.840 166.080 ;
        RECT 97.160 164.700 97.300 166.760 ;
        RECT 97.100 164.380 97.360 164.700 ;
        RECT 97.620 164.360 97.760 176.280 ;
        RECT 101.300 174.900 101.440 178.070 ;
        RECT 102.220 175.580 102.360 179.680 ;
        RECT 102.160 175.260 102.420 175.580 ;
        RECT 101.700 174.920 101.960 175.240 ;
        RECT 98.020 174.580 98.280 174.900 ;
        RECT 101.240 174.580 101.500 174.900 ;
        RECT 98.080 169.460 98.220 174.580 ;
        RECT 99.400 173.900 99.660 174.220 ;
        RECT 99.460 172.860 99.600 173.900 ;
        RECT 99.400 172.540 99.660 172.860 ;
        RECT 101.760 172.520 101.900 174.920 ;
        RECT 102.620 172.540 102.880 172.860 ;
        RECT 101.700 172.200 101.960 172.520 ;
        RECT 98.940 170.840 99.200 171.160 ;
        RECT 98.020 169.140 98.280 169.460 ;
        RECT 99.000 169.120 99.140 170.840 ;
        RECT 98.940 168.800 99.200 169.120 ;
        RECT 99.000 168.440 99.140 168.800 ;
        RECT 98.940 168.120 99.200 168.440 ;
        RECT 97.560 164.040 97.820 164.360 ;
        RECT 99.000 163.680 99.140 168.120 ;
        RECT 102.680 166.740 102.820 172.540 ;
        RECT 102.620 166.420 102.880 166.740 ;
        RECT 102.680 164.020 102.820 166.420 ;
        RECT 102.620 163.700 102.880 164.020 ;
        RECT 96.640 163.360 96.900 163.680 ;
        RECT 97.560 163.360 97.820 163.680 ;
        RECT 98.020 163.360 98.280 163.680 ;
        RECT 98.940 163.360 99.200 163.680 ;
        RECT 99.400 163.360 99.660 163.680 ;
        RECT 96.180 161.660 96.440 161.980 ;
        RECT 86.060 160.980 86.320 161.300 ;
        RECT 94.340 160.980 94.600 161.300 ;
        RECT 93.880 159.960 94.140 160.280 ;
        RECT 91.880 159.425 93.760 159.795 ;
        RECT 86.520 158.940 86.780 159.260 ;
        RECT 85.600 158.260 85.860 158.580 ;
        RECT 83.300 157.920 83.560 158.240 ;
        RECT 83.760 157.920 84.020 158.240 ;
        RECT 85.140 157.580 85.400 157.900 ;
        RECT 85.200 156.540 85.340 157.580 ;
        RECT 85.600 157.240 85.860 157.560 ;
        RECT 82.840 156.450 83.100 156.540 ;
        RECT 83.760 156.450 84.020 156.540 ;
        RECT 82.840 156.310 84.020 156.450 ;
        RECT 82.840 156.220 83.100 156.310 ;
        RECT 83.760 156.220 84.020 156.310 ;
        RECT 85.140 156.220 85.400 156.540 ;
        RECT 83.760 155.540 84.020 155.860 ;
        RECT 85.140 155.540 85.400 155.860 ;
        RECT 83.300 155.430 83.560 155.520 ;
        RECT 82.900 155.290 83.560 155.430 ;
        RECT 82.900 153.140 83.040 155.290 ;
        RECT 83.300 155.200 83.560 155.290 ;
        RECT 83.820 155.180 83.960 155.540 ;
        RECT 83.760 154.860 84.020 155.180 ;
        RECT 83.300 153.160 83.560 153.480 ;
        RECT 82.840 152.820 83.100 153.140 ;
        RECT 82.900 144.980 83.040 152.820 ;
        RECT 83.360 152.460 83.500 153.160 ;
        RECT 83.820 152.800 83.960 154.860 ;
        RECT 85.200 152.800 85.340 155.540 ;
        RECT 83.760 152.480 84.020 152.800 ;
        RECT 85.140 152.480 85.400 152.800 ;
        RECT 83.300 152.140 83.560 152.460 ;
        RECT 82.840 144.660 83.100 144.980 ;
        RECT 83.360 144.890 83.500 152.140 ;
        RECT 83.820 145.660 83.960 152.480 ;
        RECT 84.680 151.800 84.940 152.120 ;
        RECT 83.760 145.340 84.020 145.660 ;
        RECT 84.220 144.890 84.480 144.980 ;
        RECT 83.360 144.750 84.480 144.890 ;
        RECT 84.220 144.660 84.480 144.750 ;
        RECT 82.900 144.495 83.040 144.660 ;
        RECT 82.830 144.125 83.110 144.495 ;
        RECT 83.300 143.980 83.560 144.300 ;
        RECT 82.840 143.640 83.100 143.960 ;
        RECT 82.380 141.600 82.640 141.920 ;
        RECT 82.900 137.500 83.040 143.640 ;
        RECT 83.360 142.940 83.500 143.980 ;
        RECT 83.300 142.620 83.560 142.940 ;
        RECT 83.760 142.620 84.020 142.940 ;
        RECT 83.290 142.085 83.570 142.455 ;
        RECT 83.300 141.940 83.560 142.085 ;
        RECT 83.300 138.200 83.560 138.520 ;
        RECT 82.840 137.180 83.100 137.500 ;
        RECT 83.360 137.160 83.500 138.200 ;
        RECT 83.820 137.500 83.960 142.620 ;
        RECT 84.280 142.260 84.420 144.660 ;
        RECT 84.220 141.940 84.480 142.260 ;
        RECT 83.760 137.180 84.020 137.500 ;
        RECT 83.300 136.840 83.560 137.160 ;
        RECT 81.920 136.160 82.180 136.480 ;
        RECT 81.980 134.780 82.120 136.160 ;
        RECT 81.920 134.460 82.180 134.780 ;
        RECT 81.980 129.340 82.120 134.460 ;
        RECT 83.360 133.760 83.500 136.840 ;
        RECT 84.220 136.160 84.480 136.480 ;
        RECT 83.760 134.010 84.020 134.100 ;
        RECT 84.280 134.010 84.420 136.160 ;
        RECT 83.760 133.870 84.420 134.010 ;
        RECT 83.760 133.780 84.020 133.870 ;
        RECT 83.300 133.440 83.560 133.760 ;
        RECT 82.380 132.760 82.640 133.080 ;
        RECT 81.920 129.020 82.180 129.340 ;
        RECT 82.440 129.000 82.580 132.760 ;
        RECT 83.360 132.060 83.500 133.440 ;
        RECT 83.300 131.740 83.560 132.060 ;
        RECT 83.820 131.380 83.960 133.780 ;
        RECT 83.760 131.060 84.020 131.380 ;
        RECT 82.380 128.680 82.640 129.000 ;
        RECT 81.460 123.580 81.720 123.900 ;
        RECT 79.160 123.240 79.420 123.560 ;
        RECT 84.740 120.500 84.880 151.800 ;
        RECT 85.200 151.100 85.340 152.480 ;
        RECT 85.140 150.780 85.400 151.100 ;
        RECT 85.140 122.900 85.400 123.220 ;
        RECT 84.680 120.180 84.940 120.500 ;
        RECT 68.580 119.840 68.840 120.160 ;
        RECT 69.040 119.840 69.300 120.160 ;
        RECT 72.260 119.840 72.520 120.160 ;
        RECT 74.100 119.840 74.360 120.160 ;
        RECT 63.980 119.500 64.240 119.820 ;
        RECT 61.880 115.905 63.760 116.275 ;
        RECT 64.040 115.740 64.180 119.500 ;
        RECT 66.280 119.160 66.540 119.480 ;
        RECT 64.440 117.800 64.700 118.120 ;
        RECT 64.500 115.740 64.640 117.800 ;
        RECT 65.820 117.460 66.080 117.780 ;
        RECT 63.980 115.420 64.240 115.740 ;
        RECT 64.440 115.420 64.700 115.740 ;
        RECT 65.880 111.840 66.020 117.460 ;
        RECT 66.340 114.720 66.480 119.160 ;
        RECT 68.640 117.440 68.780 119.840 ;
        RECT 70.420 119.500 70.680 119.820 ;
        RECT 81.460 119.500 81.720 119.820 ;
        RECT 84.680 119.500 84.940 119.820 ;
        RECT 68.580 117.120 68.840 117.440 ;
        RECT 66.280 114.400 66.540 114.720 ;
        RECT 70.480 114.380 70.620 119.500 ;
        RECT 70.880 119.160 71.140 119.480 ;
        RECT 73.640 119.160 73.900 119.480 ;
        RECT 74.100 119.160 74.360 119.480 ;
        RECT 70.940 118.120 71.080 119.160 ;
        RECT 73.700 118.120 73.840 119.160 ;
        RECT 70.880 117.800 71.140 118.120 ;
        RECT 73.640 117.800 73.900 118.120 ;
        RECT 74.160 115.060 74.300 119.160 ;
        RECT 76.880 118.625 78.760 118.995 ;
        RECT 76.400 117.460 76.660 117.780 ;
        RECT 75.480 117.120 75.740 117.440 ;
        RECT 75.540 115.060 75.680 117.120 ;
        RECT 71.340 114.740 71.600 115.060 ;
        RECT 74.100 114.740 74.360 115.060 ;
        RECT 75.480 114.740 75.740 115.060 ;
        RECT 70.420 114.060 70.680 114.380 ;
        RECT 65.880 111.700 66.480 111.840 ;
        RECT 66.340 104.340 66.480 111.700 ;
        RECT 71.400 104.340 71.540 114.740 ;
        RECT 76.460 104.340 76.600 117.460 ;
        RECT 76.880 113.185 78.760 113.555 ;
        RECT 81.520 104.340 81.660 119.500 ;
        RECT 82.840 119.160 83.100 119.480 ;
        RECT 82.900 118.120 83.040 119.160 ;
        RECT 84.740 118.120 84.880 119.500 ;
        RECT 82.840 117.800 83.100 118.120 ;
        RECT 84.680 117.800 84.940 118.120 ;
        RECT 85.200 116.760 85.340 122.900 ;
        RECT 85.660 117.780 85.800 157.240 ;
        RECT 86.060 150.100 86.320 150.420 ;
        RECT 86.120 146.680 86.260 150.100 ;
        RECT 86.060 146.360 86.320 146.680 ;
        RECT 86.120 145.320 86.260 146.360 ;
        RECT 86.060 145.000 86.320 145.320 ;
        RECT 86.060 143.980 86.320 144.300 ;
        RECT 86.120 141.920 86.260 143.980 ;
        RECT 86.060 141.600 86.320 141.920 ;
        RECT 86.060 139.220 86.320 139.540 ;
        RECT 86.120 136.480 86.260 139.220 ;
        RECT 86.580 139.200 86.720 158.940 ;
        RECT 93.940 158.830 94.080 159.960 ;
        RECT 93.480 158.690 94.080 158.830 ;
        RECT 93.480 157.900 93.620 158.690 ;
        RECT 93.420 157.580 93.680 157.900 ;
        RECT 87.900 157.240 88.160 157.560 ;
        RECT 87.960 156.200 88.100 157.240 ;
        RECT 87.900 155.880 88.160 156.200 ;
        RECT 92.040 155.770 92.300 155.860 ;
        RECT 94.400 155.770 94.540 160.980 ;
        RECT 96.240 160.135 96.380 161.660 ;
        RECT 96.170 159.765 96.450 160.135 ;
        RECT 96.640 159.960 96.900 160.280 ;
        RECT 95.260 157.920 95.520 158.240 ;
        RECT 95.720 157.920 95.980 158.240 ;
        RECT 95.320 156.540 95.460 157.920 ;
        RECT 95.260 156.220 95.520 156.540 ;
        RECT 92.040 155.630 94.540 155.770 ;
        RECT 92.040 155.540 92.300 155.630 ;
        RECT 86.980 155.200 87.240 155.520 ;
        RECT 87.040 154.840 87.180 155.200 ;
        RECT 86.980 154.520 87.240 154.840 ;
        RECT 90.660 154.520 90.920 154.840 ;
        RECT 87.040 150.080 87.180 154.520 ;
        RECT 90.720 152.460 90.860 154.520 ;
        RECT 91.880 153.985 93.760 154.355 ;
        RECT 93.420 152.480 93.680 152.800 ;
        RECT 90.660 152.140 90.920 152.460 ;
        RECT 93.480 151.100 93.620 152.480 ;
        RECT 93.420 150.780 93.680 151.100 ;
        RECT 86.980 149.760 87.240 150.080 ;
        RECT 87.040 144.640 87.180 149.760 ;
        RECT 91.880 148.545 93.760 148.915 ;
        RECT 89.740 147.380 90.000 147.700 ;
        RECT 86.980 144.320 87.240 144.640 ;
        RECT 88.360 143.640 88.620 143.960 ;
        RECT 88.420 141.920 88.560 143.640 ;
        RECT 89.800 142.940 89.940 147.380 ;
        RECT 94.400 147.360 94.540 155.630 ;
        RECT 95.780 152.800 95.920 157.920 ;
        RECT 96.700 157.560 96.840 159.960 ;
        RECT 97.620 158.240 97.760 163.360 ;
        RECT 98.080 160.960 98.220 163.360 ;
        RECT 99.460 161.495 99.600 163.360 ;
        RECT 100.320 162.680 100.580 163.000 ;
        RECT 98.480 160.980 98.740 161.300 ;
        RECT 99.390 161.125 99.670 161.495 ;
        RECT 98.020 160.640 98.280 160.960 ;
        RECT 98.540 159.260 98.680 160.980 ;
        RECT 98.940 160.300 99.200 160.620 ;
        RECT 98.480 158.940 98.740 159.260 ;
        RECT 97.560 157.920 97.820 158.240 ;
        RECT 96.640 157.240 96.900 157.560 ;
        RECT 96.700 155.860 96.840 157.240 ;
        RECT 96.640 155.540 96.900 155.860 ;
        RECT 97.620 155.180 97.760 157.920 ;
        RECT 97.560 154.860 97.820 155.180 ;
        RECT 99.000 153.140 99.140 160.300 ;
        RECT 98.940 152.820 99.200 153.140 ;
        RECT 95.720 152.480 95.980 152.800 ;
        RECT 99.400 152.480 99.660 152.800 ;
        RECT 95.780 147.700 95.920 152.480 ;
        RECT 98.480 152.140 98.740 152.460 ;
        RECT 98.020 151.800 98.280 152.120 ;
        RECT 95.720 147.380 95.980 147.700 ;
        RECT 98.080 147.360 98.220 151.800 ;
        RECT 98.540 149.400 98.680 152.140 ;
        RECT 99.460 152.120 99.600 152.480 ;
        RECT 99.400 151.800 99.660 152.120 ;
        RECT 99.400 150.440 99.660 150.760 ;
        RECT 98.480 149.080 98.740 149.400 ;
        RECT 94.340 147.270 94.600 147.360 ;
        RECT 94.340 147.130 95.000 147.270 ;
        RECT 94.340 147.040 94.600 147.130 ;
        RECT 91.120 146.700 91.380 147.020 ;
        RECT 90.660 144.320 90.920 144.640 ;
        RECT 89.740 142.620 90.000 142.940 ;
        RECT 90.720 142.260 90.860 144.320 ;
        RECT 91.180 142.940 91.320 146.700 ;
        RECT 93.880 144.660 94.140 144.980 ;
        RECT 91.880 143.105 93.760 143.475 ;
        RECT 91.120 142.620 91.380 142.940 ;
        RECT 90.660 141.940 90.920 142.260 ;
        RECT 88.360 141.600 88.620 141.920 ;
        RECT 93.940 139.735 94.080 144.660 ;
        RECT 94.340 143.640 94.600 143.960 ;
        RECT 87.890 139.365 88.170 139.735 ;
        RECT 86.520 138.880 86.780 139.200 ;
        RECT 87.960 136.480 88.100 139.365 ;
        RECT 93.420 139.220 93.680 139.540 ;
        RECT 93.870 139.365 94.150 139.735 ;
        RECT 94.400 139.540 94.540 143.640 ;
        RECT 94.860 142.940 95.000 147.130 ;
        RECT 98.020 147.040 98.280 147.360 ;
        RECT 98.540 147.020 98.680 149.080 ;
        RECT 99.460 148.380 99.600 150.440 ;
        RECT 99.400 148.060 99.660 148.380 ;
        RECT 99.860 148.060 100.120 148.380 ;
        RECT 98.480 146.700 98.740 147.020 ;
        RECT 98.540 145.660 98.680 146.700 ;
        RECT 98.480 145.340 98.740 145.660 ;
        RECT 94.800 142.850 95.060 142.940 ;
        RECT 94.800 142.710 95.460 142.850 ;
        RECT 94.800 142.620 95.060 142.710 ;
        RECT 94.800 141.940 95.060 142.260 ;
        RECT 94.860 140.220 95.000 141.940 ;
        RECT 94.800 139.900 95.060 140.220 ;
        RECT 95.320 139.540 95.460 142.710 ;
        RECT 96.180 141.260 96.440 141.580 ;
        RECT 96.240 140.220 96.380 141.260 ;
        RECT 99.400 140.920 99.660 141.240 ;
        RECT 96.180 139.900 96.440 140.220 ;
        RECT 96.640 139.560 96.900 139.880 ;
        RECT 94.340 139.220 94.600 139.540 ;
        RECT 95.260 139.220 95.520 139.540 ;
        RECT 90.660 138.880 90.920 139.200 ;
        RECT 93.480 138.940 93.620 139.220 ;
        RECT 86.060 136.160 86.320 136.480 ;
        RECT 86.520 136.160 86.780 136.480 ;
        RECT 87.900 136.335 88.160 136.480 ;
        RECT 86.580 132.060 86.720 136.160 ;
        RECT 87.890 135.965 88.170 136.335 ;
        RECT 90.720 134.100 90.860 138.880 ;
        RECT 93.480 138.800 94.080 138.940 ;
        RECT 91.880 137.665 93.760 138.035 ;
        RECT 93.940 134.780 94.080 138.800 ;
        RECT 95.320 137.500 95.460 139.220 ;
        RECT 95.260 137.180 95.520 137.500 ;
        RECT 95.260 135.480 95.520 135.800 ;
        RECT 93.880 134.460 94.140 134.780 ;
        RECT 95.320 134.100 95.460 135.480 ;
        RECT 88.820 133.780 89.080 134.100 ;
        RECT 90.660 133.780 90.920 134.100 ;
        RECT 95.260 133.780 95.520 134.100 ;
        RECT 86.520 131.740 86.780 132.060 ;
        RECT 88.360 130.720 88.620 131.040 ;
        RECT 88.420 126.620 88.560 130.720 ;
        RECT 88.360 126.300 88.620 126.620 ;
        RECT 88.880 125.940 89.020 133.780 ;
        RECT 89.280 130.720 89.540 131.040 ;
        RECT 89.340 128.320 89.480 130.720 ;
        RECT 90.720 130.360 90.860 133.780 ;
        RECT 93.880 133.100 94.140 133.420 ;
        RECT 91.120 132.760 91.380 133.080 ;
        RECT 91.180 131.040 91.320 132.760 ;
        RECT 91.880 132.225 93.760 132.595 ;
        RECT 91.120 130.720 91.380 131.040 ;
        RECT 90.200 130.040 90.460 130.360 ;
        RECT 90.660 130.040 90.920 130.360 ;
        RECT 90.260 128.660 90.400 130.040 ;
        RECT 90.720 129.340 90.860 130.040 ;
        RECT 90.660 129.020 90.920 129.340 ;
        RECT 93.940 129.000 94.080 133.100 ;
        RECT 95.320 131.380 95.460 133.780 ;
        RECT 95.260 131.060 95.520 131.380 ;
        RECT 93.880 128.680 94.140 129.000 ;
        RECT 90.200 128.340 90.460 128.660 ;
        RECT 95.320 128.320 95.460 131.060 ;
        RECT 95.720 130.380 95.980 130.700 ;
        RECT 89.280 128.000 89.540 128.320 ;
        RECT 95.260 128.000 95.520 128.320 ;
        RECT 88.820 125.620 89.080 125.940 ;
        RECT 89.340 120.160 89.480 128.000 ;
        RECT 91.880 126.785 93.760 127.155 ;
        RECT 95.780 125.600 95.920 130.380 ;
        RECT 96.700 128.660 96.840 139.560 ;
        RECT 98.940 138.200 99.200 138.520 ;
        RECT 99.000 135.800 99.140 138.200 ;
        RECT 98.940 135.480 99.200 135.800 ;
        RECT 99.000 134.780 99.140 135.480 ;
        RECT 98.940 134.460 99.200 134.780 ;
        RECT 99.460 134.180 99.600 140.920 ;
        RECT 99.920 139.200 100.060 148.060 ;
        RECT 100.380 147.360 100.520 162.680 ;
        RECT 102.680 161.640 102.820 163.700 ;
        RECT 102.620 161.320 102.880 161.640 ;
        RECT 102.160 149.760 102.420 150.080 ;
        RECT 102.220 148.040 102.360 149.760 ;
        RECT 102.160 147.720 102.420 148.040 ;
        RECT 100.320 147.040 100.580 147.360 ;
        RECT 102.220 145.320 102.360 147.720 ;
        RECT 103.140 147.700 103.280 181.720 ;
        RECT 104.460 180.020 104.720 180.340 ;
        RECT 104.000 179.000 104.260 179.320 ;
        RECT 104.060 177.960 104.200 179.000 ;
        RECT 104.520 177.960 104.660 180.020 ;
        RECT 105.900 179.320 106.040 182.740 ;
        RECT 106.820 181.020 106.960 182.740 ;
        RECT 109.120 182.380 109.260 182.740 ;
        RECT 109.060 182.060 109.320 182.380 ;
        RECT 106.760 180.700 107.020 181.020 ;
        RECT 106.300 179.910 106.560 180.000 ;
        RECT 106.820 179.910 106.960 180.700 ;
        RECT 109.120 180.000 109.260 182.060 ;
        RECT 110.500 180.340 110.640 201.780 ;
        RECT 110.960 201.760 111.100 202.460 ;
        RECT 112.280 202.120 112.540 202.440 ;
        RECT 110.900 201.440 111.160 201.760 ;
        RECT 110.960 199.380 111.100 201.440 ;
        RECT 112.340 199.380 112.480 202.120 ;
        RECT 114.120 201.780 114.380 202.100 ;
        RECT 110.900 199.060 111.160 199.380 ;
        RECT 112.280 199.060 112.540 199.380 ;
        RECT 110.960 193.600 111.100 199.060 ;
        RECT 111.820 198.720 112.080 199.040 ;
        RECT 111.880 194.280 112.020 198.720 ;
        RECT 112.340 196.660 112.480 199.060 ;
        RECT 112.280 196.340 112.540 196.660 ;
        RECT 112.280 195.660 112.540 195.980 ;
        RECT 111.820 193.960 112.080 194.280 ;
        RECT 110.900 193.280 111.160 193.600 ;
        RECT 110.960 191.130 111.100 193.280 ;
        RECT 111.360 191.130 111.620 191.220 ;
        RECT 110.960 190.990 111.620 191.130 ;
        RECT 110.960 188.500 111.100 190.990 ;
        RECT 111.360 190.900 111.620 190.990 ;
        RECT 111.880 190.880 112.020 193.960 ;
        RECT 112.340 191.220 112.480 195.660 ;
        RECT 113.200 195.320 113.460 195.640 ;
        RECT 113.260 193.940 113.400 195.320 ;
        RECT 114.180 194.620 114.320 201.780 ;
        RECT 115.500 201.100 115.760 201.420 ;
        RECT 119.640 201.100 119.900 201.420 ;
        RECT 115.560 200.060 115.700 201.100 ;
        RECT 115.500 199.740 115.760 200.060 ;
        RECT 117.800 198.040 118.060 198.360 ;
        RECT 117.860 195.980 118.000 198.040 ;
        RECT 119.700 197.340 119.840 201.100 ;
        RECT 121.480 198.040 121.740 198.360 ;
        RECT 119.640 197.020 119.900 197.340 ;
        RECT 121.540 196.660 121.680 198.040 ;
        RECT 121.880 197.505 123.760 197.875 ;
        RECT 121.480 196.340 121.740 196.660 ;
        RECT 124.700 196.340 124.960 196.660 ;
        RECT 117.800 195.660 118.060 195.980 ;
        RECT 115.040 195.320 115.300 195.640 ;
        RECT 114.120 194.300 114.380 194.620 ;
        RECT 113.200 193.620 113.460 193.940 ;
        RECT 115.100 193.600 115.240 195.320 ;
        RECT 112.740 193.280 113.000 193.600 ;
        RECT 115.040 193.280 115.300 193.600 ;
        RECT 112.280 190.900 112.540 191.220 ;
        RECT 111.820 190.560 112.080 190.880 ;
        RECT 112.280 190.220 112.540 190.540 ;
        RECT 111.360 189.880 111.620 190.200 ;
        RECT 111.420 189.180 111.560 189.880 ;
        RECT 111.360 188.860 111.620 189.180 ;
        RECT 110.900 188.180 111.160 188.500 ;
        RECT 111.420 186.120 111.560 188.860 ;
        RECT 111.820 187.840 112.080 188.160 ;
        RECT 111.880 186.120 112.020 187.840 ;
        RECT 111.360 185.800 111.620 186.120 ;
        RECT 111.820 185.800 112.080 186.120 ;
        RECT 111.820 184.440 112.080 184.760 ;
        RECT 111.360 182.740 111.620 183.060 ;
        RECT 110.900 181.720 111.160 182.040 ;
        RECT 110.440 180.020 110.700 180.340 ;
        RECT 106.300 179.770 106.960 179.910 ;
        RECT 106.300 179.680 106.560 179.770 ;
        RECT 109.060 179.680 109.320 180.000 ;
        RECT 105.840 179.000 106.100 179.320 ;
        RECT 104.000 177.640 104.260 177.960 ;
        RECT 104.460 177.640 104.720 177.960 ;
        RECT 106.360 177.280 106.500 179.680 ;
        RECT 109.060 179.000 109.320 179.320 ;
        RECT 109.980 179.000 110.240 179.320 ;
        RECT 106.880 178.465 108.760 178.835 ;
        RECT 105.380 176.960 105.640 177.280 ;
        RECT 106.300 176.960 106.560 177.280 ;
        RECT 105.440 174.560 105.580 176.960 ;
        RECT 106.300 176.280 106.560 176.600 ;
        RECT 105.840 174.580 106.100 174.900 ;
        RECT 105.380 174.240 105.640 174.560 ;
        RECT 104.460 173.900 104.720 174.220 ;
        RECT 104.000 168.120 104.260 168.440 ;
        RECT 103.530 166.565 103.810 166.935 ;
        RECT 104.060 166.740 104.200 168.120 ;
        RECT 103.600 163.680 103.740 166.565 ;
        RECT 104.000 166.420 104.260 166.740 ;
        RECT 103.540 163.360 103.800 163.680 ;
        RECT 103.600 160.960 103.740 163.360 ;
        RECT 103.540 160.640 103.800 160.960 ;
        RECT 104.000 160.640 104.260 160.960 ;
        RECT 104.520 160.700 104.660 173.900 ;
        RECT 105.440 172.860 105.580 174.240 ;
        RECT 105.380 172.540 105.640 172.860 ;
        RECT 105.900 169.800 106.040 174.580 ;
        RECT 106.360 174.220 106.500 176.280 ;
        RECT 106.300 173.900 106.560 174.220 ;
        RECT 106.880 173.025 108.760 173.395 ;
        RECT 104.920 169.480 105.180 169.800 ;
        RECT 105.840 169.480 106.100 169.800 ;
        RECT 104.980 163.680 105.120 169.480 ;
        RECT 106.880 167.585 108.760 167.955 ;
        RECT 109.120 167.330 109.260 179.000 ;
        RECT 109.520 171.860 109.780 172.180 ;
        RECT 109.580 170.140 109.720 171.860 ;
        RECT 109.520 169.820 109.780 170.140 ;
        RECT 110.040 167.420 110.180 179.000 ;
        RECT 110.440 170.840 110.700 171.160 ;
        RECT 110.500 169.120 110.640 170.840 ;
        RECT 110.440 168.800 110.700 169.120 ;
        RECT 109.120 167.190 109.720 167.330 ;
        RECT 109.580 166.820 109.720 167.190 ;
        RECT 109.980 167.100 110.240 167.420 ;
        RECT 110.960 167.330 111.100 181.720 ;
        RECT 111.420 181.020 111.560 182.740 ;
        RECT 111.360 180.700 111.620 181.020 ;
        RECT 111.360 176.960 111.620 177.280 ;
        RECT 111.420 174.900 111.560 176.960 ;
        RECT 111.360 174.580 111.620 174.900 ;
        RECT 111.420 171.500 111.560 174.580 ;
        RECT 111.360 171.180 111.620 171.500 ;
        RECT 111.420 169.460 111.560 171.180 ;
        RECT 111.360 169.140 111.620 169.460 ;
        RECT 110.500 167.190 111.100 167.330 ;
        RECT 107.680 166.420 107.940 166.740 ;
        RECT 109.060 166.420 109.320 166.740 ;
        RECT 109.580 166.680 110.180 166.820 ;
        RECT 105.840 165.400 106.100 165.720 ;
        RECT 105.370 163.845 105.650 164.215 ;
        RECT 105.440 163.680 105.580 163.845 ;
        RECT 104.920 163.360 105.180 163.680 ;
        RECT 105.380 163.360 105.640 163.680 ;
        RECT 105.440 161.495 105.580 163.360 ;
        RECT 105.900 161.640 106.040 165.400 ;
        RECT 107.740 164.700 107.880 166.420 ;
        RECT 107.680 164.380 107.940 164.700 ;
        RECT 107.670 163.845 107.950 164.215 ;
        RECT 107.680 163.700 107.940 163.845 ;
        RECT 107.210 163.165 107.490 163.535 ;
        RECT 107.220 163.020 107.480 163.165 ;
        RECT 106.760 162.910 107.020 163.000 ;
        RECT 106.360 162.770 107.020 162.910 ;
        RECT 105.370 161.125 105.650 161.495 ;
        RECT 105.840 161.320 106.100 161.640 ;
        RECT 104.060 156.540 104.200 160.640 ;
        RECT 104.520 160.620 106.040 160.700 ;
        RECT 104.520 160.560 106.100 160.620 ;
        RECT 105.840 160.300 106.100 160.560 ;
        RECT 105.380 158.940 105.640 159.260 ;
        RECT 104.000 156.220 104.260 156.540 ;
        RECT 103.540 155.200 103.800 155.520 ;
        RECT 103.600 153.480 103.740 155.200 ;
        RECT 103.540 153.160 103.800 153.480 ;
        RECT 103.600 147.700 103.740 153.160 ;
        RECT 104.460 150.100 104.720 150.420 ;
        RECT 103.080 147.380 103.340 147.700 ;
        RECT 103.540 147.380 103.800 147.700 ;
        RECT 103.080 146.360 103.340 146.680 ;
        RECT 102.160 145.000 102.420 145.320 ;
        RECT 102.220 142.260 102.360 145.000 ;
        RECT 102.160 141.940 102.420 142.260 ;
        RECT 102.220 139.540 102.360 141.940 ;
        RECT 102.160 139.220 102.420 139.540 ;
        RECT 99.860 138.880 100.120 139.200 ;
        RECT 100.320 135.480 100.580 135.800 ;
        RECT 99.000 134.040 99.600 134.180 ;
        RECT 98.480 131.060 98.740 131.380 ;
        RECT 96.640 128.340 96.900 128.660 ;
        RECT 98.540 125.940 98.680 131.060 ;
        RECT 98.480 125.620 98.740 125.940 ;
        RECT 95.720 125.280 95.980 125.600 ;
        RECT 99.000 123.220 99.140 134.040 ;
        RECT 99.400 130.720 99.660 131.040 ;
        RECT 99.460 129.340 99.600 130.720 ;
        RECT 99.400 129.020 99.660 129.340 ;
        RECT 100.380 128.660 100.520 135.480 ;
        RECT 101.700 134.120 101.960 134.440 ;
        RECT 101.760 132.060 101.900 134.120 ;
        RECT 101.700 131.740 101.960 132.060 ;
        RECT 100.320 128.340 100.580 128.660 ;
        RECT 103.140 123.220 103.280 146.360 ;
        RECT 104.520 145.660 104.660 150.100 ;
        RECT 104.460 145.340 104.720 145.660 ;
        RECT 105.440 140.220 105.580 158.940 ;
        RECT 105.900 152.800 106.040 160.300 ;
        RECT 106.360 158.240 106.500 162.770 ;
        RECT 106.760 162.680 107.020 162.770 ;
        RECT 106.880 162.145 108.760 162.515 ;
        RECT 109.120 161.980 109.260 166.420 ;
        RECT 109.060 161.660 109.320 161.980 ;
        RECT 107.670 161.125 107.950 161.495 ;
        RECT 107.740 158.580 107.880 161.125 ;
        RECT 108.600 160.980 108.860 161.300 ;
        RECT 108.140 160.640 108.400 160.960 ;
        RECT 108.200 160.280 108.340 160.640 ;
        RECT 108.140 159.960 108.400 160.280 ;
        RECT 108.660 160.135 108.800 160.980 ;
        RECT 108.590 159.765 108.870 160.135 ;
        RECT 109.520 159.960 109.780 160.280 ;
        RECT 107.680 158.260 107.940 158.580 ;
        RECT 106.300 157.920 106.560 158.240 ;
        RECT 108.660 157.980 108.800 159.765 ;
        RECT 109.580 158.580 109.720 159.960 ;
        RECT 109.520 158.260 109.780 158.580 ;
        RECT 108.660 157.900 109.260 157.980 ;
        RECT 108.660 157.840 109.320 157.900 ;
        RECT 109.060 157.580 109.320 157.840 ;
        RECT 106.880 156.705 108.760 157.075 ;
        RECT 107.680 155.540 107.940 155.860 ;
        RECT 106.300 154.520 106.560 154.840 ;
        RECT 105.840 152.480 106.100 152.800 ;
        RECT 105.840 146.360 106.100 146.680 ;
        RECT 105.900 144.980 106.040 146.360 ;
        RECT 105.840 144.660 106.100 144.980 ;
        RECT 106.360 144.380 106.500 154.520 ;
        RECT 107.740 153.820 107.880 155.540 ;
        RECT 107.680 153.500 107.940 153.820 ;
        RECT 109.120 152.800 109.260 157.580 ;
        RECT 110.040 155.520 110.180 166.680 ;
        RECT 110.500 161.495 110.640 167.190 ;
        RECT 110.900 166.420 111.160 166.740 ;
        RECT 110.960 164.360 111.100 166.420 ;
        RECT 111.360 165.400 111.620 165.720 ;
        RECT 110.900 164.040 111.160 164.360 ;
        RECT 110.890 163.165 111.170 163.535 ;
        RECT 110.430 161.125 110.710 161.495 ;
        RECT 109.980 155.200 110.240 155.520 ;
        RECT 109.060 152.480 109.320 152.800 ;
        RECT 109.520 152.480 109.780 152.800 ;
        RECT 109.120 152.120 109.260 152.480 ;
        RECT 109.060 151.800 109.320 152.120 ;
        RECT 106.880 151.265 108.760 151.635 ;
        RECT 108.140 150.780 108.400 151.100 ;
        RECT 107.220 149.080 107.480 149.400 ;
        RECT 107.280 147.360 107.420 149.080 ;
        RECT 108.200 147.700 108.340 150.780 ;
        RECT 109.120 150.420 109.260 151.800 ;
        RECT 109.060 150.100 109.320 150.420 ;
        RECT 109.580 149.740 109.720 152.480 ;
        RECT 110.440 152.140 110.700 152.460 ;
        RECT 110.500 149.740 110.640 152.140 ;
        RECT 109.520 149.420 109.780 149.740 ;
        RECT 110.440 149.420 110.700 149.740 ;
        RECT 109.060 148.060 109.320 148.380 ;
        RECT 108.140 147.380 108.400 147.700 ;
        RECT 107.220 147.040 107.480 147.360 ;
        RECT 106.880 145.825 108.760 146.195 ;
        RECT 105.900 144.240 106.500 144.380 ;
        RECT 105.380 139.900 105.640 140.220 ;
        RECT 105.900 139.200 106.040 144.240 ;
        RECT 109.120 142.940 109.260 148.060 ;
        RECT 110.440 147.270 110.700 147.360 ;
        RECT 110.960 147.270 111.100 163.165 ;
        RECT 111.420 147.360 111.560 165.400 ;
        RECT 111.880 160.135 112.020 184.440 ;
        RECT 112.340 183.740 112.480 190.220 ;
        RECT 112.800 189.180 112.940 193.280 ;
        RECT 112.740 188.860 113.000 189.180 ;
        RECT 112.800 185.440 112.940 188.860 ;
        RECT 112.740 185.120 113.000 185.440 ;
        RECT 113.200 185.120 113.460 185.440 ;
        RECT 113.260 183.740 113.400 185.120 ;
        RECT 112.280 183.420 112.540 183.740 ;
        RECT 113.200 183.420 113.460 183.740 ;
        RECT 112.740 180.930 113.000 181.020 ;
        RECT 113.260 180.930 113.400 183.420 ;
        RECT 113.660 181.720 113.920 182.040 ;
        RECT 114.580 181.720 114.840 182.040 ;
        RECT 112.740 180.790 113.400 180.930 ;
        RECT 112.740 180.700 113.000 180.790 ;
        RECT 112.800 180.000 112.940 180.700 ;
        RECT 112.740 179.680 113.000 180.000 ;
        RECT 113.720 179.660 113.860 181.720 ;
        RECT 113.660 179.340 113.920 179.660 ;
        RECT 112.280 173.900 112.540 174.220 ;
        RECT 112.340 170.140 112.480 173.900 ;
        RECT 113.660 171.520 113.920 171.840 ;
        RECT 113.720 170.140 113.860 171.520 ;
        RECT 112.280 169.820 112.540 170.140 ;
        RECT 113.660 169.820 113.920 170.140 ;
        RECT 113.200 167.100 113.460 167.420 ;
        RECT 112.730 166.650 113.010 166.935 ;
        RECT 112.340 166.565 113.010 166.650 ;
        RECT 112.340 166.510 113.000 166.565 ;
        RECT 112.340 164.020 112.480 166.510 ;
        RECT 112.740 166.420 113.000 166.510 ;
        RECT 113.260 164.700 113.400 167.100 ;
        RECT 114.120 166.420 114.380 166.740 ;
        RECT 113.660 165.740 113.920 166.060 ;
        RECT 113.200 164.380 113.460 164.700 ;
        RECT 113.260 164.215 113.400 164.380 ;
        RECT 112.280 163.700 112.540 164.020 ;
        RECT 113.190 163.845 113.470 164.215 ;
        RECT 113.260 163.680 113.400 163.845 ;
        RECT 112.740 163.535 113.000 163.680 ;
        RECT 112.730 163.165 113.010 163.535 ;
        RECT 113.200 163.360 113.460 163.680 ;
        RECT 112.280 162.680 112.540 163.000 ;
        RECT 111.810 159.765 112.090 160.135 ;
        RECT 112.340 159.340 112.480 162.680 ;
        RECT 112.740 160.300 113.000 160.620 ;
        RECT 111.880 159.200 112.480 159.340 ;
        RECT 111.880 156.200 112.020 159.200 ;
        RECT 112.800 158.830 112.940 160.300 ;
        RECT 113.190 159.765 113.470 160.135 ;
        RECT 112.340 158.690 112.940 158.830 ;
        RECT 112.340 158.240 112.480 158.690 ;
        RECT 113.260 158.490 113.400 159.765 ;
        RECT 112.800 158.350 113.400 158.490 ;
        RECT 112.280 157.920 112.540 158.240 ;
        RECT 112.800 157.300 112.940 158.350 ;
        RECT 112.340 157.160 112.940 157.300 ;
        RECT 113.200 157.240 113.460 157.560 ;
        RECT 111.820 155.880 112.080 156.200 ;
        RECT 111.820 154.520 112.080 154.840 ;
        RECT 110.440 147.130 111.100 147.270 ;
        RECT 110.440 147.040 110.700 147.130 ;
        RECT 111.360 147.040 111.620 147.360 ;
        RECT 109.520 146.360 109.780 146.680 ;
        RECT 110.440 146.360 110.700 146.680 ;
        RECT 109.060 142.620 109.320 142.940 ;
        RECT 106.300 141.600 106.560 141.920 ;
        RECT 109.060 141.600 109.320 141.920 ;
        RECT 106.360 139.620 106.500 141.600 ;
        RECT 106.880 140.385 108.760 140.755 ;
        RECT 109.120 140.130 109.260 141.600 ;
        RECT 108.660 139.990 109.260 140.130 ;
        RECT 106.760 139.620 107.020 139.880 ;
        RECT 106.360 139.560 107.020 139.620 ;
        RECT 106.360 139.480 106.960 139.560 ;
        RECT 108.660 139.540 108.800 139.990 ;
        RECT 105.840 138.880 106.100 139.200 ;
        RECT 105.380 136.500 105.640 136.820 ;
        RECT 105.440 134.100 105.580 136.500 ;
        RECT 106.360 135.800 106.500 139.480 ;
        RECT 108.600 139.220 108.860 139.540 ;
        RECT 109.060 138.880 109.320 139.200 ;
        RECT 106.300 135.480 106.560 135.800 ;
        RECT 106.360 134.440 106.500 135.480 ;
        RECT 106.880 134.945 108.760 135.315 ;
        RECT 106.300 134.120 106.560 134.440 ;
        RECT 105.380 133.780 105.640 134.100 ;
        RECT 103.540 133.440 103.800 133.760 ;
        RECT 103.600 132.060 103.740 133.440 ;
        RECT 104.460 132.760 104.720 133.080 ;
        RECT 103.540 131.740 103.800 132.060 ;
        RECT 104.520 131.040 104.660 132.760 ;
        RECT 105.440 131.380 105.580 133.780 ;
        RECT 106.760 133.440 107.020 133.760 ;
        RECT 106.820 131.380 106.960 133.440 ;
        RECT 105.380 131.060 105.640 131.380 ;
        RECT 106.760 131.060 107.020 131.380 ;
        RECT 109.120 131.040 109.260 138.880 ;
        RECT 104.460 130.720 104.720 131.040 ;
        RECT 109.060 130.720 109.320 131.040 ;
        RECT 106.880 129.505 108.760 129.875 ;
        RECT 109.120 129.340 109.260 130.720 ;
        RECT 109.060 129.020 109.320 129.340 ;
        RECT 108.600 128.680 108.860 129.000 ;
        RECT 108.660 125.600 108.800 128.680 ;
        RECT 108.600 125.280 108.860 125.600 ;
        RECT 106.880 124.065 108.760 124.435 ;
        RECT 109.580 123.220 109.720 146.360 ;
        RECT 109.980 137.180 110.240 137.500 ;
        RECT 110.040 125.600 110.180 137.180 ;
        RECT 109.980 125.280 110.240 125.600 ;
        RECT 91.120 122.900 91.380 123.220 ;
        RECT 98.940 122.900 99.200 123.220 ;
        RECT 103.080 122.900 103.340 123.220 ;
        RECT 109.520 122.900 109.780 123.220 ;
        RECT 89.280 119.840 89.540 120.160 ;
        RECT 86.520 119.500 86.780 119.820 ;
        RECT 86.580 118.460 86.720 119.500 ;
        RECT 86.520 118.140 86.780 118.460 ;
        RECT 88.360 117.800 88.620 118.120 ;
        RECT 85.600 117.460 85.860 117.780 ;
        RECT 87.440 117.460 87.700 117.780 ;
        RECT 87.900 117.460 88.160 117.780 ;
        RECT 85.140 116.440 85.400 116.760 ;
        RECT 87.500 114.720 87.640 117.460 ;
        RECT 87.960 115.740 88.100 117.460 ;
        RECT 87.900 115.420 88.160 115.740 ;
        RECT 87.440 114.400 87.700 114.720 ;
        RECT 86.580 104.800 87.180 104.940 ;
        RECT 86.580 104.340 86.720 104.800 ;
        RECT 30.850 102.340 31.130 104.340 ;
        RECT 35.910 102.340 36.190 104.340 ;
        RECT 40.970 102.340 41.250 104.340 ;
        RECT 46.030 102.340 46.310 104.340 ;
        RECT 51.090 102.340 51.370 104.340 ;
        RECT 56.150 102.340 56.430 104.340 ;
        RECT 61.210 102.340 61.490 104.340 ;
        RECT 66.270 102.340 66.550 104.340 ;
        RECT 71.330 102.340 71.610 104.340 ;
        RECT 76.390 102.340 76.670 104.340 ;
        RECT 81.450 102.340 81.730 104.340 ;
        RECT 86.510 102.340 86.790 104.340 ;
        RECT 87.040 104.260 87.180 104.800 ;
        RECT 88.420 104.260 88.560 117.800 ;
        RECT 89.340 117.440 89.480 119.840 ;
        RECT 90.660 119.160 90.920 119.480 ;
        RECT 90.720 118.460 90.860 119.160 ;
        RECT 90.660 118.140 90.920 118.460 ;
        RECT 89.280 117.120 89.540 117.440 ;
        RECT 91.180 114.720 91.320 122.900 ;
        RECT 94.800 121.880 95.060 122.200 ;
        RECT 98.020 121.880 98.280 122.200 ;
        RECT 99.860 121.880 100.120 122.200 ;
        RECT 104.000 121.880 104.260 122.200 ;
        RECT 109.520 121.880 109.780 122.200 ;
        RECT 91.880 121.345 93.760 121.715 ;
        RECT 91.880 115.905 93.760 116.275 ;
        RECT 91.120 114.400 91.380 114.720 ;
        RECT 91.180 114.040 91.320 114.400 ;
        RECT 94.860 114.380 95.000 121.880 ;
        RECT 96.640 120.180 96.900 120.500 ;
        RECT 91.580 114.060 91.840 114.380 ;
        RECT 94.800 114.060 95.060 114.380 ;
        RECT 91.120 113.720 91.380 114.040 ;
        RECT 91.640 104.340 91.780 114.060 ;
        RECT 96.700 104.340 96.840 120.180 ;
        RECT 97.560 119.500 97.820 119.820 ;
        RECT 97.620 115.740 97.760 119.500 ;
        RECT 97.560 115.420 97.820 115.740 ;
        RECT 98.080 115.060 98.220 121.880 ;
        RECT 99.920 120.500 100.060 121.880 ;
        RECT 99.860 120.180 100.120 120.500 ;
        RECT 101.240 119.840 101.500 120.160 ;
        RECT 101.300 117.440 101.440 119.840 ;
        RECT 104.060 118.460 104.200 121.880 ;
        RECT 109.580 120.500 109.720 121.880 ;
        RECT 105.840 120.410 106.100 120.500 ;
        RECT 105.840 120.270 106.500 120.410 ;
        RECT 105.840 120.180 106.100 120.270 ;
        RECT 104.000 118.140 104.260 118.460 ;
        RECT 101.700 117.460 101.960 117.780 ;
        RECT 103.080 117.460 103.340 117.780 ;
        RECT 99.400 117.120 99.660 117.440 ;
        RECT 101.240 117.120 101.500 117.440 ;
        RECT 99.460 115.060 99.600 117.120 ;
        RECT 98.020 114.740 98.280 115.060 ;
        RECT 99.400 114.740 99.660 115.060 ;
        RECT 101.760 104.340 101.900 117.460 ;
        RECT 103.140 115.740 103.280 117.460 ;
        RECT 103.540 116.440 103.800 116.760 ;
        RECT 103.600 115.740 103.740 116.440 ;
        RECT 103.080 115.420 103.340 115.740 ;
        RECT 103.540 115.420 103.800 115.740 ;
        RECT 106.360 111.840 106.500 120.270 ;
        RECT 109.520 120.180 109.780 120.500 ;
        RECT 110.500 119.820 110.640 146.360 ;
        RECT 110.900 141.600 111.160 141.920 ;
        RECT 110.960 139.540 111.100 141.600 ;
        RECT 110.900 139.220 111.160 139.540 ;
        RECT 110.960 135.800 111.100 139.220 ;
        RECT 110.900 135.480 111.160 135.800 ;
        RECT 111.880 123.220 112.020 154.520 ;
        RECT 112.340 151.100 112.480 157.160 ;
        RECT 113.260 155.860 113.400 157.240 ;
        RECT 113.200 155.540 113.460 155.860 ;
        RECT 112.740 153.160 113.000 153.480 ;
        RECT 112.800 152.800 112.940 153.160 ;
        RECT 112.740 152.480 113.000 152.800 ;
        RECT 113.200 152.480 113.460 152.800 ;
        RECT 113.260 152.120 113.400 152.480 ;
        RECT 113.200 151.800 113.460 152.120 ;
        RECT 112.280 150.780 112.540 151.100 ;
        RECT 112.740 150.440 113.000 150.760 ;
        RECT 112.280 148.060 112.540 148.380 ;
        RECT 112.340 142.940 112.480 148.060 ;
        RECT 112.800 146.680 112.940 150.440 ;
        RECT 112.740 146.360 113.000 146.680 ;
        RECT 113.720 142.940 113.860 165.740 ;
        RECT 114.180 164.020 114.320 166.420 ;
        RECT 114.120 163.700 114.380 164.020 ;
        RECT 114.120 157.580 114.380 157.900 ;
        RECT 114.180 156.540 114.320 157.580 ;
        RECT 114.120 156.220 114.380 156.540 ;
        RECT 114.640 153.900 114.780 181.720 ;
        RECT 115.100 180.680 115.240 193.280 ;
        RECT 121.880 192.065 123.760 192.435 ;
        RECT 124.760 190.540 124.900 196.340 ;
        RECT 124.240 190.220 124.500 190.540 ;
        RECT 124.700 190.220 124.960 190.540 ;
        RECT 115.960 189.880 116.220 190.200 ;
        RECT 116.420 189.880 116.680 190.200 ;
        RECT 117.340 189.880 117.600 190.200 ;
        RECT 116.020 185.440 116.160 189.880 ;
        RECT 116.480 186.120 116.620 189.880 ;
        RECT 116.420 185.800 116.680 186.120 ;
        RECT 117.400 185.780 117.540 189.880 ;
        RECT 121.480 187.160 121.740 187.480 ;
        RECT 121.540 186.460 121.680 187.160 ;
        RECT 121.880 186.625 123.760 186.995 ;
        RECT 124.300 186.460 124.440 190.220 ;
        RECT 124.760 188.160 124.900 190.220 ;
        RECT 124.700 187.840 124.960 188.160 ;
        RECT 121.480 186.140 121.740 186.460 ;
        RECT 124.240 186.140 124.500 186.460 ;
        RECT 117.340 185.460 117.600 185.780 ;
        RECT 115.960 185.120 116.220 185.440 ;
        RECT 117.400 183.060 117.540 185.460 ;
        RECT 121.940 185.120 122.200 185.440 ;
        RECT 118.720 184.440 118.980 184.760 ;
        RECT 118.780 183.060 118.920 184.440 ;
        RECT 122.000 183.740 122.140 185.120 ;
        RECT 121.940 183.420 122.200 183.740 ;
        RECT 115.960 182.740 116.220 183.060 ;
        RECT 117.340 182.740 117.600 183.060 ;
        RECT 118.720 182.740 118.980 183.060 ;
        RECT 119.180 182.740 119.440 183.060 ;
        RECT 115.040 180.360 115.300 180.680 ;
        RECT 116.020 177.620 116.160 182.740 ;
        RECT 118.720 180.360 118.980 180.680 ;
        RECT 116.420 180.020 116.680 180.340 ;
        RECT 115.960 177.300 116.220 177.620 ;
        RECT 115.040 174.240 115.300 174.560 ;
        RECT 115.100 172.520 115.240 174.240 ;
        RECT 116.020 172.520 116.160 177.300 ;
        RECT 116.480 176.600 116.620 180.020 ;
        RECT 117.340 179.000 117.600 179.320 ;
        RECT 116.420 176.280 116.680 176.600 ;
        RECT 115.040 172.200 115.300 172.520 ;
        RECT 115.960 172.200 116.220 172.520 ;
        RECT 115.500 168.120 115.760 168.440 ;
        RECT 115.560 166.740 115.700 168.120 ;
        RECT 115.500 166.420 115.760 166.740 ;
        RECT 115.960 166.080 116.220 166.400 ;
        RECT 116.020 161.300 116.160 166.080 ;
        RECT 116.480 164.360 116.620 176.280 ;
        RECT 117.400 174.900 117.540 179.000 ;
        RECT 117.800 176.960 118.060 177.280 ;
        RECT 117.340 174.580 117.600 174.900 ;
        RECT 117.400 172.860 117.540 174.580 ;
        RECT 117.860 174.560 118.000 176.960 ;
        RECT 118.780 175.240 118.920 180.360 ;
        RECT 119.240 178.300 119.380 182.740 ;
        RECT 124.240 181.720 124.500 182.040 ;
        RECT 121.880 181.185 123.760 181.555 ;
        RECT 124.300 180.340 124.440 181.720 ;
        RECT 124.240 180.020 124.500 180.340 ;
        RECT 126.080 179.680 126.340 180.000 ;
        RECT 119.180 177.980 119.440 178.300 ;
        RECT 124.240 177.640 124.500 177.960 ;
        RECT 121.880 175.745 123.760 176.115 ;
        RECT 118.720 174.920 118.980 175.240 ;
        RECT 117.800 174.240 118.060 174.560 ;
        RECT 117.340 172.540 117.600 172.860 ;
        RECT 117.340 171.520 117.600 171.840 ;
        RECT 117.400 169.120 117.540 171.520 ;
        RECT 117.340 168.800 117.600 169.120 ;
        RECT 117.400 167.420 117.540 168.800 ;
        RECT 117.340 167.100 117.600 167.420 ;
        RECT 116.420 164.040 116.680 164.360 ;
        RECT 116.880 163.535 117.140 163.680 ;
        RECT 116.870 163.165 117.150 163.535 ;
        RECT 118.780 163.340 118.920 174.920 ;
        RECT 123.770 174.725 124.050 175.095 ;
        RECT 123.780 174.580 124.040 174.725 ;
        RECT 122.860 173.560 123.120 173.880 ;
        RECT 122.920 172.180 123.060 173.560 ;
        RECT 122.860 171.860 123.120 172.180 ;
        RECT 123.840 171.580 123.980 174.580 ;
        RECT 124.300 172.860 124.440 177.640 ;
        RECT 126.140 177.280 126.280 179.680 ;
        RECT 130.670 178.125 130.950 178.495 ;
        RECT 126.080 176.960 126.340 177.280 ;
        RECT 126.140 174.220 126.280 176.960 ;
        RECT 130.740 174.560 130.880 178.125 ;
        RECT 130.680 174.240 130.940 174.560 ;
        RECT 126.080 173.900 126.340 174.220 ;
        RECT 124.240 172.540 124.500 172.860 ;
        RECT 123.840 171.440 124.900 171.580 ;
        RECT 120.560 170.840 120.820 171.160 ;
        RECT 124.240 170.840 124.500 171.160 ;
        RECT 120.620 168.780 120.760 170.840 ;
        RECT 121.880 170.305 123.760 170.675 ;
        RECT 124.300 169.460 124.440 170.840 ;
        RECT 124.240 169.140 124.500 169.460 ;
        RECT 120.560 168.460 120.820 168.780 ;
        RECT 124.760 166.740 124.900 171.440 ;
        RECT 126.140 169.120 126.280 173.900 ;
        RECT 135.630 173.380 136.780 174.600 ;
        RECT 129.290 170.560 133.760 172.150 ;
        RECT 126.080 168.800 126.340 169.120 ;
        RECT 124.700 166.420 124.960 166.740 ;
        RECT 121.880 164.865 123.760 165.235 ;
        RECT 118.720 163.020 118.980 163.340 ;
        RECT 120.100 161.660 120.360 161.980 ;
        RECT 115.960 160.980 116.220 161.300 ;
        RECT 115.500 159.960 115.760 160.280 ;
        RECT 116.020 160.140 116.160 160.980 ;
        RECT 116.020 160.000 116.620 160.140 ;
        RECT 115.560 158.240 115.700 159.960 ;
        RECT 115.500 157.920 115.760 158.240 ;
        RECT 116.480 155.180 116.620 160.000 ;
        RECT 117.800 158.260 118.060 158.580 ;
        RECT 116.420 154.860 116.680 155.180 ;
        RECT 114.180 153.760 114.780 153.900 ;
        RECT 114.180 147.700 114.320 153.760 ;
        RECT 115.500 153.500 115.760 153.820 ;
        RECT 114.580 151.800 114.840 152.120 ;
        RECT 114.120 147.380 114.380 147.700 ;
        RECT 114.640 147.360 114.780 151.800 ;
        RECT 114.580 147.040 114.840 147.360 ;
        RECT 115.560 144.640 115.700 153.500 ;
        RECT 116.480 150.420 116.620 154.860 ;
        RECT 117.860 153.820 118.000 158.260 ;
        RECT 118.720 157.240 118.980 157.560 ;
        RECT 118.780 155.180 118.920 157.240 ;
        RECT 118.720 154.860 118.980 155.180 ;
        RECT 117.800 153.500 118.060 153.820 ;
        RECT 118.780 152.800 118.920 154.860 ;
        RECT 118.720 152.480 118.980 152.800 ;
        RECT 116.880 151.800 117.140 152.120 ;
        RECT 116.940 150.420 117.080 151.800 ;
        RECT 116.420 150.100 116.680 150.420 ;
        RECT 116.880 150.100 117.140 150.420 ;
        RECT 115.960 149.080 116.220 149.400 ;
        RECT 116.020 147.020 116.160 149.080 ;
        RECT 115.960 146.700 116.220 147.020 ;
        RECT 116.420 146.360 116.680 146.680 ;
        RECT 116.480 145.660 116.620 146.360 ;
        RECT 116.940 145.660 117.080 150.100 ;
        RECT 116.420 145.340 116.680 145.660 ;
        RECT 116.880 145.340 117.140 145.660 ;
        RECT 115.500 144.320 115.760 144.640 ;
        RECT 112.280 142.620 112.540 142.940 ;
        RECT 113.660 142.620 113.920 142.940 ;
        RECT 113.200 141.940 113.460 142.260 ;
        RECT 113.260 139.200 113.400 141.940 ;
        RECT 114.580 141.600 114.840 141.920 ;
        RECT 113.200 138.880 113.460 139.200 ;
        RECT 112.280 138.200 112.540 138.520 ;
        RECT 112.740 138.200 113.000 138.520 ;
        RECT 112.340 136.140 112.480 138.200 ;
        RECT 112.800 136.820 112.940 138.200 ;
        RECT 112.740 136.500 113.000 136.820 ;
        RECT 112.280 135.820 112.540 136.140 ;
        RECT 113.260 133.760 113.400 138.880 ;
        RECT 113.200 133.440 113.460 133.760 ;
        RECT 113.260 131.380 113.400 133.440 ;
        RECT 113.200 131.060 113.460 131.380 ;
        RECT 114.640 130.360 114.780 141.600 ;
        RECT 116.880 140.920 117.140 141.240 ;
        RECT 118.720 140.920 118.980 141.240 ;
        RECT 115.040 139.560 115.300 139.880 ;
        RECT 115.100 137.500 115.240 139.560 ;
        RECT 116.940 138.860 117.080 140.920 ;
        RECT 116.880 138.540 117.140 138.860 ;
        RECT 116.940 138.260 117.080 138.540 ;
        RECT 116.480 138.120 117.080 138.260 ;
        RECT 115.040 137.180 115.300 137.500 ;
        RECT 116.480 134.780 116.620 138.120 ;
        RECT 116.880 135.480 117.140 135.800 ;
        RECT 116.940 134.780 117.080 135.480 ;
        RECT 116.420 134.460 116.680 134.780 ;
        RECT 116.880 134.460 117.140 134.780 ;
        RECT 118.780 134.440 118.920 140.920 ;
        RECT 119.180 136.160 119.440 136.480 ;
        RECT 118.720 134.120 118.980 134.440 ;
        RECT 119.240 134.100 119.380 136.160 ;
        RECT 119.640 135.820 119.900 136.140 ;
        RECT 119.700 134.780 119.840 135.820 ;
        RECT 119.640 134.460 119.900 134.780 ;
        RECT 119.180 133.780 119.440 134.100 ;
        RECT 119.240 130.700 119.380 133.780 ;
        RECT 119.180 130.380 119.440 130.700 ;
        RECT 112.280 130.040 112.540 130.360 ;
        RECT 114.580 130.040 114.840 130.360 ;
        RECT 117.800 130.040 118.060 130.360 ;
        RECT 112.340 128.660 112.480 130.040 ;
        RECT 114.640 129.340 114.780 130.040 ;
        RECT 114.580 129.020 114.840 129.340 ;
        RECT 117.860 129.000 118.000 130.040 ;
        RECT 117.800 128.680 118.060 129.000 ;
        RECT 112.280 128.340 112.540 128.660 ;
        RECT 119.640 125.280 119.900 125.600 ;
        RECT 120.160 125.510 120.300 161.660 ;
        RECT 126.140 161.300 126.280 168.800 ;
        RECT 135.630 166.640 136.740 173.380 ;
        RECT 135.630 165.420 136.780 166.640 ;
        RECT 126.080 160.980 126.340 161.300 ;
        RECT 124.700 160.640 124.960 160.960 ;
        RECT 121.880 159.425 123.760 159.795 ;
        RECT 124.760 159.260 124.900 160.640 ;
        RECT 124.700 158.940 124.960 159.260 ;
        RECT 120.560 158.660 120.820 158.920 ;
        RECT 120.560 158.600 121.220 158.660 ;
        RECT 120.620 158.520 121.220 158.600 ;
        RECT 120.560 147.040 120.820 147.360 ;
        RECT 120.620 145.660 120.760 147.040 ;
        RECT 120.560 145.340 120.820 145.660 ;
        RECT 121.080 139.440 121.220 158.520 ;
        RECT 124.240 157.240 124.500 157.560 ;
        RECT 124.300 155.860 124.440 157.240 ;
        RECT 124.240 155.540 124.500 155.860 ;
        RECT 126.080 155.200 126.340 155.520 ;
        RECT 121.880 153.985 123.760 154.355 ;
        RECT 121.480 151.800 121.740 152.120 ;
        RECT 121.540 147.360 121.680 151.800 ;
        RECT 126.140 150.420 126.280 155.200 ;
        RECT 124.240 150.100 124.500 150.420 ;
        RECT 126.080 150.100 126.340 150.420 ;
        RECT 121.880 148.545 123.760 148.915 ;
        RECT 124.300 148.380 124.440 150.100 ;
        RECT 124.240 148.060 124.500 148.380 ;
        RECT 126.140 147.700 126.280 150.100 ;
        RECT 126.080 147.380 126.340 147.700 ;
        RECT 121.480 147.040 121.740 147.360 ;
        RECT 121.880 143.105 123.760 143.475 ;
        RECT 121.080 139.300 121.680 139.440 ;
        RECT 120.560 125.510 120.820 125.600 ;
        RECT 120.160 125.370 120.820 125.510 ;
        RECT 121.540 125.510 121.680 139.300 ;
        RECT 126.140 139.200 126.280 147.380 ;
        RECT 135.630 141.200 136.780 141.270 ;
        RECT 135.630 140.180 136.800 141.200 ;
        RECT 124.240 138.880 124.500 139.200 ;
        RECT 126.080 138.880 126.340 139.200 ;
        RECT 121.880 137.665 123.760 138.035 ;
        RECT 122.860 136.160 123.120 136.480 ;
        RECT 122.920 134.780 123.060 136.160 ;
        RECT 124.300 134.780 124.440 138.880 ;
        RECT 129.140 138.175 134.100 139.455 ;
        RECT 125.160 136.160 125.420 136.480 ;
        RECT 122.860 134.460 123.120 134.780 ;
        RECT 124.240 134.460 124.500 134.780 ;
        RECT 121.880 132.225 123.760 132.595 ;
        RECT 122.400 130.040 122.660 130.360 ;
        RECT 122.460 128.660 122.600 130.040 ;
        RECT 125.220 128.660 125.360 136.160 ;
        RECT 135.640 133.320 136.800 140.180 ;
        RECT 122.400 128.340 122.660 128.660 ;
        RECT 125.160 128.340 125.420 128.660 ;
        RECT 121.880 126.785 123.760 127.155 ;
        RECT 123.320 125.510 123.580 125.600 ;
        RECT 121.540 125.370 123.580 125.510 ;
        RECT 120.560 125.280 120.820 125.370 ;
        RECT 123.320 125.280 123.580 125.370 ;
        RECT 117.340 124.940 117.600 125.260 ;
        RECT 117.400 123.560 117.540 124.940 ;
        RECT 117.340 123.240 117.600 123.560 ;
        RECT 111.820 122.900 112.080 123.220 ;
        RECT 113.200 122.560 113.460 122.880 ;
        RECT 113.260 120.160 113.400 122.560 ;
        RECT 117.340 121.880 117.600 122.200 ;
        RECT 113.200 119.840 113.460 120.160 ;
        RECT 109.520 119.500 109.780 119.820 ;
        RECT 110.440 119.500 110.700 119.820 ;
        RECT 106.880 118.625 108.760 118.995 ;
        RECT 109.580 118.460 109.720 119.500 ;
        RECT 112.740 119.160 113.000 119.480 ;
        RECT 109.520 118.140 109.780 118.460 ;
        RECT 110.440 117.460 110.700 117.780 ;
        RECT 110.500 115.060 110.640 117.460 ;
        RECT 112.280 116.440 112.540 116.760 ;
        RECT 110.440 114.740 110.700 115.060 ;
        RECT 112.340 114.380 112.480 116.440 ;
        RECT 112.800 115.060 112.940 119.160 ;
        RECT 113.260 117.440 113.400 119.840 ;
        RECT 117.400 117.440 117.540 121.880 ;
        RECT 119.180 119.840 119.440 120.160 ;
        RECT 118.260 117.460 118.520 117.780 ;
        RECT 113.200 117.120 113.460 117.440 ;
        RECT 116.880 117.120 117.140 117.440 ;
        RECT 117.340 117.120 117.600 117.440 ;
        RECT 112.740 114.740 113.000 115.060 ;
        RECT 112.280 114.060 112.540 114.380 ;
        RECT 111.820 113.720 112.080 114.040 ;
        RECT 106.880 113.185 108.760 113.555 ;
        RECT 106.360 111.700 106.960 111.840 ;
        RECT 106.820 104.340 106.960 111.700 ;
        RECT 111.880 104.340 112.020 113.720 ;
        RECT 116.940 104.340 117.080 117.120 ;
        RECT 118.320 115.740 118.460 117.460 ;
        RECT 119.240 115.740 119.380 119.840 ;
        RECT 119.700 118.460 119.840 125.280 ;
        RECT 120.560 124.600 120.820 124.920 ;
        RECT 124.700 124.600 124.960 124.920 ;
        RECT 120.620 123.560 120.760 124.600 ;
        RECT 120.560 123.240 120.820 123.560 ;
        RECT 121.880 121.345 123.760 121.715 ;
        RECT 124.760 120.500 124.900 124.600 ;
        RECT 125.220 122.880 125.360 128.340 ;
        RECT 125.160 122.560 125.420 122.880 ;
        RECT 127.000 122.560 127.260 122.880 ;
        RECT 121.480 120.180 121.740 120.500 ;
        RECT 124.700 120.180 124.960 120.500 ;
        RECT 119.640 118.140 119.900 118.460 ;
        RECT 118.260 115.420 118.520 115.740 ;
        RECT 119.180 115.420 119.440 115.740 ;
        RECT 119.700 114.720 119.840 118.140 ;
        RECT 121.540 115.650 121.680 120.180 ;
        RECT 125.220 119.820 125.360 122.560 ;
        RECT 125.160 119.500 125.420 119.820 ;
        RECT 125.220 117.780 125.360 119.500 ;
        RECT 125.160 117.460 125.420 117.780 ;
        RECT 121.880 115.905 123.760 116.275 ;
        RECT 121.540 115.510 122.140 115.650 ;
        RECT 119.640 114.400 119.900 114.720 ;
        RECT 122.000 104.340 122.140 115.510 ;
        RECT 125.220 115.060 125.360 117.460 ;
        RECT 125.160 114.740 125.420 115.060 ;
        RECT 127.060 104.340 127.200 122.560 ;
        RECT 130.210 118.285 130.490 118.655 ;
        RECT 130.280 114.720 130.420 118.285 ;
        RECT 130.220 114.400 130.480 114.720 ;
        RECT 129.750 105.580 133.160 106.650 ;
        RECT 87.040 104.120 88.560 104.260 ;
        RECT 91.570 102.340 91.850 104.340 ;
        RECT 96.630 102.340 96.910 104.340 ;
        RECT 101.690 102.340 101.970 104.340 ;
        RECT 106.750 102.340 107.030 104.340 ;
        RECT 111.810 102.340 112.090 104.340 ;
        RECT 116.870 102.340 117.150 104.340 ;
        RECT 121.930 102.340 122.210 104.340 ;
        RECT 126.990 102.340 127.270 104.340 ;
        RECT 13.920 85.550 15.140 89.420 ;
        RECT 19.910 85.980 21.130 89.850 ;
        RECT 67.730 89.640 68.670 89.840 ;
        RECT 25.730 85.120 26.950 88.990 ;
        RECT 31.780 85.510 33.000 89.380 ;
        RECT 37.750 88.780 38.970 89.290 ;
        RECT 37.680 88.620 38.970 88.780 ;
        RECT 43.810 88.630 45.030 89.530 ;
        RECT 49.740 88.640 50.960 89.040 ;
        RECT 37.680 86.810 39.070 88.620 ;
        RECT 37.750 85.420 38.970 86.810 ;
        RECT 43.810 86.720 45.140 88.630 ;
        RECT 49.740 86.920 51.010 88.640 ;
        RECT 43.810 85.660 45.030 86.720 ;
        RECT 49.740 85.170 50.960 86.920 ;
        RECT 55.530 85.320 56.750 89.190 ;
        RECT 61.720 88.640 62.940 88.870 ;
        RECT 61.720 86.600 63.130 88.640 ;
        RECT 61.720 85.000 62.940 86.600 ;
        RECT 67.580 85.770 68.800 89.640 ;
        RECT 73.850 84.290 75.070 88.160 ;
        RECT 79.730 84.310 80.950 88.180 ;
        RECT 74.090 80.440 74.370 84.290 ;
        RECT 20.140 80.160 74.370 80.440 ;
        RECT 20.140 75.650 20.420 80.160 ;
        RECT 80.070 79.800 80.350 84.310 ;
        RECT 85.470 84.100 86.690 87.970 ;
        RECT 91.460 84.500 92.680 88.320 ;
        RECT 97.600 84.630 98.820 88.500 ;
        RECT 103.650 84.740 104.870 88.610 ;
        RECT 109.620 85.420 110.840 89.290 ;
        RECT 115.740 85.700 116.960 89.570 ;
        RECT 121.520 85.700 122.740 89.570 ;
        RECT 31.380 79.520 80.350 79.800 ;
        RECT 31.380 75.850 31.660 79.520 ;
        RECT 86.050 79.170 86.330 84.100 ;
        RECT 42.510 78.890 86.330 79.170 ;
        RECT 3.960 71.320 6.050 73.240 ;
        RECT 19.330 73.120 21.890 75.650 ;
        RECT 28.185 73.180 30.255 74.460 ;
        RECT 30.670 73.320 33.230 75.850 ;
        RECT 42.510 75.750 42.790 78.890 ;
        RECT 92.030 78.570 92.310 84.500 ;
        RECT 53.830 78.290 92.310 78.570 ;
        RECT 53.830 75.820 54.110 78.290 ;
        RECT 98.010 77.990 98.290 84.630 ;
        RECT 64.900 77.710 98.290 77.990 ;
        RECT 19.005 71.800 19.865 72.640 ;
        RECT 15.560 68.610 16.990 71.210 ;
        RECT 19.305 68.570 19.845 71.800 ;
        RECT 20.145 70.600 20.555 73.120 ;
        RECT 30.205 71.810 31.065 72.650 ;
        RECT 19.325 47.770 19.825 68.570 ;
        RECT 20.165 49.090 20.555 70.600 ;
        RECT 20.955 70.010 21.845 70.740 ;
        RECT 21.055 65.190 21.315 70.010 ;
        RECT 22.695 68.620 25.405 69.470 ;
        RECT 22.895 65.840 24.825 68.620 ;
        RECT 30.505 68.580 31.045 71.810 ;
        RECT 31.345 70.610 31.755 73.320 ;
        RECT 39.475 73.150 41.545 74.430 ;
        RECT 41.910 73.220 44.470 75.750 ;
        RECT 41.425 71.780 42.285 72.620 ;
        RECT 27.795 67.130 28.915 67.810 ;
        RECT 28.075 65.850 28.745 67.130 ;
        RECT 21.455 65.460 26.505 65.840 ;
        RECT 27.865 65.440 28.915 65.850 ;
        RECT 21.055 63.640 21.435 65.190 ;
        RECT 21.175 55.800 21.435 63.640 ;
        RECT 26.485 63.200 26.755 65.240 ;
        RECT 27.615 63.200 27.885 65.200 ;
        RECT 26.485 56.510 27.885 63.200 ;
        RECT 21.085 55.290 21.445 55.800 ;
        RECT 21.065 54.860 21.445 55.290 ;
        RECT 26.485 55.190 26.755 56.510 ;
        RECT 27.615 55.150 27.885 56.510 ;
        RECT 28.885 55.260 29.205 65.190 ;
        RECT 28.885 55.200 29.215 55.260 ;
        RECT 21.065 54.580 21.315 54.860 ;
        RECT 20.865 54.180 25.505 54.580 ;
        RECT 26.405 54.290 27.535 54.300 ;
        RECT 28.895 54.290 29.215 55.200 ;
        RECT 21.065 52.060 21.315 54.180 ;
        RECT 25.765 53.490 26.125 54.110 ;
        RECT 25.845 52.610 26.105 53.490 ;
        RECT 26.385 53.240 29.215 54.290 ;
        RECT 25.675 52.230 26.205 52.610 ;
        RECT 21.065 51.970 21.565 52.060 ;
        RECT 21.055 51.240 21.565 51.970 ;
        RECT 21.295 50.240 21.565 51.240 ;
        RECT 22.205 50.990 22.475 51.940 ;
        RECT 22.205 50.840 22.675 50.990 ;
        RECT 22.205 50.160 22.765 50.840 ;
        RECT 22.285 50.150 22.765 50.160 ;
        RECT 21.575 49.620 22.195 49.980 ;
        RECT 21.615 49.090 22.045 49.620 ;
        RECT 20.165 48.670 22.045 49.090 ;
        RECT 22.535 48.960 22.765 50.150 ;
        RECT 21.615 47.800 22.045 48.670 ;
        RECT 22.455 48.360 22.835 48.960 ;
        RECT 19.325 47.060 20.015 47.770 ;
        RECT 21.435 47.440 22.055 47.800 ;
        RECT 21.135 47.060 21.425 47.250 ;
        RECT 19.325 46.620 21.425 47.060 ;
        RECT 19.325 46.600 20.015 46.620 ;
        RECT 21.135 46.380 21.425 46.620 ;
        RECT 22.055 46.990 22.325 47.240 ;
        RECT 22.535 46.990 22.765 48.360 ;
        RECT 25.355 47.010 25.685 52.030 ;
        RECT 26.405 52.020 27.535 53.240 ;
        RECT 28.895 53.220 29.215 53.240 ;
        RECT 22.055 46.880 22.765 46.990 ;
        RECT 25.345 46.960 25.685 47.010 ;
        RECT 26.235 47.780 27.615 52.020 ;
        RECT 22.055 46.570 22.715 46.880 ;
        RECT 22.055 46.400 22.325 46.570 ;
        RECT 25.345 45.000 25.625 46.960 ;
        RECT 26.235 46.920 26.535 47.780 ;
        RECT 27.315 46.920 27.615 47.780 ;
        RECT 28.165 46.920 28.495 51.990 ;
        RECT 27.565 46.380 28.045 46.760 ;
        RECT 27.665 45.760 27.915 46.380 ;
        RECT 27.565 45.160 27.945 45.760 ;
        RECT 24.825 44.230 25.925 45.000 ;
        RECT 28.215 44.930 28.495 46.920 ;
        RECT 30.525 47.780 31.025 68.580 ;
        RECT 31.365 49.100 31.755 70.610 ;
        RECT 32.155 70.020 33.045 70.750 ;
        RECT 32.255 65.200 32.515 70.020 ;
        RECT 33.895 68.630 36.605 69.480 ;
        RECT 34.095 65.850 36.025 68.630 ;
        RECT 41.725 68.550 42.265 71.780 ;
        RECT 42.565 70.580 42.975 73.220 ;
        RECT 50.055 73.090 52.125 74.370 ;
        RECT 53.150 73.290 55.710 75.820 ;
        RECT 64.900 75.810 65.180 77.710 ;
        RECT 103.990 77.230 104.270 84.740 ;
        RECT 76.140 76.950 104.270 77.230 ;
        RECT 52.675 71.760 53.535 72.600 ;
        RECT 38.995 67.140 40.115 67.820 ;
        RECT 39.275 65.860 39.945 67.140 ;
        RECT 32.655 65.470 37.705 65.850 ;
        RECT 39.065 65.450 40.115 65.860 ;
        RECT 32.255 63.650 32.635 65.200 ;
        RECT 32.375 55.810 32.635 63.650 ;
        RECT 37.685 63.210 37.955 65.250 ;
        RECT 38.815 63.210 39.085 65.210 ;
        RECT 37.685 56.520 39.085 63.210 ;
        RECT 32.285 55.300 32.645 55.810 ;
        RECT 32.265 54.870 32.645 55.300 ;
        RECT 37.685 55.200 37.955 56.520 ;
        RECT 38.815 55.160 39.085 56.520 ;
        RECT 40.085 55.270 40.405 65.200 ;
        RECT 40.085 55.210 40.415 55.270 ;
        RECT 32.265 54.590 32.515 54.870 ;
        RECT 32.065 54.190 36.705 54.590 ;
        RECT 37.605 54.300 38.735 54.310 ;
        RECT 40.095 54.300 40.415 55.210 ;
        RECT 32.265 52.070 32.515 54.190 ;
        RECT 36.965 53.500 37.325 54.120 ;
        RECT 37.045 52.620 37.305 53.500 ;
        RECT 37.585 53.250 40.415 54.300 ;
        RECT 36.875 52.240 37.405 52.620 ;
        RECT 32.265 51.980 32.765 52.070 ;
        RECT 32.255 51.250 32.765 51.980 ;
        RECT 32.495 50.250 32.765 51.250 ;
        RECT 33.405 51.000 33.675 51.950 ;
        RECT 33.405 50.850 33.875 51.000 ;
        RECT 33.405 50.170 33.965 50.850 ;
        RECT 33.485 50.160 33.965 50.170 ;
        RECT 32.775 49.630 33.395 49.990 ;
        RECT 32.815 49.100 33.245 49.630 ;
        RECT 31.365 48.680 33.245 49.100 ;
        RECT 33.735 48.970 33.965 50.160 ;
        RECT 32.815 47.810 33.245 48.680 ;
        RECT 33.655 48.370 34.035 48.970 ;
        RECT 30.525 47.070 31.215 47.780 ;
        RECT 32.635 47.450 33.255 47.810 ;
        RECT 32.335 47.070 32.625 47.260 ;
        RECT 30.525 46.630 32.625 47.070 ;
        RECT 30.525 46.610 31.215 46.630 ;
        RECT 32.335 46.390 32.625 46.630 ;
        RECT 33.255 47.000 33.525 47.250 ;
        RECT 33.735 47.000 33.965 48.370 ;
        RECT 36.555 47.020 36.885 52.040 ;
        RECT 37.605 52.030 38.735 53.250 ;
        RECT 40.095 53.230 40.415 53.250 ;
        RECT 33.255 46.890 33.965 47.000 ;
        RECT 36.545 46.970 36.885 47.020 ;
        RECT 37.435 47.790 38.815 52.030 ;
        RECT 33.255 46.580 33.915 46.890 ;
        RECT 33.255 46.410 33.525 46.580 ;
        RECT 36.545 45.010 36.825 46.970 ;
        RECT 37.435 46.930 37.735 47.790 ;
        RECT 38.515 46.930 38.815 47.790 ;
        RECT 39.365 46.930 39.695 52.000 ;
        RECT 38.765 46.390 39.245 46.770 ;
        RECT 38.865 45.770 39.115 46.390 ;
        RECT 38.765 45.170 39.145 45.770 ;
        RECT 28.215 43.200 28.515 44.930 ;
        RECT 36.025 44.240 37.125 45.010 ;
        RECT 39.415 44.940 39.695 46.930 ;
        RECT 41.745 47.750 42.245 68.550 ;
        RECT 42.585 49.070 42.975 70.580 ;
        RECT 43.375 69.990 44.265 70.720 ;
        RECT 43.475 65.170 43.735 69.990 ;
        RECT 45.115 68.600 47.825 69.450 ;
        RECT 45.315 65.820 47.245 68.600 ;
        RECT 52.975 68.530 53.515 71.760 ;
        RECT 53.815 70.560 54.225 73.290 ;
        RECT 61.475 73.120 63.545 74.400 ;
        RECT 64.400 73.280 66.960 75.810 ;
        RECT 76.140 75.740 76.420 76.950 ;
        RECT 109.970 76.610 110.250 85.420 ;
        RECT 87.580 76.330 110.250 76.610 ;
        RECT 87.580 75.760 87.860 76.330 ;
        RECT 115.950 76.030 116.230 85.700 ;
        RECT 98.850 75.840 116.230 76.030 ;
        RECT 63.895 71.750 64.755 72.590 ;
        RECT 50.215 67.110 51.335 67.790 ;
        RECT 50.495 65.830 51.165 67.110 ;
        RECT 43.875 65.440 48.925 65.820 ;
        RECT 50.285 65.420 51.335 65.830 ;
        RECT 43.475 63.620 43.855 65.170 ;
        RECT 43.595 55.780 43.855 63.620 ;
        RECT 48.905 63.180 49.175 65.220 ;
        RECT 50.035 63.180 50.305 65.180 ;
        RECT 48.905 56.490 50.305 63.180 ;
        RECT 43.505 55.270 43.865 55.780 ;
        RECT 43.485 54.840 43.865 55.270 ;
        RECT 48.905 55.170 49.175 56.490 ;
        RECT 50.035 55.130 50.305 56.490 ;
        RECT 51.305 55.240 51.625 65.170 ;
        RECT 51.305 55.180 51.635 55.240 ;
        RECT 43.485 54.560 43.735 54.840 ;
        RECT 43.285 54.160 47.925 54.560 ;
        RECT 48.825 54.270 49.955 54.280 ;
        RECT 51.315 54.270 51.635 55.180 ;
        RECT 43.485 52.040 43.735 54.160 ;
        RECT 48.185 53.470 48.545 54.090 ;
        RECT 48.265 52.590 48.525 53.470 ;
        RECT 48.805 53.220 51.635 54.270 ;
        RECT 48.095 52.210 48.625 52.590 ;
        RECT 43.485 51.950 43.985 52.040 ;
        RECT 43.475 51.220 43.985 51.950 ;
        RECT 43.715 50.220 43.985 51.220 ;
        RECT 44.625 50.970 44.895 51.920 ;
        RECT 44.625 50.820 45.095 50.970 ;
        RECT 44.625 50.140 45.185 50.820 ;
        RECT 44.705 50.130 45.185 50.140 ;
        RECT 43.995 49.600 44.615 49.960 ;
        RECT 44.035 49.070 44.465 49.600 ;
        RECT 42.585 48.650 44.465 49.070 ;
        RECT 44.955 48.940 45.185 50.130 ;
        RECT 44.035 47.780 44.465 48.650 ;
        RECT 44.875 48.340 45.255 48.940 ;
        RECT 41.745 47.040 42.435 47.750 ;
        RECT 43.855 47.420 44.475 47.780 ;
        RECT 43.555 47.040 43.845 47.230 ;
        RECT 41.745 46.600 43.845 47.040 ;
        RECT 41.745 46.580 42.435 46.600 ;
        RECT 43.555 46.360 43.845 46.600 ;
        RECT 44.475 46.970 44.745 47.220 ;
        RECT 44.955 46.970 45.185 48.340 ;
        RECT 47.775 46.990 48.105 52.010 ;
        RECT 48.825 52.000 49.955 53.220 ;
        RECT 51.315 53.200 51.635 53.220 ;
        RECT 44.475 46.860 45.185 46.970 ;
        RECT 47.765 46.940 48.105 46.990 ;
        RECT 48.655 47.760 50.035 52.000 ;
        RECT 44.475 46.550 45.135 46.860 ;
        RECT 44.475 46.380 44.745 46.550 ;
        RECT 47.765 44.980 48.045 46.940 ;
        RECT 48.655 46.900 48.955 47.760 ;
        RECT 49.735 46.900 50.035 47.760 ;
        RECT 50.585 46.900 50.915 51.970 ;
        RECT 49.985 46.360 50.465 46.740 ;
        RECT 50.085 45.740 50.335 46.360 ;
        RECT 49.985 45.140 50.365 45.740 ;
        RECT 39.415 43.210 39.715 44.940 ;
        RECT 47.245 44.210 48.345 44.980 ;
        RECT 50.635 44.910 50.915 46.900 ;
        RECT 52.995 47.730 53.495 68.530 ;
        RECT 53.835 49.050 54.225 70.560 ;
        RECT 54.625 69.970 55.515 70.700 ;
        RECT 54.725 65.150 54.985 69.970 ;
        RECT 56.365 68.580 59.075 69.430 ;
        RECT 56.565 65.800 58.495 68.580 ;
        RECT 64.195 68.520 64.735 71.750 ;
        RECT 65.035 70.550 65.445 73.280 ;
        RECT 72.585 73.130 74.655 74.410 ;
        RECT 75.550 73.210 78.110 75.740 ;
        RECT 75.135 71.740 75.995 72.580 ;
        RECT 61.465 67.090 62.585 67.770 ;
        RECT 61.745 65.810 62.415 67.090 ;
        RECT 55.125 65.420 60.175 65.800 ;
        RECT 61.535 65.400 62.585 65.810 ;
        RECT 54.725 63.600 55.105 65.150 ;
        RECT 54.845 55.760 55.105 63.600 ;
        RECT 60.155 63.160 60.425 65.200 ;
        RECT 61.285 63.160 61.555 65.160 ;
        RECT 60.155 56.470 61.555 63.160 ;
        RECT 54.755 55.250 55.115 55.760 ;
        RECT 54.735 54.820 55.115 55.250 ;
        RECT 60.155 55.150 60.425 56.470 ;
        RECT 61.285 55.110 61.555 56.470 ;
        RECT 62.555 55.220 62.875 65.150 ;
        RECT 62.555 55.160 62.885 55.220 ;
        RECT 54.735 54.540 54.985 54.820 ;
        RECT 54.535 54.140 59.175 54.540 ;
        RECT 60.075 54.250 61.205 54.260 ;
        RECT 62.565 54.250 62.885 55.160 ;
        RECT 54.735 52.020 54.985 54.140 ;
        RECT 59.435 53.450 59.795 54.070 ;
        RECT 59.515 52.570 59.775 53.450 ;
        RECT 60.055 53.200 62.885 54.250 ;
        RECT 59.345 52.190 59.875 52.570 ;
        RECT 54.735 51.930 55.235 52.020 ;
        RECT 54.725 51.200 55.235 51.930 ;
        RECT 54.965 50.200 55.235 51.200 ;
        RECT 55.875 50.950 56.145 51.900 ;
        RECT 55.875 50.800 56.345 50.950 ;
        RECT 55.875 50.120 56.435 50.800 ;
        RECT 55.955 50.110 56.435 50.120 ;
        RECT 55.245 49.580 55.865 49.940 ;
        RECT 55.285 49.050 55.715 49.580 ;
        RECT 53.835 48.630 55.715 49.050 ;
        RECT 56.205 48.920 56.435 50.110 ;
        RECT 55.285 47.760 55.715 48.630 ;
        RECT 56.125 48.320 56.505 48.920 ;
        RECT 52.995 47.020 53.685 47.730 ;
        RECT 55.105 47.400 55.725 47.760 ;
        RECT 54.805 47.020 55.095 47.210 ;
        RECT 52.995 46.580 55.095 47.020 ;
        RECT 52.995 46.560 53.685 46.580 ;
        RECT 54.805 46.340 55.095 46.580 ;
        RECT 55.725 46.950 55.995 47.200 ;
        RECT 56.205 46.950 56.435 48.320 ;
        RECT 59.025 46.970 59.355 51.990 ;
        RECT 60.075 51.980 61.205 53.200 ;
        RECT 62.565 53.180 62.885 53.200 ;
        RECT 55.725 46.840 56.435 46.950 ;
        RECT 59.015 46.920 59.355 46.970 ;
        RECT 59.905 47.740 61.285 51.980 ;
        RECT 55.725 46.530 56.385 46.840 ;
        RECT 55.725 46.360 55.995 46.530 ;
        RECT 59.015 44.960 59.295 46.920 ;
        RECT 59.905 46.880 60.205 47.740 ;
        RECT 60.985 46.880 61.285 47.740 ;
        RECT 61.835 46.880 62.165 51.950 ;
        RECT 61.235 46.340 61.715 46.720 ;
        RECT 61.335 45.720 61.585 46.340 ;
        RECT 61.235 45.120 61.615 45.720 ;
        RECT 19.865 42.210 21.245 42.780 ;
        RECT 27.495 42.630 28.875 43.200 ;
        RECT 31.145 42.210 32.525 42.780 ;
        RECT 38.695 42.640 40.075 43.210 ;
        RECT 50.635 43.180 50.935 44.910 ;
        RECT 58.495 44.190 59.595 44.960 ;
        RECT 61.885 44.890 62.165 46.880 ;
        RECT 64.215 47.720 64.715 68.520 ;
        RECT 65.055 49.040 65.445 70.550 ;
        RECT 65.845 69.960 66.735 70.690 ;
        RECT 65.945 65.140 66.205 69.960 ;
        RECT 67.585 68.570 70.295 69.420 ;
        RECT 67.785 65.790 69.715 68.570 ;
        RECT 75.435 68.510 75.975 71.740 ;
        RECT 76.275 70.540 76.685 73.210 ;
        RECT 83.855 73.120 85.925 74.400 ;
        RECT 86.850 73.230 89.410 75.760 ;
        RECT 98.150 75.750 116.230 75.840 ;
        RECT 86.385 71.750 87.245 72.590 ;
        RECT 72.685 67.080 73.805 67.760 ;
        RECT 72.965 65.800 73.635 67.080 ;
        RECT 66.345 65.410 71.395 65.790 ;
        RECT 72.755 65.390 73.805 65.800 ;
        RECT 65.945 63.590 66.325 65.140 ;
        RECT 66.065 55.750 66.325 63.590 ;
        RECT 71.375 63.150 71.645 65.190 ;
        RECT 72.505 63.150 72.775 65.150 ;
        RECT 71.375 56.460 72.775 63.150 ;
        RECT 65.975 55.240 66.335 55.750 ;
        RECT 65.955 54.810 66.335 55.240 ;
        RECT 71.375 55.140 71.645 56.460 ;
        RECT 72.505 55.100 72.775 56.460 ;
        RECT 73.775 55.210 74.095 65.140 ;
        RECT 73.775 55.150 74.105 55.210 ;
        RECT 65.955 54.530 66.205 54.810 ;
        RECT 65.755 54.130 70.395 54.530 ;
        RECT 71.295 54.240 72.425 54.250 ;
        RECT 73.785 54.240 74.105 55.150 ;
        RECT 65.955 52.010 66.205 54.130 ;
        RECT 70.655 53.440 71.015 54.060 ;
        RECT 70.735 52.560 70.995 53.440 ;
        RECT 71.275 53.190 74.105 54.240 ;
        RECT 70.565 52.180 71.095 52.560 ;
        RECT 65.955 51.920 66.455 52.010 ;
        RECT 65.945 51.190 66.455 51.920 ;
        RECT 66.185 50.190 66.455 51.190 ;
        RECT 67.095 50.940 67.365 51.890 ;
        RECT 67.095 50.790 67.565 50.940 ;
        RECT 67.095 50.110 67.655 50.790 ;
        RECT 67.175 50.100 67.655 50.110 ;
        RECT 66.465 49.570 67.085 49.930 ;
        RECT 66.505 49.040 66.935 49.570 ;
        RECT 65.055 48.620 66.935 49.040 ;
        RECT 67.425 48.910 67.655 50.100 ;
        RECT 66.505 47.750 66.935 48.620 ;
        RECT 67.345 48.310 67.725 48.910 ;
        RECT 64.215 47.010 64.905 47.720 ;
        RECT 66.325 47.390 66.945 47.750 ;
        RECT 66.025 47.010 66.315 47.200 ;
        RECT 64.215 46.570 66.315 47.010 ;
        RECT 64.215 46.550 64.905 46.570 ;
        RECT 66.025 46.330 66.315 46.570 ;
        RECT 66.945 46.940 67.215 47.190 ;
        RECT 67.425 46.940 67.655 48.310 ;
        RECT 70.245 46.960 70.575 51.980 ;
        RECT 71.295 51.970 72.425 53.190 ;
        RECT 73.785 53.170 74.105 53.190 ;
        RECT 66.945 46.830 67.655 46.940 ;
        RECT 70.235 46.910 70.575 46.960 ;
        RECT 71.125 47.730 72.505 51.970 ;
        RECT 66.945 46.520 67.605 46.830 ;
        RECT 66.945 46.350 67.215 46.520 ;
        RECT 70.235 44.950 70.515 46.910 ;
        RECT 71.125 46.870 71.425 47.730 ;
        RECT 72.205 46.870 72.505 47.730 ;
        RECT 73.055 46.870 73.385 51.940 ;
        RECT 72.455 46.330 72.935 46.710 ;
        RECT 72.555 45.710 72.805 46.330 ;
        RECT 72.455 45.110 72.835 45.710 ;
        RECT 20.225 40.480 20.525 42.210 ;
        RECT 20.245 38.490 20.525 40.480 ;
        RECT 22.815 40.410 23.915 41.180 ;
        RECT 31.505 40.480 31.805 42.210 ;
        RECT 42.435 42.190 43.815 42.760 ;
        RECT 49.915 42.610 51.295 43.180 ;
        RECT 61.885 43.160 62.185 44.890 ;
        RECT 69.715 44.180 70.815 44.950 ;
        RECT 73.105 44.880 73.385 46.870 ;
        RECT 75.455 47.710 75.955 68.510 ;
        RECT 76.295 49.030 76.685 70.540 ;
        RECT 77.085 69.950 77.975 70.680 ;
        RECT 77.185 65.130 77.445 69.950 ;
        RECT 78.825 68.560 81.535 69.410 ;
        RECT 79.025 65.780 80.955 68.560 ;
        RECT 86.685 68.520 87.225 71.750 ;
        RECT 87.525 70.550 87.935 73.230 ;
        RECT 95.045 73.060 97.115 74.340 ;
        RECT 98.150 73.310 100.710 75.750 ;
        RECT 109.390 75.480 111.950 75.560 ;
        RECT 121.930 75.480 122.210 85.700 ;
        RECT 127.550 85.510 128.770 89.380 ;
        RECT 127.910 76.040 128.190 85.510 ;
        RECT 133.380 76.580 136.010 77.880 ;
        RECT 137.240 76.560 139.870 77.860 ;
        RECT 109.390 75.200 122.210 75.480 ;
        RECT 97.665 71.740 98.525 72.580 ;
        RECT 83.925 67.070 85.045 67.750 ;
        RECT 84.205 65.790 84.875 67.070 ;
        RECT 77.585 65.400 82.635 65.780 ;
        RECT 83.995 65.380 85.045 65.790 ;
        RECT 77.185 63.580 77.565 65.130 ;
        RECT 77.305 55.740 77.565 63.580 ;
        RECT 82.615 63.140 82.885 65.180 ;
        RECT 83.745 63.140 84.015 65.140 ;
        RECT 82.615 56.450 84.015 63.140 ;
        RECT 77.215 55.230 77.575 55.740 ;
        RECT 77.195 54.800 77.575 55.230 ;
        RECT 82.615 55.130 82.885 56.450 ;
        RECT 83.745 55.090 84.015 56.450 ;
        RECT 85.015 55.200 85.335 65.130 ;
        RECT 85.015 55.140 85.345 55.200 ;
        RECT 77.195 54.520 77.445 54.800 ;
        RECT 76.995 54.120 81.635 54.520 ;
        RECT 82.535 54.230 83.665 54.240 ;
        RECT 85.025 54.230 85.345 55.140 ;
        RECT 77.195 52.000 77.445 54.120 ;
        RECT 81.895 53.430 82.255 54.050 ;
        RECT 81.975 52.550 82.235 53.430 ;
        RECT 82.515 53.180 85.345 54.230 ;
        RECT 81.805 52.170 82.335 52.550 ;
        RECT 77.195 51.910 77.695 52.000 ;
        RECT 77.185 51.180 77.695 51.910 ;
        RECT 77.425 50.180 77.695 51.180 ;
        RECT 78.335 50.930 78.605 51.880 ;
        RECT 78.335 50.780 78.805 50.930 ;
        RECT 78.335 50.100 78.895 50.780 ;
        RECT 78.415 50.090 78.895 50.100 ;
        RECT 77.705 49.560 78.325 49.920 ;
        RECT 77.745 49.030 78.175 49.560 ;
        RECT 76.295 48.610 78.175 49.030 ;
        RECT 78.665 48.900 78.895 50.090 ;
        RECT 77.745 47.740 78.175 48.610 ;
        RECT 78.585 48.300 78.965 48.900 ;
        RECT 75.455 47.000 76.145 47.710 ;
        RECT 77.565 47.380 78.185 47.740 ;
        RECT 77.265 47.000 77.555 47.190 ;
        RECT 75.455 46.560 77.555 47.000 ;
        RECT 75.455 46.540 76.145 46.560 ;
        RECT 77.265 46.320 77.555 46.560 ;
        RECT 78.185 46.930 78.455 47.180 ;
        RECT 78.665 46.930 78.895 48.300 ;
        RECT 81.485 46.950 81.815 51.970 ;
        RECT 82.535 51.960 83.665 53.180 ;
        RECT 85.025 53.160 85.345 53.180 ;
        RECT 78.185 46.820 78.895 46.930 ;
        RECT 81.475 46.900 81.815 46.950 ;
        RECT 82.365 47.720 83.745 51.960 ;
        RECT 78.185 46.510 78.845 46.820 ;
        RECT 78.185 46.340 78.455 46.510 ;
        RECT 81.475 44.940 81.755 46.900 ;
        RECT 82.365 46.860 82.665 47.720 ;
        RECT 83.445 46.860 83.745 47.720 ;
        RECT 84.295 46.860 84.625 51.930 ;
        RECT 83.695 46.320 84.175 46.700 ;
        RECT 83.795 45.700 84.045 46.320 ;
        RECT 83.695 45.100 84.075 45.700 ;
        RECT 53.655 42.190 55.035 42.760 ;
        RECT 61.165 42.590 62.545 43.160 ;
        RECT 73.105 43.150 73.405 44.880 ;
        RECT 80.955 44.170 82.055 44.940 ;
        RECT 84.345 44.870 84.625 46.860 ;
        RECT 86.705 47.720 87.205 68.520 ;
        RECT 87.545 49.040 87.935 70.550 ;
        RECT 88.335 69.960 89.225 70.690 ;
        RECT 88.435 65.140 88.695 69.960 ;
        RECT 90.075 68.570 92.785 69.420 ;
        RECT 90.275 65.790 92.205 68.570 ;
        RECT 97.965 68.510 98.505 71.740 ;
        RECT 98.805 70.540 99.215 73.310 ;
        RECT 106.455 73.110 108.525 74.390 ;
        RECT 109.390 73.030 111.950 75.200 ;
        RECT 125.760 74.810 128.190 76.040 ;
        RECT 121.290 74.790 128.190 74.810 ;
        RECT 120.600 74.530 128.190 74.790 ;
        RECT 117.655 73.110 119.725 74.390 ;
        RECT 120.600 73.180 128.160 74.530 ;
        RECT 129.505 73.190 131.575 74.470 ;
        RECT 120.600 73.110 126.160 73.180 ;
        RECT 108.935 71.740 109.795 72.580 ;
        RECT 95.175 67.080 96.295 67.760 ;
        RECT 95.455 65.800 96.125 67.080 ;
        RECT 88.835 65.410 93.885 65.790 ;
        RECT 95.245 65.390 96.295 65.800 ;
        RECT 88.435 63.590 88.815 65.140 ;
        RECT 88.555 55.750 88.815 63.590 ;
        RECT 93.865 63.150 94.135 65.190 ;
        RECT 94.995 63.150 95.265 65.150 ;
        RECT 93.865 56.460 95.265 63.150 ;
        RECT 88.465 55.240 88.825 55.750 ;
        RECT 88.445 54.810 88.825 55.240 ;
        RECT 93.865 55.140 94.135 56.460 ;
        RECT 94.995 55.100 95.265 56.460 ;
        RECT 96.265 55.210 96.585 65.140 ;
        RECT 96.265 55.150 96.595 55.210 ;
        RECT 88.445 54.530 88.695 54.810 ;
        RECT 88.245 54.130 92.885 54.530 ;
        RECT 93.785 54.240 94.915 54.250 ;
        RECT 96.275 54.240 96.595 55.150 ;
        RECT 88.445 52.010 88.695 54.130 ;
        RECT 93.145 53.440 93.505 54.060 ;
        RECT 93.225 52.560 93.485 53.440 ;
        RECT 93.765 53.190 96.595 54.240 ;
        RECT 93.055 52.180 93.585 52.560 ;
        RECT 88.445 51.920 88.945 52.010 ;
        RECT 88.435 51.190 88.945 51.920 ;
        RECT 88.675 50.190 88.945 51.190 ;
        RECT 89.585 50.940 89.855 51.890 ;
        RECT 89.585 50.790 90.055 50.940 ;
        RECT 89.585 50.110 90.145 50.790 ;
        RECT 89.665 50.100 90.145 50.110 ;
        RECT 88.955 49.570 89.575 49.930 ;
        RECT 88.995 49.040 89.425 49.570 ;
        RECT 87.545 48.620 89.425 49.040 ;
        RECT 89.915 48.910 90.145 50.100 ;
        RECT 88.995 47.750 89.425 48.620 ;
        RECT 89.835 48.310 90.215 48.910 ;
        RECT 86.705 47.010 87.395 47.720 ;
        RECT 88.815 47.390 89.435 47.750 ;
        RECT 88.515 47.010 88.805 47.200 ;
        RECT 86.705 46.570 88.805 47.010 ;
        RECT 86.705 46.550 87.395 46.570 ;
        RECT 88.515 46.330 88.805 46.570 ;
        RECT 89.435 46.940 89.705 47.190 ;
        RECT 89.915 46.940 90.145 48.310 ;
        RECT 92.735 46.960 93.065 51.980 ;
        RECT 93.785 51.970 94.915 53.190 ;
        RECT 96.275 53.170 96.595 53.190 ;
        RECT 89.435 46.830 90.145 46.940 ;
        RECT 92.725 46.910 93.065 46.960 ;
        RECT 93.615 47.730 94.995 51.970 ;
        RECT 89.435 46.520 90.095 46.830 ;
        RECT 89.435 46.350 89.705 46.520 ;
        RECT 92.725 44.950 93.005 46.910 ;
        RECT 93.615 46.870 93.915 47.730 ;
        RECT 94.695 46.870 94.995 47.730 ;
        RECT 95.545 46.870 95.875 51.940 ;
        RECT 94.945 46.330 95.425 46.710 ;
        RECT 95.045 45.710 95.295 46.330 ;
        RECT 94.945 45.110 95.325 45.710 ;
        RECT 64.855 42.190 66.235 42.760 ;
        RECT 72.385 42.580 73.765 43.150 ;
        RECT 84.345 43.140 84.645 44.870 ;
        RECT 92.205 44.180 93.305 44.950 ;
        RECT 95.595 44.880 95.875 46.870 ;
        RECT 97.985 47.710 98.485 68.510 ;
        RECT 98.825 49.030 99.215 70.540 ;
        RECT 99.615 69.950 100.505 70.680 ;
        RECT 99.715 65.130 99.975 69.950 ;
        RECT 101.355 68.560 104.065 69.410 ;
        RECT 101.555 65.780 103.485 68.560 ;
        RECT 109.235 68.510 109.775 71.740 ;
        RECT 110.075 70.540 110.485 73.030 ;
        RECT 120.185 71.740 121.045 72.580 ;
        RECT 106.455 67.070 107.575 67.750 ;
        RECT 106.735 65.790 107.405 67.070 ;
        RECT 100.115 65.400 105.165 65.780 ;
        RECT 106.525 65.380 107.575 65.790 ;
        RECT 99.715 63.580 100.095 65.130 ;
        RECT 99.835 55.740 100.095 63.580 ;
        RECT 105.145 63.140 105.415 65.180 ;
        RECT 106.275 63.140 106.545 65.140 ;
        RECT 105.145 56.450 106.545 63.140 ;
        RECT 99.745 55.230 100.105 55.740 ;
        RECT 99.725 54.800 100.105 55.230 ;
        RECT 105.145 55.130 105.415 56.450 ;
        RECT 106.275 55.090 106.545 56.450 ;
        RECT 107.545 55.200 107.865 65.130 ;
        RECT 107.545 55.140 107.875 55.200 ;
        RECT 99.725 54.520 99.975 54.800 ;
        RECT 99.525 54.120 104.165 54.520 ;
        RECT 105.065 54.230 106.195 54.240 ;
        RECT 107.555 54.230 107.875 55.140 ;
        RECT 99.725 52.000 99.975 54.120 ;
        RECT 104.425 53.430 104.785 54.050 ;
        RECT 104.505 52.550 104.765 53.430 ;
        RECT 105.045 53.180 107.875 54.230 ;
        RECT 104.335 52.170 104.865 52.550 ;
        RECT 99.725 51.910 100.225 52.000 ;
        RECT 99.715 51.180 100.225 51.910 ;
        RECT 99.955 50.180 100.225 51.180 ;
        RECT 100.865 50.930 101.135 51.880 ;
        RECT 100.865 50.780 101.335 50.930 ;
        RECT 100.865 50.100 101.425 50.780 ;
        RECT 100.945 50.090 101.425 50.100 ;
        RECT 100.235 49.560 100.855 49.920 ;
        RECT 100.275 49.030 100.705 49.560 ;
        RECT 98.825 48.610 100.705 49.030 ;
        RECT 101.195 48.900 101.425 50.090 ;
        RECT 100.275 47.740 100.705 48.610 ;
        RECT 101.115 48.300 101.495 48.900 ;
        RECT 97.985 47.000 98.675 47.710 ;
        RECT 100.095 47.380 100.715 47.740 ;
        RECT 99.795 47.000 100.085 47.190 ;
        RECT 97.985 46.560 100.085 47.000 ;
        RECT 97.985 46.540 98.675 46.560 ;
        RECT 99.795 46.320 100.085 46.560 ;
        RECT 100.715 46.930 100.985 47.180 ;
        RECT 101.195 46.930 101.425 48.300 ;
        RECT 104.015 46.950 104.345 51.970 ;
        RECT 105.065 51.960 106.195 53.180 ;
        RECT 107.555 53.160 107.875 53.180 ;
        RECT 100.715 46.820 101.425 46.930 ;
        RECT 104.005 46.900 104.345 46.950 ;
        RECT 104.895 47.720 106.275 51.960 ;
        RECT 100.715 46.510 101.375 46.820 ;
        RECT 100.715 46.340 100.985 46.510 ;
        RECT 104.005 44.940 104.285 46.900 ;
        RECT 104.895 46.860 105.195 47.720 ;
        RECT 105.975 46.860 106.275 47.720 ;
        RECT 106.825 46.860 107.155 51.930 ;
        RECT 106.225 46.320 106.705 46.700 ;
        RECT 106.325 45.700 106.575 46.320 ;
        RECT 106.225 45.100 106.605 45.700 ;
        RECT 95.595 43.150 95.895 44.880 ;
        RECT 103.485 44.170 104.585 44.940 ;
        RECT 106.875 44.870 107.155 46.860 ;
        RECT 109.255 47.710 109.755 68.510 ;
        RECT 110.095 49.030 110.485 70.540 ;
        RECT 110.885 69.950 111.775 70.680 ;
        RECT 110.985 65.130 111.245 69.950 ;
        RECT 112.625 68.560 115.335 69.410 ;
        RECT 112.825 65.780 114.755 68.560 ;
        RECT 120.485 68.510 121.025 71.740 ;
        RECT 121.325 70.540 121.735 73.110 ;
        RECT 132.925 70.810 133.225 70.900 ;
        RECT 117.725 67.070 118.845 67.750 ;
        RECT 118.005 65.790 118.675 67.070 ;
        RECT 111.385 65.400 116.435 65.780 ;
        RECT 117.795 65.380 118.845 65.790 ;
        RECT 110.985 63.580 111.365 65.130 ;
        RECT 111.105 55.740 111.365 63.580 ;
        RECT 116.415 63.140 116.685 65.180 ;
        RECT 117.545 63.140 117.815 65.140 ;
        RECT 116.415 56.450 117.815 63.140 ;
        RECT 111.015 55.230 111.375 55.740 ;
        RECT 110.995 54.800 111.375 55.230 ;
        RECT 116.415 55.130 116.685 56.450 ;
        RECT 117.545 55.090 117.815 56.450 ;
        RECT 118.815 55.200 119.135 65.130 ;
        RECT 118.815 55.140 119.145 55.200 ;
        RECT 110.995 54.520 111.245 54.800 ;
        RECT 110.795 54.120 115.435 54.520 ;
        RECT 116.335 54.230 117.465 54.240 ;
        RECT 118.825 54.230 119.145 55.140 ;
        RECT 110.995 52.000 111.245 54.120 ;
        RECT 115.695 53.430 116.055 54.050 ;
        RECT 115.775 52.550 116.035 53.430 ;
        RECT 116.315 53.180 119.145 54.230 ;
        RECT 115.605 52.170 116.135 52.550 ;
        RECT 110.995 51.910 111.495 52.000 ;
        RECT 110.985 51.180 111.495 51.910 ;
        RECT 111.225 50.180 111.495 51.180 ;
        RECT 112.135 50.930 112.405 51.880 ;
        RECT 112.135 50.780 112.605 50.930 ;
        RECT 112.135 50.100 112.695 50.780 ;
        RECT 112.215 50.090 112.695 50.100 ;
        RECT 111.505 49.560 112.125 49.920 ;
        RECT 111.545 49.030 111.975 49.560 ;
        RECT 110.095 48.610 111.975 49.030 ;
        RECT 112.465 48.900 112.695 50.090 ;
        RECT 111.545 47.740 111.975 48.610 ;
        RECT 112.385 48.300 112.765 48.900 ;
        RECT 109.255 47.000 109.945 47.710 ;
        RECT 111.365 47.380 111.985 47.740 ;
        RECT 111.065 47.000 111.355 47.190 ;
        RECT 109.255 46.560 111.355 47.000 ;
        RECT 109.255 46.540 109.945 46.560 ;
        RECT 111.065 46.320 111.355 46.560 ;
        RECT 111.985 46.930 112.255 47.180 ;
        RECT 112.465 46.930 112.695 48.300 ;
        RECT 115.285 46.950 115.615 51.970 ;
        RECT 116.335 51.960 117.465 53.180 ;
        RECT 118.825 53.160 119.145 53.180 ;
        RECT 111.985 46.820 112.695 46.930 ;
        RECT 115.275 46.900 115.615 46.950 ;
        RECT 116.165 47.720 117.545 51.960 ;
        RECT 111.985 46.510 112.645 46.820 ;
        RECT 111.985 46.340 112.255 46.510 ;
        RECT 115.275 44.940 115.555 46.900 ;
        RECT 116.165 46.860 116.465 47.720 ;
        RECT 117.245 46.860 117.545 47.720 ;
        RECT 118.095 46.860 118.425 51.930 ;
        RECT 117.495 46.320 117.975 46.700 ;
        RECT 117.595 45.700 117.845 46.320 ;
        RECT 117.495 45.100 117.875 45.700 ;
        RECT 20.795 39.650 21.175 40.250 ;
        RECT 20.825 39.030 21.075 39.650 ;
        RECT 20.695 38.650 21.175 39.030 ;
        RECT 20.245 33.420 20.575 38.490 ;
        RECT 21.125 37.630 21.425 38.490 ;
        RECT 22.205 37.630 22.505 38.490 ;
        RECT 23.115 38.450 23.395 40.410 ;
        RECT 26.415 38.840 26.685 39.010 ;
        RECT 26.025 38.530 26.685 38.840 ;
        RECT 21.125 33.390 22.505 37.630 ;
        RECT 23.055 38.400 23.395 38.450 ;
        RECT 25.975 38.420 26.685 38.530 ;
        RECT 19.525 32.170 19.845 32.190 ;
        RECT 21.205 32.170 22.335 33.390 ;
        RECT 23.055 33.380 23.385 38.400 ;
        RECT 25.975 37.050 26.205 38.420 ;
        RECT 26.415 38.170 26.685 38.420 ;
        RECT 27.315 38.790 27.605 39.030 ;
        RECT 28.725 38.790 29.415 38.810 ;
        RECT 27.315 38.350 29.415 38.790 ;
        RECT 27.315 38.160 27.605 38.350 ;
        RECT 26.685 37.610 27.305 37.970 ;
        RECT 28.725 37.640 29.415 38.350 ;
        RECT 25.905 36.450 26.285 37.050 ;
        RECT 26.695 36.740 27.125 37.610 ;
        RECT 25.975 35.260 26.205 36.450 ;
        RECT 26.695 36.320 28.575 36.740 ;
        RECT 26.695 35.790 27.125 36.320 ;
        RECT 26.545 35.430 27.165 35.790 ;
        RECT 25.975 35.250 26.455 35.260 ;
        RECT 25.975 34.570 26.535 35.250 ;
        RECT 26.065 34.420 26.535 34.570 ;
        RECT 26.265 33.470 26.535 34.420 ;
        RECT 27.175 34.170 27.445 35.170 ;
        RECT 27.175 33.440 27.685 34.170 ;
        RECT 27.175 33.350 27.675 33.440 ;
        RECT 22.535 32.800 23.065 33.180 ;
        RECT 19.525 31.120 22.355 32.170 ;
        RECT 22.635 31.920 22.895 32.800 ;
        RECT 22.615 31.300 22.975 31.920 ;
        RECT 27.425 31.230 27.675 33.350 ;
        RECT 19.525 30.210 19.845 31.120 ;
        RECT 21.205 31.110 22.335 31.120 ;
        RECT 23.235 30.830 27.875 31.230 ;
        RECT 27.425 30.550 27.675 30.830 ;
        RECT 19.525 30.150 19.855 30.210 ;
        RECT 19.535 20.220 19.855 30.150 ;
        RECT 20.855 28.900 21.125 30.260 ;
        RECT 21.985 28.900 22.255 30.220 ;
        RECT 27.295 30.120 27.675 30.550 ;
        RECT 27.295 29.610 27.655 30.120 ;
        RECT 20.855 22.210 22.255 28.900 ;
        RECT 20.855 20.210 21.125 22.210 ;
        RECT 21.985 20.170 22.255 22.210 ;
        RECT 27.305 21.770 27.565 29.610 ;
        RECT 27.305 20.220 27.685 21.770 ;
        RECT 19.825 19.560 20.875 19.970 ;
        RECT 22.235 19.570 27.285 19.950 ;
        RECT 19.995 18.280 20.665 19.560 ;
        RECT 19.825 17.600 20.945 18.280 ;
        RECT 23.915 16.790 25.845 19.570 ;
        RECT 23.335 15.940 26.045 16.790 ;
        RECT 27.425 15.400 27.685 20.220 ;
        RECT 26.895 14.670 27.785 15.400 ;
        RECT 28.185 14.810 28.575 36.320 ;
        RECT 28.915 16.840 29.415 37.640 ;
        RECT 31.525 38.490 31.805 40.480 ;
        RECT 34.095 40.410 35.195 41.180 ;
        RECT 42.795 40.460 43.095 42.190 ;
        RECT 32.075 39.650 32.455 40.250 ;
        RECT 32.105 39.030 32.355 39.650 ;
        RECT 31.975 38.650 32.455 39.030 ;
        RECT 31.525 33.420 31.855 38.490 ;
        RECT 32.405 37.630 32.705 38.490 ;
        RECT 33.485 37.630 33.785 38.490 ;
        RECT 34.395 38.450 34.675 40.410 ;
        RECT 37.695 38.840 37.965 39.010 ;
        RECT 37.305 38.530 37.965 38.840 ;
        RECT 32.405 33.390 33.785 37.630 ;
        RECT 34.335 38.400 34.675 38.450 ;
        RECT 37.255 38.420 37.965 38.530 ;
        RECT 30.805 32.170 31.125 32.190 ;
        RECT 32.485 32.170 33.615 33.390 ;
        RECT 34.335 33.380 34.665 38.400 ;
        RECT 37.255 37.050 37.485 38.420 ;
        RECT 37.695 38.170 37.965 38.420 ;
        RECT 38.595 38.790 38.885 39.030 ;
        RECT 40.005 38.790 40.695 38.810 ;
        RECT 38.595 38.350 40.695 38.790 ;
        RECT 38.595 38.160 38.885 38.350 ;
        RECT 37.965 37.610 38.585 37.970 ;
        RECT 40.005 37.640 40.695 38.350 ;
        RECT 37.185 36.450 37.565 37.050 ;
        RECT 37.975 36.740 38.405 37.610 ;
        RECT 37.255 35.260 37.485 36.450 ;
        RECT 37.975 36.320 39.855 36.740 ;
        RECT 37.975 35.790 38.405 36.320 ;
        RECT 37.825 35.430 38.445 35.790 ;
        RECT 37.255 35.250 37.735 35.260 ;
        RECT 37.255 34.570 37.815 35.250 ;
        RECT 37.345 34.420 37.815 34.570 ;
        RECT 37.545 33.470 37.815 34.420 ;
        RECT 38.455 34.170 38.725 35.170 ;
        RECT 38.455 33.440 38.965 34.170 ;
        RECT 38.455 33.350 38.955 33.440 ;
        RECT 33.815 32.800 34.345 33.180 ;
        RECT 30.805 31.120 33.635 32.170 ;
        RECT 33.915 31.920 34.175 32.800 ;
        RECT 33.895 31.300 34.255 31.920 ;
        RECT 38.705 31.230 38.955 33.350 ;
        RECT 30.805 30.210 31.125 31.120 ;
        RECT 32.485 31.110 33.615 31.120 ;
        RECT 34.515 30.830 39.155 31.230 ;
        RECT 38.705 30.550 38.955 30.830 ;
        RECT 30.805 30.150 31.135 30.210 ;
        RECT 30.815 20.220 31.135 30.150 ;
        RECT 32.135 28.900 32.405 30.260 ;
        RECT 33.265 28.900 33.535 30.220 ;
        RECT 38.575 30.120 38.955 30.550 ;
        RECT 38.575 29.610 38.935 30.120 ;
        RECT 32.135 22.210 33.535 28.900 ;
        RECT 32.135 20.210 32.405 22.210 ;
        RECT 33.265 20.170 33.535 22.210 ;
        RECT 38.585 21.770 38.845 29.610 ;
        RECT 38.585 20.220 38.965 21.770 ;
        RECT 31.105 19.560 32.155 19.970 ;
        RECT 33.515 19.570 38.565 19.950 ;
        RECT 31.275 18.280 31.945 19.560 ;
        RECT 31.105 17.600 32.225 18.280 ;
        RECT 28.185 12.290 28.595 14.810 ;
        RECT 28.895 13.610 29.435 16.840 ;
        RECT 35.195 16.790 37.125 19.570 ;
        RECT 34.615 15.940 37.325 16.790 ;
        RECT 38.705 15.400 38.965 20.220 ;
        RECT 38.175 14.670 39.065 15.400 ;
        RECT 39.465 14.810 39.855 36.320 ;
        RECT 40.195 16.840 40.695 37.640 ;
        RECT 42.815 38.470 43.095 40.460 ;
        RECT 45.385 40.390 46.485 41.160 ;
        RECT 54.015 40.460 54.315 42.190 ;
        RECT 43.365 39.630 43.745 40.230 ;
        RECT 43.395 39.010 43.645 39.630 ;
        RECT 43.265 38.630 43.745 39.010 ;
        RECT 42.815 33.400 43.145 38.470 ;
        RECT 43.695 37.610 43.995 38.470 ;
        RECT 44.775 37.610 45.075 38.470 ;
        RECT 45.685 38.430 45.965 40.390 ;
        RECT 48.985 38.820 49.255 38.990 ;
        RECT 48.595 38.510 49.255 38.820 ;
        RECT 43.695 33.370 45.075 37.610 ;
        RECT 45.625 38.380 45.965 38.430 ;
        RECT 48.545 38.400 49.255 38.510 ;
        RECT 42.095 32.150 42.415 32.170 ;
        RECT 43.775 32.150 44.905 33.370 ;
        RECT 45.625 33.360 45.955 38.380 ;
        RECT 48.545 37.030 48.775 38.400 ;
        RECT 48.985 38.150 49.255 38.400 ;
        RECT 49.885 38.770 50.175 39.010 ;
        RECT 51.295 38.770 51.985 38.790 ;
        RECT 49.885 38.330 51.985 38.770 ;
        RECT 49.885 38.140 50.175 38.330 ;
        RECT 49.255 37.590 49.875 37.950 ;
        RECT 51.295 37.620 51.985 38.330 ;
        RECT 48.475 36.430 48.855 37.030 ;
        RECT 49.265 36.720 49.695 37.590 ;
        RECT 48.545 35.240 48.775 36.430 ;
        RECT 49.265 36.300 51.145 36.720 ;
        RECT 49.265 35.770 49.695 36.300 ;
        RECT 49.115 35.410 49.735 35.770 ;
        RECT 48.545 35.230 49.025 35.240 ;
        RECT 48.545 34.550 49.105 35.230 ;
        RECT 48.635 34.400 49.105 34.550 ;
        RECT 48.835 33.450 49.105 34.400 ;
        RECT 49.745 34.150 50.015 35.150 ;
        RECT 49.745 33.420 50.255 34.150 ;
        RECT 49.745 33.330 50.245 33.420 ;
        RECT 45.105 32.780 45.635 33.160 ;
        RECT 42.095 31.100 44.925 32.150 ;
        RECT 45.205 31.900 45.465 32.780 ;
        RECT 45.185 31.280 45.545 31.900 ;
        RECT 49.995 31.210 50.245 33.330 ;
        RECT 42.095 30.190 42.415 31.100 ;
        RECT 43.775 31.090 44.905 31.100 ;
        RECT 45.805 30.810 50.445 31.210 ;
        RECT 49.995 30.530 50.245 30.810 ;
        RECT 42.095 30.130 42.425 30.190 ;
        RECT 42.105 20.200 42.425 30.130 ;
        RECT 43.425 28.880 43.695 30.240 ;
        RECT 44.555 28.880 44.825 30.200 ;
        RECT 49.865 30.100 50.245 30.530 ;
        RECT 49.865 29.590 50.225 30.100 ;
        RECT 43.425 22.190 44.825 28.880 ;
        RECT 43.425 20.190 43.695 22.190 ;
        RECT 44.555 20.150 44.825 22.190 ;
        RECT 49.875 21.750 50.135 29.590 ;
        RECT 49.875 20.200 50.255 21.750 ;
        RECT 42.395 19.540 43.445 19.950 ;
        RECT 44.805 19.550 49.855 19.930 ;
        RECT 42.565 18.260 43.235 19.540 ;
        RECT 42.395 17.580 43.515 18.260 ;
        RECT 28.875 12.770 29.735 13.610 ;
        RECT 28.185 11.950 30.415 12.290 ;
        RECT 39.465 11.990 39.875 14.810 ;
        RECT 40.175 13.610 40.715 16.840 ;
        RECT 46.485 16.770 48.415 19.550 ;
        RECT 45.905 15.920 48.615 16.770 ;
        RECT 49.995 15.380 50.255 20.200 ;
        RECT 49.465 14.650 50.355 15.380 ;
        RECT 50.755 14.790 51.145 36.300 ;
        RECT 51.485 16.820 51.985 37.620 ;
        RECT 54.035 38.470 54.315 40.460 ;
        RECT 56.605 40.390 57.705 41.160 ;
        RECT 65.215 40.460 65.515 42.190 ;
        RECT 76.145 42.180 77.525 42.750 ;
        RECT 83.625 42.570 85.005 43.140 ;
        RECT 87.385 42.200 88.765 42.770 ;
        RECT 94.875 42.580 96.255 43.150 ;
        RECT 106.875 43.140 107.175 44.870 ;
        RECT 114.755 44.170 115.855 44.940 ;
        RECT 118.145 44.870 118.425 46.860 ;
        RECT 120.505 47.710 121.005 68.510 ;
        RECT 121.345 49.030 121.735 70.540 ;
        RECT 122.135 69.950 123.025 70.680 ;
        RECT 132.615 70.040 134.265 70.810 ;
        RECT 122.235 65.130 122.495 69.950 ;
        RECT 123.875 68.560 126.585 69.410 ;
        RECT 124.075 65.780 126.005 68.560 ;
        RECT 128.975 67.070 130.095 67.750 ;
        RECT 129.255 65.790 129.925 67.070 ;
        RECT 122.635 65.400 127.685 65.780 ;
        RECT 129.045 65.380 130.095 65.790 ;
        RECT 132.925 65.180 133.225 70.040 ;
        RECT 137.675 68.690 139.075 69.460 ;
        RECT 138.385 65.740 138.645 68.690 ;
        RECT 149.410 68.420 150.690 69.620 ;
        RECT 149.480 65.810 150.640 68.420 ;
        RECT 133.365 65.380 138.645 65.740 ;
        RECT 122.235 63.580 122.615 65.130 ;
        RECT 122.355 55.740 122.615 63.580 ;
        RECT 127.665 63.140 127.935 65.180 ;
        RECT 128.795 63.140 129.065 65.140 ;
        RECT 127.665 56.450 129.065 63.140 ;
        RECT 122.265 55.230 122.625 55.740 ;
        RECT 122.245 54.800 122.625 55.230 ;
        RECT 127.665 55.130 127.935 56.450 ;
        RECT 128.795 55.090 129.065 56.450 ;
        RECT 130.065 55.200 130.385 65.130 ;
        RECT 132.925 61.010 133.355 65.180 ;
        RECT 138.385 65.150 138.645 65.380 ;
        RECT 138.385 64.770 138.675 65.150 ;
        RECT 130.065 55.140 130.395 55.200 ;
        RECT 133.055 55.190 133.355 61.010 ;
        RECT 122.245 54.520 122.495 54.800 ;
        RECT 122.045 54.120 126.685 54.520 ;
        RECT 127.585 54.230 128.715 54.240 ;
        RECT 130.075 54.230 130.395 55.140 ;
        RECT 138.395 55.080 138.675 64.770 ;
        RECT 149.390 64.610 150.670 65.810 ;
        RECT 122.245 52.000 122.495 54.120 ;
        RECT 126.945 53.430 127.305 54.050 ;
        RECT 127.025 52.550 127.285 53.430 ;
        RECT 127.565 53.180 130.395 54.230 ;
        RECT 126.855 52.170 127.385 52.550 ;
        RECT 122.245 51.910 122.745 52.000 ;
        RECT 122.235 51.180 122.745 51.910 ;
        RECT 122.475 50.180 122.745 51.180 ;
        RECT 123.385 50.930 123.655 51.880 ;
        RECT 123.385 50.780 123.855 50.930 ;
        RECT 123.385 50.100 123.945 50.780 ;
        RECT 123.465 50.090 123.945 50.100 ;
        RECT 122.755 49.560 123.375 49.920 ;
        RECT 122.795 49.030 123.225 49.560 ;
        RECT 121.345 48.610 123.225 49.030 ;
        RECT 123.715 48.900 123.945 50.090 ;
        RECT 122.795 47.740 123.225 48.610 ;
        RECT 123.635 48.300 124.015 48.900 ;
        RECT 120.505 47.000 121.195 47.710 ;
        RECT 122.615 47.380 123.235 47.740 ;
        RECT 122.315 47.000 122.605 47.190 ;
        RECT 120.505 46.560 122.605 47.000 ;
        RECT 120.505 46.540 121.195 46.560 ;
        RECT 122.315 46.320 122.605 46.560 ;
        RECT 123.235 46.930 123.505 47.180 ;
        RECT 123.715 46.930 123.945 48.300 ;
        RECT 126.535 46.950 126.865 51.970 ;
        RECT 127.585 51.960 128.715 53.180 ;
        RECT 130.075 53.160 130.395 53.180 ;
        RECT 123.235 46.820 123.945 46.930 ;
        RECT 126.525 46.900 126.865 46.950 ;
        RECT 127.415 47.720 128.795 51.960 ;
        RECT 123.235 46.510 123.895 46.820 ;
        RECT 123.235 46.340 123.505 46.510 ;
        RECT 126.525 44.940 126.805 46.900 ;
        RECT 127.415 46.860 127.715 47.720 ;
        RECT 128.495 46.860 128.795 47.720 ;
        RECT 129.345 46.860 129.675 51.930 ;
        RECT 128.745 46.320 129.225 46.700 ;
        RECT 128.845 45.700 129.095 46.320 ;
        RECT 128.745 45.100 129.125 45.700 ;
        RECT 118.145 43.140 118.445 44.870 ;
        RECT 126.005 44.170 127.105 44.940 ;
        RECT 129.395 44.870 129.675 46.860 ;
        RECT 129.395 43.140 129.695 44.870 ;
        RECT 98.595 42.220 99.975 42.790 ;
        RECT 106.155 42.570 107.535 43.140 ;
        RECT 109.795 42.260 111.175 42.830 ;
        RECT 117.425 42.570 118.805 43.140 ;
        RECT 121.005 42.280 122.385 42.850 ;
        RECT 128.675 42.570 130.055 43.140 ;
        RECT 54.585 39.630 54.965 40.230 ;
        RECT 54.615 39.010 54.865 39.630 ;
        RECT 54.485 38.630 54.965 39.010 ;
        RECT 54.035 33.400 54.365 38.470 ;
        RECT 54.915 37.610 55.215 38.470 ;
        RECT 55.995 37.610 56.295 38.470 ;
        RECT 56.905 38.430 57.185 40.390 ;
        RECT 60.205 38.820 60.475 38.990 ;
        RECT 59.815 38.510 60.475 38.820 ;
        RECT 54.915 33.370 56.295 37.610 ;
        RECT 56.845 38.380 57.185 38.430 ;
        RECT 59.765 38.400 60.475 38.510 ;
        RECT 53.315 32.150 53.635 32.170 ;
        RECT 54.995 32.150 56.125 33.370 ;
        RECT 56.845 33.360 57.175 38.380 ;
        RECT 59.765 37.030 59.995 38.400 ;
        RECT 60.205 38.150 60.475 38.400 ;
        RECT 61.105 38.770 61.395 39.010 ;
        RECT 62.515 38.770 63.205 38.790 ;
        RECT 61.105 38.330 63.205 38.770 ;
        RECT 61.105 38.140 61.395 38.330 ;
        RECT 60.475 37.590 61.095 37.950 ;
        RECT 62.515 37.620 63.205 38.330 ;
        RECT 59.695 36.430 60.075 37.030 ;
        RECT 60.485 36.720 60.915 37.590 ;
        RECT 59.765 35.240 59.995 36.430 ;
        RECT 60.485 36.300 62.365 36.720 ;
        RECT 60.485 35.770 60.915 36.300 ;
        RECT 60.335 35.410 60.955 35.770 ;
        RECT 59.765 35.230 60.245 35.240 ;
        RECT 59.765 34.550 60.325 35.230 ;
        RECT 59.855 34.400 60.325 34.550 ;
        RECT 60.055 33.450 60.325 34.400 ;
        RECT 60.965 34.150 61.235 35.150 ;
        RECT 60.965 33.420 61.475 34.150 ;
        RECT 60.965 33.330 61.465 33.420 ;
        RECT 56.325 32.780 56.855 33.160 ;
        RECT 53.315 31.100 56.145 32.150 ;
        RECT 56.425 31.900 56.685 32.780 ;
        RECT 56.405 31.280 56.765 31.900 ;
        RECT 61.215 31.210 61.465 33.330 ;
        RECT 53.315 30.190 53.635 31.100 ;
        RECT 54.995 31.090 56.125 31.100 ;
        RECT 57.025 30.810 61.665 31.210 ;
        RECT 61.215 30.530 61.465 30.810 ;
        RECT 53.315 30.130 53.645 30.190 ;
        RECT 53.325 20.200 53.645 30.130 ;
        RECT 54.645 28.880 54.915 30.240 ;
        RECT 55.775 28.880 56.045 30.200 ;
        RECT 61.085 30.100 61.465 30.530 ;
        RECT 61.085 29.590 61.445 30.100 ;
        RECT 54.645 22.190 56.045 28.880 ;
        RECT 54.645 20.190 54.915 22.190 ;
        RECT 55.775 20.150 56.045 22.190 ;
        RECT 61.095 21.750 61.355 29.590 ;
        RECT 61.095 20.200 61.475 21.750 ;
        RECT 53.615 19.540 54.665 19.950 ;
        RECT 56.025 19.550 61.075 19.930 ;
        RECT 53.785 18.260 54.455 19.540 ;
        RECT 53.615 17.580 54.735 18.260 ;
        RECT 40.155 12.770 41.015 13.610 ;
        RECT 50.755 12.170 51.165 14.790 ;
        RECT 51.465 13.590 52.005 16.820 ;
        RECT 57.705 16.770 59.635 19.550 ;
        RECT 57.125 15.920 59.835 16.770 ;
        RECT 61.215 15.380 61.475 20.200 ;
        RECT 60.685 14.650 61.575 15.380 ;
        RECT 61.975 14.790 62.365 36.300 ;
        RECT 62.705 16.820 63.205 37.620 ;
        RECT 65.235 38.470 65.515 40.460 ;
        RECT 67.805 40.390 68.905 41.160 ;
        RECT 76.505 40.450 76.805 42.180 ;
        RECT 65.785 39.630 66.165 40.230 ;
        RECT 65.815 39.010 66.065 39.630 ;
        RECT 65.685 38.630 66.165 39.010 ;
        RECT 65.235 33.400 65.565 38.470 ;
        RECT 66.115 37.610 66.415 38.470 ;
        RECT 67.195 37.610 67.495 38.470 ;
        RECT 68.105 38.430 68.385 40.390 ;
        RECT 71.405 38.820 71.675 38.990 ;
        RECT 71.015 38.510 71.675 38.820 ;
        RECT 66.115 33.370 67.495 37.610 ;
        RECT 68.045 38.380 68.385 38.430 ;
        RECT 70.965 38.400 71.675 38.510 ;
        RECT 64.515 32.150 64.835 32.170 ;
        RECT 66.195 32.150 67.325 33.370 ;
        RECT 68.045 33.360 68.375 38.380 ;
        RECT 70.965 37.030 71.195 38.400 ;
        RECT 71.405 38.150 71.675 38.400 ;
        RECT 72.305 38.770 72.595 39.010 ;
        RECT 73.715 38.770 74.405 38.790 ;
        RECT 72.305 38.330 74.405 38.770 ;
        RECT 72.305 38.140 72.595 38.330 ;
        RECT 71.675 37.590 72.295 37.950 ;
        RECT 73.715 37.620 74.405 38.330 ;
        RECT 70.895 36.430 71.275 37.030 ;
        RECT 71.685 36.720 72.115 37.590 ;
        RECT 70.965 35.240 71.195 36.430 ;
        RECT 71.685 36.300 73.565 36.720 ;
        RECT 71.685 35.770 72.115 36.300 ;
        RECT 71.535 35.410 72.155 35.770 ;
        RECT 70.965 35.230 71.445 35.240 ;
        RECT 70.965 34.550 71.525 35.230 ;
        RECT 71.055 34.400 71.525 34.550 ;
        RECT 71.255 33.450 71.525 34.400 ;
        RECT 72.165 34.150 72.435 35.150 ;
        RECT 72.165 33.420 72.675 34.150 ;
        RECT 72.165 33.330 72.665 33.420 ;
        RECT 67.525 32.780 68.055 33.160 ;
        RECT 64.515 31.100 67.345 32.150 ;
        RECT 67.625 31.900 67.885 32.780 ;
        RECT 67.605 31.280 67.965 31.900 ;
        RECT 72.415 31.210 72.665 33.330 ;
        RECT 64.515 30.190 64.835 31.100 ;
        RECT 66.195 31.090 67.325 31.100 ;
        RECT 68.225 30.810 72.865 31.210 ;
        RECT 72.415 30.530 72.665 30.810 ;
        RECT 64.515 30.130 64.845 30.190 ;
        RECT 64.525 20.200 64.845 30.130 ;
        RECT 65.845 28.880 66.115 30.240 ;
        RECT 66.975 28.880 67.245 30.200 ;
        RECT 72.285 30.100 72.665 30.530 ;
        RECT 72.285 29.590 72.645 30.100 ;
        RECT 65.845 22.190 67.245 28.880 ;
        RECT 65.845 20.190 66.115 22.190 ;
        RECT 66.975 20.150 67.245 22.190 ;
        RECT 72.295 21.750 72.555 29.590 ;
        RECT 72.295 20.200 72.675 21.750 ;
        RECT 64.815 19.540 65.865 19.950 ;
        RECT 67.225 19.550 72.275 19.930 ;
        RECT 64.985 18.260 65.655 19.540 ;
        RECT 64.815 17.580 65.935 18.260 ;
        RECT 51.445 12.750 52.305 13.590 ;
        RECT 27.865 11.130 30.415 11.950 ;
        RECT 28.395 11.090 30.415 11.130 ;
        RECT 39.115 10.980 41.565 11.990 ;
        RECT 50.335 10.970 52.355 12.170 ;
        RECT 61.975 12.160 62.385 14.790 ;
        RECT 62.685 13.590 63.225 16.820 ;
        RECT 68.905 16.770 70.835 19.550 ;
        RECT 68.325 15.920 71.035 16.770 ;
        RECT 72.415 15.380 72.675 20.200 ;
        RECT 71.885 14.650 72.775 15.380 ;
        RECT 73.175 14.790 73.565 36.300 ;
        RECT 73.905 16.820 74.405 37.620 ;
        RECT 76.525 38.460 76.805 40.450 ;
        RECT 79.095 40.380 80.195 41.150 ;
        RECT 87.745 40.470 88.045 42.200 ;
        RECT 77.075 39.620 77.455 40.220 ;
        RECT 77.105 39.000 77.355 39.620 ;
        RECT 76.975 38.620 77.455 39.000 ;
        RECT 76.525 33.390 76.855 38.460 ;
        RECT 77.405 37.600 77.705 38.460 ;
        RECT 78.485 37.600 78.785 38.460 ;
        RECT 79.395 38.420 79.675 40.380 ;
        RECT 82.695 38.810 82.965 38.980 ;
        RECT 82.305 38.500 82.965 38.810 ;
        RECT 77.405 33.360 78.785 37.600 ;
        RECT 79.335 38.370 79.675 38.420 ;
        RECT 82.255 38.390 82.965 38.500 ;
        RECT 75.805 32.140 76.125 32.160 ;
        RECT 77.485 32.140 78.615 33.360 ;
        RECT 79.335 33.350 79.665 38.370 ;
        RECT 82.255 37.020 82.485 38.390 ;
        RECT 82.695 38.140 82.965 38.390 ;
        RECT 83.595 38.760 83.885 39.000 ;
        RECT 85.005 38.760 85.695 38.780 ;
        RECT 83.595 38.320 85.695 38.760 ;
        RECT 83.595 38.130 83.885 38.320 ;
        RECT 82.965 37.580 83.585 37.940 ;
        RECT 85.005 37.610 85.695 38.320 ;
        RECT 82.185 36.420 82.565 37.020 ;
        RECT 82.975 36.710 83.405 37.580 ;
        RECT 82.255 35.230 82.485 36.420 ;
        RECT 82.975 36.290 84.855 36.710 ;
        RECT 82.975 35.760 83.405 36.290 ;
        RECT 82.825 35.400 83.445 35.760 ;
        RECT 82.255 35.220 82.735 35.230 ;
        RECT 82.255 34.540 82.815 35.220 ;
        RECT 82.345 34.390 82.815 34.540 ;
        RECT 82.545 33.440 82.815 34.390 ;
        RECT 83.455 34.140 83.725 35.140 ;
        RECT 83.455 33.410 83.965 34.140 ;
        RECT 83.455 33.320 83.955 33.410 ;
        RECT 78.815 32.770 79.345 33.150 ;
        RECT 75.805 31.090 78.635 32.140 ;
        RECT 78.915 31.890 79.175 32.770 ;
        RECT 78.895 31.270 79.255 31.890 ;
        RECT 83.705 31.200 83.955 33.320 ;
        RECT 75.805 30.180 76.125 31.090 ;
        RECT 77.485 31.080 78.615 31.090 ;
        RECT 79.515 30.800 84.155 31.200 ;
        RECT 83.705 30.520 83.955 30.800 ;
        RECT 75.805 30.120 76.135 30.180 ;
        RECT 75.815 20.190 76.135 30.120 ;
        RECT 77.135 28.870 77.405 30.230 ;
        RECT 78.265 28.870 78.535 30.190 ;
        RECT 83.575 30.090 83.955 30.520 ;
        RECT 83.575 29.580 83.935 30.090 ;
        RECT 77.135 22.180 78.535 28.870 ;
        RECT 77.135 20.180 77.405 22.180 ;
        RECT 78.265 20.140 78.535 22.180 ;
        RECT 83.585 21.740 83.845 29.580 ;
        RECT 83.585 20.190 83.965 21.740 ;
        RECT 76.105 19.530 77.155 19.940 ;
        RECT 78.515 19.540 83.565 19.920 ;
        RECT 76.275 18.250 76.945 19.530 ;
        RECT 76.105 17.570 77.225 18.250 ;
        RECT 62.665 12.750 63.525 13.590 ;
        RECT 73.175 12.190 73.585 14.790 ;
        RECT 73.885 13.590 74.425 16.820 ;
        RECT 80.195 16.760 82.125 19.540 ;
        RECT 79.615 15.910 82.325 16.760 ;
        RECT 83.705 15.370 83.965 20.190 ;
        RECT 83.175 14.640 84.065 15.370 ;
        RECT 84.465 14.780 84.855 36.290 ;
        RECT 85.195 16.810 85.695 37.610 ;
        RECT 87.765 38.480 88.045 40.470 ;
        RECT 90.335 40.400 91.435 41.170 ;
        RECT 98.955 40.490 99.255 42.220 ;
        RECT 88.315 39.640 88.695 40.240 ;
        RECT 88.345 39.020 88.595 39.640 ;
        RECT 88.215 38.640 88.695 39.020 ;
        RECT 87.765 33.410 88.095 38.480 ;
        RECT 88.645 37.620 88.945 38.480 ;
        RECT 89.725 37.620 90.025 38.480 ;
        RECT 90.635 38.440 90.915 40.400 ;
        RECT 93.935 38.830 94.205 39.000 ;
        RECT 93.545 38.520 94.205 38.830 ;
        RECT 88.645 33.380 90.025 37.620 ;
        RECT 90.575 38.390 90.915 38.440 ;
        RECT 93.495 38.410 94.205 38.520 ;
        RECT 87.045 32.160 87.365 32.180 ;
        RECT 88.725 32.160 89.855 33.380 ;
        RECT 90.575 33.370 90.905 38.390 ;
        RECT 93.495 37.040 93.725 38.410 ;
        RECT 93.935 38.160 94.205 38.410 ;
        RECT 94.835 38.780 95.125 39.020 ;
        RECT 96.245 38.780 96.935 38.800 ;
        RECT 94.835 38.340 96.935 38.780 ;
        RECT 94.835 38.150 95.125 38.340 ;
        RECT 94.205 37.600 94.825 37.960 ;
        RECT 96.245 37.630 96.935 38.340 ;
        RECT 93.425 36.440 93.805 37.040 ;
        RECT 94.215 36.730 94.645 37.600 ;
        RECT 93.495 35.250 93.725 36.440 ;
        RECT 94.215 36.310 96.095 36.730 ;
        RECT 94.215 35.780 94.645 36.310 ;
        RECT 94.065 35.420 94.685 35.780 ;
        RECT 93.495 35.240 93.975 35.250 ;
        RECT 93.495 34.560 94.055 35.240 ;
        RECT 93.585 34.410 94.055 34.560 ;
        RECT 93.785 33.460 94.055 34.410 ;
        RECT 94.695 34.160 94.965 35.160 ;
        RECT 94.695 33.430 95.205 34.160 ;
        RECT 94.695 33.340 95.195 33.430 ;
        RECT 90.055 32.790 90.585 33.170 ;
        RECT 87.045 31.110 89.875 32.160 ;
        RECT 90.155 31.910 90.415 32.790 ;
        RECT 90.135 31.290 90.495 31.910 ;
        RECT 94.945 31.220 95.195 33.340 ;
        RECT 87.045 30.200 87.365 31.110 ;
        RECT 88.725 31.100 89.855 31.110 ;
        RECT 90.755 30.820 95.395 31.220 ;
        RECT 94.945 30.540 95.195 30.820 ;
        RECT 87.045 30.140 87.375 30.200 ;
        RECT 87.055 20.210 87.375 30.140 ;
        RECT 88.375 28.890 88.645 30.250 ;
        RECT 89.505 28.890 89.775 30.210 ;
        RECT 94.815 30.110 95.195 30.540 ;
        RECT 94.815 29.600 95.175 30.110 ;
        RECT 88.375 22.200 89.775 28.890 ;
        RECT 88.375 20.200 88.645 22.200 ;
        RECT 89.505 20.160 89.775 22.200 ;
        RECT 94.825 21.760 95.085 29.600 ;
        RECT 94.825 20.210 95.205 21.760 ;
        RECT 87.345 19.550 88.395 19.960 ;
        RECT 89.755 19.560 94.805 19.940 ;
        RECT 87.515 18.270 88.185 19.550 ;
        RECT 87.345 17.590 88.465 18.270 ;
        RECT 73.865 12.750 74.725 13.590 ;
        RECT 61.415 10.960 63.435 12.160 ;
        RECT 72.725 10.990 74.745 12.190 ;
        RECT 84.465 12.180 84.875 14.780 ;
        RECT 85.175 13.580 85.715 16.810 ;
        RECT 91.435 16.780 93.365 19.560 ;
        RECT 90.855 15.930 93.565 16.780 ;
        RECT 94.945 15.390 95.205 20.210 ;
        RECT 94.415 14.660 95.305 15.390 ;
        RECT 95.705 14.800 96.095 36.310 ;
        RECT 96.435 16.830 96.935 37.630 ;
        RECT 98.975 38.500 99.255 40.490 ;
        RECT 101.545 40.420 102.645 41.190 ;
        RECT 110.155 40.530 110.455 42.260 ;
        RECT 99.525 39.660 99.905 40.260 ;
        RECT 99.555 39.040 99.805 39.660 ;
        RECT 99.425 38.660 99.905 39.040 ;
        RECT 98.975 33.430 99.305 38.500 ;
        RECT 99.855 37.640 100.155 38.500 ;
        RECT 100.935 37.640 101.235 38.500 ;
        RECT 101.845 38.460 102.125 40.420 ;
        RECT 105.145 38.850 105.415 39.020 ;
        RECT 104.755 38.540 105.415 38.850 ;
        RECT 99.855 33.400 101.235 37.640 ;
        RECT 101.785 38.410 102.125 38.460 ;
        RECT 104.705 38.430 105.415 38.540 ;
        RECT 98.255 32.180 98.575 32.200 ;
        RECT 99.935 32.180 101.065 33.400 ;
        RECT 101.785 33.390 102.115 38.410 ;
        RECT 104.705 37.060 104.935 38.430 ;
        RECT 105.145 38.180 105.415 38.430 ;
        RECT 106.045 38.800 106.335 39.040 ;
        RECT 107.455 38.800 108.145 38.820 ;
        RECT 106.045 38.360 108.145 38.800 ;
        RECT 106.045 38.170 106.335 38.360 ;
        RECT 105.415 37.620 106.035 37.980 ;
        RECT 107.455 37.650 108.145 38.360 ;
        RECT 104.635 36.460 105.015 37.060 ;
        RECT 105.425 36.750 105.855 37.620 ;
        RECT 104.705 35.270 104.935 36.460 ;
        RECT 105.425 36.330 107.305 36.750 ;
        RECT 105.425 35.800 105.855 36.330 ;
        RECT 105.275 35.440 105.895 35.800 ;
        RECT 104.705 35.260 105.185 35.270 ;
        RECT 104.705 34.580 105.265 35.260 ;
        RECT 104.795 34.430 105.265 34.580 ;
        RECT 104.995 33.480 105.265 34.430 ;
        RECT 105.905 34.180 106.175 35.180 ;
        RECT 105.905 33.450 106.415 34.180 ;
        RECT 105.905 33.360 106.405 33.450 ;
        RECT 101.265 32.810 101.795 33.190 ;
        RECT 98.255 31.130 101.085 32.180 ;
        RECT 101.365 31.930 101.625 32.810 ;
        RECT 101.345 31.310 101.705 31.930 ;
        RECT 106.155 31.240 106.405 33.360 ;
        RECT 98.255 30.220 98.575 31.130 ;
        RECT 99.935 31.120 101.065 31.130 ;
        RECT 101.965 30.840 106.605 31.240 ;
        RECT 106.155 30.560 106.405 30.840 ;
        RECT 98.255 30.160 98.585 30.220 ;
        RECT 98.265 20.230 98.585 30.160 ;
        RECT 99.585 28.910 99.855 30.270 ;
        RECT 100.715 28.910 100.985 30.230 ;
        RECT 106.025 30.130 106.405 30.560 ;
        RECT 106.025 29.620 106.385 30.130 ;
        RECT 99.585 22.220 100.985 28.910 ;
        RECT 99.585 20.220 99.855 22.220 ;
        RECT 100.715 20.180 100.985 22.220 ;
        RECT 106.035 21.780 106.295 29.620 ;
        RECT 106.035 20.230 106.415 21.780 ;
        RECT 98.555 19.570 99.605 19.980 ;
        RECT 100.965 19.580 106.015 19.960 ;
        RECT 98.725 18.290 99.395 19.570 ;
        RECT 98.555 17.610 99.675 18.290 ;
        RECT 85.155 12.740 86.015 13.580 ;
        RECT 95.705 12.180 96.115 14.800 ;
        RECT 96.415 13.600 96.955 16.830 ;
        RECT 102.645 16.800 104.575 19.580 ;
        RECT 102.065 15.950 104.775 16.800 ;
        RECT 106.155 15.410 106.415 20.230 ;
        RECT 105.625 14.680 106.515 15.410 ;
        RECT 106.915 14.820 107.305 36.330 ;
        RECT 107.645 16.850 108.145 37.650 ;
        RECT 110.175 38.540 110.455 40.530 ;
        RECT 112.745 40.460 113.845 41.230 ;
        RECT 121.365 40.550 121.665 42.280 ;
        RECT 142.880 42.020 144.100 43.390 ;
        RECT 110.725 39.700 111.105 40.300 ;
        RECT 110.755 39.080 111.005 39.700 ;
        RECT 110.625 38.700 111.105 39.080 ;
        RECT 110.175 33.470 110.505 38.540 ;
        RECT 111.055 37.680 111.355 38.540 ;
        RECT 112.135 37.680 112.435 38.540 ;
        RECT 113.045 38.500 113.325 40.460 ;
        RECT 116.345 38.890 116.615 39.060 ;
        RECT 115.955 38.580 116.615 38.890 ;
        RECT 111.055 33.440 112.435 37.680 ;
        RECT 112.985 38.450 113.325 38.500 ;
        RECT 115.905 38.470 116.615 38.580 ;
        RECT 109.455 32.220 109.775 32.240 ;
        RECT 111.135 32.220 112.265 33.440 ;
        RECT 112.985 33.430 113.315 38.450 ;
        RECT 115.905 37.100 116.135 38.470 ;
        RECT 116.345 38.220 116.615 38.470 ;
        RECT 117.245 38.840 117.535 39.080 ;
        RECT 118.655 38.840 119.345 38.860 ;
        RECT 117.245 38.400 119.345 38.840 ;
        RECT 117.245 38.210 117.535 38.400 ;
        RECT 116.615 37.660 117.235 38.020 ;
        RECT 118.655 37.690 119.345 38.400 ;
        RECT 115.835 36.500 116.215 37.100 ;
        RECT 116.625 36.790 117.055 37.660 ;
        RECT 115.905 35.310 116.135 36.500 ;
        RECT 116.625 36.370 118.505 36.790 ;
        RECT 116.625 35.840 117.055 36.370 ;
        RECT 116.475 35.480 117.095 35.840 ;
        RECT 115.905 35.300 116.385 35.310 ;
        RECT 115.905 34.620 116.465 35.300 ;
        RECT 115.995 34.470 116.465 34.620 ;
        RECT 116.195 33.520 116.465 34.470 ;
        RECT 117.105 34.220 117.375 35.220 ;
        RECT 117.105 33.490 117.615 34.220 ;
        RECT 117.105 33.400 117.605 33.490 ;
        RECT 112.465 32.850 112.995 33.230 ;
        RECT 109.455 31.170 112.285 32.220 ;
        RECT 112.565 31.970 112.825 32.850 ;
        RECT 112.545 31.350 112.905 31.970 ;
        RECT 117.355 31.280 117.605 33.400 ;
        RECT 109.455 30.260 109.775 31.170 ;
        RECT 111.135 31.160 112.265 31.170 ;
        RECT 113.165 30.880 117.805 31.280 ;
        RECT 117.355 30.600 117.605 30.880 ;
        RECT 109.455 30.200 109.785 30.260 ;
        RECT 109.465 20.270 109.785 30.200 ;
        RECT 110.785 28.950 111.055 30.310 ;
        RECT 111.915 28.950 112.185 30.270 ;
        RECT 117.225 30.170 117.605 30.600 ;
        RECT 117.225 29.660 117.585 30.170 ;
        RECT 110.785 22.260 112.185 28.950 ;
        RECT 110.785 20.260 111.055 22.260 ;
        RECT 111.915 20.220 112.185 22.260 ;
        RECT 117.235 21.820 117.495 29.660 ;
        RECT 117.235 20.270 117.615 21.820 ;
        RECT 109.755 19.610 110.805 20.020 ;
        RECT 112.165 19.620 117.215 20.000 ;
        RECT 109.925 18.330 110.595 19.610 ;
        RECT 109.755 17.650 110.875 18.330 ;
        RECT 96.395 12.760 97.255 13.600 ;
        RECT 106.915 12.230 107.325 14.820 ;
        RECT 107.625 13.620 108.165 16.850 ;
        RECT 113.845 16.840 115.775 19.620 ;
        RECT 113.265 15.990 115.975 16.840 ;
        RECT 117.355 15.450 117.615 20.270 ;
        RECT 116.825 14.720 117.715 15.450 ;
        RECT 118.115 14.860 118.505 36.370 ;
        RECT 118.845 16.890 119.345 37.690 ;
        RECT 121.385 38.560 121.665 40.550 ;
        RECT 123.955 40.480 125.055 41.250 ;
        RECT 121.935 39.720 122.315 40.320 ;
        RECT 121.965 39.100 122.215 39.720 ;
        RECT 121.835 38.720 122.315 39.100 ;
        RECT 121.385 33.490 121.715 38.560 ;
        RECT 122.265 37.700 122.565 38.560 ;
        RECT 123.345 37.700 123.645 38.560 ;
        RECT 124.255 38.520 124.535 40.480 ;
        RECT 127.555 38.910 127.825 39.080 ;
        RECT 127.165 38.600 127.825 38.910 ;
        RECT 122.265 33.460 123.645 37.700 ;
        RECT 124.195 38.470 124.535 38.520 ;
        RECT 127.115 38.490 127.825 38.600 ;
        RECT 120.665 32.240 120.985 32.260 ;
        RECT 122.345 32.240 123.475 33.460 ;
        RECT 124.195 33.450 124.525 38.470 ;
        RECT 127.115 37.120 127.345 38.490 ;
        RECT 127.555 38.240 127.825 38.490 ;
        RECT 128.455 38.860 128.745 39.100 ;
        RECT 142.940 38.950 144.100 42.020 ;
        RECT 129.865 38.860 130.555 38.880 ;
        RECT 128.455 38.420 130.555 38.860 ;
        RECT 128.455 38.230 128.745 38.420 ;
        RECT 127.825 37.680 128.445 38.040 ;
        RECT 129.865 37.710 130.555 38.420 ;
        RECT 127.045 36.520 127.425 37.120 ;
        RECT 127.835 36.810 128.265 37.680 ;
        RECT 127.115 35.330 127.345 36.520 ;
        RECT 127.835 36.390 129.715 36.810 ;
        RECT 127.835 35.860 128.265 36.390 ;
        RECT 127.685 35.500 128.305 35.860 ;
        RECT 127.115 35.320 127.595 35.330 ;
        RECT 127.115 34.640 127.675 35.320 ;
        RECT 127.205 34.490 127.675 34.640 ;
        RECT 127.405 33.540 127.675 34.490 ;
        RECT 128.315 34.240 128.585 35.240 ;
        RECT 128.315 33.510 128.825 34.240 ;
        RECT 128.315 33.420 128.815 33.510 ;
        RECT 123.675 32.870 124.205 33.250 ;
        RECT 120.665 31.190 123.495 32.240 ;
        RECT 123.775 31.990 124.035 32.870 ;
        RECT 123.755 31.370 124.115 31.990 ;
        RECT 128.565 31.300 128.815 33.420 ;
        RECT 120.665 30.280 120.985 31.190 ;
        RECT 122.345 31.180 123.475 31.190 ;
        RECT 124.375 30.900 129.015 31.300 ;
        RECT 128.565 30.620 128.815 30.900 ;
        RECT 120.665 30.220 120.995 30.280 ;
        RECT 120.675 20.290 120.995 30.220 ;
        RECT 121.995 28.970 122.265 30.330 ;
        RECT 123.125 28.970 123.395 30.290 ;
        RECT 128.435 30.190 128.815 30.620 ;
        RECT 128.435 29.680 128.795 30.190 ;
        RECT 121.995 22.280 123.395 28.970 ;
        RECT 121.995 20.280 122.265 22.280 ;
        RECT 123.125 20.240 123.395 22.280 ;
        RECT 128.445 21.840 128.705 29.680 ;
        RECT 128.445 20.290 128.825 21.840 ;
        RECT 120.965 19.630 122.015 20.040 ;
        RECT 123.375 19.640 128.425 20.020 ;
        RECT 121.135 18.350 121.805 19.630 ;
        RECT 120.965 17.670 122.085 18.350 ;
        RECT 107.605 12.780 108.465 13.620 ;
        RECT 118.115 12.230 118.525 14.860 ;
        RECT 118.825 13.660 119.365 16.890 ;
        RECT 125.055 16.860 126.985 19.640 ;
        RECT 124.475 16.010 127.185 16.860 ;
        RECT 128.565 15.470 128.825 20.290 ;
        RECT 128.035 14.740 128.925 15.470 ;
        RECT 129.325 14.880 129.715 36.390 ;
        RECT 130.055 16.910 130.555 37.710 ;
        RECT 142.900 37.580 144.120 38.950 ;
        RECT 132.395 24.340 132.705 30.230 ;
        RECT 132.195 20.120 132.705 24.340 ;
        RECT 118.805 12.820 119.665 13.660 ;
        RECT 129.325 12.260 129.735 14.880 ;
        RECT 130.035 13.680 130.575 16.910 ;
        RECT 132.195 15.510 132.505 20.120 ;
        RECT 137.715 19.980 138.005 30.170 ;
        RECT 132.685 19.590 138.005 19.980 ;
        RECT 137.715 16.940 138.005 19.590 ;
        RECT 142.940 17.940 144.090 19.160 ;
        RECT 145.080 18.760 146.200 18.930 ;
        RECT 137.395 15.890 138.295 16.940 ;
        RECT 137.715 15.720 138.005 15.890 ;
        RECT 131.975 14.270 132.735 15.510 ;
        RECT 142.940 15.090 144.050 17.940 ;
        RECT 142.900 13.870 144.050 15.090 ;
        RECT 145.070 14.920 146.200 18.760 ;
        RECT 145.030 13.970 146.200 14.920 ;
        RECT 145.030 13.900 146.150 13.970 ;
        RECT 130.015 12.840 130.875 13.680 ;
        RECT 83.845 10.980 85.865 12.180 ;
        RECT 95.145 10.980 97.165 12.180 ;
        RECT 106.335 11.030 108.355 12.230 ;
        RECT 117.565 11.030 119.585 12.230 ;
        RECT 128.865 11.060 130.885 12.260 ;
        RECT 74.340 0.110 75.630 1.460 ;
        RECT 93.550 0.180 94.840 1.530 ;
        RECT 112.950 0.310 114.240 1.660 ;
        RECT 131.850 0.380 133.490 1.930 ;
        RECT 151.650 0.250 152.920 1.470 ;
      LAYER met3 ;
        RECT 135.340 223.855 136.790 225.205 ;
        RECT 138.130 223.785 139.580 225.135 ;
        RECT 143.180 223.815 144.630 225.165 ;
        RECT 46.830 211.125 48.810 211.455 ;
        RECT 76.830 211.125 78.810 211.455 ;
        RECT 106.830 211.125 108.810 211.455 ;
        RECT 31.830 208.405 33.810 208.735 ;
        RECT 61.830 208.405 63.810 208.735 ;
        RECT 91.830 208.405 93.810 208.735 ;
        RECT 121.830 208.405 123.810 208.735 ;
        RECT 46.830 205.685 48.810 206.015 ;
        RECT 76.830 205.685 78.810 206.015 ;
        RECT 106.830 205.685 108.810 206.015 ;
        RECT 31.830 202.965 33.810 203.295 ;
        RECT 61.830 202.965 63.810 203.295 ;
        RECT 91.830 202.965 93.810 203.295 ;
        RECT 121.830 202.965 123.810 203.295 ;
        RECT 46.830 200.245 48.810 200.575 ;
        RECT 76.830 200.245 78.810 200.575 ;
        RECT 106.830 200.245 108.810 200.575 ;
        RECT 31.830 197.525 33.810 197.855 ;
        RECT 61.830 197.525 63.810 197.855 ;
        RECT 91.830 197.525 93.810 197.855 ;
        RECT 121.830 197.525 123.810 197.855 ;
        RECT 46.830 194.805 48.810 195.135 ;
        RECT 76.830 194.805 78.810 195.135 ;
        RECT 106.830 194.805 108.810 195.135 ;
        RECT 78.665 192.740 78.995 192.755 ;
        RECT 79.330 192.740 79.710 192.750 ;
        RECT 78.665 192.440 79.710 192.740 ;
        RECT 78.665 192.425 78.995 192.440 ;
        RECT 79.330 192.430 79.710 192.440 ;
        RECT 31.830 192.085 33.810 192.415 ;
        RECT 61.830 192.085 63.810 192.415 ;
        RECT 91.830 192.085 93.810 192.415 ;
        RECT 121.830 192.085 123.810 192.415 ;
        RECT 46.830 189.365 48.810 189.695 ;
        RECT 76.830 189.365 78.810 189.695 ;
        RECT 106.830 189.365 108.810 189.695 ;
        RECT 31.830 186.645 33.810 186.975 ;
        RECT 61.830 186.645 63.810 186.975 ;
        RECT 91.830 186.645 93.810 186.975 ;
        RECT 121.830 186.645 123.810 186.975 ;
        RECT 40.485 185.940 40.815 185.955 ;
        RECT 50.605 185.940 50.935 185.955 ;
        RECT 80.045 185.940 80.375 185.955 ;
        RECT 40.485 185.640 80.375 185.940 ;
        RECT 40.485 185.625 40.815 185.640 ;
        RECT 50.605 185.625 50.935 185.640 ;
        RECT 80.045 185.625 80.375 185.640 ;
        RECT 40.945 185.260 41.275 185.275 ;
        RECT 48.765 185.260 49.095 185.275 ;
        RECT 40.945 184.960 49.095 185.260 ;
        RECT 40.945 184.945 41.275 184.960 ;
        RECT 48.765 184.945 49.095 184.960 ;
        RECT 67.625 185.260 67.955 185.275 ;
        RECT 85.105 185.270 85.435 185.275 ;
        RECT 84.850 185.260 85.435 185.270 ;
        RECT 67.625 184.960 85.640 185.260 ;
        RECT 67.625 184.945 67.955 184.960 ;
        RECT 84.850 184.950 85.435 184.960 ;
        RECT 85.105 184.945 85.435 184.950 ;
        RECT 81.425 184.580 81.755 184.595 ;
        RECT 82.090 184.580 82.470 184.590 ;
        RECT 81.425 184.280 82.470 184.580 ;
        RECT 81.425 184.265 81.755 184.280 ;
        RECT 82.090 184.270 82.470 184.280 ;
        RECT 46.830 183.925 48.810 184.255 ;
        RECT 76.830 183.925 78.810 184.255 ;
        RECT 106.830 183.925 108.810 184.255 ;
        RECT 80.045 181.870 80.375 181.875 ;
        RECT 80.045 181.860 80.630 181.870 ;
        RECT 79.820 181.560 80.630 181.860 ;
        RECT 80.045 181.550 80.630 181.560 ;
        RECT 83.010 181.860 83.390 181.870 ;
        RECT 83.725 181.860 84.055 181.875 ;
        RECT 83.010 181.560 84.055 181.860 ;
        RECT 83.010 181.550 83.390 181.560 ;
        RECT 80.045 181.545 80.375 181.550 ;
        RECT 83.725 181.545 84.055 181.560 ;
        RECT 31.830 181.205 33.810 181.535 ;
        RECT 61.830 181.205 63.810 181.535 ;
        RECT 91.830 181.205 93.810 181.535 ;
        RECT 121.830 181.205 123.810 181.535 ;
        RECT 40.025 180.500 40.355 180.515 ;
        RECT 49.225 180.500 49.555 180.515 ;
        RECT 40.025 180.200 49.555 180.500 ;
        RECT 40.025 180.185 40.355 180.200 ;
        RECT 49.225 180.185 49.555 180.200 ;
        RECT 51.065 180.500 51.395 180.515 ;
        RECT 75.445 180.500 75.775 180.515 ;
        RECT 51.065 180.200 75.775 180.500 ;
        RECT 51.065 180.185 51.395 180.200 ;
        RECT 75.445 180.185 75.775 180.200 ;
        RECT 49.685 179.820 50.015 179.835 ;
        RECT 58.885 179.820 59.215 179.835 ;
        RECT 49.685 179.520 59.215 179.820 ;
        RECT 49.685 179.505 50.015 179.520 ;
        RECT 58.885 179.505 59.215 179.520 ;
        RECT 46.830 178.485 48.810 178.815 ;
        RECT 76.830 178.485 78.810 178.815 ;
        RECT 106.830 178.485 108.810 178.815 ;
        RECT 130.645 178.460 130.975 178.475 ;
        RECT 131.340 178.460 133.340 178.610 ;
        RECT 130.645 178.160 133.340 178.460 ;
        RECT 130.645 178.145 130.975 178.160 ;
        RECT 131.340 178.010 133.340 178.160 ;
        RECT 31.830 175.765 33.810 176.095 ;
        RECT 61.830 175.765 63.810 176.095 ;
        RECT 91.830 175.765 93.810 176.095 ;
        RECT 121.830 175.765 123.810 176.095 ;
        RECT 79.125 175.060 79.455 175.075 ;
        RECT 123.745 175.060 124.075 175.075 ;
        RECT 79.125 174.760 124.075 175.060 ;
        RECT 79.125 174.745 79.455 174.760 ;
        RECT 123.745 174.745 124.075 174.760 ;
        RECT 46.830 173.045 48.810 173.375 ;
        RECT 76.830 173.045 78.810 173.375 ;
        RECT 106.830 173.045 108.810 173.375 ;
        RECT 84.850 173.020 85.230 173.030 ;
        RECT 90.165 173.020 90.495 173.035 ;
        RECT 84.850 172.720 90.495 173.020 ;
        RECT 84.850 172.710 85.230 172.720 ;
        RECT 90.165 172.705 90.495 172.720 ;
        RECT 31.830 170.325 33.810 170.655 ;
        RECT 61.830 170.325 63.810 170.655 ;
        RECT 91.830 170.325 93.810 170.655 ;
        RECT 121.830 170.325 123.810 170.655 ;
        RECT 129.240 170.585 133.810 172.125 ;
        RECT 47.845 168.940 48.175 168.955 ;
        RECT 53.825 168.940 54.155 168.955 ;
        RECT 54.745 168.940 55.075 168.955 ;
        RECT 47.845 168.640 55.075 168.940 ;
        RECT 47.845 168.625 48.175 168.640 ;
        RECT 53.825 168.625 54.155 168.640 ;
        RECT 54.745 168.625 55.075 168.640 ;
        RECT 55.665 168.260 55.995 168.275 ;
        RECT 56.330 168.260 56.710 168.270 ;
        RECT 55.665 167.960 56.710 168.260 ;
        RECT 55.665 167.945 55.995 167.960 ;
        RECT 56.330 167.950 56.710 167.960 ;
        RECT 46.830 167.605 48.810 167.935 ;
        RECT 76.830 167.605 78.810 167.935 ;
        RECT 106.830 167.605 108.810 167.935 ;
        RECT 61.185 167.580 61.515 167.595 ;
        RECT 60.970 167.265 61.515 167.580 ;
        RECT 60.970 166.910 61.270 167.265 ;
        RECT 60.930 166.900 61.310 166.910 ;
        RECT 73.145 166.900 73.475 166.915 ;
        RECT 60.930 166.600 73.475 166.900 ;
        RECT 60.930 166.590 61.310 166.600 ;
        RECT 73.145 166.585 73.475 166.600 ;
        RECT 103.505 166.900 103.835 166.915 ;
        RECT 112.705 166.900 113.035 166.915 ;
        RECT 103.505 166.600 113.035 166.900 ;
        RECT 103.505 166.585 103.835 166.600 ;
        RECT 112.705 166.585 113.035 166.600 ;
        RECT 41.865 166.220 42.195 166.235 ;
        RECT 50.605 166.220 50.935 166.235 ;
        RECT 72.225 166.220 72.555 166.235 ;
        RECT 41.865 165.920 72.555 166.220 ;
        RECT 41.865 165.905 42.195 165.920 ;
        RECT 50.605 165.905 50.935 165.920 ;
        RECT 72.225 165.905 72.555 165.920 ;
        RECT 31.830 164.885 33.810 165.215 ;
        RECT 61.830 164.885 63.810 165.215 ;
        RECT 91.830 164.885 93.810 165.215 ;
        RECT 121.830 164.885 123.810 165.215 ;
        RECT 81.425 164.180 81.755 164.195 ;
        RECT 84.185 164.180 84.515 164.195 ;
        RECT 81.425 163.880 84.515 164.180 ;
        RECT 81.425 163.865 81.755 163.880 ;
        RECT 84.185 163.865 84.515 163.880 ;
        RECT 105.345 164.180 105.675 164.195 ;
        RECT 107.645 164.180 107.975 164.195 ;
        RECT 113.165 164.180 113.495 164.195 ;
        RECT 105.345 163.880 113.495 164.180 ;
        RECT 105.345 163.865 105.675 163.880 ;
        RECT 107.645 163.865 107.975 163.880 ;
        RECT 113.165 163.865 113.495 163.880 ;
        RECT 57.045 163.500 57.375 163.515 ;
        RECT 57.965 163.500 58.295 163.515 ;
        RECT 57.045 163.200 58.295 163.500 ;
        RECT 57.045 163.185 57.375 163.200 ;
        RECT 57.965 163.185 58.295 163.200 ;
        RECT 64.865 163.500 65.195 163.515 ;
        RECT 69.465 163.500 69.795 163.515 ;
        RECT 76.365 163.500 76.695 163.515 ;
        RECT 64.865 163.200 76.695 163.500 ;
        RECT 64.865 163.185 65.195 163.200 ;
        RECT 69.465 163.185 69.795 163.200 ;
        RECT 76.365 163.185 76.695 163.200 ;
        RECT 107.185 163.500 107.515 163.515 ;
        RECT 110.865 163.500 111.195 163.515 ;
        RECT 107.185 163.200 111.195 163.500 ;
        RECT 107.185 163.185 107.515 163.200 ;
        RECT 110.865 163.185 111.195 163.200 ;
        RECT 112.705 163.500 113.035 163.515 ;
        RECT 116.845 163.500 117.175 163.515 ;
        RECT 112.705 163.200 117.175 163.500 ;
        RECT 112.705 163.185 113.035 163.200 ;
        RECT 116.845 163.185 117.175 163.200 ;
        RECT 52.905 162.820 53.235 162.835 ;
        RECT 59.805 162.820 60.135 162.835 ;
        RECT 52.905 162.520 60.135 162.820 ;
        RECT 52.905 162.505 53.235 162.520 ;
        RECT 59.805 162.505 60.135 162.520 ;
        RECT 46.830 162.165 48.810 162.495 ;
        RECT 76.830 162.165 78.810 162.495 ;
        RECT 106.830 162.165 108.810 162.495 ;
        RECT 58.425 162.140 58.755 162.155 ;
        RECT 59.090 162.140 59.470 162.150 ;
        RECT 58.425 161.840 59.470 162.140 ;
        RECT 58.425 161.825 58.755 161.840 ;
        RECT 59.090 161.830 59.470 161.840 ;
        RECT 48.305 161.460 48.635 161.475 ;
        RECT 57.505 161.460 57.835 161.475 ;
        RECT 80.045 161.460 80.375 161.475 ;
        RECT 99.365 161.460 99.695 161.475 ;
        RECT 105.345 161.460 105.675 161.475 ;
        RECT 48.305 161.160 105.675 161.460 ;
        RECT 48.305 161.145 48.635 161.160 ;
        RECT 57.505 161.145 57.835 161.160 ;
        RECT 80.045 161.145 80.375 161.160 ;
        RECT 99.365 161.145 99.695 161.160 ;
        RECT 105.345 161.145 105.675 161.160 ;
        RECT 107.645 161.460 107.975 161.475 ;
        RECT 110.405 161.460 110.735 161.475 ;
        RECT 107.645 161.160 110.735 161.460 ;
        RECT 107.645 161.145 107.975 161.160 ;
        RECT 110.405 161.145 110.735 161.160 ;
        RECT 81.885 160.780 82.215 160.795 ;
        RECT 116.130 160.780 116.510 160.790 ;
        RECT 81.885 160.480 116.510 160.780 ;
        RECT 81.885 160.465 82.215 160.480 ;
        RECT 116.130 160.470 116.510 160.480 ;
        RECT 96.145 160.100 96.475 160.115 ;
        RECT 108.565 160.100 108.895 160.115 ;
        RECT 96.145 159.800 108.895 160.100 ;
        RECT 96.145 159.785 96.475 159.800 ;
        RECT 108.565 159.785 108.895 159.800 ;
        RECT 111.785 160.100 112.115 160.115 ;
        RECT 113.165 160.100 113.495 160.115 ;
        RECT 111.785 159.800 113.495 160.100 ;
        RECT 111.785 159.785 112.115 159.800 ;
        RECT 113.165 159.785 113.495 159.800 ;
        RECT 31.830 159.445 33.810 159.775 ;
        RECT 61.830 159.445 63.810 159.775 ;
        RECT 91.830 159.445 93.810 159.775 ;
        RECT 121.830 159.445 123.810 159.775 ;
        RECT 46.830 156.725 48.810 157.055 ;
        RECT 76.830 156.725 78.810 157.055 ;
        RECT 106.830 156.725 108.810 157.055 ;
        RECT 31.830 154.005 33.810 154.335 ;
        RECT 61.830 154.005 63.810 154.335 ;
        RECT 91.830 154.005 93.810 154.335 ;
        RECT 121.830 154.005 123.810 154.335 ;
        RECT 80.505 153.310 80.835 153.315 ;
        RECT 80.250 153.300 80.835 153.310 ;
        RECT 80.050 153.000 80.835 153.300 ;
        RECT 80.250 152.990 80.835 153.000 ;
        RECT 80.505 152.985 80.835 152.990 ;
        RECT 46.830 151.285 48.810 151.615 ;
        RECT 76.830 151.285 78.810 151.615 ;
        RECT 106.830 151.285 108.810 151.615 ;
        RECT 116.130 149.900 116.510 149.910 ;
        RECT 116.130 149.600 124.750 149.900 ;
        RECT 116.130 149.590 116.510 149.600 ;
        RECT 31.830 148.565 33.810 148.895 ;
        RECT 61.830 148.565 63.810 148.895 ;
        RECT 91.830 148.565 93.810 148.895 ;
        RECT 121.830 148.565 123.810 148.895 ;
        RECT 124.450 148.540 124.750 149.600 ;
        RECT 131.340 148.540 133.340 148.690 ;
        RECT 124.450 148.240 133.340 148.540 ;
        RECT 131.340 148.090 133.340 148.240 ;
        RECT 56.585 146.500 56.915 146.515 ;
        RECT 57.250 146.500 57.630 146.510 ;
        RECT 56.585 146.200 57.630 146.500 ;
        RECT 56.585 146.185 56.915 146.200 ;
        RECT 57.250 146.190 57.630 146.200 ;
        RECT 46.830 145.845 48.810 146.175 ;
        RECT 76.830 145.845 78.810 146.175 ;
        RECT 106.830 145.845 108.810 146.175 ;
        RECT 60.930 145.820 61.310 145.830 ;
        RECT 62.565 145.820 62.895 145.835 ;
        RECT 60.930 145.520 62.895 145.820 ;
        RECT 60.930 145.510 61.310 145.520 ;
        RECT 62.565 145.505 62.895 145.520 ;
        RECT 81.885 145.820 82.215 145.835 ;
        RECT 83.010 145.820 83.390 145.830 ;
        RECT 81.885 145.520 83.390 145.820 ;
        RECT 81.885 145.505 82.215 145.520 ;
        RECT 83.010 145.510 83.390 145.520 ;
        RECT 59.090 145.140 59.470 145.150 ;
        RECT 60.725 145.140 61.055 145.155 ;
        RECT 59.090 144.840 61.055 145.140 ;
        RECT 59.090 144.830 59.470 144.840 ;
        RECT 60.725 144.825 61.055 144.840 ;
        RECT 78.665 145.140 78.995 145.155 ;
        RECT 79.330 145.140 79.710 145.150 ;
        RECT 78.665 144.840 79.710 145.140 ;
        RECT 78.665 144.825 78.995 144.840 ;
        RECT 79.330 144.830 79.710 144.840 ;
        RECT 67.625 144.460 67.955 144.475 ;
        RECT 82.805 144.460 83.135 144.475 ;
        RECT 67.625 144.160 83.135 144.460 ;
        RECT 67.625 144.145 67.955 144.160 ;
        RECT 82.805 144.145 83.135 144.160 ;
        RECT 31.830 143.125 33.810 143.455 ;
        RECT 61.830 143.125 63.810 143.455 ;
        RECT 91.830 143.125 93.810 143.455 ;
        RECT 121.830 143.125 123.810 143.455 ;
        RECT 82.090 142.420 82.470 142.430 ;
        RECT 83.265 142.420 83.595 142.435 ;
        RECT 82.090 142.120 83.595 142.420 ;
        RECT 82.090 142.110 82.470 142.120 ;
        RECT 83.265 142.105 83.595 142.120 ;
        RECT 46.830 140.405 48.810 140.735 ;
        RECT 76.830 140.405 78.810 140.735 ;
        RECT 106.830 140.405 108.810 140.735 ;
        RECT 87.865 139.700 88.195 139.715 ;
        RECT 93.845 139.700 94.175 139.715 ;
        RECT 87.865 139.400 94.175 139.700 ;
        RECT 87.865 139.385 88.195 139.400 ;
        RECT 93.845 139.385 94.175 139.400 ;
        RECT 129.090 138.200 134.150 139.430 ;
        RECT 31.830 137.685 33.810 138.015 ;
        RECT 61.830 137.685 63.810 138.015 ;
        RECT 91.830 137.685 93.810 138.015 ;
        RECT 121.830 137.685 123.810 138.015 ;
        RECT 56.330 136.980 56.710 136.990 ;
        RECT 61.645 136.980 61.975 136.995 ;
        RECT 56.330 136.680 61.975 136.980 ;
        RECT 56.330 136.670 56.710 136.680 ;
        RECT 61.645 136.665 61.975 136.680 ;
        RECT 64.405 136.300 64.735 136.315 ;
        RECT 87.865 136.300 88.195 136.315 ;
        RECT 64.405 136.000 88.195 136.300 ;
        RECT 64.405 135.985 64.735 136.000 ;
        RECT 87.865 135.985 88.195 136.000 ;
        RECT 46.830 134.965 48.810 135.295 ;
        RECT 76.830 134.965 78.810 135.295 ;
        RECT 106.830 134.965 108.810 135.295 ;
        RECT 31.830 132.245 33.810 132.575 ;
        RECT 61.830 132.245 63.810 132.575 ;
        RECT 91.830 132.245 93.810 132.575 ;
        RECT 121.830 132.245 123.810 132.575 ;
        RECT 46.830 129.525 48.810 129.855 ;
        RECT 76.830 129.525 78.810 129.855 ;
        RECT 106.830 129.525 108.810 129.855 ;
        RECT 31.830 126.805 33.810 127.135 ;
        RECT 61.830 126.805 63.810 127.135 ;
        RECT 91.830 126.805 93.810 127.135 ;
        RECT 121.830 126.805 123.810 127.135 ;
        RECT 53.365 125.420 53.695 125.435 ;
        RECT 57.250 125.420 57.630 125.430 ;
        RECT 53.365 125.120 57.630 125.420 ;
        RECT 53.365 125.105 53.695 125.120 ;
        RECT 57.250 125.110 57.630 125.120 ;
        RECT 46.830 124.085 48.810 124.415 ;
        RECT 76.830 124.085 78.810 124.415 ;
        RECT 106.830 124.085 108.810 124.415 ;
        RECT 31.830 121.365 33.810 121.695 ;
        RECT 61.830 121.365 63.810 121.695 ;
        RECT 91.830 121.365 93.810 121.695 ;
        RECT 121.830 121.365 123.810 121.695 ;
        RECT 46.830 118.645 48.810 118.975 ;
        RECT 76.830 118.645 78.810 118.975 ;
        RECT 106.830 118.645 108.810 118.975 ;
        RECT 130.185 118.620 130.515 118.635 ;
        RECT 131.340 118.620 133.340 118.770 ;
        RECT 130.185 118.320 133.340 118.620 ;
        RECT 130.185 118.305 130.515 118.320 ;
        RECT 131.340 118.170 133.340 118.320 ;
        RECT 31.830 115.925 33.810 116.255 ;
        RECT 61.830 115.925 63.810 116.255 ;
        RECT 91.830 115.925 93.810 116.255 ;
        RECT 121.830 115.925 123.810 116.255 ;
        RECT 46.830 113.205 48.810 113.535 ;
        RECT 76.830 113.205 78.810 113.535 ;
        RECT 106.830 113.205 108.810 113.535 ;
        RECT 129.700 105.605 133.210 106.625 ;
        RECT 37.630 88.620 38.970 88.755 ;
        RECT 13.950 87.980 14.980 88.515 ;
        RECT 13.950 87.500 14.990 87.980 ;
        RECT 13.950 87.175 14.980 87.500 ;
        RECT 14.070 86.570 14.810 87.175 ;
        RECT 20.050 87.105 20.920 88.515 ;
        RECT 14.070 75.715 14.700 86.570 ;
        RECT 20.170 77.115 20.800 87.105 ;
        RECT 25.910 87.055 26.860 88.515 ;
        RECT 26.070 78.385 26.700 87.055 ;
        RECT 31.730 86.965 32.910 88.585 ;
        RECT 32.005 79.615 32.635 86.965 ;
        RECT 37.630 86.835 39.120 88.620 ;
        RECT 38.060 81.125 38.690 86.835 ;
        RECT 43.790 86.745 45.190 88.605 ;
        RECT 49.710 86.945 51.060 88.615 ;
        RECT 44.175 82.625 44.805 86.745 ;
        RECT 50.070 83.875 50.700 86.945 ;
        RECT 55.530 86.785 56.750 88.545 ;
        RECT 55.825 85.115 56.455 86.785 ;
        RECT 61.670 86.625 63.180 88.615 ;
        RECT 67.680 88.305 68.720 89.815 ;
        RECT 67.885 87.225 68.515 88.305 ;
        RECT 62.110 86.175 62.740 86.625 ;
        RECT 67.885 86.595 130.605 87.225 ;
        RECT 62.110 85.545 118.855 86.175 ;
        RECT 55.825 84.485 107.605 85.115 ;
        RECT 50.070 83.245 96.285 83.875 ;
        RECT 44.175 81.995 85.055 82.625 ;
        RECT 38.060 80.495 73.765 81.125 ;
        RECT 32.005 78.985 62.635 79.615 ;
        RECT 26.070 77.755 51.245 78.385 ;
        RECT 20.170 76.485 40.645 77.115 ;
        RECT 14.070 75.660 29.295 75.715 ;
        RECT 40.015 75.710 40.645 76.485 ;
        RECT 14.070 75.085 30.410 75.660 ;
        RECT 27.850 74.670 30.410 75.085 ;
        RECT 3.910 71.345 6.100 73.215 ;
        RECT 27.850 73.120 30.450 74.670 ;
        RECT 39.060 74.510 41.620 75.710 ;
        RECT 50.615 75.580 51.245 77.755 ;
        RECT 62.005 75.690 62.635 78.985 ;
        RECT 49.930 74.650 52.490 75.580 ;
        RECT 0.970 70.330 3.070 70.430 ;
        RECT 15.510 70.330 17.040 71.185 ;
        RECT 0.960 68.750 17.040 70.330 ;
        RECT 0.970 68.710 3.070 68.750 ;
        RECT 15.510 68.635 17.040 68.750 ;
        RECT 20.145 54.060 20.605 54.135 ;
        RECT 25.715 54.060 26.175 54.085 ;
        RECT 20.145 53.620 26.175 54.060 ;
        RECT 20.145 53.565 20.605 53.620 ;
        RECT 25.715 53.515 26.175 53.620 ;
        RECT 22.405 48.870 22.885 48.935 ;
        RECT 22.405 48.550 24.205 48.870 ;
        RECT 22.405 48.385 22.885 48.550 ;
        RECT 23.635 45.710 24.195 48.550 ;
        RECT 27.515 45.710 27.995 45.735 ;
        RECT 23.635 45.290 27.995 45.710 ;
        RECT 23.635 45.280 24.195 45.290 ;
        RECT 27.515 45.185 27.995 45.290 ;
        RECT 20.745 40.120 21.225 40.225 ;
        RECT 24.545 40.120 25.105 40.130 ;
        RECT 20.745 39.700 25.105 40.120 ;
        RECT 20.745 39.675 21.225 39.700 ;
        RECT 24.545 36.860 25.105 39.700 ;
        RECT 25.855 36.860 26.335 37.025 ;
        RECT 24.535 36.540 26.335 36.860 ;
        RECT 25.855 36.475 26.335 36.540 ;
        RECT 22.565 31.790 23.025 31.895 ;
        RECT 28.135 31.790 28.595 31.845 ;
        RECT 22.565 31.350 28.595 31.790 ;
        RECT 22.565 31.325 23.025 31.350 ;
        RECT 28.135 31.275 28.595 31.350 ;
        RECT 29.765 12.265 30.255 73.120 ;
        RECT 38.960 73.080 41.730 74.510 ;
        RECT 31.345 54.070 31.805 54.145 ;
        RECT 36.915 54.070 37.375 54.095 ;
        RECT 31.345 53.630 37.375 54.070 ;
        RECT 31.345 53.575 31.805 53.630 ;
        RECT 36.915 53.525 37.375 53.630 ;
        RECT 33.605 48.880 34.085 48.945 ;
        RECT 33.605 48.560 35.405 48.880 ;
        RECT 33.605 48.395 34.085 48.560 ;
        RECT 34.835 45.720 35.395 48.560 ;
        RECT 38.715 45.720 39.195 45.745 ;
        RECT 34.835 45.300 39.195 45.720 ;
        RECT 34.835 45.290 35.395 45.300 ;
        RECT 38.715 45.195 39.195 45.300 ;
        RECT 32.025 40.120 32.505 40.225 ;
        RECT 35.825 40.120 36.385 40.130 ;
        RECT 32.025 39.700 36.385 40.120 ;
        RECT 32.025 39.675 32.505 39.700 ;
        RECT 35.825 36.860 36.385 39.700 ;
        RECT 37.135 36.860 37.615 37.025 ;
        RECT 35.815 36.540 37.615 36.860 ;
        RECT 37.135 36.475 37.615 36.540 ;
        RECT 33.845 31.790 34.305 31.895 ;
        RECT 39.415 31.790 39.875 31.845 ;
        RECT 33.845 31.350 39.875 31.790 ;
        RECT 33.845 31.325 34.305 31.350 ;
        RECT 39.415 31.275 39.875 31.350 ;
        RECT 41.055 12.360 41.545 73.080 ;
        RECT 49.930 73.030 52.530 74.650 ;
        RECT 61.330 74.530 63.890 75.690 ;
        RECT 73.135 75.580 73.765 80.495 ;
        RECT 84.425 75.690 85.055 81.995 ;
        RECT 72.340 74.980 74.900 75.580 ;
        RECT 42.565 54.040 43.025 54.115 ;
        RECT 48.135 54.040 48.595 54.065 ;
        RECT 42.565 53.600 48.595 54.040 ;
        RECT 42.565 53.545 43.025 53.600 ;
        RECT 48.135 53.495 48.595 53.600 ;
        RECT 44.825 48.850 45.305 48.915 ;
        RECT 44.825 48.530 46.625 48.850 ;
        RECT 44.825 48.365 45.305 48.530 ;
        RECT 46.055 45.690 46.615 48.530 ;
        RECT 49.935 45.690 50.415 45.715 ;
        RECT 46.055 45.270 50.415 45.690 ;
        RECT 46.055 45.260 46.615 45.270 ;
        RECT 49.935 45.165 50.415 45.270 ;
        RECT 43.315 40.100 43.795 40.205 ;
        RECT 47.115 40.100 47.675 40.110 ;
        RECT 43.315 39.680 47.675 40.100 ;
        RECT 43.315 39.655 43.795 39.680 ;
        RECT 47.115 36.840 47.675 39.680 ;
        RECT 48.425 36.840 48.905 37.005 ;
        RECT 47.105 36.520 48.905 36.840 ;
        RECT 48.425 36.455 48.905 36.520 ;
        RECT 45.135 31.770 45.595 31.875 ;
        RECT 50.705 31.770 51.165 31.825 ;
        RECT 45.135 31.330 51.165 31.770 ;
        RECT 45.135 31.305 45.595 31.330 ;
        RECT 50.705 31.255 51.165 31.330 ;
        RECT 41.055 12.350 41.555 12.360 ;
        RECT 28.345 11.115 30.465 12.265 ;
        RECT 41.065 11.965 41.555 12.350 ;
        RECT 51.635 12.145 52.125 73.030 ;
        RECT 61.260 73.010 64.060 74.530 ;
        RECT 72.340 73.050 75.020 74.980 ;
        RECT 83.730 74.540 86.290 75.690 ;
        RECT 95.655 75.580 96.285 83.245 ;
        RECT 106.975 75.640 107.605 84.485 ;
        RECT 118.225 75.650 118.855 85.545 ;
        RECT 129.975 75.650 130.605 86.595 ;
        RECT 133.330 76.605 136.060 77.855 ;
        RECT 137.190 76.585 139.920 77.835 ;
        RECT 53.815 54.020 54.275 54.095 ;
        RECT 59.385 54.020 59.845 54.045 ;
        RECT 53.815 53.580 59.845 54.020 ;
        RECT 53.815 53.525 54.275 53.580 ;
        RECT 59.385 53.475 59.845 53.580 ;
        RECT 56.075 48.830 56.555 48.895 ;
        RECT 56.075 48.510 57.875 48.830 ;
        RECT 56.075 48.345 56.555 48.510 ;
        RECT 57.305 45.670 57.865 48.510 ;
        RECT 61.185 45.670 61.665 45.695 ;
        RECT 57.305 45.250 61.665 45.670 ;
        RECT 57.305 45.240 57.865 45.250 ;
        RECT 61.185 45.145 61.665 45.250 ;
        RECT 54.535 40.100 55.015 40.205 ;
        RECT 58.335 40.100 58.895 40.110 ;
        RECT 54.535 39.680 58.895 40.100 ;
        RECT 54.535 39.655 55.015 39.680 ;
        RECT 58.335 36.840 58.895 39.680 ;
        RECT 59.645 36.840 60.125 37.005 ;
        RECT 58.325 36.520 60.125 36.840 ;
        RECT 59.645 36.455 60.125 36.520 ;
        RECT 56.355 31.770 56.815 31.875 ;
        RECT 61.925 31.770 62.385 31.825 ;
        RECT 56.355 31.330 62.385 31.770 ;
        RECT 56.355 31.305 56.815 31.330 ;
        RECT 61.925 31.255 62.385 31.330 ;
        RECT 29.765 11.100 30.255 11.115 ;
        RECT 39.065 11.005 41.615 11.965 ;
        RECT 50.285 10.995 52.405 12.145 ;
        RECT 62.915 12.135 63.405 73.010 ;
        RECT 65.035 54.010 65.495 54.085 ;
        RECT 70.605 54.010 71.065 54.035 ;
        RECT 65.035 53.570 71.065 54.010 ;
        RECT 65.035 53.515 65.495 53.570 ;
        RECT 70.605 53.465 71.065 53.570 ;
        RECT 67.295 48.820 67.775 48.885 ;
        RECT 67.295 48.500 69.095 48.820 ;
        RECT 67.295 48.335 67.775 48.500 ;
        RECT 68.525 45.660 69.085 48.500 ;
        RECT 72.405 45.660 72.885 45.685 ;
        RECT 68.525 45.240 72.885 45.660 ;
        RECT 68.525 45.230 69.085 45.240 ;
        RECT 72.405 45.135 72.885 45.240 ;
        RECT 65.735 40.100 66.215 40.205 ;
        RECT 69.535 40.100 70.095 40.110 ;
        RECT 65.735 39.680 70.095 40.100 ;
        RECT 65.735 39.655 66.215 39.680 ;
        RECT 69.535 36.840 70.095 39.680 ;
        RECT 70.845 36.840 71.325 37.005 ;
        RECT 69.525 36.520 71.325 36.840 ;
        RECT 70.845 36.455 71.325 36.520 ;
        RECT 67.555 31.770 68.015 31.875 ;
        RECT 73.125 31.770 73.585 31.825 ;
        RECT 67.555 31.330 73.585 31.770 ;
        RECT 67.555 31.305 68.015 31.330 ;
        RECT 73.125 31.255 73.585 31.330 ;
        RECT 74.055 12.165 74.545 73.050 ;
        RECT 83.690 73.000 86.290 74.540 ;
        RECT 94.960 74.710 97.520 75.580 ;
        RECT 94.960 73.020 97.570 74.710 ;
        RECT 106.340 74.460 108.900 75.640 ;
        RECT 117.470 74.720 120.030 75.650 ;
        RECT 76.275 54.000 76.735 54.075 ;
        RECT 81.845 54.000 82.305 54.025 ;
        RECT 76.275 53.560 82.305 54.000 ;
        RECT 76.275 53.505 76.735 53.560 ;
        RECT 81.845 53.455 82.305 53.560 ;
        RECT 78.535 48.810 79.015 48.875 ;
        RECT 78.535 48.490 80.335 48.810 ;
        RECT 78.535 48.325 79.015 48.490 ;
        RECT 79.765 45.650 80.325 48.490 ;
        RECT 83.645 45.650 84.125 45.675 ;
        RECT 79.765 45.230 84.125 45.650 ;
        RECT 79.765 45.220 80.325 45.230 ;
        RECT 83.645 45.125 84.125 45.230 ;
        RECT 77.025 40.090 77.505 40.195 ;
        RECT 80.825 40.090 81.385 40.100 ;
        RECT 77.025 39.670 81.385 40.090 ;
        RECT 77.025 39.645 77.505 39.670 ;
        RECT 80.825 36.830 81.385 39.670 ;
        RECT 82.135 36.830 82.615 36.995 ;
        RECT 80.815 36.510 82.615 36.830 ;
        RECT 82.135 36.445 82.615 36.510 ;
        RECT 78.845 31.760 79.305 31.865 ;
        RECT 84.415 31.760 84.875 31.815 ;
        RECT 78.845 31.320 84.875 31.760 ;
        RECT 78.845 31.295 79.305 31.320 ;
        RECT 84.415 31.245 84.875 31.320 ;
        RECT 61.365 10.985 63.485 12.135 ;
        RECT 72.675 11.015 74.795 12.165 ;
        RECT 85.375 12.155 85.865 73.000 ;
        RECT 87.525 54.010 87.985 54.085 ;
        RECT 93.095 54.010 93.555 54.035 ;
        RECT 87.525 53.570 93.555 54.010 ;
        RECT 87.525 53.515 87.985 53.570 ;
        RECT 93.095 53.465 93.555 53.570 ;
        RECT 89.785 48.820 90.265 48.885 ;
        RECT 89.785 48.500 91.585 48.820 ;
        RECT 89.785 48.335 90.265 48.500 ;
        RECT 91.015 45.660 91.575 48.500 ;
        RECT 94.895 45.660 95.375 45.685 ;
        RECT 91.015 45.240 95.375 45.660 ;
        RECT 91.015 45.230 91.575 45.240 ;
        RECT 94.895 45.135 95.375 45.240 ;
        RECT 88.265 40.110 88.745 40.215 ;
        RECT 92.065 40.110 92.625 40.120 ;
        RECT 88.265 39.690 92.625 40.110 ;
        RECT 88.265 39.665 88.745 39.690 ;
        RECT 92.065 36.850 92.625 39.690 ;
        RECT 93.375 36.850 93.855 37.015 ;
        RECT 92.055 36.530 93.855 36.850 ;
        RECT 93.375 36.465 93.855 36.530 ;
        RECT 90.085 31.780 90.545 31.885 ;
        RECT 95.655 31.780 96.115 31.835 ;
        RECT 90.085 31.340 96.115 31.780 ;
        RECT 90.085 31.315 90.545 31.340 ;
        RECT 95.655 31.265 96.115 31.340 ;
        RECT 96.605 12.155 97.095 73.020 ;
        RECT 106.150 73.000 109.060 74.460 ;
        RECT 117.470 73.070 120.000 74.720 ;
        RECT 129.290 74.650 131.850 75.650 ;
        RECT 129.300 73.140 131.820 74.650 ;
        RECT 98.805 54.000 99.265 54.075 ;
        RECT 104.375 54.000 104.835 54.025 ;
        RECT 98.805 53.560 104.835 54.000 ;
        RECT 98.805 53.505 99.265 53.560 ;
        RECT 104.375 53.455 104.835 53.560 ;
        RECT 101.065 48.810 101.545 48.875 ;
        RECT 101.065 48.490 102.865 48.810 ;
        RECT 101.065 48.325 101.545 48.490 ;
        RECT 102.295 45.650 102.855 48.490 ;
        RECT 106.175 45.650 106.655 45.675 ;
        RECT 102.295 45.230 106.655 45.650 ;
        RECT 102.295 45.220 102.855 45.230 ;
        RECT 106.175 45.125 106.655 45.230 ;
        RECT 99.475 40.130 99.955 40.235 ;
        RECT 103.275 40.130 103.835 40.140 ;
        RECT 99.475 39.710 103.835 40.130 ;
        RECT 99.475 39.685 99.955 39.710 ;
        RECT 103.275 36.870 103.835 39.710 ;
        RECT 104.585 36.870 105.065 37.035 ;
        RECT 103.265 36.550 105.065 36.870 ;
        RECT 104.585 36.485 105.065 36.550 ;
        RECT 101.295 31.800 101.755 31.905 ;
        RECT 106.865 31.800 107.325 31.855 ;
        RECT 101.295 31.360 107.325 31.800 ;
        RECT 101.295 31.335 101.755 31.360 ;
        RECT 106.865 31.285 107.325 31.360 ;
        RECT 107.865 12.205 108.355 73.000 ;
        RECT 110.075 54.000 110.535 54.075 ;
        RECT 115.645 54.000 116.105 54.025 ;
        RECT 110.075 53.560 116.105 54.000 ;
        RECT 110.075 53.505 110.535 53.560 ;
        RECT 115.645 53.455 116.105 53.560 ;
        RECT 112.335 48.810 112.815 48.875 ;
        RECT 112.335 48.490 114.135 48.810 ;
        RECT 112.335 48.325 112.815 48.490 ;
        RECT 113.565 45.650 114.125 48.490 ;
        RECT 117.445 45.650 117.925 45.675 ;
        RECT 113.565 45.230 117.925 45.650 ;
        RECT 113.565 45.220 114.125 45.230 ;
        RECT 117.445 45.125 117.925 45.230 ;
        RECT 110.675 40.170 111.155 40.275 ;
        RECT 114.475 40.170 115.035 40.180 ;
        RECT 110.675 39.750 115.035 40.170 ;
        RECT 110.675 39.725 111.155 39.750 ;
        RECT 114.475 36.910 115.035 39.750 ;
        RECT 115.785 36.910 116.265 37.075 ;
        RECT 114.465 36.590 116.265 36.910 ;
        RECT 115.785 36.525 116.265 36.590 ;
        RECT 112.495 31.840 112.955 31.945 ;
        RECT 118.065 31.840 118.525 31.895 ;
        RECT 112.495 31.400 118.525 31.840 ;
        RECT 112.495 31.375 112.955 31.400 ;
        RECT 118.065 31.325 118.525 31.400 ;
        RECT 119.085 12.205 119.575 73.070 ;
        RECT 121.325 54.000 121.785 54.075 ;
        RECT 126.895 54.000 127.355 54.025 ;
        RECT 121.325 53.560 127.355 54.000 ;
        RECT 121.325 53.505 121.785 53.560 ;
        RECT 126.895 53.455 127.355 53.560 ;
        RECT 123.585 48.810 124.065 48.875 ;
        RECT 123.585 48.490 125.385 48.810 ;
        RECT 123.585 48.325 124.065 48.490 ;
        RECT 124.815 45.650 125.375 48.490 ;
        RECT 128.695 45.650 129.175 45.675 ;
        RECT 124.815 45.230 129.175 45.650 ;
        RECT 124.815 45.220 125.375 45.230 ;
        RECT 128.695 45.125 129.175 45.230 ;
        RECT 121.885 40.190 122.365 40.295 ;
        RECT 125.685 40.190 126.245 40.200 ;
        RECT 121.885 39.770 126.245 40.190 ;
        RECT 121.885 39.745 122.365 39.770 ;
        RECT 125.685 36.930 126.245 39.770 ;
        RECT 126.995 36.930 127.475 37.095 ;
        RECT 125.675 36.610 127.475 36.930 ;
        RECT 126.995 36.545 127.475 36.610 ;
        RECT 123.705 31.860 124.165 31.965 ;
        RECT 129.275 31.860 129.735 31.915 ;
        RECT 123.705 31.420 129.735 31.860 ;
        RECT 123.705 31.395 124.165 31.420 ;
        RECT 129.275 31.345 129.735 31.420 ;
        RECT 130.335 12.235 130.825 73.140 ;
        RECT 74.055 11.010 74.545 11.015 ;
        RECT 83.795 11.005 85.915 12.155 ;
        RECT 95.095 11.005 97.215 12.155 ;
        RECT 106.285 11.055 108.405 12.205 ;
        RECT 117.515 11.055 119.635 12.205 ;
        RECT 128.815 11.085 130.935 12.235 ;
        RECT 107.865 11.010 108.355 11.055 ;
        RECT 119.085 11.050 119.575 11.055 ;
        RECT 85.375 11.000 85.865 11.005 ;
        RECT 96.605 10.980 97.095 11.005 ;
        RECT 74.290 0.135 75.680 1.435 ;
        RECT 93.500 0.205 94.890 1.505 ;
        RECT 112.900 0.335 114.290 1.635 ;
        RECT 131.800 0.405 133.540 1.905 ;
        RECT 151.600 0.275 152.970 1.445 ;
      LAYER met4 ;
        RECT 30.420 225.130 30.670 225.140 ;
        RECT 30.300 224.760 30.670 225.130 ;
        RECT 30.970 224.760 33.430 225.140 ;
        RECT 33.730 224.760 36.190 225.140 ;
        RECT 36.490 224.760 38.950 225.140 ;
        RECT 39.250 224.760 41.710 225.140 ;
        RECT 42.010 224.760 44.470 225.140 ;
        RECT 44.770 224.760 47.230 225.140 ;
        RECT 47.530 224.760 49.990 225.140 ;
        RECT 50.290 224.760 52.750 225.140 ;
        RECT 53.050 224.760 55.510 225.140 ;
        RECT 55.810 224.760 58.270 225.140 ;
        RECT 58.570 224.760 61.030 225.140 ;
        RECT 61.330 224.760 63.790 225.140 ;
        RECT 64.090 224.760 66.550 225.140 ;
        RECT 66.850 224.760 69.310 225.140 ;
        RECT 69.610 224.760 72.070 225.140 ;
        RECT 72.370 224.760 74.830 225.140 ;
        RECT 75.130 224.760 77.590 225.140 ;
        RECT 77.890 224.760 80.350 225.140 ;
        RECT 80.650 224.760 83.110 225.140 ;
        RECT 83.410 224.760 85.870 225.140 ;
        RECT 86.170 224.760 88.630 225.140 ;
        RECT 88.930 224.760 91.390 225.140 ;
        RECT 91.690 224.760 94.150 225.140 ;
        RECT 94.450 224.760 96.910 225.140 ;
        RECT 97.210 224.760 99.670 225.140 ;
        RECT 99.970 224.760 102.430 225.140 ;
        RECT 102.730 224.760 105.190 225.140 ;
        RECT 105.490 224.760 107.950 225.140 ;
        RECT 108.250 224.760 110.710 225.140 ;
        RECT 111.010 224.760 113.470 225.140 ;
        RECT 113.770 224.760 116.230 225.140 ;
        RECT 116.530 224.760 118.990 225.140 ;
        RECT 119.290 224.760 121.750 225.140 ;
        RECT 122.050 224.760 124.510 225.140 ;
        RECT 124.810 224.760 127.270 225.140 ;
        RECT 127.570 224.760 130.030 225.140 ;
        RECT 130.330 224.760 132.790 225.140 ;
        RECT 133.090 224.760 133.520 225.140 ;
        RECT 30.300 224.240 133.520 224.760 ;
        RECT 135.385 224.760 135.550 225.185 ;
        RECT 135.850 224.760 136.745 225.185 ;
        RECT 30.300 219.100 31.660 224.240 ;
        RECT 135.385 223.875 136.745 224.760 ;
        RECT 138.175 224.760 138.310 225.115 ;
        RECT 138.610 224.760 139.535 225.115 ;
        RECT 138.175 223.805 139.535 224.760 ;
        RECT 143.225 224.760 143.830 225.145 ;
        RECT 144.130 224.760 144.585 225.145 ;
        RECT 143.225 223.835 144.585 224.760 ;
        RECT 6.000 218.040 31.660 219.100 ;
        RECT 30.300 217.960 31.660 218.040 ;
        RECT 31.820 113.130 33.820 211.530 ;
        RECT 46.820 113.130 48.820 211.530 ;
        RECT 56.355 167.945 56.685 168.275 ;
        RECT 56.370 136.995 56.670 167.945 ;
        RECT 60.955 166.585 61.285 166.915 ;
        RECT 59.115 161.825 59.445 162.155 ;
        RECT 57.275 146.185 57.605 146.515 ;
        RECT 56.355 136.665 56.685 136.995 ;
        RECT 57.290 125.435 57.590 146.185 ;
        RECT 59.130 145.155 59.430 161.825 ;
        RECT 60.970 145.835 61.270 166.585 ;
        RECT 60.955 145.505 61.285 145.835 ;
        RECT 59.115 144.825 59.445 145.155 ;
        RECT 57.275 125.105 57.605 125.435 ;
        RECT 61.820 113.130 63.820 211.530 ;
        RECT 76.820 113.130 78.820 211.530 ;
        RECT 79.355 192.425 79.685 192.755 ;
        RECT 79.370 145.155 79.670 192.425 ;
        RECT 84.875 184.945 85.205 185.275 ;
        RECT 82.115 184.265 82.445 184.595 ;
        RECT 80.275 181.545 80.605 181.875 ;
        RECT 80.290 153.315 80.590 181.545 ;
        RECT 80.275 152.985 80.605 153.315 ;
        RECT 79.355 144.825 79.685 145.155 ;
        RECT 82.130 142.435 82.430 184.265 ;
        RECT 83.035 181.545 83.365 181.875 ;
        RECT 83.050 145.835 83.350 181.545 ;
        RECT 84.890 173.035 85.190 184.945 ;
        RECT 84.875 172.705 85.205 173.035 ;
        RECT 83.035 145.505 83.365 145.835 ;
        RECT 82.115 142.105 82.445 142.435 ;
        RECT 91.820 113.130 93.820 211.530 ;
        RECT 106.820 113.130 108.820 211.530 ;
        RECT 116.155 160.465 116.485 160.795 ;
        RECT 116.170 149.915 116.470 160.465 ;
        RECT 116.155 149.585 116.485 149.915 ;
        RECT 121.820 113.130 123.820 211.530 ;
        RECT 118.110 97.700 120.130 99.670 ;
        RECT 121.810 97.750 123.830 99.720 ;
        RECT 118.130 93.980 120.130 97.700 ;
        RECT 121.820 96.830 123.820 97.750 ;
        RECT 121.820 94.830 139.410 96.830 ;
        RECT 118.130 91.980 135.580 93.980 ;
        RECT 133.580 77.835 135.580 91.980 ;
        RECT 133.375 76.625 136.015 77.835 ;
        RECT 137.410 77.815 139.410 94.830 ;
        RECT 137.235 76.605 139.875 77.815 ;
        RECT 3.955 71.365 4.000 73.195 ;
        RECT 6.000 71.365 6.055 73.195 ;
        RECT 3.000 68.705 3.025 70.435 ;
        RECT 15.555 68.655 16.995 71.165 ;
        RECT 74.335 1.000 75.635 1.415 ;
        RECT 74.335 0.155 74.530 1.000 ;
        RECT 75.430 0.155 75.635 1.000 ;
        RECT 93.545 1.000 94.845 1.485 ;
        RECT 93.545 0.225 93.850 1.000 ;
        RECT 94.750 0.225 94.845 1.000 ;
        RECT 112.945 1.000 114.245 1.615 ;
        RECT 112.945 0.355 113.170 1.000 ;
        RECT 114.070 0.355 114.245 1.000 ;
        RECT 131.845 1.000 133.495 1.885 ;
        RECT 131.845 0.425 132.490 1.000 ;
        RECT 133.390 0.425 133.495 1.000 ;
        RECT 151.645 1.000 152.925 1.425 ;
        RECT 151.645 0.295 151.810 1.000 ;
        RECT 152.710 0.295 152.925 1.000 ;
  END
END tt_um_08_sws
END LIBRARY

