VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_08_sws
  CLASS BLOCK ;
  FOREIGN tt_um_08_sws ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    ANTENNAGATEAREA 200.000000 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    ANTENNAGATEAREA 550.000000 ;
    ANTENNADIFFAREA 2.900000 ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    ANTENNAGATEAREA 550.000000 ;
    ANTENNADIFFAREA 2.900000 ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    ANTENNADIFFAREA 29.000000 ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    ANTENNADIFFAREA 29.000000 ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    ANTENNADIFFAREA 394.109192 ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 11.575 214.330 11.745 214.520 ;
        RECT 13.010 214.380 13.130 214.490 ;
        RECT 14.795 214.330 14.965 214.520 ;
        RECT 16.635 214.330 16.805 214.520 ;
        RECT 22.155 214.330 22.325 214.520 ;
        RECT 27.675 214.330 27.845 214.520 ;
        RECT 29.515 214.330 29.685 214.520 ;
        RECT 35.035 214.330 35.205 214.520 ;
        RECT 40.555 214.330 40.725 214.520 ;
        RECT 42.395 214.330 42.565 214.520 ;
        RECT 47.915 214.330 48.085 214.520 ;
        RECT 53.435 214.330 53.605 214.520 ;
        RECT 55.275 214.330 55.445 214.520 ;
        RECT 60.795 214.330 60.965 214.520 ;
        RECT 66.315 214.330 66.485 214.520 ;
        RECT 68.155 214.330 68.325 214.520 ;
        RECT 73.675 214.330 73.845 214.520 ;
        RECT 79.195 214.330 79.365 214.520 ;
        RECT 81.035 214.330 81.205 214.520 ;
        RECT 86.555 214.330 86.725 214.520 ;
        RECT 92.075 214.330 92.245 214.520 ;
        RECT 93.915 214.330 94.085 214.520 ;
        RECT 99.435 214.330 99.605 214.520 ;
        RECT 104.955 214.330 105.125 214.520 ;
        RECT 105.930 214.380 106.050 214.490 ;
        RECT 111.395 214.330 111.565 214.520 ;
        RECT 116.915 214.330 117.085 214.520 ;
        RECT 118.295 214.330 118.465 214.520 ;
        RECT 11.435 213.520 12.805 214.330 ;
        RECT 13.275 213.520 15.105 214.330 ;
        RECT 15.125 213.460 15.555 214.245 ;
        RECT 15.575 213.520 16.945 214.330 ;
        RECT 16.955 213.520 22.465 214.330 ;
        RECT 22.475 213.520 27.985 214.330 ;
        RECT 28.005 213.460 28.435 214.245 ;
        RECT 28.455 213.520 29.825 214.330 ;
        RECT 29.835 213.520 35.345 214.330 ;
        RECT 35.355 213.520 40.865 214.330 ;
        RECT 40.885 213.460 41.315 214.245 ;
        RECT 41.335 213.520 42.705 214.330 ;
        RECT 42.715 213.520 48.225 214.330 ;
        RECT 48.235 213.520 53.745 214.330 ;
        RECT 53.765 213.460 54.195 214.245 ;
        RECT 54.215 213.520 55.585 214.330 ;
        RECT 55.595 213.520 61.105 214.330 ;
        RECT 61.115 213.520 66.625 214.330 ;
        RECT 66.645 213.460 67.075 214.245 ;
        RECT 67.095 213.520 68.465 214.330 ;
        RECT 68.475 213.520 73.985 214.330 ;
        RECT 73.995 213.520 79.505 214.330 ;
        RECT 79.525 213.460 79.955 214.245 ;
        RECT 79.975 213.520 81.345 214.330 ;
        RECT 81.355 213.520 86.865 214.330 ;
        RECT 86.875 213.520 92.385 214.330 ;
        RECT 92.405 213.460 92.835 214.245 ;
        RECT 92.855 213.520 94.225 214.330 ;
        RECT 94.235 213.520 99.745 214.330 ;
        RECT 99.755 213.520 105.265 214.330 ;
        RECT 105.285 213.460 105.715 214.245 ;
        RECT 106.195 213.520 111.705 214.330 ;
        RECT 111.715 213.520 117.225 214.330 ;
        RECT 117.235 213.520 118.605 214.330 ;
      LAYER nwell ;
        RECT 11.240 210.300 118.800 213.130 ;
      LAYER pwell ;
        RECT 11.435 209.100 12.805 209.910 ;
        RECT 13.275 209.100 15.105 209.910 ;
        RECT 15.125 209.185 15.555 209.970 ;
        RECT 16.035 209.100 18.785 209.910 ;
        RECT 18.795 209.100 24.305 209.910 ;
        RECT 24.315 209.100 29.825 209.910 ;
        RECT 29.835 209.100 35.345 209.910 ;
        RECT 35.355 209.100 40.865 209.910 ;
        RECT 40.885 209.185 41.315 209.970 ;
        RECT 41.795 209.100 43.625 209.910 ;
        RECT 43.635 209.100 49.145 209.910 ;
        RECT 49.155 209.100 54.665 209.910 ;
        RECT 54.675 209.780 55.595 210.010 ;
        RECT 58.425 209.780 59.355 210.000 ;
        RECT 54.675 209.100 63.865 209.780 ;
        RECT 63.875 209.100 66.625 209.910 ;
        RECT 66.645 209.185 67.075 209.970 ;
        RECT 68.025 209.100 69.375 210.010 ;
        RECT 70.315 209.100 75.825 209.910 ;
        RECT 75.835 209.100 81.345 209.910 ;
        RECT 81.355 209.100 86.865 209.910 ;
        RECT 86.875 209.100 92.385 209.910 ;
        RECT 92.405 209.185 92.835 209.970 ;
        RECT 93.315 209.100 95.145 209.910 ;
        RECT 95.155 209.100 100.665 209.910 ;
        RECT 100.675 209.100 106.185 209.910 ;
        RECT 106.195 209.100 111.705 209.910 ;
        RECT 111.715 209.100 117.225 209.910 ;
        RECT 117.235 209.100 118.605 209.910 ;
        RECT 11.575 208.890 11.745 209.100 ;
        RECT 13.010 208.940 13.130 209.050 ;
        RECT 14.795 208.910 14.965 209.100 ;
        RECT 15.770 208.940 15.890 209.050 ;
        RECT 16.635 208.890 16.805 209.080 ;
        RECT 18.475 208.910 18.645 209.100 ;
        RECT 22.155 208.890 22.325 209.080 ;
        RECT 23.995 208.910 24.165 209.100 ;
        RECT 27.675 208.890 27.845 209.080 ;
        RECT 28.650 208.940 28.770 209.050 ;
        RECT 29.515 208.910 29.685 209.100 ;
        RECT 34.115 208.890 34.285 209.080 ;
        RECT 35.035 208.910 35.205 209.100 ;
        RECT 39.635 208.890 39.805 209.080 ;
        RECT 40.555 208.910 40.725 209.100 ;
        RECT 41.530 208.940 41.650 209.050 ;
        RECT 43.315 208.910 43.485 209.100 ;
        RECT 45.155 208.890 45.325 209.080 ;
        RECT 48.835 208.910 49.005 209.100 ;
        RECT 50.675 208.890 50.845 209.080 ;
        RECT 52.055 208.890 52.225 209.080 ;
        RECT 52.515 208.890 52.685 209.080 ;
        RECT 54.355 208.910 54.525 209.100 ;
        RECT 63.095 208.890 63.265 209.080 ;
        RECT 63.555 208.910 63.725 209.100 ;
        RECT 64.475 208.890 64.645 209.080 ;
        RECT 66.315 208.910 66.485 209.100 ;
        RECT 67.695 208.945 67.855 209.055 ;
        RECT 69.075 208.910 69.245 209.100 ;
        RECT 69.995 208.945 70.155 209.055 ;
        RECT 73.675 208.890 73.845 209.080 ;
        RECT 75.515 208.910 75.685 209.100 ;
        RECT 79.195 208.890 79.365 209.080 ;
        RECT 81.035 208.890 81.205 209.100 ;
        RECT 86.555 208.890 86.725 209.100 ;
        RECT 92.075 208.890 92.245 209.100 ;
        RECT 93.050 208.940 93.170 209.050 ;
        RECT 94.835 208.910 95.005 209.100 ;
        RECT 100.355 208.910 100.525 209.100 ;
        RECT 101.275 208.890 101.445 209.080 ;
        RECT 104.955 208.890 105.125 209.080 ;
        RECT 105.875 209.050 106.045 209.100 ;
        RECT 105.875 208.940 106.050 209.050 ;
        RECT 105.875 208.910 106.045 208.940 ;
        RECT 111.395 208.890 111.565 209.100 ;
        RECT 116.915 208.890 117.085 209.100 ;
        RECT 118.295 208.890 118.465 209.100 ;
        RECT 11.435 208.080 12.805 208.890 ;
        RECT 13.275 208.080 16.945 208.890 ;
        RECT 16.955 208.080 22.465 208.890 ;
        RECT 22.475 208.080 27.985 208.890 ;
        RECT 28.005 208.020 28.435 208.805 ;
        RECT 28.915 208.080 34.425 208.890 ;
        RECT 34.435 208.080 39.945 208.890 ;
        RECT 39.955 208.080 45.465 208.890 ;
        RECT 45.475 208.080 50.985 208.890 ;
        RECT 51.005 207.980 52.355 208.890 ;
        RECT 52.385 207.980 53.735 208.890 ;
        RECT 53.765 208.020 54.195 208.805 ;
        RECT 54.215 208.210 63.405 208.890 ;
        RECT 54.215 207.980 55.135 208.210 ;
        RECT 57.965 207.990 58.895 208.210 ;
        RECT 63.415 208.080 64.785 208.890 ;
        RECT 64.795 208.210 73.985 208.890 ;
        RECT 64.795 207.980 65.715 208.210 ;
        RECT 68.545 207.990 69.475 208.210 ;
        RECT 73.995 208.080 79.505 208.890 ;
        RECT 79.525 208.020 79.955 208.805 ;
        RECT 79.975 208.080 81.345 208.890 ;
        RECT 81.355 208.080 86.865 208.890 ;
        RECT 86.875 208.080 92.385 208.890 ;
        RECT 92.395 208.210 101.585 208.890 ;
        RECT 92.395 207.980 93.315 208.210 ;
        RECT 96.145 207.990 97.075 208.210 ;
        RECT 101.595 208.080 105.265 208.890 ;
        RECT 105.285 208.020 105.715 208.805 ;
        RECT 106.195 208.080 111.705 208.890 ;
        RECT 111.715 208.080 117.225 208.890 ;
        RECT 117.235 208.080 118.605 208.890 ;
      LAYER nwell ;
        RECT 11.240 204.860 118.800 207.690 ;
      LAYER pwell ;
        RECT 11.435 203.660 12.805 204.470 ;
        RECT 13.275 203.660 15.105 204.470 ;
        RECT 15.125 203.745 15.555 204.530 ;
        RECT 16.035 203.660 18.785 204.470 ;
        RECT 18.795 203.660 24.305 204.470 ;
        RECT 24.315 203.660 29.825 204.470 ;
        RECT 29.835 203.660 35.345 204.470 ;
        RECT 35.355 203.660 40.865 204.470 ;
        RECT 40.885 203.745 41.315 204.530 ;
        RECT 41.795 203.660 47.305 204.470 ;
        RECT 47.315 203.660 52.825 204.470 ;
        RECT 52.835 204.340 54.180 204.570 ;
        RECT 54.675 204.340 56.020 204.570 ;
        RECT 56.515 204.340 57.445 204.570 ;
        RECT 61.115 204.340 62.035 204.570 ;
        RECT 52.835 203.660 54.665 204.340 ;
        RECT 54.675 203.660 56.505 204.340 ;
        RECT 56.515 203.660 60.185 204.340 ;
        RECT 61.115 203.660 63.405 204.340 ;
        RECT 63.415 203.660 66.525 204.570 ;
        RECT 66.645 203.745 67.075 204.530 ;
        RECT 67.095 203.660 68.445 204.570 ;
        RECT 69.405 203.660 70.755 204.570 ;
        RECT 71.235 203.660 73.065 204.470 ;
        RECT 73.075 203.660 78.585 204.470 ;
        RECT 78.595 203.660 84.105 204.470 ;
        RECT 84.115 203.660 85.485 204.440 ;
        RECT 85.495 203.660 91.005 204.470 ;
        RECT 91.025 203.660 92.375 204.570 ;
        RECT 92.405 203.745 92.835 204.530 ;
        RECT 92.855 204.340 93.775 204.570 ;
        RECT 96.605 204.340 97.535 204.560 ;
        RECT 92.855 203.660 102.045 204.340 ;
        RECT 102.515 203.660 106.185 204.470 ;
        RECT 106.195 203.660 111.705 204.470 ;
        RECT 111.715 203.660 117.225 204.470 ;
        RECT 117.235 203.660 118.605 204.470 ;
        RECT 11.575 203.450 11.745 203.660 ;
        RECT 13.010 203.500 13.130 203.610 ;
        RECT 14.795 203.470 14.965 203.660 ;
        RECT 15.770 203.500 15.890 203.610 ;
        RECT 16.635 203.450 16.805 203.640 ;
        RECT 18.475 203.470 18.645 203.660 ;
        RECT 22.155 203.450 22.325 203.640 ;
        RECT 23.995 203.470 24.165 203.660 ;
        RECT 27.675 203.450 27.845 203.640 ;
        RECT 28.650 203.500 28.770 203.610 ;
        RECT 29.515 203.470 29.685 203.660 ;
        RECT 31.355 203.450 31.525 203.640 ;
        RECT 35.035 203.470 35.205 203.660 ;
        RECT 36.875 203.450 37.045 203.640 ;
        RECT 40.555 203.470 40.725 203.660 ;
        RECT 41.530 203.500 41.650 203.610 ;
        RECT 42.395 203.450 42.565 203.640 ;
        RECT 46.995 203.470 47.165 203.660 ;
        RECT 47.915 203.450 48.085 203.640 ;
        RECT 52.515 203.470 52.685 203.660 ;
        RECT 53.435 203.450 53.605 203.640 ;
        RECT 54.355 203.470 54.525 203.660 ;
        RECT 55.275 203.450 55.445 203.640 ;
        RECT 55.735 203.450 55.905 203.640 ;
        RECT 56.195 203.470 56.365 203.660 ;
        RECT 57.575 203.450 57.745 203.640 ;
        RECT 59.875 203.470 60.045 203.660 ;
        RECT 60.795 203.505 60.955 203.615 ;
        RECT 62.230 203.500 62.350 203.610 ;
        RECT 63.095 203.470 63.265 203.660 ;
        RECT 63.555 203.450 63.725 203.640 ;
        RECT 64.935 203.450 65.105 203.640 ;
        RECT 66.315 203.470 66.485 203.660 ;
        RECT 67.235 203.470 67.405 203.640 ;
        RECT 68.160 203.470 68.330 203.660 ;
        RECT 67.235 203.450 67.400 203.470 ;
        RECT 68.615 203.450 68.785 203.640 ;
        RECT 69.075 203.505 69.235 203.615 ;
        RECT 69.535 203.470 69.705 203.660 ;
        RECT 70.970 203.500 71.090 203.610 ;
        RECT 72.295 203.450 72.465 203.640 ;
        RECT 72.755 203.470 72.925 203.660 ;
        RECT 77.815 203.450 77.985 203.640 ;
        RECT 78.275 203.450 78.445 203.660 ;
        RECT 83.795 203.470 83.965 203.660 ;
        RECT 84.255 203.470 84.425 203.660 ;
        RECT 88.855 203.450 89.025 203.640 ;
        RECT 89.370 203.500 89.490 203.610 ;
        RECT 90.695 203.470 90.865 203.660 ;
        RECT 91.155 203.470 91.325 203.660 ;
        RECT 92.075 203.450 92.245 203.640 ;
        RECT 92.535 203.450 92.705 203.640 ;
        RECT 97.320 203.450 97.490 203.640 ;
        RECT 98.055 203.450 98.225 203.640 ;
        RECT 99.435 203.450 99.605 203.640 ;
        RECT 101.275 203.495 101.435 203.605 ;
        RECT 101.735 203.470 101.905 203.660 ;
        RECT 102.250 203.500 102.370 203.610 ;
        RECT 104.955 203.450 105.125 203.640 ;
        RECT 105.875 203.610 106.045 203.660 ;
        RECT 105.875 203.500 106.050 203.610 ;
        RECT 105.875 203.470 106.045 203.500 ;
        RECT 111.395 203.450 111.565 203.660 ;
        RECT 116.915 203.450 117.085 203.660 ;
        RECT 118.295 203.450 118.465 203.660 ;
        RECT 11.435 202.640 12.805 203.450 ;
        RECT 13.275 202.640 16.945 203.450 ;
        RECT 16.955 202.640 22.465 203.450 ;
        RECT 22.475 202.640 27.985 203.450 ;
        RECT 28.005 202.580 28.435 203.365 ;
        RECT 28.915 202.640 31.665 203.450 ;
        RECT 31.675 202.640 37.185 203.450 ;
        RECT 37.195 202.640 42.705 203.450 ;
        RECT 42.715 202.640 48.225 203.450 ;
        RECT 48.235 202.640 53.745 203.450 ;
        RECT 53.765 202.580 54.195 203.365 ;
        RECT 54.215 202.640 55.585 203.450 ;
        RECT 55.595 202.770 57.425 203.450 ;
        RECT 57.435 203.220 59.005 203.450 ;
        RECT 61.095 203.410 62.015 203.450 ;
        RECT 61.095 203.220 62.025 203.410 ;
        RECT 57.435 202.860 62.025 203.220 ;
        RECT 57.435 202.770 62.015 202.860 ;
        RECT 59.015 202.540 62.015 202.770 ;
        RECT 62.495 202.670 63.865 203.450 ;
        RECT 63.875 202.640 65.245 203.450 ;
        RECT 65.565 202.770 67.400 203.450 ;
        RECT 65.565 202.540 66.495 202.770 ;
        RECT 67.555 202.640 68.925 203.450 ;
        RECT 68.935 202.640 72.605 203.450 ;
        RECT 72.615 202.640 78.125 203.450 ;
        RECT 78.145 202.540 79.495 203.450 ;
        RECT 79.525 202.580 79.955 203.365 ;
        RECT 79.975 202.770 89.165 203.450 ;
        RECT 79.975 202.540 80.895 202.770 ;
        RECT 83.725 202.550 84.655 202.770 ;
        RECT 89.635 202.640 92.385 203.450 ;
        RECT 92.405 202.540 93.755 203.450 ;
        RECT 94.005 202.770 97.905 203.450 ;
        RECT 96.975 202.540 97.905 202.770 ;
        RECT 97.915 202.670 99.285 203.450 ;
        RECT 99.295 202.670 100.665 203.450 ;
        RECT 101.595 202.640 105.265 203.450 ;
        RECT 105.285 202.580 105.715 203.365 ;
        RECT 106.195 202.640 111.705 203.450 ;
        RECT 111.715 202.640 117.225 203.450 ;
        RECT 117.235 202.640 118.605 203.450 ;
      LAYER nwell ;
        RECT 11.240 199.420 118.800 202.250 ;
      LAYER pwell ;
        RECT 11.435 198.220 12.805 199.030 ;
        RECT 13.275 198.220 15.105 199.030 ;
        RECT 15.125 198.305 15.555 199.090 ;
        RECT 16.035 198.220 18.785 199.030 ;
        RECT 18.795 198.220 24.305 199.030 ;
        RECT 24.315 198.220 29.825 199.030 ;
        RECT 29.835 198.220 35.345 199.030 ;
        RECT 35.355 198.220 40.865 199.030 ;
        RECT 40.885 198.305 41.315 199.090 ;
        RECT 42.265 198.220 43.615 199.130 ;
        RECT 43.635 198.220 45.005 199.030 ;
        RECT 45.015 198.220 46.385 199.000 ;
        RECT 46.405 198.220 47.755 199.130 ;
        RECT 48.695 198.220 52.365 199.030 ;
        RECT 56.885 198.900 57.815 199.120 ;
        RECT 60.535 198.900 62.745 199.130 ;
        RECT 52.375 198.220 62.745 198.900 ;
        RECT 62.955 198.220 66.625 199.030 ;
        RECT 66.645 198.305 67.075 199.090 ;
        RECT 67.095 198.220 69.845 199.030 ;
        RECT 69.855 198.220 75.365 199.030 ;
        RECT 75.745 199.020 76.665 199.130 ;
        RECT 75.745 198.900 78.080 199.020 ;
        RECT 82.745 198.900 83.665 199.120 ;
        RECT 75.745 198.220 85.025 198.900 ;
        RECT 85.035 198.220 86.865 199.030 ;
        RECT 86.875 198.220 92.385 199.030 ;
        RECT 92.405 198.305 92.835 199.090 ;
        RECT 92.855 198.220 94.685 199.030 ;
        RECT 97.895 198.900 98.825 199.130 ;
        RECT 94.925 198.220 98.825 198.900 ;
        RECT 98.835 198.220 100.665 199.030 ;
        RECT 100.675 198.220 102.045 199.000 ;
        RECT 102.515 198.220 106.185 199.030 ;
        RECT 106.195 198.220 111.705 199.030 ;
        RECT 111.715 198.220 117.225 199.030 ;
        RECT 117.235 198.220 118.605 199.030 ;
        RECT 11.575 198.010 11.745 198.220 ;
        RECT 13.010 198.060 13.130 198.170 ;
        RECT 14.795 198.030 14.965 198.220 ;
        RECT 15.770 198.060 15.890 198.170 ;
        RECT 16.635 198.010 16.805 198.200 ;
        RECT 18.475 198.030 18.645 198.220 ;
        RECT 22.155 198.010 22.325 198.200 ;
        RECT 23.995 198.030 24.165 198.220 ;
        RECT 27.675 198.010 27.845 198.200 ;
        RECT 29.055 198.055 29.215 198.165 ;
        RECT 29.515 198.030 29.685 198.220 ;
        RECT 32.735 198.010 32.905 198.200 ;
        RECT 33.195 198.010 33.365 198.200 ;
        RECT 35.035 198.030 35.205 198.220 ;
        RECT 40.555 198.030 40.725 198.220 ;
        RECT 41.935 198.065 42.095 198.175 ;
        RECT 43.315 198.030 43.485 198.220 ;
        RECT 44.695 198.030 44.865 198.220 ;
        RECT 46.075 198.030 46.245 198.220 ;
        RECT 47.455 198.030 47.625 198.220 ;
        RECT 48.375 198.065 48.535 198.175 ;
        RECT 52.055 198.010 52.225 198.220 ;
        RECT 52.515 198.030 52.685 198.220 ;
        RECT 53.435 198.010 53.605 198.200 ;
        RECT 56.655 198.010 56.825 198.200 ;
        RECT 57.115 198.010 57.285 198.200 ;
        RECT 59.415 198.010 59.585 198.200 ;
        RECT 62.630 198.010 62.800 198.200 ;
        RECT 11.435 197.200 12.805 198.010 ;
        RECT 13.275 197.200 16.945 198.010 ;
        RECT 16.955 197.200 22.465 198.010 ;
        RECT 22.475 197.200 27.985 198.010 ;
        RECT 28.005 197.140 28.435 197.925 ;
        RECT 29.375 197.200 33.045 198.010 ;
        RECT 33.055 197.330 42.335 198.010 ;
        RECT 34.415 197.110 35.335 197.330 ;
        RECT 40.000 197.210 42.335 197.330 ;
        RECT 41.415 197.100 42.335 197.210 ;
        RECT 43.085 197.330 52.365 198.010 ;
        RECT 43.085 197.210 45.420 197.330 ;
        RECT 43.085 197.100 44.005 197.210 ;
        RECT 50.085 197.110 51.005 197.330 ;
        RECT 52.375 197.200 53.745 198.010 ;
        RECT 53.765 197.140 54.195 197.925 ;
        RECT 54.215 197.200 56.965 198.010 ;
        RECT 56.985 197.100 58.335 198.010 ;
        RECT 58.355 197.230 59.725 198.010 ;
        RECT 60.025 197.100 62.945 198.010 ;
        RECT 62.955 197.980 63.900 198.010 ;
        RECT 65.855 197.980 66.025 198.200 ;
        RECT 66.315 198.030 66.485 198.220 ;
        RECT 68.155 198.010 68.325 198.200 ;
        RECT 69.535 198.030 69.705 198.220 ;
        RECT 73.675 198.010 73.845 198.200 ;
        RECT 74.135 198.010 74.305 198.200 ;
        RECT 75.055 198.030 75.225 198.220 ;
        RECT 78.920 198.010 79.090 198.200 ;
        RECT 83.520 198.010 83.690 198.200 ;
        RECT 84.715 198.030 84.885 198.220 ;
        RECT 85.175 198.010 85.345 198.200 ;
        RECT 86.555 198.030 86.725 198.220 ;
        RECT 87.935 198.010 88.105 198.200 ;
        RECT 92.075 198.030 92.245 198.220 ;
        RECT 93.455 198.010 93.625 198.200 ;
        RECT 93.915 198.010 94.085 198.200 ;
        RECT 94.375 198.030 94.545 198.220 ;
        RECT 98.240 198.030 98.410 198.220 ;
        RECT 100.355 198.030 100.525 198.220 ;
        RECT 100.815 198.030 100.985 198.220 ;
        RECT 102.250 198.060 102.370 198.170 ;
        RECT 104.035 198.010 104.205 198.200 ;
        RECT 105.875 198.170 106.045 198.220 ;
        RECT 104.955 198.055 105.115 198.165 ;
        RECT 105.875 198.060 106.050 198.170 ;
        RECT 105.875 198.030 106.045 198.060 ;
        RECT 111.395 198.010 111.565 198.220 ;
        RECT 116.915 198.010 117.085 198.220 ;
        RECT 118.295 198.010 118.465 198.220 ;
        RECT 62.955 197.780 66.025 197.980 ;
        RECT 62.955 197.300 66.165 197.780 ;
        RECT 62.955 197.100 63.900 197.300 ;
        RECT 65.235 197.100 66.165 197.300 ;
        RECT 66.175 197.330 68.465 198.010 ;
        RECT 66.175 197.100 67.095 197.330 ;
        RECT 68.475 197.200 73.985 198.010 ;
        RECT 74.005 197.100 75.355 198.010 ;
        RECT 75.605 197.330 79.505 198.010 ;
        RECT 78.575 197.100 79.505 197.330 ;
        RECT 79.525 197.140 79.955 197.925 ;
        RECT 80.205 197.330 84.105 198.010 ;
        RECT 83.175 197.100 84.105 197.330 ;
        RECT 84.115 197.230 85.485 198.010 ;
        RECT 85.495 197.200 88.245 198.010 ;
        RECT 88.255 197.200 93.765 198.010 ;
        RECT 93.785 197.100 95.135 198.010 ;
        RECT 95.155 197.330 104.345 198.010 ;
        RECT 95.155 197.100 96.075 197.330 ;
        RECT 98.905 197.110 99.835 197.330 ;
        RECT 105.285 197.140 105.715 197.925 ;
        RECT 106.195 197.200 111.705 198.010 ;
        RECT 111.715 197.200 117.225 198.010 ;
        RECT 117.235 197.200 118.605 198.010 ;
      LAYER nwell ;
        RECT 11.240 193.980 118.800 196.810 ;
      LAYER pwell ;
        RECT 11.435 192.780 12.805 193.590 ;
        RECT 13.275 192.780 15.105 193.590 ;
        RECT 15.125 192.865 15.555 193.650 ;
        RECT 15.575 192.780 16.945 193.590 ;
        RECT 16.955 192.780 22.465 193.590 ;
        RECT 22.475 192.780 27.985 193.590 ;
        RECT 27.995 193.460 28.915 193.690 ;
        RECT 31.745 193.460 32.675 193.680 ;
        RECT 27.995 192.780 37.185 193.460 ;
        RECT 37.195 192.780 38.565 193.590 ;
        RECT 38.575 192.780 39.945 193.560 ;
        RECT 40.885 192.865 41.315 193.650 ;
        RECT 45.455 193.460 46.385 193.690 ;
        RECT 42.485 192.780 46.385 193.460 ;
        RECT 46.855 192.780 48.685 193.590 ;
        RECT 48.695 192.780 50.065 193.560 ;
        RECT 50.535 192.780 54.205 193.590 ;
        RECT 54.215 192.780 59.725 193.590 ;
        RECT 62.390 193.460 63.310 193.690 ;
        RECT 59.845 192.780 63.310 193.460 ;
        RECT 63.415 193.490 64.360 193.690 ;
        RECT 65.695 193.490 66.625 193.690 ;
        RECT 63.415 193.010 66.625 193.490 ;
        RECT 63.415 192.810 66.485 193.010 ;
        RECT 66.645 192.865 67.075 193.650 ;
        RECT 63.415 192.780 64.360 192.810 ;
        RECT 11.575 192.570 11.745 192.780 ;
        RECT 13.010 192.620 13.130 192.730 ;
        RECT 14.335 192.570 14.505 192.760 ;
        RECT 14.795 192.590 14.965 192.780 ;
        RECT 16.635 192.590 16.805 192.780 ;
        RECT 19.855 192.570 20.025 192.760 ;
        RECT 20.315 192.570 20.485 192.760 ;
        RECT 22.155 192.590 22.325 192.780 ;
        RECT 27.400 192.570 27.570 192.760 ;
        RECT 27.675 192.590 27.845 192.780 ;
        RECT 29.055 192.615 29.215 192.725 ;
        RECT 29.515 192.570 29.685 192.760 ;
        RECT 30.895 192.570 31.065 192.760 ;
        RECT 36.875 192.590 37.045 192.780 ;
        RECT 38.255 192.590 38.425 192.780 ;
        RECT 38.715 192.590 38.885 192.780 ;
        RECT 40.555 192.625 40.715 192.735 ;
        RECT 41.015 192.570 41.185 192.760 ;
        RECT 41.530 192.620 41.650 192.730 ;
        RECT 41.935 192.625 42.095 192.735 ;
        RECT 45.155 192.570 45.325 192.760 ;
        RECT 45.800 192.590 45.970 192.780 ;
        RECT 46.590 192.620 46.710 192.730 ;
        RECT 48.375 192.590 48.545 192.780 ;
        RECT 48.835 192.590 49.005 192.780 ;
        RECT 49.020 192.570 49.190 192.760 ;
        RECT 49.810 192.620 49.930 192.730 ;
        RECT 50.270 192.620 50.390 192.730 ;
        RECT 51.135 192.570 51.305 192.760 ;
        RECT 51.650 192.620 51.770 192.730 ;
        RECT 52.055 192.570 52.225 192.760 ;
        RECT 53.490 192.620 53.610 192.730 ;
        RECT 53.895 192.590 54.065 192.780 ;
        RECT 54.410 192.620 54.530 192.730 ;
        RECT 56.195 192.570 56.365 192.760 ;
        RECT 56.655 192.570 56.825 192.760 ;
        RECT 59.415 192.590 59.585 192.780 ;
        RECT 59.875 192.590 60.045 192.780 ;
        RECT 66.315 192.590 66.485 192.810 ;
        RECT 67.095 192.780 69.385 193.690 ;
        RECT 69.395 192.780 71.225 193.590 ;
        RECT 71.605 193.580 72.525 193.690 ;
        RECT 71.605 193.460 73.940 193.580 ;
        RECT 78.605 193.460 79.525 193.680 ;
        RECT 71.605 192.780 80.885 193.460 ;
        RECT 80.905 192.780 82.255 193.690 ;
        RECT 82.735 192.780 88.245 193.590 ;
        RECT 88.255 193.460 89.185 193.690 ;
        RECT 88.255 192.780 92.155 193.460 ;
        RECT 92.405 192.865 92.835 193.650 ;
        RECT 92.855 192.780 94.685 193.590 ;
        RECT 97.895 193.460 98.825 193.690 ;
        RECT 102.035 193.460 102.965 193.690 ;
        RECT 94.925 192.780 98.825 193.460 ;
        RECT 99.065 192.780 102.965 193.460 ;
        RECT 103.435 192.780 106.185 193.590 ;
        RECT 106.195 192.780 111.705 193.590 ;
        RECT 111.715 192.780 117.225 193.590 ;
        RECT 117.235 192.780 118.605 193.590 ;
        RECT 66.775 192.570 66.945 192.760 ;
        RECT 67.240 192.590 67.410 192.780 ;
        RECT 69.995 192.570 70.165 192.760 ;
        RECT 70.510 192.620 70.630 192.730 ;
        RECT 70.915 192.590 71.085 192.780 ;
        RECT 73.215 192.570 73.385 192.760 ;
        RECT 77.080 192.570 77.250 192.760 ;
        RECT 77.815 192.570 77.985 192.760 ;
        RECT 79.250 192.620 79.370 192.730 ;
        RECT 80.575 192.590 80.745 192.780 ;
        RECT 81.955 192.590 82.125 192.780 ;
        RECT 82.415 192.730 82.585 192.760 ;
        RECT 82.415 192.620 82.590 192.730 ;
        RECT 82.415 192.570 82.585 192.620 ;
        RECT 82.875 192.570 83.045 192.760 ;
        RECT 87.935 192.590 88.105 192.780 ;
        RECT 88.670 192.590 88.840 192.780 ;
        RECT 92.995 192.570 93.165 192.760 ;
        RECT 94.375 192.590 94.545 192.780 ;
        RECT 98.240 192.590 98.410 192.780 ;
        RECT 102.195 192.570 102.365 192.760 ;
        RECT 102.380 192.590 102.550 192.780 ;
        RECT 103.170 192.620 103.290 192.730 ;
        RECT 104.955 192.570 105.125 192.760 ;
        RECT 105.875 192.590 106.045 192.780 ;
        RECT 108.175 192.570 108.345 192.760 ;
        RECT 109.555 192.570 109.725 192.760 ;
        RECT 111.395 192.570 111.565 192.780 ;
        RECT 116.915 192.570 117.085 192.780 ;
        RECT 118.295 192.570 118.465 192.780 ;
        RECT 11.435 191.760 12.805 192.570 ;
        RECT 12.815 191.760 14.645 192.570 ;
        RECT 14.655 191.760 20.165 192.570 ;
        RECT 20.285 191.890 23.750 192.570 ;
        RECT 24.085 191.890 27.985 192.570 ;
        RECT 22.830 191.660 23.750 191.890 ;
        RECT 27.055 191.660 27.985 191.890 ;
        RECT 28.005 191.700 28.435 192.485 ;
        RECT 29.385 191.660 30.735 192.570 ;
        RECT 30.765 191.660 32.115 192.570 ;
        RECT 32.135 191.890 41.325 192.570 ;
        RECT 32.135 191.660 33.055 191.890 ;
        RECT 35.885 191.670 36.815 191.890 ;
        RECT 41.795 191.760 45.465 192.570 ;
        RECT 45.705 191.890 49.605 192.570 ;
        RECT 48.675 191.660 49.605 191.890 ;
        RECT 50.085 191.660 51.435 192.570 ;
        RECT 51.915 191.790 53.285 192.570 ;
        RECT 53.765 191.700 54.195 192.485 ;
        RECT 54.675 191.760 56.505 192.570 ;
        RECT 56.525 191.660 57.875 192.570 ;
        RECT 57.895 191.890 67.085 192.570 ;
        RECT 57.895 191.660 58.815 191.890 ;
        RECT 61.645 191.670 62.575 191.890 ;
        RECT 67.095 191.660 70.205 192.570 ;
        RECT 70.775 191.760 73.525 192.570 ;
        RECT 73.765 191.890 77.665 192.570 ;
        RECT 76.735 191.660 77.665 191.890 ;
        RECT 77.675 191.790 79.045 192.570 ;
        RECT 79.525 191.700 79.955 192.485 ;
        RECT 79.975 191.760 82.725 192.570 ;
        RECT 82.745 191.660 84.095 192.570 ;
        RECT 84.115 191.890 93.305 192.570 ;
        RECT 93.315 191.890 102.505 192.570 ;
        RECT 84.115 191.660 85.035 191.890 ;
        RECT 87.865 191.670 88.795 191.890 ;
        RECT 93.315 191.660 94.235 191.890 ;
        RECT 97.065 191.670 97.995 191.890 ;
        RECT 102.515 191.760 105.265 192.570 ;
        RECT 105.285 191.700 105.715 192.485 ;
        RECT 105.735 191.760 108.485 192.570 ;
        RECT 108.505 191.660 109.855 192.570 ;
        RECT 109.875 191.760 111.705 192.570 ;
        RECT 111.715 191.760 117.225 192.570 ;
        RECT 117.235 191.760 118.605 192.570 ;
      LAYER nwell ;
        RECT 11.240 188.540 118.800 191.370 ;
      LAYER pwell ;
        RECT 11.435 187.340 12.805 188.150 ;
        RECT 13.275 187.340 15.105 188.150 ;
        RECT 15.125 187.425 15.555 188.210 ;
        RECT 15.575 187.340 19.245 188.150 ;
        RECT 19.265 187.340 20.615 188.250 ;
        RECT 20.635 188.020 21.555 188.250 ;
        RECT 24.385 188.020 25.315 188.240 ;
        RECT 20.635 187.340 29.825 188.020 ;
        RECT 30.755 187.340 32.125 188.120 ;
        RECT 32.135 188.020 33.065 188.250 ;
        RECT 39.475 188.020 40.405 188.250 ;
        RECT 32.135 187.340 36.035 188.020 ;
        RECT 36.505 187.340 40.405 188.020 ;
        RECT 40.885 187.425 41.315 188.210 ;
        RECT 41.335 187.340 45.005 188.150 ;
        RECT 45.025 187.340 46.375 188.250 ;
        RECT 46.765 188.140 47.685 188.250 ;
        RECT 46.765 188.020 49.100 188.140 ;
        RECT 53.765 188.020 54.685 188.240 ;
        RECT 46.765 187.340 56.045 188.020 ;
        RECT 56.515 187.340 58.345 188.150 ;
        RECT 58.355 187.340 63.865 188.150 ;
        RECT 63.875 187.340 66.485 188.250 ;
        RECT 66.645 187.425 67.075 188.210 ;
        RECT 67.095 187.340 68.465 188.150 ;
        RECT 68.475 187.340 73.985 188.150 ;
        RECT 74.005 187.340 75.355 188.250 ;
        RECT 75.835 187.340 78.585 188.150 ;
        RECT 78.605 187.340 79.955 188.250 ;
        RECT 79.975 187.340 81.345 188.120 ;
        RECT 85.475 188.020 86.405 188.250 ;
        RECT 82.505 187.340 86.405 188.020 ;
        RECT 86.875 187.340 88.245 188.120 ;
        RECT 88.350 188.020 89.270 188.250 ;
        RECT 88.350 187.340 91.815 188.020 ;
        RECT 92.405 187.425 92.835 188.210 ;
        RECT 92.855 187.340 94.225 188.150 ;
        RECT 94.245 187.340 95.595 188.250 ;
        RECT 96.075 187.340 97.905 188.150 ;
        RECT 97.915 187.340 99.285 188.120 ;
        RECT 99.295 187.340 100.665 188.150 ;
        RECT 100.685 187.340 102.035 188.250 ;
        RECT 104.710 188.020 105.630 188.250 ;
        RECT 102.165 187.340 105.630 188.020 ;
        RECT 105.735 188.020 106.655 188.250 ;
        RECT 109.485 188.020 110.415 188.240 ;
        RECT 105.735 187.340 114.925 188.020 ;
        RECT 115.395 187.340 117.225 188.150 ;
        RECT 117.235 187.340 118.605 188.150 ;
        RECT 11.575 187.130 11.745 187.340 ;
        RECT 13.010 187.180 13.130 187.290 ;
        RECT 14.795 187.150 14.965 187.340 ;
        RECT 15.255 187.130 15.425 187.320 ;
        RECT 18.935 187.150 19.105 187.340 ;
        RECT 19.395 187.150 19.565 187.340 ;
        RECT 20.775 187.130 20.945 187.320 ;
        RECT 26.295 187.130 26.465 187.320 ;
        RECT 26.755 187.130 26.925 187.320 ;
        RECT 29.055 187.175 29.215 187.285 ;
        RECT 29.515 187.150 29.685 187.340 ;
        RECT 30.435 187.185 30.595 187.295 ;
        RECT 30.895 187.150 31.065 187.340 ;
        RECT 32.550 187.150 32.720 187.340 ;
        RECT 32.735 187.130 32.905 187.320 ;
        RECT 38.255 187.130 38.425 187.320 ;
        RECT 38.715 187.130 38.885 187.320 ;
        RECT 39.820 187.150 39.990 187.340 ;
        RECT 40.610 187.180 40.730 187.290 ;
        RECT 44.695 187.150 44.865 187.340 ;
        RECT 45.155 187.150 45.325 187.340 ;
        RECT 51.320 187.130 51.490 187.320 ;
        RECT 52.055 187.130 52.225 187.320 ;
        RECT 53.490 187.180 53.610 187.290 ;
        RECT 54.410 187.180 54.530 187.290 ;
        RECT 55.735 187.150 55.905 187.340 ;
        RECT 56.250 187.180 56.370 187.290 ;
        RECT 58.035 187.130 58.205 187.340 ;
        RECT 63.555 187.130 63.725 187.340 ;
        RECT 64.020 187.320 64.190 187.340 ;
        RECT 64.015 187.150 64.190 187.320 ;
        RECT 67.290 187.180 67.410 187.290 ;
        RECT 64.115 187.130 64.185 187.150 ;
        RECT 67.700 187.130 67.870 187.320 ;
        RECT 68.155 187.150 68.325 187.340 ;
        RECT 73.675 187.150 73.845 187.340 ;
        RECT 75.055 187.150 75.225 187.340 ;
        RECT 75.570 187.180 75.690 187.290 ;
        RECT 78.275 187.150 78.445 187.340 ;
        RECT 78.735 187.150 78.905 187.340 ;
        RECT 79.195 187.130 79.365 187.320 ;
        RECT 81.035 187.150 81.205 187.340 ;
        RECT 81.955 187.185 82.115 187.295 ;
        RECT 85.820 187.150 85.990 187.340 ;
        RECT 86.610 187.180 86.730 187.290 ;
        RECT 87.015 187.150 87.185 187.340 ;
        RECT 88.855 187.130 89.025 187.320 ;
        RECT 89.775 187.175 89.935 187.285 ;
        RECT 91.615 187.150 91.785 187.340 ;
        RECT 92.130 187.180 92.250 187.290 ;
        RECT 93.455 187.130 93.625 187.320 ;
        RECT 93.915 187.150 94.085 187.340 ;
        RECT 94.375 187.150 94.545 187.340 ;
        RECT 95.810 187.180 95.930 187.290 ;
        RECT 97.595 187.150 97.765 187.340 ;
        RECT 98.055 187.150 98.225 187.340 ;
        RECT 98.975 187.130 99.145 187.320 ;
        RECT 100.355 187.130 100.525 187.340 ;
        RECT 100.815 187.290 100.985 187.340 ;
        RECT 100.815 187.180 100.990 187.290 ;
        RECT 100.815 187.150 100.985 187.180 ;
        RECT 102.195 187.150 102.365 187.340 ;
        RECT 104.680 187.130 104.850 187.320 ;
        RECT 114.615 187.130 114.785 187.340 ;
        RECT 115.130 187.180 115.250 187.290 ;
        RECT 115.995 187.130 116.165 187.320 ;
        RECT 116.915 187.150 117.085 187.340 ;
        RECT 118.295 187.130 118.465 187.340 ;
        RECT 11.435 186.320 12.805 187.130 ;
        RECT 12.815 186.320 15.565 187.130 ;
        RECT 15.575 186.320 21.085 187.130 ;
        RECT 21.095 186.320 26.605 187.130 ;
        RECT 26.615 186.350 27.985 187.130 ;
        RECT 28.005 186.260 28.435 187.045 ;
        RECT 29.375 186.320 33.045 187.130 ;
        RECT 33.055 186.320 38.565 187.130 ;
        RECT 38.575 186.450 47.680 187.130 ;
        RECT 48.005 186.450 51.905 187.130 ;
        RECT 50.975 186.220 51.905 186.450 ;
        RECT 51.915 186.350 53.285 187.130 ;
        RECT 53.765 186.260 54.195 187.045 ;
        RECT 54.675 186.320 58.345 187.130 ;
        RECT 58.355 186.320 63.865 187.130 ;
        RECT 64.115 186.900 66.385 187.130 ;
        RECT 64.115 186.220 66.870 186.900 ;
        RECT 67.555 186.220 70.165 187.130 ;
        RECT 70.315 186.450 79.505 187.130 ;
        RECT 70.315 186.220 71.235 186.450 ;
        RECT 74.065 186.230 74.995 186.450 ;
        RECT 79.525 186.260 79.955 187.045 ;
        RECT 79.975 186.450 89.165 187.130 ;
        RECT 79.975 186.220 80.895 186.450 ;
        RECT 83.725 186.230 84.655 186.450 ;
        RECT 90.095 186.320 93.765 187.130 ;
        RECT 93.775 186.320 99.285 187.130 ;
        RECT 99.305 186.220 100.655 187.130 ;
        RECT 101.365 186.450 105.265 187.130 ;
        RECT 104.335 186.220 105.265 186.450 ;
        RECT 105.285 186.260 105.715 187.045 ;
        RECT 105.735 186.450 114.925 187.130 ;
        RECT 105.735 186.220 106.655 186.450 ;
        RECT 109.485 186.230 110.415 186.450 ;
        RECT 114.935 186.350 116.305 187.130 ;
        RECT 117.235 186.320 118.605 187.130 ;
      LAYER nwell ;
        RECT 11.240 183.100 118.800 185.930 ;
      LAYER pwell ;
        RECT 11.435 181.900 12.805 182.710 ;
        RECT 13.275 181.900 15.105 182.710 ;
        RECT 15.125 181.985 15.555 182.770 ;
        RECT 16.035 181.900 18.785 182.710 ;
        RECT 18.795 181.900 24.305 182.710 ;
        RECT 24.315 182.580 25.235 182.810 ;
        RECT 28.065 182.580 28.995 182.800 ;
        RECT 24.315 181.900 33.505 182.580 ;
        RECT 33.975 181.900 36.725 182.710 ;
        RECT 39.935 182.580 40.865 182.810 ;
        RECT 36.965 181.900 40.865 182.580 ;
        RECT 40.885 181.985 41.315 182.770 ;
        RECT 41.335 181.900 42.705 182.680 ;
        RECT 42.725 181.900 44.075 182.810 ;
        RECT 46.305 182.700 47.225 182.810 ;
        RECT 46.305 182.580 48.640 182.700 ;
        RECT 53.305 182.580 54.225 182.800 ;
        RECT 44.095 181.900 45.460 182.580 ;
        RECT 46.305 181.900 55.585 182.580 ;
        RECT 56.055 181.900 58.805 182.710 ;
        RECT 59.030 182.130 61.785 182.810 ;
        RECT 63.615 182.580 66.615 182.810 ;
        RECT 59.515 181.900 61.785 182.130 ;
        RECT 62.035 182.490 66.615 182.580 ;
        RECT 62.035 182.130 66.625 182.490 ;
        RECT 62.035 181.900 63.605 182.130 ;
        RECT 65.695 181.940 66.625 182.130 ;
        RECT 66.645 181.985 67.075 182.770 ;
        RECT 67.335 182.130 70.090 182.810 ;
        RECT 65.695 181.900 66.615 181.940 ;
        RECT 67.335 181.900 69.605 182.130 ;
        RECT 70.315 181.900 71.685 182.710 ;
        RECT 74.895 182.580 75.825 182.810 ;
        RECT 71.925 181.900 75.825 182.580 ;
        RECT 75.920 181.900 85.025 182.580 ;
        RECT 85.495 181.900 87.325 182.710 ;
        RECT 87.335 181.900 88.705 182.680 ;
        RECT 89.185 181.900 90.535 182.810 ;
        RECT 91.015 181.900 92.385 182.680 ;
        RECT 92.405 181.985 92.835 182.770 ;
        RECT 93.050 181.900 96.525 182.810 ;
        RECT 96.535 182.580 97.455 182.810 ;
        RECT 100.285 182.580 101.215 182.800 ;
        RECT 108.935 182.580 109.865 182.810 ;
        RECT 96.535 181.900 105.725 182.580 ;
        RECT 105.965 181.900 109.865 182.580 ;
        RECT 110.795 181.900 112.165 182.680 ;
        RECT 112.175 181.900 113.545 182.710 ;
        RECT 113.555 181.900 117.225 182.710 ;
        RECT 117.235 181.900 118.605 182.710 ;
        RECT 11.575 181.690 11.745 181.900 ;
        RECT 13.010 181.740 13.130 181.850 ;
        RECT 14.795 181.710 14.965 181.900 ;
        RECT 15.715 181.850 15.885 181.880 ;
        RECT 15.715 181.740 15.890 181.850 ;
        RECT 15.715 181.690 15.885 181.740 ;
        RECT 16.175 181.690 16.345 181.880 ;
        RECT 18.475 181.710 18.645 181.900 ;
        RECT 23.995 181.710 24.165 181.900 ;
        RECT 26.295 181.690 26.465 181.880 ;
        RECT 27.675 181.690 27.845 181.880 ;
        RECT 32.000 181.690 32.170 181.880 ;
        RECT 33.195 181.710 33.365 181.900 ;
        RECT 33.655 181.850 33.825 181.880 ;
        RECT 33.655 181.740 33.830 181.850 ;
        RECT 34.170 181.740 34.290 181.850 ;
        RECT 33.655 181.690 33.825 181.740 ;
        RECT 36.415 181.710 36.585 181.900 ;
        RECT 36.875 181.690 37.045 181.880 ;
        RECT 37.335 181.690 37.505 181.880 ;
        RECT 40.280 181.710 40.450 181.900 ;
        RECT 42.395 181.710 42.565 181.900 ;
        RECT 43.775 181.710 43.945 181.900 ;
        RECT 45.615 181.710 45.785 181.880 ;
        RECT 47.050 181.740 47.170 181.850 ;
        RECT 50.860 181.690 51.030 181.880 ;
        RECT 51.650 181.740 51.770 181.850 ;
        RECT 53.435 181.690 53.605 181.880 ;
        RECT 55.275 181.710 55.445 181.900 ;
        RECT 55.790 181.740 55.910 181.850 ;
        RECT 56.655 181.690 56.825 181.880 ;
        RECT 58.495 181.690 58.665 181.900 ;
        RECT 61.715 181.880 61.785 181.900 ;
        RECT 61.715 181.710 61.885 181.880 ;
        RECT 62.175 181.690 62.345 181.900 ;
        RECT 67.335 181.880 67.405 181.900 ;
        RECT 62.635 181.690 62.805 181.880 ;
        RECT 66.775 181.710 66.945 181.880 ;
        RECT 67.235 181.710 67.405 181.880 ;
        RECT 66.775 181.690 66.845 181.710 ;
        RECT 68.155 181.690 68.325 181.880 ;
        RECT 68.615 181.690 68.785 181.880 ;
        RECT 71.375 181.710 71.545 181.900 ;
        RECT 73.675 181.690 73.845 181.880 ;
        RECT 75.240 181.710 75.410 181.900 ;
        RECT 79.195 181.690 79.365 181.880 ;
        RECT 80.170 181.740 80.290 181.850 ;
        RECT 81.955 181.690 82.125 181.880 ;
        RECT 84.715 181.690 84.885 181.900 ;
        RECT 85.230 181.740 85.350 181.850 ;
        RECT 85.635 181.735 85.795 181.845 ;
        RECT 87.015 181.710 87.185 181.900 ;
        RECT 88.395 181.710 88.565 181.900 ;
        RECT 88.910 181.740 89.030 181.850 ;
        RECT 90.235 181.710 90.405 181.900 ;
        RECT 90.750 181.740 90.870 181.850 ;
        RECT 91.155 181.710 91.325 181.900 ;
        RECT 94.835 181.690 95.005 181.880 ;
        RECT 96.210 181.710 96.380 181.900 ;
        RECT 104.035 181.690 104.205 181.880 ;
        RECT 104.955 181.735 105.115 181.845 ;
        RECT 105.415 181.710 105.585 181.900 ;
        RECT 109.090 181.690 109.260 181.880 ;
        RECT 109.280 181.710 109.450 181.900 ;
        RECT 110.475 181.690 110.645 181.880 ;
        RECT 110.935 181.690 111.105 181.900 ;
        RECT 112.370 181.740 112.490 181.850 ;
        RECT 112.775 181.690 112.945 181.880 ;
        RECT 113.235 181.710 113.405 181.900 ;
        RECT 114.210 181.740 114.330 181.850 ;
        RECT 116.915 181.690 117.085 181.900 ;
        RECT 118.295 181.690 118.465 181.900 ;
        RECT 11.435 180.880 12.805 181.690 ;
        RECT 13.275 180.880 16.025 181.690 ;
        RECT 16.045 180.780 17.395 181.690 ;
        RECT 17.415 181.010 26.605 181.690 ;
        RECT 17.415 180.780 18.335 181.010 ;
        RECT 21.165 180.790 22.095 181.010 ;
        RECT 26.615 180.910 27.985 181.690 ;
        RECT 28.005 180.820 28.435 181.605 ;
        RECT 28.685 181.010 32.585 181.690 ;
        RECT 31.655 180.780 32.585 181.010 ;
        RECT 32.595 180.910 33.965 181.690 ;
        RECT 34.435 180.880 37.185 181.690 ;
        RECT 37.195 181.010 46.475 181.690 ;
        RECT 47.545 181.010 51.445 181.690 ;
        RECT 38.555 180.790 39.475 181.010 ;
        RECT 44.140 180.890 46.475 181.010 ;
        RECT 45.555 180.780 46.475 180.890 ;
        RECT 50.515 180.780 51.445 181.010 ;
        RECT 51.915 180.880 53.745 181.690 ;
        RECT 53.765 180.820 54.195 181.605 ;
        RECT 54.215 180.880 56.965 181.690 ;
        RECT 56.975 181.010 58.805 181.690 ;
        RECT 56.975 180.780 58.320 181.010 ;
        RECT 58.815 180.880 62.485 181.690 ;
        RECT 62.505 180.780 63.855 181.690 ;
        RECT 64.575 181.460 66.845 181.690 ;
        RECT 64.090 180.780 66.845 181.460 ;
        RECT 67.095 180.880 68.465 181.690 ;
        RECT 68.475 181.010 71.215 181.690 ;
        RECT 71.235 180.880 73.985 181.690 ;
        RECT 73.995 180.880 79.505 181.690 ;
        RECT 79.525 180.820 79.955 181.605 ;
        RECT 80.435 180.880 82.265 181.690 ;
        RECT 82.285 181.010 85.025 181.690 ;
        RECT 85.955 181.010 95.145 181.690 ;
        RECT 95.240 181.010 104.345 181.690 ;
        RECT 85.955 180.780 86.875 181.010 ;
        RECT 89.705 180.790 90.635 181.010 ;
        RECT 105.285 180.820 105.715 181.605 ;
        RECT 105.930 180.780 109.405 181.690 ;
        RECT 109.415 180.910 110.785 181.690 ;
        RECT 110.805 180.780 112.155 181.690 ;
        RECT 112.635 180.910 114.005 181.690 ;
        RECT 114.475 180.880 117.225 181.690 ;
        RECT 117.235 180.880 118.605 181.690 ;
      LAYER nwell ;
        RECT 11.240 177.660 118.800 180.490 ;
      LAYER pwell ;
        RECT 11.435 176.460 12.805 177.270 ;
        RECT 13.275 176.460 15.105 177.270 ;
        RECT 15.125 176.545 15.555 177.330 ;
        RECT 16.495 176.460 20.165 177.270 ;
        RECT 20.185 176.460 21.535 177.370 ;
        RECT 24.210 177.140 25.130 177.370 ;
        RECT 28.435 177.140 29.365 177.370 ;
        RECT 21.665 176.460 25.130 177.140 ;
        RECT 25.465 176.460 29.365 177.140 ;
        RECT 29.375 176.460 30.745 177.270 ;
        RECT 30.755 176.460 34.425 177.270 ;
        RECT 34.435 176.460 37.910 177.370 ;
        RECT 38.115 176.460 40.865 177.270 ;
        RECT 40.885 176.545 41.315 177.330 ;
        RECT 41.335 176.460 45.005 177.270 ;
        RECT 45.015 176.460 48.490 177.370 ;
        RECT 49.155 176.460 50.985 177.270 ;
        RECT 51.005 176.460 53.745 177.140 ;
        RECT 53.755 176.460 55.125 177.270 ;
        RECT 55.135 177.140 56.480 177.370 ;
        RECT 56.975 177.140 58.320 177.370 ;
        RECT 59.300 177.140 60.645 177.370 ;
        RECT 55.135 176.460 56.965 177.140 ;
        RECT 56.975 176.460 58.805 177.140 ;
        RECT 58.815 176.460 60.645 177.140 ;
        RECT 61.575 176.460 64.295 177.370 ;
        RECT 64.795 176.460 66.165 177.240 ;
        RECT 66.645 176.545 67.075 177.330 ;
        RECT 67.095 176.460 68.465 177.240 ;
        RECT 68.475 176.460 71.225 177.270 ;
        RECT 71.235 176.460 73.975 177.140 ;
        RECT 73.995 176.460 75.825 177.270 ;
        RECT 76.205 177.260 77.125 177.370 ;
        RECT 76.205 177.140 78.540 177.260 ;
        RECT 83.205 177.140 84.125 177.360 ;
        RECT 89.615 177.140 90.545 177.370 ;
        RECT 76.205 176.460 85.485 177.140 ;
        RECT 86.645 176.460 90.545 177.140 ;
        RECT 90.555 176.460 92.385 177.270 ;
        RECT 92.405 176.545 92.835 177.330 ;
        RECT 95.510 177.140 96.430 177.370 ;
        RECT 100.655 177.140 101.585 177.370 ;
        RECT 92.965 176.460 96.430 177.140 ;
        RECT 97.685 176.460 101.585 177.140 ;
        RECT 101.595 176.460 105.070 177.370 ;
        RECT 107.575 177.140 108.495 177.370 ;
        RECT 111.325 177.140 112.255 177.360 ;
        RECT 105.275 176.460 106.640 177.140 ;
        RECT 107.575 176.460 116.765 177.140 ;
        RECT 117.235 176.460 118.605 177.270 ;
        RECT 11.575 176.250 11.745 176.460 ;
        RECT 13.010 176.300 13.130 176.410 ;
        RECT 14.335 176.250 14.505 176.440 ;
        RECT 14.795 176.270 14.965 176.460 ;
        RECT 16.175 176.305 16.335 176.415 ;
        RECT 19.855 176.250 20.025 176.460 ;
        RECT 20.315 176.250 20.485 176.460 ;
        RECT 21.695 176.270 21.865 176.460 ;
        RECT 22.615 176.250 22.785 176.440 ;
        RECT 26.295 176.250 26.465 176.440 ;
        RECT 26.755 176.250 26.925 176.440 ;
        RECT 28.650 176.300 28.770 176.410 ;
        RECT 28.780 176.270 28.950 176.460 ;
        RECT 30.435 176.270 30.605 176.460 ;
        RECT 32.270 176.250 32.440 176.440 ;
        RECT 34.115 176.270 34.285 176.460 ;
        RECT 34.580 176.270 34.750 176.460 ;
        RECT 35.950 176.250 36.120 176.440 ;
        RECT 36.420 176.250 36.590 176.440 ;
        RECT 40.150 176.300 40.270 176.410 ;
        RECT 40.555 176.270 40.725 176.460 ;
        RECT 41.935 176.250 42.105 176.440 ;
        RECT 44.695 176.270 44.865 176.460 ;
        RECT 45.160 176.270 45.330 176.460 ;
        RECT 45.610 176.250 45.780 176.440 ;
        RECT 46.080 176.250 46.250 176.440 ;
        RECT 48.890 176.300 49.010 176.410 ;
        RECT 49.810 176.300 49.930 176.410 ;
        RECT 50.675 176.270 50.845 176.460 ;
        RECT 53.435 176.250 53.605 176.460 ;
        RECT 54.410 176.300 54.530 176.410 ;
        RECT 54.815 176.270 54.985 176.460 ;
        RECT 56.655 176.270 56.825 176.460 ;
        RECT 58.035 176.250 58.205 176.440 ;
        RECT 58.495 176.250 58.665 176.460 ;
        RECT 58.955 176.270 59.125 176.460 ;
        RECT 59.875 176.250 60.045 176.440 ;
        RECT 61.255 176.305 61.415 176.415 ;
        RECT 61.715 176.270 61.885 176.460 ;
        RECT 62.175 176.250 62.345 176.440 ;
        RECT 64.015 176.250 64.185 176.440 ;
        RECT 64.530 176.300 64.650 176.410 ;
        RECT 64.935 176.270 65.105 176.460 ;
        RECT 66.370 176.300 66.490 176.410 ;
        RECT 68.155 176.270 68.325 176.460 ;
        RECT 68.615 176.250 68.785 176.440 ;
        RECT 70.455 176.250 70.625 176.440 ;
        RECT 70.915 176.270 71.085 176.460 ;
        RECT 71.375 176.270 71.545 176.460 ;
        RECT 75.055 176.250 75.225 176.440 ;
        RECT 75.515 176.270 75.685 176.460 ;
        RECT 78.920 176.250 79.090 176.440 ;
        RECT 80.170 176.300 80.290 176.410 ;
        RECT 81.495 176.250 81.665 176.440 ;
        RECT 81.955 176.250 82.125 176.440 ;
        RECT 83.335 176.250 83.505 176.440 ;
        RECT 85.175 176.270 85.345 176.460 ;
        RECT 86.095 176.305 86.255 176.415 ;
        RECT 88.855 176.250 89.025 176.440 ;
        RECT 89.960 176.270 90.130 176.460 ;
        RECT 92.075 176.270 92.245 176.460 ;
        RECT 92.995 176.270 93.165 176.460 ;
        RECT 97.135 176.305 97.295 176.415 ;
        RECT 98.515 176.250 98.685 176.440 ;
        RECT 99.895 176.250 100.065 176.440 ;
        RECT 100.360 176.250 100.530 176.440 ;
        RECT 101.000 176.270 101.170 176.460 ;
        RECT 101.740 176.270 101.910 176.460 ;
        RECT 104.955 176.250 105.125 176.440 ;
        RECT 106.335 176.295 106.495 176.405 ;
        RECT 106.795 176.270 106.965 176.440 ;
        RECT 107.310 176.300 107.430 176.410 ;
        RECT 110.200 176.250 110.370 176.440 ;
        RECT 111.395 176.295 111.555 176.405 ;
        RECT 116.455 176.270 116.625 176.460 ;
        RECT 116.915 176.410 117.085 176.440 ;
        RECT 116.915 176.300 117.090 176.410 ;
        RECT 116.915 176.250 117.085 176.300 ;
        RECT 118.295 176.250 118.465 176.460 ;
        RECT 11.435 175.440 12.805 176.250 ;
        RECT 12.815 175.440 14.645 176.250 ;
        RECT 14.655 175.440 20.165 176.250 ;
        RECT 20.175 175.470 21.545 176.250 ;
        RECT 21.555 175.440 22.925 176.250 ;
        RECT 22.935 175.440 26.605 176.250 ;
        RECT 26.625 175.340 27.975 176.250 ;
        RECT 28.005 175.380 28.435 176.165 ;
        RECT 29.110 175.340 32.585 176.250 ;
        RECT 32.790 175.340 36.265 176.250 ;
        RECT 36.275 175.340 39.750 176.250 ;
        RECT 40.415 175.440 42.245 176.250 ;
        RECT 42.450 175.340 45.925 176.250 ;
        RECT 45.935 175.340 49.410 176.250 ;
        RECT 50.075 175.440 53.745 176.250 ;
        RECT 53.765 175.380 54.195 176.165 ;
        RECT 54.675 175.440 58.345 176.250 ;
        RECT 58.355 175.470 59.725 176.250 ;
        RECT 59.735 175.470 61.105 176.250 ;
        RECT 61.115 175.470 62.485 176.250 ;
        RECT 62.495 175.570 64.325 176.250 ;
        RECT 62.495 175.340 63.840 175.570 ;
        RECT 64.375 175.340 68.925 176.250 ;
        RECT 68.935 175.570 70.765 176.250 ;
        RECT 68.935 175.340 70.280 175.570 ;
        RECT 71.695 175.440 75.365 176.250 ;
        RECT 75.605 175.570 79.505 176.250 ;
        RECT 78.575 175.340 79.505 175.570 ;
        RECT 79.525 175.380 79.955 176.165 ;
        RECT 80.445 175.340 81.795 176.250 ;
        RECT 81.815 175.470 83.185 176.250 ;
        RECT 83.195 175.470 84.565 176.250 ;
        RECT 85.495 175.440 89.165 176.250 ;
        RECT 89.545 175.570 98.825 176.250 ;
        RECT 89.545 175.450 91.880 175.570 ;
        RECT 89.545 175.340 90.465 175.450 ;
        RECT 96.545 175.350 97.465 175.570 ;
        RECT 98.835 175.440 100.205 176.250 ;
        RECT 100.215 175.340 103.690 176.250 ;
        RECT 103.895 175.440 105.265 176.250 ;
        RECT 105.285 175.380 105.715 176.165 ;
        RECT 106.885 175.570 110.785 176.250 ;
        RECT 109.855 175.340 110.785 175.570 ;
        RECT 111.715 175.440 117.225 176.250 ;
        RECT 117.235 175.440 118.605 176.250 ;
      LAYER nwell ;
        RECT 11.240 172.220 118.800 175.050 ;
      LAYER pwell ;
        RECT 11.435 171.020 12.805 171.830 ;
        RECT 13.745 171.020 15.095 171.930 ;
        RECT 15.125 171.105 15.555 171.890 ;
        RECT 15.575 171.700 16.495 171.930 ;
        RECT 19.325 171.700 20.255 171.920 ;
        RECT 25.235 171.700 26.155 171.930 ;
        RECT 28.985 171.700 29.915 171.920 ;
        RECT 15.575 171.020 24.765 171.700 ;
        RECT 25.235 171.020 34.425 171.700 ;
        RECT 35.355 171.020 38.830 171.930 ;
        RECT 39.035 171.020 40.865 171.830 ;
        RECT 40.885 171.105 41.315 171.890 ;
        RECT 41.335 171.020 44.085 171.830 ;
        RECT 44.095 171.020 47.570 171.930 ;
        RECT 47.775 171.020 49.605 171.830 ;
        RECT 49.625 171.020 50.975 171.930 ;
        RECT 51.915 171.020 55.585 171.830 ;
        RECT 55.595 171.020 61.105 171.830 ;
        RECT 61.115 171.020 66.625 171.830 ;
        RECT 66.645 171.105 67.075 171.890 ;
        RECT 67.095 171.020 68.465 171.830 ;
        RECT 68.670 171.020 72.145 171.930 ;
        RECT 72.155 171.020 75.630 171.930 ;
        RECT 75.835 171.020 77.665 171.830 ;
        RECT 77.685 171.020 79.035 171.930 ;
        RECT 82.255 171.700 83.185 171.930 ;
        RECT 79.285 171.020 83.185 171.700 ;
        RECT 83.205 171.020 84.555 171.930 ;
        RECT 84.575 171.020 85.945 171.800 ;
        RECT 85.955 171.020 88.705 171.830 ;
        RECT 88.715 171.020 92.190 171.930 ;
        RECT 92.405 171.105 92.835 171.890 ;
        RECT 96.055 171.700 96.985 171.930 ;
        RECT 93.085 171.020 96.985 171.700 ;
        RECT 96.995 171.020 100.470 171.930 ;
        RECT 103.875 171.700 104.805 171.930 ;
        RECT 100.905 171.020 104.805 171.700 ;
        RECT 105.185 171.820 106.105 171.930 ;
        RECT 105.185 171.700 107.520 171.820 ;
        RECT 112.185 171.700 113.105 171.920 ;
        RECT 105.185 171.020 114.465 171.700 ;
        RECT 114.475 171.020 116.305 171.700 ;
        RECT 117.235 171.020 118.605 171.830 ;
        RECT 11.575 170.810 11.745 171.020 ;
        RECT 13.010 170.860 13.130 170.970 ;
        RECT 13.415 170.865 13.575 170.975 ;
        RECT 14.335 170.810 14.505 171.000 ;
        RECT 14.795 170.830 14.965 171.020 ;
        RECT 18.200 170.810 18.370 171.000 ;
        RECT 24.455 170.830 24.625 171.020 ;
        RECT 24.970 170.860 25.090 170.970 ;
        RECT 27.675 170.810 27.845 171.000 ;
        RECT 29.975 170.830 30.145 171.000 ;
        RECT 30.435 170.810 30.605 171.000 ;
        RECT 32.275 170.855 32.435 170.965 ;
        RECT 34.115 170.830 34.285 171.020 ;
        RECT 35.035 170.810 35.205 171.000 ;
        RECT 35.500 170.830 35.670 171.020 ;
        RECT 37.790 170.810 37.960 171.000 ;
        RECT 40.555 170.810 40.725 171.020 ;
        RECT 41.020 170.810 41.190 171.000 ;
        RECT 43.775 170.830 43.945 171.020 ;
        RECT 44.240 170.830 44.410 171.020 ;
        RECT 44.695 170.810 44.865 171.000 ;
        RECT 49.295 170.830 49.465 171.020 ;
        RECT 49.755 170.830 49.925 171.020 ;
        RECT 51.595 170.865 51.755 170.975 ;
        RECT 54.410 170.860 54.530 170.970 ;
        RECT 55.275 170.830 55.445 171.020 ;
        RECT 58.035 170.810 58.205 171.000 ;
        RECT 59.415 170.810 59.585 171.000 ;
        RECT 60.335 170.855 60.495 170.965 ;
        RECT 60.795 170.810 60.965 171.020 ;
        RECT 64.935 170.810 65.105 171.000 ;
        RECT 66.315 170.810 66.485 171.020 ;
        RECT 67.695 170.810 67.865 171.000 ;
        RECT 68.155 170.830 68.325 171.020 ;
        RECT 71.830 171.000 72.000 171.020 ;
        RECT 71.370 170.810 71.540 171.000 ;
        RECT 71.830 170.830 72.010 171.000 ;
        RECT 72.300 170.830 72.470 171.020 ;
        RECT 77.355 170.830 77.525 171.020 ;
        RECT 78.735 170.830 78.905 171.020 ;
        RECT 71.840 170.810 72.010 170.830 ;
        RECT 78.920 170.810 79.090 171.000 ;
        RECT 82.600 170.830 82.770 171.020 ;
        RECT 83.335 170.830 83.505 171.020 ;
        RECT 84.715 170.830 84.885 171.020 ;
        RECT 88.395 170.830 88.565 171.020 ;
        RECT 88.860 170.830 89.030 171.020 ;
        RECT 89.315 170.810 89.485 171.000 ;
        RECT 89.830 170.860 89.950 170.970 ;
        RECT 92.535 170.810 92.705 171.000 ;
        RECT 93.915 170.810 94.085 171.000 ;
        RECT 95.755 170.810 95.925 171.000 ;
        RECT 96.215 170.810 96.385 171.000 ;
        RECT 96.400 170.830 96.570 171.020 ;
        RECT 97.140 170.830 97.310 171.020 ;
        RECT 97.650 170.860 97.770 170.970 ;
        RECT 99.435 170.810 99.605 171.000 ;
        RECT 104.220 170.830 104.390 171.020 ;
        RECT 104.955 170.810 105.125 171.000 ;
        RECT 105.930 170.860 106.050 170.970 ;
        RECT 106.335 170.810 106.505 171.000 ;
        RECT 110.010 170.810 110.180 171.000 ;
        RECT 110.475 170.810 110.645 171.000 ;
        RECT 114.155 170.830 114.325 171.020 ;
        RECT 115.995 170.830 116.165 171.020 ;
        RECT 116.915 170.810 117.085 171.000 ;
        RECT 118.295 170.810 118.465 171.020 ;
        RECT 11.435 170.000 12.805 170.810 ;
        RECT 13.285 169.900 14.635 170.810 ;
        RECT 14.885 170.130 18.785 170.810 ;
        RECT 18.880 170.130 27.985 170.810 ;
        RECT 17.855 169.900 18.785 170.130 ;
        RECT 28.005 169.940 28.435 170.725 ;
        RECT 28.455 170.130 29.820 170.810 ;
        RECT 30.305 169.900 31.655 170.810 ;
        RECT 32.605 170.130 35.345 170.810 ;
        RECT 35.495 169.900 38.105 170.810 ;
        RECT 38.115 170.000 40.865 170.810 ;
        RECT 40.875 169.900 44.350 170.810 ;
        RECT 44.555 170.130 53.745 170.810 ;
        RECT 49.065 169.910 49.995 170.130 ;
        RECT 52.825 169.900 53.745 170.130 ;
        RECT 53.765 169.940 54.195 170.725 ;
        RECT 54.675 170.000 58.345 170.810 ;
        RECT 58.365 169.900 59.715 170.810 ;
        RECT 60.655 170.130 62.485 170.810 ;
        RECT 62.505 170.130 65.245 170.810 ;
        RECT 61.140 169.900 62.485 170.130 ;
        RECT 65.255 170.000 66.625 170.810 ;
        RECT 66.645 169.900 67.995 170.810 ;
        RECT 68.210 169.900 71.685 170.810 ;
        RECT 71.695 169.900 75.170 170.810 ;
        RECT 75.605 170.130 79.505 170.810 ;
        RECT 78.575 169.900 79.505 170.130 ;
        RECT 79.525 169.940 79.955 170.725 ;
        RECT 80.345 170.130 89.625 170.810 ;
        RECT 80.345 170.010 82.680 170.130 ;
        RECT 80.345 169.900 81.265 170.010 ;
        RECT 87.345 169.910 88.265 170.130 ;
        RECT 90.095 170.000 92.845 170.810 ;
        RECT 92.865 169.900 94.215 170.810 ;
        RECT 94.235 170.000 96.065 170.810 ;
        RECT 96.075 170.030 97.445 170.810 ;
        RECT 97.915 170.000 99.745 170.810 ;
        RECT 99.755 170.000 105.265 170.810 ;
        RECT 105.285 169.940 105.715 170.725 ;
        RECT 106.205 169.900 107.555 170.810 ;
        RECT 107.715 169.900 110.325 170.810 ;
        RECT 110.335 170.030 111.705 170.810 ;
        RECT 111.715 170.000 117.225 170.810 ;
        RECT 117.235 170.000 118.605 170.810 ;
      LAYER nwell ;
        RECT 11.240 166.780 118.800 169.610 ;
      LAYER pwell ;
        RECT 11.435 165.580 12.805 166.390 ;
        RECT 13.735 165.580 15.105 166.360 ;
        RECT 15.125 165.665 15.555 166.450 ;
        RECT 15.575 166.260 16.495 166.490 ;
        RECT 19.325 166.260 20.255 166.480 ;
        RECT 28.895 166.260 29.825 166.490 ;
        RECT 33.035 166.260 33.965 166.490 ;
        RECT 15.575 165.580 24.765 166.260 ;
        RECT 25.925 165.580 29.825 166.260 ;
        RECT 30.065 165.580 33.965 166.260 ;
        RECT 33.975 165.580 35.345 166.360 ;
        RECT 35.355 165.580 40.865 166.390 ;
        RECT 40.885 165.665 41.315 166.450 ;
        RECT 41.335 165.580 45.005 166.390 ;
        RECT 45.155 165.580 47.765 166.490 ;
        RECT 47.775 165.580 49.145 166.390 ;
        RECT 49.155 166.260 50.085 166.490 ;
        RECT 53.665 166.380 54.585 166.490 ;
        RECT 53.665 166.260 56.000 166.380 ;
        RECT 60.665 166.260 61.585 166.480 ;
        RECT 64.360 166.260 65.705 166.490 ;
        RECT 49.155 165.580 53.055 166.260 ;
        RECT 53.665 165.580 62.945 166.260 ;
        RECT 63.875 165.580 65.705 166.260 ;
        RECT 66.645 165.665 67.075 166.450 ;
        RECT 67.580 166.260 68.925 166.490 ;
        RECT 69.420 166.260 70.765 166.490 ;
        RECT 67.095 165.580 68.925 166.260 ;
        RECT 68.935 165.580 70.765 166.260 ;
        RECT 71.235 165.580 76.745 166.390 ;
        RECT 77.125 166.380 78.045 166.490 ;
        RECT 77.125 166.260 79.460 166.380 ;
        RECT 84.125 166.260 85.045 166.480 ;
        RECT 77.125 165.580 86.405 166.260 ;
        RECT 86.875 165.580 92.385 166.390 ;
        RECT 92.405 165.665 92.835 166.450 ;
        RECT 93.970 165.580 97.445 166.490 ;
        RECT 97.915 165.580 100.665 166.390 ;
        RECT 100.675 165.580 106.185 166.390 ;
        RECT 106.195 165.580 111.705 166.390 ;
        RECT 111.715 165.580 117.225 166.390 ;
        RECT 117.235 165.580 118.605 166.390 ;
        RECT 11.575 165.370 11.745 165.580 ;
        RECT 13.415 165.425 13.575 165.535 ;
        RECT 13.875 165.390 14.045 165.580 ;
        RECT 15.255 165.370 15.425 165.560 ;
        RECT 15.715 165.370 15.885 165.560 ;
        RECT 17.095 165.370 17.265 165.560 ;
        RECT 18.750 165.370 18.920 165.560 ;
        RECT 24.455 165.390 24.625 165.580 ;
        RECT 25.375 165.425 25.535 165.535 ;
        RECT 27.675 165.370 27.845 165.560 ;
        RECT 28.595 165.370 28.765 165.560 ;
        RECT 29.240 165.390 29.410 165.580 ;
        RECT 33.380 165.390 33.550 165.580 ;
        RECT 35.035 165.390 35.205 165.580 ;
        RECT 39.635 165.370 39.805 165.560 ;
        RECT 40.555 165.390 40.725 165.580 ;
        RECT 43.310 165.370 43.480 165.560 ;
        RECT 44.695 165.390 44.865 165.580 ;
        RECT 46.990 165.370 47.160 165.560 ;
        RECT 47.450 165.390 47.620 165.580 ;
        RECT 48.375 165.370 48.545 165.560 ;
        RECT 48.835 165.390 49.005 165.580 ;
        RECT 49.570 165.390 49.740 165.580 ;
        RECT 52.055 165.370 52.225 165.560 ;
        RECT 53.435 165.370 53.605 165.560 ;
        RECT 54.410 165.420 54.530 165.530 ;
        RECT 54.820 165.370 54.990 165.560 ;
        RECT 61.900 165.370 62.070 165.560 ;
        RECT 62.635 165.390 62.805 165.580 ;
        RECT 63.555 165.425 63.715 165.535 ;
        RECT 64.015 165.390 64.185 165.580 ;
        RECT 66.315 165.425 66.475 165.535 ;
        RECT 67.235 165.390 67.405 165.580 ;
        RECT 69.075 165.390 69.245 165.580 ;
        RECT 70.970 165.420 71.090 165.530 ;
        RECT 71.835 165.370 72.005 165.560 ;
        RECT 73.215 165.370 73.385 165.560 ;
        RECT 73.730 165.420 73.850 165.530 ;
        RECT 76.435 165.390 76.605 165.580 ;
        RECT 79.195 165.370 79.365 165.560 ;
        RECT 80.170 165.420 80.290 165.530 ;
        RECT 82.875 165.370 83.045 165.560 ;
        RECT 86.095 165.390 86.265 165.580 ;
        RECT 92.075 165.560 92.245 165.580 ;
        RECT 86.610 165.420 86.730 165.530 ;
        RECT 88.395 165.370 88.565 165.560 ;
        RECT 92.070 165.390 92.245 165.560 ;
        RECT 93.455 165.425 93.615 165.535 ;
        RECT 92.070 165.370 92.240 165.390 ;
        RECT 95.750 165.370 95.920 165.560 ;
        RECT 97.130 165.390 97.300 165.580 ;
        RECT 97.650 165.420 97.770 165.530 ;
        RECT 99.430 165.370 99.600 165.560 ;
        RECT 11.435 164.560 12.805 165.370 ;
        RECT 12.815 164.560 15.565 165.370 ;
        RECT 15.585 164.460 16.935 165.370 ;
        RECT 16.955 164.590 18.325 165.370 ;
        RECT 18.335 164.690 22.235 165.370 ;
        RECT 18.335 164.460 19.265 164.690 ;
        RECT 22.475 164.560 27.985 165.370 ;
        RECT 28.005 164.500 28.435 165.285 ;
        RECT 28.455 164.690 37.735 165.370 ;
        RECT 29.815 164.470 30.735 164.690 ;
        RECT 35.400 164.570 37.735 164.690 ;
        RECT 36.815 164.460 37.735 164.570 ;
        RECT 38.115 164.560 39.945 165.370 ;
        RECT 40.150 164.460 43.625 165.370 ;
        RECT 43.830 164.460 47.305 165.370 ;
        RECT 47.315 164.590 48.685 165.370 ;
        RECT 48.790 164.690 52.255 165.370 ;
        RECT 48.790 164.460 49.710 164.690 ;
        RECT 52.375 164.560 53.745 165.370 ;
        RECT 53.765 164.500 54.195 165.285 ;
        RECT 54.675 164.460 58.150 165.370 ;
        RECT 58.585 164.690 62.485 165.370 ;
        RECT 61.555 164.460 62.485 164.690 ;
        RECT 62.865 164.690 72.145 165.370 ;
        RECT 62.865 164.570 65.200 164.690 ;
        RECT 62.865 164.460 63.785 164.570 ;
        RECT 69.865 164.470 70.785 164.690 ;
        RECT 72.155 164.590 73.525 165.370 ;
        RECT 73.995 164.560 79.505 165.370 ;
        RECT 79.525 164.500 79.955 165.285 ;
        RECT 80.435 164.560 83.185 165.370 ;
        RECT 83.195 164.560 88.705 165.370 ;
        RECT 88.910 164.460 92.385 165.370 ;
        RECT 92.590 164.460 96.065 165.370 ;
        RECT 96.270 164.460 99.745 165.370 ;
        RECT 99.900 165.340 100.070 165.560 ;
        RECT 100.355 165.390 100.525 165.580 ;
        RECT 104.955 165.370 105.125 165.560 ;
        RECT 105.875 165.370 106.045 165.580 ;
        RECT 111.395 165.390 111.565 165.580 ;
        RECT 115.995 165.370 116.165 165.560 ;
        RECT 116.915 165.390 117.085 165.580 ;
        RECT 118.295 165.370 118.465 165.580 ;
        RECT 101.560 165.340 102.505 165.370 ;
        RECT 99.755 164.660 102.505 165.340 ;
        RECT 101.560 164.460 102.505 164.660 ;
        RECT 102.515 164.560 105.265 165.370 ;
        RECT 105.285 164.500 105.715 165.285 ;
        RECT 105.745 164.460 107.095 165.370 ;
        RECT 107.115 164.690 116.305 165.370 ;
        RECT 107.115 164.460 108.035 164.690 ;
        RECT 110.865 164.470 111.795 164.690 ;
        RECT 117.235 164.560 118.605 165.370 ;
      LAYER nwell ;
        RECT 11.240 161.340 118.800 164.170 ;
      LAYER pwell ;
        RECT 11.435 160.140 12.805 160.950 ;
        RECT 13.275 160.140 15.105 160.950 ;
        RECT 15.125 160.225 15.555 161.010 ;
        RECT 15.575 160.820 16.495 161.050 ;
        RECT 19.325 160.820 20.255 161.040 ;
        RECT 15.575 160.140 24.765 160.820 ;
        RECT 25.235 160.140 27.985 160.950 ;
        RECT 27.995 160.140 33.505 160.950 ;
        RECT 33.515 160.140 34.885 160.920 ;
        RECT 35.355 160.140 37.185 160.950 ;
        RECT 37.390 160.140 40.865 161.050 ;
        RECT 40.885 160.225 41.315 161.010 ;
        RECT 42.255 160.140 45.730 161.050 ;
        RECT 45.935 160.140 47.305 160.950 ;
        RECT 47.315 160.140 50.525 161.050 ;
        RECT 50.535 160.140 54.010 161.050 ;
        RECT 54.215 160.140 57.690 161.050 ;
        RECT 57.895 160.140 59.725 160.950 ;
        RECT 62.935 160.820 63.865 161.050 ;
        RECT 59.965 160.140 63.865 160.820 ;
        RECT 63.875 160.140 66.625 160.950 ;
        RECT 66.645 160.225 67.075 161.010 ;
        RECT 68.015 160.820 69.360 161.050 ;
        RECT 68.015 160.140 69.845 160.820 ;
        RECT 69.855 160.140 73.525 160.950 ;
        RECT 73.535 160.140 79.045 160.950 ;
        RECT 79.055 160.140 84.565 160.950 ;
        RECT 84.575 160.140 85.945 160.920 ;
        RECT 85.955 160.140 88.705 160.950 ;
        RECT 88.910 160.140 92.385 161.050 ;
        RECT 92.405 160.225 92.835 161.010 ;
        RECT 93.510 160.140 96.985 161.050 ;
        RECT 96.995 160.140 98.825 160.950 ;
        RECT 100.640 160.850 101.585 161.050 ;
        RECT 98.835 160.170 101.585 160.850 ;
        RECT 11.575 159.930 11.745 160.140 ;
        RECT 13.010 159.980 13.130 160.090 ;
        RECT 14.795 159.950 14.965 160.140 ;
        RECT 18.015 159.930 18.185 160.120 ;
        RECT 18.750 159.930 18.920 160.120 ;
        RECT 24.455 159.950 24.625 160.140 ;
        RECT 24.970 159.980 25.090 160.090 ;
        RECT 27.675 159.930 27.845 160.140 ;
        RECT 29.975 159.930 30.145 160.120 ;
        RECT 33.195 159.950 33.365 160.140 ;
        RECT 33.840 159.930 34.010 160.120 ;
        RECT 34.575 159.950 34.745 160.140 ;
        RECT 35.090 159.980 35.210 160.090 ;
        RECT 35.495 159.930 35.665 160.120 ;
        RECT 36.875 159.950 37.045 160.140 ;
        RECT 37.335 159.930 37.505 160.120 ;
        RECT 11.435 159.120 12.805 159.930 ;
        RECT 12.815 159.120 18.325 159.930 ;
        RECT 18.335 159.250 22.235 159.930 ;
        RECT 18.335 159.020 19.265 159.250 ;
        RECT 22.475 159.120 27.985 159.930 ;
        RECT 28.005 159.060 28.435 159.845 ;
        RECT 28.455 159.120 30.285 159.930 ;
        RECT 30.525 159.250 34.425 159.930 ;
        RECT 33.495 159.020 34.425 159.250 ;
        RECT 34.435 159.150 35.805 159.930 ;
        RECT 35.815 159.120 37.645 159.930 ;
        RECT 37.655 159.900 38.600 159.930 ;
        RECT 40.090 159.900 40.260 160.120 ;
        RECT 40.550 159.950 40.720 160.140 ;
        RECT 41.935 159.985 42.095 160.095 ;
        RECT 42.400 159.950 42.570 160.140 ;
        RECT 40.415 159.900 41.360 159.930 ;
        RECT 42.850 159.900 43.020 160.120 ;
        RECT 46.530 159.930 46.700 160.120 ;
        RECT 46.995 159.950 47.165 160.140 ;
        RECT 47.455 159.950 47.625 160.140 ;
        RECT 37.655 159.220 40.405 159.900 ;
        RECT 40.415 159.220 43.165 159.900 ;
        RECT 37.655 159.020 38.600 159.220 ;
        RECT 40.415 159.020 41.360 159.220 ;
        RECT 43.370 159.020 46.845 159.930 ;
        RECT 46.855 159.900 47.800 159.930 ;
        RECT 49.290 159.900 49.460 160.120 ;
        RECT 49.810 159.980 49.930 160.090 ;
        RECT 50.680 159.950 50.850 160.140 ;
        RECT 53.435 159.930 53.605 160.120 ;
        RECT 54.360 159.950 54.530 160.140 ;
        RECT 55.735 159.930 55.905 160.120 ;
        RECT 59.415 159.950 59.585 160.140 ;
        RECT 63.280 159.950 63.450 160.140 ;
        RECT 64.935 159.930 65.105 160.120 ;
        RECT 66.315 159.950 66.485 160.140 ;
        RECT 66.775 159.930 66.945 160.120 ;
        RECT 67.695 159.975 67.855 160.095 ;
        RECT 69.535 159.930 69.705 160.140 ;
        RECT 70.915 159.930 71.085 160.120 ;
        RECT 72.295 159.930 72.465 160.120 ;
        RECT 73.215 159.950 73.385 160.140 ;
        RECT 75.970 159.930 76.140 160.120 ;
        RECT 77.815 159.930 77.985 160.120 ;
        RECT 78.735 159.950 78.905 160.140 ;
        RECT 79.195 159.930 79.365 160.120 ;
        RECT 84.255 159.950 84.425 160.140 ;
        RECT 84.715 159.950 84.885 160.140 ;
        RECT 88.395 159.950 88.565 160.140 ;
        RECT 88.855 159.930 89.025 160.120 ;
        RECT 90.235 159.930 90.405 160.120 ;
        RECT 92.070 159.950 92.240 160.140 ;
        RECT 93.050 159.980 93.170 160.090 ;
        RECT 93.915 159.930 94.085 160.120 ;
        RECT 46.855 159.220 49.605 159.900 ;
        RECT 46.855 159.020 47.800 159.220 ;
        RECT 50.075 159.120 53.745 159.930 ;
        RECT 53.765 159.060 54.195 159.845 ;
        RECT 54.215 159.120 56.045 159.930 ;
        RECT 56.140 159.250 65.245 159.930 ;
        RECT 65.255 159.250 67.085 159.930 ;
        RECT 68.015 159.250 69.845 159.930 ;
        RECT 65.255 159.020 66.600 159.250 ;
        RECT 68.015 159.020 69.360 159.250 ;
        RECT 69.855 159.150 71.225 159.930 ;
        RECT 71.235 159.120 72.605 159.930 ;
        RECT 72.810 159.020 76.285 159.930 ;
        RECT 76.295 159.120 78.125 159.930 ;
        RECT 78.145 159.020 79.495 159.930 ;
        RECT 79.525 159.060 79.955 159.845 ;
        RECT 79.975 159.250 89.165 159.930 ;
        RECT 79.975 159.020 80.895 159.250 ;
        RECT 83.725 159.030 84.655 159.250 ;
        RECT 89.175 159.120 90.545 159.930 ;
        RECT 90.555 159.120 94.225 159.930 ;
        RECT 94.235 159.900 95.180 159.930 ;
        RECT 96.670 159.900 96.840 160.140 ;
        RECT 97.140 159.930 97.310 160.120 ;
        RECT 98.515 159.950 98.685 160.140 ;
        RECT 98.980 159.950 99.150 160.170 ;
        RECT 100.640 160.140 101.585 160.170 ;
        RECT 101.595 160.140 105.070 161.050 ;
        RECT 108.935 160.820 109.865 161.050 ;
        RECT 105.965 160.140 109.865 160.820 ;
        RECT 110.345 160.140 111.695 161.050 ;
        RECT 112.635 160.140 114.005 160.920 ;
        RECT 114.015 160.140 115.385 160.920 ;
        RECT 115.395 160.140 117.225 160.950 ;
        RECT 117.235 160.140 118.605 160.950 ;
        RECT 101.275 159.975 101.435 160.085 ;
        RECT 101.740 159.930 101.910 160.140 ;
        RECT 105.470 159.980 105.590 160.090 ;
        RECT 106.795 159.930 106.965 160.120 ;
        RECT 109.280 159.950 109.450 160.140 ;
        RECT 110.070 159.980 110.190 160.090 ;
        RECT 110.475 159.950 110.645 160.140 ;
        RECT 112.315 159.985 112.475 160.095 ;
        RECT 112.775 159.950 112.945 160.140 ;
        RECT 114.155 159.950 114.325 160.140 ;
        RECT 116.455 159.930 116.625 160.120 ;
        RECT 116.915 160.090 117.085 160.140 ;
        RECT 116.915 159.980 117.090 160.090 ;
        RECT 116.915 159.950 117.085 159.980 ;
        RECT 118.295 159.930 118.465 160.140 ;
        RECT 94.235 159.220 96.985 159.900 ;
        RECT 94.235 159.020 95.180 159.220 ;
        RECT 96.995 159.020 100.470 159.930 ;
        RECT 101.595 159.020 105.070 159.930 ;
        RECT 105.285 159.060 105.715 159.845 ;
        RECT 105.735 159.120 107.105 159.930 ;
        RECT 107.485 159.250 116.765 159.930 ;
        RECT 107.485 159.130 109.820 159.250 ;
        RECT 107.485 159.020 108.405 159.130 ;
        RECT 114.485 159.030 115.405 159.250 ;
        RECT 117.235 159.120 118.605 159.930 ;
      LAYER nwell ;
        RECT 11.240 155.900 118.800 158.730 ;
      LAYER pwell ;
        RECT 11.435 154.700 12.805 155.510 ;
        RECT 13.275 154.700 15.105 155.510 ;
        RECT 15.125 154.785 15.555 155.570 ;
        RECT 15.575 154.700 17.405 155.510 ;
        RECT 17.425 154.700 18.775 155.610 ;
        RECT 18.795 154.700 22.465 155.510 ;
        RECT 22.475 154.700 23.845 155.480 ;
        RECT 23.855 154.700 25.225 155.510 ;
        RECT 25.245 154.700 26.595 155.610 ;
        RECT 26.615 155.380 27.535 155.610 ;
        RECT 30.365 155.380 31.295 155.600 ;
        RECT 26.615 154.700 35.805 155.380 ;
        RECT 35.815 154.700 37.185 155.510 ;
        RECT 37.195 154.700 40.865 155.510 ;
        RECT 40.885 154.785 41.315 155.570 ;
        RECT 41.795 154.700 44.545 155.510 ;
        RECT 44.555 155.410 45.500 155.610 ;
        RECT 44.555 154.730 47.305 155.410 ;
        RECT 44.555 154.700 45.500 154.730 ;
        RECT 11.575 154.490 11.745 154.700 ;
        RECT 13.010 154.540 13.130 154.650 ;
        RECT 14.795 154.510 14.965 154.700 ;
        RECT 17.095 154.510 17.265 154.700 ;
        RECT 18.475 154.510 18.645 154.700 ;
        RECT 22.155 154.490 22.325 154.700 ;
        RECT 22.615 154.490 22.785 154.680 ;
        RECT 23.535 154.510 23.705 154.700 ;
        RECT 24.915 154.510 25.085 154.700 ;
        RECT 25.375 154.510 25.545 154.700 ;
        RECT 27.675 154.490 27.845 154.680 ;
        RECT 28.870 154.490 29.040 154.680 ;
        RECT 32.790 154.540 32.910 154.650 ;
        RECT 35.495 154.490 35.665 154.700 ;
        RECT 35.960 154.490 36.130 154.680 ;
        RECT 36.875 154.510 37.045 154.700 ;
        RECT 39.640 154.490 39.810 154.680 ;
        RECT 40.555 154.510 40.725 154.700 ;
        RECT 41.530 154.540 41.650 154.650 ;
        RECT 43.775 154.490 43.945 154.680 ;
        RECT 44.235 154.510 44.405 154.700 ;
        RECT 46.990 154.510 47.160 154.730 ;
        RECT 47.785 154.700 49.135 155.610 ;
        RECT 52.355 155.380 53.285 155.610 ;
        RECT 49.385 154.700 53.285 155.380 ;
        RECT 53.295 154.700 56.770 155.610 ;
        RECT 57.345 155.500 58.265 155.610 ;
        RECT 57.345 155.380 59.680 155.500 ;
        RECT 64.345 155.380 65.265 155.600 ;
        RECT 57.345 154.700 66.625 155.380 ;
        RECT 66.645 154.785 67.075 155.570 ;
        RECT 67.095 154.700 69.815 155.610 ;
        RECT 69.855 154.700 72.595 155.380 ;
        RECT 72.810 154.700 76.285 155.610 ;
        RECT 76.755 154.700 80.425 155.510 ;
        RECT 83.635 155.380 84.565 155.610 ;
        RECT 80.665 154.700 84.565 155.380 ;
        RECT 85.035 154.700 86.865 155.510 ;
        RECT 86.875 154.700 92.385 155.510 ;
        RECT 92.405 154.785 92.835 155.570 ;
        RECT 92.855 154.700 96.525 155.510 ;
        RECT 96.535 155.410 97.480 155.610 ;
        RECT 96.535 154.730 99.285 155.410 ;
        RECT 96.535 154.700 97.480 154.730 ;
        RECT 47.510 154.540 47.630 154.650 ;
        RECT 48.835 154.510 49.005 154.700 ;
        RECT 52.700 154.510 52.870 154.700 ;
        RECT 53.440 154.680 53.610 154.700 ;
        RECT 53.435 154.510 53.610 154.680 ;
        RECT 53.435 154.490 53.605 154.510 ;
        RECT 55.275 154.490 55.445 154.680 ;
        RECT 58.955 154.490 59.125 154.680 ;
        RECT 59.415 154.490 59.585 154.680 ;
        RECT 61.255 154.490 61.425 154.680 ;
        RECT 63.150 154.540 63.270 154.650 ;
        RECT 65.855 154.490 66.025 154.680 ;
        RECT 66.315 154.490 66.485 154.700 ;
        RECT 67.235 154.510 67.405 154.700 ;
        RECT 68.155 154.490 68.325 154.680 ;
        RECT 69.995 154.490 70.165 154.700 ;
        RECT 75.050 154.490 75.220 154.680 ;
        RECT 75.570 154.540 75.690 154.650 ;
        RECT 75.970 154.510 76.140 154.700 ;
        RECT 76.490 154.540 76.610 154.650 ;
        RECT 79.195 154.490 79.365 154.680 ;
        RECT 80.115 154.510 80.285 154.700 ;
        RECT 83.980 154.510 84.150 154.700 ;
        RECT 84.770 154.540 84.890 154.650 ;
        RECT 86.555 154.510 86.725 154.700 ;
        RECT 89.315 154.490 89.485 154.680 ;
        RECT 89.830 154.540 89.950 154.650 ;
        RECT 92.075 154.510 92.245 154.700 ;
        RECT 11.435 153.680 12.805 154.490 ;
        RECT 13.275 153.810 22.465 154.490 ;
        RECT 22.585 153.810 26.050 154.490 ;
        RECT 13.275 153.580 14.195 153.810 ;
        RECT 17.025 153.590 17.955 153.810 ;
        RECT 25.130 153.580 26.050 153.810 ;
        RECT 26.155 153.680 27.985 154.490 ;
        RECT 28.005 153.620 28.435 154.405 ;
        RECT 28.455 153.810 32.355 154.490 ;
        RECT 28.455 153.580 29.385 153.810 ;
        RECT 33.055 153.680 35.805 154.490 ;
        RECT 35.815 153.580 39.290 154.490 ;
        RECT 39.495 153.580 42.105 154.490 ;
        RECT 42.255 153.680 44.085 154.490 ;
        RECT 44.465 153.810 53.745 154.490 ;
        RECT 44.465 153.690 46.800 153.810 ;
        RECT 44.465 153.580 45.385 153.690 ;
        RECT 51.465 153.590 52.385 153.810 ;
        RECT 53.765 153.620 54.195 154.405 ;
        RECT 54.215 153.710 55.585 154.490 ;
        RECT 55.595 153.680 59.265 154.490 ;
        RECT 59.275 153.810 61.105 154.490 ;
        RECT 61.115 153.810 62.945 154.490 ;
        RECT 63.425 153.810 66.165 154.490 ;
        RECT 66.175 153.810 68.005 154.490 ;
        RECT 68.015 153.810 69.845 154.490 ;
        RECT 69.855 153.810 71.685 154.490 ;
        RECT 59.760 153.580 61.105 153.810 ;
        RECT 61.600 153.580 62.945 153.810 ;
        RECT 66.660 153.580 68.005 153.810 ;
        RECT 68.500 153.580 69.845 153.810 ;
        RECT 70.340 153.580 71.685 153.810 ;
        RECT 71.890 153.580 75.365 154.490 ;
        RECT 75.835 153.680 79.505 154.490 ;
        RECT 79.525 153.620 79.955 154.405 ;
        RECT 80.345 153.810 89.625 154.490 ;
        RECT 90.095 154.460 91.040 154.490 ;
        RECT 92.530 154.460 92.700 154.680 ;
        RECT 93.000 154.490 93.170 154.680 ;
        RECT 96.215 154.510 96.385 154.700 ;
        RECT 98.970 154.680 99.140 154.730 ;
        RECT 99.295 154.700 101.125 155.510 ;
        RECT 101.135 154.700 104.610 155.610 ;
        RECT 105.275 154.700 107.105 155.510 ;
        RECT 110.315 155.380 111.245 155.610 ;
        RECT 107.345 154.700 111.245 155.380 ;
        RECT 111.715 154.700 117.225 155.510 ;
        RECT 117.235 154.700 118.605 155.510 ;
        RECT 96.730 154.540 96.850 154.650 ;
        RECT 98.515 154.490 98.685 154.680 ;
        RECT 98.970 154.510 99.150 154.680 ;
        RECT 100.815 154.510 100.985 154.700 ;
        RECT 101.280 154.510 101.450 154.700 ;
        RECT 104.955 154.650 105.125 154.680 ;
        RECT 104.955 154.540 105.130 154.650 ;
        RECT 98.980 154.490 99.150 154.510 ;
        RECT 104.955 154.490 105.125 154.540 ;
        RECT 106.795 154.490 106.965 154.700 ;
        RECT 110.660 154.490 110.830 154.700 ;
        RECT 111.450 154.540 111.570 154.650 ;
        RECT 113.690 154.490 113.860 154.680 ;
        RECT 114.210 154.540 114.330 154.650 ;
        RECT 116.915 154.490 117.085 154.700 ;
        RECT 118.295 154.490 118.465 154.700 ;
        RECT 80.345 153.690 82.680 153.810 ;
        RECT 80.345 153.580 81.265 153.690 ;
        RECT 87.345 153.590 88.265 153.810 ;
        RECT 90.095 153.780 92.845 154.460 ;
        RECT 90.095 153.580 91.040 153.780 ;
        RECT 92.855 153.580 96.330 154.490 ;
        RECT 96.995 153.680 98.825 154.490 ;
        RECT 98.835 153.580 102.310 154.490 ;
        RECT 102.515 153.680 105.265 154.490 ;
        RECT 105.285 153.620 105.715 154.405 ;
        RECT 105.735 153.680 107.105 154.490 ;
        RECT 107.345 153.810 111.245 154.490 ;
        RECT 110.315 153.580 111.245 153.810 ;
        RECT 111.395 153.580 114.005 154.490 ;
        RECT 114.475 153.680 117.225 154.490 ;
        RECT 117.235 153.680 118.605 154.490 ;
      LAYER nwell ;
        RECT 11.240 150.460 118.800 153.290 ;
      LAYER pwell ;
        RECT 11.435 149.260 12.805 150.070 ;
        RECT 13.275 149.260 15.105 150.070 ;
        RECT 15.125 149.345 15.555 150.130 ;
        RECT 16.035 149.260 17.865 150.070 ;
        RECT 21.075 149.940 22.005 150.170 ;
        RECT 18.105 149.260 22.005 149.940 ;
        RECT 22.025 149.260 23.375 150.170 ;
        RECT 23.395 149.940 24.315 150.170 ;
        RECT 27.145 149.940 28.075 150.160 ;
        RECT 23.395 149.260 32.585 149.940 ;
        RECT 33.055 149.260 34.885 150.070 ;
        RECT 34.895 149.260 38.370 150.170 ;
        RECT 39.035 149.260 40.865 150.070 ;
        RECT 40.885 149.345 41.315 150.130 ;
        RECT 41.335 149.260 44.085 150.070 ;
        RECT 44.095 149.260 47.570 150.170 ;
        RECT 47.775 149.260 49.605 150.070 ;
        RECT 52.815 149.940 53.745 150.170 ;
        RECT 49.845 149.260 53.745 149.940 ;
        RECT 53.755 149.260 57.425 150.070 ;
        RECT 57.435 149.260 62.945 150.070 ;
        RECT 62.965 149.260 64.315 150.170 ;
        RECT 64.795 149.260 66.625 150.070 ;
        RECT 66.645 149.345 67.075 150.130 ;
        RECT 67.555 149.260 71.225 150.070 ;
        RECT 71.430 149.260 74.905 150.170 ;
        RECT 74.915 149.260 78.390 150.170 ;
        RECT 78.595 149.260 80.425 150.070 ;
        RECT 83.635 149.940 84.565 150.170 ;
        RECT 80.665 149.260 84.565 149.940 ;
        RECT 85.045 149.260 86.395 150.170 ;
        RECT 86.415 149.260 87.785 150.040 ;
        RECT 88.715 149.260 92.385 150.070 ;
        RECT 92.405 149.345 92.835 150.130 ;
        RECT 93.775 149.260 99.285 150.070 ;
        RECT 101.100 149.970 102.045 150.170 ;
        RECT 99.295 149.290 102.045 149.970 ;
        RECT 11.575 149.050 11.745 149.260 ;
        RECT 13.010 149.100 13.130 149.210 ;
        RECT 13.415 149.095 13.575 149.205 ;
        RECT 14.795 149.070 14.965 149.260 ;
        RECT 15.770 149.100 15.890 149.210 ;
        RECT 17.555 149.070 17.725 149.260 ;
        RECT 21.420 149.070 21.590 149.260 ;
        RECT 22.155 149.070 22.325 149.260 ;
        RECT 22.615 149.050 22.785 149.240 ;
        RECT 23.130 149.100 23.250 149.210 ;
        RECT 23.810 149.050 23.980 149.240 ;
        RECT 27.730 149.100 27.850 149.210 ;
        RECT 29.515 149.050 29.685 149.240 ;
        RECT 29.975 149.050 30.145 149.240 ;
        RECT 32.275 149.070 32.445 149.260 ;
        RECT 34.575 149.240 34.745 149.260 ;
        RECT 32.790 149.100 32.910 149.210 ;
        RECT 34.570 149.070 34.745 149.240 ;
        RECT 35.040 149.070 35.210 149.260 ;
        RECT 40.555 149.240 40.725 149.260 ;
        RECT 34.570 149.050 34.740 149.070 ;
        RECT 38.250 149.050 38.420 149.240 ;
        RECT 38.770 149.100 38.890 149.210 ;
        RECT 40.095 149.050 40.265 149.240 ;
        RECT 40.555 149.070 40.730 149.240 ;
        RECT 43.775 149.070 43.945 149.260 ;
        RECT 44.240 149.070 44.410 149.260 ;
        RECT 49.295 149.070 49.465 149.260 ;
        RECT 53.160 149.070 53.330 149.260 ;
        RECT 40.560 149.050 40.730 149.070 ;
        RECT 53.435 149.050 53.605 149.240 ;
        RECT 55.275 149.050 55.445 149.240 ;
        RECT 57.115 149.050 57.285 149.260 ;
        RECT 57.575 149.050 57.745 149.240 ;
        RECT 59.415 149.095 59.575 149.205 ;
        RECT 62.635 149.070 62.805 149.260 ;
        RECT 64.015 149.070 64.185 149.260 ;
        RECT 66.315 149.240 66.485 149.260 ;
        RECT 64.530 149.100 64.650 149.210 ;
        RECT 64.935 149.050 65.105 149.240 ;
        RECT 66.305 149.070 66.485 149.240 ;
        RECT 67.290 149.100 67.410 149.210 ;
        RECT 70.915 149.070 71.085 149.260 ;
        RECT 66.305 149.050 66.475 149.070 ;
        RECT 71.835 149.050 72.005 149.240 ;
        RECT 11.435 148.240 12.805 149.050 ;
        RECT 13.735 148.370 22.925 149.050 ;
        RECT 23.395 148.370 27.295 149.050 ;
        RECT 13.735 148.140 14.655 148.370 ;
        RECT 17.485 148.150 18.415 148.370 ;
        RECT 23.395 148.140 24.325 148.370 ;
        RECT 28.005 148.180 28.435 148.965 ;
        RECT 28.455 148.240 29.825 149.050 ;
        RECT 29.835 148.270 31.205 149.050 ;
        RECT 31.410 148.140 34.885 149.050 ;
        RECT 35.090 148.140 38.565 149.050 ;
        RECT 38.575 148.240 40.405 149.050 ;
        RECT 40.415 148.140 43.890 149.050 ;
        RECT 44.465 148.370 53.745 149.050 ;
        RECT 44.465 148.250 46.800 148.370 ;
        RECT 44.465 148.140 45.385 148.250 ;
        RECT 51.465 148.150 52.385 148.370 ;
        RECT 53.765 148.180 54.195 148.965 ;
        RECT 54.215 148.270 55.585 149.050 ;
        RECT 55.595 148.240 57.425 149.050 ;
        RECT 57.445 148.140 58.795 149.050 ;
        RECT 59.735 148.240 65.245 149.050 ;
        RECT 65.255 148.270 66.625 149.050 ;
        RECT 66.635 148.240 72.145 149.050 ;
        RECT 72.155 149.020 73.100 149.050 ;
        RECT 74.590 149.020 74.760 149.260 ;
        RECT 75.060 149.070 75.230 149.260 ;
        RECT 75.515 149.095 75.675 149.205 ;
        RECT 79.195 149.050 79.365 149.240 ;
        RECT 80.115 149.070 80.285 149.260 ;
        RECT 80.575 149.095 80.735 149.205 ;
        RECT 83.980 149.070 84.150 149.260 ;
        RECT 84.770 149.100 84.890 149.210 ;
        RECT 86.095 149.070 86.265 149.260 ;
        RECT 86.555 149.070 86.725 149.260 ;
        RECT 88.395 149.105 88.555 149.215 ;
        RECT 90.235 149.050 90.405 149.240 ;
        RECT 92.075 149.070 92.245 149.260 ;
        RECT 93.455 149.105 93.615 149.215 ;
        RECT 93.915 149.050 94.085 149.240 ;
        RECT 97.780 149.050 97.950 149.240 ;
        RECT 98.975 149.070 99.145 149.260 ;
        RECT 99.440 149.070 99.610 149.290 ;
        RECT 101.100 149.260 102.045 149.290 ;
        RECT 102.055 149.260 104.805 150.070 ;
        RECT 104.825 149.260 106.175 150.170 ;
        RECT 106.565 150.060 107.485 150.170 ;
        RECT 106.565 149.940 108.900 150.060 ;
        RECT 113.565 149.940 114.485 150.160 ;
        RECT 106.565 149.260 115.845 149.940 ;
        RECT 115.855 149.260 117.225 150.040 ;
        RECT 117.235 149.260 118.605 150.070 ;
        RECT 101.920 149.050 102.090 149.240 ;
        RECT 104.495 149.070 104.665 149.260 ;
        RECT 104.955 149.050 105.125 149.260 ;
        RECT 105.930 149.100 106.050 149.210 ;
        RECT 106.335 149.050 106.505 149.240 ;
        RECT 115.535 149.070 115.705 149.260 ;
        RECT 116.915 149.050 117.085 149.260 ;
        RECT 118.295 149.050 118.465 149.260 ;
        RECT 72.155 148.340 74.905 149.020 ;
        RECT 72.155 148.140 73.100 148.340 ;
        RECT 75.835 148.240 79.505 149.050 ;
        RECT 79.525 148.180 79.955 148.965 ;
        RECT 81.265 148.370 90.545 149.050 ;
        RECT 81.265 148.250 83.600 148.370 ;
        RECT 81.265 148.140 82.185 148.250 ;
        RECT 88.265 148.150 89.185 148.370 ;
        RECT 90.555 148.240 94.225 149.050 ;
        RECT 94.465 148.370 98.365 149.050 ;
        RECT 98.605 148.370 102.505 149.050 ;
        RECT 97.435 148.140 98.365 148.370 ;
        RECT 101.575 148.140 102.505 148.370 ;
        RECT 102.515 148.240 105.265 149.050 ;
        RECT 105.285 148.180 105.715 148.965 ;
        RECT 106.205 148.140 107.555 149.050 ;
        RECT 107.945 148.370 117.225 149.050 ;
        RECT 107.945 148.250 110.280 148.370 ;
        RECT 107.945 148.140 108.865 148.250 ;
        RECT 114.945 148.150 115.865 148.370 ;
        RECT 117.235 148.240 118.605 149.050 ;
      LAYER nwell ;
        RECT 11.240 145.020 118.800 147.850 ;
      LAYER pwell ;
        RECT 11.435 143.820 12.805 144.630 ;
        RECT 13.745 143.820 15.095 144.730 ;
        RECT 15.125 143.905 15.555 144.690 ;
        RECT 15.585 143.820 16.935 144.730 ;
        RECT 16.955 143.820 18.325 144.600 ;
        RECT 18.335 144.500 19.255 144.730 ;
        RECT 22.085 144.500 23.015 144.720 ;
        RECT 18.335 143.820 27.525 144.500 ;
        RECT 28.455 143.820 32.125 144.630 ;
        RECT 32.135 144.530 33.080 144.730 ;
        RECT 32.135 143.850 34.885 144.530 ;
        RECT 32.135 143.820 33.080 143.850 ;
        RECT 11.575 143.610 11.745 143.820 ;
        RECT 13.010 143.660 13.130 143.770 ;
        RECT 13.415 143.610 13.585 143.800 ;
        RECT 14.795 143.630 14.965 143.820 ;
        RECT 15.715 143.630 15.885 143.820 ;
        RECT 17.095 143.630 17.265 143.820 ;
        RECT 18.475 143.610 18.645 143.800 ;
        RECT 19.210 143.610 19.380 143.800 ;
        RECT 23.995 143.610 24.165 143.800 ;
        RECT 24.455 143.610 24.625 143.800 ;
        RECT 25.890 143.660 26.010 143.770 ;
        RECT 27.215 143.630 27.385 143.820 ;
        RECT 27.675 143.610 27.845 143.800 ;
        RECT 28.135 143.665 28.295 143.775 ;
        RECT 28.650 143.660 28.770 143.770 ;
        RECT 31.815 143.630 31.985 143.820 ;
        RECT 32.275 143.610 32.445 143.800 ;
        RECT 11.435 142.800 12.805 143.610 ;
        RECT 13.385 142.930 16.850 143.610 ;
        RECT 15.930 142.700 16.850 142.930 ;
        RECT 16.955 142.800 18.785 143.610 ;
        RECT 18.795 142.930 22.695 143.610 ;
        RECT 18.795 142.700 19.725 142.930 ;
        RECT 22.935 142.800 24.305 143.610 ;
        RECT 24.315 142.830 25.685 143.610 ;
        RECT 26.155 142.800 27.985 143.610 ;
        RECT 28.005 142.740 28.435 143.525 ;
        RECT 28.915 142.800 32.585 143.610 ;
        RECT 32.740 143.580 32.910 143.800 ;
        RECT 34.570 143.630 34.740 143.850 ;
        RECT 34.895 143.820 38.370 144.730 ;
        RECT 39.035 143.820 40.865 144.630 ;
        RECT 40.885 143.905 41.315 144.690 ;
        RECT 41.795 143.820 44.545 144.630 ;
        RECT 44.555 143.820 48.030 144.730 ;
        RECT 48.695 143.820 50.525 144.630 ;
        RECT 50.545 143.820 51.895 144.730 ;
        RECT 52.375 143.820 54.205 144.630 ;
        RECT 54.225 143.820 55.575 144.730 ;
        RECT 55.965 144.620 56.885 144.730 ;
        RECT 55.965 144.500 58.300 144.620 ;
        RECT 62.965 144.500 63.885 144.720 ;
        RECT 55.965 143.820 65.245 144.500 ;
        RECT 65.255 143.820 66.625 144.630 ;
        RECT 66.645 143.905 67.075 144.690 ;
        RECT 67.555 143.820 71.225 144.630 ;
        RECT 71.235 144.530 72.180 144.730 ;
        RECT 71.235 143.850 73.985 144.530 ;
        RECT 71.235 143.820 72.180 143.850 ;
        RECT 35.040 143.630 35.210 143.820 ;
        RECT 34.400 143.580 35.345 143.610 ;
        RECT 32.595 142.900 35.345 143.580 ;
        RECT 34.400 142.700 35.345 142.900 ;
        RECT 35.355 143.580 36.300 143.610 ;
        RECT 37.790 143.580 37.960 143.800 ;
        RECT 38.310 143.660 38.430 143.770 ;
        RECT 38.770 143.660 38.890 143.770 ;
        RECT 40.095 143.610 40.265 143.800 ;
        RECT 40.555 143.630 40.725 143.820 ;
        RECT 41.530 143.660 41.650 143.770 ;
        RECT 44.235 143.630 44.405 143.820 ;
        RECT 44.700 143.630 44.870 143.820 ;
        RECT 45.615 143.610 45.785 143.800 ;
        RECT 46.080 143.610 46.250 143.800 ;
        RECT 48.430 143.660 48.550 143.770 ;
        RECT 50.215 143.630 50.385 143.820 ;
        RECT 51.595 143.630 51.765 143.820 ;
        RECT 52.110 143.660 52.230 143.770 ;
        RECT 53.160 143.610 53.330 143.800 ;
        RECT 53.895 143.630 54.065 143.820 ;
        RECT 54.355 143.630 54.525 143.820 ;
        RECT 55.275 143.610 55.445 143.800 ;
        RECT 64.935 143.610 65.105 143.820 ;
        RECT 66.315 143.630 66.485 143.820 ;
        RECT 67.290 143.660 67.410 143.770 ;
        RECT 70.455 143.610 70.625 143.800 ;
        RECT 70.915 143.630 71.085 143.820 ;
        RECT 73.670 143.630 73.840 143.850 ;
        RECT 73.995 143.820 77.470 144.730 ;
        RECT 77.675 143.820 81.345 144.630 ;
        RECT 84.555 144.500 85.485 144.730 ;
        RECT 81.585 143.820 85.485 144.500 ;
        RECT 85.505 143.820 86.855 144.730 ;
        RECT 86.875 143.820 88.245 144.600 ;
        RECT 88.715 143.820 92.385 144.630 ;
        RECT 92.405 143.905 92.835 144.690 ;
        RECT 93.785 143.820 95.135 144.730 ;
        RECT 95.525 144.620 96.445 144.730 ;
        RECT 95.525 144.500 97.860 144.620 ;
        RECT 102.525 144.500 103.445 144.720 ;
        RECT 95.525 143.820 104.805 144.500 ;
        RECT 104.815 143.820 106.185 144.630 ;
        RECT 109.395 144.500 110.325 144.730 ;
        RECT 106.425 143.820 110.325 144.500 ;
        RECT 111.255 143.820 112.625 144.600 ;
        RECT 113.555 143.820 117.225 144.630 ;
        RECT 117.235 143.820 118.605 144.630 ;
        RECT 74.140 143.800 74.310 143.820 ;
        RECT 74.130 143.630 74.310 143.800 ;
        RECT 74.130 143.610 74.300 143.630 ;
        RECT 74.600 143.610 74.770 143.800 ;
        RECT 79.195 143.610 79.365 143.800 ;
        RECT 81.035 143.630 81.205 143.820 ;
        RECT 82.415 143.610 82.585 143.800 ;
        RECT 84.900 143.630 85.070 143.820 ;
        RECT 86.280 143.610 86.450 143.800 ;
        RECT 86.555 143.630 86.725 143.820 ;
        RECT 87.015 143.610 87.185 143.820 ;
        RECT 88.450 143.660 88.570 143.770 ;
        RECT 91.615 143.610 91.785 143.800 ;
        RECT 92.075 143.630 92.245 143.820 ;
        RECT 93.455 143.665 93.615 143.775 ;
        RECT 93.915 143.630 94.085 143.820 ;
        RECT 101.275 143.610 101.445 143.800 ;
        RECT 101.735 143.610 101.905 143.800 ;
        RECT 103.170 143.660 103.290 143.770 ;
        RECT 104.495 143.630 104.665 143.820 ;
        RECT 104.955 143.610 105.125 143.800 ;
        RECT 105.875 143.770 106.045 143.820 ;
        RECT 105.875 143.660 106.050 143.770 ;
        RECT 105.875 143.630 106.045 143.660 ;
        RECT 109.740 143.630 109.910 143.820 ;
        RECT 110.935 143.665 111.095 143.775 ;
        RECT 111.395 143.610 111.565 143.820 ;
        RECT 113.235 143.665 113.395 143.775 ;
        RECT 116.915 143.610 117.085 143.820 ;
        RECT 118.295 143.610 118.465 143.820 ;
        RECT 35.355 142.900 38.105 143.580 ;
        RECT 35.355 142.700 36.300 142.900 ;
        RECT 38.575 142.800 40.405 143.610 ;
        RECT 40.415 142.800 45.925 143.610 ;
        RECT 45.935 142.700 49.410 143.610 ;
        RECT 49.845 142.930 53.745 143.610 ;
        RECT 52.815 142.700 53.745 142.930 ;
        RECT 53.765 142.740 54.195 143.525 ;
        RECT 54.215 142.800 55.585 143.610 ;
        RECT 55.965 142.930 65.245 143.610 ;
        RECT 55.965 142.810 58.300 142.930 ;
        RECT 55.965 142.700 56.885 142.810 ;
        RECT 62.965 142.710 63.885 142.930 ;
        RECT 65.255 142.800 70.765 143.610 ;
        RECT 70.970 142.700 74.445 143.610 ;
        RECT 74.455 142.700 77.930 143.610 ;
        RECT 78.135 142.800 79.505 143.610 ;
        RECT 79.525 142.740 79.955 143.525 ;
        RECT 79.975 142.800 82.725 143.610 ;
        RECT 82.965 142.930 86.865 143.610 ;
        RECT 85.935 142.700 86.865 142.930 ;
        RECT 86.875 142.830 88.245 143.610 ;
        RECT 88.255 142.800 91.925 143.610 ;
        RECT 92.305 142.930 101.585 143.610 ;
        RECT 92.305 142.810 94.640 142.930 ;
        RECT 92.305 142.700 93.225 142.810 ;
        RECT 99.305 142.710 100.225 142.930 ;
        RECT 101.595 142.830 102.965 143.610 ;
        RECT 103.435 142.800 105.265 143.610 ;
        RECT 105.285 142.740 105.715 143.525 ;
        RECT 106.195 142.800 111.705 143.610 ;
        RECT 111.715 142.800 117.225 143.610 ;
        RECT 117.235 142.800 118.605 143.610 ;
      LAYER nwell ;
        RECT 11.240 139.580 118.800 142.410 ;
      LAYER pwell ;
        RECT 11.435 138.380 12.805 139.190 ;
        RECT 13.275 138.380 15.105 139.190 ;
        RECT 15.125 138.465 15.555 139.250 ;
        RECT 16.035 138.380 21.545 139.190 ;
        RECT 21.555 138.380 27.065 139.190 ;
        RECT 27.075 138.380 32.585 139.190 ;
        RECT 32.595 139.090 33.540 139.290 ;
        RECT 35.355 139.090 36.300 139.290 ;
        RECT 32.595 138.410 35.345 139.090 ;
        RECT 35.355 138.410 38.105 139.090 ;
        RECT 32.595 138.380 33.540 138.410 ;
        RECT 11.575 138.170 11.745 138.380 ;
        RECT 13.010 138.220 13.130 138.330 ;
        RECT 14.795 138.190 14.965 138.380 ;
        RECT 15.770 138.220 15.890 138.330 ;
        RECT 21.235 138.190 21.405 138.380 ;
        RECT 22.615 138.170 22.785 138.360 ;
        RECT 23.130 138.220 23.250 138.330 ;
        RECT 25.835 138.170 26.005 138.360 ;
        RECT 26.755 138.190 26.925 138.380 ;
        RECT 27.215 138.170 27.385 138.360 ;
        RECT 27.730 138.220 27.850 138.330 ;
        RECT 29.515 138.170 29.685 138.360 ;
        RECT 29.975 138.190 30.145 138.360 ;
        RECT 32.275 138.190 32.445 138.380 ;
        RECT 35.030 138.190 35.200 138.410 ;
        RECT 35.355 138.380 36.300 138.410 ;
        RECT 36.415 138.190 36.585 138.360 ;
        RECT 36.875 138.190 37.045 138.360 ;
        RECT 37.790 138.190 37.960 138.410 ;
        RECT 38.115 138.380 40.865 139.190 ;
        RECT 40.885 138.465 41.315 139.250 ;
        RECT 41.335 138.380 43.165 139.190 ;
        RECT 43.175 139.090 44.120 139.290 ;
        RECT 43.175 138.410 45.925 139.090 ;
        RECT 43.175 138.380 44.120 138.410 ;
        RECT 40.555 138.190 40.725 138.380 ;
        RECT 29.995 138.170 30.145 138.190 ;
        RECT 32.295 138.170 32.445 138.190 ;
        RECT 36.415 138.170 36.565 138.190 ;
        RECT 11.435 137.360 12.805 138.170 ;
        RECT 13.645 137.490 22.925 138.170 ;
        RECT 13.645 137.370 15.980 137.490 ;
        RECT 13.645 137.260 14.565 137.370 ;
        RECT 20.645 137.270 21.565 137.490 ;
        RECT 23.395 137.360 26.145 138.170 ;
        RECT 26.155 137.390 27.525 138.170 ;
        RECT 28.005 137.300 28.435 138.085 ;
        RECT 28.455 137.360 29.825 138.170 ;
        RECT 29.995 137.350 31.925 138.170 ;
        RECT 32.295 137.350 34.225 138.170 ;
        RECT 30.975 137.260 31.925 137.350 ;
        RECT 33.275 137.260 34.225 137.350 ;
        RECT 34.635 137.350 36.565 138.170 ;
        RECT 36.895 138.170 37.045 138.190 ;
        RECT 42.395 138.170 42.565 138.360 ;
        RECT 42.855 138.190 43.025 138.380 ;
        RECT 45.610 138.190 45.780 138.410 ;
        RECT 45.935 138.380 49.410 139.290 ;
        RECT 49.615 138.380 53.090 139.290 ;
        RECT 53.295 138.380 56.045 139.190 ;
        RECT 59.255 139.060 60.185 139.290 ;
        RECT 56.285 138.380 60.185 139.060 ;
        RECT 60.195 138.380 61.565 139.160 ;
        RECT 61.575 138.380 62.945 139.160 ;
        RECT 62.955 138.380 66.625 139.190 ;
        RECT 66.645 138.465 67.075 139.250 ;
        RECT 67.555 138.380 69.385 139.190 ;
        RECT 69.395 139.090 70.340 139.290 ;
        RECT 72.155 139.090 73.100 139.290 ;
        RECT 69.395 138.410 72.145 139.090 ;
        RECT 72.155 138.410 74.905 139.090 ;
        RECT 69.395 138.380 70.340 138.410 ;
        RECT 46.080 138.190 46.250 138.380 ;
        RECT 47.915 138.170 48.085 138.360 ;
        RECT 49.760 138.190 49.930 138.380 ;
        RECT 53.435 138.170 53.605 138.360 ;
        RECT 54.410 138.220 54.530 138.330 ;
        RECT 55.735 138.190 55.905 138.380 ;
        RECT 57.115 138.170 57.285 138.360 ;
        RECT 59.600 138.190 59.770 138.380 ;
        RECT 60.335 138.190 60.505 138.380 ;
        RECT 60.980 138.170 61.150 138.360 ;
        RECT 61.715 138.190 61.885 138.380 ;
        RECT 62.175 138.215 62.335 138.325 ;
        RECT 62.635 138.170 62.805 138.360 ;
        RECT 64.070 138.220 64.190 138.330 ;
        RECT 64.475 138.170 64.645 138.360 ;
        RECT 65.855 138.170 66.025 138.360 ;
        RECT 66.315 138.190 66.485 138.380 ;
        RECT 67.290 138.220 67.410 138.330 ;
        RECT 69.075 138.190 69.245 138.380 ;
        RECT 69.995 138.170 70.165 138.360 ;
        RECT 70.455 138.190 70.625 138.360 ;
        RECT 71.830 138.190 72.000 138.410 ;
        RECT 72.155 138.380 73.100 138.410 ;
        RECT 74.590 138.360 74.760 138.410 ;
        RECT 75.375 138.380 80.885 139.190 ;
        RECT 81.265 139.180 82.185 139.290 ;
        RECT 81.265 139.060 83.600 139.180 ;
        RECT 88.265 139.060 89.185 139.280 ;
        RECT 81.265 138.380 90.545 139.060 ;
        RECT 90.555 138.380 92.385 139.190 ;
        RECT 92.405 138.465 92.835 139.250 ;
        RECT 92.855 138.380 95.605 139.190 ;
        RECT 95.625 138.380 96.975 139.290 ;
        RECT 97.915 138.380 99.285 139.160 ;
        RECT 100.215 138.380 103.885 139.190 ;
        RECT 103.895 138.380 109.405 139.190 ;
        RECT 109.425 138.380 110.775 139.290 ;
        RECT 110.795 138.380 112.165 139.160 ;
        RECT 112.175 138.380 113.545 139.190 ;
        RECT 113.555 138.380 117.225 139.190 ;
        RECT 117.235 138.380 118.605 139.190 ;
        RECT 74.590 138.190 74.765 138.360 ;
        RECT 75.110 138.220 75.230 138.330 ;
        RECT 75.515 138.215 75.675 138.325 ;
        RECT 70.475 138.170 70.625 138.190 ;
        RECT 74.595 138.170 74.745 138.190 ;
        RECT 79.195 138.170 79.365 138.360 ;
        RECT 80.170 138.220 80.290 138.330 ;
        RECT 80.575 138.190 80.745 138.380 ;
        RECT 82.875 138.170 83.045 138.360 ;
        RECT 84.255 138.170 84.425 138.360 ;
        RECT 85.175 138.215 85.335 138.325 ;
        RECT 86.555 138.170 86.725 138.360 ;
        RECT 90.235 138.170 90.405 138.380 ;
        RECT 92.075 138.190 92.245 138.380 ;
        RECT 94.100 138.170 94.270 138.360 ;
        RECT 95.295 138.190 95.465 138.380 ;
        RECT 96.675 138.170 96.845 138.380 ;
        RECT 97.595 138.225 97.755 138.335 ;
        RECT 98.055 138.190 98.225 138.380 ;
        RECT 98.975 138.190 99.145 138.360 ;
        RECT 99.895 138.225 100.055 138.335 ;
        RECT 98.975 138.170 99.125 138.190 ;
        RECT 101.735 138.170 101.905 138.360 ;
        RECT 103.575 138.190 103.745 138.380 ;
        RECT 104.035 138.190 104.205 138.360 ;
        RECT 104.955 138.215 105.115 138.325 ;
        RECT 105.930 138.220 106.050 138.330 ;
        RECT 109.095 138.190 109.265 138.380 ;
        RECT 109.555 138.190 109.725 138.380 ;
        RECT 110.935 138.190 111.105 138.380 ;
        RECT 113.235 138.190 113.405 138.380 ;
        RECT 104.035 138.170 104.185 138.190 ;
        RECT 115.535 138.170 115.705 138.360 ;
        RECT 116.915 138.170 117.085 138.380 ;
        RECT 118.295 138.170 118.465 138.380 ;
        RECT 36.895 137.350 38.825 138.170 ;
        RECT 39.035 137.360 42.705 138.170 ;
        RECT 42.715 137.360 48.225 138.170 ;
        RECT 48.235 137.360 53.745 138.170 ;
        RECT 34.635 137.260 35.585 137.350 ;
        RECT 37.875 137.260 38.825 137.350 ;
        RECT 53.765 137.300 54.195 138.085 ;
        RECT 54.675 137.360 57.425 138.170 ;
        RECT 57.665 137.490 61.565 138.170 ;
        RECT 60.635 137.260 61.565 137.490 ;
        RECT 62.495 137.390 63.865 138.170 ;
        RECT 64.335 137.390 65.705 138.170 ;
        RECT 65.715 137.490 67.545 138.170 ;
        RECT 67.555 137.360 70.305 138.170 ;
        RECT 70.475 137.350 72.405 138.170 ;
        RECT 71.455 137.260 72.405 137.350 ;
        RECT 72.815 137.350 74.745 138.170 ;
        RECT 75.835 137.360 79.505 138.170 ;
        RECT 72.815 137.260 73.765 137.350 ;
        RECT 79.525 137.300 79.955 138.085 ;
        RECT 80.435 137.360 83.185 138.170 ;
        RECT 83.205 137.260 84.555 138.170 ;
        RECT 85.505 137.260 86.855 138.170 ;
        RECT 86.875 137.360 90.545 138.170 ;
        RECT 90.785 137.490 94.685 138.170 ;
        RECT 93.755 137.260 94.685 137.490 ;
        RECT 95.615 137.390 96.985 138.170 ;
        RECT 97.195 137.350 99.125 138.170 ;
        RECT 99.295 137.360 102.045 138.170 ;
        RECT 102.255 137.350 104.185 138.170 ;
        RECT 97.195 137.260 98.145 137.350 ;
        RECT 102.255 137.260 103.205 137.350 ;
        RECT 105.285 137.300 105.715 138.085 ;
        RECT 106.565 137.490 115.845 138.170 ;
        RECT 106.565 137.370 108.900 137.490 ;
        RECT 106.565 137.260 107.485 137.370 ;
        RECT 113.565 137.270 114.485 137.490 ;
        RECT 115.855 137.360 117.225 138.170 ;
        RECT 117.235 137.360 118.605 138.170 ;
      LAYER nwell ;
        RECT 11.240 134.140 118.800 136.970 ;
      LAYER pwell ;
        RECT 11.435 132.940 12.805 133.750 ;
        RECT 13.745 132.940 15.095 133.850 ;
        RECT 15.125 133.025 15.555 133.810 ;
        RECT 15.585 132.940 16.935 133.850 ;
        RECT 18.705 133.740 19.625 133.850 ;
        RECT 16.955 132.940 18.325 133.720 ;
        RECT 18.705 133.620 21.040 133.740 ;
        RECT 25.705 133.620 26.625 133.840 ;
        RECT 27.995 133.620 28.925 133.850 ;
        RECT 35.795 133.620 36.725 133.850 ;
        RECT 38.775 133.760 39.725 133.850 ;
        RECT 18.705 132.940 27.985 133.620 ;
        RECT 27.995 132.940 31.895 133.620 ;
        RECT 32.825 132.940 36.725 133.620 ;
        RECT 36.735 132.940 38.565 133.750 ;
        RECT 38.775 132.940 40.705 133.760 ;
        RECT 40.885 133.025 41.315 133.810 ;
        RECT 42.475 133.760 43.425 133.850 ;
        RECT 44.775 133.760 45.725 133.850 ;
        RECT 11.575 132.730 11.745 132.940 ;
        RECT 13.415 132.785 13.575 132.895 ;
        RECT 13.875 132.730 14.045 132.920 ;
        RECT 14.795 132.750 14.965 132.940 ;
        RECT 15.715 132.750 15.885 132.940 ;
        RECT 17.095 132.750 17.265 132.940 ;
        RECT 17.740 132.730 17.910 132.920 ;
        RECT 18.750 132.730 18.920 132.920 ;
        RECT 22.670 132.780 22.790 132.890 ;
        RECT 26.295 132.730 26.465 132.920 ;
        RECT 26.755 132.730 26.925 132.920 ;
        RECT 27.675 132.750 27.845 132.940 ;
        RECT 28.410 132.750 28.580 132.940 ;
        RECT 32.330 132.780 32.450 132.890 ;
        RECT 36.140 132.750 36.310 132.940 ;
        RECT 37.795 132.730 37.965 132.920 ;
        RECT 38.255 132.750 38.425 132.940 ;
        RECT 40.555 132.920 40.705 132.940 ;
        RECT 41.495 132.940 43.425 133.760 ;
        RECT 43.795 132.940 45.725 133.760 ;
        RECT 46.135 133.760 47.085 133.850 ;
        RECT 46.135 132.940 48.065 133.760 ;
        RECT 48.235 132.940 50.065 133.750 ;
        RECT 50.075 132.940 55.585 133.750 ;
        RECT 55.605 132.940 56.955 133.850 ;
        RECT 57.345 133.740 58.265 133.850 ;
        RECT 57.345 133.620 59.680 133.740 ;
        RECT 64.345 133.620 65.265 133.840 ;
        RECT 57.345 132.940 66.625 133.620 ;
        RECT 66.645 133.025 67.075 133.810 ;
        RECT 70.975 133.760 71.925 133.850 ;
        RECT 73.275 133.760 74.225 133.850 ;
        RECT 67.095 132.940 68.925 133.620 ;
        RECT 68.935 132.940 70.765 133.750 ;
        RECT 70.975 132.940 72.905 133.760 ;
        RECT 73.275 132.940 75.205 133.760 ;
        RECT 78.575 133.620 79.505 133.850 ;
        RECT 75.605 132.940 79.505 133.620 ;
        RECT 79.885 133.740 80.805 133.850 ;
        RECT 79.885 133.620 82.220 133.740 ;
        RECT 86.885 133.620 87.805 133.840 ;
        RECT 79.885 132.940 89.165 133.620 ;
        RECT 89.175 132.940 91.005 133.750 ;
        RECT 91.025 132.940 92.375 133.850 ;
        RECT 92.405 133.025 92.835 133.810 ;
        RECT 94.215 133.620 95.135 133.840 ;
        RECT 101.215 133.740 102.135 133.850 ;
        RECT 99.800 133.620 102.135 133.740 ;
        RECT 92.855 132.940 102.135 133.620 ;
        RECT 102.515 132.940 104.345 133.750 ;
        RECT 107.555 133.620 108.485 133.850 ;
        RECT 111.695 133.620 112.625 133.850 ;
        RECT 104.585 132.940 108.485 133.620 ;
        RECT 108.725 132.940 112.625 133.620 ;
        RECT 113.555 132.940 117.225 133.750 ;
        RECT 117.235 132.940 118.605 133.750 ;
        RECT 41.495 132.920 41.645 132.940 ;
        RECT 43.795 132.920 43.945 132.940 ;
        RECT 39.175 132.730 39.345 132.920 ;
        RECT 39.690 132.780 39.810 132.890 ;
        RECT 40.555 132.750 40.725 132.920 ;
        RECT 41.475 132.750 41.645 132.920 ;
        RECT 42.395 132.730 42.565 132.920 ;
        RECT 43.775 132.750 43.945 132.920 ;
        RECT 47.915 132.920 48.065 132.940 ;
        RECT 47.915 132.730 48.085 132.920 ;
        RECT 49.755 132.750 49.925 132.940 ;
        RECT 50.215 132.750 50.385 132.920 ;
        RECT 50.730 132.780 50.850 132.890 ;
        RECT 50.215 132.730 50.365 132.750 ;
        RECT 53.435 132.730 53.605 132.920 ;
        RECT 54.410 132.780 54.530 132.890 ;
        RECT 55.275 132.750 55.445 132.940 ;
        RECT 56.195 132.730 56.365 132.920 ;
        RECT 56.655 132.750 56.825 132.940 ;
        RECT 58.955 132.730 59.125 132.920 ;
        RECT 62.820 132.730 62.990 132.920 ;
        RECT 64.015 132.775 64.175 132.885 ;
        RECT 64.475 132.730 64.645 132.920 ;
        RECT 65.855 132.750 66.025 132.920 ;
        RECT 66.315 132.750 66.485 132.940 ;
        RECT 67.235 132.750 67.405 132.940 ;
        RECT 68.210 132.780 68.330 132.890 ;
        RECT 65.875 132.730 66.025 132.750 ;
        RECT 68.615 132.730 68.785 132.920 ;
        RECT 70.455 132.750 70.625 132.940 ;
        RECT 72.755 132.920 72.905 132.940 ;
        RECT 75.055 132.920 75.205 132.940 ;
        RECT 71.430 132.780 71.550 132.890 ;
        RECT 72.755 132.750 72.925 132.920 ;
        RECT 73.215 132.730 73.385 132.920 ;
        RECT 75.055 132.750 75.225 132.920 ;
        RECT 77.080 132.730 77.250 132.920 ;
        RECT 78.920 132.750 79.090 132.940 ;
        RECT 79.195 132.730 79.365 132.920 ;
        RECT 81.035 132.730 81.205 132.920 ;
        RECT 83.795 132.730 83.965 132.920 ;
        RECT 84.255 132.730 84.425 132.920 ;
        RECT 88.855 132.750 89.025 132.940 ;
        RECT 90.695 132.730 90.865 132.940 ;
        RECT 91.155 132.750 91.325 132.940 ;
        RECT 92.995 132.750 93.165 132.940 ;
        RECT 92.995 132.730 93.145 132.750 ;
        RECT 96.860 132.730 97.030 132.920 ;
        RECT 97.650 132.780 97.770 132.890 ;
        RECT 99.895 132.750 100.065 132.920 ;
        RECT 102.195 132.750 102.365 132.920 ;
        RECT 104.035 132.750 104.205 132.940 ;
        RECT 104.495 132.750 104.665 132.920 ;
        RECT 105.010 132.780 105.130 132.890 ;
        RECT 106.335 132.775 106.495 132.885 ;
        RECT 107.900 132.750 108.070 132.940 ;
        RECT 112.040 132.750 112.210 132.940 ;
        RECT 113.235 132.785 113.395 132.895 ;
        RECT 99.895 132.730 100.045 132.750 ;
        RECT 102.195 132.730 102.345 132.750 ;
        RECT 104.495 132.730 104.645 132.750 ;
        RECT 115.995 132.730 116.165 132.920 ;
        RECT 116.915 132.750 117.085 132.940 ;
        RECT 118.295 132.730 118.465 132.940 ;
        RECT 11.435 131.920 12.805 132.730 ;
        RECT 12.815 131.920 14.185 132.730 ;
        RECT 14.425 132.050 18.325 132.730 ;
        RECT 17.395 131.820 18.325 132.050 ;
        RECT 18.335 132.050 22.235 132.730 ;
        RECT 18.335 131.820 19.265 132.050 ;
        RECT 22.935 131.920 26.605 132.730 ;
        RECT 26.625 131.820 27.975 132.730 ;
        RECT 28.005 131.860 28.435 132.645 ;
        RECT 28.825 132.050 38.105 132.730 ;
        RECT 28.825 131.930 31.160 132.050 ;
        RECT 28.825 131.820 29.745 131.930 ;
        RECT 35.825 131.830 36.745 132.050 ;
        RECT 38.115 131.950 39.485 132.730 ;
        RECT 39.955 131.920 42.705 132.730 ;
        RECT 42.715 131.920 48.225 132.730 ;
        RECT 48.435 131.910 50.365 132.730 ;
        RECT 50.995 131.920 53.745 132.730 ;
        RECT 48.435 131.820 49.385 131.910 ;
        RECT 53.765 131.860 54.195 132.645 ;
        RECT 54.675 131.920 56.505 132.730 ;
        RECT 56.525 132.050 59.265 132.730 ;
        RECT 59.505 132.050 63.405 132.730 ;
        RECT 62.475 131.820 63.405 132.050 ;
        RECT 64.335 131.950 65.705 132.730 ;
        RECT 65.875 131.910 67.805 132.730 ;
        RECT 68.475 132.050 71.215 132.730 ;
        RECT 71.695 131.920 73.525 132.730 ;
        RECT 73.765 132.050 77.665 132.730 ;
        RECT 66.855 131.820 67.805 131.910 ;
        RECT 76.735 131.820 77.665 132.050 ;
        RECT 77.675 131.920 79.505 132.730 ;
        RECT 79.525 131.860 79.955 132.645 ;
        RECT 79.975 131.950 81.345 132.730 ;
        RECT 81.355 131.920 84.105 132.730 ;
        RECT 84.115 131.950 85.485 132.730 ;
        RECT 85.495 131.920 91.005 132.730 ;
        RECT 91.215 131.910 93.145 132.730 ;
        RECT 93.545 132.050 97.445 132.730 ;
        RECT 91.215 131.820 92.165 131.910 ;
        RECT 96.515 131.820 97.445 132.050 ;
        RECT 98.115 131.910 100.045 132.730 ;
        RECT 100.415 131.910 102.345 132.730 ;
        RECT 102.715 131.910 104.645 132.730 ;
        RECT 98.115 131.820 99.065 131.910 ;
        RECT 100.415 131.820 101.365 131.910 ;
        RECT 102.715 131.820 103.665 131.910 ;
        RECT 105.285 131.860 105.715 132.645 ;
        RECT 107.025 132.050 116.305 132.730 ;
        RECT 107.025 131.930 109.360 132.050 ;
        RECT 107.025 131.820 107.945 131.930 ;
        RECT 114.025 131.830 114.945 132.050 ;
        RECT 117.235 131.920 118.605 132.730 ;
      LAYER nwell ;
        RECT 11.240 128.700 118.800 131.530 ;
      LAYER pwell ;
        RECT 11.435 127.500 12.805 128.310 ;
        RECT 13.745 127.500 15.095 128.410 ;
        RECT 15.125 127.585 15.555 128.370 ;
        RECT 16.495 127.500 17.865 128.280 ;
        RECT 17.875 128.180 18.805 128.410 ;
        RECT 35.115 128.320 36.065 128.410 ;
        RECT 17.875 127.500 21.775 128.180 ;
        RECT 22.935 127.500 28.445 128.310 ;
        RECT 28.455 127.500 33.965 128.310 ;
        RECT 34.135 127.500 36.065 128.320 ;
        RECT 39.935 128.180 40.865 128.410 ;
        RECT 36.965 127.500 40.865 128.180 ;
        RECT 40.885 127.585 41.315 128.370 ;
        RECT 42.165 128.300 43.085 128.410 ;
        RECT 42.165 128.180 44.500 128.300 ;
        RECT 49.165 128.180 50.085 128.400 ;
        RECT 42.165 127.500 51.445 128.180 ;
        RECT 51.465 127.500 52.815 128.410 ;
        RECT 57.345 128.300 58.265 128.410 ;
        RECT 53.295 127.500 54.665 128.280 ;
        RECT 57.345 128.180 59.680 128.300 ;
        RECT 64.345 128.180 65.265 128.400 ;
        RECT 55.135 127.500 56.090 128.180 ;
        RECT 57.345 127.500 66.625 128.180 ;
        RECT 66.645 127.585 67.075 128.370 ;
        RECT 67.555 127.500 70.305 128.310 ;
        RECT 70.685 128.300 71.605 128.410 ;
        RECT 70.685 128.180 73.020 128.300 ;
        RECT 77.685 128.180 78.605 128.400 ;
        RECT 70.685 127.500 79.965 128.180 ;
        RECT 80.060 127.500 89.165 128.180 ;
        RECT 89.185 127.500 90.535 128.410 ;
        RECT 90.555 127.500 92.385 128.310 ;
        RECT 92.405 127.585 92.835 128.370 ;
        RECT 93.315 127.500 95.145 128.310 ;
        RECT 95.155 127.500 96.525 128.280 ;
        RECT 108.935 128.180 109.865 128.410 ;
        RECT 96.535 127.500 105.640 128.180 ;
        RECT 105.965 127.500 109.865 128.180 ;
        RECT 109.875 127.500 110.830 128.180 ;
        RECT 111.265 127.500 112.615 128.410 ;
        RECT 112.635 127.500 114.005 128.280 ;
        RECT 114.475 127.500 117.225 128.310 ;
        RECT 117.235 127.500 118.605 128.310 ;
        RECT 11.575 127.290 11.745 127.500 ;
        RECT 13.415 127.335 13.575 127.455 ;
        RECT 14.795 127.310 14.965 127.500 ;
        RECT 16.175 127.345 16.335 127.455 ;
        RECT 16.635 127.310 16.805 127.500 ;
        RECT 18.290 127.310 18.460 127.500 ;
        RECT 22.615 127.345 22.775 127.455 ;
        RECT 23.075 127.290 23.245 127.480 ;
        RECT 23.590 127.340 23.710 127.450 ;
        RECT 23.995 127.290 24.165 127.480 ;
        RECT 27.675 127.290 27.845 127.480 ;
        RECT 28.135 127.310 28.305 127.500 ;
        RECT 32.000 127.290 32.170 127.480 ;
        RECT 33.655 127.290 33.825 127.500 ;
        RECT 34.135 127.480 34.285 127.500 ;
        RECT 34.115 127.310 34.285 127.480 ;
        RECT 36.470 127.340 36.590 127.450 ;
        RECT 40.280 127.310 40.450 127.500 ;
        RECT 41.530 127.340 41.650 127.450 ;
        RECT 43.315 127.290 43.485 127.480 ;
        RECT 43.830 127.340 43.950 127.450 ;
        RECT 51.135 127.310 51.305 127.500 ;
        RECT 52.515 127.310 52.685 127.500 ;
        RECT 53.030 127.340 53.150 127.450 ;
        RECT 53.435 127.290 53.605 127.480 ;
        RECT 54.355 127.310 54.525 127.500 ;
        RECT 54.630 127.290 54.800 127.480 ;
        RECT 54.870 127.340 54.990 127.450 ;
        RECT 56.195 127.310 56.365 127.480 ;
        RECT 56.710 127.340 56.830 127.450 ;
        RECT 58.955 127.335 59.115 127.445 ;
        RECT 62.635 127.290 62.805 127.480 ;
        RECT 64.015 127.290 64.185 127.480 ;
        RECT 64.530 127.340 64.650 127.450 ;
        RECT 66.315 127.290 66.485 127.500 ;
        RECT 67.290 127.340 67.410 127.450 ;
        RECT 69.995 127.310 70.165 127.500 ;
        RECT 71.835 127.290 72.005 127.480 ;
        RECT 72.295 127.290 72.465 127.480 ;
        RECT 73.675 127.290 73.845 127.480 ;
        RECT 75.110 127.340 75.230 127.450 ;
        RECT 78.920 127.290 79.090 127.480 ;
        RECT 79.655 127.310 79.825 127.500 ;
        RECT 81.495 127.290 81.665 127.480 ;
        RECT 81.955 127.290 82.125 127.480 ;
        RECT 86.740 127.290 86.910 127.480 ;
        RECT 88.855 127.310 89.025 127.500 ;
        RECT 89.315 127.310 89.485 127.500 ;
        RECT 92.075 127.310 92.245 127.500 ;
        RECT 93.050 127.340 93.170 127.450 ;
        RECT 94.835 127.310 95.005 127.500 ;
        RECT 95.295 127.310 95.465 127.500 ;
        RECT 96.675 127.290 96.845 127.500 ;
        RECT 97.190 127.340 97.310 127.450 ;
        RECT 98.975 127.290 99.145 127.480 ;
        RECT 99.435 127.290 99.605 127.480 ;
        RECT 101.090 127.290 101.260 127.480 ;
        RECT 105.010 127.340 105.130 127.450 ;
        RECT 109.280 127.310 109.450 127.500 ;
        RECT 110.935 127.310 111.105 127.480 ;
        RECT 112.315 127.310 112.485 127.500 ;
        RECT 112.775 127.310 112.945 127.500 ;
        RECT 114.210 127.340 114.330 127.450 ;
        RECT 115.075 127.290 115.245 127.480 ;
        RECT 116.915 127.290 117.085 127.500 ;
        RECT 118.295 127.290 118.465 127.500 ;
        RECT 11.435 126.480 12.805 127.290 ;
        RECT 14.105 126.610 23.385 127.290 ;
        RECT 14.105 126.490 16.440 126.610 ;
        RECT 14.105 126.380 15.025 126.490 ;
        RECT 21.105 126.390 22.025 126.610 ;
        RECT 23.865 126.380 25.215 127.290 ;
        RECT 25.245 126.610 27.985 127.290 ;
        RECT 28.005 126.420 28.435 127.205 ;
        RECT 28.685 126.610 32.585 127.290 ;
        RECT 31.655 126.380 32.585 126.610 ;
        RECT 32.595 126.480 33.965 127.290 ;
        RECT 34.345 126.610 43.625 127.290 ;
        RECT 44.465 126.610 53.745 127.290 ;
        RECT 34.345 126.490 36.680 126.610 ;
        RECT 34.345 126.380 35.265 126.490 ;
        RECT 41.345 126.390 42.265 126.610 ;
        RECT 44.465 126.490 46.800 126.610 ;
        RECT 44.465 126.380 45.385 126.490 ;
        RECT 51.465 126.390 52.385 126.610 ;
        RECT 53.765 126.420 54.195 127.205 ;
        RECT 54.215 126.610 58.115 127.290 ;
        RECT 54.215 126.380 55.145 126.610 ;
        RECT 59.275 126.480 62.945 127.290 ;
        RECT 62.965 126.380 64.315 127.290 ;
        RECT 64.795 126.480 66.625 127.290 ;
        RECT 66.635 126.480 72.145 127.290 ;
        RECT 72.165 126.380 73.515 127.290 ;
        RECT 73.545 126.380 74.895 127.290 ;
        RECT 75.605 126.610 79.505 127.290 ;
        RECT 78.575 126.380 79.505 126.610 ;
        RECT 79.525 126.420 79.955 127.205 ;
        RECT 79.975 126.480 81.805 127.290 ;
        RECT 81.825 126.380 83.175 127.290 ;
        RECT 83.425 126.610 87.325 127.290 ;
        RECT 86.395 126.380 87.325 126.610 ;
        RECT 87.705 126.610 96.985 127.290 ;
        RECT 87.705 126.490 90.040 126.610 ;
        RECT 87.705 126.380 88.625 126.490 ;
        RECT 94.705 126.390 95.625 126.610 ;
        RECT 97.455 126.480 99.285 127.290 ;
        RECT 99.305 126.380 100.655 127.290 ;
        RECT 100.675 126.610 104.575 127.290 ;
        RECT 100.675 126.380 101.605 126.610 ;
        RECT 105.285 126.420 105.715 127.205 ;
        RECT 106.105 126.610 115.385 127.290 ;
        RECT 106.105 126.490 108.440 126.610 ;
        RECT 106.105 126.380 107.025 126.490 ;
        RECT 113.105 126.390 114.025 126.610 ;
        RECT 115.395 126.480 117.225 127.290 ;
        RECT 117.235 126.480 118.605 127.290 ;
      LAYER nwell ;
        RECT 11.240 123.260 118.800 126.090 ;
      LAYER pwell ;
        RECT 11.435 122.060 12.805 122.870 ;
        RECT 13.745 122.060 15.095 122.970 ;
        RECT 15.125 122.145 15.555 122.930 ;
        RECT 15.945 122.860 16.865 122.970 ;
        RECT 15.945 122.740 18.280 122.860 ;
        RECT 22.945 122.740 23.865 122.960 ;
        RECT 25.605 122.860 26.525 122.970 ;
        RECT 25.605 122.740 27.940 122.860 ;
        RECT 32.605 122.740 33.525 122.960 ;
        RECT 15.945 122.060 25.225 122.740 ;
        RECT 25.605 122.060 34.885 122.740 ;
        RECT 35.355 122.060 37.185 122.870 ;
        RECT 37.205 122.060 38.555 122.970 ;
        RECT 39.035 122.060 40.865 122.870 ;
        RECT 40.885 122.145 41.315 122.930 ;
        RECT 41.335 122.060 42.705 122.840 ;
        RECT 42.725 122.060 44.075 122.970 ;
        RECT 53.665 122.860 54.585 122.970 ;
        RECT 53.665 122.740 56.000 122.860 ;
        RECT 60.665 122.740 61.585 122.960 ;
        RECT 44.180 122.060 53.285 122.740 ;
        RECT 53.665 122.060 62.945 122.740 ;
        RECT 62.955 122.060 66.625 122.870 ;
        RECT 66.645 122.145 67.075 122.930 ;
        RECT 67.555 122.060 70.305 122.870 ;
        RECT 70.325 122.060 71.675 122.970 ;
        RECT 72.525 122.860 73.445 122.970 ;
        RECT 72.525 122.740 74.860 122.860 ;
        RECT 79.525 122.740 80.445 122.960 ;
        RECT 82.185 122.860 83.105 122.970 ;
        RECT 82.185 122.740 84.520 122.860 ;
        RECT 89.185 122.740 90.105 122.960 ;
        RECT 72.525 122.060 81.805 122.740 ;
        RECT 82.185 122.060 91.465 122.740 ;
        RECT 92.405 122.145 92.835 122.930 ;
        RECT 93.315 122.060 95.145 122.870 ;
        RECT 96.905 122.860 97.825 122.970 ;
        RECT 95.155 122.060 96.525 122.840 ;
        RECT 96.905 122.740 99.240 122.860 ;
        RECT 103.905 122.740 104.825 122.960 ;
        RECT 96.905 122.060 106.185 122.740 ;
        RECT 106.195 122.060 108.945 122.870 ;
        RECT 108.965 122.060 110.315 122.970 ;
        RECT 110.795 122.060 112.165 122.840 ;
        RECT 112.175 122.060 113.545 122.870 ;
        RECT 113.555 122.060 117.225 122.870 ;
        RECT 117.235 122.060 118.605 122.870 ;
        RECT 11.575 121.850 11.745 122.060 ;
        RECT 13.415 121.895 13.575 122.015 ;
        RECT 14.795 121.870 14.965 122.060 ;
        RECT 17.095 121.850 17.265 122.040 ;
        RECT 17.555 121.850 17.725 122.040 ;
        RECT 24.915 121.870 25.085 122.060 ;
        RECT 27.675 121.850 27.845 122.040 ;
        RECT 28.650 121.900 28.770 122.010 ;
        RECT 31.355 121.850 31.525 122.040 ;
        RECT 31.815 121.850 31.985 122.040 ;
        RECT 33.250 121.900 33.370 122.010 ;
        RECT 34.575 121.870 34.745 122.060 ;
        RECT 35.090 121.900 35.210 122.010 ;
        RECT 36.875 121.870 37.045 122.060 ;
        RECT 37.335 121.870 37.505 122.060 ;
        RECT 38.715 122.010 38.885 122.040 ;
        RECT 38.715 121.900 38.890 122.010 ;
        RECT 38.715 121.850 38.885 121.900 ;
        RECT 40.555 121.870 40.725 122.060 ;
        RECT 41.475 121.870 41.645 122.060 ;
        RECT 42.855 121.870 43.025 122.060 ;
        RECT 44.235 121.850 44.405 122.040 ;
        RECT 48.100 121.850 48.270 122.040 ;
        RECT 48.890 121.900 49.010 122.010 ;
        RECT 52.700 121.850 52.870 122.040 ;
        RECT 52.975 121.870 53.145 122.060 ;
        RECT 53.490 121.900 53.610 122.010 ;
        RECT 54.355 121.850 54.525 122.040 ;
        RECT 55.735 121.850 55.905 122.040 ;
        RECT 59.410 121.850 59.580 122.040 ;
        RECT 60.795 121.850 60.965 122.040 ;
        RECT 62.635 121.870 62.805 122.060 ;
        RECT 66.315 121.850 66.485 122.060 ;
        RECT 67.290 121.900 67.410 122.010 ;
        RECT 69.995 121.870 70.165 122.060 ;
        RECT 71.375 121.870 71.545 122.060 ;
        RECT 71.835 122.010 72.005 122.040 ;
        RECT 71.835 121.900 72.010 122.010 ;
        RECT 71.835 121.850 72.005 121.900 ;
        RECT 73.215 121.850 73.385 122.040 ;
        RECT 74.135 121.895 74.295 122.005 ;
        RECT 77.815 121.850 77.985 122.040 ;
        RECT 78.275 121.850 78.445 122.040 ;
        RECT 81.495 121.870 81.665 122.060 ;
        RECT 82.415 121.850 82.585 122.040 ;
        RECT 87.935 121.850 88.105 122.040 ;
        RECT 88.395 121.850 88.565 122.040 ;
        RECT 90.235 121.895 90.395 122.005 ;
        RECT 91.155 121.870 91.325 122.060 ;
        RECT 92.075 121.905 92.235 122.015 ;
        RECT 93.050 121.900 93.170 122.010 ;
        RECT 93.915 121.850 94.085 122.040 ;
        RECT 94.835 121.870 95.005 122.060 ;
        RECT 96.215 121.870 96.385 122.060 ;
        RECT 99.435 121.850 99.605 122.040 ;
        RECT 104.955 121.850 105.125 122.040 ;
        RECT 105.875 121.870 106.045 122.060 ;
        RECT 106.795 121.850 106.965 122.040 ;
        RECT 108.635 121.870 108.805 122.060 ;
        RECT 109.095 121.870 109.265 122.060 ;
        RECT 110.475 122.010 110.645 122.040 ;
        RECT 110.475 121.900 110.650 122.010 ;
        RECT 110.475 121.850 110.645 121.900 ;
        RECT 110.935 121.850 111.105 122.060 ;
        RECT 112.775 121.895 112.935 122.005 ;
        RECT 113.235 121.850 113.405 122.060 ;
        RECT 116.915 122.040 117.085 122.060 ;
        RECT 115.535 121.850 115.705 122.040 ;
        RECT 116.905 121.870 117.085 122.040 ;
        RECT 116.905 121.850 117.075 121.870 ;
        RECT 118.295 121.850 118.465 122.060 ;
        RECT 11.435 121.040 12.805 121.850 ;
        RECT 13.735 121.040 17.405 121.850 ;
        RECT 17.415 121.070 18.785 121.850 ;
        RECT 18.880 121.170 27.985 121.850 ;
        RECT 28.005 120.980 28.435 121.765 ;
        RECT 28.915 121.040 31.665 121.850 ;
        RECT 31.675 121.070 33.045 121.850 ;
        RECT 33.515 121.040 39.025 121.850 ;
        RECT 39.035 121.040 44.545 121.850 ;
        RECT 44.785 121.170 48.685 121.850 ;
        RECT 49.385 121.170 53.285 121.850 ;
        RECT 47.755 120.940 48.685 121.170 ;
        RECT 52.355 120.940 53.285 121.170 ;
        RECT 53.765 120.980 54.195 121.765 ;
        RECT 54.225 120.940 55.575 121.850 ;
        RECT 55.595 121.070 56.965 121.850 ;
        RECT 57.115 120.940 59.725 121.850 ;
        RECT 59.735 121.040 61.105 121.850 ;
        RECT 61.115 121.040 66.625 121.850 ;
        RECT 66.635 121.040 72.145 121.850 ;
        RECT 72.165 120.940 73.515 121.850 ;
        RECT 74.455 121.040 78.125 121.850 ;
        RECT 78.135 121.070 79.505 121.850 ;
        RECT 79.525 120.980 79.955 121.765 ;
        RECT 79.975 121.040 82.725 121.850 ;
        RECT 82.735 121.040 88.245 121.850 ;
        RECT 88.255 121.070 89.625 121.850 ;
        RECT 90.555 121.040 94.225 121.850 ;
        RECT 94.235 121.040 99.745 121.850 ;
        RECT 99.755 121.040 105.265 121.850 ;
        RECT 105.285 120.980 105.715 121.765 ;
        RECT 105.735 121.040 107.105 121.850 ;
        RECT 107.115 121.040 110.785 121.850 ;
        RECT 110.805 120.940 112.155 121.850 ;
        RECT 113.095 121.070 114.465 121.850 ;
        RECT 114.475 121.040 115.845 121.850 ;
        RECT 115.855 121.070 117.225 121.850 ;
        RECT 117.235 121.040 118.605 121.850 ;
      LAYER nwell ;
        RECT 11.240 117.820 118.800 120.650 ;
      LAYER pwell ;
        RECT 11.435 116.620 12.805 117.430 ;
        RECT 13.275 116.620 15.105 117.430 ;
        RECT 15.125 116.705 15.555 117.490 ;
        RECT 15.575 116.620 18.325 117.430 ;
        RECT 18.335 116.620 23.845 117.430 ;
        RECT 23.855 116.620 25.225 117.400 ;
        RECT 25.235 116.620 26.605 117.430 ;
        RECT 26.615 116.620 30.285 117.430 ;
        RECT 30.495 117.300 32.705 117.530 ;
        RECT 35.425 117.300 36.355 117.520 ;
        RECT 30.495 116.620 40.865 117.300 ;
        RECT 40.885 116.705 41.315 117.490 ;
        RECT 41.335 116.620 42.705 117.400 ;
        RECT 42.715 116.620 44.085 117.400 ;
        RECT 44.095 116.620 46.845 117.430 ;
        RECT 46.855 116.620 48.225 117.400 ;
        RECT 48.235 116.620 49.605 117.400 ;
        RECT 50.075 116.620 51.905 117.430 ;
        RECT 51.915 116.620 57.425 117.430 ;
        RECT 57.445 116.620 58.795 117.530 ;
        RECT 58.955 116.620 61.565 117.530 ;
        RECT 61.575 116.620 63.405 117.430 ;
        RECT 63.415 116.620 64.785 117.400 ;
        RECT 64.795 116.620 66.625 117.430 ;
        RECT 66.645 116.705 67.075 117.490 ;
        RECT 67.095 116.620 68.465 117.430 ;
        RECT 68.485 116.620 69.835 117.530 ;
        RECT 69.855 116.620 72.465 117.530 ;
        RECT 72.615 116.620 73.985 117.400 ;
        RECT 73.995 116.620 75.365 117.400 ;
        RECT 75.835 116.620 77.665 117.430 ;
        RECT 77.675 116.620 79.045 117.400 ;
        RECT 79.515 116.620 85.025 117.430 ;
        RECT 85.035 116.620 86.405 117.400 ;
        RECT 86.875 116.620 92.385 117.430 ;
        RECT 92.405 116.705 92.835 117.490 ;
        RECT 92.855 116.620 94.225 117.430 ;
        RECT 94.235 116.620 97.905 117.430 ;
        RECT 97.915 116.620 99.285 117.400 ;
        RECT 99.765 116.620 101.115 117.530 ;
        RECT 101.135 116.620 102.505 117.400 ;
        RECT 102.515 116.620 103.885 117.430 ;
        RECT 103.905 116.620 105.255 117.530 ;
        RECT 105.275 116.620 106.645 117.400 ;
        RECT 111.165 117.300 112.095 117.520 ;
        RECT 114.815 117.300 117.025 117.530 ;
        RECT 106.655 116.620 117.025 117.300 ;
        RECT 117.235 116.620 118.605 117.430 ;
        RECT 11.575 116.410 11.745 116.620 ;
        RECT 13.010 116.460 13.130 116.570 ;
        RECT 14.795 116.430 14.965 116.620 ;
        RECT 15.715 116.410 15.885 116.600 ;
        RECT 18.015 116.430 18.185 116.620 ;
        RECT 23.535 116.430 23.705 116.620 ;
        RECT 24.915 116.430 25.085 116.620 ;
        RECT 26.295 116.410 26.465 116.620 ;
        RECT 27.675 116.410 27.845 116.600 ;
        RECT 28.595 116.410 28.765 116.600 ;
        RECT 29.975 116.410 30.145 116.620 ;
        RECT 32.275 116.410 32.445 116.600 ;
        RECT 40.555 116.430 40.725 116.620 ;
        RECT 42.395 116.430 42.565 116.620 ;
        RECT 42.855 116.410 43.025 116.600 ;
        RECT 43.775 116.430 43.945 116.620 ;
        RECT 46.535 116.430 46.705 116.620 ;
        RECT 46.995 116.430 47.165 116.620 ;
        RECT 48.375 116.430 48.545 116.620 ;
        RECT 49.810 116.460 49.930 116.570 ;
        RECT 51.595 116.430 51.765 116.620 ;
        RECT 53.435 116.410 53.605 116.600 ;
        RECT 55.275 116.410 55.445 116.600 ;
        RECT 55.790 116.460 55.910 116.570 ;
        RECT 56.195 116.410 56.365 116.600 ;
        RECT 57.115 116.430 57.285 116.620 ;
        RECT 57.575 116.430 57.745 116.620 ;
        RECT 61.250 116.430 61.420 116.620 ;
        RECT 63.095 116.430 63.265 116.620 ;
        RECT 63.555 116.430 63.725 116.620 ;
        RECT 66.315 116.430 66.485 116.620 ;
        RECT 67.695 116.410 67.865 116.600 ;
        RECT 68.155 116.430 68.325 116.620 ;
        RECT 69.535 116.430 69.705 116.620 ;
        RECT 70.000 116.430 70.170 116.620 ;
        RECT 72.755 116.430 72.925 116.620 ;
        RECT 74.135 116.430 74.305 116.620 ;
        RECT 75.570 116.460 75.690 116.570 ;
        RECT 77.355 116.430 77.525 116.620 ;
        RECT 77.815 116.430 77.985 116.620 ;
        RECT 78.275 116.410 78.445 116.600 ;
        RECT 79.250 116.565 79.370 116.570 ;
        RECT 79.195 116.460 79.370 116.565 ;
        RECT 79.195 116.455 79.355 116.460 ;
        RECT 84.715 116.430 84.885 116.620 ;
        RECT 85.175 116.430 85.345 116.620 ;
        RECT 86.610 116.460 86.730 116.570 ;
        RECT 90.235 116.410 90.405 116.600 ;
        RECT 91.615 116.410 91.785 116.600 ;
        RECT 92.075 116.430 92.245 116.620 ;
        RECT 92.995 116.410 93.165 116.600 ;
        RECT 93.455 116.410 93.625 116.600 ;
        RECT 93.915 116.430 94.085 116.620 ;
        RECT 97.595 116.430 97.765 116.620 ;
        RECT 98.055 116.430 98.225 116.620 ;
        RECT 99.490 116.460 99.610 116.570 ;
        RECT 100.815 116.430 100.985 116.620 ;
        RECT 101.275 116.430 101.445 116.620 ;
        RECT 103.575 116.430 103.745 116.620 ;
        RECT 104.035 116.430 104.205 116.620 ;
        RECT 104.955 116.410 105.125 116.600 ;
        RECT 105.415 116.430 105.585 116.620 ;
        RECT 106.335 116.455 106.495 116.565 ;
        RECT 106.795 116.430 106.965 116.620 ;
        RECT 116.915 116.410 117.085 116.600 ;
        RECT 118.295 116.410 118.465 116.620 ;
        RECT 11.435 115.600 12.805 116.410 ;
        RECT 13.275 115.600 16.025 116.410 ;
        RECT 16.235 115.730 26.605 116.410 ;
        RECT 16.235 115.500 18.445 115.730 ;
        RECT 21.165 115.510 22.095 115.730 ;
        RECT 26.615 115.630 27.985 116.410 ;
        RECT 28.005 115.540 28.435 116.325 ;
        RECT 28.465 115.500 29.815 116.410 ;
        RECT 29.845 115.500 31.195 116.410 ;
        RECT 31.215 115.630 32.585 116.410 ;
        RECT 32.795 115.730 43.165 116.410 ;
        RECT 43.375 115.730 53.745 116.410 ;
        RECT 32.795 115.500 35.005 115.730 ;
        RECT 37.725 115.510 38.655 115.730 ;
        RECT 43.375 115.500 45.585 115.730 ;
        RECT 48.305 115.510 49.235 115.730 ;
        RECT 53.765 115.540 54.195 116.325 ;
        RECT 54.215 115.630 55.585 116.410 ;
        RECT 56.055 115.630 57.425 116.410 ;
        RECT 57.635 115.730 68.005 116.410 ;
        RECT 68.215 115.730 78.585 116.410 ;
        RECT 57.635 115.500 59.845 115.730 ;
        RECT 62.565 115.510 63.495 115.730 ;
        RECT 68.215 115.500 70.425 115.730 ;
        RECT 73.145 115.510 74.075 115.730 ;
        RECT 79.525 115.540 79.955 116.325 ;
        RECT 80.175 115.730 90.545 116.410 ;
        RECT 80.175 115.500 82.385 115.730 ;
        RECT 85.105 115.510 86.035 115.730 ;
        RECT 90.555 115.600 91.925 116.410 ;
        RECT 91.935 115.630 93.305 116.410 ;
        RECT 93.325 115.500 94.675 116.410 ;
        RECT 94.895 115.730 105.265 116.410 ;
        RECT 94.895 115.500 97.105 115.730 ;
        RECT 99.825 115.510 100.755 115.730 ;
        RECT 105.285 115.540 105.715 116.325 ;
        RECT 106.855 115.730 117.225 116.410 ;
        RECT 106.855 115.500 109.065 115.730 ;
        RECT 111.785 115.510 112.715 115.730 ;
        RECT 117.235 115.600 118.605 116.410 ;
      LAYER nwell ;
        RECT 11.240 112.380 118.800 115.210 ;
      LAYER pwell ;
        RECT 11.435 111.180 12.805 111.990 ;
        RECT 13.745 111.180 15.095 112.090 ;
        RECT 15.125 111.265 15.555 112.050 ;
        RECT 15.585 111.180 16.935 112.090 ;
        RECT 17.155 111.860 19.365 112.090 ;
        RECT 22.085 111.860 23.015 112.080 ;
        RECT 27.735 111.860 29.945 112.090 ;
        RECT 32.665 111.860 33.595 112.080 ;
        RECT 17.155 111.180 27.525 111.860 ;
        RECT 27.735 111.180 38.105 111.860 ;
        RECT 38.125 111.180 39.475 112.090 ;
        RECT 39.495 111.180 40.865 111.960 ;
        RECT 40.885 111.265 41.315 112.050 ;
        RECT 41.795 111.180 43.625 111.990 ;
        RECT 43.835 111.860 46.045 112.090 ;
        RECT 48.765 111.860 49.695 112.080 ;
        RECT 54.415 111.860 56.625 112.090 ;
        RECT 59.345 111.860 60.275 112.080 ;
        RECT 43.835 111.180 54.205 111.860 ;
        RECT 54.415 111.180 64.785 111.860 ;
        RECT 64.795 111.180 66.625 111.990 ;
        RECT 66.645 111.265 67.075 112.050 ;
        RECT 67.755 111.860 69.965 112.090 ;
        RECT 72.685 111.860 73.615 112.080 ;
        RECT 78.335 111.860 80.545 112.090 ;
        RECT 83.265 111.860 84.195 112.080 ;
        RECT 67.755 111.180 78.125 111.860 ;
        RECT 78.335 111.180 88.705 111.860 ;
        RECT 88.725 111.180 90.075 112.090 ;
        RECT 90.105 111.180 91.455 112.090 ;
        RECT 92.405 111.265 92.835 112.050 ;
        RECT 93.055 111.860 95.265 112.090 ;
        RECT 97.985 111.860 98.915 112.080 ;
        RECT 103.635 111.860 105.845 112.090 ;
        RECT 108.565 111.860 109.495 112.080 ;
        RECT 93.055 111.180 103.425 111.860 ;
        RECT 103.635 111.180 114.005 111.860 ;
        RECT 114.015 111.180 115.385 111.960 ;
        RECT 115.395 111.180 117.225 111.990 ;
        RECT 117.235 111.180 118.605 111.990 ;
        RECT 11.575 110.970 11.745 111.180 ;
        RECT 13.010 111.020 13.130 111.130 ;
        RECT 13.415 111.025 13.575 111.135 ;
        RECT 14.795 110.970 14.965 111.180 ;
        RECT 15.715 110.990 15.885 111.180 ;
        RECT 25.835 110.970 26.005 111.160 ;
        RECT 27.215 110.970 27.385 111.180 ;
        RECT 27.730 111.020 27.850 111.130 ;
        RECT 29.515 110.970 29.685 111.160 ;
        RECT 35.035 110.970 35.205 111.160 ;
        RECT 37.795 110.990 37.965 111.180 ;
        RECT 39.175 110.990 39.345 111.180 ;
        RECT 40.555 110.970 40.725 111.180 ;
        RECT 41.530 111.020 41.650 111.130 ;
        RECT 43.315 110.990 43.485 111.180 ;
        RECT 46.995 110.970 47.165 111.160 ;
        RECT 48.375 110.970 48.545 111.160 ;
        RECT 51.135 110.970 51.305 111.160 ;
        RECT 52.515 110.970 52.685 111.160 ;
        RECT 53.435 111.015 53.595 111.125 ;
        RECT 53.895 110.990 54.065 111.180 ;
        RECT 54.410 111.020 54.530 111.130 ;
        RECT 58.035 110.970 58.205 111.160 ;
        RECT 59.415 110.970 59.585 111.160 ;
        RECT 60.795 110.970 60.965 111.160 ;
        RECT 64.475 110.990 64.645 111.180 ;
        RECT 66.315 110.970 66.485 111.180 ;
        RECT 67.290 111.020 67.410 111.130 ;
        RECT 72.295 110.970 72.465 111.160 ;
        RECT 77.815 110.970 77.985 111.180 ;
        RECT 78.275 110.970 78.445 111.160 ;
        RECT 81.495 110.970 81.665 111.160 ;
        RECT 88.395 110.990 88.565 111.180 ;
        RECT 89.775 110.990 89.945 111.180 ;
        RECT 91.155 110.990 91.325 111.180 ;
        RECT 92.075 110.970 92.245 111.160 ;
        RECT 93.915 110.970 94.085 111.160 ;
        RECT 99.435 110.970 99.605 111.160 ;
        RECT 103.115 110.990 103.285 111.180 ;
        RECT 104.955 110.970 105.125 111.160 ;
        RECT 106.335 111.015 106.495 111.125 ;
        RECT 110.015 110.970 110.185 111.160 ;
        RECT 110.475 110.970 110.645 111.160 ;
        RECT 113.695 110.990 113.865 111.180 ;
        RECT 114.155 110.990 114.325 111.180 ;
        RECT 116.915 110.970 117.085 111.180 ;
        RECT 118.295 110.970 118.465 111.180 ;
        RECT 11.435 110.160 12.805 110.970 ;
        RECT 13.275 110.160 15.105 110.970 ;
        RECT 15.125 110.100 15.555 110.885 ;
        RECT 15.775 110.290 26.145 110.970 ;
        RECT 15.775 110.060 17.985 110.290 ;
        RECT 20.705 110.070 21.635 110.290 ;
        RECT 26.165 110.060 27.515 110.970 ;
        RECT 28.005 110.100 28.435 110.885 ;
        RECT 28.455 110.160 29.825 110.970 ;
        RECT 29.835 110.160 35.345 110.970 ;
        RECT 35.355 110.160 40.865 110.970 ;
        RECT 40.885 110.100 41.315 110.885 ;
        RECT 41.795 110.160 47.305 110.970 ;
        RECT 47.325 110.060 48.675 110.970 ;
        RECT 48.695 110.160 51.445 110.970 ;
        RECT 51.465 110.060 52.815 110.970 ;
        RECT 53.765 110.100 54.195 110.885 ;
        RECT 54.675 110.160 58.345 110.970 ;
        RECT 58.365 110.060 59.715 110.970 ;
        RECT 59.735 110.160 61.105 110.970 ;
        RECT 61.115 110.160 66.625 110.970 ;
        RECT 66.645 110.100 67.075 110.885 ;
        RECT 67.095 110.160 72.605 110.970 ;
        RECT 72.615 110.160 78.125 110.970 ;
        RECT 78.145 110.060 79.495 110.970 ;
        RECT 79.525 110.100 79.955 110.885 ;
        RECT 79.975 110.160 81.805 110.970 ;
        RECT 82.015 110.290 92.385 110.970 ;
        RECT 82.015 110.060 84.225 110.290 ;
        RECT 86.945 110.070 87.875 110.290 ;
        RECT 92.405 110.100 92.835 110.885 ;
        RECT 92.855 110.160 94.225 110.970 ;
        RECT 94.235 110.160 99.745 110.970 ;
        RECT 99.755 110.160 105.265 110.970 ;
        RECT 105.285 110.100 105.715 110.885 ;
        RECT 106.655 110.160 110.325 110.970 ;
        RECT 110.345 110.060 111.695 110.970 ;
        RECT 111.715 110.160 117.225 110.970 ;
        RECT 117.235 110.160 118.605 110.970 ;
      LAYER nwell ;
        RECT 11.240 108.165 118.800 109.770 ;
        RECT 20.485 54.580 29.875 66.420 ;
        RECT 31.685 54.590 41.075 66.430 ;
        RECT 42.905 54.560 52.295 66.400 ;
        RECT 54.155 54.540 63.545 66.380 ;
        RECT 65.375 54.530 74.765 66.370 ;
        RECT 76.615 54.520 86.005 66.360 ;
        RECT 87.865 54.530 97.255 66.370 ;
        RECT 99.145 54.520 108.535 66.360 ;
        RECT 110.415 54.520 119.805 66.360 ;
        RECT 121.665 54.520 131.055 66.360 ;
        RECT 132.415 54.490 139.375 66.330 ;
        RECT 20.655 49.020 23.115 53.210 ;
      LAYER pwell ;
        RECT 20.555 45.340 22.915 48.340 ;
      LAYER nwell ;
        RECT 24.735 45.940 29.125 53.130 ;
        RECT 31.855 49.030 34.315 53.220 ;
      LAYER pwell ;
        RECT 31.755 45.350 34.115 48.350 ;
      LAYER nwell ;
        RECT 35.935 45.950 40.325 53.140 ;
        RECT 43.075 49.000 45.535 53.190 ;
      LAYER pwell ;
        RECT 42.975 45.320 45.335 48.320 ;
      LAYER nwell ;
        RECT 47.155 45.920 51.545 53.110 ;
        RECT 54.325 48.980 56.785 53.170 ;
      LAYER pwell ;
        RECT 54.225 45.300 56.585 48.300 ;
      LAYER nwell ;
        RECT 58.405 45.900 62.795 53.090 ;
        RECT 65.545 48.970 68.005 53.160 ;
      LAYER pwell ;
        RECT 65.445 45.290 67.805 48.290 ;
      LAYER nwell ;
        RECT 69.625 45.890 74.015 53.080 ;
        RECT 76.785 48.960 79.245 53.150 ;
      LAYER pwell ;
        RECT 76.685 45.280 79.045 48.280 ;
      LAYER nwell ;
        RECT 80.865 45.880 85.255 53.070 ;
        RECT 88.035 48.970 90.495 53.160 ;
      LAYER pwell ;
        RECT 87.935 45.290 90.295 48.290 ;
      LAYER nwell ;
        RECT 92.115 45.890 96.505 53.080 ;
        RECT 99.315 48.960 101.775 53.150 ;
      LAYER pwell ;
        RECT 99.215 45.280 101.575 48.280 ;
      LAYER nwell ;
        RECT 103.395 45.880 107.785 53.070 ;
        RECT 110.585 48.960 113.045 53.150 ;
      LAYER pwell ;
        RECT 110.485 45.280 112.845 48.280 ;
      LAYER nwell ;
        RECT 114.665 45.880 119.055 53.070 ;
        RECT 121.835 48.960 124.295 53.150 ;
      LAYER pwell ;
        RECT 121.735 45.280 124.095 48.280 ;
      LAYER nwell ;
        RECT 125.915 45.880 130.305 53.070 ;
        RECT 19.615 32.280 24.005 39.470 ;
      LAYER pwell ;
        RECT 25.825 37.070 28.185 40.070 ;
      LAYER nwell ;
        RECT 25.625 32.200 28.085 36.390 ;
        RECT 30.895 32.280 35.285 39.470 ;
      LAYER pwell ;
        RECT 37.105 37.070 39.465 40.070 ;
      LAYER nwell ;
        RECT 36.905 32.200 39.365 36.390 ;
        RECT 42.185 32.260 46.575 39.450 ;
      LAYER pwell ;
        RECT 48.395 37.050 50.755 40.050 ;
      LAYER nwell ;
        RECT 48.195 32.180 50.655 36.370 ;
        RECT 53.405 32.260 57.795 39.450 ;
      LAYER pwell ;
        RECT 59.615 37.050 61.975 40.050 ;
      LAYER nwell ;
        RECT 59.415 32.180 61.875 36.370 ;
        RECT 64.605 32.260 68.995 39.450 ;
      LAYER pwell ;
        RECT 70.815 37.050 73.175 40.050 ;
      LAYER nwell ;
        RECT 70.615 32.180 73.075 36.370 ;
        RECT 75.895 32.250 80.285 39.440 ;
      LAYER pwell ;
        RECT 82.105 37.040 84.465 40.040 ;
      LAYER nwell ;
        RECT 81.905 32.170 84.365 36.360 ;
        RECT 87.135 32.270 91.525 39.460 ;
      LAYER pwell ;
        RECT 93.345 37.060 95.705 40.060 ;
      LAYER nwell ;
        RECT 93.145 32.190 95.605 36.380 ;
        RECT 98.345 32.290 102.735 39.480 ;
      LAYER pwell ;
        RECT 104.555 37.080 106.915 40.080 ;
      LAYER nwell ;
        RECT 104.355 32.210 106.815 36.400 ;
        RECT 109.545 32.330 113.935 39.520 ;
      LAYER pwell ;
        RECT 115.755 37.120 118.115 40.120 ;
      LAYER nwell ;
        RECT 115.555 32.250 118.015 36.440 ;
        RECT 120.755 32.350 125.145 39.540 ;
      LAYER pwell ;
        RECT 126.965 37.140 129.325 40.140 ;
      LAYER nwell ;
        RECT 126.765 32.270 129.225 36.460 ;
        RECT 18.865 18.990 28.255 30.830 ;
        RECT 30.145 18.990 39.535 30.830 ;
        RECT 41.435 18.970 50.825 30.810 ;
        RECT 52.655 18.970 62.045 30.810 ;
        RECT 63.855 18.970 73.245 30.810 ;
        RECT 75.145 18.960 84.535 30.800 ;
        RECT 86.385 18.980 95.775 30.820 ;
        RECT 97.595 19.000 106.985 30.840 ;
        RECT 108.795 19.040 118.185 30.880 ;
        RECT 120.005 19.060 129.395 30.900 ;
        RECT 131.725 19.030 138.685 30.870 ;
      LAYER li1 ;
        RECT 11.430 214.350 118.610 214.520 ;
        RECT 11.515 213.600 12.725 214.350 ;
        RECT 11.515 213.060 12.035 213.600 ;
        RECT 13.355 213.580 15.025 214.350 ;
        RECT 15.195 213.625 15.485 214.350 ;
        RECT 15.655 213.600 16.865 214.350 ;
        RECT 17.040 213.805 22.385 214.350 ;
        RECT 22.560 213.805 27.905 214.350 ;
        RECT 12.205 212.890 12.725 213.430 ;
        RECT 11.515 211.800 12.725 212.890 ;
        RECT 13.355 212.890 14.105 213.410 ;
        RECT 14.275 213.060 15.025 213.580 ;
        RECT 13.355 211.800 15.025 212.890 ;
        RECT 15.195 211.800 15.485 212.965 ;
        RECT 15.655 212.890 16.175 213.430 ;
        RECT 16.345 213.060 16.865 213.600 ;
        RECT 15.655 211.800 16.865 212.890 ;
        RECT 18.630 212.235 18.980 213.485 ;
        RECT 20.460 212.975 20.800 213.805 ;
        RECT 24.150 212.235 24.500 213.485 ;
        RECT 25.980 212.975 26.320 213.805 ;
        RECT 28.075 213.625 28.365 214.350 ;
        RECT 28.535 213.600 29.745 214.350 ;
        RECT 29.920 213.805 35.265 214.350 ;
        RECT 35.440 213.805 40.785 214.350 ;
        RECT 17.040 211.800 22.385 212.235 ;
        RECT 22.560 211.800 27.905 212.235 ;
        RECT 28.075 211.800 28.365 212.965 ;
        RECT 28.535 212.890 29.055 213.430 ;
        RECT 29.225 213.060 29.745 213.600 ;
        RECT 28.535 211.800 29.745 212.890 ;
        RECT 31.510 212.235 31.860 213.485 ;
        RECT 33.340 212.975 33.680 213.805 ;
        RECT 37.030 212.235 37.380 213.485 ;
        RECT 38.860 212.975 39.200 213.805 ;
        RECT 40.955 213.625 41.245 214.350 ;
        RECT 41.415 213.600 42.625 214.350 ;
        RECT 42.800 213.805 48.145 214.350 ;
        RECT 48.320 213.805 53.665 214.350 ;
        RECT 29.920 211.800 35.265 212.235 ;
        RECT 35.440 211.800 40.785 212.235 ;
        RECT 40.955 211.800 41.245 212.965 ;
        RECT 41.415 212.890 41.935 213.430 ;
        RECT 42.105 213.060 42.625 213.600 ;
        RECT 41.415 211.800 42.625 212.890 ;
        RECT 44.390 212.235 44.740 213.485 ;
        RECT 46.220 212.975 46.560 213.805 ;
        RECT 49.910 212.235 50.260 213.485 ;
        RECT 51.740 212.975 52.080 213.805 ;
        RECT 53.835 213.625 54.125 214.350 ;
        RECT 54.295 213.600 55.505 214.350 ;
        RECT 55.680 213.805 61.025 214.350 ;
        RECT 61.200 213.805 66.545 214.350 ;
        RECT 42.800 211.800 48.145 212.235 ;
        RECT 48.320 211.800 53.665 212.235 ;
        RECT 53.835 211.800 54.125 212.965 ;
        RECT 54.295 212.890 54.815 213.430 ;
        RECT 54.985 213.060 55.505 213.600 ;
        RECT 54.295 211.800 55.505 212.890 ;
        RECT 57.270 212.235 57.620 213.485 ;
        RECT 59.100 212.975 59.440 213.805 ;
        RECT 62.790 212.235 63.140 213.485 ;
        RECT 64.620 212.975 64.960 213.805 ;
        RECT 66.715 213.625 67.005 214.350 ;
        RECT 67.175 213.600 68.385 214.350 ;
        RECT 68.560 213.805 73.905 214.350 ;
        RECT 74.080 213.805 79.425 214.350 ;
        RECT 55.680 211.800 61.025 212.235 ;
        RECT 61.200 211.800 66.545 212.235 ;
        RECT 66.715 211.800 67.005 212.965 ;
        RECT 67.175 212.890 67.695 213.430 ;
        RECT 67.865 213.060 68.385 213.600 ;
        RECT 67.175 211.800 68.385 212.890 ;
        RECT 70.150 212.235 70.500 213.485 ;
        RECT 71.980 212.975 72.320 213.805 ;
        RECT 75.670 212.235 76.020 213.485 ;
        RECT 77.500 212.975 77.840 213.805 ;
        RECT 79.595 213.625 79.885 214.350 ;
        RECT 80.055 213.600 81.265 214.350 ;
        RECT 81.440 213.805 86.785 214.350 ;
        RECT 86.960 213.805 92.305 214.350 ;
        RECT 68.560 211.800 73.905 212.235 ;
        RECT 74.080 211.800 79.425 212.235 ;
        RECT 79.595 211.800 79.885 212.965 ;
        RECT 80.055 212.890 80.575 213.430 ;
        RECT 80.745 213.060 81.265 213.600 ;
        RECT 80.055 211.800 81.265 212.890 ;
        RECT 83.030 212.235 83.380 213.485 ;
        RECT 84.860 212.975 85.200 213.805 ;
        RECT 88.550 212.235 88.900 213.485 ;
        RECT 90.380 212.975 90.720 213.805 ;
        RECT 92.475 213.625 92.765 214.350 ;
        RECT 92.935 213.600 94.145 214.350 ;
        RECT 94.320 213.805 99.665 214.350 ;
        RECT 99.840 213.805 105.185 214.350 ;
        RECT 81.440 211.800 86.785 212.235 ;
        RECT 86.960 211.800 92.305 212.235 ;
        RECT 92.475 211.800 92.765 212.965 ;
        RECT 92.935 212.890 93.455 213.430 ;
        RECT 93.625 213.060 94.145 213.600 ;
        RECT 92.935 211.800 94.145 212.890 ;
        RECT 95.910 212.235 96.260 213.485 ;
        RECT 97.740 212.975 98.080 213.805 ;
        RECT 101.430 212.235 101.780 213.485 ;
        RECT 103.260 212.975 103.600 213.805 ;
        RECT 105.355 213.625 105.645 214.350 ;
        RECT 106.280 213.805 111.625 214.350 ;
        RECT 111.800 213.805 117.145 214.350 ;
        RECT 94.320 211.800 99.665 212.235 ;
        RECT 99.840 211.800 105.185 212.235 ;
        RECT 105.355 211.800 105.645 212.965 ;
        RECT 107.870 212.235 108.220 213.485 ;
        RECT 109.700 212.975 110.040 213.805 ;
        RECT 113.390 212.235 113.740 213.485 ;
        RECT 115.220 212.975 115.560 213.805 ;
        RECT 117.315 213.600 118.525 214.350 ;
        RECT 117.315 212.890 117.835 213.430 ;
        RECT 118.005 213.060 118.525 213.600 ;
        RECT 106.280 211.800 111.625 212.235 ;
        RECT 111.800 211.800 117.145 212.235 ;
        RECT 117.315 211.800 118.525 212.890 ;
        RECT 11.430 211.630 118.610 211.800 ;
        RECT 11.515 210.540 12.725 211.630 ;
        RECT 11.515 209.830 12.035 210.370 ;
        RECT 12.205 210.000 12.725 210.540 ;
        RECT 13.355 210.540 15.025 211.630 ;
        RECT 13.355 210.020 14.105 210.540 ;
        RECT 15.195 210.465 15.485 211.630 ;
        RECT 16.115 210.540 18.705 211.630 ;
        RECT 18.880 211.195 24.225 211.630 ;
        RECT 24.400 211.195 29.745 211.630 ;
        RECT 29.920 211.195 35.265 211.630 ;
        RECT 35.440 211.195 40.785 211.630 ;
        RECT 14.275 209.850 15.025 210.370 ;
        RECT 16.115 210.020 17.325 210.540 ;
        RECT 17.495 209.850 18.705 210.370 ;
        RECT 20.470 209.945 20.820 211.195 ;
        RECT 11.515 209.080 12.725 209.830 ;
        RECT 13.355 209.080 15.025 209.850 ;
        RECT 15.195 209.080 15.485 209.805 ;
        RECT 16.115 209.080 18.705 209.850 ;
        RECT 22.300 209.625 22.640 210.455 ;
        RECT 25.990 209.945 26.340 211.195 ;
        RECT 27.820 209.625 28.160 210.455 ;
        RECT 31.510 209.945 31.860 211.195 ;
        RECT 33.340 209.625 33.680 210.455 ;
        RECT 37.030 209.945 37.380 211.195 ;
        RECT 40.955 210.465 41.245 211.630 ;
        RECT 41.875 210.540 43.545 211.630 ;
        RECT 43.720 211.195 49.065 211.630 ;
        RECT 49.240 211.195 54.585 211.630 ;
        RECT 38.860 209.625 39.200 210.455 ;
        RECT 41.875 210.020 42.625 210.540 ;
        RECT 42.795 209.850 43.545 210.370 ;
        RECT 45.310 209.945 45.660 211.195 ;
        RECT 18.880 209.080 24.225 209.625 ;
        RECT 24.400 209.080 29.745 209.625 ;
        RECT 29.920 209.080 35.265 209.625 ;
        RECT 35.440 209.080 40.785 209.625 ;
        RECT 40.955 209.080 41.245 209.805 ;
        RECT 41.875 209.080 43.545 209.850 ;
        RECT 47.140 209.625 47.480 210.455 ;
        RECT 50.830 209.945 51.180 211.195 ;
        RECT 52.660 209.625 53.000 210.455 ;
        RECT 54.760 210.440 55.015 211.320 ;
        RECT 55.185 210.490 55.490 211.630 ;
        RECT 55.830 211.250 56.160 211.630 ;
        RECT 56.340 211.080 56.510 211.370 ;
        RECT 56.680 211.170 56.930 211.630 ;
        RECT 55.710 210.910 56.510 211.080 ;
        RECT 57.100 211.120 57.970 211.460 ;
        RECT 54.760 209.790 54.970 210.440 ;
        RECT 55.710 210.320 55.880 210.910 ;
        RECT 57.100 210.740 57.270 211.120 ;
        RECT 58.205 211.000 58.375 211.460 ;
        RECT 58.545 211.170 58.915 211.630 ;
        RECT 59.210 211.030 59.380 211.370 ;
        RECT 59.550 211.200 59.880 211.630 ;
        RECT 60.115 211.030 60.285 211.370 ;
        RECT 56.050 210.570 57.270 210.740 ;
        RECT 57.440 210.660 57.900 210.950 ;
        RECT 58.205 210.830 58.765 211.000 ;
        RECT 59.210 210.860 60.285 211.030 ;
        RECT 60.455 211.130 61.135 211.460 ;
        RECT 61.350 211.130 61.600 211.460 ;
        RECT 61.770 211.170 62.020 211.630 ;
        RECT 58.595 210.690 58.765 210.830 ;
        RECT 57.440 210.650 58.405 210.660 ;
        RECT 57.100 210.480 57.270 210.570 ;
        RECT 57.730 210.490 58.405 210.650 ;
        RECT 55.140 210.290 55.880 210.320 ;
        RECT 55.140 209.990 56.055 210.290 ;
        RECT 55.730 209.815 56.055 209.990 ;
        RECT 43.720 209.080 49.065 209.625 ;
        RECT 49.240 209.080 54.585 209.625 ;
        RECT 54.760 209.260 55.015 209.790 ;
        RECT 55.185 209.080 55.490 209.540 ;
        RECT 55.735 209.460 56.055 209.815 ;
        RECT 56.225 210.030 56.765 210.400 ;
        RECT 57.100 210.310 57.505 210.480 ;
        RECT 56.225 209.630 56.465 210.030 ;
        RECT 56.945 209.860 57.165 210.140 ;
        RECT 56.635 209.690 57.165 209.860 ;
        RECT 56.635 209.460 56.805 209.690 ;
        RECT 57.335 209.530 57.505 210.310 ;
        RECT 57.675 209.700 58.025 210.320 ;
        RECT 58.195 209.700 58.405 210.490 ;
        RECT 58.595 210.520 60.095 210.690 ;
        RECT 58.595 209.830 58.765 210.520 ;
        RECT 60.455 210.350 60.625 211.130 ;
        RECT 61.430 211.000 61.600 211.130 ;
        RECT 58.935 210.180 60.625 210.350 ;
        RECT 60.795 210.570 61.260 210.960 ;
        RECT 61.430 210.830 61.825 211.000 ;
        RECT 58.935 210.000 59.105 210.180 ;
        RECT 55.735 209.290 56.805 209.460 ;
        RECT 56.975 209.080 57.165 209.520 ;
        RECT 57.335 209.250 58.285 209.530 ;
        RECT 58.595 209.440 58.855 209.830 ;
        RECT 59.275 209.760 60.065 210.010 ;
        RECT 58.505 209.270 58.855 209.440 ;
        RECT 59.065 209.080 59.395 209.540 ;
        RECT 60.270 209.470 60.440 210.180 ;
        RECT 60.795 209.980 60.965 210.570 ;
        RECT 60.610 209.760 60.965 209.980 ;
        RECT 61.135 209.760 61.485 210.380 ;
        RECT 61.655 209.470 61.825 210.830 ;
        RECT 62.190 210.660 62.515 211.445 ;
        RECT 61.995 209.610 62.455 210.660 ;
        RECT 60.270 209.300 61.125 209.470 ;
        RECT 61.330 209.300 61.825 209.470 ;
        RECT 61.995 209.080 62.325 209.440 ;
        RECT 62.685 209.340 62.855 211.460 ;
        RECT 63.025 211.130 63.355 211.630 ;
        RECT 63.525 210.960 63.780 211.460 ;
        RECT 63.030 210.790 63.780 210.960 ;
        RECT 63.030 209.800 63.260 210.790 ;
        RECT 63.430 209.970 63.780 210.620 ;
        RECT 63.955 210.540 66.545 211.630 ;
        RECT 63.955 210.020 65.165 210.540 ;
        RECT 66.715 210.465 67.005 211.630 ;
        RECT 68.155 210.490 68.365 211.630 ;
        RECT 68.535 210.480 68.865 211.460 ;
        RECT 69.035 210.490 69.265 211.630 ;
        RECT 70.400 211.195 75.745 211.630 ;
        RECT 75.920 211.195 81.265 211.630 ;
        RECT 81.440 211.195 86.785 211.630 ;
        RECT 86.960 211.195 92.305 211.630 ;
        RECT 65.335 209.850 66.545 210.370 ;
        RECT 63.030 209.630 63.780 209.800 ;
        RECT 63.025 209.080 63.355 209.460 ;
        RECT 63.525 209.340 63.780 209.630 ;
        RECT 63.955 209.080 66.545 209.850 ;
        RECT 66.715 209.080 67.005 209.805 ;
        RECT 68.155 209.080 68.365 209.900 ;
        RECT 68.535 209.880 68.785 210.480 ;
        RECT 68.955 210.070 69.285 210.320 ;
        RECT 71.990 209.945 72.340 211.195 ;
        RECT 68.535 209.250 68.865 209.880 ;
        RECT 69.035 209.080 69.265 209.900 ;
        RECT 73.820 209.625 74.160 210.455 ;
        RECT 77.510 209.945 77.860 211.195 ;
        RECT 79.340 209.625 79.680 210.455 ;
        RECT 83.030 209.945 83.380 211.195 ;
        RECT 84.860 209.625 85.200 210.455 ;
        RECT 88.550 209.945 88.900 211.195 ;
        RECT 92.475 210.465 92.765 211.630 ;
        RECT 93.395 210.540 95.065 211.630 ;
        RECT 95.240 211.195 100.585 211.630 ;
        RECT 100.760 211.195 106.105 211.630 ;
        RECT 106.280 211.195 111.625 211.630 ;
        RECT 111.800 211.195 117.145 211.630 ;
        RECT 90.380 209.625 90.720 210.455 ;
        RECT 93.395 210.020 94.145 210.540 ;
        RECT 94.315 209.850 95.065 210.370 ;
        RECT 96.830 209.945 97.180 211.195 ;
        RECT 70.400 209.080 75.745 209.625 ;
        RECT 75.920 209.080 81.265 209.625 ;
        RECT 81.440 209.080 86.785 209.625 ;
        RECT 86.960 209.080 92.305 209.625 ;
        RECT 92.475 209.080 92.765 209.805 ;
        RECT 93.395 209.080 95.065 209.850 ;
        RECT 98.660 209.625 99.000 210.455 ;
        RECT 102.350 209.945 102.700 211.195 ;
        RECT 104.180 209.625 104.520 210.455 ;
        RECT 107.870 209.945 108.220 211.195 ;
        RECT 109.700 209.625 110.040 210.455 ;
        RECT 113.390 209.945 113.740 211.195 ;
        RECT 117.315 210.540 118.525 211.630 ;
        RECT 115.220 209.625 115.560 210.455 ;
        RECT 117.315 210.000 117.835 210.540 ;
        RECT 118.005 209.830 118.525 210.370 ;
        RECT 95.240 209.080 100.585 209.625 ;
        RECT 100.760 209.080 106.105 209.625 ;
        RECT 106.280 209.080 111.625 209.625 ;
        RECT 111.800 209.080 117.145 209.625 ;
        RECT 117.315 209.080 118.525 209.830 ;
        RECT 11.430 208.910 118.610 209.080 ;
        RECT 11.515 208.160 12.725 208.910 ;
        RECT 11.515 207.620 12.035 208.160 ;
        RECT 13.355 208.140 16.865 208.910 ;
        RECT 17.040 208.365 22.385 208.910 ;
        RECT 22.560 208.365 27.905 208.910 ;
        RECT 12.205 207.450 12.725 207.990 ;
        RECT 11.515 206.360 12.725 207.450 ;
        RECT 13.355 207.450 15.045 207.970 ;
        RECT 15.215 207.620 16.865 208.140 ;
        RECT 13.355 206.360 16.865 207.450 ;
        RECT 18.630 206.795 18.980 208.045 ;
        RECT 20.460 207.535 20.800 208.365 ;
        RECT 24.150 206.795 24.500 208.045 ;
        RECT 25.980 207.535 26.320 208.365 ;
        RECT 28.075 208.185 28.365 208.910 ;
        RECT 29.000 208.365 34.345 208.910 ;
        RECT 34.520 208.365 39.865 208.910 ;
        RECT 40.040 208.365 45.385 208.910 ;
        RECT 45.560 208.365 50.905 208.910 ;
        RECT 17.040 206.360 22.385 206.795 ;
        RECT 22.560 206.360 27.905 206.795 ;
        RECT 28.075 206.360 28.365 207.525 ;
        RECT 30.590 206.795 30.940 208.045 ;
        RECT 32.420 207.535 32.760 208.365 ;
        RECT 36.110 206.795 36.460 208.045 ;
        RECT 37.940 207.535 38.280 208.365 ;
        RECT 41.630 206.795 41.980 208.045 ;
        RECT 43.460 207.535 43.800 208.365 ;
        RECT 47.150 206.795 47.500 208.045 ;
        RECT 48.980 207.535 49.320 208.365 ;
        RECT 51.135 208.090 51.345 208.910 ;
        RECT 51.515 208.110 51.845 208.740 ;
        RECT 51.515 207.510 51.765 208.110 ;
        RECT 52.015 208.090 52.245 208.910 ;
        RECT 52.495 208.090 52.725 208.910 ;
        RECT 52.895 208.110 53.225 208.740 ;
        RECT 51.935 207.670 52.265 207.920 ;
        RECT 52.475 207.670 52.805 207.920 ;
        RECT 52.975 207.510 53.225 208.110 ;
        RECT 53.395 208.090 53.605 208.910 ;
        RECT 53.835 208.185 54.125 208.910 ;
        RECT 54.300 208.200 54.555 208.730 ;
        RECT 54.725 208.450 55.030 208.910 ;
        RECT 55.275 208.530 56.345 208.700 ;
        RECT 54.300 207.550 54.510 208.200 ;
        RECT 55.275 208.175 55.595 208.530 ;
        RECT 55.270 208.000 55.595 208.175 ;
        RECT 54.680 207.700 55.595 208.000 ;
        RECT 55.765 207.960 56.005 208.360 ;
        RECT 56.175 208.300 56.345 208.530 ;
        RECT 56.515 208.470 56.705 208.910 ;
        RECT 56.875 208.460 57.825 208.740 ;
        RECT 58.045 208.550 58.395 208.720 ;
        RECT 56.175 208.130 56.705 208.300 ;
        RECT 54.680 207.670 55.420 207.700 ;
        RECT 29.000 206.360 34.345 206.795 ;
        RECT 34.520 206.360 39.865 206.795 ;
        RECT 40.040 206.360 45.385 206.795 ;
        RECT 45.560 206.360 50.905 206.795 ;
        RECT 51.135 206.360 51.345 207.500 ;
        RECT 51.515 206.530 51.845 207.510 ;
        RECT 52.015 206.360 52.245 207.500 ;
        RECT 52.495 206.360 52.725 207.500 ;
        RECT 52.895 206.530 53.225 207.510 ;
        RECT 53.395 206.360 53.605 207.500 ;
        RECT 53.835 206.360 54.125 207.525 ;
        RECT 54.300 206.670 54.555 207.550 ;
        RECT 54.725 206.360 55.030 207.500 ;
        RECT 55.250 207.080 55.420 207.670 ;
        RECT 55.765 207.590 56.305 207.960 ;
        RECT 56.485 207.850 56.705 208.130 ;
        RECT 56.875 207.680 57.045 208.460 ;
        RECT 56.640 207.510 57.045 207.680 ;
        RECT 57.215 207.670 57.565 208.290 ;
        RECT 56.640 207.420 56.810 207.510 ;
        RECT 57.735 207.500 57.945 208.290 ;
        RECT 55.590 207.250 56.810 207.420 ;
        RECT 57.270 207.340 57.945 207.500 ;
        RECT 55.250 206.910 56.050 207.080 ;
        RECT 55.370 206.360 55.700 206.740 ;
        RECT 55.880 206.620 56.050 206.910 ;
        RECT 56.640 206.870 56.810 207.250 ;
        RECT 56.980 207.330 57.945 207.340 ;
        RECT 58.135 208.160 58.395 208.550 ;
        RECT 58.605 208.450 58.935 208.910 ;
        RECT 59.810 208.520 60.665 208.690 ;
        RECT 60.870 208.520 61.365 208.690 ;
        RECT 61.535 208.550 61.865 208.910 ;
        RECT 58.135 207.470 58.305 208.160 ;
        RECT 58.475 207.810 58.645 207.990 ;
        RECT 58.815 207.980 59.605 208.230 ;
        RECT 59.810 207.810 59.980 208.520 ;
        RECT 60.150 208.010 60.505 208.230 ;
        RECT 58.475 207.640 60.165 207.810 ;
        RECT 56.980 207.040 57.440 207.330 ;
        RECT 58.135 207.300 59.635 207.470 ;
        RECT 58.135 207.160 58.305 207.300 ;
        RECT 57.745 206.990 58.305 207.160 ;
        RECT 56.220 206.360 56.470 206.820 ;
        RECT 56.640 206.530 57.510 206.870 ;
        RECT 57.745 206.530 57.915 206.990 ;
        RECT 58.750 206.960 59.825 207.130 ;
        RECT 58.085 206.360 58.455 206.820 ;
        RECT 58.750 206.620 58.920 206.960 ;
        RECT 59.090 206.360 59.420 206.790 ;
        RECT 59.655 206.620 59.825 206.960 ;
        RECT 59.995 206.860 60.165 207.640 ;
        RECT 60.335 207.420 60.505 208.010 ;
        RECT 60.675 207.610 61.025 208.230 ;
        RECT 60.335 207.030 60.800 207.420 ;
        RECT 61.195 207.160 61.365 208.520 ;
        RECT 61.535 207.330 61.995 208.380 ;
        RECT 60.970 206.990 61.365 207.160 ;
        RECT 60.970 206.860 61.140 206.990 ;
        RECT 59.995 206.530 60.675 206.860 ;
        RECT 60.890 206.530 61.140 206.860 ;
        RECT 61.310 206.360 61.560 206.820 ;
        RECT 61.730 206.545 62.055 207.330 ;
        RECT 62.225 206.530 62.395 208.650 ;
        RECT 62.565 208.530 62.895 208.910 ;
        RECT 63.065 208.360 63.320 208.650 ;
        RECT 62.570 208.190 63.320 208.360 ;
        RECT 62.570 207.200 62.800 208.190 ;
        RECT 63.495 208.160 64.705 208.910 ;
        RECT 62.970 207.370 63.320 208.020 ;
        RECT 63.495 207.450 64.015 207.990 ;
        RECT 64.185 207.620 64.705 208.160 ;
        RECT 64.880 208.200 65.135 208.730 ;
        RECT 65.305 208.450 65.610 208.910 ;
        RECT 65.855 208.530 66.925 208.700 ;
        RECT 64.880 207.550 65.090 208.200 ;
        RECT 65.855 208.175 66.175 208.530 ;
        RECT 65.850 208.000 66.175 208.175 ;
        RECT 65.260 207.700 66.175 208.000 ;
        RECT 66.345 207.960 66.585 208.360 ;
        RECT 66.755 208.300 66.925 208.530 ;
        RECT 67.095 208.470 67.285 208.910 ;
        RECT 67.455 208.460 68.405 208.740 ;
        RECT 68.625 208.550 68.975 208.720 ;
        RECT 66.755 208.130 67.285 208.300 ;
        RECT 65.260 207.670 66.000 207.700 ;
        RECT 62.570 207.030 63.320 207.200 ;
        RECT 62.565 206.360 62.895 206.860 ;
        RECT 63.065 206.530 63.320 207.030 ;
        RECT 63.495 206.360 64.705 207.450 ;
        RECT 64.880 206.670 65.135 207.550 ;
        RECT 65.305 206.360 65.610 207.500 ;
        RECT 65.830 207.080 66.000 207.670 ;
        RECT 66.345 207.590 66.885 207.960 ;
        RECT 67.065 207.850 67.285 208.130 ;
        RECT 67.455 207.680 67.625 208.460 ;
        RECT 67.220 207.510 67.625 207.680 ;
        RECT 67.795 207.670 68.145 208.290 ;
        RECT 67.220 207.420 67.390 207.510 ;
        RECT 68.315 207.500 68.525 208.290 ;
        RECT 66.170 207.250 67.390 207.420 ;
        RECT 67.850 207.340 68.525 207.500 ;
        RECT 65.830 206.910 66.630 207.080 ;
        RECT 65.950 206.360 66.280 206.740 ;
        RECT 66.460 206.620 66.630 206.910 ;
        RECT 67.220 206.870 67.390 207.250 ;
        RECT 67.560 207.330 68.525 207.340 ;
        RECT 68.715 208.160 68.975 208.550 ;
        RECT 69.185 208.450 69.515 208.910 ;
        RECT 70.390 208.520 71.245 208.690 ;
        RECT 71.450 208.520 71.945 208.690 ;
        RECT 72.115 208.550 72.445 208.910 ;
        RECT 68.715 207.470 68.885 208.160 ;
        RECT 69.055 207.810 69.225 207.990 ;
        RECT 69.395 207.980 70.185 208.230 ;
        RECT 70.390 207.810 70.560 208.520 ;
        RECT 70.730 208.010 71.085 208.230 ;
        RECT 69.055 207.640 70.745 207.810 ;
        RECT 67.560 207.040 68.020 207.330 ;
        RECT 68.715 207.300 70.215 207.470 ;
        RECT 68.715 207.160 68.885 207.300 ;
        RECT 68.325 206.990 68.885 207.160 ;
        RECT 66.800 206.360 67.050 206.820 ;
        RECT 67.220 206.530 68.090 206.870 ;
        RECT 68.325 206.530 68.495 206.990 ;
        RECT 69.330 206.960 70.405 207.130 ;
        RECT 68.665 206.360 69.035 206.820 ;
        RECT 69.330 206.620 69.500 206.960 ;
        RECT 69.670 206.360 70.000 206.790 ;
        RECT 70.235 206.620 70.405 206.960 ;
        RECT 70.575 206.860 70.745 207.640 ;
        RECT 70.915 207.420 71.085 208.010 ;
        RECT 71.255 207.610 71.605 208.230 ;
        RECT 70.915 207.030 71.380 207.420 ;
        RECT 71.775 207.160 71.945 208.520 ;
        RECT 72.115 207.330 72.575 208.380 ;
        RECT 71.550 206.990 71.945 207.160 ;
        RECT 71.550 206.860 71.720 206.990 ;
        RECT 70.575 206.530 71.255 206.860 ;
        RECT 71.470 206.530 71.720 206.860 ;
        RECT 71.890 206.360 72.140 206.820 ;
        RECT 72.310 206.545 72.635 207.330 ;
        RECT 72.805 206.530 72.975 208.650 ;
        RECT 73.145 208.530 73.475 208.910 ;
        RECT 73.645 208.360 73.900 208.650 ;
        RECT 74.080 208.365 79.425 208.910 ;
        RECT 73.150 208.190 73.900 208.360 ;
        RECT 73.150 207.200 73.380 208.190 ;
        RECT 73.550 207.370 73.900 208.020 ;
        RECT 73.150 207.030 73.900 207.200 ;
        RECT 73.145 206.360 73.475 206.860 ;
        RECT 73.645 206.530 73.900 207.030 ;
        RECT 75.670 206.795 76.020 208.045 ;
        RECT 77.500 207.535 77.840 208.365 ;
        RECT 79.595 208.185 79.885 208.910 ;
        RECT 80.055 208.160 81.265 208.910 ;
        RECT 81.440 208.365 86.785 208.910 ;
        RECT 86.960 208.365 92.305 208.910 ;
        RECT 74.080 206.360 79.425 206.795 ;
        RECT 79.595 206.360 79.885 207.525 ;
        RECT 80.055 207.450 80.575 207.990 ;
        RECT 80.745 207.620 81.265 208.160 ;
        RECT 80.055 206.360 81.265 207.450 ;
        RECT 83.030 206.795 83.380 208.045 ;
        RECT 84.860 207.535 85.200 208.365 ;
        RECT 88.550 206.795 88.900 208.045 ;
        RECT 90.380 207.535 90.720 208.365 ;
        RECT 92.480 208.200 92.735 208.730 ;
        RECT 92.905 208.450 93.210 208.910 ;
        RECT 93.455 208.530 94.525 208.700 ;
        RECT 92.480 207.550 92.690 208.200 ;
        RECT 93.455 208.175 93.775 208.530 ;
        RECT 93.450 208.000 93.775 208.175 ;
        RECT 92.860 207.700 93.775 208.000 ;
        RECT 93.945 207.960 94.185 208.360 ;
        RECT 94.355 208.300 94.525 208.530 ;
        RECT 94.695 208.470 94.885 208.910 ;
        RECT 95.055 208.460 96.005 208.740 ;
        RECT 96.225 208.550 96.575 208.720 ;
        RECT 94.355 208.130 94.885 208.300 ;
        RECT 92.860 207.670 93.600 207.700 ;
        RECT 81.440 206.360 86.785 206.795 ;
        RECT 86.960 206.360 92.305 206.795 ;
        RECT 92.480 206.670 92.735 207.550 ;
        RECT 92.905 206.360 93.210 207.500 ;
        RECT 93.430 207.080 93.600 207.670 ;
        RECT 93.945 207.590 94.485 207.960 ;
        RECT 94.665 207.850 94.885 208.130 ;
        RECT 95.055 207.680 95.225 208.460 ;
        RECT 94.820 207.510 95.225 207.680 ;
        RECT 95.395 207.670 95.745 208.290 ;
        RECT 94.820 207.420 94.990 207.510 ;
        RECT 95.915 207.500 96.125 208.290 ;
        RECT 93.770 207.250 94.990 207.420 ;
        RECT 95.450 207.340 96.125 207.500 ;
        RECT 93.430 206.910 94.230 207.080 ;
        RECT 93.550 206.360 93.880 206.740 ;
        RECT 94.060 206.620 94.230 206.910 ;
        RECT 94.820 206.870 94.990 207.250 ;
        RECT 95.160 207.330 96.125 207.340 ;
        RECT 96.315 208.160 96.575 208.550 ;
        RECT 96.785 208.450 97.115 208.910 ;
        RECT 97.990 208.520 98.845 208.690 ;
        RECT 99.050 208.520 99.545 208.690 ;
        RECT 99.715 208.550 100.045 208.910 ;
        RECT 96.315 207.470 96.485 208.160 ;
        RECT 96.655 207.810 96.825 207.990 ;
        RECT 96.995 207.980 97.785 208.230 ;
        RECT 97.990 207.810 98.160 208.520 ;
        RECT 98.330 208.010 98.685 208.230 ;
        RECT 96.655 207.640 98.345 207.810 ;
        RECT 95.160 207.040 95.620 207.330 ;
        RECT 96.315 207.300 97.815 207.470 ;
        RECT 96.315 207.160 96.485 207.300 ;
        RECT 95.925 206.990 96.485 207.160 ;
        RECT 94.400 206.360 94.650 206.820 ;
        RECT 94.820 206.530 95.690 206.870 ;
        RECT 95.925 206.530 96.095 206.990 ;
        RECT 96.930 206.960 98.005 207.130 ;
        RECT 96.265 206.360 96.635 206.820 ;
        RECT 96.930 206.620 97.100 206.960 ;
        RECT 97.270 206.360 97.600 206.790 ;
        RECT 97.835 206.620 98.005 206.960 ;
        RECT 98.175 206.860 98.345 207.640 ;
        RECT 98.515 207.420 98.685 208.010 ;
        RECT 98.855 207.610 99.205 208.230 ;
        RECT 98.515 207.030 98.980 207.420 ;
        RECT 99.375 207.160 99.545 208.520 ;
        RECT 99.715 207.330 100.175 208.380 ;
        RECT 99.150 206.990 99.545 207.160 ;
        RECT 99.150 206.860 99.320 206.990 ;
        RECT 98.175 206.530 98.855 206.860 ;
        RECT 99.070 206.530 99.320 206.860 ;
        RECT 99.490 206.360 99.740 206.820 ;
        RECT 99.910 206.545 100.235 207.330 ;
        RECT 100.405 206.530 100.575 208.650 ;
        RECT 100.745 208.530 101.075 208.910 ;
        RECT 101.245 208.360 101.500 208.650 ;
        RECT 100.750 208.190 101.500 208.360 ;
        RECT 100.750 207.200 100.980 208.190 ;
        RECT 101.675 208.140 105.185 208.910 ;
        RECT 105.355 208.185 105.645 208.910 ;
        RECT 106.280 208.365 111.625 208.910 ;
        RECT 111.800 208.365 117.145 208.910 ;
        RECT 101.150 207.370 101.500 208.020 ;
        RECT 101.675 207.450 103.365 207.970 ;
        RECT 103.535 207.620 105.185 208.140 ;
        RECT 100.750 207.030 101.500 207.200 ;
        RECT 100.745 206.360 101.075 206.860 ;
        RECT 101.245 206.530 101.500 207.030 ;
        RECT 101.675 206.360 105.185 207.450 ;
        RECT 105.355 206.360 105.645 207.525 ;
        RECT 107.870 206.795 108.220 208.045 ;
        RECT 109.700 207.535 110.040 208.365 ;
        RECT 113.390 206.795 113.740 208.045 ;
        RECT 115.220 207.535 115.560 208.365 ;
        RECT 117.315 208.160 118.525 208.910 ;
        RECT 117.315 207.450 117.835 207.990 ;
        RECT 118.005 207.620 118.525 208.160 ;
        RECT 106.280 206.360 111.625 206.795 ;
        RECT 111.800 206.360 117.145 206.795 ;
        RECT 117.315 206.360 118.525 207.450 ;
        RECT 11.430 206.190 118.610 206.360 ;
        RECT 11.515 205.100 12.725 206.190 ;
        RECT 11.515 204.390 12.035 204.930 ;
        RECT 12.205 204.560 12.725 205.100 ;
        RECT 13.355 205.100 15.025 206.190 ;
        RECT 13.355 204.580 14.105 205.100 ;
        RECT 15.195 205.025 15.485 206.190 ;
        RECT 16.115 205.100 18.705 206.190 ;
        RECT 18.880 205.755 24.225 206.190 ;
        RECT 24.400 205.755 29.745 206.190 ;
        RECT 29.920 205.755 35.265 206.190 ;
        RECT 35.440 205.755 40.785 206.190 ;
        RECT 14.275 204.410 15.025 204.930 ;
        RECT 16.115 204.580 17.325 205.100 ;
        RECT 17.495 204.410 18.705 204.930 ;
        RECT 20.470 204.505 20.820 205.755 ;
        RECT 11.515 203.640 12.725 204.390 ;
        RECT 13.355 203.640 15.025 204.410 ;
        RECT 15.195 203.640 15.485 204.365 ;
        RECT 16.115 203.640 18.705 204.410 ;
        RECT 22.300 204.185 22.640 205.015 ;
        RECT 25.990 204.505 26.340 205.755 ;
        RECT 27.820 204.185 28.160 205.015 ;
        RECT 31.510 204.505 31.860 205.755 ;
        RECT 33.340 204.185 33.680 205.015 ;
        RECT 37.030 204.505 37.380 205.755 ;
        RECT 40.955 205.025 41.245 206.190 ;
        RECT 41.880 205.755 47.225 206.190 ;
        RECT 47.400 205.755 52.745 206.190 ;
        RECT 38.860 204.185 39.200 205.015 ;
        RECT 43.470 204.505 43.820 205.755 ;
        RECT 18.880 203.640 24.225 204.185 ;
        RECT 24.400 203.640 29.745 204.185 ;
        RECT 29.920 203.640 35.265 204.185 ;
        RECT 35.440 203.640 40.785 204.185 ;
        RECT 40.955 203.640 41.245 204.365 ;
        RECT 45.300 204.185 45.640 205.015 ;
        RECT 48.990 204.505 49.340 205.755 ;
        RECT 52.920 205.040 53.180 206.190 ;
        RECT 53.355 205.115 53.610 206.020 ;
        RECT 53.780 205.430 54.110 206.190 ;
        RECT 54.325 205.260 54.495 206.020 ;
        RECT 50.820 204.185 51.160 205.015 ;
        RECT 41.880 203.640 47.225 204.185 ;
        RECT 47.400 203.640 52.745 204.185 ;
        RECT 52.920 203.640 53.180 204.480 ;
        RECT 53.355 204.385 53.525 205.115 ;
        RECT 53.780 205.090 54.495 205.260 ;
        RECT 53.780 204.880 53.950 205.090 ;
        RECT 54.760 205.040 55.020 206.190 ;
        RECT 55.195 205.115 55.450 206.020 ;
        RECT 55.620 205.430 55.950 206.190 ;
        RECT 56.165 205.260 56.335 206.020 ;
        RECT 53.695 204.550 53.950 204.880 ;
        RECT 53.355 203.810 53.610 204.385 ;
        RECT 53.780 204.360 53.950 204.550 ;
        RECT 54.230 204.540 54.585 204.910 ;
        RECT 53.780 204.190 54.495 204.360 ;
        RECT 53.780 203.640 54.110 204.020 ;
        RECT 54.325 203.810 54.495 204.190 ;
        RECT 54.760 203.640 55.020 204.480 ;
        RECT 55.195 204.385 55.365 205.115 ;
        RECT 55.620 205.090 56.335 205.260 ;
        RECT 55.620 204.880 55.790 205.090 ;
        RECT 56.595 205.050 56.855 206.020 ;
        RECT 57.050 205.780 57.380 206.190 ;
        RECT 57.580 205.600 57.750 206.020 ;
        RECT 57.965 205.780 58.635 206.190 ;
        RECT 58.870 205.600 59.040 206.020 ;
        RECT 59.345 205.750 59.675 206.190 ;
        RECT 57.025 205.430 59.040 205.600 ;
        RECT 59.845 205.570 60.020 206.020 ;
        RECT 55.535 204.550 55.790 204.880 ;
        RECT 55.195 203.810 55.450 204.385 ;
        RECT 55.620 204.360 55.790 204.550 ;
        RECT 56.070 204.540 56.425 204.910 ;
        RECT 56.595 204.360 56.765 205.050 ;
        RECT 57.025 204.880 57.195 205.430 ;
        RECT 56.935 204.550 57.195 204.880 ;
        RECT 55.620 204.190 56.335 204.360 ;
        RECT 55.620 203.640 55.950 204.020 ;
        RECT 56.165 203.810 56.335 204.190 ;
        RECT 56.595 203.895 56.935 204.360 ;
        RECT 57.365 204.220 57.705 205.250 ;
        RECT 57.895 204.830 58.165 205.250 ;
        RECT 57.895 204.660 58.205 204.830 ;
        RECT 56.600 203.850 56.935 203.895 ;
        RECT 57.105 203.640 57.435 204.020 ;
        RECT 57.895 203.975 58.165 204.660 ;
        RECT 58.390 203.975 58.670 205.250 ;
        RECT 58.870 204.140 59.040 205.430 ;
        RECT 59.390 205.400 60.020 205.570 ;
        RECT 59.390 204.880 59.560 205.400 ;
        RECT 61.195 205.320 61.470 206.020 ;
        RECT 61.640 205.645 61.895 206.190 ;
        RECT 62.065 205.680 62.545 206.020 ;
        RECT 62.720 205.635 63.325 206.190 ;
        RECT 63.515 205.680 63.815 206.190 ;
        RECT 63.985 205.680 64.365 205.850 ;
        RECT 64.945 205.680 65.575 206.190 ;
        RECT 62.710 205.535 63.325 205.635 ;
        RECT 62.710 205.510 62.895 205.535 ;
        RECT 63.985 205.510 64.155 205.680 ;
        RECT 65.745 205.510 66.075 206.020 ;
        RECT 66.245 205.680 66.545 206.190 ;
        RECT 59.210 204.550 59.560 204.880 ;
        RECT 59.740 204.550 60.105 205.230 ;
        RECT 59.390 204.380 59.560 204.550 ;
        RECT 59.390 204.210 60.020 204.380 ;
        RECT 58.870 203.810 59.100 204.140 ;
        RECT 59.345 203.640 59.675 204.020 ;
        RECT 59.845 203.810 60.020 204.210 ;
        RECT 61.195 204.290 61.365 205.320 ;
        RECT 61.640 205.190 62.395 205.440 ;
        RECT 62.565 205.265 62.895 205.510 ;
        RECT 61.640 205.155 62.410 205.190 ;
        RECT 61.640 205.145 62.425 205.155 ;
        RECT 61.535 205.130 62.430 205.145 ;
        RECT 61.535 205.115 62.450 205.130 ;
        RECT 61.535 205.105 62.470 205.115 ;
        RECT 61.535 205.095 62.495 205.105 ;
        RECT 61.535 205.065 62.565 205.095 ;
        RECT 61.535 205.035 62.585 205.065 ;
        RECT 61.535 205.005 62.605 205.035 ;
        RECT 61.535 204.980 62.635 205.005 ;
        RECT 61.535 204.945 62.670 204.980 ;
        RECT 61.535 204.940 62.700 204.945 ;
        RECT 61.535 204.545 61.765 204.940 ;
        RECT 62.310 204.935 62.700 204.940 ;
        RECT 62.335 204.925 62.700 204.935 ;
        RECT 62.350 204.920 62.700 204.925 ;
        RECT 62.365 204.915 62.700 204.920 ;
        RECT 63.065 204.915 63.325 205.365 ;
        RECT 62.365 204.910 63.325 204.915 ;
        RECT 62.375 204.900 63.325 204.910 ;
        RECT 62.385 204.895 63.325 204.900 ;
        RECT 62.395 204.885 63.325 204.895 ;
        RECT 62.400 204.875 63.325 204.885 ;
        RECT 62.405 204.870 63.325 204.875 ;
        RECT 62.415 204.855 63.325 204.870 ;
        RECT 62.420 204.840 63.325 204.855 ;
        RECT 62.430 204.815 63.325 204.840 ;
        RECT 61.935 204.345 62.265 204.770 ;
        RECT 61.195 203.810 61.455 204.290 ;
        RECT 61.625 203.640 61.875 204.180 ;
        RECT 62.045 203.860 62.265 204.345 ;
        RECT 62.435 204.745 63.325 204.815 ;
        RECT 63.495 205.310 64.155 205.510 ;
        RECT 64.325 205.340 66.545 205.510 ;
        RECT 62.435 204.020 62.605 204.745 ;
        RECT 62.775 204.190 63.325 204.575 ;
        RECT 63.495 204.380 63.665 205.310 ;
        RECT 64.325 205.140 64.495 205.340 ;
        RECT 63.835 204.970 64.495 205.140 ;
        RECT 64.665 205.000 66.205 205.170 ;
        RECT 63.835 204.550 64.005 204.970 ;
        RECT 64.665 204.800 64.835 205.000 ;
        RECT 64.235 204.630 64.835 204.800 ;
        RECT 65.005 204.630 65.700 204.830 ;
        RECT 65.960 204.550 66.205 205.000 ;
        RECT 64.325 204.380 65.235 204.460 ;
        RECT 62.435 203.850 63.325 204.020 ;
        RECT 63.495 203.900 63.815 204.380 ;
        RECT 63.985 204.290 65.235 204.380 ;
        RECT 63.985 204.210 64.495 204.290 ;
        RECT 63.985 203.810 64.215 204.210 ;
        RECT 64.385 203.640 64.735 204.030 ;
        RECT 64.905 203.810 65.235 204.290 ;
        RECT 65.405 203.640 65.575 204.460 ;
        RECT 66.375 204.380 66.545 205.340 ;
        RECT 66.715 205.025 67.005 206.190 ;
        RECT 67.175 205.050 67.435 206.190 ;
        RECT 67.605 205.040 67.935 206.020 ;
        RECT 68.105 205.050 68.385 206.190 ;
        RECT 69.515 205.050 69.745 206.190 ;
        RECT 69.915 205.040 70.245 206.020 ;
        RECT 70.415 205.050 70.625 206.190 ;
        RECT 71.315 205.100 72.985 206.190 ;
        RECT 73.160 205.755 78.505 206.190 ;
        RECT 78.680 205.755 84.025 206.190 ;
        RECT 67.695 205.000 67.870 205.040 ;
        RECT 67.195 204.630 67.530 204.880 ;
        RECT 67.700 204.440 67.870 205.000 ;
        RECT 68.040 204.610 68.375 204.880 ;
        RECT 69.495 204.630 69.825 204.880 ;
        RECT 66.080 203.835 66.545 204.380 ;
        RECT 66.715 203.640 67.005 204.365 ;
        RECT 67.175 203.810 67.870 204.440 ;
        RECT 68.075 203.640 68.385 204.440 ;
        RECT 69.515 203.640 69.745 204.460 ;
        RECT 69.995 204.440 70.245 205.040 ;
        RECT 71.315 204.580 72.065 205.100 ;
        RECT 69.915 203.810 70.245 204.440 ;
        RECT 70.415 203.640 70.625 204.460 ;
        RECT 72.235 204.410 72.985 204.930 ;
        RECT 74.750 204.505 75.100 205.755 ;
        RECT 71.315 203.640 72.985 204.410 ;
        RECT 76.580 204.185 76.920 205.015 ;
        RECT 80.270 204.505 80.620 205.755 ;
        RECT 84.285 205.260 84.455 206.020 ;
        RECT 84.635 205.430 84.965 206.190 ;
        RECT 84.285 205.090 84.950 205.260 ;
        RECT 85.135 205.115 85.405 206.020 ;
        RECT 85.580 205.755 90.925 206.190 ;
        RECT 82.100 204.185 82.440 205.015 ;
        RECT 84.780 204.945 84.950 205.090 ;
        RECT 84.215 204.540 84.545 204.910 ;
        RECT 84.780 204.615 85.065 204.945 ;
        RECT 84.780 204.360 84.950 204.615 ;
        RECT 84.285 204.190 84.950 204.360 ;
        RECT 85.235 204.315 85.405 205.115 ;
        RECT 87.170 204.505 87.520 205.755 ;
        RECT 91.135 205.050 91.365 206.190 ;
        RECT 91.535 205.040 91.865 206.020 ;
        RECT 92.035 205.050 92.245 206.190 ;
        RECT 73.160 203.640 78.505 204.185 ;
        RECT 78.680 203.640 84.025 204.185 ;
        RECT 84.285 203.810 84.455 204.190 ;
        RECT 84.635 203.640 84.965 204.020 ;
        RECT 85.145 203.810 85.405 204.315 ;
        RECT 89.000 204.185 89.340 205.015 ;
        RECT 91.115 204.630 91.445 204.880 ;
        RECT 85.580 203.640 90.925 204.185 ;
        RECT 91.135 203.640 91.365 204.460 ;
        RECT 91.615 204.440 91.865 205.040 ;
        RECT 92.475 205.025 92.765 206.190 ;
        RECT 92.940 205.000 93.195 205.880 ;
        RECT 93.365 205.050 93.670 206.190 ;
        RECT 94.010 205.810 94.340 206.190 ;
        RECT 94.520 205.640 94.690 205.930 ;
        RECT 94.860 205.730 95.110 206.190 ;
        RECT 93.890 205.470 94.690 205.640 ;
        RECT 95.280 205.680 96.150 206.020 ;
        RECT 91.535 203.810 91.865 204.440 ;
        RECT 92.035 203.640 92.245 204.460 ;
        RECT 92.475 203.640 92.765 204.365 ;
        RECT 92.940 204.350 93.150 205.000 ;
        RECT 93.890 204.880 94.060 205.470 ;
        RECT 95.280 205.300 95.450 205.680 ;
        RECT 96.385 205.560 96.555 206.020 ;
        RECT 96.725 205.730 97.095 206.190 ;
        RECT 97.390 205.590 97.560 205.930 ;
        RECT 97.730 205.760 98.060 206.190 ;
        RECT 98.295 205.590 98.465 205.930 ;
        RECT 94.230 205.130 95.450 205.300 ;
        RECT 95.620 205.220 96.080 205.510 ;
        RECT 96.385 205.390 96.945 205.560 ;
        RECT 97.390 205.420 98.465 205.590 ;
        RECT 98.635 205.690 99.315 206.020 ;
        RECT 99.530 205.690 99.780 206.020 ;
        RECT 99.950 205.730 100.200 206.190 ;
        RECT 96.775 205.250 96.945 205.390 ;
        RECT 95.620 205.210 96.585 205.220 ;
        RECT 95.280 205.040 95.450 205.130 ;
        RECT 95.910 205.050 96.585 205.210 ;
        RECT 93.320 204.850 94.060 204.880 ;
        RECT 93.320 204.550 94.235 204.850 ;
        RECT 93.910 204.375 94.235 204.550 ;
        RECT 92.940 203.820 93.195 204.350 ;
        RECT 93.365 203.640 93.670 204.100 ;
        RECT 93.915 204.020 94.235 204.375 ;
        RECT 94.405 204.590 94.945 204.960 ;
        RECT 95.280 204.870 95.685 205.040 ;
        RECT 94.405 204.190 94.645 204.590 ;
        RECT 95.125 204.420 95.345 204.700 ;
        RECT 94.815 204.250 95.345 204.420 ;
        RECT 94.815 204.020 94.985 204.250 ;
        RECT 95.515 204.090 95.685 204.870 ;
        RECT 95.855 204.260 96.205 204.880 ;
        RECT 96.375 204.260 96.585 205.050 ;
        RECT 96.775 205.080 98.275 205.250 ;
        RECT 96.775 204.390 96.945 205.080 ;
        RECT 98.635 204.910 98.805 205.690 ;
        RECT 99.610 205.560 99.780 205.690 ;
        RECT 97.115 204.740 98.805 204.910 ;
        RECT 98.975 205.130 99.440 205.520 ;
        RECT 99.610 205.390 100.005 205.560 ;
        RECT 97.115 204.560 97.285 204.740 ;
        RECT 93.915 203.850 94.985 204.020 ;
        RECT 95.155 203.640 95.345 204.080 ;
        RECT 95.515 203.810 96.465 204.090 ;
        RECT 96.775 204.000 97.035 204.390 ;
        RECT 97.455 204.320 98.245 204.570 ;
        RECT 96.685 203.830 97.035 204.000 ;
        RECT 97.245 203.640 97.575 204.100 ;
        RECT 98.450 204.030 98.620 204.740 ;
        RECT 98.975 204.540 99.145 205.130 ;
        RECT 98.790 204.320 99.145 204.540 ;
        RECT 99.315 204.320 99.665 204.940 ;
        RECT 99.835 204.030 100.005 205.390 ;
        RECT 100.370 205.220 100.695 206.005 ;
        RECT 100.175 204.170 100.635 205.220 ;
        RECT 98.450 203.860 99.305 204.030 ;
        RECT 99.510 203.860 100.005 204.030 ;
        RECT 100.175 203.640 100.505 204.000 ;
        RECT 100.865 203.900 101.035 206.020 ;
        RECT 101.205 205.690 101.535 206.190 ;
        RECT 101.705 205.520 101.960 206.020 ;
        RECT 101.210 205.350 101.960 205.520 ;
        RECT 101.210 204.360 101.440 205.350 ;
        RECT 101.610 204.530 101.960 205.180 ;
        RECT 102.595 205.100 106.105 206.190 ;
        RECT 106.280 205.755 111.625 206.190 ;
        RECT 111.800 205.755 117.145 206.190 ;
        RECT 102.595 204.580 104.285 205.100 ;
        RECT 104.455 204.410 106.105 204.930 ;
        RECT 107.870 204.505 108.220 205.755 ;
        RECT 101.210 204.190 101.960 204.360 ;
        RECT 101.205 203.640 101.535 204.020 ;
        RECT 101.705 203.900 101.960 204.190 ;
        RECT 102.595 203.640 106.105 204.410 ;
        RECT 109.700 204.185 110.040 205.015 ;
        RECT 113.390 204.505 113.740 205.755 ;
        RECT 117.315 205.100 118.525 206.190 ;
        RECT 115.220 204.185 115.560 205.015 ;
        RECT 117.315 204.560 117.835 205.100 ;
        RECT 118.005 204.390 118.525 204.930 ;
        RECT 106.280 203.640 111.625 204.185 ;
        RECT 111.800 203.640 117.145 204.185 ;
        RECT 117.315 203.640 118.525 204.390 ;
        RECT 11.430 203.470 118.610 203.640 ;
        RECT 11.515 202.720 12.725 203.470 ;
        RECT 11.515 202.180 12.035 202.720 ;
        RECT 13.355 202.700 16.865 203.470 ;
        RECT 17.040 202.925 22.385 203.470 ;
        RECT 22.560 202.925 27.905 203.470 ;
        RECT 12.205 202.010 12.725 202.550 ;
        RECT 11.515 200.920 12.725 202.010 ;
        RECT 13.355 202.010 15.045 202.530 ;
        RECT 15.215 202.180 16.865 202.700 ;
        RECT 13.355 200.920 16.865 202.010 ;
        RECT 18.630 201.355 18.980 202.605 ;
        RECT 20.460 202.095 20.800 202.925 ;
        RECT 24.150 201.355 24.500 202.605 ;
        RECT 25.980 202.095 26.320 202.925 ;
        RECT 28.075 202.745 28.365 203.470 ;
        RECT 28.995 202.700 31.585 203.470 ;
        RECT 31.760 202.925 37.105 203.470 ;
        RECT 37.280 202.925 42.625 203.470 ;
        RECT 42.800 202.925 48.145 203.470 ;
        RECT 48.320 202.925 53.665 203.470 ;
        RECT 17.040 200.920 22.385 201.355 ;
        RECT 22.560 200.920 27.905 201.355 ;
        RECT 28.075 200.920 28.365 202.085 ;
        RECT 28.995 202.010 30.205 202.530 ;
        RECT 30.375 202.180 31.585 202.700 ;
        RECT 28.995 200.920 31.585 202.010 ;
        RECT 33.350 201.355 33.700 202.605 ;
        RECT 35.180 202.095 35.520 202.925 ;
        RECT 38.870 201.355 39.220 202.605 ;
        RECT 40.700 202.095 41.040 202.925 ;
        RECT 44.390 201.355 44.740 202.605 ;
        RECT 46.220 202.095 46.560 202.925 ;
        RECT 49.910 201.355 50.260 202.605 ;
        RECT 51.740 202.095 52.080 202.925 ;
        RECT 53.835 202.745 54.125 203.470 ;
        RECT 54.295 202.720 55.505 203.470 ;
        RECT 31.760 200.920 37.105 201.355 ;
        RECT 37.280 200.920 42.625 201.355 ;
        RECT 42.800 200.920 48.145 201.355 ;
        RECT 48.320 200.920 53.665 201.355 ;
        RECT 53.835 200.920 54.125 202.085 ;
        RECT 54.295 202.010 54.815 202.550 ;
        RECT 54.985 202.180 55.505 202.720 ;
        RECT 55.675 202.970 55.935 203.300 ;
        RECT 56.145 202.990 56.420 203.470 ;
        RECT 55.675 202.060 55.845 202.970 ;
        RECT 56.630 202.900 56.835 203.300 ;
        RECT 57.005 203.070 57.340 203.470 ;
        RECT 57.515 202.970 57.775 203.300 ;
        RECT 58.085 203.090 58.415 203.470 ;
        RECT 58.595 203.130 60.075 203.300 ;
        RECT 56.015 202.230 56.375 202.810 ;
        RECT 56.630 202.730 57.315 202.900 ;
        RECT 56.555 202.060 56.805 202.560 ;
        RECT 54.295 200.920 55.505 202.010 ;
        RECT 55.675 201.890 56.805 202.060 ;
        RECT 55.675 201.120 55.945 201.890 ;
        RECT 56.975 201.700 57.315 202.730 ;
        RECT 56.115 200.920 56.445 201.700 ;
        RECT 56.650 201.525 57.315 201.700 ;
        RECT 57.515 202.270 57.685 202.970 ;
        RECT 58.595 202.800 58.995 203.130 ;
        RECT 58.035 202.610 58.245 202.790 ;
        RECT 58.035 202.440 58.655 202.610 ;
        RECT 58.825 202.320 58.995 202.800 ;
        RECT 59.185 202.630 59.735 202.960 ;
        RECT 57.515 202.100 58.645 202.270 ;
        RECT 58.825 202.150 59.395 202.320 ;
        RECT 56.650 201.120 56.835 201.525 ;
        RECT 57.515 201.420 57.685 202.100 ;
        RECT 58.475 201.980 58.645 202.100 ;
        RECT 57.855 201.600 58.205 201.930 ;
        RECT 58.475 201.810 59.055 201.980 ;
        RECT 59.225 201.640 59.395 202.150 ;
        RECT 58.655 201.470 59.395 201.640 ;
        RECT 59.565 201.640 59.735 202.630 ;
        RECT 59.905 202.230 60.075 203.130 ;
        RECT 60.325 202.560 60.510 203.140 ;
        RECT 60.780 202.560 60.975 203.135 ;
        RECT 61.185 203.090 61.515 203.470 ;
        RECT 60.325 202.230 60.555 202.560 ;
        RECT 60.780 202.230 61.035 202.560 ;
        RECT 60.325 201.920 60.510 202.230 ;
        RECT 60.780 201.920 60.975 202.230 ;
        RECT 61.345 201.640 61.515 202.560 ;
        RECT 59.565 201.470 61.515 201.640 ;
        RECT 57.005 200.920 57.340 201.345 ;
        RECT 57.515 201.090 57.775 201.420 ;
        RECT 58.085 200.920 58.415 201.300 ;
        RECT 58.655 201.090 58.845 201.470 ;
        RECT 59.095 200.920 59.425 201.300 ;
        RECT 59.635 201.090 59.805 201.470 ;
        RECT 60.000 200.920 60.330 201.300 ;
        RECT 60.590 201.090 60.760 201.470 ;
        RECT 61.185 200.920 61.515 201.300 ;
        RECT 61.685 201.090 61.945 203.300 ;
        RECT 62.575 202.795 62.835 203.300 ;
        RECT 63.015 203.090 63.345 203.470 ;
        RECT 63.525 202.920 63.695 203.300 ;
        RECT 62.575 201.995 62.745 202.795 ;
        RECT 63.030 202.750 63.695 202.920 ;
        RECT 63.030 202.495 63.200 202.750 ;
        RECT 63.955 202.720 65.165 203.470 ;
        RECT 62.915 202.165 63.200 202.495 ;
        RECT 63.435 202.200 63.765 202.570 ;
        RECT 63.030 202.020 63.200 202.165 ;
        RECT 62.575 201.090 62.845 201.995 ;
        RECT 63.030 201.850 63.695 202.020 ;
        RECT 63.015 200.920 63.345 201.680 ;
        RECT 63.525 201.090 63.695 201.850 ;
        RECT 63.955 202.010 64.475 202.550 ;
        RECT 64.645 202.180 65.165 202.720 ;
        RECT 65.370 202.730 65.985 203.300 ;
        RECT 66.155 202.960 66.370 203.470 ;
        RECT 66.600 202.960 66.880 203.290 ;
        RECT 67.060 202.960 67.300 203.470 ;
        RECT 63.955 200.920 65.165 202.010 ;
        RECT 65.370 201.710 65.685 202.730 ;
        RECT 65.855 202.060 66.025 202.560 ;
        RECT 66.275 202.230 66.540 202.790 ;
        RECT 66.710 202.060 66.880 202.960 ;
        RECT 67.050 202.230 67.405 202.790 ;
        RECT 67.635 202.720 68.845 203.470 ;
        RECT 65.855 201.890 67.280 202.060 ;
        RECT 65.370 201.090 65.905 201.710 ;
        RECT 66.075 200.920 66.405 201.720 ;
        RECT 66.890 201.715 67.280 201.890 ;
        RECT 67.635 202.010 68.155 202.550 ;
        RECT 68.325 202.180 68.845 202.720 ;
        RECT 69.015 202.700 72.525 203.470 ;
        RECT 72.700 202.925 78.045 203.470 ;
        RECT 69.015 202.010 70.705 202.530 ;
        RECT 70.875 202.180 72.525 202.700 ;
        RECT 67.635 200.920 68.845 202.010 ;
        RECT 69.015 200.920 72.525 202.010 ;
        RECT 74.290 201.355 74.640 202.605 ;
        RECT 76.120 202.095 76.460 202.925 ;
        RECT 78.255 202.650 78.485 203.470 ;
        RECT 78.655 202.670 78.985 203.300 ;
        RECT 78.235 202.230 78.565 202.480 ;
        RECT 78.735 202.070 78.985 202.670 ;
        RECT 79.155 202.650 79.365 203.470 ;
        RECT 79.595 202.745 79.885 203.470 ;
        RECT 80.060 202.760 80.315 203.290 ;
        RECT 80.485 203.010 80.790 203.470 ;
        RECT 81.035 203.090 82.105 203.260 ;
        RECT 80.060 202.110 80.270 202.760 ;
        RECT 81.035 202.735 81.355 203.090 ;
        RECT 81.030 202.560 81.355 202.735 ;
        RECT 80.440 202.260 81.355 202.560 ;
        RECT 81.525 202.520 81.765 202.920 ;
        RECT 81.935 202.860 82.105 203.090 ;
        RECT 82.275 203.030 82.465 203.470 ;
        RECT 82.635 203.020 83.585 203.300 ;
        RECT 83.805 203.110 84.155 203.280 ;
        RECT 81.935 202.690 82.465 202.860 ;
        RECT 80.440 202.230 81.180 202.260 ;
        RECT 72.700 200.920 78.045 201.355 ;
        RECT 78.255 200.920 78.485 202.060 ;
        RECT 78.655 201.090 78.985 202.070 ;
        RECT 79.155 200.920 79.365 202.060 ;
        RECT 79.595 200.920 79.885 202.085 ;
        RECT 80.060 201.230 80.315 202.110 ;
        RECT 80.485 200.920 80.790 202.060 ;
        RECT 81.010 201.640 81.180 202.230 ;
        RECT 81.525 202.150 82.065 202.520 ;
        RECT 82.245 202.410 82.465 202.690 ;
        RECT 82.635 202.240 82.805 203.020 ;
        RECT 82.400 202.070 82.805 202.240 ;
        RECT 82.975 202.230 83.325 202.850 ;
        RECT 82.400 201.980 82.570 202.070 ;
        RECT 83.495 202.060 83.705 202.850 ;
        RECT 81.350 201.810 82.570 201.980 ;
        RECT 83.030 201.900 83.705 202.060 ;
        RECT 81.010 201.470 81.810 201.640 ;
        RECT 81.130 200.920 81.460 201.300 ;
        RECT 81.640 201.180 81.810 201.470 ;
        RECT 82.400 201.430 82.570 201.810 ;
        RECT 82.740 201.890 83.705 201.900 ;
        RECT 83.895 202.720 84.155 203.110 ;
        RECT 84.365 203.010 84.695 203.470 ;
        RECT 85.570 203.080 86.425 203.250 ;
        RECT 86.630 203.080 87.125 203.250 ;
        RECT 87.295 203.110 87.625 203.470 ;
        RECT 83.895 202.030 84.065 202.720 ;
        RECT 84.235 202.370 84.405 202.550 ;
        RECT 84.575 202.540 85.365 202.790 ;
        RECT 85.570 202.370 85.740 203.080 ;
        RECT 85.910 202.570 86.265 202.790 ;
        RECT 84.235 202.200 85.925 202.370 ;
        RECT 82.740 201.600 83.200 201.890 ;
        RECT 83.895 201.860 85.395 202.030 ;
        RECT 83.895 201.720 84.065 201.860 ;
        RECT 83.505 201.550 84.065 201.720 ;
        RECT 81.980 200.920 82.230 201.380 ;
        RECT 82.400 201.090 83.270 201.430 ;
        RECT 83.505 201.090 83.675 201.550 ;
        RECT 84.510 201.520 85.585 201.690 ;
        RECT 83.845 200.920 84.215 201.380 ;
        RECT 84.510 201.180 84.680 201.520 ;
        RECT 84.850 200.920 85.180 201.350 ;
        RECT 85.415 201.180 85.585 201.520 ;
        RECT 85.755 201.420 85.925 202.200 ;
        RECT 86.095 201.980 86.265 202.570 ;
        RECT 86.435 202.170 86.785 202.790 ;
        RECT 86.095 201.590 86.560 201.980 ;
        RECT 86.955 201.720 87.125 203.080 ;
        RECT 87.295 201.890 87.755 202.940 ;
        RECT 86.730 201.550 87.125 201.720 ;
        RECT 86.730 201.420 86.900 201.550 ;
        RECT 85.755 201.090 86.435 201.420 ;
        RECT 86.650 201.090 86.900 201.420 ;
        RECT 87.070 200.920 87.320 201.380 ;
        RECT 87.490 201.105 87.815 201.890 ;
        RECT 87.985 201.090 88.155 203.210 ;
        RECT 88.325 203.090 88.655 203.470 ;
        RECT 88.825 202.920 89.080 203.210 ;
        RECT 88.330 202.750 89.080 202.920 ;
        RECT 88.330 201.760 88.560 202.750 ;
        RECT 89.715 202.700 92.305 203.470 ;
        RECT 88.730 201.930 89.080 202.580 ;
        RECT 89.715 202.010 90.925 202.530 ;
        RECT 91.095 202.180 92.305 202.700 ;
        RECT 92.515 202.650 92.745 203.470 ;
        RECT 92.915 202.670 93.245 203.300 ;
        RECT 92.495 202.230 92.825 202.480 ;
        RECT 92.995 202.070 93.245 202.670 ;
        RECT 93.415 202.650 93.625 203.470 ;
        RECT 94.130 202.660 94.375 203.265 ;
        RECT 94.595 202.935 95.105 203.470 ;
        RECT 88.330 201.590 89.080 201.760 ;
        RECT 88.325 200.920 88.655 201.420 ;
        RECT 88.825 201.090 89.080 201.590 ;
        RECT 89.715 200.920 92.305 202.010 ;
        RECT 92.515 200.920 92.745 202.060 ;
        RECT 92.915 201.090 93.245 202.070 ;
        RECT 93.855 202.490 95.085 202.660 ;
        RECT 93.415 200.920 93.625 202.060 ;
        RECT 93.855 201.680 94.195 202.490 ;
        RECT 94.365 201.925 95.115 202.115 ;
        RECT 93.855 201.270 94.370 201.680 ;
        RECT 94.605 200.920 94.775 201.680 ;
        RECT 94.945 201.260 95.115 201.925 ;
        RECT 95.285 201.940 95.475 203.300 ;
        RECT 95.645 202.790 95.920 203.300 ;
        RECT 96.110 202.935 96.640 203.300 ;
        RECT 97.065 203.070 97.395 203.470 ;
        RECT 96.465 202.900 96.640 202.935 ;
        RECT 95.645 202.620 95.925 202.790 ;
        RECT 95.645 202.140 95.920 202.620 ;
        RECT 96.125 201.940 96.295 202.740 ;
        RECT 95.285 201.770 96.295 201.940 ;
        RECT 96.465 202.730 97.395 202.900 ;
        RECT 97.565 202.730 97.820 203.300 ;
        RECT 98.085 202.920 98.255 203.300 ;
        RECT 98.435 203.090 98.765 203.470 ;
        RECT 98.085 202.750 98.750 202.920 ;
        RECT 98.945 202.795 99.205 203.300 ;
        RECT 96.465 201.600 96.635 202.730 ;
        RECT 97.225 202.560 97.395 202.730 ;
        RECT 95.510 201.430 96.635 201.600 ;
        RECT 96.805 202.230 97.000 202.560 ;
        RECT 97.225 202.230 97.480 202.560 ;
        RECT 96.805 201.260 96.975 202.230 ;
        RECT 97.650 202.060 97.820 202.730 ;
        RECT 98.015 202.200 98.345 202.570 ;
        RECT 98.580 202.495 98.750 202.750 ;
        RECT 94.945 201.090 96.975 201.260 ;
        RECT 97.145 200.920 97.315 202.060 ;
        RECT 97.485 201.090 97.820 202.060 ;
        RECT 98.580 202.165 98.865 202.495 ;
        RECT 98.580 202.020 98.750 202.165 ;
        RECT 98.085 201.850 98.750 202.020 ;
        RECT 99.035 201.995 99.205 202.795 ;
        RECT 99.465 202.920 99.635 203.300 ;
        RECT 99.815 203.090 100.145 203.470 ;
        RECT 99.465 202.750 100.130 202.920 ;
        RECT 100.325 202.795 100.585 203.300 ;
        RECT 99.395 202.200 99.725 202.570 ;
        RECT 99.960 202.495 100.130 202.750 ;
        RECT 99.960 202.165 100.245 202.495 ;
        RECT 99.960 202.020 100.130 202.165 ;
        RECT 98.085 201.090 98.255 201.850 ;
        RECT 98.435 200.920 98.765 201.680 ;
        RECT 98.935 201.090 99.205 201.995 ;
        RECT 99.465 201.850 100.130 202.020 ;
        RECT 100.415 201.995 100.585 202.795 ;
        RECT 101.675 202.700 105.185 203.470 ;
        RECT 105.355 202.745 105.645 203.470 ;
        RECT 106.280 202.925 111.625 203.470 ;
        RECT 111.800 202.925 117.145 203.470 ;
        RECT 99.465 201.090 99.635 201.850 ;
        RECT 99.815 200.920 100.145 201.680 ;
        RECT 100.315 201.090 100.585 201.995 ;
        RECT 101.675 202.010 103.365 202.530 ;
        RECT 103.535 202.180 105.185 202.700 ;
        RECT 101.675 200.920 105.185 202.010 ;
        RECT 105.355 200.920 105.645 202.085 ;
        RECT 107.870 201.355 108.220 202.605 ;
        RECT 109.700 202.095 110.040 202.925 ;
        RECT 113.390 201.355 113.740 202.605 ;
        RECT 115.220 202.095 115.560 202.925 ;
        RECT 117.315 202.720 118.525 203.470 ;
        RECT 117.315 202.010 117.835 202.550 ;
        RECT 118.005 202.180 118.525 202.720 ;
        RECT 106.280 200.920 111.625 201.355 ;
        RECT 111.800 200.920 117.145 201.355 ;
        RECT 117.315 200.920 118.525 202.010 ;
        RECT 11.430 200.750 118.610 200.920 ;
        RECT 11.515 199.660 12.725 200.750 ;
        RECT 11.515 198.950 12.035 199.490 ;
        RECT 12.205 199.120 12.725 199.660 ;
        RECT 13.355 199.660 15.025 200.750 ;
        RECT 13.355 199.140 14.105 199.660 ;
        RECT 15.195 199.585 15.485 200.750 ;
        RECT 16.115 199.660 18.705 200.750 ;
        RECT 18.880 200.315 24.225 200.750 ;
        RECT 24.400 200.315 29.745 200.750 ;
        RECT 29.920 200.315 35.265 200.750 ;
        RECT 35.440 200.315 40.785 200.750 ;
        RECT 14.275 198.970 15.025 199.490 ;
        RECT 16.115 199.140 17.325 199.660 ;
        RECT 17.495 198.970 18.705 199.490 ;
        RECT 20.470 199.065 20.820 200.315 ;
        RECT 11.515 198.200 12.725 198.950 ;
        RECT 13.355 198.200 15.025 198.970 ;
        RECT 15.195 198.200 15.485 198.925 ;
        RECT 16.115 198.200 18.705 198.970 ;
        RECT 22.300 198.745 22.640 199.575 ;
        RECT 25.990 199.065 26.340 200.315 ;
        RECT 27.820 198.745 28.160 199.575 ;
        RECT 31.510 199.065 31.860 200.315 ;
        RECT 33.340 198.745 33.680 199.575 ;
        RECT 37.030 199.065 37.380 200.315 ;
        RECT 40.955 199.585 41.245 200.750 ;
        RECT 42.395 199.610 42.605 200.750 ;
        RECT 42.775 199.600 43.105 200.580 ;
        RECT 43.275 199.610 43.505 200.750 ;
        RECT 43.715 199.660 44.925 200.750 ;
        RECT 45.095 199.675 45.365 200.580 ;
        RECT 45.535 199.990 45.865 200.750 ;
        RECT 46.045 199.820 46.215 200.580 ;
        RECT 38.860 198.745 39.200 199.575 ;
        RECT 18.880 198.200 24.225 198.745 ;
        RECT 24.400 198.200 29.745 198.745 ;
        RECT 29.920 198.200 35.265 198.745 ;
        RECT 35.440 198.200 40.785 198.745 ;
        RECT 40.955 198.200 41.245 198.925 ;
        RECT 42.395 198.200 42.605 199.020 ;
        RECT 42.775 199.000 43.025 199.600 ;
        RECT 43.195 199.190 43.525 199.440 ;
        RECT 43.715 199.120 44.235 199.660 ;
        RECT 42.775 198.370 43.105 199.000 ;
        RECT 43.275 198.200 43.505 199.020 ;
        RECT 44.405 198.950 44.925 199.490 ;
        RECT 43.715 198.200 44.925 198.950 ;
        RECT 45.095 198.875 45.265 199.675 ;
        RECT 45.550 199.650 46.215 199.820 ;
        RECT 45.550 199.505 45.720 199.650 ;
        RECT 46.535 199.610 46.745 200.750 ;
        RECT 45.435 199.175 45.720 199.505 ;
        RECT 46.915 199.600 47.245 200.580 ;
        RECT 47.415 199.610 47.645 200.750 ;
        RECT 48.775 199.660 52.285 200.750 ;
        RECT 52.460 200.080 52.715 200.580 ;
        RECT 52.885 200.250 53.215 200.750 ;
        RECT 52.460 199.910 53.210 200.080 ;
        RECT 45.550 198.920 45.720 199.175 ;
        RECT 45.955 199.100 46.285 199.470 ;
        RECT 45.095 198.370 45.355 198.875 ;
        RECT 45.550 198.750 46.215 198.920 ;
        RECT 45.535 198.200 45.865 198.580 ;
        RECT 46.045 198.370 46.215 198.750 ;
        RECT 46.535 198.200 46.745 199.020 ;
        RECT 46.915 199.000 47.165 199.600 ;
        RECT 47.335 199.190 47.665 199.440 ;
        RECT 48.775 199.140 50.465 199.660 ;
        RECT 46.915 198.370 47.245 199.000 ;
        RECT 47.415 198.200 47.645 199.020 ;
        RECT 50.635 198.970 52.285 199.490 ;
        RECT 52.460 199.090 52.810 199.740 ;
        RECT 48.775 198.200 52.285 198.970 ;
        RECT 52.980 198.920 53.210 199.910 ;
        RECT 52.460 198.750 53.210 198.920 ;
        RECT 52.460 198.460 52.715 198.750 ;
        RECT 52.885 198.200 53.215 198.580 ;
        RECT 53.385 198.460 53.555 200.580 ;
        RECT 53.725 199.780 54.050 200.565 ;
        RECT 54.220 200.290 54.470 200.750 ;
        RECT 54.640 200.250 54.890 200.580 ;
        RECT 55.105 200.250 55.785 200.580 ;
        RECT 54.640 200.120 54.810 200.250 ;
        RECT 54.415 199.950 54.810 200.120 ;
        RECT 53.785 198.730 54.245 199.780 ;
        RECT 54.415 198.590 54.585 199.950 ;
        RECT 54.980 199.690 55.445 200.080 ;
        RECT 54.755 198.880 55.105 199.500 ;
        RECT 55.275 199.100 55.445 199.690 ;
        RECT 55.615 199.470 55.785 200.250 ;
        RECT 55.955 200.150 56.125 200.490 ;
        RECT 56.360 200.320 56.690 200.750 ;
        RECT 56.860 200.150 57.030 200.490 ;
        RECT 57.325 200.290 57.695 200.750 ;
        RECT 55.955 199.980 57.030 200.150 ;
        RECT 57.865 200.120 58.035 200.580 ;
        RECT 58.270 200.240 59.140 200.580 ;
        RECT 59.310 200.290 59.560 200.750 ;
        RECT 57.475 199.950 58.035 200.120 ;
        RECT 57.475 199.810 57.645 199.950 ;
        RECT 56.145 199.640 57.645 199.810 ;
        RECT 58.340 199.780 58.800 200.070 ;
        RECT 55.615 199.300 57.305 199.470 ;
        RECT 55.275 198.880 55.630 199.100 ;
        RECT 55.800 198.590 55.970 199.300 ;
        RECT 56.175 198.880 56.965 199.130 ;
        RECT 57.135 199.120 57.305 199.300 ;
        RECT 57.475 198.950 57.645 199.640 ;
        RECT 53.915 198.200 54.245 198.560 ;
        RECT 54.415 198.420 54.910 198.590 ;
        RECT 55.115 198.420 55.970 198.590 ;
        RECT 56.845 198.200 57.175 198.660 ;
        RECT 57.385 198.560 57.645 198.950 ;
        RECT 57.835 199.770 58.800 199.780 ;
        RECT 58.970 199.860 59.140 200.240 ;
        RECT 59.730 200.200 59.900 200.490 ;
        RECT 60.080 200.370 60.410 200.750 ;
        RECT 59.730 200.030 60.530 200.200 ;
        RECT 57.835 199.610 58.510 199.770 ;
        RECT 58.970 199.690 60.190 199.860 ;
        RECT 57.835 198.820 58.045 199.610 ;
        RECT 58.970 199.600 59.140 199.690 ;
        RECT 58.215 198.820 58.565 199.440 ;
        RECT 58.735 199.430 59.140 199.600 ;
        RECT 58.735 198.650 58.905 199.430 ;
        RECT 59.075 198.980 59.295 199.260 ;
        RECT 59.475 199.150 60.015 199.520 ;
        RECT 60.360 199.410 60.530 200.030 ;
        RECT 60.705 199.690 60.875 200.750 ;
        RECT 61.085 199.740 61.375 200.580 ;
        RECT 61.545 199.910 61.715 200.750 ;
        RECT 61.925 199.740 62.175 200.580 ;
        RECT 62.385 199.910 62.555 200.750 ;
        RECT 61.085 199.570 62.810 199.740 ;
        RECT 59.075 198.810 59.605 198.980 ;
        RECT 57.385 198.390 57.735 198.560 ;
        RECT 57.955 198.370 58.905 198.650 ;
        RECT 59.075 198.200 59.265 198.640 ;
        RECT 59.435 198.580 59.605 198.810 ;
        RECT 59.775 198.750 60.015 199.150 ;
        RECT 60.185 199.400 60.530 199.410 ;
        RECT 60.185 199.190 62.215 199.400 ;
        RECT 60.185 198.935 60.510 199.190 ;
        RECT 62.400 199.020 62.810 199.570 ;
        RECT 63.035 199.660 66.545 200.750 ;
        RECT 63.035 199.140 64.725 199.660 ;
        RECT 66.715 199.585 67.005 200.750 ;
        RECT 67.175 199.660 69.765 200.750 ;
        RECT 69.940 200.315 75.285 200.750 ;
        RECT 60.185 198.580 60.505 198.935 ;
        RECT 59.435 198.410 60.505 198.580 ;
        RECT 60.705 198.200 60.875 199.010 ;
        RECT 61.045 198.850 62.810 199.020 ;
        RECT 64.895 198.970 66.545 199.490 ;
        RECT 67.175 199.140 68.385 199.660 ;
        RECT 68.555 198.970 69.765 199.490 ;
        RECT 71.530 199.065 71.880 200.315 ;
        RECT 75.830 199.770 76.085 200.440 ;
        RECT 76.265 199.950 76.550 200.750 ;
        RECT 76.730 200.030 77.060 200.540 ;
        RECT 61.045 198.370 61.375 198.850 ;
        RECT 61.545 198.200 61.715 198.670 ;
        RECT 61.885 198.370 62.215 198.850 ;
        RECT 62.385 198.200 62.555 198.670 ;
        RECT 63.035 198.200 66.545 198.970 ;
        RECT 66.715 198.200 67.005 198.925 ;
        RECT 67.175 198.200 69.765 198.970 ;
        RECT 73.360 198.745 73.700 199.575 ;
        RECT 75.830 198.910 76.010 199.770 ;
        RECT 76.730 199.440 76.980 200.030 ;
        RECT 77.330 199.880 77.500 200.490 ;
        RECT 77.670 200.060 78.000 200.750 ;
        RECT 78.230 200.200 78.470 200.490 ;
        RECT 78.670 200.370 79.090 200.750 ;
        RECT 79.270 200.280 79.900 200.530 ;
        RECT 80.370 200.370 80.700 200.750 ;
        RECT 79.270 200.200 79.440 200.280 ;
        RECT 80.870 200.200 81.040 200.490 ;
        RECT 81.220 200.370 81.600 200.750 ;
        RECT 81.840 200.365 82.670 200.535 ;
        RECT 78.230 200.030 79.440 200.200 ;
        RECT 76.180 199.110 76.980 199.440 ;
        RECT 69.940 198.200 75.285 198.745 ;
        RECT 75.830 198.710 76.085 198.910 ;
        RECT 75.745 198.540 76.085 198.710 ;
        RECT 75.830 198.380 76.085 198.540 ;
        RECT 76.265 198.200 76.550 198.660 ;
        RECT 76.730 198.460 76.980 199.110 ;
        RECT 77.180 199.860 77.500 199.880 ;
        RECT 77.180 199.690 79.100 199.860 ;
        RECT 77.180 198.795 77.370 199.690 ;
        RECT 79.270 199.520 79.440 200.030 ;
        RECT 79.610 199.770 80.130 200.080 ;
        RECT 77.540 199.350 79.440 199.520 ;
        RECT 77.540 199.290 77.870 199.350 ;
        RECT 78.020 199.120 78.350 199.180 ;
        RECT 77.690 198.850 78.350 199.120 ;
        RECT 77.180 198.465 77.500 198.795 ;
        RECT 77.680 198.200 78.340 198.680 ;
        RECT 78.540 198.590 78.710 199.350 ;
        RECT 79.610 199.180 79.790 199.590 ;
        RECT 78.880 199.010 79.210 199.130 ;
        RECT 79.960 199.010 80.130 199.770 ;
        RECT 78.880 198.840 80.130 199.010 ;
        RECT 80.300 199.950 81.670 200.200 ;
        RECT 80.300 199.180 80.490 199.950 ;
        RECT 81.420 199.690 81.670 199.950 ;
        RECT 80.660 199.520 80.910 199.680 ;
        RECT 81.840 199.520 82.010 200.365 ;
        RECT 82.905 200.080 83.075 200.580 ;
        RECT 83.245 200.250 83.575 200.750 ;
        RECT 82.180 199.690 82.680 200.070 ;
        RECT 82.905 199.910 83.600 200.080 ;
        RECT 80.660 199.350 82.010 199.520 ;
        RECT 81.590 199.310 82.010 199.350 ;
        RECT 80.300 198.840 80.720 199.180 ;
        RECT 81.010 198.850 81.420 199.180 ;
        RECT 78.540 198.420 79.390 198.590 ;
        RECT 79.950 198.200 80.270 198.660 ;
        RECT 80.470 198.410 80.720 198.840 ;
        RECT 81.010 198.200 81.420 198.640 ;
        RECT 81.590 198.580 81.760 199.310 ;
        RECT 81.930 198.760 82.280 199.130 ;
        RECT 82.460 198.820 82.680 199.690 ;
        RECT 82.850 199.120 83.260 199.740 ;
        RECT 83.430 198.940 83.600 199.910 ;
        RECT 82.905 198.750 83.600 198.940 ;
        RECT 81.590 198.380 82.605 198.580 ;
        RECT 82.905 198.420 83.075 198.750 ;
        RECT 83.245 198.200 83.575 198.580 ;
        RECT 83.790 198.460 84.015 200.580 ;
        RECT 84.185 200.250 84.515 200.750 ;
        RECT 84.685 200.080 84.855 200.580 ;
        RECT 84.190 199.910 84.855 200.080 ;
        RECT 84.190 198.920 84.420 199.910 ;
        RECT 84.590 199.090 84.940 199.740 ;
        RECT 85.115 199.660 86.785 200.750 ;
        RECT 86.960 200.315 92.305 200.750 ;
        RECT 85.115 199.140 85.865 199.660 ;
        RECT 86.035 198.970 86.785 199.490 ;
        RECT 88.550 199.065 88.900 200.315 ;
        RECT 92.475 199.585 92.765 200.750 ;
        RECT 92.935 199.660 94.605 200.750 ;
        RECT 94.775 199.990 95.290 200.400 ;
        RECT 95.525 199.990 95.695 200.750 ;
        RECT 95.865 200.410 97.895 200.580 ;
        RECT 84.190 198.750 84.855 198.920 ;
        RECT 84.185 198.200 84.515 198.580 ;
        RECT 84.685 198.460 84.855 198.750 ;
        RECT 85.115 198.200 86.785 198.970 ;
        RECT 90.380 198.745 90.720 199.575 ;
        RECT 92.935 199.140 93.685 199.660 ;
        RECT 93.855 198.970 94.605 199.490 ;
        RECT 94.775 199.180 95.115 199.990 ;
        RECT 95.865 199.745 96.035 200.410 ;
        RECT 96.430 200.070 97.555 200.240 ;
        RECT 95.285 199.555 96.035 199.745 ;
        RECT 96.205 199.730 97.215 199.900 ;
        RECT 94.775 199.010 96.005 199.180 ;
        RECT 86.960 198.200 92.305 198.745 ;
        RECT 92.475 198.200 92.765 198.925 ;
        RECT 92.935 198.200 94.605 198.970 ;
        RECT 95.050 198.405 95.295 199.010 ;
        RECT 95.515 198.200 96.025 198.735 ;
        RECT 96.205 198.370 96.395 199.730 ;
        RECT 96.565 198.710 96.840 199.530 ;
        RECT 97.045 198.930 97.215 199.730 ;
        RECT 97.385 198.940 97.555 200.070 ;
        RECT 97.725 199.440 97.895 200.410 ;
        RECT 98.065 199.610 98.235 200.750 ;
        RECT 98.405 199.610 98.740 200.580 ;
        RECT 97.725 199.110 97.920 199.440 ;
        RECT 98.145 199.110 98.400 199.440 ;
        RECT 98.145 198.940 98.315 199.110 ;
        RECT 98.570 198.940 98.740 199.610 ;
        RECT 98.915 199.660 100.585 200.750 ;
        RECT 100.845 199.820 101.015 200.580 ;
        RECT 101.195 199.990 101.525 200.750 ;
        RECT 98.915 199.140 99.665 199.660 ;
        RECT 100.845 199.650 101.510 199.820 ;
        RECT 101.695 199.675 101.965 200.580 ;
        RECT 101.340 199.505 101.510 199.650 ;
        RECT 99.835 198.970 100.585 199.490 ;
        RECT 100.775 199.100 101.105 199.470 ;
        RECT 101.340 199.175 101.625 199.505 ;
        RECT 97.385 198.770 98.315 198.940 ;
        RECT 97.385 198.735 97.560 198.770 ;
        RECT 96.565 198.540 96.845 198.710 ;
        RECT 96.565 198.370 96.840 198.540 ;
        RECT 97.030 198.370 97.560 198.735 ;
        RECT 97.985 198.200 98.315 198.600 ;
        RECT 98.485 198.370 98.740 198.940 ;
        RECT 98.915 198.200 100.585 198.970 ;
        RECT 101.340 198.920 101.510 199.175 ;
        RECT 100.845 198.750 101.510 198.920 ;
        RECT 101.795 198.875 101.965 199.675 ;
        RECT 102.595 199.660 106.105 200.750 ;
        RECT 106.280 200.315 111.625 200.750 ;
        RECT 111.800 200.315 117.145 200.750 ;
        RECT 102.595 199.140 104.285 199.660 ;
        RECT 104.455 198.970 106.105 199.490 ;
        RECT 107.870 199.065 108.220 200.315 ;
        RECT 100.845 198.370 101.015 198.750 ;
        RECT 101.195 198.200 101.525 198.580 ;
        RECT 101.705 198.370 101.965 198.875 ;
        RECT 102.595 198.200 106.105 198.970 ;
        RECT 109.700 198.745 110.040 199.575 ;
        RECT 113.390 199.065 113.740 200.315 ;
        RECT 117.315 199.660 118.525 200.750 ;
        RECT 115.220 198.745 115.560 199.575 ;
        RECT 117.315 199.120 117.835 199.660 ;
        RECT 118.005 198.950 118.525 199.490 ;
        RECT 106.280 198.200 111.625 198.745 ;
        RECT 111.800 198.200 117.145 198.745 ;
        RECT 117.315 198.200 118.525 198.950 ;
        RECT 11.430 198.030 118.610 198.200 ;
        RECT 11.515 197.280 12.725 198.030 ;
        RECT 11.515 196.740 12.035 197.280 ;
        RECT 13.355 197.260 16.865 198.030 ;
        RECT 17.040 197.485 22.385 198.030 ;
        RECT 22.560 197.485 27.905 198.030 ;
        RECT 12.205 196.570 12.725 197.110 ;
        RECT 11.515 195.480 12.725 196.570 ;
        RECT 13.355 196.570 15.045 197.090 ;
        RECT 15.215 196.740 16.865 197.260 ;
        RECT 13.355 195.480 16.865 196.570 ;
        RECT 18.630 195.915 18.980 197.165 ;
        RECT 20.460 196.655 20.800 197.485 ;
        RECT 24.150 195.915 24.500 197.165 ;
        RECT 25.980 196.655 26.320 197.485 ;
        RECT 28.075 197.305 28.365 198.030 ;
        RECT 29.455 197.260 32.965 198.030 ;
        RECT 33.225 197.480 33.395 197.770 ;
        RECT 33.565 197.650 33.895 198.030 ;
        RECT 33.225 197.310 33.890 197.480 ;
        RECT 17.040 195.480 22.385 195.915 ;
        RECT 22.560 195.480 27.905 195.915 ;
        RECT 28.075 195.480 28.365 196.645 ;
        RECT 29.455 196.570 31.145 197.090 ;
        RECT 31.315 196.740 32.965 197.260 ;
        RECT 29.455 195.480 32.965 196.570 ;
        RECT 33.140 196.490 33.490 197.140 ;
        RECT 33.660 196.320 33.890 197.310 ;
        RECT 33.225 196.150 33.890 196.320 ;
        RECT 33.225 195.650 33.395 196.150 ;
        RECT 33.565 195.480 33.895 195.980 ;
        RECT 34.065 195.650 34.290 197.770 ;
        RECT 34.505 197.650 34.835 198.030 ;
        RECT 35.005 197.480 35.175 197.810 ;
        RECT 35.475 197.650 36.490 197.850 ;
        RECT 34.480 197.290 35.175 197.480 ;
        RECT 34.480 196.320 34.650 197.290 ;
        RECT 34.820 196.490 35.230 197.110 ;
        RECT 35.400 196.540 35.620 197.410 ;
        RECT 35.800 197.100 36.150 197.470 ;
        RECT 36.320 196.920 36.490 197.650 ;
        RECT 36.660 197.590 37.070 198.030 ;
        RECT 37.360 197.390 37.610 197.820 ;
        RECT 37.810 197.570 38.130 198.030 ;
        RECT 38.690 197.640 39.540 197.810 ;
        RECT 36.660 197.050 37.070 197.380 ;
        RECT 37.360 197.050 37.780 197.390 ;
        RECT 36.070 196.880 36.490 196.920 ;
        RECT 36.070 196.710 37.420 196.880 ;
        RECT 34.480 196.150 35.175 196.320 ;
        RECT 35.400 196.160 35.900 196.540 ;
        RECT 34.505 195.480 34.835 195.980 ;
        RECT 35.005 195.650 35.175 196.150 ;
        RECT 36.070 195.865 36.240 196.710 ;
        RECT 37.170 196.550 37.420 196.710 ;
        RECT 36.410 196.280 36.660 196.540 ;
        RECT 37.590 196.280 37.780 197.050 ;
        RECT 36.410 196.030 37.780 196.280 ;
        RECT 37.950 197.220 39.200 197.390 ;
        RECT 37.950 196.460 38.120 197.220 ;
        RECT 38.870 197.100 39.200 197.220 ;
        RECT 38.290 196.640 38.470 197.050 ;
        RECT 39.370 196.880 39.540 197.640 ;
        RECT 39.740 197.550 40.400 198.030 ;
        RECT 40.580 197.435 40.900 197.765 ;
        RECT 39.730 197.110 40.390 197.380 ;
        RECT 39.730 197.050 40.060 197.110 ;
        RECT 40.210 196.880 40.540 196.940 ;
        RECT 38.640 196.710 40.540 196.880 ;
        RECT 37.950 196.150 38.470 196.460 ;
        RECT 38.640 196.200 38.810 196.710 ;
        RECT 40.710 196.540 40.900 197.435 ;
        RECT 38.980 196.370 40.900 196.540 ;
        RECT 40.580 196.350 40.900 196.370 ;
        RECT 41.100 197.120 41.350 197.770 ;
        RECT 41.530 197.570 41.815 198.030 ;
        RECT 41.995 197.320 42.250 197.850 ;
        RECT 41.100 196.790 41.900 197.120 ;
        RECT 38.640 196.030 39.850 196.200 ;
        RECT 35.410 195.695 36.240 195.865 ;
        RECT 36.480 195.480 36.860 195.860 ;
        RECT 37.040 195.740 37.210 196.030 ;
        RECT 38.640 195.950 38.810 196.030 ;
        RECT 37.380 195.480 37.710 195.860 ;
        RECT 38.180 195.700 38.810 195.950 ;
        RECT 38.990 195.480 39.410 195.860 ;
        RECT 39.610 195.740 39.850 196.030 ;
        RECT 40.080 195.480 40.410 196.170 ;
        RECT 40.580 195.740 40.750 196.350 ;
        RECT 41.100 196.200 41.350 196.790 ;
        RECT 42.070 196.460 42.250 197.320 ;
        RECT 41.995 196.330 42.250 196.460 ;
        RECT 43.170 197.320 43.425 197.850 ;
        RECT 43.605 197.570 43.890 198.030 ;
        RECT 43.170 196.460 43.350 197.320 ;
        RECT 44.070 197.120 44.320 197.770 ;
        RECT 43.520 196.790 44.320 197.120 ;
        RECT 41.020 195.690 41.350 196.200 ;
        RECT 41.530 195.480 41.815 196.280 ;
        RECT 41.995 196.160 42.335 196.330 ;
        RECT 41.995 195.790 42.250 196.160 ;
        RECT 43.170 195.990 43.425 196.460 ;
        RECT 43.085 195.820 43.425 195.990 ;
        RECT 43.170 195.790 43.425 195.820 ;
        RECT 43.605 195.480 43.890 196.280 ;
        RECT 44.070 196.200 44.320 196.790 ;
        RECT 44.520 197.435 44.840 197.765 ;
        RECT 45.020 197.550 45.680 198.030 ;
        RECT 45.880 197.640 46.730 197.810 ;
        RECT 44.520 196.540 44.710 197.435 ;
        RECT 45.030 197.110 45.690 197.380 ;
        RECT 45.360 197.050 45.690 197.110 ;
        RECT 44.880 196.880 45.210 196.940 ;
        RECT 45.880 196.880 46.050 197.640 ;
        RECT 47.290 197.570 47.610 198.030 ;
        RECT 47.810 197.390 48.060 197.820 ;
        RECT 48.350 197.590 48.760 198.030 ;
        RECT 48.930 197.650 49.945 197.850 ;
        RECT 46.220 197.220 47.470 197.390 ;
        RECT 46.220 197.100 46.550 197.220 ;
        RECT 44.880 196.710 46.780 196.880 ;
        RECT 44.520 196.370 46.440 196.540 ;
        RECT 44.520 196.350 44.840 196.370 ;
        RECT 44.070 195.690 44.400 196.200 ;
        RECT 44.670 195.740 44.840 196.350 ;
        RECT 46.610 196.200 46.780 196.710 ;
        RECT 46.950 196.640 47.130 197.050 ;
        RECT 47.300 196.460 47.470 197.220 ;
        RECT 45.010 195.480 45.340 196.170 ;
        RECT 45.570 196.030 46.780 196.200 ;
        RECT 46.950 196.150 47.470 196.460 ;
        RECT 47.640 197.050 48.060 197.390 ;
        RECT 48.350 197.050 48.760 197.380 ;
        RECT 47.640 196.280 47.830 197.050 ;
        RECT 48.930 196.920 49.100 197.650 ;
        RECT 50.245 197.480 50.415 197.810 ;
        RECT 50.585 197.650 50.915 198.030 ;
        RECT 49.270 197.100 49.620 197.470 ;
        RECT 48.930 196.880 49.350 196.920 ;
        RECT 48.000 196.710 49.350 196.880 ;
        RECT 48.000 196.550 48.250 196.710 ;
        RECT 48.760 196.280 49.010 196.540 ;
        RECT 47.640 196.030 49.010 196.280 ;
        RECT 45.570 195.740 45.810 196.030 ;
        RECT 46.610 195.950 46.780 196.030 ;
        RECT 46.010 195.480 46.430 195.860 ;
        RECT 46.610 195.700 47.240 195.950 ;
        RECT 47.710 195.480 48.040 195.860 ;
        RECT 48.210 195.740 48.380 196.030 ;
        RECT 49.180 195.865 49.350 196.710 ;
        RECT 49.800 196.540 50.020 197.410 ;
        RECT 50.245 197.290 50.940 197.480 ;
        RECT 49.520 196.160 50.020 196.540 ;
        RECT 50.190 196.490 50.600 197.110 ;
        RECT 50.770 196.320 50.940 197.290 ;
        RECT 50.245 196.150 50.940 196.320 ;
        RECT 48.560 195.480 48.940 195.860 ;
        RECT 49.180 195.695 50.010 195.865 ;
        RECT 50.245 195.650 50.415 196.150 ;
        RECT 50.585 195.480 50.915 195.980 ;
        RECT 51.130 195.650 51.355 197.770 ;
        RECT 51.525 197.650 51.855 198.030 ;
        RECT 52.025 197.480 52.195 197.770 ;
        RECT 51.530 197.310 52.195 197.480 ;
        RECT 51.530 196.320 51.760 197.310 ;
        RECT 52.455 197.280 53.665 198.030 ;
        RECT 53.835 197.305 54.125 198.030 ;
        RECT 51.930 196.490 52.280 197.140 ;
        RECT 52.455 196.570 52.975 197.110 ;
        RECT 53.145 196.740 53.665 197.280 ;
        RECT 54.295 197.260 56.885 198.030 ;
        RECT 51.530 196.150 52.195 196.320 ;
        RECT 51.525 195.480 51.855 195.980 ;
        RECT 52.025 195.650 52.195 196.150 ;
        RECT 52.455 195.480 53.665 196.570 ;
        RECT 53.835 195.480 54.125 196.645 ;
        RECT 54.295 196.570 55.505 197.090 ;
        RECT 55.675 196.740 56.885 197.260 ;
        RECT 57.095 197.210 57.325 198.030 ;
        RECT 57.495 197.230 57.825 197.860 ;
        RECT 57.075 196.790 57.405 197.040 ;
        RECT 57.575 196.630 57.825 197.230 ;
        RECT 57.995 197.210 58.205 198.030 ;
        RECT 58.435 197.355 58.695 197.860 ;
        RECT 58.875 197.650 59.205 198.030 ;
        RECT 59.385 197.480 59.555 197.860 ;
        RECT 60.145 197.630 60.475 198.030 ;
        RECT 54.295 195.480 56.885 196.570 ;
        RECT 57.095 195.480 57.325 196.620 ;
        RECT 57.495 195.650 57.825 196.630 ;
        RECT 57.995 195.480 58.205 196.620 ;
        RECT 58.435 196.555 58.605 197.355 ;
        RECT 58.890 197.310 59.555 197.480 ;
        RECT 60.645 197.460 60.975 197.800 ;
        RECT 62.025 197.630 62.355 198.030 ;
        RECT 58.890 197.055 59.060 197.310 ;
        RECT 59.990 197.290 62.355 197.460 ;
        RECT 62.525 197.305 62.855 197.815 ;
        RECT 58.775 196.725 59.060 197.055 ;
        RECT 59.295 196.760 59.625 197.130 ;
        RECT 58.890 196.580 59.060 196.725 ;
        RECT 58.435 195.650 58.705 196.555 ;
        RECT 58.890 196.410 59.555 196.580 ;
        RECT 58.875 195.480 59.205 196.240 ;
        RECT 59.385 195.650 59.555 196.410 ;
        RECT 59.990 196.290 60.160 197.290 ;
        RECT 62.185 197.120 62.355 197.290 ;
        RECT 60.330 196.460 60.575 197.120 ;
        RECT 60.790 196.460 61.055 197.120 ;
        RECT 61.250 196.460 61.535 197.120 ;
        RECT 61.710 196.790 62.015 197.120 ;
        RECT 62.185 196.790 62.495 197.120 ;
        RECT 61.710 196.460 61.925 196.790 ;
        RECT 59.990 196.120 60.445 196.290 ;
        RECT 60.115 195.690 60.445 196.120 ;
        RECT 60.625 196.120 61.915 196.290 ;
        RECT 60.625 195.700 60.875 196.120 ;
        RECT 61.105 195.480 61.435 195.950 ;
        RECT 61.665 195.700 61.915 196.120 ;
        RECT 62.105 195.480 62.355 196.620 ;
        RECT 62.665 196.540 62.855 197.305 ;
        RECT 62.525 195.690 62.855 196.540 ;
        RECT 63.035 197.355 63.310 197.700 ;
        RECT 63.500 197.630 63.875 198.030 ;
        RECT 64.045 197.460 64.215 197.810 ;
        RECT 64.385 197.630 64.715 198.030 ;
        RECT 64.885 197.460 65.145 197.860 ;
        RECT 63.035 196.620 63.205 197.355 ;
        RECT 63.480 197.290 65.145 197.460 ;
        RECT 63.480 197.120 63.650 197.290 ;
        RECT 65.325 197.210 65.655 197.630 ;
        RECT 65.825 197.210 66.085 198.030 ;
        RECT 66.255 197.380 66.515 197.860 ;
        RECT 66.685 197.490 66.935 198.030 ;
        RECT 65.325 197.120 65.575 197.210 ;
        RECT 63.375 196.790 63.650 197.120 ;
        RECT 63.820 196.790 64.645 197.120 ;
        RECT 64.860 196.790 65.575 197.120 ;
        RECT 65.745 196.790 66.080 197.040 ;
        RECT 63.480 196.620 63.650 196.790 ;
        RECT 63.035 195.650 63.310 196.620 ;
        RECT 63.480 196.450 64.140 196.620 ;
        RECT 64.400 196.500 64.645 196.790 ;
        RECT 63.970 196.330 64.140 196.450 ;
        RECT 64.815 196.330 65.145 196.620 ;
        RECT 63.520 195.480 63.800 196.280 ;
        RECT 63.970 196.160 65.145 196.330 ;
        RECT 65.405 196.230 65.575 196.790 ;
        RECT 63.970 195.660 65.585 195.990 ;
        RECT 65.825 195.480 66.085 196.620 ;
        RECT 66.255 196.350 66.425 197.380 ;
        RECT 67.105 197.350 67.325 197.810 ;
        RECT 67.075 197.325 67.325 197.350 ;
        RECT 66.595 196.730 66.825 197.125 ;
        RECT 66.995 196.900 67.325 197.325 ;
        RECT 67.495 197.650 68.385 197.820 ;
        RECT 67.495 196.925 67.665 197.650 ;
        RECT 68.560 197.485 73.905 198.030 ;
        RECT 67.835 197.095 68.385 197.480 ;
        RECT 67.495 196.855 68.385 196.925 ;
        RECT 67.490 196.830 68.385 196.855 ;
        RECT 67.480 196.815 68.385 196.830 ;
        RECT 67.475 196.800 68.385 196.815 ;
        RECT 67.465 196.795 68.385 196.800 ;
        RECT 67.460 196.785 68.385 196.795 ;
        RECT 67.455 196.775 68.385 196.785 ;
        RECT 67.445 196.770 68.385 196.775 ;
        RECT 67.435 196.760 68.385 196.770 ;
        RECT 67.425 196.755 68.385 196.760 ;
        RECT 67.425 196.750 67.760 196.755 ;
        RECT 67.410 196.745 67.760 196.750 ;
        RECT 67.395 196.735 67.760 196.745 ;
        RECT 67.370 196.730 67.760 196.735 ;
        RECT 66.595 196.725 67.760 196.730 ;
        RECT 66.595 196.690 67.730 196.725 ;
        RECT 66.595 196.665 67.695 196.690 ;
        RECT 66.595 196.635 67.665 196.665 ;
        RECT 66.595 196.605 67.645 196.635 ;
        RECT 66.595 196.575 67.625 196.605 ;
        RECT 66.595 196.565 67.555 196.575 ;
        RECT 66.595 196.555 67.530 196.565 ;
        RECT 66.595 196.540 67.510 196.555 ;
        RECT 66.595 196.525 67.490 196.540 ;
        RECT 66.700 196.515 67.485 196.525 ;
        RECT 66.700 196.480 67.470 196.515 ;
        RECT 66.255 195.650 66.530 196.350 ;
        RECT 66.700 196.230 67.455 196.480 ;
        RECT 67.625 196.160 67.955 196.405 ;
        RECT 68.125 196.305 68.385 196.755 ;
        RECT 67.770 196.135 67.955 196.160 ;
        RECT 67.770 196.035 68.385 196.135 ;
        RECT 66.700 195.480 66.955 196.025 ;
        RECT 67.125 195.650 67.605 195.990 ;
        RECT 67.780 195.480 68.385 196.035 ;
        RECT 70.150 195.915 70.500 197.165 ;
        RECT 71.980 196.655 72.320 197.485 ;
        RECT 74.115 197.210 74.345 198.030 ;
        RECT 74.515 197.230 74.845 197.860 ;
        RECT 74.095 196.790 74.425 197.040 ;
        RECT 74.595 196.630 74.845 197.230 ;
        RECT 75.015 197.210 75.225 198.030 ;
        RECT 75.730 197.220 75.975 197.825 ;
        RECT 76.195 197.495 76.705 198.030 ;
        RECT 68.560 195.480 73.905 195.915 ;
        RECT 74.115 195.480 74.345 196.620 ;
        RECT 74.515 195.650 74.845 196.630 ;
        RECT 75.455 197.050 76.685 197.220 ;
        RECT 75.015 195.480 75.225 196.620 ;
        RECT 75.455 196.240 75.795 197.050 ;
        RECT 75.965 196.485 76.715 196.675 ;
        RECT 75.455 195.830 75.970 196.240 ;
        RECT 76.205 195.480 76.375 196.240 ;
        RECT 76.545 195.820 76.715 196.485 ;
        RECT 76.885 196.500 77.075 197.860 ;
        RECT 77.245 197.010 77.520 197.860 ;
        RECT 77.710 197.495 78.240 197.860 ;
        RECT 78.665 197.630 78.995 198.030 ;
        RECT 78.065 197.460 78.240 197.495 ;
        RECT 77.245 196.840 77.525 197.010 ;
        RECT 77.245 196.700 77.520 196.840 ;
        RECT 77.725 196.500 77.895 197.300 ;
        RECT 76.885 196.330 77.895 196.500 ;
        RECT 78.065 197.290 78.995 197.460 ;
        RECT 79.165 197.290 79.420 197.860 ;
        RECT 79.595 197.305 79.885 198.030 ;
        RECT 78.065 196.160 78.235 197.290 ;
        RECT 78.825 197.120 78.995 197.290 ;
        RECT 77.110 195.990 78.235 196.160 ;
        RECT 78.405 196.790 78.600 197.120 ;
        RECT 78.825 196.790 79.080 197.120 ;
        RECT 78.405 195.820 78.575 196.790 ;
        RECT 79.250 196.620 79.420 197.290 ;
        RECT 80.330 197.220 80.575 197.825 ;
        RECT 80.795 197.495 81.305 198.030 ;
        RECT 80.055 197.050 81.285 197.220 ;
        RECT 76.545 195.650 78.575 195.820 ;
        RECT 78.745 195.480 78.915 196.620 ;
        RECT 79.085 195.650 79.420 196.620 ;
        RECT 79.595 195.480 79.885 196.645 ;
        RECT 80.055 196.240 80.395 197.050 ;
        RECT 80.565 196.485 81.315 196.675 ;
        RECT 80.055 195.830 80.570 196.240 ;
        RECT 80.805 195.480 80.975 196.240 ;
        RECT 81.145 195.820 81.315 196.485 ;
        RECT 81.485 196.500 81.675 197.860 ;
        RECT 81.845 197.350 82.120 197.860 ;
        RECT 82.310 197.495 82.840 197.860 ;
        RECT 83.265 197.630 83.595 198.030 ;
        RECT 82.665 197.460 82.840 197.495 ;
        RECT 81.845 197.180 82.125 197.350 ;
        RECT 81.845 196.700 82.120 197.180 ;
        RECT 82.325 196.500 82.495 197.300 ;
        RECT 81.485 196.330 82.495 196.500 ;
        RECT 82.665 197.290 83.595 197.460 ;
        RECT 83.765 197.290 84.020 197.860 ;
        RECT 82.665 196.160 82.835 197.290 ;
        RECT 83.425 197.120 83.595 197.290 ;
        RECT 81.710 195.990 82.835 196.160 ;
        RECT 83.005 196.790 83.200 197.120 ;
        RECT 83.425 196.790 83.680 197.120 ;
        RECT 83.005 195.820 83.175 196.790 ;
        RECT 83.850 196.620 84.020 197.290 ;
        RECT 81.145 195.650 83.175 195.820 ;
        RECT 83.345 195.480 83.515 196.620 ;
        RECT 83.685 195.650 84.020 196.620 ;
        RECT 84.195 197.355 84.455 197.860 ;
        RECT 84.635 197.650 84.965 198.030 ;
        RECT 85.145 197.480 85.315 197.860 ;
        RECT 84.195 196.555 84.365 197.355 ;
        RECT 84.650 197.310 85.315 197.480 ;
        RECT 84.650 197.055 84.820 197.310 ;
        RECT 85.575 197.260 88.165 198.030 ;
        RECT 88.340 197.485 93.685 198.030 ;
        RECT 84.535 196.725 84.820 197.055 ;
        RECT 85.055 196.760 85.385 197.130 ;
        RECT 84.650 196.580 84.820 196.725 ;
        RECT 84.195 195.650 84.465 196.555 ;
        RECT 84.650 196.410 85.315 196.580 ;
        RECT 84.635 195.480 84.965 196.240 ;
        RECT 85.145 195.650 85.315 196.410 ;
        RECT 85.575 196.570 86.785 197.090 ;
        RECT 86.955 196.740 88.165 197.260 ;
        RECT 85.575 195.480 88.165 196.570 ;
        RECT 89.930 195.915 90.280 197.165 ;
        RECT 91.760 196.655 92.100 197.485 ;
        RECT 93.895 197.210 94.125 198.030 ;
        RECT 94.295 197.230 94.625 197.860 ;
        RECT 93.875 196.790 94.205 197.040 ;
        RECT 94.375 196.630 94.625 197.230 ;
        RECT 94.795 197.210 95.005 198.030 ;
        RECT 95.240 197.320 95.495 197.850 ;
        RECT 95.665 197.570 95.970 198.030 ;
        RECT 96.215 197.650 97.285 197.820 ;
        RECT 88.340 195.480 93.685 195.915 ;
        RECT 93.895 195.480 94.125 196.620 ;
        RECT 94.295 195.650 94.625 196.630 ;
        RECT 95.240 196.670 95.450 197.320 ;
        RECT 96.215 197.295 96.535 197.650 ;
        RECT 96.210 197.120 96.535 197.295 ;
        RECT 95.620 196.820 96.535 197.120 ;
        RECT 96.705 197.080 96.945 197.480 ;
        RECT 97.115 197.420 97.285 197.650 ;
        RECT 97.455 197.590 97.645 198.030 ;
        RECT 97.815 197.580 98.765 197.860 ;
        RECT 98.985 197.670 99.335 197.840 ;
        RECT 97.115 197.250 97.645 197.420 ;
        RECT 95.620 196.790 96.360 196.820 ;
        RECT 94.795 195.480 95.005 196.620 ;
        RECT 95.240 195.790 95.495 196.670 ;
        RECT 95.665 195.480 95.970 196.620 ;
        RECT 96.190 196.200 96.360 196.790 ;
        RECT 96.705 196.710 97.245 197.080 ;
        RECT 97.425 196.970 97.645 197.250 ;
        RECT 97.815 196.800 97.985 197.580 ;
        RECT 97.580 196.630 97.985 196.800 ;
        RECT 98.155 196.790 98.505 197.410 ;
        RECT 97.580 196.540 97.750 196.630 ;
        RECT 98.675 196.620 98.885 197.410 ;
        RECT 96.530 196.370 97.750 196.540 ;
        RECT 98.210 196.460 98.885 196.620 ;
        RECT 96.190 196.030 96.990 196.200 ;
        RECT 96.310 195.480 96.640 195.860 ;
        RECT 96.820 195.740 96.990 196.030 ;
        RECT 97.580 195.990 97.750 196.370 ;
        RECT 97.920 196.450 98.885 196.460 ;
        RECT 99.075 197.280 99.335 197.670 ;
        RECT 99.545 197.570 99.875 198.030 ;
        RECT 100.750 197.640 101.605 197.810 ;
        RECT 101.810 197.640 102.305 197.810 ;
        RECT 102.475 197.670 102.805 198.030 ;
        RECT 99.075 196.590 99.245 197.280 ;
        RECT 99.415 196.930 99.585 197.110 ;
        RECT 99.755 197.100 100.545 197.350 ;
        RECT 100.750 196.930 100.920 197.640 ;
        RECT 101.090 197.130 101.445 197.350 ;
        RECT 99.415 196.760 101.105 196.930 ;
        RECT 97.920 196.160 98.380 196.450 ;
        RECT 99.075 196.420 100.575 196.590 ;
        RECT 99.075 196.280 99.245 196.420 ;
        RECT 98.685 196.110 99.245 196.280 ;
        RECT 97.160 195.480 97.410 195.940 ;
        RECT 97.580 195.650 98.450 195.990 ;
        RECT 98.685 195.650 98.855 196.110 ;
        RECT 99.690 196.080 100.765 196.250 ;
        RECT 99.025 195.480 99.395 195.940 ;
        RECT 99.690 195.740 99.860 196.080 ;
        RECT 100.030 195.480 100.360 195.910 ;
        RECT 100.595 195.740 100.765 196.080 ;
        RECT 100.935 195.980 101.105 196.760 ;
        RECT 101.275 196.540 101.445 197.130 ;
        RECT 101.615 196.730 101.965 197.350 ;
        RECT 101.275 196.150 101.740 196.540 ;
        RECT 102.135 196.280 102.305 197.640 ;
        RECT 102.475 196.450 102.935 197.500 ;
        RECT 101.910 196.110 102.305 196.280 ;
        RECT 101.910 195.980 102.080 196.110 ;
        RECT 100.935 195.650 101.615 195.980 ;
        RECT 101.830 195.650 102.080 195.980 ;
        RECT 102.250 195.480 102.500 195.940 ;
        RECT 102.670 195.665 102.995 196.450 ;
        RECT 103.165 195.650 103.335 197.770 ;
        RECT 103.505 197.650 103.835 198.030 ;
        RECT 104.005 197.480 104.260 197.770 ;
        RECT 103.510 197.310 104.260 197.480 ;
        RECT 103.510 196.320 103.740 197.310 ;
        RECT 105.355 197.305 105.645 198.030 ;
        RECT 106.280 197.485 111.625 198.030 ;
        RECT 111.800 197.485 117.145 198.030 ;
        RECT 103.910 196.490 104.260 197.140 ;
        RECT 103.510 196.150 104.260 196.320 ;
        RECT 103.505 195.480 103.835 195.980 ;
        RECT 104.005 195.650 104.260 196.150 ;
        RECT 105.355 195.480 105.645 196.645 ;
        RECT 107.870 195.915 108.220 197.165 ;
        RECT 109.700 196.655 110.040 197.485 ;
        RECT 113.390 195.915 113.740 197.165 ;
        RECT 115.220 196.655 115.560 197.485 ;
        RECT 117.315 197.280 118.525 198.030 ;
        RECT 117.315 196.570 117.835 197.110 ;
        RECT 118.005 196.740 118.525 197.280 ;
        RECT 106.280 195.480 111.625 195.915 ;
        RECT 111.800 195.480 117.145 195.915 ;
        RECT 117.315 195.480 118.525 196.570 ;
        RECT 11.430 195.310 118.610 195.480 ;
        RECT 11.515 194.220 12.725 195.310 ;
        RECT 11.515 193.510 12.035 194.050 ;
        RECT 12.205 193.680 12.725 194.220 ;
        RECT 13.355 194.220 15.025 195.310 ;
        RECT 13.355 193.700 14.105 194.220 ;
        RECT 15.195 194.145 15.485 195.310 ;
        RECT 15.655 194.220 16.865 195.310 ;
        RECT 17.040 194.875 22.385 195.310 ;
        RECT 22.560 194.875 27.905 195.310 ;
        RECT 14.275 193.530 15.025 194.050 ;
        RECT 15.655 193.680 16.175 194.220 ;
        RECT 11.515 192.760 12.725 193.510 ;
        RECT 13.355 192.760 15.025 193.530 ;
        RECT 16.345 193.510 16.865 194.050 ;
        RECT 18.630 193.625 18.980 194.875 ;
        RECT 15.195 192.760 15.485 193.485 ;
        RECT 15.655 192.760 16.865 193.510 ;
        RECT 20.460 193.305 20.800 194.135 ;
        RECT 24.150 193.625 24.500 194.875 ;
        RECT 25.980 193.305 26.320 194.135 ;
        RECT 28.080 194.120 28.335 195.000 ;
        RECT 28.505 194.170 28.810 195.310 ;
        RECT 29.150 194.930 29.480 195.310 ;
        RECT 29.660 194.760 29.830 195.050 ;
        RECT 30.000 194.850 30.250 195.310 ;
        RECT 29.030 194.590 29.830 194.760 ;
        RECT 30.420 194.800 31.290 195.140 ;
        RECT 28.080 193.470 28.290 194.120 ;
        RECT 29.030 194.000 29.200 194.590 ;
        RECT 30.420 194.420 30.590 194.800 ;
        RECT 31.525 194.680 31.695 195.140 ;
        RECT 31.865 194.850 32.235 195.310 ;
        RECT 32.530 194.710 32.700 195.050 ;
        RECT 32.870 194.880 33.200 195.310 ;
        RECT 33.435 194.710 33.605 195.050 ;
        RECT 29.370 194.250 30.590 194.420 ;
        RECT 30.760 194.340 31.220 194.630 ;
        RECT 31.525 194.510 32.085 194.680 ;
        RECT 32.530 194.540 33.605 194.710 ;
        RECT 33.775 194.810 34.455 195.140 ;
        RECT 34.670 194.810 34.920 195.140 ;
        RECT 35.090 194.850 35.340 195.310 ;
        RECT 31.915 194.370 32.085 194.510 ;
        RECT 30.760 194.330 31.725 194.340 ;
        RECT 30.420 194.160 30.590 194.250 ;
        RECT 31.050 194.170 31.725 194.330 ;
        RECT 28.460 193.970 29.200 194.000 ;
        RECT 28.460 193.670 29.375 193.970 ;
        RECT 29.050 193.495 29.375 193.670 ;
        RECT 17.040 192.760 22.385 193.305 ;
        RECT 22.560 192.760 27.905 193.305 ;
        RECT 28.080 192.940 28.335 193.470 ;
        RECT 28.505 192.760 28.810 193.220 ;
        RECT 29.055 193.140 29.375 193.495 ;
        RECT 29.545 193.710 30.085 194.080 ;
        RECT 30.420 193.990 30.825 194.160 ;
        RECT 29.545 193.310 29.785 193.710 ;
        RECT 30.265 193.540 30.485 193.820 ;
        RECT 29.955 193.370 30.485 193.540 ;
        RECT 29.955 193.140 30.125 193.370 ;
        RECT 30.655 193.210 30.825 193.990 ;
        RECT 30.995 193.380 31.345 194.000 ;
        RECT 31.515 193.380 31.725 194.170 ;
        RECT 31.915 194.200 33.415 194.370 ;
        RECT 31.915 193.510 32.085 194.200 ;
        RECT 33.775 194.030 33.945 194.810 ;
        RECT 34.750 194.680 34.920 194.810 ;
        RECT 32.255 193.860 33.945 194.030 ;
        RECT 34.115 194.250 34.580 194.640 ;
        RECT 34.750 194.510 35.145 194.680 ;
        RECT 32.255 193.680 32.425 193.860 ;
        RECT 29.055 192.970 30.125 193.140 ;
        RECT 30.295 192.760 30.485 193.200 ;
        RECT 30.655 192.930 31.605 193.210 ;
        RECT 31.915 193.120 32.175 193.510 ;
        RECT 32.595 193.440 33.385 193.690 ;
        RECT 31.825 192.950 32.175 193.120 ;
        RECT 32.385 192.760 32.715 193.220 ;
        RECT 33.590 193.150 33.760 193.860 ;
        RECT 34.115 193.660 34.285 194.250 ;
        RECT 33.930 193.440 34.285 193.660 ;
        RECT 34.455 193.440 34.805 194.060 ;
        RECT 34.975 193.150 35.145 194.510 ;
        RECT 35.510 194.340 35.835 195.125 ;
        RECT 35.315 193.290 35.775 194.340 ;
        RECT 33.590 192.980 34.445 193.150 ;
        RECT 34.650 192.980 35.145 193.150 ;
        RECT 35.315 192.760 35.645 193.120 ;
        RECT 36.005 193.020 36.175 195.140 ;
        RECT 36.345 194.810 36.675 195.310 ;
        RECT 36.845 194.640 37.100 195.140 ;
        RECT 36.350 194.470 37.100 194.640 ;
        RECT 36.350 193.480 36.580 194.470 ;
        RECT 36.750 193.650 37.100 194.300 ;
        RECT 37.275 194.220 38.485 195.310 ;
        RECT 38.745 194.380 38.915 195.140 ;
        RECT 39.095 194.550 39.425 195.310 ;
        RECT 37.275 193.680 37.795 194.220 ;
        RECT 38.745 194.210 39.410 194.380 ;
        RECT 39.595 194.235 39.865 195.140 ;
        RECT 39.240 194.065 39.410 194.210 ;
        RECT 37.965 193.510 38.485 194.050 ;
        RECT 38.675 193.660 39.005 194.030 ;
        RECT 39.240 193.735 39.525 194.065 ;
        RECT 36.350 193.310 37.100 193.480 ;
        RECT 36.345 192.760 36.675 193.140 ;
        RECT 36.845 193.020 37.100 193.310 ;
        RECT 37.275 192.760 38.485 193.510 ;
        RECT 39.240 193.480 39.410 193.735 ;
        RECT 38.745 193.310 39.410 193.480 ;
        RECT 39.695 193.435 39.865 194.235 ;
        RECT 40.955 194.145 41.245 195.310 ;
        RECT 42.335 194.550 42.850 194.960 ;
        RECT 43.085 194.550 43.255 195.310 ;
        RECT 43.425 194.970 45.455 195.140 ;
        RECT 42.335 193.740 42.675 194.550 ;
        RECT 43.425 194.305 43.595 194.970 ;
        RECT 43.990 194.630 45.115 194.800 ;
        RECT 42.845 194.115 43.595 194.305 ;
        RECT 43.765 194.290 44.775 194.460 ;
        RECT 42.335 193.570 43.565 193.740 ;
        RECT 38.745 192.930 38.915 193.310 ;
        RECT 39.095 192.760 39.425 193.140 ;
        RECT 39.605 192.930 39.865 193.435 ;
        RECT 40.955 192.760 41.245 193.485 ;
        RECT 42.610 192.965 42.855 193.570 ;
        RECT 43.075 192.760 43.585 193.295 ;
        RECT 43.765 192.930 43.955 194.290 ;
        RECT 44.125 193.270 44.400 194.090 ;
        RECT 44.605 193.490 44.775 194.290 ;
        RECT 44.945 193.500 45.115 194.630 ;
        RECT 45.285 194.000 45.455 194.970 ;
        RECT 45.625 194.170 45.795 195.310 ;
        RECT 45.965 194.170 46.300 195.140 ;
        RECT 45.285 193.670 45.480 194.000 ;
        RECT 45.705 193.670 45.960 194.000 ;
        RECT 45.705 193.500 45.875 193.670 ;
        RECT 46.130 193.500 46.300 194.170 ;
        RECT 46.935 194.220 48.605 195.310 ;
        RECT 48.865 194.380 49.035 195.140 ;
        RECT 49.215 194.550 49.545 195.310 ;
        RECT 46.935 193.700 47.685 194.220 ;
        RECT 48.865 194.210 49.530 194.380 ;
        RECT 49.715 194.235 49.985 195.140 ;
        RECT 49.360 194.065 49.530 194.210 ;
        RECT 47.855 193.530 48.605 194.050 ;
        RECT 48.795 193.660 49.125 194.030 ;
        RECT 49.360 193.735 49.645 194.065 ;
        RECT 44.945 193.330 45.875 193.500 ;
        RECT 44.945 193.295 45.120 193.330 ;
        RECT 44.125 193.100 44.405 193.270 ;
        RECT 44.125 192.930 44.400 193.100 ;
        RECT 44.590 192.930 45.120 193.295 ;
        RECT 45.545 192.760 45.875 193.160 ;
        RECT 46.045 192.930 46.300 193.500 ;
        RECT 46.935 192.760 48.605 193.530 ;
        RECT 49.360 193.480 49.530 193.735 ;
        RECT 48.865 193.310 49.530 193.480 ;
        RECT 49.815 193.435 49.985 194.235 ;
        RECT 50.615 194.220 54.125 195.310 ;
        RECT 54.300 194.875 59.645 195.310 ;
        RECT 50.615 193.700 52.305 194.220 ;
        RECT 52.475 193.530 54.125 194.050 ;
        RECT 55.890 193.625 56.240 194.875 ;
        RECT 59.930 194.680 60.215 195.140 ;
        RECT 60.385 194.850 60.655 195.310 ;
        RECT 59.930 194.460 60.885 194.680 ;
        RECT 48.865 192.930 49.035 193.310 ;
        RECT 49.215 192.760 49.545 193.140 ;
        RECT 49.725 192.930 49.985 193.435 ;
        RECT 50.615 192.760 54.125 193.530 ;
        RECT 57.720 193.305 58.060 194.135 ;
        RECT 59.815 193.730 60.505 194.290 ;
        RECT 60.675 193.560 60.885 194.460 ;
        RECT 59.930 193.390 60.885 193.560 ;
        RECT 61.055 194.290 61.455 195.140 ;
        RECT 61.645 194.680 61.925 195.140 ;
        RECT 62.445 194.850 62.770 195.310 ;
        RECT 61.645 194.460 62.770 194.680 ;
        RECT 61.055 193.730 62.150 194.290 ;
        RECT 62.320 194.000 62.770 194.460 ;
        RECT 62.940 194.170 63.325 195.140 ;
        RECT 54.300 192.760 59.645 193.305 ;
        RECT 59.930 192.930 60.215 193.390 ;
        RECT 60.385 192.760 60.655 193.220 ;
        RECT 61.055 192.930 61.455 193.730 ;
        RECT 62.320 193.670 62.875 194.000 ;
        RECT 62.320 193.560 62.770 193.670 ;
        RECT 61.645 193.390 62.770 193.560 ;
        RECT 63.045 193.500 63.325 194.170 ;
        RECT 61.645 192.930 61.925 193.390 ;
        RECT 62.445 192.760 62.770 193.220 ;
        RECT 62.940 192.930 63.325 193.500 ;
        RECT 63.495 194.170 63.770 195.140 ;
        RECT 63.980 194.510 64.260 195.310 ;
        RECT 64.430 194.800 66.045 195.130 ;
        RECT 64.430 194.460 65.605 194.630 ;
        RECT 64.430 194.340 64.600 194.460 ;
        RECT 63.940 194.170 64.600 194.340 ;
        RECT 63.495 193.435 63.665 194.170 ;
        RECT 63.940 194.000 64.110 194.170 ;
        RECT 64.860 194.000 65.105 194.290 ;
        RECT 65.275 194.170 65.605 194.460 ;
        RECT 65.865 194.000 66.035 194.560 ;
        RECT 66.285 194.170 66.545 195.310 ;
        RECT 66.715 194.145 67.005 195.310 ;
        RECT 67.175 194.170 67.435 195.310 ;
        RECT 67.605 194.340 67.935 195.140 ;
        RECT 68.105 194.510 68.275 195.310 ;
        RECT 68.475 194.340 68.805 195.140 ;
        RECT 69.005 194.510 69.285 195.310 ;
        RECT 67.605 194.170 68.885 194.340 ;
        RECT 63.835 193.670 64.110 194.000 ;
        RECT 64.280 193.670 65.105 194.000 ;
        RECT 65.320 193.670 66.035 194.000 ;
        RECT 66.205 193.750 66.540 194.000 ;
        RECT 67.200 193.670 67.485 194.000 ;
        RECT 67.685 193.670 68.065 194.000 ;
        RECT 68.235 193.670 68.545 194.000 ;
        RECT 63.940 193.500 64.110 193.670 ;
        RECT 65.785 193.580 66.035 193.670 ;
        RECT 63.495 193.090 63.770 193.435 ;
        RECT 63.940 193.330 65.605 193.500 ;
        RECT 63.960 192.760 64.335 193.160 ;
        RECT 64.505 192.980 64.675 193.330 ;
        RECT 64.845 192.760 65.175 193.160 ;
        RECT 65.345 192.930 65.605 193.330 ;
        RECT 65.785 193.160 66.115 193.580 ;
        RECT 66.285 192.760 66.545 193.580 ;
        RECT 66.715 192.760 67.005 193.485 ;
        RECT 67.180 192.760 67.515 193.500 ;
        RECT 67.685 192.975 67.900 193.670 ;
        RECT 68.235 193.500 68.440 193.670 ;
        RECT 68.715 193.500 68.885 194.170 ;
        RECT 69.065 193.670 69.305 194.340 ;
        RECT 69.475 194.220 71.145 195.310 ;
        RECT 71.690 194.330 71.945 195.000 ;
        RECT 72.125 194.510 72.410 195.310 ;
        RECT 72.590 194.590 72.920 195.100 ;
        RECT 69.475 193.700 70.225 194.220 ;
        RECT 70.395 193.530 71.145 194.050 ;
        RECT 68.090 192.975 68.440 193.500 ;
        RECT 68.610 192.930 69.305 193.500 ;
        RECT 69.475 192.760 71.145 193.530 ;
        RECT 71.690 193.470 71.870 194.330 ;
        RECT 72.590 194.000 72.840 194.590 ;
        RECT 73.190 194.440 73.360 195.050 ;
        RECT 73.530 194.620 73.860 195.310 ;
        RECT 74.090 194.760 74.330 195.050 ;
        RECT 74.530 194.930 74.950 195.310 ;
        RECT 75.130 194.840 75.760 195.090 ;
        RECT 76.230 194.930 76.560 195.310 ;
        RECT 75.130 194.760 75.300 194.840 ;
        RECT 76.730 194.760 76.900 195.050 ;
        RECT 77.080 194.930 77.460 195.310 ;
        RECT 77.700 194.925 78.530 195.095 ;
        RECT 74.090 194.590 75.300 194.760 ;
        RECT 72.040 193.670 72.840 194.000 ;
        RECT 71.690 193.270 71.945 193.470 ;
        RECT 71.605 193.100 71.945 193.270 ;
        RECT 71.690 192.940 71.945 193.100 ;
        RECT 72.125 192.760 72.410 193.220 ;
        RECT 72.590 193.020 72.840 193.670 ;
        RECT 73.040 194.420 73.360 194.440 ;
        RECT 73.040 194.250 74.960 194.420 ;
        RECT 73.040 193.355 73.230 194.250 ;
        RECT 75.130 194.080 75.300 194.590 ;
        RECT 75.470 194.330 75.990 194.640 ;
        RECT 73.400 193.910 75.300 194.080 ;
        RECT 73.400 193.850 73.730 193.910 ;
        RECT 73.880 193.680 74.210 193.740 ;
        RECT 73.550 193.410 74.210 193.680 ;
        RECT 73.040 193.025 73.360 193.355 ;
        RECT 73.540 192.760 74.200 193.240 ;
        RECT 74.400 193.150 74.570 193.910 ;
        RECT 75.470 193.740 75.650 194.150 ;
        RECT 74.740 193.570 75.070 193.690 ;
        RECT 75.820 193.570 75.990 194.330 ;
        RECT 74.740 193.400 75.990 193.570 ;
        RECT 76.160 194.510 77.530 194.760 ;
        RECT 76.160 193.740 76.350 194.510 ;
        RECT 77.280 194.250 77.530 194.510 ;
        RECT 76.520 194.080 76.770 194.240 ;
        RECT 77.700 194.080 77.870 194.925 ;
        RECT 78.765 194.640 78.935 195.140 ;
        RECT 79.105 194.810 79.435 195.310 ;
        RECT 78.040 194.250 78.540 194.630 ;
        RECT 78.765 194.470 79.460 194.640 ;
        RECT 76.520 193.910 77.870 194.080 ;
        RECT 77.450 193.870 77.870 193.910 ;
        RECT 76.160 193.400 76.580 193.740 ;
        RECT 76.870 193.410 77.280 193.740 ;
        RECT 74.400 192.980 75.250 193.150 ;
        RECT 75.810 192.760 76.130 193.220 ;
        RECT 76.330 192.970 76.580 193.400 ;
        RECT 76.870 192.760 77.280 193.200 ;
        RECT 77.450 193.140 77.620 193.870 ;
        RECT 77.790 193.320 78.140 193.690 ;
        RECT 78.320 193.380 78.540 194.250 ;
        RECT 78.710 193.680 79.120 194.300 ;
        RECT 79.290 193.500 79.460 194.470 ;
        RECT 78.765 193.310 79.460 193.500 ;
        RECT 77.450 192.940 78.465 193.140 ;
        RECT 78.765 192.980 78.935 193.310 ;
        RECT 79.105 192.760 79.435 193.140 ;
        RECT 79.650 193.020 79.875 195.140 ;
        RECT 80.045 194.810 80.375 195.310 ;
        RECT 80.545 194.640 80.715 195.140 ;
        RECT 80.050 194.470 80.715 194.640 ;
        RECT 80.050 193.480 80.280 194.470 ;
        RECT 80.450 193.650 80.800 194.300 ;
        RECT 81.035 194.170 81.245 195.310 ;
        RECT 81.415 194.160 81.745 195.140 ;
        RECT 81.915 194.170 82.145 195.310 ;
        RECT 82.820 194.875 88.165 195.310 ;
        RECT 80.050 193.310 80.715 193.480 ;
        RECT 80.045 192.760 80.375 193.140 ;
        RECT 80.545 193.020 80.715 193.310 ;
        RECT 81.035 192.760 81.245 193.580 ;
        RECT 81.415 193.560 81.665 194.160 ;
        RECT 81.835 193.750 82.165 194.000 ;
        RECT 84.410 193.625 84.760 194.875 ;
        RECT 88.340 194.170 88.675 195.140 ;
        RECT 88.845 194.170 89.015 195.310 ;
        RECT 89.185 194.970 91.215 195.140 ;
        RECT 81.415 192.930 81.745 193.560 ;
        RECT 81.915 192.760 82.145 193.580 ;
        RECT 86.240 193.305 86.580 194.135 ;
        RECT 88.340 193.500 88.510 194.170 ;
        RECT 89.185 194.000 89.355 194.970 ;
        RECT 88.680 193.670 88.935 194.000 ;
        RECT 89.160 193.670 89.355 194.000 ;
        RECT 89.525 194.630 90.650 194.800 ;
        RECT 88.765 193.500 88.935 193.670 ;
        RECT 89.525 193.500 89.695 194.630 ;
        RECT 82.820 192.760 88.165 193.305 ;
        RECT 88.340 192.930 88.595 193.500 ;
        RECT 88.765 193.330 89.695 193.500 ;
        RECT 89.865 194.290 90.875 194.460 ;
        RECT 89.865 193.490 90.035 194.290 ;
        RECT 89.520 193.295 89.695 193.330 ;
        RECT 88.765 192.760 89.095 193.160 ;
        RECT 89.520 192.930 90.050 193.295 ;
        RECT 90.240 193.270 90.515 194.090 ;
        RECT 90.235 193.100 90.515 193.270 ;
        RECT 90.240 192.930 90.515 193.100 ;
        RECT 90.685 192.930 90.875 194.290 ;
        RECT 91.045 194.305 91.215 194.970 ;
        RECT 91.385 194.550 91.555 195.310 ;
        RECT 91.790 194.550 92.305 194.960 ;
        RECT 91.045 194.115 91.795 194.305 ;
        RECT 91.965 193.740 92.305 194.550 ;
        RECT 92.475 194.145 92.765 195.310 ;
        RECT 92.935 194.220 94.605 195.310 ;
        RECT 94.775 194.550 95.290 194.960 ;
        RECT 95.525 194.550 95.695 195.310 ;
        RECT 95.865 194.970 97.895 195.140 ;
        RECT 91.075 193.570 92.305 193.740 ;
        RECT 92.935 193.700 93.685 194.220 ;
        RECT 91.055 192.760 91.565 193.295 ;
        RECT 91.785 192.965 92.030 193.570 ;
        RECT 93.855 193.530 94.605 194.050 ;
        RECT 94.775 193.740 95.115 194.550 ;
        RECT 95.865 194.305 96.035 194.970 ;
        RECT 96.430 194.630 97.555 194.800 ;
        RECT 95.285 194.115 96.035 194.305 ;
        RECT 96.205 194.290 97.215 194.460 ;
        RECT 94.775 193.570 96.005 193.740 ;
        RECT 92.475 192.760 92.765 193.485 ;
        RECT 92.935 192.760 94.605 193.530 ;
        RECT 95.050 192.965 95.295 193.570 ;
        RECT 95.515 192.760 96.025 193.295 ;
        RECT 96.205 192.930 96.395 194.290 ;
        RECT 96.565 193.270 96.840 194.090 ;
        RECT 97.045 193.490 97.215 194.290 ;
        RECT 97.385 193.500 97.555 194.630 ;
        RECT 97.725 194.000 97.895 194.970 ;
        RECT 98.065 194.170 98.235 195.310 ;
        RECT 98.405 194.170 98.740 195.140 ;
        RECT 97.725 193.670 97.920 194.000 ;
        RECT 98.145 193.670 98.400 194.000 ;
        RECT 98.145 193.500 98.315 193.670 ;
        RECT 98.570 193.500 98.740 194.170 ;
        RECT 98.915 194.550 99.430 194.960 ;
        RECT 99.665 194.550 99.835 195.310 ;
        RECT 100.005 194.970 102.035 195.140 ;
        RECT 98.915 193.740 99.255 194.550 ;
        RECT 100.005 194.305 100.175 194.970 ;
        RECT 100.570 194.630 101.695 194.800 ;
        RECT 99.425 194.115 100.175 194.305 ;
        RECT 100.345 194.290 101.355 194.460 ;
        RECT 98.915 193.570 100.145 193.740 ;
        RECT 97.385 193.330 98.315 193.500 ;
        RECT 97.385 193.295 97.560 193.330 ;
        RECT 96.565 193.100 96.845 193.270 ;
        RECT 96.565 192.930 96.840 193.100 ;
        RECT 97.030 192.930 97.560 193.295 ;
        RECT 97.985 192.760 98.315 193.160 ;
        RECT 98.485 192.930 98.740 193.500 ;
        RECT 99.190 192.965 99.435 193.570 ;
        RECT 99.655 192.760 100.165 193.295 ;
        RECT 100.345 192.930 100.535 194.290 ;
        RECT 100.705 193.270 100.980 194.090 ;
        RECT 101.185 193.490 101.355 194.290 ;
        RECT 101.525 193.500 101.695 194.630 ;
        RECT 101.865 194.000 102.035 194.970 ;
        RECT 102.205 194.170 102.375 195.310 ;
        RECT 102.545 194.170 102.880 195.140 ;
        RECT 101.865 193.670 102.060 194.000 ;
        RECT 102.285 193.670 102.540 194.000 ;
        RECT 102.285 193.500 102.455 193.670 ;
        RECT 102.710 193.500 102.880 194.170 ;
        RECT 103.515 194.220 106.105 195.310 ;
        RECT 106.280 194.875 111.625 195.310 ;
        RECT 111.800 194.875 117.145 195.310 ;
        RECT 103.515 193.700 104.725 194.220 ;
        RECT 104.895 193.530 106.105 194.050 ;
        RECT 107.870 193.625 108.220 194.875 ;
        RECT 101.525 193.330 102.455 193.500 ;
        RECT 101.525 193.295 101.700 193.330 ;
        RECT 100.705 193.100 100.985 193.270 ;
        RECT 100.705 192.930 100.980 193.100 ;
        RECT 101.170 192.930 101.700 193.295 ;
        RECT 102.125 192.760 102.455 193.160 ;
        RECT 102.625 192.930 102.880 193.500 ;
        RECT 103.515 192.760 106.105 193.530 ;
        RECT 109.700 193.305 110.040 194.135 ;
        RECT 113.390 193.625 113.740 194.875 ;
        RECT 117.315 194.220 118.525 195.310 ;
        RECT 115.220 193.305 115.560 194.135 ;
        RECT 117.315 193.680 117.835 194.220 ;
        RECT 118.005 193.510 118.525 194.050 ;
        RECT 106.280 192.760 111.625 193.305 ;
        RECT 111.800 192.760 117.145 193.305 ;
        RECT 117.315 192.760 118.525 193.510 ;
        RECT 11.430 192.590 118.610 192.760 ;
        RECT 11.515 191.840 12.725 192.590 ;
        RECT 11.515 191.300 12.035 191.840 ;
        RECT 12.895 191.820 14.565 192.590 ;
        RECT 14.740 192.045 20.085 192.590 ;
        RECT 12.205 191.130 12.725 191.670 ;
        RECT 11.515 190.040 12.725 191.130 ;
        RECT 12.895 191.130 13.645 191.650 ;
        RECT 13.815 191.300 14.565 191.820 ;
        RECT 12.895 190.040 14.565 191.130 ;
        RECT 16.330 190.475 16.680 191.725 ;
        RECT 18.160 191.215 18.500 192.045 ;
        RECT 20.370 191.960 20.655 192.420 ;
        RECT 20.825 192.130 21.095 192.590 ;
        RECT 20.370 191.790 21.325 191.960 ;
        RECT 20.255 191.060 20.945 191.620 ;
        RECT 21.115 190.890 21.325 191.790 ;
        RECT 20.370 190.670 21.325 190.890 ;
        RECT 21.495 191.620 21.895 192.420 ;
        RECT 22.085 191.960 22.365 192.420 ;
        RECT 22.885 192.130 23.210 192.590 ;
        RECT 22.085 191.790 23.210 191.960 ;
        RECT 23.380 191.850 23.765 192.420 ;
        RECT 22.760 191.680 23.210 191.790 ;
        RECT 21.495 191.060 22.590 191.620 ;
        RECT 22.760 191.350 23.315 191.680 ;
        RECT 14.740 190.040 20.085 190.475 ;
        RECT 20.370 190.210 20.655 190.670 ;
        RECT 20.825 190.040 21.095 190.500 ;
        RECT 21.495 190.210 21.895 191.060 ;
        RECT 22.760 190.890 23.210 191.350 ;
        RECT 23.485 191.180 23.765 191.850 ;
        RECT 24.210 191.780 24.455 192.385 ;
        RECT 24.675 192.055 25.185 192.590 ;
        RECT 22.085 190.670 23.210 190.890 ;
        RECT 22.085 190.210 22.365 190.670 ;
        RECT 22.885 190.040 23.210 190.500 ;
        RECT 23.380 190.210 23.765 191.180 ;
        RECT 23.935 191.610 25.165 191.780 ;
        RECT 23.935 190.800 24.275 191.610 ;
        RECT 24.445 191.045 25.195 191.235 ;
        RECT 23.935 190.390 24.450 190.800 ;
        RECT 24.685 190.040 24.855 190.800 ;
        RECT 25.025 190.380 25.195 191.045 ;
        RECT 25.365 191.060 25.555 192.420 ;
        RECT 25.725 191.910 26.000 192.420 ;
        RECT 26.190 192.055 26.720 192.420 ;
        RECT 27.145 192.190 27.475 192.590 ;
        RECT 26.545 192.020 26.720 192.055 ;
        RECT 25.725 191.740 26.005 191.910 ;
        RECT 25.725 191.260 26.000 191.740 ;
        RECT 26.205 191.060 26.375 191.860 ;
        RECT 25.365 190.890 26.375 191.060 ;
        RECT 26.545 191.850 27.475 192.020 ;
        RECT 27.645 191.850 27.900 192.420 ;
        RECT 28.075 191.865 28.365 192.590 ;
        RECT 26.545 190.720 26.715 191.850 ;
        RECT 27.305 191.680 27.475 191.850 ;
        RECT 25.590 190.550 26.715 190.720 ;
        RECT 26.885 191.350 27.080 191.680 ;
        RECT 27.305 191.350 27.560 191.680 ;
        RECT 26.885 190.380 27.055 191.350 ;
        RECT 27.730 191.180 27.900 191.850 ;
        RECT 29.495 191.770 29.725 192.590 ;
        RECT 29.895 191.790 30.225 192.420 ;
        RECT 29.475 191.350 29.805 191.600 ;
        RECT 25.025 190.210 27.055 190.380 ;
        RECT 27.225 190.040 27.395 191.180 ;
        RECT 27.565 190.210 27.900 191.180 ;
        RECT 28.075 190.040 28.365 191.205 ;
        RECT 29.975 191.190 30.225 191.790 ;
        RECT 30.395 191.770 30.605 192.590 ;
        RECT 30.875 191.770 31.105 192.590 ;
        RECT 31.275 191.790 31.605 192.420 ;
        RECT 30.855 191.350 31.185 191.600 ;
        RECT 31.355 191.190 31.605 191.790 ;
        RECT 31.775 191.770 31.985 192.590 ;
        RECT 32.220 191.880 32.475 192.410 ;
        RECT 32.645 192.130 32.950 192.590 ;
        RECT 33.195 192.210 34.265 192.380 ;
        RECT 29.495 190.040 29.725 191.180 ;
        RECT 29.895 190.210 30.225 191.190 ;
        RECT 30.395 190.040 30.605 191.180 ;
        RECT 30.875 190.040 31.105 191.180 ;
        RECT 31.275 190.210 31.605 191.190 ;
        RECT 32.220 191.230 32.430 191.880 ;
        RECT 33.195 191.855 33.515 192.210 ;
        RECT 33.190 191.680 33.515 191.855 ;
        RECT 32.600 191.380 33.515 191.680 ;
        RECT 33.685 191.640 33.925 192.040 ;
        RECT 34.095 191.980 34.265 192.210 ;
        RECT 34.435 192.150 34.625 192.590 ;
        RECT 34.795 192.140 35.745 192.420 ;
        RECT 35.965 192.230 36.315 192.400 ;
        RECT 34.095 191.810 34.625 191.980 ;
        RECT 32.600 191.350 33.340 191.380 ;
        RECT 31.775 190.040 31.985 191.180 ;
        RECT 32.220 190.350 32.475 191.230 ;
        RECT 32.645 190.040 32.950 191.180 ;
        RECT 33.170 190.760 33.340 191.350 ;
        RECT 33.685 191.270 34.225 191.640 ;
        RECT 34.405 191.530 34.625 191.810 ;
        RECT 34.795 191.360 34.965 192.140 ;
        RECT 34.560 191.190 34.965 191.360 ;
        RECT 35.135 191.350 35.485 191.970 ;
        RECT 34.560 191.100 34.730 191.190 ;
        RECT 35.655 191.180 35.865 191.970 ;
        RECT 33.510 190.930 34.730 191.100 ;
        RECT 35.190 191.020 35.865 191.180 ;
        RECT 33.170 190.590 33.970 190.760 ;
        RECT 33.290 190.040 33.620 190.420 ;
        RECT 33.800 190.300 33.970 190.590 ;
        RECT 34.560 190.550 34.730 190.930 ;
        RECT 34.900 191.010 35.865 191.020 ;
        RECT 36.055 191.840 36.315 192.230 ;
        RECT 36.525 192.130 36.855 192.590 ;
        RECT 37.730 192.200 38.585 192.370 ;
        RECT 38.790 192.200 39.285 192.370 ;
        RECT 39.455 192.230 39.785 192.590 ;
        RECT 36.055 191.150 36.225 191.840 ;
        RECT 36.395 191.490 36.565 191.670 ;
        RECT 36.735 191.660 37.525 191.910 ;
        RECT 37.730 191.490 37.900 192.200 ;
        RECT 38.070 191.690 38.425 191.910 ;
        RECT 36.395 191.320 38.085 191.490 ;
        RECT 34.900 190.720 35.360 191.010 ;
        RECT 36.055 190.980 37.555 191.150 ;
        RECT 36.055 190.840 36.225 190.980 ;
        RECT 35.665 190.670 36.225 190.840 ;
        RECT 34.140 190.040 34.390 190.500 ;
        RECT 34.560 190.210 35.430 190.550 ;
        RECT 35.665 190.210 35.835 190.670 ;
        RECT 36.670 190.640 37.745 190.810 ;
        RECT 36.005 190.040 36.375 190.500 ;
        RECT 36.670 190.300 36.840 190.640 ;
        RECT 37.010 190.040 37.340 190.470 ;
        RECT 37.575 190.300 37.745 190.640 ;
        RECT 37.915 190.540 38.085 191.320 ;
        RECT 38.255 191.100 38.425 191.690 ;
        RECT 38.595 191.290 38.945 191.910 ;
        RECT 38.255 190.710 38.720 191.100 ;
        RECT 39.115 190.840 39.285 192.200 ;
        RECT 39.455 191.010 39.915 192.060 ;
        RECT 38.890 190.670 39.285 190.840 ;
        RECT 38.890 190.540 39.060 190.670 ;
        RECT 37.915 190.210 38.595 190.540 ;
        RECT 38.810 190.210 39.060 190.540 ;
        RECT 39.230 190.040 39.480 190.500 ;
        RECT 39.650 190.225 39.975 191.010 ;
        RECT 40.145 190.210 40.315 192.330 ;
        RECT 40.485 192.210 40.815 192.590 ;
        RECT 40.985 192.040 41.240 192.330 ;
        RECT 40.490 191.870 41.240 192.040 ;
        RECT 40.490 190.880 40.720 191.870 ;
        RECT 41.875 191.820 45.385 192.590 ;
        RECT 40.890 191.050 41.240 191.700 ;
        RECT 41.875 191.130 43.565 191.650 ;
        RECT 43.735 191.300 45.385 191.820 ;
        RECT 45.830 191.780 46.075 192.385 ;
        RECT 46.295 192.055 46.805 192.590 ;
        RECT 45.555 191.610 46.785 191.780 ;
        RECT 40.490 190.710 41.240 190.880 ;
        RECT 40.485 190.040 40.815 190.540 ;
        RECT 40.985 190.210 41.240 190.710 ;
        RECT 41.875 190.040 45.385 191.130 ;
        RECT 45.555 190.800 45.895 191.610 ;
        RECT 46.065 191.045 46.815 191.235 ;
        RECT 45.555 190.390 46.070 190.800 ;
        RECT 46.305 190.040 46.475 190.800 ;
        RECT 46.645 190.380 46.815 191.045 ;
        RECT 46.985 191.060 47.175 192.420 ;
        RECT 47.345 191.570 47.620 192.420 ;
        RECT 47.810 192.055 48.340 192.420 ;
        RECT 48.765 192.190 49.095 192.590 ;
        RECT 48.165 192.020 48.340 192.055 ;
        RECT 47.345 191.400 47.625 191.570 ;
        RECT 47.345 191.260 47.620 191.400 ;
        RECT 47.825 191.060 47.995 191.860 ;
        RECT 46.985 190.890 47.995 191.060 ;
        RECT 48.165 191.850 49.095 192.020 ;
        RECT 49.265 191.850 49.520 192.420 ;
        RECT 48.165 190.720 48.335 191.850 ;
        RECT 48.925 191.680 49.095 191.850 ;
        RECT 47.210 190.550 48.335 190.720 ;
        RECT 48.505 191.350 48.700 191.680 ;
        RECT 48.925 191.350 49.180 191.680 ;
        RECT 48.505 190.380 48.675 191.350 ;
        RECT 49.350 191.180 49.520 191.850 ;
        RECT 50.215 191.770 50.425 192.590 ;
        RECT 50.595 191.790 50.925 192.420 ;
        RECT 50.595 191.190 50.845 191.790 ;
        RECT 51.095 191.770 51.325 192.590 ;
        RECT 52.085 192.040 52.255 192.420 ;
        RECT 52.435 192.210 52.765 192.590 ;
        RECT 52.085 191.870 52.750 192.040 ;
        RECT 52.945 191.915 53.205 192.420 ;
        RECT 51.015 191.350 51.345 191.600 ;
        RECT 52.015 191.320 52.345 191.690 ;
        RECT 52.580 191.615 52.750 191.870 ;
        RECT 52.580 191.285 52.865 191.615 ;
        RECT 46.645 190.210 48.675 190.380 ;
        RECT 48.845 190.040 49.015 191.180 ;
        RECT 49.185 190.210 49.520 191.180 ;
        RECT 50.215 190.040 50.425 191.180 ;
        RECT 50.595 190.210 50.925 191.190 ;
        RECT 51.095 190.040 51.325 191.180 ;
        RECT 52.580 191.140 52.750 191.285 ;
        RECT 52.085 190.970 52.750 191.140 ;
        RECT 53.035 191.115 53.205 191.915 ;
        RECT 53.835 191.865 54.125 192.590 ;
        RECT 54.755 191.820 56.425 192.590 ;
        RECT 52.085 190.210 52.255 190.970 ;
        RECT 52.435 190.040 52.765 190.800 ;
        RECT 52.935 190.210 53.205 191.115 ;
        RECT 53.835 190.040 54.125 191.205 ;
        RECT 54.755 191.130 55.505 191.650 ;
        RECT 55.675 191.300 56.425 191.820 ;
        RECT 56.635 191.770 56.865 192.590 ;
        RECT 57.035 191.790 57.365 192.420 ;
        RECT 56.615 191.350 56.945 191.600 ;
        RECT 57.115 191.190 57.365 191.790 ;
        RECT 57.535 191.770 57.745 192.590 ;
        RECT 57.980 191.880 58.235 192.410 ;
        RECT 58.405 192.130 58.710 192.590 ;
        RECT 58.955 192.210 60.025 192.380 ;
        RECT 54.755 190.040 56.425 191.130 ;
        RECT 56.635 190.040 56.865 191.180 ;
        RECT 57.035 190.210 57.365 191.190 ;
        RECT 57.980 191.230 58.190 191.880 ;
        RECT 58.955 191.855 59.275 192.210 ;
        RECT 58.950 191.680 59.275 191.855 ;
        RECT 58.360 191.380 59.275 191.680 ;
        RECT 59.445 191.640 59.685 192.040 ;
        RECT 59.855 191.980 60.025 192.210 ;
        RECT 60.195 192.150 60.385 192.590 ;
        RECT 60.555 192.140 61.505 192.420 ;
        RECT 61.725 192.230 62.075 192.400 ;
        RECT 59.855 191.810 60.385 191.980 ;
        RECT 58.360 191.350 59.100 191.380 ;
        RECT 57.535 190.040 57.745 191.180 ;
        RECT 57.980 190.350 58.235 191.230 ;
        RECT 58.405 190.040 58.710 191.180 ;
        RECT 58.930 190.760 59.100 191.350 ;
        RECT 59.445 191.270 59.985 191.640 ;
        RECT 60.165 191.530 60.385 191.810 ;
        RECT 60.555 191.360 60.725 192.140 ;
        RECT 60.320 191.190 60.725 191.360 ;
        RECT 60.895 191.350 61.245 191.970 ;
        RECT 60.320 191.100 60.490 191.190 ;
        RECT 61.415 191.180 61.625 191.970 ;
        RECT 59.270 190.930 60.490 191.100 ;
        RECT 60.950 191.020 61.625 191.180 ;
        RECT 58.930 190.590 59.730 190.760 ;
        RECT 59.050 190.040 59.380 190.420 ;
        RECT 59.560 190.300 59.730 190.590 ;
        RECT 60.320 190.550 60.490 190.930 ;
        RECT 60.660 191.010 61.625 191.020 ;
        RECT 61.815 191.840 62.075 192.230 ;
        RECT 62.285 192.130 62.615 192.590 ;
        RECT 63.490 192.200 64.345 192.370 ;
        RECT 64.550 192.200 65.045 192.370 ;
        RECT 65.215 192.230 65.545 192.590 ;
        RECT 61.815 191.150 61.985 191.840 ;
        RECT 62.155 191.490 62.325 191.670 ;
        RECT 62.495 191.660 63.285 191.910 ;
        RECT 63.490 191.490 63.660 192.200 ;
        RECT 63.830 191.690 64.185 191.910 ;
        RECT 62.155 191.320 63.845 191.490 ;
        RECT 60.660 190.720 61.120 191.010 ;
        RECT 61.815 190.980 63.315 191.150 ;
        RECT 61.815 190.840 61.985 190.980 ;
        RECT 61.425 190.670 61.985 190.840 ;
        RECT 59.900 190.040 60.150 190.500 ;
        RECT 60.320 190.210 61.190 190.550 ;
        RECT 61.425 190.210 61.595 190.670 ;
        RECT 62.430 190.640 63.505 190.810 ;
        RECT 61.765 190.040 62.135 190.500 ;
        RECT 62.430 190.300 62.600 190.640 ;
        RECT 62.770 190.040 63.100 190.470 ;
        RECT 63.335 190.300 63.505 190.640 ;
        RECT 63.675 190.540 63.845 191.320 ;
        RECT 64.015 191.100 64.185 191.690 ;
        RECT 64.355 191.290 64.705 191.910 ;
        RECT 64.015 190.710 64.480 191.100 ;
        RECT 64.875 190.840 65.045 192.200 ;
        RECT 65.215 191.010 65.675 192.060 ;
        RECT 64.650 190.670 65.045 190.840 ;
        RECT 64.650 190.540 64.820 190.670 ;
        RECT 63.675 190.210 64.355 190.540 ;
        RECT 64.570 190.210 64.820 190.540 ;
        RECT 64.990 190.040 65.240 190.500 ;
        RECT 65.410 190.225 65.735 191.010 ;
        RECT 65.905 190.210 66.075 192.330 ;
        RECT 66.245 192.210 66.575 192.590 ;
        RECT 66.745 192.040 67.000 192.330 ;
        RECT 66.250 191.870 67.000 192.040 ;
        RECT 66.250 190.880 66.480 191.870 ;
        RECT 67.175 191.850 67.495 192.330 ;
        RECT 67.665 192.020 67.895 192.420 ;
        RECT 68.065 192.200 68.415 192.590 ;
        RECT 67.665 191.940 68.175 192.020 ;
        RECT 68.585 191.940 68.915 192.420 ;
        RECT 67.665 191.850 68.915 191.940 ;
        RECT 66.650 191.050 67.000 191.700 ;
        RECT 67.175 190.920 67.345 191.850 ;
        RECT 68.005 191.770 68.915 191.850 ;
        RECT 69.085 191.770 69.255 192.590 ;
        RECT 69.760 191.850 70.225 192.395 ;
        RECT 67.515 191.260 67.685 191.680 ;
        RECT 67.915 191.430 68.515 191.600 ;
        RECT 67.515 191.090 68.175 191.260 ;
        RECT 66.250 190.710 67.000 190.880 ;
        RECT 67.175 190.720 67.835 190.920 ;
        RECT 68.005 190.890 68.175 191.090 ;
        RECT 68.345 191.230 68.515 191.430 ;
        RECT 68.685 191.400 69.380 191.600 ;
        RECT 69.640 191.230 69.885 191.680 ;
        RECT 68.345 191.060 69.885 191.230 ;
        RECT 70.055 190.890 70.225 191.850 ;
        RECT 70.855 191.820 73.445 192.590 ;
        RECT 68.005 190.720 70.225 190.890 ;
        RECT 70.855 191.130 72.065 191.650 ;
        RECT 72.235 191.300 73.445 191.820 ;
        RECT 73.890 191.780 74.135 192.385 ;
        RECT 74.355 192.055 74.865 192.590 ;
        RECT 73.615 191.610 74.845 191.780 ;
        RECT 66.245 190.040 66.575 190.540 ;
        RECT 66.745 190.210 67.000 190.710 ;
        RECT 67.665 190.550 67.835 190.720 ;
        RECT 67.195 190.040 67.495 190.550 ;
        RECT 67.665 190.380 68.045 190.550 ;
        RECT 68.625 190.040 69.255 190.550 ;
        RECT 69.425 190.210 69.755 190.720 ;
        RECT 69.925 190.040 70.225 190.550 ;
        RECT 70.855 190.040 73.445 191.130 ;
        RECT 73.615 190.800 73.955 191.610 ;
        RECT 74.125 191.045 74.875 191.235 ;
        RECT 73.615 190.390 74.130 190.800 ;
        RECT 74.365 190.040 74.535 190.800 ;
        RECT 74.705 190.380 74.875 191.045 ;
        RECT 75.045 191.060 75.235 192.420 ;
        RECT 75.405 191.570 75.680 192.420 ;
        RECT 75.870 192.055 76.400 192.420 ;
        RECT 76.825 192.190 77.155 192.590 ;
        RECT 76.225 192.020 76.400 192.055 ;
        RECT 75.405 191.400 75.685 191.570 ;
        RECT 75.405 191.260 75.680 191.400 ;
        RECT 75.885 191.060 76.055 191.860 ;
        RECT 75.045 190.890 76.055 191.060 ;
        RECT 76.225 191.850 77.155 192.020 ;
        RECT 77.325 191.850 77.580 192.420 ;
        RECT 77.845 192.040 78.015 192.420 ;
        RECT 78.195 192.210 78.525 192.590 ;
        RECT 77.845 191.870 78.510 192.040 ;
        RECT 78.705 191.915 78.965 192.420 ;
        RECT 76.225 190.720 76.395 191.850 ;
        RECT 76.985 191.680 77.155 191.850 ;
        RECT 75.270 190.550 76.395 190.720 ;
        RECT 76.565 191.350 76.760 191.680 ;
        RECT 76.985 191.350 77.240 191.680 ;
        RECT 76.565 190.380 76.735 191.350 ;
        RECT 77.410 191.180 77.580 191.850 ;
        RECT 77.775 191.320 78.105 191.690 ;
        RECT 78.340 191.615 78.510 191.870 ;
        RECT 74.705 190.210 76.735 190.380 ;
        RECT 76.905 190.040 77.075 191.180 ;
        RECT 77.245 190.210 77.580 191.180 ;
        RECT 78.340 191.285 78.625 191.615 ;
        RECT 78.340 191.140 78.510 191.285 ;
        RECT 77.845 190.970 78.510 191.140 ;
        RECT 78.795 191.115 78.965 191.915 ;
        RECT 79.595 191.865 79.885 192.590 ;
        RECT 80.055 191.820 82.645 192.590 ;
        RECT 77.845 190.210 78.015 190.970 ;
        RECT 78.195 190.040 78.525 190.800 ;
        RECT 78.695 190.210 78.965 191.115 ;
        RECT 79.595 190.040 79.885 191.205 ;
        RECT 80.055 191.130 81.265 191.650 ;
        RECT 81.435 191.300 82.645 191.820 ;
        RECT 82.855 191.770 83.085 192.590 ;
        RECT 83.255 191.790 83.585 192.420 ;
        RECT 82.835 191.350 83.165 191.600 ;
        RECT 83.335 191.190 83.585 191.790 ;
        RECT 83.755 191.770 83.965 192.590 ;
        RECT 84.200 191.880 84.455 192.410 ;
        RECT 84.625 192.130 84.930 192.590 ;
        RECT 85.175 192.210 86.245 192.380 ;
        RECT 80.055 190.040 82.645 191.130 ;
        RECT 82.855 190.040 83.085 191.180 ;
        RECT 83.255 190.210 83.585 191.190 ;
        RECT 84.200 191.230 84.410 191.880 ;
        RECT 85.175 191.855 85.495 192.210 ;
        RECT 85.170 191.680 85.495 191.855 ;
        RECT 84.580 191.380 85.495 191.680 ;
        RECT 85.665 191.640 85.905 192.040 ;
        RECT 86.075 191.980 86.245 192.210 ;
        RECT 86.415 192.150 86.605 192.590 ;
        RECT 86.775 192.140 87.725 192.420 ;
        RECT 87.945 192.230 88.295 192.400 ;
        RECT 86.075 191.810 86.605 191.980 ;
        RECT 84.580 191.350 85.320 191.380 ;
        RECT 83.755 190.040 83.965 191.180 ;
        RECT 84.200 190.350 84.455 191.230 ;
        RECT 84.625 190.040 84.930 191.180 ;
        RECT 85.150 190.760 85.320 191.350 ;
        RECT 85.665 191.270 86.205 191.640 ;
        RECT 86.385 191.530 86.605 191.810 ;
        RECT 86.775 191.360 86.945 192.140 ;
        RECT 86.540 191.190 86.945 191.360 ;
        RECT 87.115 191.350 87.465 191.970 ;
        RECT 86.540 191.100 86.710 191.190 ;
        RECT 87.635 191.180 87.845 191.970 ;
        RECT 85.490 190.930 86.710 191.100 ;
        RECT 87.170 191.020 87.845 191.180 ;
        RECT 85.150 190.590 85.950 190.760 ;
        RECT 85.270 190.040 85.600 190.420 ;
        RECT 85.780 190.300 85.950 190.590 ;
        RECT 86.540 190.550 86.710 190.930 ;
        RECT 86.880 191.010 87.845 191.020 ;
        RECT 88.035 191.840 88.295 192.230 ;
        RECT 88.505 192.130 88.835 192.590 ;
        RECT 89.710 192.200 90.565 192.370 ;
        RECT 90.770 192.200 91.265 192.370 ;
        RECT 91.435 192.230 91.765 192.590 ;
        RECT 88.035 191.150 88.205 191.840 ;
        RECT 88.375 191.490 88.545 191.670 ;
        RECT 88.715 191.660 89.505 191.910 ;
        RECT 89.710 191.490 89.880 192.200 ;
        RECT 90.050 191.690 90.405 191.910 ;
        RECT 88.375 191.320 90.065 191.490 ;
        RECT 86.880 190.720 87.340 191.010 ;
        RECT 88.035 190.980 89.535 191.150 ;
        RECT 88.035 190.840 88.205 190.980 ;
        RECT 87.645 190.670 88.205 190.840 ;
        RECT 86.120 190.040 86.370 190.500 ;
        RECT 86.540 190.210 87.410 190.550 ;
        RECT 87.645 190.210 87.815 190.670 ;
        RECT 88.650 190.640 89.725 190.810 ;
        RECT 87.985 190.040 88.355 190.500 ;
        RECT 88.650 190.300 88.820 190.640 ;
        RECT 88.990 190.040 89.320 190.470 ;
        RECT 89.555 190.300 89.725 190.640 ;
        RECT 89.895 190.540 90.065 191.320 ;
        RECT 90.235 191.100 90.405 191.690 ;
        RECT 90.575 191.290 90.925 191.910 ;
        RECT 90.235 190.710 90.700 191.100 ;
        RECT 91.095 190.840 91.265 192.200 ;
        RECT 91.435 191.010 91.895 192.060 ;
        RECT 90.870 190.670 91.265 190.840 ;
        RECT 90.870 190.540 91.040 190.670 ;
        RECT 89.895 190.210 90.575 190.540 ;
        RECT 90.790 190.210 91.040 190.540 ;
        RECT 91.210 190.040 91.460 190.500 ;
        RECT 91.630 190.225 91.955 191.010 ;
        RECT 92.125 190.210 92.295 192.330 ;
        RECT 92.465 192.210 92.795 192.590 ;
        RECT 92.965 192.040 93.220 192.330 ;
        RECT 92.470 191.870 93.220 192.040 ;
        RECT 93.400 191.880 93.655 192.410 ;
        RECT 93.825 192.130 94.130 192.590 ;
        RECT 94.375 192.210 95.445 192.380 ;
        RECT 92.470 190.880 92.700 191.870 ;
        RECT 92.870 191.050 93.220 191.700 ;
        RECT 93.400 191.230 93.610 191.880 ;
        RECT 94.375 191.855 94.695 192.210 ;
        RECT 94.370 191.680 94.695 191.855 ;
        RECT 93.780 191.380 94.695 191.680 ;
        RECT 94.865 191.640 95.105 192.040 ;
        RECT 95.275 191.980 95.445 192.210 ;
        RECT 95.615 192.150 95.805 192.590 ;
        RECT 95.975 192.140 96.925 192.420 ;
        RECT 97.145 192.230 97.495 192.400 ;
        RECT 95.275 191.810 95.805 191.980 ;
        RECT 93.780 191.350 94.520 191.380 ;
        RECT 92.470 190.710 93.220 190.880 ;
        RECT 92.465 190.040 92.795 190.540 ;
        RECT 92.965 190.210 93.220 190.710 ;
        RECT 93.400 190.350 93.655 191.230 ;
        RECT 93.825 190.040 94.130 191.180 ;
        RECT 94.350 190.760 94.520 191.350 ;
        RECT 94.865 191.270 95.405 191.640 ;
        RECT 95.585 191.530 95.805 191.810 ;
        RECT 95.975 191.360 96.145 192.140 ;
        RECT 95.740 191.190 96.145 191.360 ;
        RECT 96.315 191.350 96.665 191.970 ;
        RECT 95.740 191.100 95.910 191.190 ;
        RECT 96.835 191.180 97.045 191.970 ;
        RECT 94.690 190.930 95.910 191.100 ;
        RECT 96.370 191.020 97.045 191.180 ;
        RECT 94.350 190.590 95.150 190.760 ;
        RECT 94.470 190.040 94.800 190.420 ;
        RECT 94.980 190.300 95.150 190.590 ;
        RECT 95.740 190.550 95.910 190.930 ;
        RECT 96.080 191.010 97.045 191.020 ;
        RECT 97.235 191.840 97.495 192.230 ;
        RECT 97.705 192.130 98.035 192.590 ;
        RECT 98.910 192.200 99.765 192.370 ;
        RECT 99.970 192.200 100.465 192.370 ;
        RECT 100.635 192.230 100.965 192.590 ;
        RECT 97.235 191.150 97.405 191.840 ;
        RECT 97.575 191.490 97.745 191.670 ;
        RECT 97.915 191.660 98.705 191.910 ;
        RECT 98.910 191.490 99.080 192.200 ;
        RECT 99.250 191.690 99.605 191.910 ;
        RECT 97.575 191.320 99.265 191.490 ;
        RECT 96.080 190.720 96.540 191.010 ;
        RECT 97.235 190.980 98.735 191.150 ;
        RECT 97.235 190.840 97.405 190.980 ;
        RECT 96.845 190.670 97.405 190.840 ;
        RECT 95.320 190.040 95.570 190.500 ;
        RECT 95.740 190.210 96.610 190.550 ;
        RECT 96.845 190.210 97.015 190.670 ;
        RECT 97.850 190.640 98.925 190.810 ;
        RECT 97.185 190.040 97.555 190.500 ;
        RECT 97.850 190.300 98.020 190.640 ;
        RECT 98.190 190.040 98.520 190.470 ;
        RECT 98.755 190.300 98.925 190.640 ;
        RECT 99.095 190.540 99.265 191.320 ;
        RECT 99.435 191.100 99.605 191.690 ;
        RECT 99.775 191.290 100.125 191.910 ;
        RECT 99.435 190.710 99.900 191.100 ;
        RECT 100.295 190.840 100.465 192.200 ;
        RECT 100.635 191.010 101.095 192.060 ;
        RECT 100.070 190.670 100.465 190.840 ;
        RECT 100.070 190.540 100.240 190.670 ;
        RECT 99.095 190.210 99.775 190.540 ;
        RECT 99.990 190.210 100.240 190.540 ;
        RECT 100.410 190.040 100.660 190.500 ;
        RECT 100.830 190.225 101.155 191.010 ;
        RECT 101.325 190.210 101.495 192.330 ;
        RECT 101.665 192.210 101.995 192.590 ;
        RECT 102.165 192.040 102.420 192.330 ;
        RECT 101.670 191.870 102.420 192.040 ;
        RECT 101.670 190.880 101.900 191.870 ;
        RECT 102.595 191.820 105.185 192.590 ;
        RECT 105.355 191.865 105.645 192.590 ;
        RECT 105.815 191.820 108.405 192.590 ;
        RECT 102.070 191.050 102.420 191.700 ;
        RECT 102.595 191.130 103.805 191.650 ;
        RECT 103.975 191.300 105.185 191.820 ;
        RECT 101.670 190.710 102.420 190.880 ;
        RECT 101.665 190.040 101.995 190.540 ;
        RECT 102.165 190.210 102.420 190.710 ;
        RECT 102.595 190.040 105.185 191.130 ;
        RECT 105.355 190.040 105.645 191.205 ;
        RECT 105.815 191.130 107.025 191.650 ;
        RECT 107.195 191.300 108.405 191.820 ;
        RECT 108.635 191.770 108.845 192.590 ;
        RECT 109.015 191.790 109.345 192.420 ;
        RECT 109.015 191.190 109.265 191.790 ;
        RECT 109.515 191.770 109.745 192.590 ;
        RECT 109.955 191.820 111.625 192.590 ;
        RECT 111.800 192.045 117.145 192.590 ;
        RECT 109.435 191.350 109.765 191.600 ;
        RECT 105.815 190.040 108.405 191.130 ;
        RECT 108.635 190.040 108.845 191.180 ;
        RECT 109.015 190.210 109.345 191.190 ;
        RECT 109.515 190.040 109.745 191.180 ;
        RECT 109.955 191.130 110.705 191.650 ;
        RECT 110.875 191.300 111.625 191.820 ;
        RECT 109.955 190.040 111.625 191.130 ;
        RECT 113.390 190.475 113.740 191.725 ;
        RECT 115.220 191.215 115.560 192.045 ;
        RECT 117.315 191.840 118.525 192.590 ;
        RECT 117.315 191.130 117.835 191.670 ;
        RECT 118.005 191.300 118.525 191.840 ;
        RECT 111.800 190.040 117.145 190.475 ;
        RECT 117.315 190.040 118.525 191.130 ;
        RECT 11.430 189.870 118.610 190.040 ;
        RECT 11.515 188.780 12.725 189.870 ;
        RECT 11.515 188.070 12.035 188.610 ;
        RECT 12.205 188.240 12.725 188.780 ;
        RECT 13.355 188.780 15.025 189.870 ;
        RECT 13.355 188.260 14.105 188.780 ;
        RECT 15.195 188.705 15.485 189.870 ;
        RECT 15.655 188.780 19.165 189.870 ;
        RECT 14.275 188.090 15.025 188.610 ;
        RECT 15.655 188.260 17.345 188.780 ;
        RECT 19.375 188.730 19.605 189.870 ;
        RECT 19.775 188.720 20.105 189.700 ;
        RECT 20.275 188.730 20.485 189.870 ;
        RECT 17.515 188.090 19.165 188.610 ;
        RECT 19.355 188.310 19.685 188.560 ;
        RECT 11.515 187.320 12.725 188.070 ;
        RECT 13.355 187.320 15.025 188.090 ;
        RECT 15.195 187.320 15.485 188.045 ;
        RECT 15.655 187.320 19.165 188.090 ;
        RECT 19.375 187.320 19.605 188.140 ;
        RECT 19.855 188.120 20.105 188.720 ;
        RECT 20.720 188.680 20.975 189.560 ;
        RECT 21.145 188.730 21.450 189.870 ;
        RECT 21.790 189.490 22.120 189.870 ;
        RECT 22.300 189.320 22.470 189.610 ;
        RECT 22.640 189.410 22.890 189.870 ;
        RECT 21.670 189.150 22.470 189.320 ;
        RECT 23.060 189.360 23.930 189.700 ;
        RECT 19.775 187.490 20.105 188.120 ;
        RECT 20.275 187.320 20.485 188.140 ;
        RECT 20.720 188.030 20.930 188.680 ;
        RECT 21.670 188.560 21.840 189.150 ;
        RECT 23.060 188.980 23.230 189.360 ;
        RECT 24.165 189.240 24.335 189.700 ;
        RECT 24.505 189.410 24.875 189.870 ;
        RECT 25.170 189.270 25.340 189.610 ;
        RECT 25.510 189.440 25.840 189.870 ;
        RECT 26.075 189.270 26.245 189.610 ;
        RECT 22.010 188.810 23.230 188.980 ;
        RECT 23.400 188.900 23.860 189.190 ;
        RECT 24.165 189.070 24.725 189.240 ;
        RECT 25.170 189.100 26.245 189.270 ;
        RECT 26.415 189.370 27.095 189.700 ;
        RECT 27.310 189.370 27.560 189.700 ;
        RECT 27.730 189.410 27.980 189.870 ;
        RECT 24.555 188.930 24.725 189.070 ;
        RECT 23.400 188.890 24.365 188.900 ;
        RECT 23.060 188.720 23.230 188.810 ;
        RECT 23.690 188.730 24.365 188.890 ;
        RECT 21.100 188.530 21.840 188.560 ;
        RECT 21.100 188.230 22.015 188.530 ;
        RECT 21.690 188.055 22.015 188.230 ;
        RECT 20.720 187.500 20.975 188.030 ;
        RECT 21.145 187.320 21.450 187.780 ;
        RECT 21.695 187.700 22.015 188.055 ;
        RECT 22.185 188.270 22.725 188.640 ;
        RECT 23.060 188.550 23.465 188.720 ;
        RECT 22.185 187.870 22.425 188.270 ;
        RECT 22.905 188.100 23.125 188.380 ;
        RECT 22.595 187.930 23.125 188.100 ;
        RECT 22.595 187.700 22.765 187.930 ;
        RECT 23.295 187.770 23.465 188.550 ;
        RECT 23.635 187.940 23.985 188.560 ;
        RECT 24.155 187.940 24.365 188.730 ;
        RECT 24.555 188.760 26.055 188.930 ;
        RECT 24.555 188.070 24.725 188.760 ;
        RECT 26.415 188.590 26.585 189.370 ;
        RECT 27.390 189.240 27.560 189.370 ;
        RECT 24.895 188.420 26.585 188.590 ;
        RECT 26.755 188.810 27.220 189.200 ;
        RECT 27.390 189.070 27.785 189.240 ;
        RECT 24.895 188.240 25.065 188.420 ;
        RECT 21.695 187.530 22.765 187.700 ;
        RECT 22.935 187.320 23.125 187.760 ;
        RECT 23.295 187.490 24.245 187.770 ;
        RECT 24.555 187.680 24.815 188.070 ;
        RECT 25.235 188.000 26.025 188.250 ;
        RECT 24.465 187.510 24.815 187.680 ;
        RECT 25.025 187.320 25.355 187.780 ;
        RECT 26.230 187.710 26.400 188.420 ;
        RECT 26.755 188.220 26.925 188.810 ;
        RECT 26.570 188.000 26.925 188.220 ;
        RECT 27.095 188.000 27.445 188.620 ;
        RECT 27.615 187.710 27.785 189.070 ;
        RECT 28.150 188.900 28.475 189.685 ;
        RECT 27.955 187.850 28.415 188.900 ;
        RECT 26.230 187.540 27.085 187.710 ;
        RECT 27.290 187.540 27.785 187.710 ;
        RECT 27.955 187.320 28.285 187.680 ;
        RECT 28.645 187.580 28.815 189.700 ;
        RECT 28.985 189.370 29.315 189.870 ;
        RECT 29.485 189.200 29.740 189.700 ;
        RECT 28.990 189.030 29.740 189.200 ;
        RECT 28.990 188.040 29.220 189.030 ;
        RECT 30.925 188.940 31.095 189.700 ;
        RECT 31.275 189.110 31.605 189.870 ;
        RECT 29.390 188.210 29.740 188.860 ;
        RECT 30.925 188.770 31.590 188.940 ;
        RECT 31.775 188.795 32.045 189.700 ;
        RECT 31.420 188.625 31.590 188.770 ;
        RECT 30.855 188.220 31.185 188.590 ;
        RECT 31.420 188.295 31.705 188.625 ;
        RECT 31.420 188.040 31.590 188.295 ;
        RECT 28.990 187.870 29.740 188.040 ;
        RECT 28.985 187.320 29.315 187.700 ;
        RECT 29.485 187.580 29.740 187.870 ;
        RECT 30.925 187.870 31.590 188.040 ;
        RECT 31.875 187.995 32.045 188.795 ;
        RECT 30.925 187.490 31.095 187.870 ;
        RECT 31.275 187.320 31.605 187.700 ;
        RECT 31.785 187.490 32.045 187.995 ;
        RECT 32.220 188.730 32.555 189.700 ;
        RECT 32.725 188.730 32.895 189.870 ;
        RECT 33.065 189.530 35.095 189.700 ;
        RECT 32.220 188.060 32.390 188.730 ;
        RECT 33.065 188.560 33.235 189.530 ;
        RECT 32.560 188.230 32.815 188.560 ;
        RECT 33.040 188.230 33.235 188.560 ;
        RECT 33.405 189.190 34.530 189.360 ;
        RECT 32.645 188.060 32.815 188.230 ;
        RECT 33.405 188.060 33.575 189.190 ;
        RECT 32.220 187.490 32.475 188.060 ;
        RECT 32.645 187.890 33.575 188.060 ;
        RECT 33.745 188.850 34.755 189.020 ;
        RECT 33.745 188.050 33.915 188.850 ;
        RECT 33.400 187.855 33.575 187.890 ;
        RECT 32.645 187.320 32.975 187.720 ;
        RECT 33.400 187.490 33.930 187.855 ;
        RECT 34.120 187.830 34.395 188.650 ;
        RECT 34.115 187.660 34.395 187.830 ;
        RECT 34.120 187.490 34.395 187.660 ;
        RECT 34.565 187.490 34.755 188.850 ;
        RECT 34.925 188.865 35.095 189.530 ;
        RECT 35.265 189.110 35.435 189.870 ;
        RECT 35.670 189.110 36.185 189.520 ;
        RECT 34.925 188.675 35.675 188.865 ;
        RECT 35.845 188.300 36.185 189.110 ;
        RECT 34.955 188.130 36.185 188.300 ;
        RECT 36.355 189.110 36.870 189.520 ;
        RECT 37.105 189.110 37.275 189.870 ;
        RECT 37.445 189.530 39.475 189.700 ;
        RECT 36.355 188.300 36.695 189.110 ;
        RECT 37.445 188.865 37.615 189.530 ;
        RECT 38.010 189.190 39.135 189.360 ;
        RECT 36.865 188.675 37.615 188.865 ;
        RECT 37.785 188.850 38.795 189.020 ;
        RECT 36.355 188.130 37.585 188.300 ;
        RECT 34.935 187.320 35.445 187.855 ;
        RECT 35.665 187.525 35.910 188.130 ;
        RECT 36.630 187.525 36.875 188.130 ;
        RECT 37.095 187.320 37.605 187.855 ;
        RECT 37.785 187.490 37.975 188.850 ;
        RECT 38.145 188.170 38.420 188.650 ;
        RECT 38.145 188.000 38.425 188.170 ;
        RECT 38.625 188.050 38.795 188.850 ;
        RECT 38.965 188.060 39.135 189.190 ;
        RECT 39.305 188.560 39.475 189.530 ;
        RECT 39.645 188.730 39.815 189.870 ;
        RECT 39.985 188.730 40.320 189.700 ;
        RECT 39.305 188.230 39.500 188.560 ;
        RECT 39.725 188.230 39.980 188.560 ;
        RECT 39.725 188.060 39.895 188.230 ;
        RECT 40.150 188.060 40.320 188.730 ;
        RECT 40.955 188.705 41.245 189.870 ;
        RECT 41.415 188.780 44.925 189.870 ;
        RECT 41.415 188.260 43.105 188.780 ;
        RECT 45.135 188.730 45.365 189.870 ;
        RECT 45.535 188.720 45.865 189.700 ;
        RECT 46.035 188.730 46.245 189.870 ;
        RECT 46.850 188.890 47.105 189.560 ;
        RECT 47.285 189.070 47.570 189.870 ;
        RECT 47.750 189.150 48.080 189.660 ;
        RECT 43.275 188.090 44.925 188.610 ;
        RECT 45.115 188.310 45.445 188.560 ;
        RECT 38.145 187.490 38.420 188.000 ;
        RECT 38.965 187.890 39.895 188.060 ;
        RECT 38.965 187.855 39.140 187.890 ;
        RECT 38.610 187.490 39.140 187.855 ;
        RECT 39.565 187.320 39.895 187.720 ;
        RECT 40.065 187.490 40.320 188.060 ;
        RECT 40.955 187.320 41.245 188.045 ;
        RECT 41.415 187.320 44.925 188.090 ;
        RECT 45.135 187.320 45.365 188.140 ;
        RECT 45.615 188.120 45.865 188.720 ;
        RECT 46.850 188.170 47.030 188.890 ;
        RECT 47.750 188.560 48.000 189.150 ;
        RECT 48.350 189.000 48.520 189.610 ;
        RECT 48.690 189.180 49.020 189.870 ;
        RECT 49.250 189.320 49.490 189.610 ;
        RECT 49.690 189.490 50.110 189.870 ;
        RECT 50.290 189.400 50.920 189.650 ;
        RECT 51.390 189.490 51.720 189.870 ;
        RECT 50.290 189.320 50.460 189.400 ;
        RECT 51.890 189.320 52.060 189.610 ;
        RECT 52.240 189.490 52.620 189.870 ;
        RECT 52.860 189.485 53.690 189.655 ;
        RECT 49.250 189.150 50.460 189.320 ;
        RECT 47.200 188.230 48.000 188.560 ;
        RECT 45.535 187.490 45.865 188.120 ;
        RECT 46.035 187.320 46.245 188.140 ;
        RECT 46.765 188.030 47.030 188.170 ;
        RECT 46.765 188.000 47.105 188.030 ;
        RECT 46.850 187.500 47.105 188.000 ;
        RECT 47.285 187.320 47.570 187.780 ;
        RECT 47.750 187.580 48.000 188.230 ;
        RECT 48.200 188.980 48.520 189.000 ;
        RECT 48.200 188.810 50.120 188.980 ;
        RECT 48.200 187.915 48.390 188.810 ;
        RECT 50.290 188.640 50.460 189.150 ;
        RECT 50.630 188.890 51.150 189.200 ;
        RECT 48.560 188.470 50.460 188.640 ;
        RECT 48.560 188.410 48.890 188.470 ;
        RECT 49.040 188.240 49.370 188.300 ;
        RECT 48.710 187.970 49.370 188.240 ;
        RECT 48.200 187.585 48.520 187.915 ;
        RECT 48.700 187.320 49.360 187.800 ;
        RECT 49.560 187.710 49.730 188.470 ;
        RECT 50.630 188.300 50.810 188.710 ;
        RECT 49.900 188.130 50.230 188.250 ;
        RECT 50.980 188.130 51.150 188.890 ;
        RECT 49.900 187.960 51.150 188.130 ;
        RECT 51.320 189.070 52.690 189.320 ;
        RECT 51.320 188.300 51.510 189.070 ;
        RECT 52.440 188.810 52.690 189.070 ;
        RECT 51.680 188.640 51.930 188.800 ;
        RECT 52.860 188.640 53.030 189.485 ;
        RECT 53.925 189.200 54.095 189.700 ;
        RECT 54.265 189.370 54.595 189.870 ;
        RECT 53.200 188.810 53.700 189.190 ;
        RECT 53.925 189.030 54.620 189.200 ;
        RECT 51.680 188.470 53.030 188.640 ;
        RECT 52.610 188.430 53.030 188.470 ;
        RECT 51.320 187.960 51.740 188.300 ;
        RECT 52.030 187.970 52.440 188.300 ;
        RECT 49.560 187.540 50.410 187.710 ;
        RECT 50.970 187.320 51.290 187.780 ;
        RECT 51.490 187.530 51.740 187.960 ;
        RECT 52.030 187.320 52.440 187.760 ;
        RECT 52.610 187.700 52.780 188.430 ;
        RECT 52.950 187.880 53.300 188.250 ;
        RECT 53.480 187.940 53.700 188.810 ;
        RECT 53.870 188.240 54.280 188.860 ;
        RECT 54.450 188.060 54.620 189.030 ;
        RECT 53.925 187.870 54.620 188.060 ;
        RECT 52.610 187.500 53.625 187.700 ;
        RECT 53.925 187.540 54.095 187.870 ;
        RECT 54.265 187.320 54.595 187.700 ;
        RECT 54.810 187.580 55.035 189.700 ;
        RECT 55.205 189.370 55.535 189.870 ;
        RECT 55.705 189.200 55.875 189.700 ;
        RECT 55.210 189.030 55.875 189.200 ;
        RECT 55.210 188.040 55.440 189.030 ;
        RECT 55.610 188.210 55.960 188.860 ;
        RECT 56.595 188.780 58.265 189.870 ;
        RECT 58.440 189.435 63.785 189.870 ;
        RECT 56.595 188.260 57.345 188.780 ;
        RECT 57.515 188.090 58.265 188.610 ;
        RECT 60.030 188.185 60.380 189.435 ;
        RECT 63.965 188.890 64.295 189.700 ;
        RECT 64.465 189.070 64.705 189.870 ;
        RECT 63.965 188.720 64.680 188.890 ;
        RECT 55.210 187.870 55.875 188.040 ;
        RECT 55.205 187.320 55.535 187.700 ;
        RECT 55.705 187.580 55.875 187.870 ;
        RECT 56.595 187.320 58.265 188.090 ;
        RECT 61.860 187.865 62.200 188.695 ;
        RECT 63.960 188.310 64.340 188.550 ;
        RECT 64.510 188.480 64.680 188.720 ;
        RECT 64.885 188.850 65.055 189.700 ;
        RECT 65.225 189.070 65.555 189.870 ;
        RECT 65.725 188.850 65.895 189.700 ;
        RECT 64.885 188.680 65.895 188.850 ;
        RECT 66.065 188.720 66.395 189.870 ;
        RECT 66.715 188.705 67.005 189.870 ;
        RECT 67.175 188.780 68.385 189.870 ;
        RECT 68.560 189.435 73.905 189.870 ;
        RECT 64.510 188.310 65.010 188.480 ;
        RECT 64.510 188.140 64.680 188.310 ;
        RECT 65.400 188.140 65.895 188.680 ;
        RECT 67.175 188.240 67.695 188.780 ;
        RECT 64.045 187.970 64.680 188.140 ;
        RECT 64.885 187.970 65.895 188.140 ;
        RECT 58.440 187.320 63.785 187.865 ;
        RECT 64.045 187.490 64.215 187.970 ;
        RECT 64.395 187.320 64.635 187.800 ;
        RECT 64.885 187.490 65.055 187.970 ;
        RECT 65.225 187.320 65.555 187.800 ;
        RECT 65.725 187.490 65.895 187.970 ;
        RECT 66.065 187.320 66.395 188.120 ;
        RECT 67.865 188.070 68.385 188.610 ;
        RECT 70.150 188.185 70.500 189.435 ;
        RECT 74.135 188.730 74.345 189.870 ;
        RECT 74.515 188.720 74.845 189.700 ;
        RECT 75.015 188.730 75.245 189.870 ;
        RECT 75.915 188.780 78.505 189.870 ;
        RECT 66.715 187.320 67.005 188.045 ;
        RECT 67.175 187.320 68.385 188.070 ;
        RECT 71.980 187.865 72.320 188.695 ;
        RECT 68.560 187.320 73.905 187.865 ;
        RECT 74.135 187.320 74.345 188.140 ;
        RECT 74.515 188.120 74.765 188.720 ;
        RECT 74.935 188.310 75.265 188.560 ;
        RECT 75.915 188.260 77.125 188.780 ;
        RECT 78.715 188.730 78.945 189.870 ;
        RECT 79.115 188.720 79.445 189.700 ;
        RECT 79.615 188.730 79.825 189.870 ;
        RECT 80.055 188.795 80.325 189.700 ;
        RECT 80.495 189.110 80.825 189.870 ;
        RECT 81.005 188.940 81.175 189.700 ;
        RECT 74.515 187.490 74.845 188.120 ;
        RECT 75.015 187.320 75.245 188.140 ;
        RECT 77.295 188.090 78.505 188.610 ;
        RECT 78.695 188.310 79.025 188.560 ;
        RECT 75.915 187.320 78.505 188.090 ;
        RECT 78.715 187.320 78.945 188.140 ;
        RECT 79.195 188.120 79.445 188.720 ;
        RECT 79.115 187.490 79.445 188.120 ;
        RECT 79.615 187.320 79.825 188.140 ;
        RECT 80.055 187.995 80.225 188.795 ;
        RECT 80.510 188.770 81.175 188.940 ;
        RECT 82.355 189.110 82.870 189.520 ;
        RECT 83.105 189.110 83.275 189.870 ;
        RECT 83.445 189.530 85.475 189.700 ;
        RECT 80.510 188.625 80.680 188.770 ;
        RECT 80.395 188.295 80.680 188.625 ;
        RECT 80.510 188.040 80.680 188.295 ;
        RECT 80.915 188.220 81.245 188.590 ;
        RECT 82.355 188.300 82.695 189.110 ;
        RECT 83.445 188.865 83.615 189.530 ;
        RECT 84.010 189.190 85.135 189.360 ;
        RECT 82.865 188.675 83.615 188.865 ;
        RECT 83.785 188.850 84.795 189.020 ;
        RECT 82.355 188.130 83.585 188.300 ;
        RECT 80.055 187.490 80.315 187.995 ;
        RECT 80.510 187.870 81.175 188.040 ;
        RECT 80.495 187.320 80.825 187.700 ;
        RECT 81.005 187.490 81.175 187.870 ;
        RECT 82.630 187.525 82.875 188.130 ;
        RECT 83.095 187.320 83.605 187.855 ;
        RECT 83.785 187.490 83.975 188.850 ;
        RECT 84.145 187.830 84.420 188.650 ;
        RECT 84.625 188.050 84.795 188.850 ;
        RECT 84.965 188.060 85.135 189.190 ;
        RECT 85.305 188.560 85.475 189.530 ;
        RECT 85.645 188.730 85.815 189.870 ;
        RECT 85.985 188.730 86.320 189.700 ;
        RECT 87.045 188.940 87.215 189.700 ;
        RECT 87.395 189.110 87.725 189.870 ;
        RECT 87.045 188.770 87.710 188.940 ;
        RECT 87.895 188.795 88.165 189.700 ;
        RECT 85.305 188.230 85.500 188.560 ;
        RECT 85.725 188.230 85.980 188.560 ;
        RECT 85.725 188.060 85.895 188.230 ;
        RECT 86.150 188.060 86.320 188.730 ;
        RECT 87.540 188.625 87.710 188.770 ;
        RECT 86.975 188.220 87.305 188.590 ;
        RECT 87.540 188.295 87.825 188.625 ;
        RECT 84.965 187.890 85.895 188.060 ;
        RECT 84.965 187.855 85.140 187.890 ;
        RECT 84.145 187.660 84.425 187.830 ;
        RECT 84.145 187.490 84.420 187.660 ;
        RECT 84.610 187.490 85.140 187.855 ;
        RECT 85.565 187.320 85.895 187.720 ;
        RECT 86.065 187.490 86.320 188.060 ;
        RECT 87.540 188.040 87.710 188.295 ;
        RECT 87.045 187.870 87.710 188.040 ;
        RECT 87.995 187.995 88.165 188.795 ;
        RECT 87.045 187.490 87.215 187.870 ;
        RECT 87.395 187.320 87.725 187.700 ;
        RECT 87.905 187.490 88.165 187.995 ;
        RECT 88.335 188.730 88.720 189.700 ;
        RECT 88.890 189.410 89.215 189.870 ;
        RECT 89.735 189.240 90.015 189.700 ;
        RECT 88.890 189.020 90.015 189.240 ;
        RECT 88.335 188.060 88.615 188.730 ;
        RECT 88.890 188.560 89.340 189.020 ;
        RECT 90.205 188.850 90.605 189.700 ;
        RECT 91.005 189.410 91.275 189.870 ;
        RECT 91.445 189.240 91.730 189.700 ;
        RECT 88.785 188.230 89.340 188.560 ;
        RECT 89.510 188.290 90.605 188.850 ;
        RECT 88.890 188.120 89.340 188.230 ;
        RECT 88.335 187.490 88.720 188.060 ;
        RECT 88.890 187.950 90.015 188.120 ;
        RECT 88.890 187.320 89.215 187.780 ;
        RECT 89.735 187.490 90.015 187.950 ;
        RECT 90.205 187.490 90.605 188.290 ;
        RECT 90.775 189.020 91.730 189.240 ;
        RECT 90.775 188.120 90.985 189.020 ;
        RECT 91.155 188.290 91.845 188.850 ;
        RECT 92.475 188.705 92.765 189.870 ;
        RECT 92.935 188.780 94.145 189.870 ;
        RECT 92.935 188.240 93.455 188.780 ;
        RECT 94.355 188.730 94.585 189.870 ;
        RECT 94.755 188.720 95.085 189.700 ;
        RECT 95.255 188.730 95.465 189.870 ;
        RECT 96.155 188.780 97.825 189.870 ;
        RECT 98.085 188.940 98.255 189.700 ;
        RECT 98.435 189.110 98.765 189.870 ;
        RECT 90.775 187.950 91.730 188.120 ;
        RECT 93.625 188.070 94.145 188.610 ;
        RECT 94.335 188.310 94.665 188.560 ;
        RECT 91.005 187.320 91.275 187.780 ;
        RECT 91.445 187.490 91.730 187.950 ;
        RECT 92.475 187.320 92.765 188.045 ;
        RECT 92.935 187.320 94.145 188.070 ;
        RECT 94.355 187.320 94.585 188.140 ;
        RECT 94.835 188.120 95.085 188.720 ;
        RECT 96.155 188.260 96.905 188.780 ;
        RECT 98.085 188.770 98.750 188.940 ;
        RECT 98.935 188.795 99.205 189.700 ;
        RECT 98.580 188.625 98.750 188.770 ;
        RECT 94.755 187.490 95.085 188.120 ;
        RECT 95.255 187.320 95.465 188.140 ;
        RECT 97.075 188.090 97.825 188.610 ;
        RECT 98.015 188.220 98.345 188.590 ;
        RECT 98.580 188.295 98.865 188.625 ;
        RECT 96.155 187.320 97.825 188.090 ;
        RECT 98.580 188.040 98.750 188.295 ;
        RECT 98.085 187.870 98.750 188.040 ;
        RECT 99.035 187.995 99.205 188.795 ;
        RECT 99.375 188.780 100.585 189.870 ;
        RECT 99.375 188.240 99.895 188.780 ;
        RECT 100.795 188.730 101.025 189.870 ;
        RECT 101.195 188.720 101.525 189.700 ;
        RECT 101.695 188.730 101.905 189.870 ;
        RECT 102.250 189.240 102.535 189.700 ;
        RECT 102.705 189.410 102.975 189.870 ;
        RECT 102.250 189.020 103.205 189.240 ;
        RECT 100.065 188.070 100.585 188.610 ;
        RECT 100.775 188.310 101.105 188.560 ;
        RECT 98.085 187.490 98.255 187.870 ;
        RECT 98.435 187.320 98.765 187.700 ;
        RECT 98.945 187.490 99.205 187.995 ;
        RECT 99.375 187.320 100.585 188.070 ;
        RECT 100.795 187.320 101.025 188.140 ;
        RECT 101.275 188.120 101.525 188.720 ;
        RECT 102.135 188.290 102.825 188.850 ;
        RECT 101.195 187.490 101.525 188.120 ;
        RECT 101.695 187.320 101.905 188.140 ;
        RECT 102.995 188.120 103.205 189.020 ;
        RECT 102.250 187.950 103.205 188.120 ;
        RECT 103.375 188.850 103.775 189.700 ;
        RECT 103.965 189.240 104.245 189.700 ;
        RECT 104.765 189.410 105.090 189.870 ;
        RECT 103.965 189.020 105.090 189.240 ;
        RECT 103.375 188.290 104.470 188.850 ;
        RECT 104.640 188.560 105.090 189.020 ;
        RECT 105.260 188.730 105.645 189.700 ;
        RECT 102.250 187.490 102.535 187.950 ;
        RECT 102.705 187.320 102.975 187.780 ;
        RECT 103.375 187.490 103.775 188.290 ;
        RECT 104.640 188.230 105.195 188.560 ;
        RECT 104.640 188.120 105.090 188.230 ;
        RECT 103.965 187.950 105.090 188.120 ;
        RECT 105.365 188.060 105.645 188.730 ;
        RECT 103.965 187.490 104.245 187.950 ;
        RECT 104.765 187.320 105.090 187.780 ;
        RECT 105.260 187.490 105.645 188.060 ;
        RECT 105.820 188.680 106.075 189.560 ;
        RECT 106.245 188.730 106.550 189.870 ;
        RECT 106.890 189.490 107.220 189.870 ;
        RECT 107.400 189.320 107.570 189.610 ;
        RECT 107.740 189.410 107.990 189.870 ;
        RECT 106.770 189.150 107.570 189.320 ;
        RECT 108.160 189.360 109.030 189.700 ;
        RECT 105.820 188.030 106.030 188.680 ;
        RECT 106.770 188.560 106.940 189.150 ;
        RECT 108.160 188.980 108.330 189.360 ;
        RECT 109.265 189.240 109.435 189.700 ;
        RECT 109.605 189.410 109.975 189.870 ;
        RECT 110.270 189.270 110.440 189.610 ;
        RECT 110.610 189.440 110.940 189.870 ;
        RECT 111.175 189.270 111.345 189.610 ;
        RECT 107.110 188.810 108.330 188.980 ;
        RECT 108.500 188.900 108.960 189.190 ;
        RECT 109.265 189.070 109.825 189.240 ;
        RECT 110.270 189.100 111.345 189.270 ;
        RECT 111.515 189.370 112.195 189.700 ;
        RECT 112.410 189.370 112.660 189.700 ;
        RECT 112.830 189.410 113.080 189.870 ;
        RECT 109.655 188.930 109.825 189.070 ;
        RECT 108.500 188.890 109.465 188.900 ;
        RECT 108.160 188.720 108.330 188.810 ;
        RECT 108.790 188.730 109.465 188.890 ;
        RECT 106.200 188.530 106.940 188.560 ;
        RECT 106.200 188.230 107.115 188.530 ;
        RECT 106.790 188.055 107.115 188.230 ;
        RECT 105.820 187.500 106.075 188.030 ;
        RECT 106.245 187.320 106.550 187.780 ;
        RECT 106.795 187.700 107.115 188.055 ;
        RECT 107.285 188.270 107.825 188.640 ;
        RECT 108.160 188.550 108.565 188.720 ;
        RECT 107.285 187.870 107.525 188.270 ;
        RECT 108.005 188.100 108.225 188.380 ;
        RECT 107.695 187.930 108.225 188.100 ;
        RECT 107.695 187.700 107.865 187.930 ;
        RECT 108.395 187.770 108.565 188.550 ;
        RECT 108.735 187.940 109.085 188.560 ;
        RECT 109.255 187.940 109.465 188.730 ;
        RECT 109.655 188.760 111.155 188.930 ;
        RECT 109.655 188.070 109.825 188.760 ;
        RECT 111.515 188.590 111.685 189.370 ;
        RECT 112.490 189.240 112.660 189.370 ;
        RECT 109.995 188.420 111.685 188.590 ;
        RECT 111.855 188.810 112.320 189.200 ;
        RECT 112.490 189.070 112.885 189.240 ;
        RECT 109.995 188.240 110.165 188.420 ;
        RECT 106.795 187.530 107.865 187.700 ;
        RECT 108.035 187.320 108.225 187.760 ;
        RECT 108.395 187.490 109.345 187.770 ;
        RECT 109.655 187.680 109.915 188.070 ;
        RECT 110.335 188.000 111.125 188.250 ;
        RECT 109.565 187.510 109.915 187.680 ;
        RECT 110.125 187.320 110.455 187.780 ;
        RECT 111.330 187.710 111.500 188.420 ;
        RECT 111.855 188.220 112.025 188.810 ;
        RECT 111.670 188.000 112.025 188.220 ;
        RECT 112.195 188.000 112.545 188.620 ;
        RECT 112.715 187.710 112.885 189.070 ;
        RECT 113.250 188.900 113.575 189.685 ;
        RECT 113.055 187.850 113.515 188.900 ;
        RECT 111.330 187.540 112.185 187.710 ;
        RECT 112.390 187.540 112.885 187.710 ;
        RECT 113.055 187.320 113.385 187.680 ;
        RECT 113.745 187.580 113.915 189.700 ;
        RECT 114.085 189.370 114.415 189.870 ;
        RECT 114.585 189.200 114.840 189.700 ;
        RECT 114.090 189.030 114.840 189.200 ;
        RECT 114.090 188.040 114.320 189.030 ;
        RECT 114.490 188.210 114.840 188.860 ;
        RECT 115.475 188.780 117.145 189.870 ;
        RECT 117.315 188.780 118.525 189.870 ;
        RECT 115.475 188.260 116.225 188.780 ;
        RECT 116.395 188.090 117.145 188.610 ;
        RECT 117.315 188.240 117.835 188.780 ;
        RECT 114.090 187.870 114.840 188.040 ;
        RECT 114.085 187.320 114.415 187.700 ;
        RECT 114.585 187.580 114.840 187.870 ;
        RECT 115.475 187.320 117.145 188.090 ;
        RECT 118.005 188.070 118.525 188.610 ;
        RECT 117.315 187.320 118.525 188.070 ;
        RECT 11.430 187.150 118.610 187.320 ;
        RECT 11.515 186.400 12.725 187.150 ;
        RECT 11.515 185.860 12.035 186.400 ;
        RECT 12.895 186.380 15.485 187.150 ;
        RECT 15.660 186.605 21.005 187.150 ;
        RECT 21.180 186.605 26.525 187.150 ;
        RECT 12.205 185.690 12.725 186.230 ;
        RECT 11.515 184.600 12.725 185.690 ;
        RECT 12.895 185.690 14.105 186.210 ;
        RECT 14.275 185.860 15.485 186.380 ;
        RECT 12.895 184.600 15.485 185.690 ;
        RECT 17.250 185.035 17.600 186.285 ;
        RECT 19.080 185.775 19.420 186.605 ;
        RECT 22.770 185.035 23.120 186.285 ;
        RECT 24.600 185.775 24.940 186.605 ;
        RECT 26.785 186.600 26.955 186.980 ;
        RECT 27.135 186.770 27.465 187.150 ;
        RECT 26.785 186.430 27.450 186.600 ;
        RECT 27.645 186.475 27.905 186.980 ;
        RECT 26.715 185.880 27.045 186.250 ;
        RECT 27.280 186.175 27.450 186.430 ;
        RECT 27.280 185.845 27.565 186.175 ;
        RECT 27.280 185.700 27.450 185.845 ;
        RECT 26.785 185.530 27.450 185.700 ;
        RECT 27.735 185.675 27.905 186.475 ;
        RECT 28.075 186.425 28.365 187.150 ;
        RECT 29.455 186.380 32.965 187.150 ;
        RECT 33.140 186.605 38.485 187.150 ;
        RECT 38.655 186.640 38.960 187.150 ;
        RECT 15.660 184.600 21.005 185.035 ;
        RECT 21.180 184.600 26.525 185.035 ;
        RECT 26.785 184.770 26.955 185.530 ;
        RECT 27.135 184.600 27.465 185.360 ;
        RECT 27.635 184.770 27.905 185.675 ;
        RECT 28.075 184.600 28.365 185.765 ;
        RECT 29.455 185.690 31.145 186.210 ;
        RECT 31.315 185.860 32.965 186.380 ;
        RECT 29.455 184.600 32.965 185.690 ;
        RECT 34.730 185.035 35.080 186.285 ;
        RECT 36.560 185.775 36.900 186.605 ;
        RECT 38.655 185.910 38.970 186.470 ;
        RECT 39.140 186.160 39.390 186.970 ;
        RECT 39.560 186.625 39.820 187.150 ;
        RECT 40.000 186.160 40.250 186.970 ;
        RECT 40.420 186.590 40.680 187.150 ;
        RECT 40.850 186.500 41.110 186.955 ;
        RECT 41.280 186.670 41.540 187.150 ;
        RECT 41.710 186.500 41.970 186.955 ;
        RECT 42.140 186.670 42.400 187.150 ;
        RECT 42.570 186.500 42.830 186.955 ;
        RECT 43.000 186.670 43.245 187.150 ;
        RECT 43.415 186.500 43.690 186.955 ;
        RECT 43.860 186.670 44.105 187.150 ;
        RECT 44.275 186.500 44.535 186.955 ;
        RECT 44.715 186.670 44.965 187.150 ;
        RECT 45.135 186.500 45.395 186.955 ;
        RECT 45.575 186.670 45.825 187.150 ;
        RECT 45.995 186.500 46.255 186.955 ;
        RECT 46.435 186.670 46.695 187.150 ;
        RECT 46.865 186.500 47.125 186.955 ;
        RECT 47.295 186.670 47.595 187.150 ;
        RECT 40.850 186.330 47.595 186.500 ;
        RECT 48.130 186.340 48.375 186.945 ;
        RECT 48.595 186.615 49.105 187.150 ;
        RECT 39.140 185.910 46.260 186.160 ;
        RECT 33.140 184.600 38.485 185.035 ;
        RECT 38.665 184.600 38.960 185.410 ;
        RECT 39.140 184.770 39.385 185.910 ;
        RECT 39.560 184.600 39.820 185.410 ;
        RECT 40.000 184.775 40.250 185.910 ;
        RECT 46.430 185.740 47.595 186.330 ;
        RECT 40.850 185.515 47.595 185.740 ;
        RECT 47.855 186.170 49.085 186.340 ;
        RECT 40.850 185.500 46.255 185.515 ;
        RECT 40.420 184.605 40.680 185.400 ;
        RECT 40.850 184.775 41.110 185.500 ;
        RECT 41.280 184.605 41.540 185.330 ;
        RECT 41.710 184.775 41.970 185.500 ;
        RECT 42.140 184.605 42.400 185.330 ;
        RECT 42.570 184.775 42.830 185.500 ;
        RECT 43.000 184.605 43.260 185.330 ;
        RECT 43.430 184.775 43.690 185.500 ;
        RECT 43.860 184.605 44.105 185.330 ;
        RECT 44.275 184.775 44.535 185.500 ;
        RECT 44.720 184.605 44.965 185.330 ;
        RECT 45.135 184.775 45.395 185.500 ;
        RECT 45.580 184.605 45.825 185.330 ;
        RECT 45.995 184.775 46.255 185.500 ;
        RECT 46.440 184.605 46.695 185.330 ;
        RECT 46.865 184.775 47.155 185.515 ;
        RECT 47.855 185.360 48.195 186.170 ;
        RECT 48.365 185.605 49.115 185.795 ;
        RECT 40.420 184.600 46.695 184.605 ;
        RECT 47.325 184.600 47.595 185.345 ;
        RECT 47.855 184.950 48.370 185.360 ;
        RECT 48.605 184.600 48.775 185.360 ;
        RECT 48.945 184.940 49.115 185.605 ;
        RECT 49.285 185.620 49.475 186.980 ;
        RECT 49.645 186.470 49.920 186.980 ;
        RECT 50.110 186.615 50.640 186.980 ;
        RECT 51.065 186.750 51.395 187.150 ;
        RECT 50.465 186.580 50.640 186.615 ;
        RECT 49.645 186.300 49.925 186.470 ;
        RECT 49.645 185.820 49.920 186.300 ;
        RECT 50.125 185.620 50.295 186.420 ;
        RECT 49.285 185.450 50.295 185.620 ;
        RECT 50.465 186.410 51.395 186.580 ;
        RECT 51.565 186.410 51.820 186.980 ;
        RECT 52.085 186.600 52.255 186.980 ;
        RECT 52.435 186.770 52.765 187.150 ;
        RECT 52.085 186.430 52.750 186.600 ;
        RECT 52.945 186.475 53.205 186.980 ;
        RECT 50.465 185.280 50.635 186.410 ;
        RECT 51.225 186.240 51.395 186.410 ;
        RECT 49.510 185.110 50.635 185.280 ;
        RECT 50.805 185.910 51.000 186.240 ;
        RECT 51.225 185.910 51.480 186.240 ;
        RECT 50.805 184.940 50.975 185.910 ;
        RECT 51.650 185.740 51.820 186.410 ;
        RECT 52.015 185.880 52.345 186.250 ;
        RECT 52.580 186.175 52.750 186.430 ;
        RECT 48.945 184.770 50.975 184.940 ;
        RECT 51.145 184.600 51.315 185.740 ;
        RECT 51.485 184.770 51.820 185.740 ;
        RECT 52.580 185.845 52.865 186.175 ;
        RECT 52.580 185.700 52.750 185.845 ;
        RECT 52.085 185.530 52.750 185.700 ;
        RECT 53.035 185.675 53.205 186.475 ;
        RECT 53.835 186.425 54.125 187.150 ;
        RECT 54.755 186.380 58.265 187.150 ;
        RECT 58.440 186.605 63.785 187.150 ;
        RECT 64.225 186.755 64.555 187.150 ;
        RECT 52.085 184.770 52.255 185.530 ;
        RECT 52.435 184.600 52.765 185.360 ;
        RECT 52.935 184.770 53.205 185.675 ;
        RECT 53.835 184.600 54.125 185.765 ;
        RECT 54.755 185.690 56.445 186.210 ;
        RECT 56.615 185.860 58.265 186.380 ;
        RECT 54.755 184.600 58.265 185.690 ;
        RECT 60.030 185.035 60.380 186.285 ;
        RECT 61.860 185.775 62.200 186.605 ;
        RECT 64.725 186.580 64.925 186.935 ;
        RECT 65.095 186.750 65.425 187.150 ;
        RECT 65.595 186.580 65.795 186.925 ;
        RECT 63.955 186.410 65.795 186.580 ;
        RECT 65.965 186.410 66.295 187.150 ;
        RECT 66.530 186.580 66.700 186.830 ;
        RECT 66.530 186.410 67.005 186.580 ;
        RECT 58.440 184.600 63.785 185.035 ;
        RECT 63.955 184.785 64.215 186.410 ;
        RECT 64.395 185.440 64.615 186.240 ;
        RECT 64.855 185.620 65.155 186.240 ;
        RECT 65.325 185.620 65.655 186.240 ;
        RECT 65.825 185.620 66.145 186.240 ;
        RECT 66.315 185.620 66.665 186.240 ;
        RECT 66.835 185.440 67.005 186.410 ;
        RECT 67.725 186.500 67.895 186.980 ;
        RECT 68.075 186.670 68.315 187.150 ;
        RECT 68.565 186.500 68.735 186.980 ;
        RECT 68.905 186.670 69.235 187.150 ;
        RECT 69.405 186.500 69.575 186.980 ;
        RECT 67.725 186.330 68.360 186.500 ;
        RECT 68.565 186.330 69.575 186.500 ;
        RECT 69.745 186.350 70.075 187.150 ;
        RECT 70.400 186.440 70.655 186.970 ;
        RECT 70.825 186.690 71.130 187.150 ;
        RECT 71.375 186.770 72.445 186.940 ;
        RECT 68.190 186.160 68.360 186.330 ;
        RECT 67.640 185.920 68.020 186.160 ;
        RECT 68.190 185.990 68.690 186.160 ;
        RECT 68.190 185.750 68.360 185.990 ;
        RECT 69.080 185.790 69.575 186.330 ;
        RECT 64.395 185.230 67.005 185.440 ;
        RECT 67.645 185.580 68.360 185.750 ;
        RECT 68.565 185.620 69.575 185.790 ;
        RECT 70.400 185.790 70.610 186.440 ;
        RECT 71.375 186.415 71.695 186.770 ;
        RECT 71.370 186.240 71.695 186.415 ;
        RECT 70.780 185.940 71.695 186.240 ;
        RECT 71.865 186.200 72.105 186.600 ;
        RECT 72.275 186.540 72.445 186.770 ;
        RECT 72.615 186.710 72.805 187.150 ;
        RECT 72.975 186.700 73.925 186.980 ;
        RECT 74.145 186.790 74.495 186.960 ;
        RECT 72.275 186.370 72.805 186.540 ;
        RECT 70.780 185.910 71.520 185.940 ;
        RECT 65.965 184.600 66.295 185.050 ;
        RECT 67.645 184.770 67.975 185.580 ;
        RECT 68.145 184.600 68.385 185.400 ;
        RECT 68.565 184.770 68.735 185.620 ;
        RECT 68.905 184.600 69.235 185.400 ;
        RECT 69.405 184.770 69.575 185.620 ;
        RECT 69.745 184.600 70.075 185.750 ;
        RECT 70.400 184.910 70.655 185.790 ;
        RECT 70.825 184.600 71.130 185.740 ;
        RECT 71.350 185.320 71.520 185.910 ;
        RECT 71.865 185.830 72.405 186.200 ;
        RECT 72.585 186.090 72.805 186.370 ;
        RECT 72.975 185.920 73.145 186.700 ;
        RECT 72.740 185.750 73.145 185.920 ;
        RECT 73.315 185.910 73.665 186.530 ;
        RECT 72.740 185.660 72.910 185.750 ;
        RECT 73.835 185.740 74.045 186.530 ;
        RECT 71.690 185.490 72.910 185.660 ;
        RECT 73.370 185.580 74.045 185.740 ;
        RECT 71.350 185.150 72.150 185.320 ;
        RECT 71.470 184.600 71.800 184.980 ;
        RECT 71.980 184.860 72.150 185.150 ;
        RECT 72.740 185.110 72.910 185.490 ;
        RECT 73.080 185.570 74.045 185.580 ;
        RECT 74.235 186.400 74.495 186.790 ;
        RECT 74.705 186.690 75.035 187.150 ;
        RECT 75.910 186.760 76.765 186.930 ;
        RECT 76.970 186.760 77.465 186.930 ;
        RECT 77.635 186.790 77.965 187.150 ;
        RECT 74.235 185.710 74.405 186.400 ;
        RECT 74.575 186.050 74.745 186.230 ;
        RECT 74.915 186.220 75.705 186.470 ;
        RECT 75.910 186.050 76.080 186.760 ;
        RECT 76.250 186.250 76.605 186.470 ;
        RECT 74.575 185.880 76.265 186.050 ;
        RECT 73.080 185.280 73.540 185.570 ;
        RECT 74.235 185.540 75.735 185.710 ;
        RECT 74.235 185.400 74.405 185.540 ;
        RECT 73.845 185.230 74.405 185.400 ;
        RECT 72.320 184.600 72.570 185.060 ;
        RECT 72.740 184.770 73.610 185.110 ;
        RECT 73.845 184.770 74.015 185.230 ;
        RECT 74.850 185.200 75.925 185.370 ;
        RECT 74.185 184.600 74.555 185.060 ;
        RECT 74.850 184.860 75.020 185.200 ;
        RECT 75.190 184.600 75.520 185.030 ;
        RECT 75.755 184.860 75.925 185.200 ;
        RECT 76.095 185.100 76.265 185.880 ;
        RECT 76.435 185.660 76.605 186.250 ;
        RECT 76.775 185.850 77.125 186.470 ;
        RECT 76.435 185.270 76.900 185.660 ;
        RECT 77.295 185.400 77.465 186.760 ;
        RECT 77.635 185.570 78.095 186.620 ;
        RECT 77.070 185.230 77.465 185.400 ;
        RECT 77.070 185.100 77.240 185.230 ;
        RECT 76.095 184.770 76.775 185.100 ;
        RECT 76.990 184.770 77.240 185.100 ;
        RECT 77.410 184.600 77.660 185.060 ;
        RECT 77.830 184.785 78.155 185.570 ;
        RECT 78.325 184.770 78.495 186.890 ;
        RECT 78.665 186.770 78.995 187.150 ;
        RECT 79.165 186.600 79.420 186.890 ;
        RECT 78.670 186.430 79.420 186.600 ;
        RECT 78.670 185.440 78.900 186.430 ;
        RECT 79.595 186.425 79.885 187.150 ;
        RECT 80.060 186.440 80.315 186.970 ;
        RECT 80.485 186.690 80.790 187.150 ;
        RECT 81.035 186.770 82.105 186.940 ;
        RECT 79.070 185.610 79.420 186.260 ;
        RECT 80.060 185.790 80.270 186.440 ;
        RECT 81.035 186.415 81.355 186.770 ;
        RECT 81.030 186.240 81.355 186.415 ;
        RECT 80.440 185.940 81.355 186.240 ;
        RECT 81.525 186.200 81.765 186.600 ;
        RECT 81.935 186.540 82.105 186.770 ;
        RECT 82.275 186.710 82.465 187.150 ;
        RECT 82.635 186.700 83.585 186.980 ;
        RECT 83.805 186.790 84.155 186.960 ;
        RECT 81.935 186.370 82.465 186.540 ;
        RECT 80.440 185.910 81.180 185.940 ;
        RECT 78.670 185.270 79.420 185.440 ;
        RECT 78.665 184.600 78.995 185.100 ;
        RECT 79.165 184.770 79.420 185.270 ;
        RECT 79.595 184.600 79.885 185.765 ;
        RECT 80.060 184.910 80.315 185.790 ;
        RECT 80.485 184.600 80.790 185.740 ;
        RECT 81.010 185.320 81.180 185.910 ;
        RECT 81.525 185.830 82.065 186.200 ;
        RECT 82.245 186.090 82.465 186.370 ;
        RECT 82.635 185.920 82.805 186.700 ;
        RECT 82.400 185.750 82.805 185.920 ;
        RECT 82.975 185.910 83.325 186.530 ;
        RECT 82.400 185.660 82.570 185.750 ;
        RECT 83.495 185.740 83.705 186.530 ;
        RECT 81.350 185.490 82.570 185.660 ;
        RECT 83.030 185.580 83.705 185.740 ;
        RECT 81.010 185.150 81.810 185.320 ;
        RECT 81.130 184.600 81.460 184.980 ;
        RECT 81.640 184.860 81.810 185.150 ;
        RECT 82.400 185.110 82.570 185.490 ;
        RECT 82.740 185.570 83.705 185.580 ;
        RECT 83.895 186.400 84.155 186.790 ;
        RECT 84.365 186.690 84.695 187.150 ;
        RECT 85.570 186.760 86.425 186.930 ;
        RECT 86.630 186.760 87.125 186.930 ;
        RECT 87.295 186.790 87.625 187.150 ;
        RECT 83.895 185.710 84.065 186.400 ;
        RECT 84.235 186.050 84.405 186.230 ;
        RECT 84.575 186.220 85.365 186.470 ;
        RECT 85.570 186.050 85.740 186.760 ;
        RECT 85.910 186.250 86.265 186.470 ;
        RECT 84.235 185.880 85.925 186.050 ;
        RECT 82.740 185.280 83.200 185.570 ;
        RECT 83.895 185.540 85.395 185.710 ;
        RECT 83.895 185.400 84.065 185.540 ;
        RECT 83.505 185.230 84.065 185.400 ;
        RECT 81.980 184.600 82.230 185.060 ;
        RECT 82.400 184.770 83.270 185.110 ;
        RECT 83.505 184.770 83.675 185.230 ;
        RECT 84.510 185.200 85.585 185.370 ;
        RECT 83.845 184.600 84.215 185.060 ;
        RECT 84.510 184.860 84.680 185.200 ;
        RECT 84.850 184.600 85.180 185.030 ;
        RECT 85.415 184.860 85.585 185.200 ;
        RECT 85.755 185.100 85.925 185.880 ;
        RECT 86.095 185.660 86.265 186.250 ;
        RECT 86.435 185.850 86.785 186.470 ;
        RECT 86.095 185.270 86.560 185.660 ;
        RECT 86.955 185.400 87.125 186.760 ;
        RECT 87.295 185.570 87.755 186.620 ;
        RECT 86.730 185.230 87.125 185.400 ;
        RECT 86.730 185.100 86.900 185.230 ;
        RECT 85.755 184.770 86.435 185.100 ;
        RECT 86.650 184.770 86.900 185.100 ;
        RECT 87.070 184.600 87.320 185.060 ;
        RECT 87.490 184.785 87.815 185.570 ;
        RECT 87.985 184.770 88.155 186.890 ;
        RECT 88.325 186.770 88.655 187.150 ;
        RECT 88.825 186.600 89.080 186.890 ;
        RECT 88.330 186.430 89.080 186.600 ;
        RECT 88.330 185.440 88.560 186.430 ;
        RECT 90.175 186.380 93.685 187.150 ;
        RECT 93.860 186.605 99.205 187.150 ;
        RECT 88.730 185.610 89.080 186.260 ;
        RECT 90.175 185.690 91.865 186.210 ;
        RECT 92.035 185.860 93.685 186.380 ;
        RECT 88.330 185.270 89.080 185.440 ;
        RECT 88.325 184.600 88.655 185.100 ;
        RECT 88.825 184.770 89.080 185.270 ;
        RECT 90.175 184.600 93.685 185.690 ;
        RECT 95.450 185.035 95.800 186.285 ;
        RECT 97.280 185.775 97.620 186.605 ;
        RECT 99.435 186.330 99.645 187.150 ;
        RECT 99.815 186.350 100.145 186.980 ;
        RECT 99.815 185.750 100.065 186.350 ;
        RECT 100.315 186.330 100.545 187.150 ;
        RECT 101.490 186.340 101.735 186.945 ;
        RECT 101.955 186.615 102.465 187.150 ;
        RECT 101.215 186.170 102.445 186.340 ;
        RECT 100.235 185.910 100.565 186.160 ;
        RECT 93.860 184.600 99.205 185.035 ;
        RECT 99.435 184.600 99.645 185.740 ;
        RECT 99.815 184.770 100.145 185.750 ;
        RECT 100.315 184.600 100.545 185.740 ;
        RECT 101.215 185.360 101.555 186.170 ;
        RECT 101.725 185.605 102.475 185.795 ;
        RECT 101.215 184.950 101.730 185.360 ;
        RECT 101.965 184.600 102.135 185.360 ;
        RECT 102.305 184.940 102.475 185.605 ;
        RECT 102.645 185.620 102.835 186.980 ;
        RECT 103.005 186.470 103.280 186.980 ;
        RECT 103.470 186.615 104.000 186.980 ;
        RECT 104.425 186.750 104.755 187.150 ;
        RECT 103.825 186.580 104.000 186.615 ;
        RECT 103.005 186.300 103.285 186.470 ;
        RECT 103.005 185.820 103.280 186.300 ;
        RECT 103.485 185.620 103.655 186.420 ;
        RECT 102.645 185.450 103.655 185.620 ;
        RECT 103.825 186.410 104.755 186.580 ;
        RECT 104.925 186.410 105.180 186.980 ;
        RECT 105.355 186.425 105.645 187.150 ;
        RECT 105.820 186.440 106.075 186.970 ;
        RECT 106.245 186.690 106.550 187.150 ;
        RECT 106.795 186.770 107.865 186.940 ;
        RECT 103.825 185.280 103.995 186.410 ;
        RECT 104.585 186.240 104.755 186.410 ;
        RECT 102.870 185.110 103.995 185.280 ;
        RECT 104.165 185.910 104.360 186.240 ;
        RECT 104.585 185.910 104.840 186.240 ;
        RECT 104.165 184.940 104.335 185.910 ;
        RECT 105.010 185.740 105.180 186.410 ;
        RECT 105.820 185.790 106.030 186.440 ;
        RECT 106.795 186.415 107.115 186.770 ;
        RECT 106.790 186.240 107.115 186.415 ;
        RECT 106.200 185.940 107.115 186.240 ;
        RECT 107.285 186.200 107.525 186.600 ;
        RECT 107.695 186.540 107.865 186.770 ;
        RECT 108.035 186.710 108.225 187.150 ;
        RECT 108.395 186.700 109.345 186.980 ;
        RECT 109.565 186.790 109.915 186.960 ;
        RECT 107.695 186.370 108.225 186.540 ;
        RECT 106.200 185.910 106.940 185.940 ;
        RECT 102.305 184.770 104.335 184.940 ;
        RECT 104.505 184.600 104.675 185.740 ;
        RECT 104.845 184.770 105.180 185.740 ;
        RECT 105.355 184.600 105.645 185.765 ;
        RECT 105.820 184.910 106.075 185.790 ;
        RECT 106.245 184.600 106.550 185.740 ;
        RECT 106.770 185.320 106.940 185.910 ;
        RECT 107.285 185.830 107.825 186.200 ;
        RECT 108.005 186.090 108.225 186.370 ;
        RECT 108.395 185.920 108.565 186.700 ;
        RECT 108.160 185.750 108.565 185.920 ;
        RECT 108.735 185.910 109.085 186.530 ;
        RECT 108.160 185.660 108.330 185.750 ;
        RECT 109.255 185.740 109.465 186.530 ;
        RECT 107.110 185.490 108.330 185.660 ;
        RECT 108.790 185.580 109.465 185.740 ;
        RECT 106.770 185.150 107.570 185.320 ;
        RECT 106.890 184.600 107.220 184.980 ;
        RECT 107.400 184.860 107.570 185.150 ;
        RECT 108.160 185.110 108.330 185.490 ;
        RECT 108.500 185.570 109.465 185.580 ;
        RECT 109.655 186.400 109.915 186.790 ;
        RECT 110.125 186.690 110.455 187.150 ;
        RECT 111.330 186.760 112.185 186.930 ;
        RECT 112.390 186.760 112.885 186.930 ;
        RECT 113.055 186.790 113.385 187.150 ;
        RECT 109.655 185.710 109.825 186.400 ;
        RECT 109.995 186.050 110.165 186.230 ;
        RECT 110.335 186.220 111.125 186.470 ;
        RECT 111.330 186.050 111.500 186.760 ;
        RECT 111.670 186.250 112.025 186.470 ;
        RECT 109.995 185.880 111.685 186.050 ;
        RECT 108.500 185.280 108.960 185.570 ;
        RECT 109.655 185.540 111.155 185.710 ;
        RECT 109.655 185.400 109.825 185.540 ;
        RECT 109.265 185.230 109.825 185.400 ;
        RECT 107.740 184.600 107.990 185.060 ;
        RECT 108.160 184.770 109.030 185.110 ;
        RECT 109.265 184.770 109.435 185.230 ;
        RECT 110.270 185.200 111.345 185.370 ;
        RECT 109.605 184.600 109.975 185.060 ;
        RECT 110.270 184.860 110.440 185.200 ;
        RECT 110.610 184.600 110.940 185.030 ;
        RECT 111.175 184.860 111.345 185.200 ;
        RECT 111.515 185.100 111.685 185.880 ;
        RECT 111.855 185.660 112.025 186.250 ;
        RECT 112.195 185.850 112.545 186.470 ;
        RECT 111.855 185.270 112.320 185.660 ;
        RECT 112.715 185.400 112.885 186.760 ;
        RECT 113.055 185.570 113.515 186.620 ;
        RECT 112.490 185.230 112.885 185.400 ;
        RECT 112.490 185.100 112.660 185.230 ;
        RECT 111.515 184.770 112.195 185.100 ;
        RECT 112.410 184.770 112.660 185.100 ;
        RECT 112.830 184.600 113.080 185.060 ;
        RECT 113.250 184.785 113.575 185.570 ;
        RECT 113.745 184.770 113.915 186.890 ;
        RECT 114.085 186.770 114.415 187.150 ;
        RECT 114.585 186.600 114.840 186.890 ;
        RECT 114.090 186.430 114.840 186.600 ;
        RECT 115.015 186.475 115.275 186.980 ;
        RECT 115.455 186.770 115.785 187.150 ;
        RECT 115.965 186.600 116.135 186.980 ;
        RECT 114.090 185.440 114.320 186.430 ;
        RECT 114.490 185.610 114.840 186.260 ;
        RECT 115.015 185.675 115.185 186.475 ;
        RECT 115.470 186.430 116.135 186.600 ;
        RECT 115.470 186.175 115.640 186.430 ;
        RECT 117.315 186.400 118.525 187.150 ;
        RECT 115.355 185.845 115.640 186.175 ;
        RECT 115.875 185.880 116.205 186.250 ;
        RECT 115.470 185.700 115.640 185.845 ;
        RECT 114.090 185.270 114.840 185.440 ;
        RECT 114.085 184.600 114.415 185.100 ;
        RECT 114.585 184.770 114.840 185.270 ;
        RECT 115.015 184.770 115.285 185.675 ;
        RECT 115.470 185.530 116.135 185.700 ;
        RECT 115.455 184.600 115.785 185.360 ;
        RECT 115.965 184.770 116.135 185.530 ;
        RECT 117.315 185.690 117.835 186.230 ;
        RECT 118.005 185.860 118.525 186.400 ;
        RECT 117.315 184.600 118.525 185.690 ;
        RECT 11.430 184.430 118.610 184.600 ;
        RECT 11.515 183.340 12.725 184.430 ;
        RECT 11.515 182.630 12.035 183.170 ;
        RECT 12.205 182.800 12.725 183.340 ;
        RECT 13.355 183.340 15.025 184.430 ;
        RECT 13.355 182.820 14.105 183.340 ;
        RECT 15.195 183.265 15.485 184.430 ;
        RECT 16.115 183.340 18.705 184.430 ;
        RECT 18.880 183.995 24.225 184.430 ;
        RECT 14.275 182.650 15.025 183.170 ;
        RECT 16.115 182.820 17.325 183.340 ;
        RECT 17.495 182.650 18.705 183.170 ;
        RECT 20.470 182.745 20.820 183.995 ;
        RECT 11.515 181.880 12.725 182.630 ;
        RECT 13.355 181.880 15.025 182.650 ;
        RECT 15.195 181.880 15.485 182.605 ;
        RECT 16.115 181.880 18.705 182.650 ;
        RECT 22.300 182.425 22.640 183.255 ;
        RECT 24.400 183.240 24.655 184.120 ;
        RECT 24.825 183.290 25.130 184.430 ;
        RECT 25.470 184.050 25.800 184.430 ;
        RECT 25.980 183.880 26.150 184.170 ;
        RECT 26.320 183.970 26.570 184.430 ;
        RECT 25.350 183.710 26.150 183.880 ;
        RECT 26.740 183.920 27.610 184.260 ;
        RECT 24.400 182.590 24.610 183.240 ;
        RECT 25.350 183.120 25.520 183.710 ;
        RECT 26.740 183.540 26.910 183.920 ;
        RECT 27.845 183.800 28.015 184.260 ;
        RECT 28.185 183.970 28.555 184.430 ;
        RECT 28.850 183.830 29.020 184.170 ;
        RECT 29.190 184.000 29.520 184.430 ;
        RECT 29.755 183.830 29.925 184.170 ;
        RECT 25.690 183.370 26.910 183.540 ;
        RECT 27.080 183.460 27.540 183.750 ;
        RECT 27.845 183.630 28.405 183.800 ;
        RECT 28.850 183.660 29.925 183.830 ;
        RECT 30.095 183.930 30.775 184.260 ;
        RECT 30.990 183.930 31.240 184.260 ;
        RECT 31.410 183.970 31.660 184.430 ;
        RECT 28.235 183.490 28.405 183.630 ;
        RECT 27.080 183.450 28.045 183.460 ;
        RECT 26.740 183.280 26.910 183.370 ;
        RECT 27.370 183.290 28.045 183.450 ;
        RECT 24.780 183.090 25.520 183.120 ;
        RECT 24.780 182.790 25.695 183.090 ;
        RECT 25.370 182.615 25.695 182.790 ;
        RECT 18.880 181.880 24.225 182.425 ;
        RECT 24.400 182.060 24.655 182.590 ;
        RECT 24.825 181.880 25.130 182.340 ;
        RECT 25.375 182.260 25.695 182.615 ;
        RECT 25.865 182.830 26.405 183.200 ;
        RECT 26.740 183.110 27.145 183.280 ;
        RECT 25.865 182.430 26.105 182.830 ;
        RECT 26.585 182.660 26.805 182.940 ;
        RECT 26.275 182.490 26.805 182.660 ;
        RECT 26.275 182.260 26.445 182.490 ;
        RECT 26.975 182.330 27.145 183.110 ;
        RECT 27.315 182.500 27.665 183.120 ;
        RECT 27.835 182.500 28.045 183.290 ;
        RECT 28.235 183.320 29.735 183.490 ;
        RECT 28.235 182.630 28.405 183.320 ;
        RECT 30.095 183.150 30.265 183.930 ;
        RECT 31.070 183.800 31.240 183.930 ;
        RECT 28.575 182.980 30.265 183.150 ;
        RECT 30.435 183.370 30.900 183.760 ;
        RECT 31.070 183.630 31.465 183.800 ;
        RECT 28.575 182.800 28.745 182.980 ;
        RECT 25.375 182.090 26.445 182.260 ;
        RECT 26.615 181.880 26.805 182.320 ;
        RECT 26.975 182.050 27.925 182.330 ;
        RECT 28.235 182.240 28.495 182.630 ;
        RECT 28.915 182.560 29.705 182.810 ;
        RECT 28.145 182.070 28.495 182.240 ;
        RECT 28.705 181.880 29.035 182.340 ;
        RECT 29.910 182.270 30.080 182.980 ;
        RECT 30.435 182.780 30.605 183.370 ;
        RECT 30.250 182.560 30.605 182.780 ;
        RECT 30.775 182.560 31.125 183.180 ;
        RECT 31.295 182.270 31.465 183.630 ;
        RECT 31.830 183.460 32.155 184.245 ;
        RECT 31.635 182.410 32.095 183.460 ;
        RECT 29.910 182.100 30.765 182.270 ;
        RECT 30.970 182.100 31.465 182.270 ;
        RECT 31.635 181.880 31.965 182.240 ;
        RECT 32.325 182.140 32.495 184.260 ;
        RECT 32.665 183.930 32.995 184.430 ;
        RECT 33.165 183.760 33.420 184.260 ;
        RECT 32.670 183.590 33.420 183.760 ;
        RECT 32.670 182.600 32.900 183.590 ;
        RECT 33.070 182.770 33.420 183.420 ;
        RECT 34.055 183.340 36.645 184.430 ;
        RECT 36.815 183.670 37.330 184.080 ;
        RECT 37.565 183.670 37.735 184.430 ;
        RECT 37.905 184.090 39.935 184.260 ;
        RECT 34.055 182.820 35.265 183.340 ;
        RECT 35.435 182.650 36.645 183.170 ;
        RECT 36.815 182.860 37.155 183.670 ;
        RECT 37.905 183.425 38.075 184.090 ;
        RECT 38.470 183.750 39.595 183.920 ;
        RECT 37.325 183.235 38.075 183.425 ;
        RECT 38.245 183.410 39.255 183.580 ;
        RECT 36.815 182.690 38.045 182.860 ;
        RECT 32.670 182.430 33.420 182.600 ;
        RECT 32.665 181.880 32.995 182.260 ;
        RECT 33.165 182.140 33.420 182.430 ;
        RECT 34.055 181.880 36.645 182.650 ;
        RECT 37.090 182.085 37.335 182.690 ;
        RECT 37.555 181.880 38.065 182.415 ;
        RECT 38.245 182.050 38.435 183.410 ;
        RECT 38.605 182.390 38.880 183.210 ;
        RECT 39.085 182.610 39.255 183.410 ;
        RECT 39.425 182.620 39.595 183.750 ;
        RECT 39.765 183.120 39.935 184.090 ;
        RECT 40.105 183.290 40.275 184.430 ;
        RECT 40.445 183.290 40.780 184.260 ;
        RECT 39.765 182.790 39.960 183.120 ;
        RECT 40.185 182.790 40.440 183.120 ;
        RECT 40.185 182.620 40.355 182.790 ;
        RECT 40.610 182.620 40.780 183.290 ;
        RECT 40.955 183.265 41.245 184.430 ;
        RECT 41.415 183.355 41.685 184.260 ;
        RECT 41.855 183.670 42.185 184.430 ;
        RECT 42.365 183.500 42.535 184.260 ;
        RECT 39.425 182.450 40.355 182.620 ;
        RECT 39.425 182.415 39.600 182.450 ;
        RECT 38.605 182.220 38.885 182.390 ;
        RECT 38.605 182.050 38.880 182.220 ;
        RECT 39.070 182.050 39.600 182.415 ;
        RECT 40.025 181.880 40.355 182.280 ;
        RECT 40.525 182.050 40.780 182.620 ;
        RECT 40.955 181.880 41.245 182.605 ;
        RECT 41.415 182.555 41.585 183.355 ;
        RECT 41.870 183.330 42.535 183.500 ;
        RECT 41.870 183.185 42.040 183.330 ;
        RECT 42.855 183.290 43.065 184.430 ;
        RECT 41.755 182.855 42.040 183.185 ;
        RECT 43.235 183.280 43.565 184.260 ;
        RECT 43.735 183.290 43.965 184.430 ;
        RECT 44.235 183.595 44.490 184.430 ;
        RECT 44.660 183.425 44.920 184.230 ;
        RECT 45.090 183.595 45.350 184.430 ;
        RECT 45.520 183.425 45.775 184.230 ;
        RECT 41.870 182.600 42.040 182.855 ;
        RECT 42.275 182.780 42.605 183.150 ;
        RECT 41.415 182.050 41.675 182.555 ;
        RECT 41.870 182.430 42.535 182.600 ;
        RECT 41.855 181.880 42.185 182.260 ;
        RECT 42.365 182.050 42.535 182.430 ;
        RECT 42.855 181.880 43.065 182.700 ;
        RECT 43.235 182.680 43.485 183.280 ;
        RECT 44.175 183.255 45.775 183.425 ;
        RECT 46.390 183.450 46.645 184.120 ;
        RECT 46.825 183.630 47.110 184.430 ;
        RECT 47.290 183.710 47.620 184.220 ;
        RECT 43.655 182.870 43.985 183.120 ;
        RECT 43.235 182.050 43.565 182.680 ;
        RECT 43.735 181.880 43.965 182.700 ;
        RECT 44.175 182.690 44.455 183.255 ;
        RECT 44.625 182.860 45.845 183.085 ;
        RECT 44.175 182.520 44.905 182.690 ;
        RECT 44.180 181.880 44.510 182.350 ;
        RECT 44.680 182.075 44.905 182.520 ;
        RECT 46.390 182.590 46.570 183.450 ;
        RECT 47.290 183.120 47.540 183.710 ;
        RECT 47.890 183.560 48.060 184.170 ;
        RECT 48.230 183.740 48.560 184.430 ;
        RECT 48.790 183.880 49.030 184.170 ;
        RECT 49.230 184.050 49.650 184.430 ;
        RECT 49.830 183.960 50.460 184.210 ;
        RECT 50.930 184.050 51.260 184.430 ;
        RECT 49.830 183.880 50.000 183.960 ;
        RECT 51.430 183.880 51.600 184.170 ;
        RECT 51.780 184.050 52.160 184.430 ;
        RECT 52.400 184.045 53.230 184.215 ;
        RECT 48.790 183.710 50.000 183.880 ;
        RECT 46.740 182.790 47.540 183.120 ;
        RECT 45.075 181.880 45.370 182.405 ;
        RECT 46.390 182.390 46.645 182.590 ;
        RECT 46.305 182.220 46.645 182.390 ;
        RECT 46.390 182.060 46.645 182.220 ;
        RECT 46.825 181.880 47.110 182.340 ;
        RECT 47.290 182.140 47.540 182.790 ;
        RECT 47.740 183.540 48.060 183.560 ;
        RECT 47.740 183.370 49.660 183.540 ;
        RECT 47.740 182.475 47.930 183.370 ;
        RECT 49.830 183.200 50.000 183.710 ;
        RECT 50.170 183.450 50.690 183.760 ;
        RECT 48.100 183.030 50.000 183.200 ;
        RECT 48.100 182.970 48.430 183.030 ;
        RECT 48.580 182.800 48.910 182.860 ;
        RECT 48.250 182.530 48.910 182.800 ;
        RECT 47.740 182.145 48.060 182.475 ;
        RECT 48.240 181.880 48.900 182.360 ;
        RECT 49.100 182.270 49.270 183.030 ;
        RECT 50.170 182.860 50.350 183.270 ;
        RECT 49.440 182.690 49.770 182.810 ;
        RECT 50.520 182.690 50.690 183.450 ;
        RECT 49.440 182.520 50.690 182.690 ;
        RECT 50.860 183.630 52.230 183.880 ;
        RECT 50.860 182.860 51.050 183.630 ;
        RECT 51.980 183.370 52.230 183.630 ;
        RECT 51.220 183.200 51.470 183.360 ;
        RECT 52.400 183.200 52.570 184.045 ;
        RECT 53.465 183.760 53.635 184.260 ;
        RECT 53.805 183.930 54.135 184.430 ;
        RECT 52.740 183.370 53.240 183.750 ;
        RECT 53.465 183.590 54.160 183.760 ;
        RECT 51.220 183.030 52.570 183.200 ;
        RECT 52.150 182.990 52.570 183.030 ;
        RECT 50.860 182.520 51.280 182.860 ;
        RECT 51.570 182.530 51.980 182.860 ;
        RECT 49.100 182.100 49.950 182.270 ;
        RECT 50.510 181.880 50.830 182.340 ;
        RECT 51.030 182.090 51.280 182.520 ;
        RECT 51.570 181.880 51.980 182.320 ;
        RECT 52.150 182.260 52.320 182.990 ;
        RECT 52.490 182.440 52.840 182.810 ;
        RECT 53.020 182.500 53.240 183.370 ;
        RECT 53.410 182.800 53.820 183.420 ;
        RECT 53.990 182.620 54.160 183.590 ;
        RECT 53.465 182.430 54.160 182.620 ;
        RECT 52.150 182.060 53.165 182.260 ;
        RECT 53.465 182.100 53.635 182.430 ;
        RECT 53.805 181.880 54.135 182.260 ;
        RECT 54.350 182.140 54.575 184.260 ;
        RECT 54.745 183.930 55.075 184.430 ;
        RECT 55.245 183.760 55.415 184.260 ;
        RECT 54.750 183.590 55.415 183.760 ;
        RECT 54.750 182.600 54.980 183.590 ;
        RECT 55.150 182.770 55.500 183.420 ;
        RECT 56.135 183.340 58.725 184.430 ;
        RECT 59.605 183.980 59.935 184.430 ;
        RECT 58.895 183.590 61.505 183.800 ;
        RECT 56.135 182.820 57.345 183.340 ;
        RECT 57.515 182.650 58.725 183.170 ;
        RECT 54.750 182.430 55.415 182.600 ;
        RECT 54.745 181.880 55.075 182.260 ;
        RECT 55.245 182.140 55.415 182.430 ;
        RECT 56.135 181.880 58.725 182.650 ;
        RECT 58.895 182.620 59.065 183.590 ;
        RECT 59.235 182.790 59.585 183.410 ;
        RECT 59.755 182.790 60.075 183.410 ;
        RECT 60.245 182.790 60.575 183.410 ;
        RECT 60.745 182.790 61.045 183.410 ;
        RECT 61.285 182.790 61.505 183.590 ;
        RECT 61.685 182.620 61.945 184.245 ;
        RECT 58.895 182.450 59.370 182.620 ;
        RECT 59.200 182.200 59.370 182.450 ;
        RECT 59.605 181.880 59.935 182.620 ;
        RECT 60.105 182.450 61.945 182.620 ;
        RECT 62.115 183.930 62.375 184.260 ;
        RECT 62.685 184.050 63.015 184.430 ;
        RECT 62.115 183.250 62.285 183.930 ;
        RECT 63.255 183.880 63.445 184.260 ;
        RECT 63.695 184.050 64.025 184.430 ;
        RECT 64.235 183.880 64.405 184.260 ;
        RECT 64.600 184.050 64.930 184.430 ;
        RECT 65.190 183.880 65.360 184.260 ;
        RECT 65.785 184.050 66.115 184.430 ;
        RECT 62.455 183.420 62.805 183.750 ;
        RECT 63.255 183.710 63.995 183.880 ;
        RECT 63.075 183.370 63.655 183.540 ;
        RECT 63.075 183.250 63.245 183.370 ;
        RECT 62.115 183.080 63.245 183.250 ;
        RECT 63.825 183.200 63.995 183.710 ;
        RECT 60.105 182.105 60.305 182.450 ;
        RECT 60.475 181.880 60.805 182.280 ;
        RECT 60.975 182.095 61.175 182.450 ;
        RECT 62.115 182.380 62.285 183.080 ;
        RECT 63.425 183.030 63.995 183.200 ;
        RECT 64.165 183.710 66.115 183.880 ;
        RECT 62.635 182.740 63.255 182.910 ;
        RECT 62.635 182.560 62.845 182.740 ;
        RECT 63.425 182.550 63.595 183.030 ;
        RECT 64.165 182.720 64.335 183.710 ;
        RECT 64.925 183.120 65.110 183.430 ;
        RECT 65.380 183.120 65.575 183.430 ;
        RECT 61.345 181.880 61.675 182.275 ;
        RECT 62.115 182.050 62.375 182.380 ;
        RECT 62.685 181.880 63.015 182.260 ;
        RECT 63.195 182.220 63.595 182.550 ;
        RECT 63.785 182.390 64.335 182.720 ;
        RECT 64.505 182.220 64.675 183.120 ;
        RECT 63.195 182.050 64.675 182.220 ;
        RECT 64.925 182.790 65.155 183.120 ;
        RECT 65.380 182.790 65.635 183.120 ;
        RECT 65.945 182.790 66.115 183.710 ;
        RECT 64.925 182.210 65.110 182.790 ;
        RECT 65.380 182.215 65.575 182.790 ;
        RECT 65.785 181.880 66.115 182.260 ;
        RECT 66.285 182.050 66.545 184.260 ;
        RECT 66.715 183.265 67.005 184.430 ;
        RECT 67.175 182.620 67.435 184.245 ;
        RECT 69.185 183.980 69.515 184.430 ;
        RECT 67.615 183.590 70.225 183.800 ;
        RECT 67.615 182.790 67.835 183.590 ;
        RECT 68.075 182.790 68.375 183.410 ;
        RECT 68.545 182.790 68.875 183.410 ;
        RECT 69.045 182.790 69.365 183.410 ;
        RECT 69.535 182.790 69.885 183.410 ;
        RECT 70.055 182.620 70.225 183.590 ;
        RECT 70.395 183.340 71.605 184.430 ;
        RECT 71.775 183.670 72.290 184.080 ;
        RECT 72.525 183.670 72.695 184.430 ;
        RECT 72.865 184.090 74.895 184.260 ;
        RECT 70.395 182.800 70.915 183.340 ;
        RECT 71.085 182.630 71.605 183.170 ;
        RECT 71.775 182.860 72.115 183.670 ;
        RECT 72.865 183.425 73.035 184.090 ;
        RECT 73.430 183.750 74.555 183.920 ;
        RECT 72.285 183.235 73.035 183.425 ;
        RECT 73.205 183.410 74.215 183.580 ;
        RECT 71.775 182.690 73.005 182.860 ;
        RECT 66.715 181.880 67.005 182.605 ;
        RECT 67.175 182.450 69.015 182.620 ;
        RECT 67.445 181.880 67.775 182.275 ;
        RECT 67.945 182.095 68.145 182.450 ;
        RECT 68.315 181.880 68.645 182.280 ;
        RECT 68.815 182.105 69.015 182.450 ;
        RECT 69.185 181.880 69.515 182.620 ;
        RECT 69.750 182.450 70.225 182.620 ;
        RECT 69.750 182.200 69.920 182.450 ;
        RECT 70.395 181.880 71.605 182.630 ;
        RECT 72.050 182.085 72.295 182.690 ;
        RECT 72.515 181.880 73.025 182.415 ;
        RECT 73.205 182.050 73.395 183.410 ;
        RECT 73.565 182.390 73.840 183.210 ;
        RECT 74.045 182.610 74.215 183.410 ;
        RECT 74.385 182.620 74.555 183.750 ;
        RECT 74.725 183.120 74.895 184.090 ;
        RECT 75.065 183.290 75.235 184.430 ;
        RECT 75.405 183.290 75.740 184.260 ;
        RECT 76.005 183.685 76.275 184.430 ;
        RECT 76.905 184.425 83.180 184.430 ;
        RECT 76.445 183.515 76.735 184.255 ;
        RECT 76.905 183.700 77.160 184.425 ;
        RECT 77.345 183.530 77.605 184.255 ;
        RECT 77.775 183.700 78.020 184.425 ;
        RECT 78.205 183.530 78.465 184.255 ;
        RECT 78.635 183.700 78.880 184.425 ;
        RECT 79.065 183.530 79.325 184.255 ;
        RECT 79.495 183.700 79.740 184.425 ;
        RECT 79.910 183.530 80.170 184.255 ;
        RECT 80.340 183.700 80.600 184.425 ;
        RECT 80.770 183.530 81.030 184.255 ;
        RECT 81.200 183.700 81.460 184.425 ;
        RECT 81.630 183.530 81.890 184.255 ;
        RECT 82.060 183.700 82.320 184.425 ;
        RECT 82.490 183.530 82.750 184.255 ;
        RECT 82.920 183.630 83.180 184.425 ;
        RECT 77.345 183.515 82.750 183.530 ;
        RECT 74.725 182.790 74.920 183.120 ;
        RECT 75.145 182.790 75.400 183.120 ;
        RECT 75.145 182.620 75.315 182.790 ;
        RECT 75.570 182.620 75.740 183.290 ;
        RECT 74.385 182.450 75.315 182.620 ;
        RECT 74.385 182.415 74.560 182.450 ;
        RECT 73.565 182.220 73.845 182.390 ;
        RECT 73.565 182.050 73.840 182.220 ;
        RECT 74.030 182.050 74.560 182.415 ;
        RECT 74.985 181.880 75.315 182.280 ;
        RECT 75.485 182.050 75.740 182.620 ;
        RECT 76.005 183.290 82.750 183.515 ;
        RECT 76.005 182.700 77.170 183.290 ;
        RECT 83.350 183.120 83.600 184.255 ;
        RECT 83.780 183.620 84.040 184.430 ;
        RECT 84.215 183.120 84.460 184.260 ;
        RECT 84.640 183.620 84.935 184.430 ;
        RECT 85.575 183.340 87.245 184.430 ;
        RECT 87.415 183.355 87.685 184.260 ;
        RECT 87.855 183.670 88.185 184.430 ;
        RECT 88.365 183.500 88.535 184.260 ;
        RECT 77.340 182.870 84.460 183.120 ;
        RECT 76.005 182.530 82.750 182.700 ;
        RECT 76.005 181.880 76.305 182.360 ;
        RECT 76.475 182.075 76.735 182.530 ;
        RECT 76.905 181.880 77.165 182.360 ;
        RECT 77.345 182.075 77.605 182.530 ;
        RECT 77.775 181.880 78.025 182.360 ;
        RECT 78.205 182.075 78.465 182.530 ;
        RECT 78.635 181.880 78.885 182.360 ;
        RECT 79.065 182.075 79.325 182.530 ;
        RECT 79.495 181.880 79.740 182.360 ;
        RECT 79.910 182.075 80.185 182.530 ;
        RECT 80.355 181.880 80.600 182.360 ;
        RECT 80.770 182.075 81.030 182.530 ;
        RECT 81.200 181.880 81.460 182.360 ;
        RECT 81.630 182.075 81.890 182.530 ;
        RECT 82.060 181.880 82.320 182.360 ;
        RECT 82.490 182.075 82.750 182.530 ;
        RECT 82.920 181.880 83.180 182.440 ;
        RECT 83.350 182.060 83.600 182.870 ;
        RECT 83.780 181.880 84.040 182.405 ;
        RECT 84.210 182.060 84.460 182.870 ;
        RECT 84.630 182.560 84.945 183.120 ;
        RECT 85.575 182.820 86.325 183.340 ;
        RECT 86.495 182.650 87.245 183.170 ;
        RECT 84.640 181.880 84.945 182.390 ;
        RECT 85.575 181.880 87.245 182.650 ;
        RECT 87.415 182.555 87.585 183.355 ;
        RECT 87.870 183.330 88.535 183.500 ;
        RECT 87.870 183.185 88.040 183.330 ;
        RECT 89.315 183.290 89.525 184.430 ;
        RECT 87.755 182.855 88.040 183.185 ;
        RECT 89.695 183.280 90.025 184.260 ;
        RECT 90.195 183.290 90.425 184.430 ;
        RECT 91.185 183.500 91.355 184.260 ;
        RECT 91.535 183.670 91.865 184.430 ;
        RECT 91.185 183.330 91.850 183.500 ;
        RECT 92.035 183.355 92.305 184.260 ;
        RECT 87.870 182.600 88.040 182.855 ;
        RECT 88.275 182.780 88.605 183.150 ;
        RECT 87.415 182.050 87.675 182.555 ;
        RECT 87.870 182.430 88.535 182.600 ;
        RECT 87.855 181.880 88.185 182.260 ;
        RECT 88.365 182.050 88.535 182.430 ;
        RECT 89.315 181.880 89.525 182.700 ;
        RECT 89.695 182.680 89.945 183.280 ;
        RECT 91.680 183.185 91.850 183.330 ;
        RECT 90.115 182.870 90.445 183.120 ;
        RECT 91.115 182.780 91.445 183.150 ;
        RECT 91.680 182.855 91.965 183.185 ;
        RECT 89.695 182.050 90.025 182.680 ;
        RECT 90.195 181.880 90.425 182.700 ;
        RECT 91.680 182.600 91.850 182.855 ;
        RECT 91.185 182.430 91.850 182.600 ;
        RECT 92.135 182.555 92.305 183.355 ;
        RECT 92.475 183.265 92.765 184.430 ;
        RECT 93.140 183.460 93.470 184.260 ;
        RECT 93.640 183.630 93.970 184.430 ;
        RECT 94.270 183.460 94.600 184.260 ;
        RECT 95.245 183.630 95.495 184.430 ;
        RECT 93.140 183.290 95.575 183.460 ;
        RECT 95.765 183.290 95.935 184.430 ;
        RECT 96.105 183.290 96.445 184.260 ;
        RECT 92.935 182.870 93.285 183.120 ;
        RECT 93.470 182.660 93.640 183.290 ;
        RECT 93.810 182.870 94.140 183.070 ;
        RECT 94.310 182.870 94.640 183.070 ;
        RECT 94.810 182.870 95.230 183.070 ;
        RECT 95.405 183.040 95.575 183.290 ;
        RECT 96.215 183.240 96.445 183.290 ;
        RECT 95.405 182.870 96.100 183.040 ;
        RECT 91.185 182.050 91.355 182.430 ;
        RECT 91.535 181.880 91.865 182.260 ;
        RECT 92.045 182.050 92.305 182.555 ;
        RECT 92.475 181.880 92.765 182.605 ;
        RECT 93.140 182.050 93.640 182.660 ;
        RECT 94.270 182.530 95.495 182.700 ;
        RECT 96.270 182.680 96.445 183.240 ;
        RECT 94.270 182.050 94.600 182.530 ;
        RECT 94.770 181.880 94.995 182.340 ;
        RECT 95.165 182.050 95.495 182.530 ;
        RECT 95.685 181.880 95.935 182.680 ;
        RECT 96.105 182.050 96.445 182.680 ;
        RECT 96.620 183.240 96.875 184.120 ;
        RECT 97.045 183.290 97.350 184.430 ;
        RECT 97.690 184.050 98.020 184.430 ;
        RECT 98.200 183.880 98.370 184.170 ;
        RECT 98.540 183.970 98.790 184.430 ;
        RECT 97.570 183.710 98.370 183.880 ;
        RECT 98.960 183.920 99.830 184.260 ;
        RECT 96.620 182.590 96.830 183.240 ;
        RECT 97.570 183.120 97.740 183.710 ;
        RECT 98.960 183.540 99.130 183.920 ;
        RECT 100.065 183.800 100.235 184.260 ;
        RECT 100.405 183.970 100.775 184.430 ;
        RECT 101.070 183.830 101.240 184.170 ;
        RECT 101.410 184.000 101.740 184.430 ;
        RECT 101.975 183.830 102.145 184.170 ;
        RECT 97.910 183.370 99.130 183.540 ;
        RECT 99.300 183.460 99.760 183.750 ;
        RECT 100.065 183.630 100.625 183.800 ;
        RECT 101.070 183.660 102.145 183.830 ;
        RECT 102.315 183.930 102.995 184.260 ;
        RECT 103.210 183.930 103.460 184.260 ;
        RECT 103.630 183.970 103.880 184.430 ;
        RECT 100.455 183.490 100.625 183.630 ;
        RECT 99.300 183.450 100.265 183.460 ;
        RECT 98.960 183.280 99.130 183.370 ;
        RECT 99.590 183.290 100.265 183.450 ;
        RECT 97.000 183.090 97.740 183.120 ;
        RECT 97.000 182.790 97.915 183.090 ;
        RECT 97.590 182.615 97.915 182.790 ;
        RECT 96.620 182.060 96.875 182.590 ;
        RECT 97.045 181.880 97.350 182.340 ;
        RECT 97.595 182.260 97.915 182.615 ;
        RECT 98.085 182.830 98.625 183.200 ;
        RECT 98.960 183.110 99.365 183.280 ;
        RECT 98.085 182.430 98.325 182.830 ;
        RECT 98.805 182.660 99.025 182.940 ;
        RECT 98.495 182.490 99.025 182.660 ;
        RECT 98.495 182.260 98.665 182.490 ;
        RECT 99.195 182.330 99.365 183.110 ;
        RECT 99.535 182.500 99.885 183.120 ;
        RECT 100.055 182.500 100.265 183.290 ;
        RECT 100.455 183.320 101.955 183.490 ;
        RECT 100.455 182.630 100.625 183.320 ;
        RECT 102.315 183.150 102.485 183.930 ;
        RECT 103.290 183.800 103.460 183.930 ;
        RECT 100.795 182.980 102.485 183.150 ;
        RECT 102.655 183.370 103.120 183.760 ;
        RECT 103.290 183.630 103.685 183.800 ;
        RECT 100.795 182.800 100.965 182.980 ;
        RECT 97.595 182.090 98.665 182.260 ;
        RECT 98.835 181.880 99.025 182.320 ;
        RECT 99.195 182.050 100.145 182.330 ;
        RECT 100.455 182.240 100.715 182.630 ;
        RECT 101.135 182.560 101.925 182.810 ;
        RECT 100.365 182.070 100.715 182.240 ;
        RECT 100.925 181.880 101.255 182.340 ;
        RECT 102.130 182.270 102.300 182.980 ;
        RECT 102.655 182.780 102.825 183.370 ;
        RECT 102.470 182.560 102.825 182.780 ;
        RECT 102.995 182.560 103.345 183.180 ;
        RECT 103.515 182.270 103.685 183.630 ;
        RECT 104.050 183.460 104.375 184.245 ;
        RECT 103.855 182.410 104.315 183.460 ;
        RECT 102.130 182.100 102.985 182.270 ;
        RECT 103.190 182.100 103.685 182.270 ;
        RECT 103.855 181.880 104.185 182.240 ;
        RECT 104.545 182.140 104.715 184.260 ;
        RECT 104.885 183.930 105.215 184.430 ;
        RECT 105.385 183.760 105.640 184.260 ;
        RECT 104.890 183.590 105.640 183.760 ;
        RECT 105.815 183.670 106.330 184.080 ;
        RECT 106.565 183.670 106.735 184.430 ;
        RECT 106.905 184.090 108.935 184.260 ;
        RECT 104.890 182.600 105.120 183.590 ;
        RECT 105.290 182.770 105.640 183.420 ;
        RECT 105.815 182.860 106.155 183.670 ;
        RECT 106.905 183.425 107.075 184.090 ;
        RECT 107.470 183.750 108.595 183.920 ;
        RECT 106.325 183.235 107.075 183.425 ;
        RECT 107.245 183.410 108.255 183.580 ;
        RECT 105.815 182.690 107.045 182.860 ;
        RECT 104.890 182.430 105.640 182.600 ;
        RECT 104.885 181.880 105.215 182.260 ;
        RECT 105.385 182.140 105.640 182.430 ;
        RECT 106.090 182.085 106.335 182.690 ;
        RECT 106.555 181.880 107.065 182.415 ;
        RECT 107.245 182.050 107.435 183.410 ;
        RECT 107.605 182.390 107.880 183.210 ;
        RECT 108.085 182.610 108.255 183.410 ;
        RECT 108.425 182.620 108.595 183.750 ;
        RECT 108.765 183.120 108.935 184.090 ;
        RECT 109.105 183.290 109.275 184.430 ;
        RECT 109.445 183.290 109.780 184.260 ;
        RECT 110.965 183.500 111.135 184.260 ;
        RECT 111.315 183.670 111.645 184.430 ;
        RECT 110.965 183.330 111.630 183.500 ;
        RECT 111.815 183.355 112.085 184.260 ;
        RECT 108.765 182.790 108.960 183.120 ;
        RECT 109.185 182.790 109.440 183.120 ;
        RECT 109.185 182.620 109.355 182.790 ;
        RECT 109.610 182.620 109.780 183.290 ;
        RECT 111.460 183.185 111.630 183.330 ;
        RECT 110.895 182.780 111.225 183.150 ;
        RECT 111.460 182.855 111.745 183.185 ;
        RECT 108.425 182.450 109.355 182.620 ;
        RECT 108.425 182.415 108.600 182.450 ;
        RECT 107.605 182.220 107.885 182.390 ;
        RECT 107.605 182.050 107.880 182.220 ;
        RECT 108.070 182.050 108.600 182.415 ;
        RECT 109.025 181.880 109.355 182.280 ;
        RECT 109.525 182.050 109.780 182.620 ;
        RECT 111.460 182.600 111.630 182.855 ;
        RECT 110.965 182.430 111.630 182.600 ;
        RECT 111.915 182.555 112.085 183.355 ;
        RECT 112.255 183.340 113.465 184.430 ;
        RECT 113.635 183.340 117.145 184.430 ;
        RECT 117.315 183.340 118.525 184.430 ;
        RECT 112.255 182.800 112.775 183.340 ;
        RECT 112.945 182.630 113.465 183.170 ;
        RECT 113.635 182.820 115.325 183.340 ;
        RECT 115.495 182.650 117.145 183.170 ;
        RECT 117.315 182.800 117.835 183.340 ;
        RECT 110.965 182.050 111.135 182.430 ;
        RECT 111.315 181.880 111.645 182.260 ;
        RECT 111.825 182.050 112.085 182.555 ;
        RECT 112.255 181.880 113.465 182.630 ;
        RECT 113.635 181.880 117.145 182.650 ;
        RECT 118.005 182.630 118.525 183.170 ;
        RECT 117.315 181.880 118.525 182.630 ;
        RECT 11.430 181.710 118.610 181.880 ;
        RECT 11.515 180.960 12.725 181.710 ;
        RECT 11.515 180.420 12.035 180.960 ;
        RECT 13.355 180.940 15.945 181.710 ;
        RECT 12.205 180.250 12.725 180.790 ;
        RECT 11.515 179.160 12.725 180.250 ;
        RECT 13.355 180.250 14.565 180.770 ;
        RECT 14.735 180.420 15.945 180.940 ;
        RECT 16.155 180.890 16.385 181.710 ;
        RECT 16.555 180.910 16.885 181.540 ;
        RECT 16.135 180.470 16.465 180.720 ;
        RECT 16.635 180.310 16.885 180.910 ;
        RECT 17.055 180.890 17.265 181.710 ;
        RECT 17.500 181.000 17.755 181.530 ;
        RECT 17.925 181.250 18.230 181.710 ;
        RECT 18.475 181.330 19.545 181.500 ;
        RECT 13.355 179.160 15.945 180.250 ;
        RECT 16.155 179.160 16.385 180.300 ;
        RECT 16.555 179.330 16.885 180.310 ;
        RECT 17.500 180.350 17.710 181.000 ;
        RECT 18.475 180.975 18.795 181.330 ;
        RECT 18.470 180.800 18.795 180.975 ;
        RECT 17.880 180.500 18.795 180.800 ;
        RECT 18.965 180.760 19.205 181.160 ;
        RECT 19.375 181.100 19.545 181.330 ;
        RECT 19.715 181.270 19.905 181.710 ;
        RECT 20.075 181.260 21.025 181.540 ;
        RECT 21.245 181.350 21.595 181.520 ;
        RECT 19.375 180.930 19.905 181.100 ;
        RECT 17.880 180.470 18.620 180.500 ;
        RECT 17.055 179.160 17.265 180.300 ;
        RECT 17.500 179.470 17.755 180.350 ;
        RECT 17.925 179.160 18.230 180.300 ;
        RECT 18.450 179.880 18.620 180.470 ;
        RECT 18.965 180.390 19.505 180.760 ;
        RECT 19.685 180.650 19.905 180.930 ;
        RECT 20.075 180.480 20.245 181.260 ;
        RECT 19.840 180.310 20.245 180.480 ;
        RECT 20.415 180.470 20.765 181.090 ;
        RECT 19.840 180.220 20.010 180.310 ;
        RECT 20.935 180.300 21.145 181.090 ;
        RECT 18.790 180.050 20.010 180.220 ;
        RECT 20.470 180.140 21.145 180.300 ;
        RECT 18.450 179.710 19.250 179.880 ;
        RECT 18.570 179.160 18.900 179.540 ;
        RECT 19.080 179.420 19.250 179.710 ;
        RECT 19.840 179.670 20.010 180.050 ;
        RECT 20.180 180.130 21.145 180.140 ;
        RECT 21.335 180.960 21.595 181.350 ;
        RECT 21.805 181.250 22.135 181.710 ;
        RECT 23.010 181.320 23.865 181.490 ;
        RECT 24.070 181.320 24.565 181.490 ;
        RECT 24.735 181.350 25.065 181.710 ;
        RECT 21.335 180.270 21.505 180.960 ;
        RECT 21.675 180.610 21.845 180.790 ;
        RECT 22.015 180.780 22.805 181.030 ;
        RECT 23.010 180.610 23.180 181.320 ;
        RECT 23.350 180.810 23.705 181.030 ;
        RECT 21.675 180.440 23.365 180.610 ;
        RECT 20.180 179.840 20.640 180.130 ;
        RECT 21.335 180.100 22.835 180.270 ;
        RECT 21.335 179.960 21.505 180.100 ;
        RECT 20.945 179.790 21.505 179.960 ;
        RECT 19.420 179.160 19.670 179.620 ;
        RECT 19.840 179.330 20.710 179.670 ;
        RECT 20.945 179.330 21.115 179.790 ;
        RECT 21.950 179.760 23.025 179.930 ;
        RECT 21.285 179.160 21.655 179.620 ;
        RECT 21.950 179.420 22.120 179.760 ;
        RECT 22.290 179.160 22.620 179.590 ;
        RECT 22.855 179.420 23.025 179.760 ;
        RECT 23.195 179.660 23.365 180.440 ;
        RECT 23.535 180.220 23.705 180.810 ;
        RECT 23.875 180.410 24.225 181.030 ;
        RECT 23.535 179.830 24.000 180.220 ;
        RECT 24.395 179.960 24.565 181.320 ;
        RECT 24.735 180.130 25.195 181.180 ;
        RECT 24.170 179.790 24.565 179.960 ;
        RECT 24.170 179.660 24.340 179.790 ;
        RECT 23.195 179.330 23.875 179.660 ;
        RECT 24.090 179.330 24.340 179.660 ;
        RECT 24.510 179.160 24.760 179.620 ;
        RECT 24.930 179.345 25.255 180.130 ;
        RECT 25.425 179.330 25.595 181.450 ;
        RECT 25.765 181.330 26.095 181.710 ;
        RECT 26.265 181.160 26.520 181.450 ;
        RECT 25.770 180.990 26.520 181.160 ;
        RECT 26.695 181.035 26.955 181.540 ;
        RECT 27.135 181.330 27.465 181.710 ;
        RECT 27.645 181.160 27.815 181.540 ;
        RECT 25.770 180.000 26.000 180.990 ;
        RECT 26.170 180.170 26.520 180.820 ;
        RECT 26.695 180.235 26.865 181.035 ;
        RECT 27.150 180.990 27.815 181.160 ;
        RECT 27.150 180.735 27.320 180.990 ;
        RECT 28.075 180.985 28.365 181.710 ;
        RECT 28.810 180.900 29.055 181.505 ;
        RECT 29.275 181.175 29.785 181.710 ;
        RECT 27.035 180.405 27.320 180.735 ;
        RECT 27.555 180.440 27.885 180.810 ;
        RECT 28.535 180.730 29.765 180.900 ;
        RECT 27.150 180.260 27.320 180.405 ;
        RECT 25.770 179.830 26.520 180.000 ;
        RECT 25.765 179.160 26.095 179.660 ;
        RECT 26.265 179.330 26.520 179.830 ;
        RECT 26.695 179.330 26.965 180.235 ;
        RECT 27.150 180.090 27.815 180.260 ;
        RECT 27.135 179.160 27.465 179.920 ;
        RECT 27.645 179.330 27.815 180.090 ;
        RECT 28.075 179.160 28.365 180.325 ;
        RECT 28.535 179.920 28.875 180.730 ;
        RECT 29.045 180.165 29.795 180.355 ;
        RECT 28.535 179.510 29.050 179.920 ;
        RECT 29.285 179.160 29.455 179.920 ;
        RECT 29.625 179.500 29.795 180.165 ;
        RECT 29.965 180.180 30.155 181.540 ;
        RECT 30.325 180.690 30.600 181.540 ;
        RECT 30.790 181.175 31.320 181.540 ;
        RECT 31.745 181.310 32.075 181.710 ;
        RECT 31.145 181.140 31.320 181.175 ;
        RECT 30.325 180.520 30.605 180.690 ;
        RECT 30.325 180.380 30.600 180.520 ;
        RECT 30.805 180.180 30.975 180.980 ;
        RECT 29.965 180.010 30.975 180.180 ;
        RECT 31.145 180.970 32.075 181.140 ;
        RECT 32.245 180.970 32.500 181.540 ;
        RECT 31.145 179.840 31.315 180.970 ;
        RECT 31.905 180.800 32.075 180.970 ;
        RECT 30.190 179.670 31.315 179.840 ;
        RECT 31.485 180.470 31.680 180.800 ;
        RECT 31.905 180.470 32.160 180.800 ;
        RECT 31.485 179.500 31.655 180.470 ;
        RECT 32.330 180.300 32.500 180.970 ;
        RECT 29.625 179.330 31.655 179.500 ;
        RECT 31.825 179.160 31.995 180.300 ;
        RECT 32.165 179.330 32.500 180.300 ;
        RECT 32.675 181.035 32.935 181.540 ;
        RECT 33.115 181.330 33.445 181.710 ;
        RECT 33.625 181.160 33.795 181.540 ;
        RECT 32.675 180.235 32.845 181.035 ;
        RECT 33.130 180.990 33.795 181.160 ;
        RECT 33.130 180.735 33.300 180.990 ;
        RECT 34.515 180.940 37.105 181.710 ;
        RECT 37.365 181.160 37.535 181.450 ;
        RECT 37.705 181.330 38.035 181.710 ;
        RECT 37.365 180.990 38.030 181.160 ;
        RECT 33.015 180.405 33.300 180.735 ;
        RECT 33.535 180.440 33.865 180.810 ;
        RECT 33.130 180.260 33.300 180.405 ;
        RECT 32.675 179.330 32.945 180.235 ;
        RECT 33.130 180.090 33.795 180.260 ;
        RECT 33.115 179.160 33.445 179.920 ;
        RECT 33.625 179.330 33.795 180.090 ;
        RECT 34.515 180.250 35.725 180.770 ;
        RECT 35.895 180.420 37.105 180.940 ;
        RECT 34.515 179.160 37.105 180.250 ;
        RECT 37.280 180.170 37.630 180.820 ;
        RECT 37.800 180.000 38.030 180.990 ;
        RECT 37.365 179.830 38.030 180.000 ;
        RECT 37.365 179.330 37.535 179.830 ;
        RECT 37.705 179.160 38.035 179.660 ;
        RECT 38.205 179.330 38.430 181.450 ;
        RECT 38.645 181.330 38.975 181.710 ;
        RECT 39.145 181.160 39.315 181.490 ;
        RECT 39.615 181.330 40.630 181.530 ;
        RECT 38.620 180.970 39.315 181.160 ;
        RECT 38.620 180.000 38.790 180.970 ;
        RECT 38.960 180.170 39.370 180.790 ;
        RECT 39.540 180.220 39.760 181.090 ;
        RECT 39.940 180.780 40.290 181.150 ;
        RECT 40.460 180.600 40.630 181.330 ;
        RECT 40.800 181.270 41.210 181.710 ;
        RECT 41.500 181.070 41.750 181.500 ;
        RECT 41.950 181.250 42.270 181.710 ;
        RECT 42.830 181.320 43.680 181.490 ;
        RECT 40.800 180.730 41.210 181.060 ;
        RECT 41.500 180.730 41.920 181.070 ;
        RECT 40.210 180.560 40.630 180.600 ;
        RECT 40.210 180.390 41.560 180.560 ;
        RECT 38.620 179.830 39.315 180.000 ;
        RECT 39.540 179.840 40.040 180.220 ;
        RECT 38.645 179.160 38.975 179.660 ;
        RECT 39.145 179.330 39.315 179.830 ;
        RECT 40.210 179.545 40.380 180.390 ;
        RECT 41.310 180.230 41.560 180.390 ;
        RECT 40.550 179.960 40.800 180.220 ;
        RECT 41.730 179.960 41.920 180.730 ;
        RECT 40.550 179.710 41.920 179.960 ;
        RECT 42.090 180.900 43.340 181.070 ;
        RECT 42.090 180.140 42.260 180.900 ;
        RECT 43.010 180.780 43.340 180.900 ;
        RECT 42.430 180.320 42.610 180.730 ;
        RECT 43.510 180.560 43.680 181.320 ;
        RECT 43.880 181.230 44.540 181.710 ;
        RECT 44.720 181.115 45.040 181.445 ;
        RECT 43.870 180.790 44.530 181.060 ;
        RECT 43.870 180.730 44.200 180.790 ;
        RECT 44.350 180.560 44.680 180.620 ;
        RECT 42.780 180.390 44.680 180.560 ;
        RECT 42.090 179.830 42.610 180.140 ;
        RECT 42.780 179.880 42.950 180.390 ;
        RECT 44.850 180.220 45.040 181.115 ;
        RECT 43.120 180.050 45.040 180.220 ;
        RECT 44.720 180.030 45.040 180.050 ;
        RECT 45.240 180.800 45.490 181.450 ;
        RECT 45.670 181.250 45.955 181.710 ;
        RECT 46.135 181.370 46.390 181.530 ;
        RECT 46.135 181.200 46.475 181.370 ;
        RECT 46.135 181.000 46.390 181.200 ;
        RECT 45.240 180.470 46.040 180.800 ;
        RECT 42.780 179.710 43.990 179.880 ;
        RECT 39.550 179.375 40.380 179.545 ;
        RECT 40.620 179.160 41.000 179.540 ;
        RECT 41.180 179.420 41.350 179.710 ;
        RECT 42.780 179.630 42.950 179.710 ;
        RECT 41.520 179.160 41.850 179.540 ;
        RECT 42.320 179.380 42.950 179.630 ;
        RECT 43.130 179.160 43.550 179.540 ;
        RECT 43.750 179.420 43.990 179.710 ;
        RECT 44.220 179.160 44.550 179.850 ;
        RECT 44.720 179.420 44.890 180.030 ;
        RECT 45.240 179.880 45.490 180.470 ;
        RECT 46.210 180.140 46.390 181.000 ;
        RECT 47.670 180.900 47.915 181.505 ;
        RECT 48.135 181.175 48.645 181.710 ;
        RECT 45.160 179.370 45.490 179.880 ;
        RECT 45.670 179.160 45.955 179.960 ;
        RECT 46.135 179.470 46.390 180.140 ;
        RECT 47.395 180.730 48.625 180.900 ;
        RECT 47.395 179.920 47.735 180.730 ;
        RECT 47.905 180.165 48.655 180.355 ;
        RECT 47.395 179.510 47.910 179.920 ;
        RECT 48.145 179.160 48.315 179.920 ;
        RECT 48.485 179.500 48.655 180.165 ;
        RECT 48.825 180.180 49.015 181.540 ;
        RECT 49.185 181.030 49.460 181.540 ;
        RECT 49.650 181.175 50.180 181.540 ;
        RECT 50.605 181.310 50.935 181.710 ;
        RECT 50.005 181.140 50.180 181.175 ;
        RECT 49.185 180.860 49.465 181.030 ;
        RECT 49.185 180.380 49.460 180.860 ;
        RECT 49.665 180.180 49.835 180.980 ;
        RECT 48.825 180.010 49.835 180.180 ;
        RECT 50.005 180.970 50.935 181.140 ;
        RECT 51.105 180.970 51.360 181.540 ;
        RECT 50.005 179.840 50.175 180.970 ;
        RECT 50.765 180.800 50.935 180.970 ;
        RECT 49.050 179.670 50.175 179.840 ;
        RECT 50.345 180.470 50.540 180.800 ;
        RECT 50.765 180.470 51.020 180.800 ;
        RECT 50.345 179.500 50.515 180.470 ;
        RECT 51.190 180.300 51.360 180.970 ;
        RECT 51.995 180.940 53.665 181.710 ;
        RECT 53.835 180.985 54.125 181.710 ;
        RECT 54.295 180.940 56.885 181.710 ;
        RECT 48.485 179.330 50.515 179.500 ;
        RECT 50.685 179.160 50.855 180.300 ;
        RECT 51.025 179.330 51.360 180.300 ;
        RECT 51.995 180.250 52.745 180.770 ;
        RECT 52.915 180.420 53.665 180.940 ;
        RECT 51.995 179.160 53.665 180.250 ;
        RECT 53.835 179.160 54.125 180.325 ;
        RECT 54.295 180.250 55.505 180.770 ;
        RECT 55.675 180.420 56.885 180.940 ;
        RECT 57.060 180.870 57.320 181.710 ;
        RECT 57.495 180.965 57.750 181.540 ;
        RECT 57.920 181.330 58.250 181.710 ;
        RECT 58.465 181.160 58.635 181.540 ;
        RECT 57.920 180.990 58.635 181.160 ;
        RECT 54.295 179.160 56.885 180.250 ;
        RECT 57.060 179.160 57.320 180.310 ;
        RECT 57.495 180.235 57.665 180.965 ;
        RECT 57.920 180.800 58.090 180.990 ;
        RECT 58.895 180.940 62.405 181.710 ;
        RECT 57.835 180.470 58.090 180.800 ;
        RECT 57.920 180.260 58.090 180.470 ;
        RECT 58.370 180.440 58.725 180.810 ;
        RECT 57.495 179.330 57.750 180.235 ;
        RECT 57.920 180.090 58.635 180.260 ;
        RECT 57.920 179.160 58.250 179.920 ;
        RECT 58.465 179.330 58.635 180.090 ;
        RECT 58.895 180.250 60.585 180.770 ;
        RECT 60.755 180.420 62.405 180.940 ;
        RECT 62.615 180.890 62.845 181.710 ;
        RECT 63.015 180.910 63.345 181.540 ;
        RECT 62.595 180.470 62.925 180.720 ;
        RECT 63.095 180.310 63.345 180.910 ;
        RECT 63.515 180.890 63.725 181.710 ;
        RECT 64.260 181.140 64.430 181.390 ;
        RECT 63.955 180.970 64.430 181.140 ;
        RECT 64.665 180.970 64.995 181.710 ;
        RECT 65.165 181.140 65.365 181.485 ;
        RECT 65.535 181.310 65.865 181.710 ;
        RECT 66.035 181.140 66.235 181.495 ;
        RECT 66.405 181.315 66.735 181.710 ;
        RECT 65.165 180.970 67.005 181.140 ;
        RECT 58.895 179.160 62.405 180.250 ;
        RECT 62.615 179.160 62.845 180.300 ;
        RECT 63.015 179.330 63.345 180.310 ;
        RECT 63.515 179.160 63.725 180.300 ;
        RECT 63.955 180.000 64.125 180.970 ;
        RECT 64.295 180.180 64.645 180.800 ;
        RECT 64.815 180.180 65.135 180.800 ;
        RECT 65.305 180.180 65.635 180.800 ;
        RECT 65.805 180.180 66.105 180.800 ;
        RECT 66.345 180.000 66.565 180.800 ;
        RECT 63.955 179.790 66.565 180.000 ;
        RECT 64.665 179.160 64.995 179.610 ;
        RECT 66.745 179.345 67.005 180.970 ;
        RECT 67.175 180.960 68.385 181.710 ;
        RECT 67.175 180.250 67.695 180.790 ;
        RECT 67.865 180.420 68.385 180.960 ;
        RECT 68.555 181.210 68.855 181.540 ;
        RECT 69.025 181.230 69.300 181.710 ;
        RECT 68.555 180.300 68.725 181.210 ;
        RECT 69.480 181.060 69.775 181.450 ;
        RECT 69.945 181.230 70.200 181.710 ;
        RECT 70.375 181.060 70.635 181.450 ;
        RECT 70.805 181.230 71.085 181.710 ;
        RECT 68.895 180.470 69.245 181.040 ;
        RECT 69.480 180.890 71.130 181.060 ;
        RECT 71.315 180.940 73.905 181.710 ;
        RECT 74.080 181.165 79.425 181.710 ;
        RECT 69.415 180.550 70.555 180.720 ;
        RECT 69.415 180.300 69.585 180.550 ;
        RECT 70.725 180.380 71.130 180.890 ;
        RECT 67.175 179.160 68.385 180.250 ;
        RECT 68.555 180.130 69.585 180.300 ;
        RECT 70.375 180.210 71.130 180.380 ;
        RECT 71.315 180.250 72.525 180.770 ;
        RECT 72.695 180.420 73.905 180.940 ;
        RECT 68.555 179.330 68.865 180.130 ;
        RECT 70.375 179.960 70.635 180.210 ;
        RECT 69.035 179.160 69.345 179.960 ;
        RECT 69.515 179.790 70.635 179.960 ;
        RECT 69.515 179.330 69.775 179.790 ;
        RECT 69.945 179.160 70.200 179.620 ;
        RECT 70.375 179.330 70.635 179.790 ;
        RECT 70.805 179.160 71.090 180.030 ;
        RECT 71.315 179.160 73.905 180.250 ;
        RECT 75.670 179.595 76.020 180.845 ;
        RECT 77.500 180.335 77.840 181.165 ;
        RECT 79.595 180.985 79.885 181.710 ;
        RECT 80.515 180.940 82.185 181.710 ;
        RECT 82.415 181.230 82.695 181.710 ;
        RECT 82.865 181.060 83.125 181.450 ;
        RECT 83.300 181.230 83.555 181.710 ;
        RECT 83.725 181.060 84.020 181.450 ;
        RECT 84.200 181.230 84.475 181.710 ;
        RECT 84.645 181.210 84.945 181.540 ;
        RECT 74.080 179.160 79.425 179.595 ;
        RECT 79.595 179.160 79.885 180.325 ;
        RECT 80.515 180.250 81.265 180.770 ;
        RECT 81.435 180.420 82.185 180.940 ;
        RECT 82.370 180.890 84.020 181.060 ;
        RECT 82.370 180.380 82.775 180.890 ;
        RECT 82.945 180.550 84.085 180.720 ;
        RECT 80.515 179.160 82.185 180.250 ;
        RECT 82.370 180.210 83.125 180.380 ;
        RECT 82.410 179.160 82.695 180.030 ;
        RECT 82.865 179.960 83.125 180.210 ;
        RECT 83.915 180.300 84.085 180.550 ;
        RECT 84.255 180.470 84.605 181.040 ;
        RECT 84.775 180.300 84.945 181.210 ;
        RECT 83.915 180.130 84.945 180.300 ;
        RECT 82.865 179.790 83.985 179.960 ;
        RECT 82.865 179.330 83.125 179.790 ;
        RECT 83.300 179.160 83.555 179.620 ;
        RECT 83.725 179.330 83.985 179.790 ;
        RECT 84.155 179.160 84.465 179.960 ;
        RECT 84.635 179.330 84.945 180.130 ;
        RECT 86.040 181.000 86.295 181.530 ;
        RECT 86.465 181.250 86.770 181.710 ;
        RECT 87.015 181.330 88.085 181.500 ;
        RECT 86.040 180.350 86.250 181.000 ;
        RECT 87.015 180.975 87.335 181.330 ;
        RECT 87.010 180.800 87.335 180.975 ;
        RECT 86.420 180.500 87.335 180.800 ;
        RECT 87.505 180.760 87.745 181.160 ;
        RECT 87.915 181.100 88.085 181.330 ;
        RECT 88.255 181.270 88.445 181.710 ;
        RECT 88.615 181.260 89.565 181.540 ;
        RECT 89.785 181.350 90.135 181.520 ;
        RECT 87.915 180.930 88.445 181.100 ;
        RECT 86.420 180.470 87.160 180.500 ;
        RECT 86.040 179.470 86.295 180.350 ;
        RECT 86.465 179.160 86.770 180.300 ;
        RECT 86.990 179.880 87.160 180.470 ;
        RECT 87.505 180.390 88.045 180.760 ;
        RECT 88.225 180.650 88.445 180.930 ;
        RECT 88.615 180.480 88.785 181.260 ;
        RECT 88.380 180.310 88.785 180.480 ;
        RECT 88.955 180.470 89.305 181.090 ;
        RECT 88.380 180.220 88.550 180.310 ;
        RECT 89.475 180.300 89.685 181.090 ;
        RECT 87.330 180.050 88.550 180.220 ;
        RECT 89.010 180.140 89.685 180.300 ;
        RECT 86.990 179.710 87.790 179.880 ;
        RECT 87.110 179.160 87.440 179.540 ;
        RECT 87.620 179.420 87.790 179.710 ;
        RECT 88.380 179.670 88.550 180.050 ;
        RECT 88.720 180.130 89.685 180.140 ;
        RECT 89.875 180.960 90.135 181.350 ;
        RECT 90.345 181.250 90.675 181.710 ;
        RECT 91.550 181.320 92.405 181.490 ;
        RECT 92.610 181.320 93.105 181.490 ;
        RECT 93.275 181.350 93.605 181.710 ;
        RECT 89.875 180.270 90.045 180.960 ;
        RECT 90.215 180.610 90.385 180.790 ;
        RECT 90.555 180.780 91.345 181.030 ;
        RECT 91.550 180.610 91.720 181.320 ;
        RECT 91.890 180.810 92.245 181.030 ;
        RECT 90.215 180.440 91.905 180.610 ;
        RECT 88.720 179.840 89.180 180.130 ;
        RECT 89.875 180.100 91.375 180.270 ;
        RECT 89.875 179.960 90.045 180.100 ;
        RECT 89.485 179.790 90.045 179.960 ;
        RECT 87.960 179.160 88.210 179.620 ;
        RECT 88.380 179.330 89.250 179.670 ;
        RECT 89.485 179.330 89.655 179.790 ;
        RECT 90.490 179.760 91.565 179.930 ;
        RECT 89.825 179.160 90.195 179.620 ;
        RECT 90.490 179.420 90.660 179.760 ;
        RECT 90.830 179.160 91.160 179.590 ;
        RECT 91.395 179.420 91.565 179.760 ;
        RECT 91.735 179.660 91.905 180.440 ;
        RECT 92.075 180.220 92.245 180.810 ;
        RECT 92.415 180.410 92.765 181.030 ;
        RECT 92.075 179.830 92.540 180.220 ;
        RECT 92.935 179.960 93.105 181.320 ;
        RECT 93.275 180.130 93.735 181.180 ;
        RECT 92.710 179.790 93.105 179.960 ;
        RECT 92.710 179.660 92.880 179.790 ;
        RECT 91.735 179.330 92.415 179.660 ;
        RECT 92.630 179.330 92.880 179.660 ;
        RECT 93.050 179.160 93.300 179.620 ;
        RECT 93.470 179.345 93.795 180.130 ;
        RECT 93.965 179.330 94.135 181.450 ;
        RECT 94.305 181.330 94.635 181.710 ;
        RECT 94.805 181.160 95.060 181.450 ;
        RECT 95.325 181.230 95.625 181.710 ;
        RECT 94.310 180.990 95.060 181.160 ;
        RECT 95.795 181.060 96.055 181.515 ;
        RECT 96.225 181.230 96.485 181.710 ;
        RECT 96.665 181.060 96.925 181.515 ;
        RECT 97.095 181.230 97.345 181.710 ;
        RECT 97.525 181.060 97.785 181.515 ;
        RECT 97.955 181.230 98.205 181.710 ;
        RECT 98.385 181.060 98.645 181.515 ;
        RECT 98.815 181.230 99.060 181.710 ;
        RECT 99.230 181.060 99.505 181.515 ;
        RECT 99.675 181.230 99.920 181.710 ;
        RECT 100.090 181.060 100.350 181.515 ;
        RECT 100.520 181.230 100.780 181.710 ;
        RECT 100.950 181.060 101.210 181.515 ;
        RECT 101.380 181.230 101.640 181.710 ;
        RECT 101.810 181.060 102.070 181.515 ;
        RECT 102.240 181.150 102.500 181.710 ;
        RECT 94.310 180.000 94.540 180.990 ;
        RECT 95.325 180.890 102.070 181.060 ;
        RECT 94.710 180.170 95.060 180.820 ;
        RECT 95.325 180.300 96.490 180.890 ;
        RECT 102.670 180.720 102.920 181.530 ;
        RECT 103.100 181.185 103.360 181.710 ;
        RECT 103.530 180.720 103.780 181.530 ;
        RECT 103.960 181.200 104.265 181.710 ;
        RECT 96.660 180.470 103.780 180.720 ;
        RECT 103.950 180.470 104.265 181.030 ;
        RECT 105.355 180.985 105.645 181.710 ;
        RECT 106.020 180.930 106.520 181.540 ;
        RECT 105.815 180.470 106.165 180.720 ;
        RECT 95.325 180.075 102.070 180.300 ;
        RECT 94.310 179.830 95.060 180.000 ;
        RECT 94.305 179.160 94.635 179.660 ;
        RECT 94.805 179.330 95.060 179.830 ;
        RECT 95.325 179.160 95.595 179.905 ;
        RECT 95.765 179.335 96.055 180.075 ;
        RECT 96.665 180.060 102.070 180.075 ;
        RECT 96.225 179.165 96.480 179.890 ;
        RECT 96.665 179.335 96.925 180.060 ;
        RECT 97.095 179.165 97.340 179.890 ;
        RECT 97.525 179.335 97.785 180.060 ;
        RECT 97.955 179.165 98.200 179.890 ;
        RECT 98.385 179.335 98.645 180.060 ;
        RECT 98.815 179.165 99.060 179.890 ;
        RECT 99.230 179.335 99.490 180.060 ;
        RECT 99.660 179.165 99.920 179.890 ;
        RECT 100.090 179.335 100.350 180.060 ;
        RECT 100.520 179.165 100.780 179.890 ;
        RECT 100.950 179.335 101.210 180.060 ;
        RECT 101.380 179.165 101.640 179.890 ;
        RECT 101.810 179.335 102.070 180.060 ;
        RECT 102.240 179.165 102.500 179.960 ;
        RECT 102.670 179.335 102.920 180.470 ;
        RECT 96.225 179.160 102.500 179.165 ;
        RECT 103.100 179.160 103.360 179.970 ;
        RECT 103.535 179.330 103.780 180.470 ;
        RECT 103.960 179.160 104.255 179.970 ;
        RECT 105.355 179.160 105.645 180.325 ;
        RECT 106.350 180.300 106.520 180.930 ;
        RECT 107.150 181.060 107.480 181.540 ;
        RECT 107.650 181.250 107.875 181.710 ;
        RECT 108.045 181.060 108.375 181.540 ;
        RECT 107.150 180.890 108.375 181.060 ;
        RECT 108.565 180.910 108.815 181.710 ;
        RECT 108.985 180.910 109.325 181.540 ;
        RECT 106.690 180.520 107.020 180.720 ;
        RECT 107.190 180.520 107.520 180.720 ;
        RECT 107.690 180.520 108.110 180.720 ;
        RECT 108.285 180.550 108.980 180.720 ;
        RECT 108.285 180.300 108.455 180.550 ;
        RECT 109.150 180.300 109.325 180.910 ;
        RECT 106.020 180.130 108.455 180.300 ;
        RECT 106.020 179.330 106.350 180.130 ;
        RECT 106.520 179.160 106.850 179.960 ;
        RECT 107.150 179.330 107.480 180.130 ;
        RECT 108.125 179.160 108.375 179.960 ;
        RECT 108.645 179.160 108.815 180.300 ;
        RECT 108.985 179.330 109.325 180.300 ;
        RECT 109.495 181.035 109.755 181.540 ;
        RECT 109.935 181.330 110.265 181.710 ;
        RECT 110.445 181.160 110.615 181.540 ;
        RECT 109.495 180.235 109.665 181.035 ;
        RECT 109.950 180.990 110.615 181.160 ;
        RECT 109.950 180.735 110.120 180.990 ;
        RECT 110.915 180.890 111.145 181.710 ;
        RECT 111.315 180.910 111.645 181.540 ;
        RECT 109.835 180.405 110.120 180.735 ;
        RECT 110.355 180.440 110.685 180.810 ;
        RECT 110.895 180.470 111.225 180.720 ;
        RECT 109.950 180.260 110.120 180.405 ;
        RECT 111.395 180.310 111.645 180.910 ;
        RECT 111.815 180.890 112.025 181.710 ;
        RECT 112.805 181.160 112.975 181.540 ;
        RECT 113.155 181.330 113.485 181.710 ;
        RECT 112.805 180.990 113.470 181.160 ;
        RECT 113.665 181.035 113.925 181.540 ;
        RECT 112.735 180.440 113.065 180.810 ;
        RECT 113.300 180.735 113.470 180.990 ;
        RECT 109.495 179.330 109.765 180.235 ;
        RECT 109.950 180.090 110.615 180.260 ;
        RECT 109.935 179.160 110.265 179.920 ;
        RECT 110.445 179.330 110.615 180.090 ;
        RECT 110.915 179.160 111.145 180.300 ;
        RECT 111.315 179.330 111.645 180.310 ;
        RECT 113.300 180.405 113.585 180.735 ;
        RECT 111.815 179.160 112.025 180.300 ;
        RECT 113.300 180.260 113.470 180.405 ;
        RECT 112.805 180.090 113.470 180.260 ;
        RECT 113.755 180.235 113.925 181.035 ;
        RECT 114.555 180.940 117.145 181.710 ;
        RECT 117.315 180.960 118.525 181.710 ;
        RECT 112.805 179.330 112.975 180.090 ;
        RECT 113.155 179.160 113.485 179.920 ;
        RECT 113.655 179.330 113.925 180.235 ;
        RECT 114.555 180.250 115.765 180.770 ;
        RECT 115.935 180.420 117.145 180.940 ;
        RECT 117.315 180.250 117.835 180.790 ;
        RECT 118.005 180.420 118.525 180.960 ;
        RECT 114.555 179.160 117.145 180.250 ;
        RECT 117.315 179.160 118.525 180.250 ;
        RECT 11.430 178.990 118.610 179.160 ;
        RECT 11.515 177.900 12.725 178.990 ;
        RECT 11.515 177.190 12.035 177.730 ;
        RECT 12.205 177.360 12.725 177.900 ;
        RECT 13.355 177.900 15.025 178.990 ;
        RECT 13.355 177.380 14.105 177.900 ;
        RECT 15.195 177.825 15.485 178.990 ;
        RECT 16.575 177.900 20.085 178.990 ;
        RECT 14.275 177.210 15.025 177.730 ;
        RECT 16.575 177.380 18.265 177.900 ;
        RECT 20.295 177.850 20.525 178.990 ;
        RECT 20.695 177.840 21.025 178.820 ;
        RECT 21.195 177.850 21.405 178.990 ;
        RECT 21.750 178.360 22.035 178.820 ;
        RECT 22.205 178.530 22.475 178.990 ;
        RECT 21.750 178.140 22.705 178.360 ;
        RECT 18.435 177.210 20.085 177.730 ;
        RECT 20.275 177.430 20.605 177.680 ;
        RECT 11.515 176.440 12.725 177.190 ;
        RECT 13.355 176.440 15.025 177.210 ;
        RECT 15.195 176.440 15.485 177.165 ;
        RECT 16.575 176.440 20.085 177.210 ;
        RECT 20.295 176.440 20.525 177.260 ;
        RECT 20.775 177.240 21.025 177.840 ;
        RECT 21.635 177.410 22.325 177.970 ;
        RECT 20.695 176.610 21.025 177.240 ;
        RECT 21.195 176.440 21.405 177.260 ;
        RECT 22.495 177.240 22.705 178.140 ;
        RECT 21.750 177.070 22.705 177.240 ;
        RECT 22.875 177.970 23.275 178.820 ;
        RECT 23.465 178.360 23.745 178.820 ;
        RECT 24.265 178.530 24.590 178.990 ;
        RECT 23.465 178.140 24.590 178.360 ;
        RECT 22.875 177.410 23.970 177.970 ;
        RECT 24.140 177.680 24.590 178.140 ;
        RECT 24.760 177.850 25.145 178.820 ;
        RECT 21.750 176.610 22.035 177.070 ;
        RECT 22.205 176.440 22.475 176.900 ;
        RECT 22.875 176.610 23.275 177.410 ;
        RECT 24.140 177.350 24.695 177.680 ;
        RECT 24.140 177.240 24.590 177.350 ;
        RECT 23.465 177.070 24.590 177.240 ;
        RECT 24.865 177.180 25.145 177.850 ;
        RECT 25.315 178.230 25.830 178.640 ;
        RECT 26.065 178.230 26.235 178.990 ;
        RECT 26.405 178.650 28.435 178.820 ;
        RECT 25.315 177.420 25.655 178.230 ;
        RECT 26.405 177.985 26.575 178.650 ;
        RECT 26.970 178.310 28.095 178.480 ;
        RECT 25.825 177.795 26.575 177.985 ;
        RECT 26.745 177.970 27.755 178.140 ;
        RECT 25.315 177.250 26.545 177.420 ;
        RECT 23.465 176.610 23.745 177.070 ;
        RECT 24.265 176.440 24.590 176.900 ;
        RECT 24.760 176.610 25.145 177.180 ;
        RECT 25.590 176.645 25.835 177.250 ;
        RECT 26.055 176.440 26.565 176.975 ;
        RECT 26.745 176.610 26.935 177.970 ;
        RECT 27.105 177.630 27.380 177.770 ;
        RECT 27.105 177.460 27.385 177.630 ;
        RECT 27.105 176.610 27.380 177.460 ;
        RECT 27.585 177.170 27.755 177.970 ;
        RECT 27.925 177.180 28.095 178.310 ;
        RECT 28.265 177.680 28.435 178.650 ;
        RECT 28.605 177.850 28.775 178.990 ;
        RECT 28.945 177.850 29.280 178.820 ;
        RECT 28.265 177.350 28.460 177.680 ;
        RECT 28.685 177.350 28.940 177.680 ;
        RECT 28.685 177.180 28.855 177.350 ;
        RECT 29.110 177.180 29.280 177.850 ;
        RECT 29.455 177.900 30.665 178.990 ;
        RECT 30.835 177.900 34.345 178.990 ;
        RECT 29.455 177.360 29.975 177.900 ;
        RECT 30.145 177.190 30.665 177.730 ;
        RECT 30.835 177.380 32.525 177.900 ;
        RECT 34.515 177.850 34.855 178.820 ;
        RECT 35.025 177.850 35.195 178.990 ;
        RECT 35.465 178.190 35.715 178.990 ;
        RECT 36.360 178.020 36.690 178.820 ;
        RECT 36.990 178.190 37.320 178.990 ;
        RECT 37.490 178.020 37.820 178.820 ;
        RECT 35.385 177.850 37.820 178.020 ;
        RECT 38.195 177.900 40.785 178.990 ;
        RECT 32.695 177.210 34.345 177.730 ;
        RECT 27.925 177.010 28.855 177.180 ;
        RECT 27.925 176.975 28.100 177.010 ;
        RECT 27.570 176.610 28.100 176.975 ;
        RECT 28.525 176.440 28.855 176.840 ;
        RECT 29.025 176.610 29.280 177.180 ;
        RECT 29.455 176.440 30.665 177.190 ;
        RECT 30.835 176.440 34.345 177.210 ;
        RECT 34.515 177.240 34.690 177.850 ;
        RECT 35.385 177.600 35.555 177.850 ;
        RECT 34.860 177.430 35.555 177.600 ;
        RECT 35.730 177.430 36.150 177.630 ;
        RECT 36.320 177.430 36.650 177.630 ;
        RECT 36.820 177.430 37.150 177.630 ;
        RECT 34.515 176.610 34.855 177.240 ;
        RECT 35.025 176.440 35.275 177.240 ;
        RECT 35.465 177.090 36.690 177.260 ;
        RECT 35.465 176.610 35.795 177.090 ;
        RECT 35.965 176.440 36.190 176.900 ;
        RECT 36.360 176.610 36.690 177.090 ;
        RECT 37.320 177.220 37.490 177.850 ;
        RECT 37.675 177.430 38.025 177.680 ;
        RECT 38.195 177.380 39.405 177.900 ;
        RECT 40.955 177.825 41.245 178.990 ;
        RECT 41.415 177.900 44.925 178.990 ;
        RECT 37.320 176.610 37.820 177.220 ;
        RECT 39.575 177.210 40.785 177.730 ;
        RECT 41.415 177.380 43.105 177.900 ;
        RECT 45.095 177.850 45.435 178.820 ;
        RECT 45.605 177.850 45.775 178.990 ;
        RECT 46.045 178.190 46.295 178.990 ;
        RECT 46.940 178.020 47.270 178.820 ;
        RECT 47.570 178.190 47.900 178.990 ;
        RECT 48.070 178.020 48.400 178.820 ;
        RECT 45.965 177.850 48.400 178.020 ;
        RECT 49.235 177.900 50.905 178.990 ;
        RECT 51.130 178.120 51.415 178.990 ;
        RECT 51.585 178.360 51.845 178.820 ;
        RECT 52.020 178.530 52.275 178.990 ;
        RECT 52.445 178.360 52.705 178.820 ;
        RECT 51.585 178.190 52.705 178.360 ;
        RECT 52.875 178.190 53.185 178.990 ;
        RECT 51.585 177.940 51.845 178.190 ;
        RECT 53.355 178.020 53.665 178.820 ;
        RECT 43.275 177.210 44.925 177.730 ;
        RECT 38.195 176.440 40.785 177.210 ;
        RECT 40.955 176.440 41.245 177.165 ;
        RECT 41.415 176.440 44.925 177.210 ;
        RECT 45.095 177.240 45.270 177.850 ;
        RECT 45.965 177.600 46.135 177.850 ;
        RECT 45.440 177.430 46.135 177.600 ;
        RECT 46.310 177.430 46.730 177.630 ;
        RECT 46.900 177.430 47.230 177.630 ;
        RECT 47.400 177.430 47.730 177.630 ;
        RECT 45.095 176.610 45.435 177.240 ;
        RECT 45.605 176.440 45.855 177.240 ;
        RECT 46.045 177.090 47.270 177.260 ;
        RECT 46.045 176.610 46.375 177.090 ;
        RECT 46.545 176.440 46.770 176.900 ;
        RECT 46.940 176.610 47.270 177.090 ;
        RECT 47.900 177.220 48.070 177.850 ;
        RECT 48.255 177.430 48.605 177.680 ;
        RECT 49.235 177.380 49.985 177.900 ;
        RECT 51.090 177.770 51.845 177.940 ;
        RECT 52.635 177.850 53.665 178.020 ;
        RECT 47.900 176.610 48.400 177.220 ;
        RECT 50.155 177.210 50.905 177.730 ;
        RECT 49.235 176.440 50.905 177.210 ;
        RECT 51.090 177.260 51.495 177.770 ;
        RECT 52.635 177.600 52.805 177.850 ;
        RECT 51.665 177.430 52.805 177.600 ;
        RECT 51.090 177.090 52.740 177.260 ;
        RECT 52.975 177.110 53.325 177.680 ;
        RECT 51.135 176.440 51.415 176.920 ;
        RECT 51.585 176.700 51.845 177.090 ;
        RECT 52.020 176.440 52.275 176.920 ;
        RECT 52.445 176.700 52.740 177.090 ;
        RECT 53.495 176.940 53.665 177.850 ;
        RECT 53.835 177.900 55.045 178.990 ;
        RECT 53.835 177.360 54.355 177.900 ;
        RECT 55.220 177.840 55.480 178.990 ;
        RECT 55.655 177.915 55.910 178.820 ;
        RECT 56.080 178.230 56.410 178.990 ;
        RECT 56.625 178.060 56.795 178.820 ;
        RECT 54.525 177.190 55.045 177.730 ;
        RECT 52.920 176.440 53.195 176.920 ;
        RECT 53.365 176.610 53.665 176.940 ;
        RECT 53.835 176.440 55.045 177.190 ;
        RECT 55.220 176.440 55.480 177.280 ;
        RECT 55.655 177.185 55.825 177.915 ;
        RECT 56.080 177.890 56.795 178.060 ;
        RECT 56.080 177.680 56.250 177.890 ;
        RECT 57.060 177.840 57.320 178.990 ;
        RECT 57.495 177.915 57.750 178.820 ;
        RECT 57.920 178.230 58.250 178.990 ;
        RECT 58.465 178.060 58.635 178.820 ;
        RECT 55.995 177.350 56.250 177.680 ;
        RECT 55.655 176.610 55.910 177.185 ;
        RECT 56.080 177.160 56.250 177.350 ;
        RECT 56.530 177.340 56.885 177.710 ;
        RECT 56.080 176.990 56.795 177.160 ;
        RECT 56.080 176.440 56.410 176.820 ;
        RECT 56.625 176.610 56.795 176.990 ;
        RECT 57.060 176.440 57.320 177.280 ;
        RECT 57.495 177.185 57.665 177.915 ;
        RECT 57.920 177.890 58.635 178.060 ;
        RECT 58.985 178.060 59.155 178.820 ;
        RECT 59.370 178.230 59.700 178.990 ;
        RECT 58.985 177.890 59.700 178.060 ;
        RECT 59.870 177.915 60.125 178.820 ;
        RECT 57.920 177.680 58.090 177.890 ;
        RECT 57.835 177.350 58.090 177.680 ;
        RECT 57.495 176.610 57.750 177.185 ;
        RECT 57.920 177.160 58.090 177.350 ;
        RECT 58.370 177.340 58.725 177.710 ;
        RECT 58.895 177.340 59.250 177.710 ;
        RECT 59.530 177.680 59.700 177.890 ;
        RECT 59.530 177.350 59.785 177.680 ;
        RECT 59.530 177.160 59.700 177.350 ;
        RECT 59.955 177.185 60.125 177.915 ;
        RECT 60.300 177.840 60.560 178.990 ;
        RECT 61.665 177.930 61.995 178.990 ;
        RECT 62.175 177.680 62.345 178.605 ;
        RECT 62.515 178.400 62.845 178.800 ;
        RECT 63.015 178.630 63.345 178.990 ;
        RECT 63.545 178.400 64.245 178.820 ;
        RECT 62.515 178.170 64.245 178.400 ;
        RECT 62.515 177.950 62.845 178.170 ;
        RECT 63.040 177.680 63.365 177.970 ;
        RECT 61.655 177.350 61.965 177.680 ;
        RECT 62.175 177.350 62.550 177.680 ;
        RECT 62.870 177.350 63.365 177.680 ;
        RECT 63.540 177.430 63.870 177.970 ;
        RECT 64.040 177.290 64.245 178.170 ;
        RECT 64.965 178.060 65.135 178.820 ;
        RECT 65.315 178.230 65.645 178.990 ;
        RECT 64.965 177.890 65.630 178.060 ;
        RECT 65.815 177.915 66.085 178.820 ;
        RECT 65.460 177.745 65.630 177.890 ;
        RECT 64.895 177.340 65.225 177.710 ;
        RECT 65.460 177.415 65.745 177.745 ;
        RECT 57.920 176.990 58.635 177.160 ;
        RECT 57.920 176.440 58.250 176.820 ;
        RECT 58.465 176.610 58.635 176.990 ;
        RECT 58.985 176.990 59.700 177.160 ;
        RECT 58.985 176.610 59.155 176.990 ;
        RECT 59.370 176.440 59.700 176.820 ;
        RECT 59.870 176.610 60.125 177.185 ;
        RECT 60.300 176.440 60.560 177.280 ;
        RECT 64.015 177.200 64.245 177.290 ;
        RECT 61.665 176.970 63.025 177.180 ;
        RECT 61.665 176.610 61.995 176.970 ;
        RECT 62.165 176.440 62.495 176.800 ;
        RECT 62.695 176.610 63.025 176.970 ;
        RECT 63.535 176.610 64.245 177.200 ;
        RECT 65.460 177.160 65.630 177.415 ;
        RECT 64.965 176.990 65.630 177.160 ;
        RECT 65.915 177.115 66.085 177.915 ;
        RECT 66.715 177.825 67.005 178.990 ;
        RECT 67.175 177.915 67.445 178.820 ;
        RECT 67.615 178.230 67.945 178.990 ;
        RECT 68.125 178.060 68.295 178.820 ;
        RECT 64.965 176.610 65.135 176.990 ;
        RECT 65.315 176.440 65.645 176.820 ;
        RECT 65.825 176.610 66.085 177.115 ;
        RECT 66.715 176.440 67.005 177.165 ;
        RECT 67.175 177.115 67.345 177.915 ;
        RECT 67.630 177.890 68.295 178.060 ;
        RECT 68.555 177.900 71.145 178.990 ;
        RECT 71.315 178.020 71.625 178.820 ;
        RECT 71.795 178.190 72.105 178.990 ;
        RECT 72.275 178.360 72.535 178.820 ;
        RECT 72.705 178.530 72.960 178.990 ;
        RECT 73.135 178.360 73.395 178.820 ;
        RECT 72.275 178.190 73.395 178.360 ;
        RECT 67.630 177.745 67.800 177.890 ;
        RECT 67.515 177.415 67.800 177.745 ;
        RECT 67.630 177.160 67.800 177.415 ;
        RECT 68.035 177.340 68.365 177.710 ;
        RECT 68.555 177.380 69.765 177.900 ;
        RECT 71.315 177.850 72.345 178.020 ;
        RECT 69.935 177.210 71.145 177.730 ;
        RECT 67.175 176.610 67.435 177.115 ;
        RECT 67.630 176.990 68.295 177.160 ;
        RECT 67.615 176.440 67.945 176.820 ;
        RECT 68.125 176.610 68.295 176.990 ;
        RECT 68.555 176.440 71.145 177.210 ;
        RECT 71.315 176.940 71.485 177.850 ;
        RECT 71.655 177.110 72.005 177.680 ;
        RECT 72.175 177.600 72.345 177.850 ;
        RECT 73.135 177.940 73.395 178.190 ;
        RECT 73.565 178.120 73.850 178.990 ;
        RECT 73.135 177.770 73.890 177.940 ;
        RECT 72.175 177.430 73.315 177.600 ;
        RECT 73.485 177.260 73.890 177.770 ;
        RECT 74.075 177.900 75.745 178.990 ;
        RECT 76.290 178.010 76.545 178.680 ;
        RECT 76.725 178.190 77.010 178.990 ;
        RECT 77.190 178.270 77.520 178.780 ;
        RECT 74.075 177.380 74.825 177.900 ;
        RECT 72.240 177.090 73.890 177.260 ;
        RECT 74.995 177.210 75.745 177.730 ;
        RECT 71.315 176.610 71.615 176.940 ;
        RECT 71.785 176.440 72.060 176.920 ;
        RECT 72.240 176.700 72.535 177.090 ;
        RECT 72.705 176.440 72.960 176.920 ;
        RECT 73.135 176.700 73.395 177.090 ;
        RECT 73.565 176.440 73.845 176.920 ;
        RECT 74.075 176.440 75.745 177.210 ;
        RECT 76.290 177.150 76.470 178.010 ;
        RECT 77.190 177.680 77.440 178.270 ;
        RECT 77.790 178.120 77.960 178.730 ;
        RECT 78.130 178.300 78.460 178.990 ;
        RECT 78.690 178.440 78.930 178.730 ;
        RECT 79.130 178.610 79.550 178.990 ;
        RECT 79.730 178.520 80.360 178.770 ;
        RECT 80.830 178.610 81.160 178.990 ;
        RECT 79.730 178.440 79.900 178.520 ;
        RECT 81.330 178.440 81.500 178.730 ;
        RECT 81.680 178.610 82.060 178.990 ;
        RECT 82.300 178.605 83.130 178.775 ;
        RECT 78.690 178.270 79.900 178.440 ;
        RECT 76.640 177.350 77.440 177.680 ;
        RECT 76.290 176.950 76.545 177.150 ;
        RECT 76.205 176.780 76.545 176.950 ;
        RECT 76.290 176.620 76.545 176.780 ;
        RECT 76.725 176.440 77.010 176.900 ;
        RECT 77.190 176.700 77.440 177.350 ;
        RECT 77.640 178.100 77.960 178.120 ;
        RECT 77.640 177.930 79.560 178.100 ;
        RECT 77.640 177.035 77.830 177.930 ;
        RECT 79.730 177.760 79.900 178.270 ;
        RECT 80.070 178.010 80.590 178.320 ;
        RECT 78.000 177.590 79.900 177.760 ;
        RECT 78.000 177.530 78.330 177.590 ;
        RECT 78.480 177.360 78.810 177.420 ;
        RECT 78.150 177.090 78.810 177.360 ;
        RECT 77.640 176.705 77.960 177.035 ;
        RECT 78.140 176.440 78.800 176.920 ;
        RECT 79.000 176.830 79.170 177.590 ;
        RECT 80.070 177.420 80.250 177.830 ;
        RECT 79.340 177.250 79.670 177.370 ;
        RECT 80.420 177.250 80.590 178.010 ;
        RECT 79.340 177.080 80.590 177.250 ;
        RECT 80.760 178.190 82.130 178.440 ;
        RECT 80.760 177.420 80.950 178.190 ;
        RECT 81.880 177.930 82.130 178.190 ;
        RECT 81.120 177.760 81.370 177.920 ;
        RECT 82.300 177.760 82.470 178.605 ;
        RECT 83.365 178.320 83.535 178.820 ;
        RECT 83.705 178.490 84.035 178.990 ;
        RECT 82.640 177.930 83.140 178.310 ;
        RECT 83.365 178.150 84.060 178.320 ;
        RECT 81.120 177.590 82.470 177.760 ;
        RECT 82.050 177.550 82.470 177.590 ;
        RECT 80.760 177.080 81.180 177.420 ;
        RECT 81.470 177.090 81.880 177.420 ;
        RECT 79.000 176.660 79.850 176.830 ;
        RECT 80.410 176.440 80.730 176.900 ;
        RECT 80.930 176.650 81.180 177.080 ;
        RECT 81.470 176.440 81.880 176.880 ;
        RECT 82.050 176.820 82.220 177.550 ;
        RECT 82.390 177.000 82.740 177.370 ;
        RECT 82.920 177.060 83.140 177.930 ;
        RECT 83.310 177.360 83.720 177.980 ;
        RECT 83.890 177.180 84.060 178.150 ;
        RECT 83.365 176.990 84.060 177.180 ;
        RECT 82.050 176.620 83.065 176.820 ;
        RECT 83.365 176.660 83.535 176.990 ;
        RECT 83.705 176.440 84.035 176.820 ;
        RECT 84.250 176.700 84.475 178.820 ;
        RECT 84.645 178.490 84.975 178.990 ;
        RECT 85.145 178.320 85.315 178.820 ;
        RECT 84.650 178.150 85.315 178.320 ;
        RECT 86.495 178.230 87.010 178.640 ;
        RECT 87.245 178.230 87.415 178.990 ;
        RECT 87.585 178.650 89.615 178.820 ;
        RECT 84.650 177.160 84.880 178.150 ;
        RECT 85.050 177.330 85.400 177.980 ;
        RECT 86.495 177.420 86.835 178.230 ;
        RECT 87.585 177.985 87.755 178.650 ;
        RECT 88.150 178.310 89.275 178.480 ;
        RECT 87.005 177.795 87.755 177.985 ;
        RECT 87.925 177.970 88.935 178.140 ;
        RECT 86.495 177.250 87.725 177.420 ;
        RECT 84.650 176.990 85.315 177.160 ;
        RECT 84.645 176.440 84.975 176.820 ;
        RECT 85.145 176.700 85.315 176.990 ;
        RECT 86.770 176.645 87.015 177.250 ;
        RECT 87.235 176.440 87.745 176.975 ;
        RECT 87.925 176.610 88.115 177.970 ;
        RECT 88.285 176.950 88.560 177.770 ;
        RECT 88.765 177.170 88.935 177.970 ;
        RECT 89.105 177.180 89.275 178.310 ;
        RECT 89.445 177.680 89.615 178.650 ;
        RECT 89.785 177.850 89.955 178.990 ;
        RECT 90.125 177.850 90.460 178.820 ;
        RECT 89.445 177.350 89.640 177.680 ;
        RECT 89.865 177.350 90.120 177.680 ;
        RECT 89.865 177.180 90.035 177.350 ;
        RECT 90.290 177.180 90.460 177.850 ;
        RECT 90.635 177.900 92.305 178.990 ;
        RECT 90.635 177.380 91.385 177.900 ;
        RECT 92.475 177.825 92.765 178.990 ;
        RECT 93.050 178.360 93.335 178.820 ;
        RECT 93.505 178.530 93.775 178.990 ;
        RECT 93.050 178.140 94.005 178.360 ;
        RECT 91.555 177.210 92.305 177.730 ;
        RECT 92.935 177.410 93.625 177.970 ;
        RECT 93.795 177.240 94.005 178.140 ;
        RECT 89.105 177.010 90.035 177.180 ;
        RECT 89.105 176.975 89.280 177.010 ;
        RECT 88.285 176.780 88.565 176.950 ;
        RECT 88.285 176.610 88.560 176.780 ;
        RECT 88.750 176.610 89.280 176.975 ;
        RECT 89.705 176.440 90.035 176.840 ;
        RECT 90.205 176.610 90.460 177.180 ;
        RECT 90.635 176.440 92.305 177.210 ;
        RECT 92.475 176.440 92.765 177.165 ;
        RECT 93.050 177.070 94.005 177.240 ;
        RECT 94.175 177.970 94.575 178.820 ;
        RECT 94.765 178.360 95.045 178.820 ;
        RECT 95.565 178.530 95.890 178.990 ;
        RECT 94.765 178.140 95.890 178.360 ;
        RECT 94.175 177.410 95.270 177.970 ;
        RECT 95.440 177.680 95.890 178.140 ;
        RECT 96.060 177.850 96.445 178.820 ;
        RECT 93.050 176.610 93.335 177.070 ;
        RECT 93.505 176.440 93.775 176.900 ;
        RECT 94.175 176.610 94.575 177.410 ;
        RECT 95.440 177.350 95.995 177.680 ;
        RECT 95.440 177.240 95.890 177.350 ;
        RECT 94.765 177.070 95.890 177.240 ;
        RECT 96.165 177.180 96.445 177.850 ;
        RECT 97.535 178.230 98.050 178.640 ;
        RECT 98.285 178.230 98.455 178.990 ;
        RECT 98.625 178.650 100.655 178.820 ;
        RECT 97.535 177.420 97.875 178.230 ;
        RECT 98.625 177.985 98.795 178.650 ;
        RECT 99.190 178.310 100.315 178.480 ;
        RECT 98.045 177.795 98.795 177.985 ;
        RECT 98.965 177.970 99.975 178.140 ;
        RECT 97.535 177.250 98.765 177.420 ;
        RECT 94.765 176.610 95.045 177.070 ;
        RECT 95.565 176.440 95.890 176.900 ;
        RECT 96.060 176.610 96.445 177.180 ;
        RECT 97.810 176.645 98.055 177.250 ;
        RECT 98.275 176.440 98.785 176.975 ;
        RECT 98.965 176.610 99.155 177.970 ;
        RECT 99.325 177.630 99.600 177.770 ;
        RECT 99.325 177.460 99.605 177.630 ;
        RECT 99.325 176.610 99.600 177.460 ;
        RECT 99.805 177.170 99.975 177.970 ;
        RECT 100.145 177.180 100.315 178.310 ;
        RECT 100.485 177.680 100.655 178.650 ;
        RECT 100.825 177.850 100.995 178.990 ;
        RECT 101.165 177.850 101.500 178.820 ;
        RECT 100.485 177.350 100.680 177.680 ;
        RECT 100.905 177.350 101.160 177.680 ;
        RECT 100.905 177.180 101.075 177.350 ;
        RECT 101.330 177.180 101.500 177.850 ;
        RECT 100.145 177.010 101.075 177.180 ;
        RECT 100.145 176.975 100.320 177.010 ;
        RECT 99.790 176.610 100.320 176.975 ;
        RECT 100.745 176.440 101.075 176.840 ;
        RECT 101.245 176.610 101.500 177.180 ;
        RECT 101.675 177.850 102.015 178.820 ;
        RECT 102.185 177.850 102.355 178.990 ;
        RECT 102.625 178.190 102.875 178.990 ;
        RECT 103.520 178.020 103.850 178.820 ;
        RECT 104.150 178.190 104.480 178.990 ;
        RECT 104.650 178.020 104.980 178.820 ;
        RECT 105.415 178.155 105.670 178.990 ;
        RECT 102.545 177.850 104.980 178.020 ;
        RECT 105.840 177.985 106.100 178.790 ;
        RECT 106.270 178.155 106.530 178.990 ;
        RECT 106.700 177.985 106.955 178.790 ;
        RECT 101.675 177.240 101.850 177.850 ;
        RECT 102.545 177.600 102.715 177.850 ;
        RECT 102.020 177.430 102.715 177.600 ;
        RECT 102.890 177.430 103.310 177.630 ;
        RECT 103.480 177.430 103.810 177.630 ;
        RECT 103.980 177.430 104.310 177.630 ;
        RECT 101.675 176.610 102.015 177.240 ;
        RECT 102.185 176.440 102.435 177.240 ;
        RECT 102.625 177.090 103.850 177.260 ;
        RECT 102.625 176.610 102.955 177.090 ;
        RECT 103.125 176.440 103.350 176.900 ;
        RECT 103.520 176.610 103.850 177.090 ;
        RECT 104.480 177.220 104.650 177.850 ;
        RECT 105.355 177.815 106.955 177.985 ;
        RECT 104.835 177.430 105.185 177.680 ;
        RECT 105.355 177.250 105.635 177.815 ;
        RECT 107.660 177.800 107.915 178.680 ;
        RECT 108.085 177.850 108.390 178.990 ;
        RECT 108.730 178.610 109.060 178.990 ;
        RECT 109.240 178.440 109.410 178.730 ;
        RECT 109.580 178.530 109.830 178.990 ;
        RECT 108.610 178.270 109.410 178.440 ;
        RECT 110.000 178.480 110.870 178.820 ;
        RECT 105.805 177.420 107.025 177.645 ;
        RECT 104.480 176.610 104.980 177.220 ;
        RECT 105.355 177.080 106.085 177.250 ;
        RECT 105.360 176.440 105.690 176.910 ;
        RECT 105.860 176.635 106.085 177.080 ;
        RECT 107.660 177.150 107.870 177.800 ;
        RECT 108.610 177.680 108.780 178.270 ;
        RECT 110.000 178.100 110.170 178.480 ;
        RECT 111.105 178.360 111.275 178.820 ;
        RECT 111.445 178.530 111.815 178.990 ;
        RECT 112.110 178.390 112.280 178.730 ;
        RECT 112.450 178.560 112.780 178.990 ;
        RECT 113.015 178.390 113.185 178.730 ;
        RECT 108.950 177.930 110.170 178.100 ;
        RECT 110.340 178.020 110.800 178.310 ;
        RECT 111.105 178.190 111.665 178.360 ;
        RECT 112.110 178.220 113.185 178.390 ;
        RECT 113.355 178.490 114.035 178.820 ;
        RECT 114.250 178.490 114.500 178.820 ;
        RECT 114.670 178.530 114.920 178.990 ;
        RECT 111.495 178.050 111.665 178.190 ;
        RECT 110.340 178.010 111.305 178.020 ;
        RECT 110.000 177.840 110.170 177.930 ;
        RECT 110.630 177.850 111.305 178.010 ;
        RECT 108.040 177.650 108.780 177.680 ;
        RECT 108.040 177.350 108.955 177.650 ;
        RECT 108.630 177.175 108.955 177.350 ;
        RECT 106.255 176.440 106.550 176.965 ;
        RECT 107.660 176.620 107.915 177.150 ;
        RECT 108.085 176.440 108.390 176.900 ;
        RECT 108.635 176.820 108.955 177.175 ;
        RECT 109.125 177.390 109.665 177.760 ;
        RECT 110.000 177.670 110.405 177.840 ;
        RECT 109.125 176.990 109.365 177.390 ;
        RECT 109.845 177.220 110.065 177.500 ;
        RECT 109.535 177.050 110.065 177.220 ;
        RECT 109.535 176.820 109.705 177.050 ;
        RECT 110.235 176.890 110.405 177.670 ;
        RECT 110.575 177.060 110.925 177.680 ;
        RECT 111.095 177.060 111.305 177.850 ;
        RECT 111.495 177.880 112.995 178.050 ;
        RECT 111.495 177.190 111.665 177.880 ;
        RECT 113.355 177.710 113.525 178.490 ;
        RECT 114.330 178.360 114.500 178.490 ;
        RECT 111.835 177.540 113.525 177.710 ;
        RECT 113.695 177.930 114.160 178.320 ;
        RECT 114.330 178.190 114.725 178.360 ;
        RECT 111.835 177.360 112.005 177.540 ;
        RECT 108.635 176.650 109.705 176.820 ;
        RECT 109.875 176.440 110.065 176.880 ;
        RECT 110.235 176.610 111.185 176.890 ;
        RECT 111.495 176.800 111.755 177.190 ;
        RECT 112.175 177.120 112.965 177.370 ;
        RECT 111.405 176.630 111.755 176.800 ;
        RECT 111.965 176.440 112.295 176.900 ;
        RECT 113.170 176.830 113.340 177.540 ;
        RECT 113.695 177.340 113.865 177.930 ;
        RECT 113.510 177.120 113.865 177.340 ;
        RECT 114.035 177.120 114.385 177.740 ;
        RECT 114.555 176.830 114.725 178.190 ;
        RECT 115.090 178.020 115.415 178.805 ;
        RECT 114.895 176.970 115.355 178.020 ;
        RECT 113.170 176.660 114.025 176.830 ;
        RECT 114.230 176.660 114.725 176.830 ;
        RECT 114.895 176.440 115.225 176.800 ;
        RECT 115.585 176.700 115.755 178.820 ;
        RECT 115.925 178.490 116.255 178.990 ;
        RECT 116.425 178.320 116.680 178.820 ;
        RECT 115.930 178.150 116.680 178.320 ;
        RECT 115.930 177.160 116.160 178.150 ;
        RECT 116.330 177.330 116.680 177.980 ;
        RECT 117.315 177.900 118.525 178.990 ;
        RECT 117.315 177.360 117.835 177.900 ;
        RECT 118.005 177.190 118.525 177.730 ;
        RECT 115.930 176.990 116.680 177.160 ;
        RECT 115.925 176.440 116.255 176.820 ;
        RECT 116.425 176.700 116.680 176.990 ;
        RECT 117.315 176.440 118.525 177.190 ;
        RECT 11.430 176.270 118.610 176.440 ;
        RECT 11.515 175.520 12.725 176.270 ;
        RECT 11.515 174.980 12.035 175.520 ;
        RECT 12.895 175.500 14.565 176.270 ;
        RECT 14.740 175.725 20.085 176.270 ;
        RECT 12.205 174.810 12.725 175.350 ;
        RECT 11.515 173.720 12.725 174.810 ;
        RECT 12.895 174.810 13.645 175.330 ;
        RECT 13.815 174.980 14.565 175.500 ;
        RECT 12.895 173.720 14.565 174.810 ;
        RECT 16.330 174.155 16.680 175.405 ;
        RECT 18.160 174.895 18.500 175.725 ;
        RECT 20.345 175.720 20.515 176.100 ;
        RECT 20.695 175.890 21.025 176.270 ;
        RECT 20.345 175.550 21.010 175.720 ;
        RECT 21.205 175.595 21.465 176.100 ;
        RECT 20.275 175.000 20.605 175.370 ;
        RECT 20.840 175.295 21.010 175.550 ;
        RECT 20.840 174.965 21.125 175.295 ;
        RECT 20.840 174.820 21.010 174.965 ;
        RECT 20.345 174.650 21.010 174.820 ;
        RECT 21.295 174.795 21.465 175.595 ;
        RECT 21.635 175.520 22.845 176.270 ;
        RECT 14.740 173.720 20.085 174.155 ;
        RECT 20.345 173.890 20.515 174.650 ;
        RECT 20.695 173.720 21.025 174.480 ;
        RECT 21.195 173.890 21.465 174.795 ;
        RECT 21.635 174.810 22.155 175.350 ;
        RECT 22.325 174.980 22.845 175.520 ;
        RECT 23.015 175.500 26.525 176.270 ;
        RECT 23.015 174.810 24.705 175.330 ;
        RECT 24.875 174.980 26.525 175.500 ;
        RECT 26.735 175.450 26.965 176.270 ;
        RECT 27.135 175.470 27.465 176.100 ;
        RECT 26.715 175.030 27.045 175.280 ;
        RECT 27.215 174.870 27.465 175.470 ;
        RECT 27.635 175.450 27.845 176.270 ;
        RECT 28.075 175.545 28.365 176.270 ;
        RECT 29.200 175.490 29.700 176.100 ;
        RECT 28.995 175.030 29.345 175.280 ;
        RECT 21.635 173.720 22.845 174.810 ;
        RECT 23.015 173.720 26.525 174.810 ;
        RECT 26.735 173.720 26.965 174.860 ;
        RECT 27.135 173.890 27.465 174.870 ;
        RECT 27.635 173.720 27.845 174.860 ;
        RECT 28.075 173.720 28.365 174.885 ;
        RECT 29.530 174.860 29.700 175.490 ;
        RECT 30.330 175.620 30.660 176.100 ;
        RECT 30.830 175.810 31.055 176.270 ;
        RECT 31.225 175.620 31.555 176.100 ;
        RECT 30.330 175.450 31.555 175.620 ;
        RECT 31.745 175.470 31.995 176.270 ;
        RECT 32.165 175.470 32.505 176.100 ;
        RECT 32.880 175.490 33.380 176.100 ;
        RECT 29.870 175.080 30.200 175.280 ;
        RECT 30.370 175.080 30.700 175.280 ;
        RECT 30.870 175.080 31.290 175.280 ;
        RECT 31.465 175.110 32.160 175.280 ;
        RECT 31.465 174.860 31.635 175.110 ;
        RECT 32.330 174.860 32.505 175.470 ;
        RECT 32.675 175.030 33.025 175.280 ;
        RECT 33.210 174.860 33.380 175.490 ;
        RECT 34.010 175.620 34.340 176.100 ;
        RECT 34.510 175.810 34.735 176.270 ;
        RECT 34.905 175.620 35.235 176.100 ;
        RECT 34.010 175.450 35.235 175.620 ;
        RECT 35.425 175.470 35.675 176.270 ;
        RECT 35.845 175.470 36.185 176.100 ;
        RECT 33.550 175.080 33.880 175.280 ;
        RECT 34.050 175.080 34.380 175.280 ;
        RECT 34.550 175.080 34.970 175.280 ;
        RECT 35.145 175.110 35.840 175.280 ;
        RECT 35.145 174.860 35.315 175.110 ;
        RECT 36.010 174.860 36.185 175.470 ;
        RECT 29.200 174.690 31.635 174.860 ;
        RECT 29.200 173.890 29.530 174.690 ;
        RECT 29.700 173.720 30.030 174.520 ;
        RECT 30.330 173.890 30.660 174.690 ;
        RECT 31.305 173.720 31.555 174.520 ;
        RECT 31.825 173.720 31.995 174.860 ;
        RECT 32.165 173.890 32.505 174.860 ;
        RECT 32.880 174.690 35.315 174.860 ;
        RECT 32.880 173.890 33.210 174.690 ;
        RECT 33.380 173.720 33.710 174.520 ;
        RECT 34.010 173.890 34.340 174.690 ;
        RECT 34.985 173.720 35.235 174.520 ;
        RECT 35.505 173.720 35.675 174.860 ;
        RECT 35.845 173.890 36.185 174.860 ;
        RECT 36.355 175.470 36.695 176.100 ;
        RECT 36.865 175.470 37.115 176.270 ;
        RECT 37.305 175.620 37.635 176.100 ;
        RECT 37.805 175.810 38.030 176.270 ;
        RECT 38.200 175.620 38.530 176.100 ;
        RECT 36.355 174.910 36.530 175.470 ;
        RECT 37.305 175.450 38.530 175.620 ;
        RECT 39.160 175.490 39.660 176.100 ;
        RECT 40.495 175.500 42.165 176.270 ;
        RECT 36.700 175.110 37.395 175.280 ;
        RECT 36.355 174.860 36.585 174.910 ;
        RECT 37.225 174.860 37.395 175.110 ;
        RECT 37.570 175.080 37.990 175.280 ;
        RECT 38.160 175.080 38.490 175.280 ;
        RECT 38.660 175.080 38.990 175.280 ;
        RECT 39.160 174.860 39.330 175.490 ;
        RECT 39.515 175.030 39.865 175.280 ;
        RECT 36.355 173.890 36.695 174.860 ;
        RECT 36.865 173.720 37.035 174.860 ;
        RECT 37.225 174.690 39.660 174.860 ;
        RECT 37.305 173.720 37.555 174.520 ;
        RECT 38.200 173.890 38.530 174.690 ;
        RECT 38.830 173.720 39.160 174.520 ;
        RECT 39.330 173.890 39.660 174.690 ;
        RECT 40.495 174.810 41.245 175.330 ;
        RECT 41.415 174.980 42.165 175.500 ;
        RECT 42.540 175.490 43.040 176.100 ;
        RECT 42.335 175.030 42.685 175.280 ;
        RECT 42.870 174.860 43.040 175.490 ;
        RECT 43.670 175.620 44.000 176.100 ;
        RECT 44.170 175.810 44.395 176.270 ;
        RECT 44.565 175.620 44.895 176.100 ;
        RECT 43.670 175.450 44.895 175.620 ;
        RECT 45.085 175.470 45.335 176.270 ;
        RECT 45.505 175.470 45.845 176.100 ;
        RECT 43.210 175.080 43.540 175.280 ;
        RECT 43.710 175.080 44.040 175.280 ;
        RECT 44.210 175.080 44.630 175.280 ;
        RECT 44.805 175.110 45.500 175.280 ;
        RECT 44.805 174.860 44.975 175.110 ;
        RECT 45.670 174.910 45.845 175.470 ;
        RECT 45.615 174.860 45.845 174.910 ;
        RECT 40.495 173.720 42.165 174.810 ;
        RECT 42.540 174.690 44.975 174.860 ;
        RECT 42.540 173.890 42.870 174.690 ;
        RECT 43.040 173.720 43.370 174.520 ;
        RECT 43.670 173.890 44.000 174.690 ;
        RECT 44.645 173.720 44.895 174.520 ;
        RECT 45.165 173.720 45.335 174.860 ;
        RECT 45.505 173.890 45.845 174.860 ;
        RECT 46.015 175.470 46.355 176.100 ;
        RECT 46.525 175.470 46.775 176.270 ;
        RECT 46.965 175.620 47.295 176.100 ;
        RECT 47.465 175.810 47.690 176.270 ;
        RECT 47.860 175.620 48.190 176.100 ;
        RECT 46.015 174.860 46.190 175.470 ;
        RECT 46.965 175.450 48.190 175.620 ;
        RECT 48.820 175.490 49.320 176.100 ;
        RECT 50.155 175.500 53.665 176.270 ;
        RECT 53.835 175.545 54.125 176.270 ;
        RECT 54.755 175.500 58.265 176.270 ;
        RECT 58.525 175.720 58.695 176.100 ;
        RECT 58.875 175.890 59.205 176.270 ;
        RECT 58.525 175.550 59.190 175.720 ;
        RECT 59.385 175.595 59.645 176.100 ;
        RECT 46.360 175.110 47.055 175.280 ;
        RECT 46.885 174.860 47.055 175.110 ;
        RECT 47.230 175.080 47.650 175.280 ;
        RECT 47.820 175.080 48.150 175.280 ;
        RECT 48.320 175.080 48.650 175.280 ;
        RECT 48.820 174.860 48.990 175.490 ;
        RECT 49.175 175.030 49.525 175.280 ;
        RECT 46.015 173.890 46.355 174.860 ;
        RECT 46.525 173.720 46.695 174.860 ;
        RECT 46.885 174.690 49.320 174.860 ;
        RECT 46.965 173.720 47.215 174.520 ;
        RECT 47.860 173.890 48.190 174.690 ;
        RECT 48.490 173.720 48.820 174.520 ;
        RECT 48.990 173.890 49.320 174.690 ;
        RECT 50.155 174.810 51.845 175.330 ;
        RECT 52.015 174.980 53.665 175.500 ;
        RECT 50.155 173.720 53.665 174.810 ;
        RECT 53.835 173.720 54.125 174.885 ;
        RECT 54.755 174.810 56.445 175.330 ;
        RECT 56.615 174.980 58.265 175.500 ;
        RECT 58.455 175.000 58.785 175.370 ;
        RECT 59.020 175.295 59.190 175.550 ;
        RECT 59.020 174.965 59.305 175.295 ;
        RECT 59.020 174.820 59.190 174.965 ;
        RECT 54.755 173.720 58.265 174.810 ;
        RECT 58.525 174.650 59.190 174.820 ;
        RECT 59.475 174.795 59.645 175.595 ;
        RECT 59.905 175.720 60.075 176.100 ;
        RECT 60.255 175.890 60.585 176.270 ;
        RECT 59.905 175.550 60.570 175.720 ;
        RECT 60.765 175.595 61.025 176.100 ;
        RECT 59.835 175.000 60.165 175.370 ;
        RECT 60.400 175.295 60.570 175.550 ;
        RECT 60.400 174.965 60.685 175.295 ;
        RECT 60.400 174.820 60.570 174.965 ;
        RECT 58.525 173.890 58.695 174.650 ;
        RECT 58.875 173.720 59.205 174.480 ;
        RECT 59.375 173.890 59.645 174.795 ;
        RECT 59.905 174.650 60.570 174.820 ;
        RECT 60.855 174.795 61.025 175.595 ;
        RECT 59.905 173.890 60.075 174.650 ;
        RECT 60.255 173.720 60.585 174.480 ;
        RECT 60.755 173.890 61.025 174.795 ;
        RECT 61.195 175.595 61.455 176.100 ;
        RECT 61.635 175.890 61.965 176.270 ;
        RECT 62.145 175.720 62.315 176.100 ;
        RECT 61.195 174.795 61.365 175.595 ;
        RECT 61.650 175.550 62.315 175.720 ;
        RECT 61.650 175.295 61.820 175.550 ;
        RECT 62.580 175.430 62.840 176.270 ;
        RECT 63.015 175.525 63.270 176.100 ;
        RECT 63.440 175.890 63.770 176.270 ;
        RECT 63.985 175.720 64.155 176.100 ;
        RECT 64.485 175.910 64.815 176.270 ;
        RECT 65.345 175.910 65.675 176.270 ;
        RECT 66.205 175.910 66.535 176.270 ;
        RECT 66.765 175.910 68.835 176.100 ;
        RECT 66.765 175.890 67.885 175.910 ;
        RECT 63.440 175.550 64.155 175.720 ;
        RECT 64.985 175.720 65.175 175.840 ;
        RECT 61.535 174.965 61.820 175.295 ;
        RECT 62.055 175.000 62.385 175.370 ;
        RECT 61.650 174.820 61.820 174.965 ;
        RECT 61.195 173.890 61.465 174.795 ;
        RECT 61.650 174.650 62.315 174.820 ;
        RECT 61.635 173.720 61.965 174.480 ;
        RECT 62.145 173.890 62.315 174.650 ;
        RECT 62.580 173.720 62.840 174.870 ;
        RECT 63.015 174.795 63.185 175.525 ;
        RECT 63.440 175.360 63.610 175.550 ;
        RECT 63.355 175.030 63.610 175.360 ;
        RECT 63.440 174.820 63.610 175.030 ;
        RECT 63.890 175.000 64.245 175.370 ;
        RECT 64.475 175.280 64.815 175.590 ;
        RECT 64.985 175.510 67.525 175.720 ;
        RECT 67.695 175.465 67.885 175.890 ;
        RECT 64.475 175.110 65.425 175.280 ;
        RECT 64.475 175.060 65.370 175.110 ;
        RECT 65.595 175.000 66.565 175.280 ;
        RECT 67.025 174.990 67.885 175.280 ;
        RECT 63.015 173.890 63.270 174.795 ;
        RECT 63.440 174.650 64.155 174.820 ;
        RECT 63.440 173.720 63.770 174.480 ;
        RECT 63.985 173.890 64.155 174.650 ;
        RECT 64.485 174.660 65.605 174.830 ;
        RECT 68.055 174.815 68.385 175.685 ;
        RECT 69.020 175.430 69.280 176.270 ;
        RECT 69.455 175.525 69.710 176.100 ;
        RECT 69.880 175.890 70.210 176.270 ;
        RECT 70.425 175.720 70.595 176.100 ;
        RECT 69.880 175.550 70.595 175.720 ;
        RECT 64.485 173.890 64.745 174.660 ;
        RECT 64.915 173.720 65.245 174.490 ;
        RECT 65.415 174.060 65.605 174.660 ;
        RECT 65.775 174.645 68.385 174.815 ;
        RECT 65.775 174.230 66.105 174.645 ;
        RECT 66.275 174.060 66.535 174.255 ;
        RECT 65.415 173.890 66.535 174.060 ;
        RECT 66.765 173.720 67.095 174.440 ;
        RECT 67.265 173.890 67.455 174.645 ;
        RECT 67.625 173.720 67.955 174.440 ;
        RECT 68.125 173.890 68.385 174.645 ;
        RECT 68.555 174.385 68.845 175.360 ;
        RECT 68.555 173.720 68.815 174.180 ;
        RECT 69.020 173.720 69.280 174.870 ;
        RECT 69.455 174.795 69.625 175.525 ;
        RECT 69.880 175.360 70.050 175.550 ;
        RECT 71.775 175.500 75.285 176.270 ;
        RECT 69.795 175.030 70.050 175.360 ;
        RECT 69.880 174.820 70.050 175.030 ;
        RECT 70.330 175.000 70.685 175.370 ;
        RECT 69.455 173.890 69.710 174.795 ;
        RECT 69.880 174.650 70.595 174.820 ;
        RECT 69.880 173.720 70.210 174.480 ;
        RECT 70.425 173.890 70.595 174.650 ;
        RECT 71.775 174.810 73.465 175.330 ;
        RECT 73.635 174.980 75.285 175.500 ;
        RECT 75.730 175.460 75.975 176.065 ;
        RECT 76.195 175.735 76.705 176.270 ;
        RECT 75.455 175.290 76.685 175.460 ;
        RECT 71.775 173.720 75.285 174.810 ;
        RECT 75.455 174.480 75.795 175.290 ;
        RECT 75.965 174.725 76.715 174.915 ;
        RECT 75.455 174.070 75.970 174.480 ;
        RECT 76.205 173.720 76.375 174.480 ;
        RECT 76.545 174.060 76.715 174.725 ;
        RECT 76.885 174.740 77.075 176.100 ;
        RECT 77.245 175.250 77.520 176.100 ;
        RECT 77.710 175.735 78.240 176.100 ;
        RECT 78.665 175.870 78.995 176.270 ;
        RECT 78.065 175.700 78.240 175.735 ;
        RECT 77.245 175.080 77.525 175.250 ;
        RECT 77.245 174.940 77.520 175.080 ;
        RECT 77.725 174.740 77.895 175.540 ;
        RECT 76.885 174.570 77.895 174.740 ;
        RECT 78.065 175.530 78.995 175.700 ;
        RECT 79.165 175.530 79.420 176.100 ;
        RECT 79.595 175.545 79.885 176.270 ;
        RECT 78.065 174.400 78.235 175.530 ;
        RECT 78.825 175.360 78.995 175.530 ;
        RECT 77.110 174.230 78.235 174.400 ;
        RECT 78.405 175.030 78.600 175.360 ;
        RECT 78.825 175.030 79.080 175.360 ;
        RECT 78.405 174.060 78.575 175.030 ;
        RECT 79.250 174.860 79.420 175.530 ;
        RECT 80.575 175.450 80.785 176.270 ;
        RECT 80.955 175.470 81.285 176.100 ;
        RECT 76.545 173.890 78.575 174.060 ;
        RECT 78.745 173.720 78.915 174.860 ;
        RECT 79.085 173.890 79.420 174.860 ;
        RECT 79.595 173.720 79.885 174.885 ;
        RECT 80.955 174.870 81.205 175.470 ;
        RECT 81.455 175.450 81.685 176.270 ;
        RECT 81.985 175.720 82.155 176.100 ;
        RECT 82.335 175.890 82.665 176.270 ;
        RECT 81.985 175.550 82.650 175.720 ;
        RECT 82.845 175.595 83.105 176.100 ;
        RECT 81.375 175.030 81.705 175.280 ;
        RECT 81.915 175.000 82.245 175.370 ;
        RECT 82.480 175.295 82.650 175.550 ;
        RECT 82.480 174.965 82.765 175.295 ;
        RECT 80.575 173.720 80.785 174.860 ;
        RECT 80.955 173.890 81.285 174.870 ;
        RECT 81.455 173.720 81.685 174.860 ;
        RECT 82.480 174.820 82.650 174.965 ;
        RECT 81.985 174.650 82.650 174.820 ;
        RECT 82.935 174.795 83.105 175.595 ;
        RECT 83.365 175.720 83.535 176.100 ;
        RECT 83.715 175.890 84.045 176.270 ;
        RECT 83.365 175.550 84.030 175.720 ;
        RECT 84.225 175.595 84.485 176.100 ;
        RECT 83.295 175.000 83.625 175.370 ;
        RECT 83.860 175.295 84.030 175.550 ;
        RECT 83.860 174.965 84.145 175.295 ;
        RECT 83.860 174.820 84.030 174.965 ;
        RECT 81.985 173.890 82.155 174.650 ;
        RECT 82.335 173.720 82.665 174.480 ;
        RECT 82.835 173.890 83.105 174.795 ;
        RECT 83.365 174.650 84.030 174.820 ;
        RECT 84.315 174.795 84.485 175.595 ;
        RECT 85.575 175.500 89.085 176.270 ;
        RECT 83.365 173.890 83.535 174.650 ;
        RECT 83.715 173.720 84.045 174.480 ;
        RECT 84.215 173.890 84.485 174.795 ;
        RECT 85.575 174.810 87.265 175.330 ;
        RECT 87.435 174.980 89.085 175.500 ;
        RECT 89.630 175.560 89.885 176.090 ;
        RECT 90.065 175.810 90.350 176.270 ;
        RECT 85.575 173.720 89.085 174.810 ;
        RECT 89.630 174.700 89.810 175.560 ;
        RECT 90.530 175.360 90.780 176.010 ;
        RECT 89.980 175.030 90.780 175.360 ;
        RECT 89.630 174.230 89.885 174.700 ;
        RECT 89.545 174.060 89.885 174.230 ;
        RECT 89.630 174.030 89.885 174.060 ;
        RECT 90.065 173.720 90.350 174.520 ;
        RECT 90.530 174.440 90.780 175.030 ;
        RECT 90.980 175.675 91.300 176.005 ;
        RECT 91.480 175.790 92.140 176.270 ;
        RECT 92.340 175.880 93.190 176.050 ;
        RECT 90.980 174.780 91.170 175.675 ;
        RECT 91.490 175.350 92.150 175.620 ;
        RECT 91.820 175.290 92.150 175.350 ;
        RECT 91.340 175.120 91.670 175.180 ;
        RECT 92.340 175.120 92.510 175.880 ;
        RECT 93.750 175.810 94.070 176.270 ;
        RECT 94.270 175.630 94.520 176.060 ;
        RECT 94.810 175.830 95.220 176.270 ;
        RECT 95.390 175.890 96.405 176.090 ;
        RECT 92.680 175.460 93.930 175.630 ;
        RECT 92.680 175.340 93.010 175.460 ;
        RECT 91.340 174.950 93.240 175.120 ;
        RECT 90.980 174.610 92.900 174.780 ;
        RECT 90.980 174.590 91.300 174.610 ;
        RECT 90.530 173.930 90.860 174.440 ;
        RECT 91.130 173.980 91.300 174.590 ;
        RECT 93.070 174.440 93.240 174.950 ;
        RECT 93.410 174.880 93.590 175.290 ;
        RECT 93.760 174.700 93.930 175.460 ;
        RECT 91.470 173.720 91.800 174.410 ;
        RECT 92.030 174.270 93.240 174.440 ;
        RECT 93.410 174.390 93.930 174.700 ;
        RECT 94.100 175.290 94.520 175.630 ;
        RECT 94.810 175.290 95.220 175.620 ;
        RECT 94.100 174.520 94.290 175.290 ;
        RECT 95.390 175.160 95.560 175.890 ;
        RECT 96.705 175.720 96.875 176.050 ;
        RECT 97.045 175.890 97.375 176.270 ;
        RECT 95.730 175.340 96.080 175.710 ;
        RECT 95.390 175.120 95.810 175.160 ;
        RECT 94.460 174.950 95.810 175.120 ;
        RECT 94.460 174.790 94.710 174.950 ;
        RECT 95.220 174.520 95.470 174.780 ;
        RECT 94.100 174.270 95.470 174.520 ;
        RECT 92.030 173.980 92.270 174.270 ;
        RECT 93.070 174.190 93.240 174.270 ;
        RECT 92.470 173.720 92.890 174.100 ;
        RECT 93.070 173.940 93.700 174.190 ;
        RECT 94.170 173.720 94.500 174.100 ;
        RECT 94.670 173.980 94.840 174.270 ;
        RECT 95.640 174.105 95.810 174.950 ;
        RECT 96.260 174.780 96.480 175.650 ;
        RECT 96.705 175.530 97.400 175.720 ;
        RECT 95.980 174.400 96.480 174.780 ;
        RECT 96.650 174.730 97.060 175.350 ;
        RECT 97.230 174.560 97.400 175.530 ;
        RECT 96.705 174.390 97.400 174.560 ;
        RECT 95.020 173.720 95.400 174.100 ;
        RECT 95.640 173.935 96.470 174.105 ;
        RECT 96.705 173.890 96.875 174.390 ;
        RECT 97.045 173.720 97.375 174.220 ;
        RECT 97.590 173.890 97.815 176.010 ;
        RECT 97.985 175.890 98.315 176.270 ;
        RECT 98.485 175.720 98.655 176.010 ;
        RECT 97.990 175.550 98.655 175.720 ;
        RECT 97.990 174.560 98.220 175.550 ;
        RECT 98.915 175.520 100.125 176.270 ;
        RECT 98.390 174.730 98.740 175.380 ;
        RECT 98.915 174.810 99.435 175.350 ;
        RECT 99.605 174.980 100.125 175.520 ;
        RECT 100.295 175.470 100.635 176.100 ;
        RECT 100.805 175.470 101.055 176.270 ;
        RECT 101.245 175.620 101.575 176.100 ;
        RECT 101.745 175.810 101.970 176.270 ;
        RECT 102.140 175.620 102.470 176.100 ;
        RECT 100.295 174.860 100.470 175.470 ;
        RECT 101.245 175.450 102.470 175.620 ;
        RECT 103.100 175.490 103.600 176.100 ;
        RECT 103.975 175.520 105.185 176.270 ;
        RECT 105.355 175.545 105.645 176.270 ;
        RECT 100.640 175.110 101.335 175.280 ;
        RECT 101.165 174.860 101.335 175.110 ;
        RECT 101.510 175.080 101.930 175.280 ;
        RECT 102.100 175.080 102.430 175.280 ;
        RECT 102.600 175.080 102.930 175.280 ;
        RECT 103.100 174.860 103.270 175.490 ;
        RECT 103.455 175.030 103.805 175.280 ;
        RECT 97.990 174.390 98.655 174.560 ;
        RECT 97.985 173.720 98.315 174.220 ;
        RECT 98.485 173.890 98.655 174.390 ;
        RECT 98.915 173.720 100.125 174.810 ;
        RECT 100.295 173.890 100.635 174.860 ;
        RECT 100.805 173.720 100.975 174.860 ;
        RECT 101.165 174.690 103.600 174.860 ;
        RECT 101.245 173.720 101.495 174.520 ;
        RECT 102.140 173.890 102.470 174.690 ;
        RECT 102.770 173.720 103.100 174.520 ;
        RECT 103.270 173.890 103.600 174.690 ;
        RECT 103.975 174.810 104.495 175.350 ;
        RECT 104.665 174.980 105.185 175.520 ;
        RECT 107.010 175.460 107.255 176.065 ;
        RECT 107.475 175.735 107.985 176.270 ;
        RECT 106.735 175.290 107.965 175.460 ;
        RECT 103.975 173.720 105.185 174.810 ;
        RECT 105.355 173.720 105.645 174.885 ;
        RECT 106.735 174.480 107.075 175.290 ;
        RECT 107.245 174.725 107.995 174.915 ;
        RECT 106.735 174.070 107.250 174.480 ;
        RECT 107.485 173.720 107.655 174.480 ;
        RECT 107.825 174.060 107.995 174.725 ;
        RECT 108.165 174.740 108.355 176.100 ;
        RECT 108.525 175.250 108.800 176.100 ;
        RECT 108.990 175.735 109.520 176.100 ;
        RECT 109.945 175.870 110.275 176.270 ;
        RECT 109.345 175.700 109.520 175.735 ;
        RECT 108.525 175.080 108.805 175.250 ;
        RECT 108.525 174.940 108.800 175.080 ;
        RECT 109.005 174.740 109.175 175.540 ;
        RECT 108.165 174.570 109.175 174.740 ;
        RECT 109.345 175.530 110.275 175.700 ;
        RECT 110.445 175.530 110.700 176.100 ;
        RECT 111.800 175.725 117.145 176.270 ;
        RECT 109.345 174.400 109.515 175.530 ;
        RECT 110.105 175.360 110.275 175.530 ;
        RECT 108.390 174.230 109.515 174.400 ;
        RECT 109.685 175.030 109.880 175.360 ;
        RECT 110.105 175.030 110.360 175.360 ;
        RECT 109.685 174.060 109.855 175.030 ;
        RECT 110.530 174.860 110.700 175.530 ;
        RECT 107.825 173.890 109.855 174.060 ;
        RECT 110.025 173.720 110.195 174.860 ;
        RECT 110.365 173.890 110.700 174.860 ;
        RECT 113.390 174.155 113.740 175.405 ;
        RECT 115.220 174.895 115.560 175.725 ;
        RECT 117.315 175.520 118.525 176.270 ;
        RECT 117.315 174.810 117.835 175.350 ;
        RECT 118.005 174.980 118.525 175.520 ;
        RECT 111.800 173.720 117.145 174.155 ;
        RECT 117.315 173.720 118.525 174.810 ;
        RECT 11.430 173.550 118.610 173.720 ;
        RECT 11.515 172.460 12.725 173.550 ;
        RECT 11.515 171.750 12.035 172.290 ;
        RECT 12.205 171.920 12.725 172.460 ;
        RECT 13.875 172.410 14.085 173.550 ;
        RECT 14.255 172.400 14.585 173.380 ;
        RECT 14.755 172.410 14.985 173.550 ;
        RECT 11.515 171.000 12.725 171.750 ;
        RECT 13.875 171.000 14.085 171.820 ;
        RECT 14.255 171.800 14.505 172.400 ;
        RECT 15.195 172.385 15.485 173.550 ;
        RECT 15.660 172.360 15.915 173.240 ;
        RECT 16.085 172.410 16.390 173.550 ;
        RECT 16.730 173.170 17.060 173.550 ;
        RECT 17.240 173.000 17.410 173.290 ;
        RECT 17.580 173.090 17.830 173.550 ;
        RECT 16.610 172.830 17.410 173.000 ;
        RECT 18.000 173.040 18.870 173.380 ;
        RECT 14.675 171.990 15.005 172.240 ;
        RECT 14.255 171.170 14.585 171.800 ;
        RECT 14.755 171.000 14.985 171.820 ;
        RECT 15.195 171.000 15.485 171.725 ;
        RECT 15.660 171.710 15.870 172.360 ;
        RECT 16.610 172.240 16.780 172.830 ;
        RECT 18.000 172.660 18.170 173.040 ;
        RECT 19.105 172.920 19.275 173.380 ;
        RECT 19.445 173.090 19.815 173.550 ;
        RECT 20.110 172.950 20.280 173.290 ;
        RECT 20.450 173.120 20.780 173.550 ;
        RECT 21.015 172.950 21.185 173.290 ;
        RECT 16.950 172.490 18.170 172.660 ;
        RECT 18.340 172.580 18.800 172.870 ;
        RECT 19.105 172.750 19.665 172.920 ;
        RECT 20.110 172.780 21.185 172.950 ;
        RECT 21.355 173.050 22.035 173.380 ;
        RECT 22.250 173.050 22.500 173.380 ;
        RECT 22.670 173.090 22.920 173.550 ;
        RECT 19.495 172.610 19.665 172.750 ;
        RECT 18.340 172.570 19.305 172.580 ;
        RECT 18.000 172.400 18.170 172.490 ;
        RECT 18.630 172.410 19.305 172.570 ;
        RECT 16.040 172.210 16.780 172.240 ;
        RECT 16.040 171.910 16.955 172.210 ;
        RECT 16.630 171.735 16.955 171.910 ;
        RECT 15.660 171.180 15.915 171.710 ;
        RECT 16.085 171.000 16.390 171.460 ;
        RECT 16.635 171.380 16.955 171.735 ;
        RECT 17.125 171.950 17.665 172.320 ;
        RECT 18.000 172.230 18.405 172.400 ;
        RECT 17.125 171.550 17.365 171.950 ;
        RECT 17.845 171.780 18.065 172.060 ;
        RECT 17.535 171.610 18.065 171.780 ;
        RECT 17.535 171.380 17.705 171.610 ;
        RECT 18.235 171.450 18.405 172.230 ;
        RECT 18.575 171.620 18.925 172.240 ;
        RECT 19.095 171.620 19.305 172.410 ;
        RECT 19.495 172.440 20.995 172.610 ;
        RECT 19.495 171.750 19.665 172.440 ;
        RECT 21.355 172.270 21.525 173.050 ;
        RECT 22.330 172.920 22.500 173.050 ;
        RECT 19.835 172.100 21.525 172.270 ;
        RECT 21.695 172.490 22.160 172.880 ;
        RECT 22.330 172.750 22.725 172.920 ;
        RECT 19.835 171.920 20.005 172.100 ;
        RECT 16.635 171.210 17.705 171.380 ;
        RECT 17.875 171.000 18.065 171.440 ;
        RECT 18.235 171.170 19.185 171.450 ;
        RECT 19.495 171.360 19.755 171.750 ;
        RECT 20.175 171.680 20.965 171.930 ;
        RECT 19.405 171.190 19.755 171.360 ;
        RECT 19.965 171.000 20.295 171.460 ;
        RECT 21.170 171.390 21.340 172.100 ;
        RECT 21.695 171.900 21.865 172.490 ;
        RECT 21.510 171.680 21.865 171.900 ;
        RECT 22.035 171.680 22.385 172.300 ;
        RECT 22.555 171.390 22.725 172.750 ;
        RECT 23.090 172.580 23.415 173.365 ;
        RECT 22.895 171.530 23.355 172.580 ;
        RECT 21.170 171.220 22.025 171.390 ;
        RECT 22.230 171.220 22.725 171.390 ;
        RECT 22.895 171.000 23.225 171.360 ;
        RECT 23.585 171.260 23.755 173.380 ;
        RECT 23.925 173.050 24.255 173.550 ;
        RECT 24.425 172.880 24.680 173.380 ;
        RECT 23.930 172.710 24.680 172.880 ;
        RECT 23.930 171.720 24.160 172.710 ;
        RECT 24.330 171.890 24.680 172.540 ;
        RECT 25.320 172.360 25.575 173.240 ;
        RECT 25.745 172.410 26.050 173.550 ;
        RECT 26.390 173.170 26.720 173.550 ;
        RECT 26.900 173.000 27.070 173.290 ;
        RECT 27.240 173.090 27.490 173.550 ;
        RECT 26.270 172.830 27.070 173.000 ;
        RECT 27.660 173.040 28.530 173.380 ;
        RECT 23.930 171.550 24.680 171.720 ;
        RECT 23.925 171.000 24.255 171.380 ;
        RECT 24.425 171.260 24.680 171.550 ;
        RECT 25.320 171.710 25.530 172.360 ;
        RECT 26.270 172.240 26.440 172.830 ;
        RECT 27.660 172.660 27.830 173.040 ;
        RECT 28.765 172.920 28.935 173.380 ;
        RECT 29.105 173.090 29.475 173.550 ;
        RECT 29.770 172.950 29.940 173.290 ;
        RECT 30.110 173.120 30.440 173.550 ;
        RECT 30.675 172.950 30.845 173.290 ;
        RECT 26.610 172.490 27.830 172.660 ;
        RECT 28.000 172.580 28.460 172.870 ;
        RECT 28.765 172.750 29.325 172.920 ;
        RECT 29.770 172.780 30.845 172.950 ;
        RECT 31.015 173.050 31.695 173.380 ;
        RECT 31.910 173.050 32.160 173.380 ;
        RECT 32.330 173.090 32.580 173.550 ;
        RECT 29.155 172.610 29.325 172.750 ;
        RECT 28.000 172.570 28.965 172.580 ;
        RECT 27.660 172.400 27.830 172.490 ;
        RECT 28.290 172.410 28.965 172.570 ;
        RECT 25.700 172.210 26.440 172.240 ;
        RECT 25.700 171.910 26.615 172.210 ;
        RECT 26.290 171.735 26.615 171.910 ;
        RECT 25.320 171.180 25.575 171.710 ;
        RECT 25.745 171.000 26.050 171.460 ;
        RECT 26.295 171.380 26.615 171.735 ;
        RECT 26.785 171.950 27.325 172.320 ;
        RECT 27.660 172.230 28.065 172.400 ;
        RECT 26.785 171.550 27.025 171.950 ;
        RECT 27.505 171.780 27.725 172.060 ;
        RECT 27.195 171.610 27.725 171.780 ;
        RECT 27.195 171.380 27.365 171.610 ;
        RECT 27.895 171.450 28.065 172.230 ;
        RECT 28.235 171.620 28.585 172.240 ;
        RECT 28.755 171.620 28.965 172.410 ;
        RECT 29.155 172.440 30.655 172.610 ;
        RECT 29.155 171.750 29.325 172.440 ;
        RECT 31.015 172.270 31.185 173.050 ;
        RECT 31.990 172.920 32.160 173.050 ;
        RECT 29.495 172.100 31.185 172.270 ;
        RECT 31.355 172.490 31.820 172.880 ;
        RECT 31.990 172.750 32.385 172.920 ;
        RECT 29.495 171.920 29.665 172.100 ;
        RECT 26.295 171.210 27.365 171.380 ;
        RECT 27.535 171.000 27.725 171.440 ;
        RECT 27.895 171.170 28.845 171.450 ;
        RECT 29.155 171.360 29.415 171.750 ;
        RECT 29.835 171.680 30.625 171.930 ;
        RECT 29.065 171.190 29.415 171.360 ;
        RECT 29.625 171.000 29.955 171.460 ;
        RECT 30.830 171.390 31.000 172.100 ;
        RECT 31.355 171.900 31.525 172.490 ;
        RECT 31.170 171.680 31.525 171.900 ;
        RECT 31.695 171.680 32.045 172.300 ;
        RECT 32.215 171.390 32.385 172.750 ;
        RECT 32.750 172.580 33.075 173.365 ;
        RECT 32.555 171.530 33.015 172.580 ;
        RECT 30.830 171.220 31.685 171.390 ;
        RECT 31.890 171.220 32.385 171.390 ;
        RECT 32.555 171.000 32.885 171.360 ;
        RECT 33.245 171.260 33.415 173.380 ;
        RECT 33.585 173.050 33.915 173.550 ;
        RECT 34.085 172.880 34.340 173.380 ;
        RECT 33.590 172.710 34.340 172.880 ;
        RECT 33.590 171.720 33.820 172.710 ;
        RECT 33.990 171.890 34.340 172.540 ;
        RECT 35.435 172.410 35.775 173.380 ;
        RECT 35.945 172.410 36.115 173.550 ;
        RECT 36.385 172.750 36.635 173.550 ;
        RECT 37.280 172.580 37.610 173.380 ;
        RECT 37.910 172.750 38.240 173.550 ;
        RECT 38.410 172.580 38.740 173.380 ;
        RECT 36.305 172.410 38.740 172.580 ;
        RECT 39.115 172.460 40.785 173.550 ;
        RECT 35.435 171.800 35.610 172.410 ;
        RECT 36.305 172.160 36.475 172.410 ;
        RECT 35.780 171.990 36.475 172.160 ;
        RECT 36.650 171.990 37.070 172.190 ;
        RECT 37.240 171.990 37.570 172.190 ;
        RECT 37.740 171.990 38.070 172.190 ;
        RECT 33.590 171.550 34.340 171.720 ;
        RECT 33.585 171.000 33.915 171.380 ;
        RECT 34.085 171.260 34.340 171.550 ;
        RECT 35.435 171.170 35.775 171.800 ;
        RECT 35.945 171.000 36.195 171.800 ;
        RECT 36.385 171.650 37.610 171.820 ;
        RECT 36.385 171.170 36.715 171.650 ;
        RECT 36.885 171.000 37.110 171.460 ;
        RECT 37.280 171.170 37.610 171.650 ;
        RECT 38.240 171.780 38.410 172.410 ;
        RECT 38.595 171.990 38.945 172.240 ;
        RECT 39.115 171.940 39.865 172.460 ;
        RECT 40.955 172.385 41.245 173.550 ;
        RECT 41.415 172.460 44.005 173.550 ;
        RECT 38.240 171.170 38.740 171.780 ;
        RECT 40.035 171.770 40.785 172.290 ;
        RECT 41.415 171.940 42.625 172.460 ;
        RECT 44.175 172.410 44.515 173.380 ;
        RECT 44.685 172.410 44.855 173.550 ;
        RECT 45.125 172.750 45.375 173.550 ;
        RECT 46.020 172.580 46.350 173.380 ;
        RECT 46.650 172.750 46.980 173.550 ;
        RECT 47.150 172.580 47.480 173.380 ;
        RECT 45.045 172.410 47.480 172.580 ;
        RECT 47.855 172.460 49.525 173.550 ;
        RECT 42.795 171.770 44.005 172.290 ;
        RECT 39.115 171.000 40.785 171.770 ;
        RECT 40.955 171.000 41.245 171.725 ;
        RECT 41.415 171.000 44.005 171.770 ;
        RECT 44.175 171.800 44.350 172.410 ;
        RECT 45.045 172.160 45.215 172.410 ;
        RECT 44.520 171.990 45.215 172.160 ;
        RECT 45.390 171.990 45.810 172.190 ;
        RECT 45.980 171.990 46.310 172.190 ;
        RECT 46.480 171.990 46.810 172.190 ;
        RECT 44.175 171.170 44.515 171.800 ;
        RECT 44.685 171.000 44.935 171.800 ;
        RECT 45.125 171.650 46.350 171.820 ;
        RECT 45.125 171.170 45.455 171.650 ;
        RECT 45.625 171.000 45.850 171.460 ;
        RECT 46.020 171.170 46.350 171.650 ;
        RECT 46.980 171.780 47.150 172.410 ;
        RECT 47.335 171.990 47.685 172.240 ;
        RECT 47.855 171.940 48.605 172.460 ;
        RECT 49.735 172.410 49.965 173.550 ;
        RECT 50.135 172.400 50.465 173.380 ;
        RECT 50.635 172.410 50.845 173.550 ;
        RECT 51.995 172.460 55.505 173.550 ;
        RECT 55.680 173.115 61.025 173.550 ;
        RECT 61.200 173.115 66.545 173.550 ;
        RECT 46.980 171.170 47.480 171.780 ;
        RECT 48.775 171.770 49.525 172.290 ;
        RECT 49.715 171.990 50.045 172.240 ;
        RECT 47.855 171.000 49.525 171.770 ;
        RECT 49.735 171.000 49.965 171.820 ;
        RECT 50.215 171.800 50.465 172.400 ;
        RECT 51.995 171.940 53.685 172.460 ;
        RECT 50.135 171.170 50.465 171.800 ;
        RECT 50.635 171.000 50.845 171.820 ;
        RECT 53.855 171.770 55.505 172.290 ;
        RECT 57.270 171.865 57.620 173.115 ;
        RECT 51.995 171.000 55.505 171.770 ;
        RECT 59.100 171.545 59.440 172.375 ;
        RECT 62.790 171.865 63.140 173.115 ;
        RECT 66.715 172.385 67.005 173.550 ;
        RECT 67.175 172.460 68.385 173.550 ;
        RECT 68.760 172.580 69.090 173.380 ;
        RECT 69.260 172.750 69.590 173.550 ;
        RECT 69.890 172.580 70.220 173.380 ;
        RECT 70.865 172.750 71.115 173.550 ;
        RECT 64.620 171.545 64.960 172.375 ;
        RECT 67.175 171.920 67.695 172.460 ;
        RECT 68.760 172.410 71.195 172.580 ;
        RECT 71.385 172.410 71.555 173.550 ;
        RECT 71.725 172.410 72.065 173.380 ;
        RECT 67.865 171.750 68.385 172.290 ;
        RECT 68.555 171.990 68.905 172.240 ;
        RECT 69.090 171.780 69.260 172.410 ;
        RECT 69.430 171.990 69.760 172.190 ;
        RECT 69.930 171.990 70.260 172.190 ;
        RECT 70.430 171.990 70.850 172.190 ;
        RECT 71.025 172.160 71.195 172.410 ;
        RECT 71.025 171.990 71.720 172.160 ;
        RECT 71.890 171.850 72.065 172.410 ;
        RECT 55.680 171.000 61.025 171.545 ;
        RECT 61.200 171.000 66.545 171.545 ;
        RECT 66.715 171.000 67.005 171.725 ;
        RECT 67.175 171.000 68.385 171.750 ;
        RECT 68.760 171.170 69.260 171.780 ;
        RECT 69.890 171.650 71.115 171.820 ;
        RECT 71.835 171.800 72.065 171.850 ;
        RECT 69.890 171.170 70.220 171.650 ;
        RECT 70.390 171.000 70.615 171.460 ;
        RECT 70.785 171.170 71.115 171.650 ;
        RECT 71.305 171.000 71.555 171.800 ;
        RECT 71.725 171.170 72.065 171.800 ;
        RECT 72.235 172.410 72.575 173.380 ;
        RECT 72.745 172.410 72.915 173.550 ;
        RECT 73.185 172.750 73.435 173.550 ;
        RECT 74.080 172.580 74.410 173.380 ;
        RECT 74.710 172.750 75.040 173.550 ;
        RECT 75.210 172.580 75.540 173.380 ;
        RECT 73.105 172.410 75.540 172.580 ;
        RECT 75.915 172.460 77.585 173.550 ;
        RECT 72.235 171.800 72.410 172.410 ;
        RECT 73.105 172.160 73.275 172.410 ;
        RECT 72.580 171.990 73.275 172.160 ;
        RECT 73.450 171.990 73.870 172.190 ;
        RECT 74.040 171.990 74.370 172.190 ;
        RECT 74.540 171.990 74.870 172.190 ;
        RECT 72.235 171.170 72.575 171.800 ;
        RECT 72.745 171.000 72.995 171.800 ;
        RECT 73.185 171.650 74.410 171.820 ;
        RECT 73.185 171.170 73.515 171.650 ;
        RECT 73.685 171.000 73.910 171.460 ;
        RECT 74.080 171.170 74.410 171.650 ;
        RECT 75.040 171.780 75.210 172.410 ;
        RECT 75.395 171.990 75.745 172.240 ;
        RECT 75.915 171.940 76.665 172.460 ;
        RECT 77.815 172.410 78.025 173.550 ;
        RECT 78.195 172.400 78.525 173.380 ;
        RECT 78.695 172.410 78.925 173.550 ;
        RECT 79.135 172.790 79.650 173.200 ;
        RECT 79.885 172.790 80.055 173.550 ;
        RECT 80.225 173.210 82.255 173.380 ;
        RECT 75.040 171.170 75.540 171.780 ;
        RECT 76.835 171.770 77.585 172.290 ;
        RECT 75.915 171.000 77.585 171.770 ;
        RECT 77.815 171.000 78.025 171.820 ;
        RECT 78.195 171.800 78.445 172.400 ;
        RECT 78.615 171.990 78.945 172.240 ;
        RECT 79.135 171.980 79.475 172.790 ;
        RECT 80.225 172.545 80.395 173.210 ;
        RECT 80.790 172.870 81.915 173.040 ;
        RECT 79.645 172.355 80.395 172.545 ;
        RECT 80.565 172.530 81.575 172.700 ;
        RECT 78.195 171.170 78.525 171.800 ;
        RECT 78.695 171.000 78.925 171.820 ;
        RECT 79.135 171.810 80.365 171.980 ;
        RECT 79.410 171.205 79.655 171.810 ;
        RECT 79.875 171.000 80.385 171.535 ;
        RECT 80.565 171.170 80.755 172.530 ;
        RECT 80.925 171.850 81.200 172.330 ;
        RECT 80.925 171.680 81.205 171.850 ;
        RECT 81.405 171.730 81.575 172.530 ;
        RECT 81.745 171.740 81.915 172.870 ;
        RECT 82.085 172.240 82.255 173.210 ;
        RECT 82.425 172.410 82.595 173.550 ;
        RECT 82.765 172.410 83.100 173.380 ;
        RECT 83.315 172.410 83.545 173.550 ;
        RECT 82.085 171.910 82.280 172.240 ;
        RECT 82.505 171.910 82.760 172.240 ;
        RECT 82.505 171.740 82.675 171.910 ;
        RECT 82.930 171.740 83.100 172.410 ;
        RECT 83.715 172.400 84.045 173.380 ;
        RECT 84.215 172.410 84.425 173.550 ;
        RECT 84.745 172.620 84.915 173.380 ;
        RECT 85.095 172.790 85.425 173.550 ;
        RECT 84.745 172.450 85.410 172.620 ;
        RECT 85.595 172.475 85.865 173.380 ;
        RECT 83.295 171.990 83.625 172.240 ;
        RECT 80.925 171.170 81.200 171.680 ;
        RECT 81.745 171.570 82.675 171.740 ;
        RECT 81.745 171.535 81.920 171.570 ;
        RECT 81.390 171.170 81.920 171.535 ;
        RECT 82.345 171.000 82.675 171.400 ;
        RECT 82.845 171.170 83.100 171.740 ;
        RECT 83.315 171.000 83.545 171.820 ;
        RECT 83.795 171.800 84.045 172.400 ;
        RECT 85.240 172.305 85.410 172.450 ;
        RECT 84.675 171.900 85.005 172.270 ;
        RECT 85.240 171.975 85.525 172.305 ;
        RECT 83.715 171.170 84.045 171.800 ;
        RECT 84.215 171.000 84.425 171.820 ;
        RECT 85.240 171.720 85.410 171.975 ;
        RECT 84.745 171.550 85.410 171.720 ;
        RECT 85.695 171.675 85.865 172.475 ;
        RECT 86.035 172.460 88.625 173.550 ;
        RECT 86.035 171.940 87.245 172.460 ;
        RECT 88.795 172.410 89.135 173.380 ;
        RECT 89.305 172.410 89.475 173.550 ;
        RECT 89.745 172.750 89.995 173.550 ;
        RECT 90.640 172.580 90.970 173.380 ;
        RECT 91.270 172.750 91.600 173.550 ;
        RECT 91.770 172.580 92.100 173.380 ;
        RECT 89.665 172.410 92.100 172.580 ;
        RECT 87.415 171.770 88.625 172.290 ;
        RECT 84.745 171.170 84.915 171.550 ;
        RECT 85.095 171.000 85.425 171.380 ;
        RECT 85.605 171.170 85.865 171.675 ;
        RECT 86.035 171.000 88.625 171.770 ;
        RECT 88.795 171.800 88.970 172.410 ;
        RECT 89.665 172.160 89.835 172.410 ;
        RECT 89.140 171.990 89.835 172.160 ;
        RECT 90.010 171.990 90.430 172.190 ;
        RECT 90.600 171.990 90.930 172.190 ;
        RECT 91.100 171.990 91.430 172.190 ;
        RECT 88.795 171.170 89.135 171.800 ;
        RECT 89.305 171.000 89.555 171.800 ;
        RECT 89.745 171.650 90.970 171.820 ;
        RECT 89.745 171.170 90.075 171.650 ;
        RECT 90.245 171.000 90.470 171.460 ;
        RECT 90.640 171.170 90.970 171.650 ;
        RECT 91.600 171.780 91.770 172.410 ;
        RECT 92.475 172.385 92.765 173.550 ;
        RECT 92.935 172.790 93.450 173.200 ;
        RECT 93.685 172.790 93.855 173.550 ;
        RECT 94.025 173.210 96.055 173.380 ;
        RECT 91.955 171.990 92.305 172.240 ;
        RECT 92.935 171.980 93.275 172.790 ;
        RECT 94.025 172.545 94.195 173.210 ;
        RECT 94.590 172.870 95.715 173.040 ;
        RECT 93.445 172.355 94.195 172.545 ;
        RECT 94.365 172.530 95.375 172.700 ;
        RECT 92.935 171.810 94.165 171.980 ;
        RECT 91.600 171.170 92.100 171.780 ;
        RECT 92.475 171.000 92.765 171.725 ;
        RECT 93.210 171.205 93.455 171.810 ;
        RECT 93.675 171.000 94.185 171.535 ;
        RECT 94.365 171.170 94.555 172.530 ;
        RECT 94.725 172.190 95.000 172.330 ;
        RECT 94.725 172.020 95.005 172.190 ;
        RECT 94.725 171.170 95.000 172.020 ;
        RECT 95.205 171.730 95.375 172.530 ;
        RECT 95.545 171.740 95.715 172.870 ;
        RECT 95.885 172.240 96.055 173.210 ;
        RECT 96.225 172.410 96.395 173.550 ;
        RECT 96.565 172.410 96.900 173.380 ;
        RECT 95.885 171.910 96.080 172.240 ;
        RECT 96.305 171.910 96.560 172.240 ;
        RECT 96.305 171.740 96.475 171.910 ;
        RECT 96.730 171.740 96.900 172.410 ;
        RECT 95.545 171.570 96.475 171.740 ;
        RECT 95.545 171.535 95.720 171.570 ;
        RECT 95.190 171.170 95.720 171.535 ;
        RECT 96.145 171.000 96.475 171.400 ;
        RECT 96.645 171.170 96.900 171.740 ;
        RECT 97.075 172.410 97.415 173.380 ;
        RECT 97.585 172.410 97.755 173.550 ;
        RECT 98.025 172.750 98.275 173.550 ;
        RECT 98.920 172.580 99.250 173.380 ;
        RECT 99.550 172.750 99.880 173.550 ;
        RECT 100.050 172.580 100.380 173.380 ;
        RECT 97.945 172.410 100.380 172.580 ;
        RECT 100.755 172.790 101.270 173.200 ;
        RECT 101.505 172.790 101.675 173.550 ;
        RECT 101.845 173.210 103.875 173.380 ;
        RECT 97.075 171.800 97.250 172.410 ;
        RECT 97.945 172.160 98.115 172.410 ;
        RECT 97.420 171.990 98.115 172.160 ;
        RECT 98.290 171.990 98.710 172.190 ;
        RECT 98.880 171.990 99.210 172.190 ;
        RECT 99.380 171.990 99.710 172.190 ;
        RECT 97.075 171.170 97.415 171.800 ;
        RECT 97.585 171.000 97.835 171.800 ;
        RECT 98.025 171.650 99.250 171.820 ;
        RECT 98.025 171.170 98.355 171.650 ;
        RECT 98.525 171.000 98.750 171.460 ;
        RECT 98.920 171.170 99.250 171.650 ;
        RECT 99.880 171.780 100.050 172.410 ;
        RECT 100.235 171.990 100.585 172.240 ;
        RECT 100.755 171.980 101.095 172.790 ;
        RECT 101.845 172.545 102.015 173.210 ;
        RECT 102.410 172.870 103.535 173.040 ;
        RECT 101.265 172.355 102.015 172.545 ;
        RECT 102.185 172.530 103.195 172.700 ;
        RECT 100.755 171.810 101.985 171.980 ;
        RECT 99.880 171.170 100.380 171.780 ;
        RECT 101.030 171.205 101.275 171.810 ;
        RECT 101.495 171.000 102.005 171.535 ;
        RECT 102.185 171.170 102.375 172.530 ;
        RECT 102.545 172.190 102.820 172.330 ;
        RECT 102.545 172.020 102.825 172.190 ;
        RECT 102.545 171.170 102.820 172.020 ;
        RECT 103.025 171.730 103.195 172.530 ;
        RECT 103.365 171.740 103.535 172.870 ;
        RECT 103.705 172.240 103.875 173.210 ;
        RECT 104.045 172.410 104.215 173.550 ;
        RECT 104.385 172.410 104.720 173.380 ;
        RECT 105.270 172.570 105.525 173.240 ;
        RECT 105.705 172.750 105.990 173.550 ;
        RECT 106.170 172.830 106.500 173.340 ;
        RECT 105.270 172.530 105.450 172.570 ;
        RECT 103.705 171.910 103.900 172.240 ;
        RECT 104.125 171.910 104.380 172.240 ;
        RECT 104.125 171.740 104.295 171.910 ;
        RECT 104.550 171.740 104.720 172.410 ;
        RECT 105.185 172.360 105.450 172.530 ;
        RECT 103.365 171.570 104.295 171.740 ;
        RECT 103.365 171.535 103.540 171.570 ;
        RECT 103.010 171.170 103.540 171.535 ;
        RECT 103.965 171.000 104.295 171.400 ;
        RECT 104.465 171.170 104.720 171.740 ;
        RECT 105.270 171.710 105.450 172.360 ;
        RECT 106.170 172.240 106.420 172.830 ;
        RECT 106.770 172.680 106.940 173.290 ;
        RECT 107.110 172.860 107.440 173.550 ;
        RECT 107.670 173.000 107.910 173.290 ;
        RECT 108.110 173.170 108.530 173.550 ;
        RECT 108.710 173.080 109.340 173.330 ;
        RECT 109.810 173.170 110.140 173.550 ;
        RECT 108.710 173.000 108.880 173.080 ;
        RECT 110.310 173.000 110.480 173.290 ;
        RECT 110.660 173.170 111.040 173.550 ;
        RECT 111.280 173.165 112.110 173.335 ;
        RECT 107.670 172.830 108.880 173.000 ;
        RECT 105.620 171.910 106.420 172.240 ;
        RECT 105.270 171.180 105.525 171.710 ;
        RECT 105.705 171.000 105.990 171.460 ;
        RECT 106.170 171.260 106.420 171.910 ;
        RECT 106.620 172.660 106.940 172.680 ;
        RECT 106.620 172.490 108.540 172.660 ;
        RECT 106.620 171.595 106.810 172.490 ;
        RECT 108.710 172.320 108.880 172.830 ;
        RECT 109.050 172.570 109.570 172.880 ;
        RECT 106.980 172.150 108.880 172.320 ;
        RECT 106.980 172.090 107.310 172.150 ;
        RECT 107.460 171.920 107.790 171.980 ;
        RECT 107.130 171.650 107.790 171.920 ;
        RECT 106.620 171.265 106.940 171.595 ;
        RECT 107.120 171.000 107.780 171.480 ;
        RECT 107.980 171.390 108.150 172.150 ;
        RECT 109.050 171.980 109.230 172.390 ;
        RECT 108.320 171.810 108.650 171.930 ;
        RECT 109.400 171.810 109.570 172.570 ;
        RECT 108.320 171.640 109.570 171.810 ;
        RECT 109.740 172.750 111.110 173.000 ;
        RECT 109.740 171.980 109.930 172.750 ;
        RECT 110.860 172.490 111.110 172.750 ;
        RECT 110.100 172.320 110.350 172.480 ;
        RECT 111.280 172.320 111.450 173.165 ;
        RECT 112.345 172.880 112.515 173.380 ;
        RECT 112.685 173.050 113.015 173.550 ;
        RECT 111.620 172.490 112.120 172.870 ;
        RECT 112.345 172.710 113.040 172.880 ;
        RECT 110.100 172.150 111.450 172.320 ;
        RECT 111.030 172.110 111.450 172.150 ;
        RECT 109.740 171.640 110.160 171.980 ;
        RECT 110.450 171.650 110.860 171.980 ;
        RECT 107.980 171.220 108.830 171.390 ;
        RECT 109.390 171.000 109.710 171.460 ;
        RECT 109.910 171.210 110.160 171.640 ;
        RECT 110.450 171.000 110.860 171.440 ;
        RECT 111.030 171.380 111.200 172.110 ;
        RECT 111.370 171.560 111.720 171.930 ;
        RECT 111.900 171.620 112.120 172.490 ;
        RECT 112.290 171.920 112.700 172.540 ;
        RECT 112.870 171.740 113.040 172.710 ;
        RECT 112.345 171.550 113.040 171.740 ;
        RECT 111.030 171.180 112.045 171.380 ;
        RECT 112.345 171.220 112.515 171.550 ;
        RECT 112.685 171.000 113.015 171.380 ;
        RECT 113.230 171.260 113.455 173.380 ;
        RECT 113.625 173.050 113.955 173.550 ;
        RECT 114.125 172.880 114.295 173.380 ;
        RECT 114.560 173.125 114.895 173.550 ;
        RECT 115.065 172.945 115.250 173.350 ;
        RECT 113.630 172.710 114.295 172.880 ;
        RECT 114.585 172.770 115.250 172.945 ;
        RECT 115.455 172.770 115.785 173.550 ;
        RECT 113.630 171.720 113.860 172.710 ;
        RECT 114.030 171.890 114.380 172.540 ;
        RECT 114.585 171.740 114.925 172.770 ;
        RECT 115.955 172.580 116.225 173.350 ;
        RECT 115.095 172.410 116.225 172.580 ;
        RECT 115.095 171.910 115.345 172.410 ;
        RECT 113.630 171.550 114.295 171.720 ;
        RECT 114.585 171.570 115.270 171.740 ;
        RECT 115.525 171.660 115.885 172.240 ;
        RECT 113.625 171.000 113.955 171.380 ;
        RECT 114.125 171.260 114.295 171.550 ;
        RECT 114.560 171.000 114.895 171.400 ;
        RECT 115.065 171.170 115.270 171.570 ;
        RECT 116.055 171.500 116.225 172.410 ;
        RECT 117.315 172.460 118.525 173.550 ;
        RECT 117.315 171.920 117.835 172.460 ;
        RECT 118.005 171.750 118.525 172.290 ;
        RECT 115.480 171.000 115.755 171.480 ;
        RECT 115.965 171.170 116.225 171.500 ;
        RECT 117.315 171.000 118.525 171.750 ;
        RECT 11.430 170.830 118.610 171.000 ;
        RECT 11.515 170.080 12.725 170.830 ;
        RECT 11.515 169.540 12.035 170.080 ;
        RECT 13.415 170.010 13.625 170.830 ;
        RECT 13.795 170.030 14.125 170.660 ;
        RECT 12.205 169.370 12.725 169.910 ;
        RECT 13.795 169.430 14.045 170.030 ;
        RECT 14.295 170.010 14.525 170.830 ;
        RECT 15.010 170.020 15.255 170.625 ;
        RECT 15.475 170.295 15.985 170.830 ;
        RECT 14.735 169.850 15.965 170.020 ;
        RECT 14.215 169.590 14.545 169.840 ;
        RECT 11.515 168.280 12.725 169.370 ;
        RECT 13.415 168.280 13.625 169.420 ;
        RECT 13.795 168.450 14.125 169.430 ;
        RECT 14.295 168.280 14.525 169.420 ;
        RECT 14.735 169.040 15.075 169.850 ;
        RECT 15.245 169.285 15.995 169.475 ;
        RECT 14.735 168.630 15.250 169.040 ;
        RECT 15.485 168.280 15.655 169.040 ;
        RECT 15.825 168.620 15.995 169.285 ;
        RECT 16.165 169.300 16.355 170.660 ;
        RECT 16.525 170.150 16.800 170.660 ;
        RECT 16.990 170.295 17.520 170.660 ;
        RECT 17.945 170.430 18.275 170.830 ;
        RECT 17.345 170.260 17.520 170.295 ;
        RECT 16.525 169.980 16.805 170.150 ;
        RECT 16.525 169.500 16.800 169.980 ;
        RECT 17.005 169.300 17.175 170.100 ;
        RECT 16.165 169.130 17.175 169.300 ;
        RECT 17.345 170.090 18.275 170.260 ;
        RECT 18.445 170.090 18.700 170.660 ;
        RECT 18.965 170.350 19.265 170.830 ;
        RECT 19.435 170.180 19.695 170.635 ;
        RECT 19.865 170.350 20.125 170.830 ;
        RECT 20.305 170.180 20.565 170.635 ;
        RECT 20.735 170.350 20.985 170.830 ;
        RECT 21.165 170.180 21.425 170.635 ;
        RECT 21.595 170.350 21.845 170.830 ;
        RECT 22.025 170.180 22.285 170.635 ;
        RECT 22.455 170.350 22.700 170.830 ;
        RECT 22.870 170.180 23.145 170.635 ;
        RECT 23.315 170.350 23.560 170.830 ;
        RECT 23.730 170.180 23.990 170.635 ;
        RECT 24.160 170.350 24.420 170.830 ;
        RECT 24.590 170.180 24.850 170.635 ;
        RECT 25.020 170.350 25.280 170.830 ;
        RECT 25.450 170.180 25.710 170.635 ;
        RECT 25.880 170.270 26.140 170.830 ;
        RECT 17.345 168.960 17.515 170.090 ;
        RECT 18.105 169.920 18.275 170.090 ;
        RECT 16.390 168.790 17.515 168.960 ;
        RECT 17.685 169.590 17.880 169.920 ;
        RECT 18.105 169.590 18.360 169.920 ;
        RECT 17.685 168.620 17.855 169.590 ;
        RECT 18.530 169.420 18.700 170.090 ;
        RECT 15.825 168.450 17.855 168.620 ;
        RECT 18.025 168.280 18.195 169.420 ;
        RECT 18.365 168.450 18.700 169.420 ;
        RECT 18.965 170.010 25.710 170.180 ;
        RECT 18.965 169.420 20.130 170.010 ;
        RECT 26.310 169.840 26.560 170.650 ;
        RECT 26.740 170.305 27.000 170.830 ;
        RECT 27.170 169.840 27.420 170.650 ;
        RECT 27.600 170.320 27.905 170.830 ;
        RECT 20.300 169.590 27.420 169.840 ;
        RECT 27.590 169.590 27.905 170.150 ;
        RECT 28.075 170.105 28.365 170.830 ;
        RECT 28.540 170.360 28.870 170.830 ;
        RECT 29.040 170.190 29.265 170.635 ;
        RECT 29.435 170.305 29.730 170.830 ;
        RECT 28.535 170.020 29.265 170.190 ;
        RECT 18.965 169.195 25.710 169.420 ;
        RECT 18.965 168.280 19.235 169.025 ;
        RECT 19.405 168.455 19.695 169.195 ;
        RECT 20.305 169.180 25.710 169.195 ;
        RECT 19.865 168.285 20.120 169.010 ;
        RECT 20.305 168.455 20.565 169.180 ;
        RECT 20.735 168.285 20.980 169.010 ;
        RECT 21.165 168.455 21.425 169.180 ;
        RECT 21.595 168.285 21.840 169.010 ;
        RECT 22.025 168.455 22.285 169.180 ;
        RECT 22.455 168.285 22.700 169.010 ;
        RECT 22.870 168.455 23.130 169.180 ;
        RECT 23.300 168.285 23.560 169.010 ;
        RECT 23.730 168.455 23.990 169.180 ;
        RECT 24.160 168.285 24.420 169.010 ;
        RECT 24.590 168.455 24.850 169.180 ;
        RECT 25.020 168.285 25.280 169.010 ;
        RECT 25.450 168.455 25.710 169.180 ;
        RECT 25.880 168.285 26.140 169.080 ;
        RECT 26.310 168.455 26.560 169.590 ;
        RECT 19.865 168.280 26.140 168.285 ;
        RECT 26.740 168.280 27.000 169.090 ;
        RECT 27.175 168.450 27.420 169.590 ;
        RECT 28.535 169.455 28.815 170.020 ;
        RECT 30.415 170.010 30.645 170.830 ;
        RECT 30.815 170.030 31.145 170.660 ;
        RECT 28.985 169.625 30.205 169.850 ;
        RECT 30.395 169.590 30.725 169.840 ;
        RECT 27.600 168.280 27.895 169.090 ;
        RECT 28.075 168.280 28.365 169.445 ;
        RECT 28.535 169.285 30.135 169.455 ;
        RECT 30.895 169.430 31.145 170.030 ;
        RECT 31.315 170.010 31.525 170.830 ;
        RECT 32.735 170.350 33.015 170.830 ;
        RECT 33.185 170.180 33.445 170.570 ;
        RECT 33.620 170.350 33.875 170.830 ;
        RECT 34.045 170.180 34.340 170.570 ;
        RECT 34.520 170.350 34.795 170.830 ;
        RECT 34.965 170.330 35.265 170.660 ;
        RECT 32.690 170.010 34.340 170.180 ;
        RECT 28.595 168.280 28.850 169.115 ;
        RECT 29.020 168.480 29.280 169.285 ;
        RECT 29.450 168.280 29.710 169.115 ;
        RECT 29.880 168.480 30.135 169.285 ;
        RECT 30.415 168.280 30.645 169.420 ;
        RECT 30.815 168.450 31.145 169.430 ;
        RECT 32.690 169.500 33.095 170.010 ;
        RECT 33.265 169.670 34.405 169.840 ;
        RECT 31.315 168.280 31.525 169.420 ;
        RECT 32.690 169.330 33.445 169.500 ;
        RECT 32.730 168.280 33.015 169.150 ;
        RECT 33.185 169.080 33.445 169.330 ;
        RECT 34.235 169.420 34.405 169.670 ;
        RECT 34.575 169.590 34.925 170.160 ;
        RECT 35.095 169.420 35.265 170.330 ;
        RECT 35.585 170.030 35.915 170.830 ;
        RECT 36.085 170.180 36.255 170.660 ;
        RECT 36.425 170.350 36.755 170.830 ;
        RECT 36.925 170.180 37.095 170.660 ;
        RECT 37.345 170.350 37.585 170.830 ;
        RECT 37.765 170.180 37.935 170.660 ;
        RECT 36.085 170.010 37.095 170.180 ;
        RECT 37.300 170.010 37.935 170.180 ;
        RECT 38.195 170.060 40.785 170.830 ;
        RECT 36.085 169.810 36.580 170.010 ;
        RECT 37.300 169.840 37.470 170.010 ;
        RECT 36.085 169.640 36.585 169.810 ;
        RECT 36.970 169.670 37.470 169.840 ;
        RECT 36.085 169.470 36.580 169.640 ;
        RECT 34.235 169.250 35.265 169.420 ;
        RECT 33.185 168.910 34.305 169.080 ;
        RECT 33.185 168.450 33.445 168.910 ;
        RECT 33.620 168.280 33.875 168.740 ;
        RECT 34.045 168.450 34.305 168.910 ;
        RECT 34.475 168.280 34.785 169.080 ;
        RECT 34.955 168.450 35.265 169.250 ;
        RECT 35.585 168.280 35.915 169.430 ;
        RECT 36.085 169.300 37.095 169.470 ;
        RECT 36.085 168.450 36.255 169.300 ;
        RECT 36.425 168.280 36.755 169.080 ;
        RECT 36.925 168.450 37.095 169.300 ;
        RECT 37.300 169.430 37.470 169.670 ;
        RECT 37.640 169.600 38.020 169.840 ;
        RECT 37.300 169.260 38.015 169.430 ;
        RECT 37.275 168.280 37.515 169.080 ;
        RECT 37.685 168.450 38.015 169.260 ;
        RECT 38.195 169.370 39.405 169.890 ;
        RECT 39.575 169.540 40.785 170.060 ;
        RECT 40.955 170.030 41.295 170.660 ;
        RECT 41.465 170.030 41.715 170.830 ;
        RECT 41.905 170.180 42.235 170.660 ;
        RECT 42.405 170.370 42.630 170.830 ;
        RECT 42.800 170.180 43.130 170.660 ;
        RECT 40.955 169.420 41.130 170.030 ;
        RECT 41.905 170.010 43.130 170.180 ;
        RECT 43.760 170.050 44.260 170.660 ;
        RECT 44.640 170.280 44.895 170.570 ;
        RECT 45.065 170.450 45.395 170.830 ;
        RECT 44.640 170.110 45.390 170.280 ;
        RECT 41.300 169.670 41.995 169.840 ;
        RECT 41.825 169.420 41.995 169.670 ;
        RECT 42.170 169.640 42.590 169.840 ;
        RECT 42.760 169.640 43.090 169.840 ;
        RECT 43.260 169.640 43.590 169.840 ;
        RECT 43.760 169.420 43.930 170.050 ;
        RECT 44.115 169.590 44.465 169.840 ;
        RECT 38.195 168.280 40.785 169.370 ;
        RECT 40.955 168.450 41.295 169.420 ;
        RECT 41.465 168.280 41.635 169.420 ;
        RECT 41.825 169.250 44.260 169.420 ;
        RECT 44.640 169.290 44.990 169.940 ;
        RECT 41.905 168.280 42.155 169.080 ;
        RECT 42.800 168.450 43.130 169.250 ;
        RECT 43.430 168.280 43.760 169.080 ;
        RECT 43.930 168.450 44.260 169.250 ;
        RECT 45.160 169.120 45.390 170.110 ;
        RECT 44.640 168.950 45.390 169.120 ;
        RECT 44.640 168.450 44.895 168.950 ;
        RECT 45.065 168.280 45.395 168.780 ;
        RECT 45.565 168.450 45.735 170.570 ;
        RECT 46.095 170.470 46.425 170.830 ;
        RECT 46.595 170.440 47.090 170.610 ;
        RECT 47.295 170.440 48.150 170.610 ;
        RECT 45.965 169.250 46.425 170.300 ;
        RECT 45.905 168.465 46.230 169.250 ;
        RECT 46.595 169.080 46.765 170.440 ;
        RECT 46.935 169.530 47.285 170.150 ;
        RECT 47.455 169.930 47.810 170.150 ;
        RECT 47.455 169.340 47.625 169.930 ;
        RECT 47.980 169.730 48.150 170.440 ;
        RECT 49.025 170.370 49.355 170.830 ;
        RECT 49.565 170.470 49.915 170.640 ;
        RECT 48.355 169.900 49.145 170.150 ;
        RECT 49.565 170.080 49.825 170.470 ;
        RECT 50.135 170.380 51.085 170.660 ;
        RECT 51.255 170.390 51.445 170.830 ;
        RECT 51.615 170.450 52.685 170.620 ;
        RECT 49.315 169.730 49.485 169.910 ;
        RECT 46.595 168.910 46.990 169.080 ;
        RECT 47.160 168.950 47.625 169.340 ;
        RECT 47.795 169.560 49.485 169.730 ;
        RECT 46.820 168.780 46.990 168.910 ;
        RECT 47.795 168.780 47.965 169.560 ;
        RECT 49.655 169.390 49.825 170.080 ;
        RECT 48.325 169.220 49.825 169.390 ;
        RECT 50.015 169.420 50.225 170.210 ;
        RECT 50.395 169.590 50.745 170.210 ;
        RECT 50.915 169.600 51.085 170.380 ;
        RECT 51.615 170.220 51.785 170.450 ;
        RECT 51.255 170.050 51.785 170.220 ;
        RECT 51.255 169.770 51.475 170.050 ;
        RECT 51.955 169.880 52.195 170.280 ;
        RECT 50.915 169.430 51.320 169.600 ;
        RECT 51.655 169.510 52.195 169.880 ;
        RECT 52.365 170.095 52.685 170.450 ;
        RECT 52.930 170.370 53.235 170.830 ;
        RECT 53.405 170.120 53.660 170.650 ;
        RECT 52.365 169.920 52.690 170.095 ;
        RECT 52.365 169.620 53.280 169.920 ;
        RECT 52.540 169.590 53.280 169.620 ;
        RECT 50.015 169.260 50.690 169.420 ;
        RECT 51.150 169.340 51.320 169.430 ;
        RECT 50.015 169.250 50.980 169.260 ;
        RECT 49.655 169.080 49.825 169.220 ;
        RECT 46.400 168.280 46.650 168.740 ;
        RECT 46.820 168.450 47.070 168.780 ;
        RECT 47.285 168.450 47.965 168.780 ;
        RECT 48.135 168.880 49.210 169.050 ;
        RECT 49.655 168.910 50.215 169.080 ;
        RECT 50.520 168.960 50.980 169.250 ;
        RECT 51.150 169.170 52.370 169.340 ;
        RECT 48.135 168.540 48.305 168.880 ;
        RECT 48.540 168.280 48.870 168.710 ;
        RECT 49.040 168.540 49.210 168.880 ;
        RECT 49.505 168.280 49.875 168.740 ;
        RECT 50.045 168.450 50.215 168.910 ;
        RECT 51.150 168.790 51.320 169.170 ;
        RECT 52.540 169.000 52.710 169.590 ;
        RECT 53.450 169.470 53.660 170.120 ;
        RECT 53.835 170.105 54.125 170.830 ;
        RECT 54.755 170.060 58.265 170.830 ;
        RECT 50.450 168.450 51.320 168.790 ;
        RECT 51.910 168.830 52.710 169.000 ;
        RECT 51.490 168.280 51.740 168.740 ;
        RECT 51.910 168.540 52.080 168.830 ;
        RECT 52.260 168.280 52.590 168.660 ;
        RECT 52.930 168.280 53.235 169.420 ;
        RECT 53.405 168.590 53.660 169.470 ;
        RECT 53.835 168.280 54.125 169.445 ;
        RECT 54.755 169.370 56.445 169.890 ;
        RECT 56.615 169.540 58.265 170.060 ;
        RECT 58.495 170.010 58.705 170.830 ;
        RECT 58.875 170.030 59.205 170.660 ;
        RECT 58.875 169.430 59.125 170.030 ;
        RECT 59.375 170.010 59.605 170.830 ;
        RECT 60.825 170.280 60.995 170.660 ;
        RECT 61.210 170.450 61.540 170.830 ;
        RECT 60.825 170.110 61.540 170.280 ;
        RECT 59.295 169.590 59.625 169.840 ;
        RECT 60.735 169.560 61.090 169.930 ;
        RECT 61.370 169.920 61.540 170.110 ;
        RECT 61.710 170.085 61.965 170.660 ;
        RECT 61.370 169.590 61.625 169.920 ;
        RECT 54.755 168.280 58.265 169.370 ;
        RECT 58.495 168.280 58.705 169.420 ;
        RECT 58.875 168.450 59.205 169.430 ;
        RECT 59.375 168.280 59.605 169.420 ;
        RECT 61.370 169.380 61.540 169.590 ;
        RECT 60.825 169.210 61.540 169.380 ;
        RECT 61.795 169.355 61.965 170.085 ;
        RECT 62.140 169.990 62.400 170.830 ;
        RECT 62.635 170.350 62.915 170.830 ;
        RECT 63.085 170.180 63.345 170.570 ;
        RECT 63.520 170.350 63.775 170.830 ;
        RECT 63.945 170.180 64.240 170.570 ;
        RECT 64.420 170.350 64.695 170.830 ;
        RECT 64.865 170.330 65.165 170.660 ;
        RECT 62.590 170.010 64.240 170.180 ;
        RECT 62.590 169.500 62.995 170.010 ;
        RECT 63.165 169.670 64.305 169.840 ;
        RECT 60.825 168.450 60.995 169.210 ;
        RECT 61.210 168.280 61.540 169.040 ;
        RECT 61.710 168.450 61.965 169.355 ;
        RECT 62.140 168.280 62.400 169.430 ;
        RECT 62.590 169.330 63.345 169.500 ;
        RECT 62.630 168.280 62.915 169.150 ;
        RECT 63.085 169.080 63.345 169.330 ;
        RECT 64.135 169.420 64.305 169.670 ;
        RECT 64.475 169.590 64.825 170.160 ;
        RECT 64.995 169.420 65.165 170.330 ;
        RECT 65.335 170.080 66.545 170.830 ;
        RECT 64.135 169.250 65.165 169.420 ;
        RECT 63.085 168.910 64.205 169.080 ;
        RECT 63.085 168.450 63.345 168.910 ;
        RECT 63.520 168.280 63.775 168.740 ;
        RECT 63.945 168.450 64.205 168.910 ;
        RECT 64.375 168.280 64.685 169.080 ;
        RECT 64.855 168.450 65.165 169.250 ;
        RECT 65.335 169.370 65.855 169.910 ;
        RECT 66.025 169.540 66.545 170.080 ;
        RECT 66.775 170.010 66.985 170.830 ;
        RECT 67.155 170.030 67.485 170.660 ;
        RECT 67.155 169.430 67.405 170.030 ;
        RECT 67.655 170.010 67.885 170.830 ;
        RECT 68.300 170.050 68.800 170.660 ;
        RECT 67.575 169.590 67.905 169.840 ;
        RECT 68.095 169.590 68.445 169.840 ;
        RECT 65.335 168.280 66.545 169.370 ;
        RECT 66.775 168.280 66.985 169.420 ;
        RECT 67.155 168.450 67.485 169.430 ;
        RECT 68.630 169.420 68.800 170.050 ;
        RECT 69.430 170.180 69.760 170.660 ;
        RECT 69.930 170.370 70.155 170.830 ;
        RECT 70.325 170.180 70.655 170.660 ;
        RECT 69.430 170.010 70.655 170.180 ;
        RECT 70.845 170.030 71.095 170.830 ;
        RECT 71.265 170.030 71.605 170.660 ;
        RECT 68.970 169.640 69.300 169.840 ;
        RECT 69.470 169.640 69.800 169.840 ;
        RECT 69.970 169.640 70.390 169.840 ;
        RECT 70.565 169.670 71.260 169.840 ;
        RECT 70.565 169.420 70.735 169.670 ;
        RECT 71.430 169.420 71.605 170.030 ;
        RECT 67.655 168.280 67.885 169.420 ;
        RECT 68.300 169.250 70.735 169.420 ;
        RECT 68.300 168.450 68.630 169.250 ;
        RECT 68.800 168.280 69.130 169.080 ;
        RECT 69.430 168.450 69.760 169.250 ;
        RECT 70.405 168.280 70.655 169.080 ;
        RECT 70.925 168.280 71.095 169.420 ;
        RECT 71.265 168.450 71.605 169.420 ;
        RECT 71.775 170.030 72.115 170.660 ;
        RECT 72.285 170.030 72.535 170.830 ;
        RECT 72.725 170.180 73.055 170.660 ;
        RECT 73.225 170.370 73.450 170.830 ;
        RECT 73.620 170.180 73.950 170.660 ;
        RECT 71.775 169.420 71.950 170.030 ;
        RECT 72.725 170.010 73.950 170.180 ;
        RECT 74.580 170.050 75.080 170.660 ;
        RECT 72.120 169.670 72.815 169.840 ;
        RECT 72.645 169.420 72.815 169.670 ;
        RECT 72.990 169.640 73.410 169.840 ;
        RECT 73.580 169.640 73.910 169.840 ;
        RECT 74.080 169.640 74.410 169.840 ;
        RECT 74.580 169.420 74.750 170.050 ;
        RECT 75.730 170.020 75.975 170.625 ;
        RECT 76.195 170.295 76.705 170.830 ;
        RECT 75.455 169.850 76.685 170.020 ;
        RECT 74.935 169.590 75.285 169.840 ;
        RECT 71.775 168.450 72.115 169.420 ;
        RECT 72.285 168.280 72.455 169.420 ;
        RECT 72.645 169.250 75.080 169.420 ;
        RECT 72.725 168.280 72.975 169.080 ;
        RECT 73.620 168.450 73.950 169.250 ;
        RECT 74.250 168.280 74.580 169.080 ;
        RECT 74.750 168.450 75.080 169.250 ;
        RECT 75.455 169.040 75.795 169.850 ;
        RECT 75.965 169.285 76.715 169.475 ;
        RECT 75.455 168.630 75.970 169.040 ;
        RECT 76.205 168.280 76.375 169.040 ;
        RECT 76.545 168.620 76.715 169.285 ;
        RECT 76.885 169.300 77.075 170.660 ;
        RECT 77.245 169.810 77.520 170.660 ;
        RECT 77.710 170.295 78.240 170.660 ;
        RECT 78.665 170.430 78.995 170.830 ;
        RECT 78.065 170.260 78.240 170.295 ;
        RECT 77.245 169.640 77.525 169.810 ;
        RECT 77.245 169.500 77.520 169.640 ;
        RECT 77.725 169.300 77.895 170.100 ;
        RECT 76.885 169.130 77.895 169.300 ;
        RECT 78.065 170.090 78.995 170.260 ;
        RECT 79.165 170.090 79.420 170.660 ;
        RECT 79.595 170.105 79.885 170.830 ;
        RECT 80.430 170.120 80.685 170.650 ;
        RECT 80.865 170.370 81.150 170.830 ;
        RECT 78.065 168.960 78.235 170.090 ;
        RECT 78.825 169.920 78.995 170.090 ;
        RECT 77.110 168.790 78.235 168.960 ;
        RECT 78.405 169.590 78.600 169.920 ;
        RECT 78.825 169.590 79.080 169.920 ;
        RECT 78.405 168.620 78.575 169.590 ;
        RECT 79.250 169.420 79.420 170.090 ;
        RECT 80.430 169.810 80.610 170.120 ;
        RECT 81.330 169.920 81.580 170.570 ;
        RECT 80.345 169.640 80.610 169.810 ;
        RECT 76.545 168.450 78.575 168.620 ;
        RECT 78.745 168.280 78.915 169.420 ;
        RECT 79.085 168.450 79.420 169.420 ;
        RECT 79.595 168.280 79.885 169.445 ;
        RECT 80.430 169.260 80.610 169.640 ;
        RECT 80.780 169.590 81.580 169.920 ;
        RECT 80.430 168.590 80.685 169.260 ;
        RECT 80.865 168.280 81.150 169.080 ;
        RECT 81.330 169.000 81.580 169.590 ;
        RECT 81.780 170.235 82.100 170.565 ;
        RECT 82.280 170.350 82.940 170.830 ;
        RECT 83.140 170.440 83.990 170.610 ;
        RECT 81.780 169.340 81.970 170.235 ;
        RECT 82.290 169.910 82.950 170.180 ;
        RECT 82.620 169.850 82.950 169.910 ;
        RECT 82.140 169.680 82.470 169.740 ;
        RECT 83.140 169.680 83.310 170.440 ;
        RECT 84.550 170.370 84.870 170.830 ;
        RECT 85.070 170.190 85.320 170.620 ;
        RECT 85.610 170.390 86.020 170.830 ;
        RECT 86.190 170.450 87.205 170.650 ;
        RECT 83.480 170.020 84.730 170.190 ;
        RECT 83.480 169.900 83.810 170.020 ;
        RECT 82.140 169.510 84.040 169.680 ;
        RECT 81.780 169.170 83.700 169.340 ;
        RECT 81.780 169.150 82.100 169.170 ;
        RECT 81.330 168.490 81.660 169.000 ;
        RECT 81.930 168.540 82.100 169.150 ;
        RECT 83.870 169.000 84.040 169.510 ;
        RECT 84.210 169.440 84.390 169.850 ;
        RECT 84.560 169.260 84.730 170.020 ;
        RECT 82.270 168.280 82.600 168.970 ;
        RECT 82.830 168.830 84.040 169.000 ;
        RECT 84.210 168.950 84.730 169.260 ;
        RECT 84.900 169.850 85.320 170.190 ;
        RECT 85.610 169.850 86.020 170.180 ;
        RECT 84.900 169.080 85.090 169.850 ;
        RECT 86.190 169.720 86.360 170.450 ;
        RECT 87.505 170.280 87.675 170.610 ;
        RECT 87.845 170.450 88.175 170.830 ;
        RECT 86.530 169.900 86.880 170.270 ;
        RECT 86.190 169.680 86.610 169.720 ;
        RECT 85.260 169.510 86.610 169.680 ;
        RECT 85.260 169.350 85.510 169.510 ;
        RECT 86.020 169.080 86.270 169.340 ;
        RECT 84.900 168.830 86.270 169.080 ;
        RECT 82.830 168.540 83.070 168.830 ;
        RECT 83.870 168.750 84.040 168.830 ;
        RECT 83.270 168.280 83.690 168.660 ;
        RECT 83.870 168.500 84.500 168.750 ;
        RECT 84.970 168.280 85.300 168.660 ;
        RECT 85.470 168.540 85.640 168.830 ;
        RECT 86.440 168.665 86.610 169.510 ;
        RECT 87.060 169.340 87.280 170.210 ;
        RECT 87.505 170.090 88.200 170.280 ;
        RECT 86.780 168.960 87.280 169.340 ;
        RECT 87.450 169.290 87.860 169.910 ;
        RECT 88.030 169.120 88.200 170.090 ;
        RECT 87.505 168.950 88.200 169.120 ;
        RECT 85.820 168.280 86.200 168.660 ;
        RECT 86.440 168.495 87.270 168.665 ;
        RECT 87.505 168.450 87.675 168.950 ;
        RECT 87.845 168.280 88.175 168.780 ;
        RECT 88.390 168.450 88.615 170.570 ;
        RECT 88.785 170.450 89.115 170.830 ;
        RECT 89.285 170.280 89.455 170.570 ;
        RECT 88.790 170.110 89.455 170.280 ;
        RECT 88.790 169.120 89.020 170.110 ;
        RECT 90.175 170.060 92.765 170.830 ;
        RECT 89.190 169.290 89.540 169.940 ;
        RECT 90.175 169.370 91.385 169.890 ;
        RECT 91.555 169.540 92.765 170.060 ;
        RECT 92.995 170.010 93.205 170.830 ;
        RECT 93.375 170.030 93.705 170.660 ;
        RECT 93.375 169.430 93.625 170.030 ;
        RECT 93.875 170.010 94.105 170.830 ;
        RECT 94.315 170.060 95.985 170.830 ;
        RECT 96.245 170.280 96.415 170.660 ;
        RECT 96.595 170.450 96.925 170.830 ;
        RECT 96.245 170.110 96.910 170.280 ;
        RECT 97.105 170.155 97.365 170.660 ;
        RECT 93.795 169.590 94.125 169.840 ;
        RECT 88.790 168.950 89.455 169.120 ;
        RECT 88.785 168.280 89.115 168.780 ;
        RECT 89.285 168.450 89.455 168.950 ;
        RECT 90.175 168.280 92.765 169.370 ;
        RECT 92.995 168.280 93.205 169.420 ;
        RECT 93.375 168.450 93.705 169.430 ;
        RECT 93.875 168.280 94.105 169.420 ;
        RECT 94.315 169.370 95.065 169.890 ;
        RECT 95.235 169.540 95.985 170.060 ;
        RECT 96.175 169.560 96.505 169.930 ;
        RECT 96.740 169.855 96.910 170.110 ;
        RECT 96.740 169.525 97.025 169.855 ;
        RECT 96.740 169.380 96.910 169.525 ;
        RECT 94.315 168.280 95.985 169.370 ;
        RECT 96.245 169.210 96.910 169.380 ;
        RECT 97.195 169.355 97.365 170.155 ;
        RECT 97.995 170.060 99.665 170.830 ;
        RECT 99.840 170.285 105.185 170.830 ;
        RECT 96.245 168.450 96.415 169.210 ;
        RECT 96.595 168.280 96.925 169.040 ;
        RECT 97.095 168.450 97.365 169.355 ;
        RECT 97.995 169.370 98.745 169.890 ;
        RECT 98.915 169.540 99.665 170.060 ;
        RECT 97.995 168.280 99.665 169.370 ;
        RECT 101.430 168.715 101.780 169.965 ;
        RECT 103.260 169.455 103.600 170.285 ;
        RECT 105.355 170.105 105.645 170.830 ;
        RECT 106.315 170.010 106.545 170.830 ;
        RECT 106.715 170.030 107.045 170.660 ;
        RECT 106.295 169.590 106.625 169.840 ;
        RECT 99.840 168.280 105.185 168.715 ;
        RECT 105.355 168.280 105.645 169.445 ;
        RECT 106.795 169.430 107.045 170.030 ;
        RECT 107.215 170.010 107.425 170.830 ;
        RECT 107.805 170.030 108.135 170.830 ;
        RECT 108.305 170.180 108.475 170.660 ;
        RECT 108.645 170.350 108.975 170.830 ;
        RECT 109.145 170.180 109.315 170.660 ;
        RECT 109.565 170.350 109.805 170.830 ;
        RECT 109.985 170.180 110.155 170.660 ;
        RECT 108.305 170.010 109.315 170.180 ;
        RECT 109.520 170.010 110.155 170.180 ;
        RECT 110.505 170.280 110.675 170.660 ;
        RECT 110.855 170.450 111.185 170.830 ;
        RECT 110.505 170.110 111.170 170.280 ;
        RECT 111.365 170.155 111.625 170.660 ;
        RECT 111.800 170.285 117.145 170.830 ;
        RECT 108.305 169.810 108.800 170.010 ;
        RECT 109.520 169.840 109.690 170.010 ;
        RECT 108.305 169.640 108.805 169.810 ;
        RECT 109.190 169.670 109.690 169.840 ;
        RECT 108.305 169.470 108.800 169.640 ;
        RECT 106.315 168.280 106.545 169.420 ;
        RECT 106.715 168.450 107.045 169.430 ;
        RECT 107.215 168.280 107.425 169.420 ;
        RECT 107.805 168.280 108.135 169.430 ;
        RECT 108.305 169.300 109.315 169.470 ;
        RECT 108.305 168.450 108.475 169.300 ;
        RECT 108.645 168.280 108.975 169.080 ;
        RECT 109.145 168.450 109.315 169.300 ;
        RECT 109.520 169.430 109.690 169.670 ;
        RECT 109.860 169.600 110.240 169.840 ;
        RECT 110.435 169.560 110.765 169.930 ;
        RECT 111.000 169.855 111.170 170.110 ;
        RECT 111.000 169.525 111.285 169.855 ;
        RECT 109.520 169.260 110.235 169.430 ;
        RECT 111.000 169.380 111.170 169.525 ;
        RECT 109.495 168.280 109.735 169.080 ;
        RECT 109.905 168.450 110.235 169.260 ;
        RECT 110.505 169.210 111.170 169.380 ;
        RECT 111.455 169.355 111.625 170.155 ;
        RECT 110.505 168.450 110.675 169.210 ;
        RECT 110.855 168.280 111.185 169.040 ;
        RECT 111.355 168.450 111.625 169.355 ;
        RECT 113.390 168.715 113.740 169.965 ;
        RECT 115.220 169.455 115.560 170.285 ;
        RECT 117.315 170.080 118.525 170.830 ;
        RECT 117.315 169.370 117.835 169.910 ;
        RECT 118.005 169.540 118.525 170.080 ;
        RECT 111.800 168.280 117.145 168.715 ;
        RECT 117.315 168.280 118.525 169.370 ;
        RECT 11.430 168.110 118.610 168.280 ;
        RECT 11.515 167.020 12.725 168.110 ;
        RECT 11.515 166.310 12.035 166.850 ;
        RECT 12.205 166.480 12.725 167.020 ;
        RECT 13.905 167.180 14.075 167.940 ;
        RECT 14.255 167.350 14.585 168.110 ;
        RECT 13.905 167.010 14.570 167.180 ;
        RECT 14.755 167.035 15.025 167.940 ;
        RECT 14.400 166.865 14.570 167.010 ;
        RECT 13.835 166.460 14.165 166.830 ;
        RECT 14.400 166.535 14.685 166.865 ;
        RECT 11.515 165.560 12.725 166.310 ;
        RECT 14.400 166.280 14.570 166.535 ;
        RECT 13.905 166.110 14.570 166.280 ;
        RECT 14.855 166.235 15.025 167.035 ;
        RECT 15.195 166.945 15.485 168.110 ;
        RECT 15.660 166.920 15.915 167.800 ;
        RECT 16.085 166.970 16.390 168.110 ;
        RECT 16.730 167.730 17.060 168.110 ;
        RECT 17.240 167.560 17.410 167.850 ;
        RECT 17.580 167.650 17.830 168.110 ;
        RECT 16.610 167.390 17.410 167.560 ;
        RECT 18.000 167.600 18.870 167.940 ;
        RECT 13.905 165.730 14.075 166.110 ;
        RECT 14.255 165.560 14.585 165.940 ;
        RECT 14.765 165.730 15.025 166.235 ;
        RECT 15.195 165.560 15.485 166.285 ;
        RECT 15.660 166.270 15.870 166.920 ;
        RECT 16.610 166.800 16.780 167.390 ;
        RECT 18.000 167.220 18.170 167.600 ;
        RECT 19.105 167.480 19.275 167.940 ;
        RECT 19.445 167.650 19.815 168.110 ;
        RECT 20.110 167.510 20.280 167.850 ;
        RECT 20.450 167.680 20.780 168.110 ;
        RECT 21.015 167.510 21.185 167.850 ;
        RECT 16.950 167.050 18.170 167.220 ;
        RECT 18.340 167.140 18.800 167.430 ;
        RECT 19.105 167.310 19.665 167.480 ;
        RECT 20.110 167.340 21.185 167.510 ;
        RECT 21.355 167.610 22.035 167.940 ;
        RECT 22.250 167.610 22.500 167.940 ;
        RECT 22.670 167.650 22.920 168.110 ;
        RECT 19.495 167.170 19.665 167.310 ;
        RECT 18.340 167.130 19.305 167.140 ;
        RECT 18.000 166.960 18.170 167.050 ;
        RECT 18.630 166.970 19.305 167.130 ;
        RECT 16.040 166.770 16.780 166.800 ;
        RECT 16.040 166.470 16.955 166.770 ;
        RECT 16.630 166.295 16.955 166.470 ;
        RECT 15.660 165.740 15.915 166.270 ;
        RECT 16.085 165.560 16.390 166.020 ;
        RECT 16.635 165.940 16.955 166.295 ;
        RECT 17.125 166.510 17.665 166.880 ;
        RECT 18.000 166.790 18.405 166.960 ;
        RECT 17.125 166.110 17.365 166.510 ;
        RECT 17.845 166.340 18.065 166.620 ;
        RECT 17.535 166.170 18.065 166.340 ;
        RECT 17.535 165.940 17.705 166.170 ;
        RECT 18.235 166.010 18.405 166.790 ;
        RECT 18.575 166.180 18.925 166.800 ;
        RECT 19.095 166.180 19.305 166.970 ;
        RECT 19.495 167.000 20.995 167.170 ;
        RECT 19.495 166.310 19.665 167.000 ;
        RECT 21.355 166.830 21.525 167.610 ;
        RECT 22.330 167.480 22.500 167.610 ;
        RECT 19.835 166.660 21.525 166.830 ;
        RECT 21.695 167.050 22.160 167.440 ;
        RECT 22.330 167.310 22.725 167.480 ;
        RECT 19.835 166.480 20.005 166.660 ;
        RECT 16.635 165.770 17.705 165.940 ;
        RECT 17.875 165.560 18.065 166.000 ;
        RECT 18.235 165.730 19.185 166.010 ;
        RECT 19.495 165.920 19.755 166.310 ;
        RECT 20.175 166.240 20.965 166.490 ;
        RECT 19.405 165.750 19.755 165.920 ;
        RECT 19.965 165.560 20.295 166.020 ;
        RECT 21.170 165.950 21.340 166.660 ;
        RECT 21.695 166.460 21.865 167.050 ;
        RECT 21.510 166.240 21.865 166.460 ;
        RECT 22.035 166.240 22.385 166.860 ;
        RECT 22.555 165.950 22.725 167.310 ;
        RECT 23.090 167.140 23.415 167.925 ;
        RECT 22.895 166.090 23.355 167.140 ;
        RECT 21.170 165.780 22.025 165.950 ;
        RECT 22.230 165.780 22.725 165.950 ;
        RECT 22.895 165.560 23.225 165.920 ;
        RECT 23.585 165.820 23.755 167.940 ;
        RECT 23.925 167.610 24.255 168.110 ;
        RECT 24.425 167.440 24.680 167.940 ;
        RECT 23.930 167.270 24.680 167.440 ;
        RECT 25.775 167.350 26.290 167.760 ;
        RECT 26.525 167.350 26.695 168.110 ;
        RECT 26.865 167.770 28.895 167.940 ;
        RECT 23.930 166.280 24.160 167.270 ;
        RECT 24.330 166.450 24.680 167.100 ;
        RECT 25.775 166.540 26.115 167.350 ;
        RECT 26.865 167.105 27.035 167.770 ;
        RECT 27.430 167.430 28.555 167.600 ;
        RECT 26.285 166.915 27.035 167.105 ;
        RECT 27.205 167.090 28.215 167.260 ;
        RECT 25.775 166.370 27.005 166.540 ;
        RECT 23.930 166.110 24.680 166.280 ;
        RECT 23.925 165.560 24.255 165.940 ;
        RECT 24.425 165.820 24.680 166.110 ;
        RECT 26.050 165.765 26.295 166.370 ;
        RECT 26.515 165.560 27.025 166.095 ;
        RECT 27.205 165.730 27.395 167.090 ;
        RECT 27.565 166.750 27.840 166.890 ;
        RECT 27.565 166.580 27.845 166.750 ;
        RECT 27.565 165.730 27.840 166.580 ;
        RECT 28.045 166.290 28.215 167.090 ;
        RECT 28.385 166.300 28.555 167.430 ;
        RECT 28.725 166.800 28.895 167.770 ;
        RECT 29.065 166.970 29.235 168.110 ;
        RECT 29.405 166.970 29.740 167.940 ;
        RECT 28.725 166.470 28.920 166.800 ;
        RECT 29.145 166.470 29.400 166.800 ;
        RECT 29.145 166.300 29.315 166.470 ;
        RECT 29.570 166.300 29.740 166.970 ;
        RECT 29.915 167.350 30.430 167.760 ;
        RECT 30.665 167.350 30.835 168.110 ;
        RECT 31.005 167.770 33.035 167.940 ;
        RECT 29.915 166.540 30.255 167.350 ;
        RECT 31.005 167.105 31.175 167.770 ;
        RECT 31.570 167.430 32.695 167.600 ;
        RECT 30.425 166.915 31.175 167.105 ;
        RECT 31.345 167.090 32.355 167.260 ;
        RECT 29.915 166.370 31.145 166.540 ;
        RECT 28.385 166.130 29.315 166.300 ;
        RECT 28.385 166.095 28.560 166.130 ;
        RECT 28.030 165.730 28.560 166.095 ;
        RECT 28.985 165.560 29.315 165.960 ;
        RECT 29.485 165.730 29.740 166.300 ;
        RECT 30.190 165.765 30.435 166.370 ;
        RECT 30.655 165.560 31.165 166.095 ;
        RECT 31.345 165.730 31.535 167.090 ;
        RECT 31.705 166.410 31.980 166.890 ;
        RECT 31.705 166.240 31.985 166.410 ;
        RECT 32.185 166.290 32.355 167.090 ;
        RECT 32.525 166.300 32.695 167.430 ;
        RECT 32.865 166.800 33.035 167.770 ;
        RECT 33.205 166.970 33.375 168.110 ;
        RECT 33.545 166.970 33.880 167.940 ;
        RECT 32.865 166.470 33.060 166.800 ;
        RECT 33.285 166.470 33.540 166.800 ;
        RECT 33.285 166.300 33.455 166.470 ;
        RECT 33.710 166.300 33.880 166.970 ;
        RECT 31.705 165.730 31.980 166.240 ;
        RECT 32.525 166.130 33.455 166.300 ;
        RECT 32.525 166.095 32.700 166.130 ;
        RECT 32.170 165.730 32.700 166.095 ;
        RECT 33.125 165.560 33.455 165.960 ;
        RECT 33.625 165.730 33.880 166.300 ;
        RECT 34.055 167.035 34.325 167.940 ;
        RECT 34.495 167.350 34.825 168.110 ;
        RECT 35.005 167.180 35.175 167.940 ;
        RECT 35.440 167.675 40.785 168.110 ;
        RECT 34.055 166.235 34.225 167.035 ;
        RECT 34.510 167.010 35.175 167.180 ;
        RECT 34.510 166.865 34.680 167.010 ;
        RECT 34.395 166.535 34.680 166.865 ;
        RECT 34.510 166.280 34.680 166.535 ;
        RECT 34.915 166.460 35.245 166.830 ;
        RECT 37.030 166.425 37.380 167.675 ;
        RECT 40.955 166.945 41.245 168.110 ;
        RECT 41.415 167.020 44.925 168.110 ;
        RECT 34.055 165.730 34.315 166.235 ;
        RECT 34.510 166.110 35.175 166.280 ;
        RECT 34.495 165.560 34.825 165.940 ;
        RECT 35.005 165.730 35.175 166.110 ;
        RECT 38.860 166.105 39.200 166.935 ;
        RECT 41.415 166.500 43.105 167.020 ;
        RECT 45.245 166.960 45.575 168.110 ;
        RECT 45.745 167.090 45.915 167.940 ;
        RECT 46.085 167.310 46.415 168.110 ;
        RECT 46.585 167.090 46.755 167.940 ;
        RECT 46.935 167.310 47.175 168.110 ;
        RECT 47.345 167.130 47.675 167.940 ;
        RECT 45.745 166.920 46.755 167.090 ;
        RECT 46.960 166.960 47.675 167.130 ;
        RECT 47.855 167.020 49.065 168.110 ;
        RECT 43.275 166.330 44.925 166.850 ;
        RECT 45.745 166.410 46.240 166.920 ;
        RECT 46.960 166.720 47.130 166.960 ;
        RECT 46.630 166.550 47.130 166.720 ;
        RECT 47.300 166.550 47.680 166.790 ;
        RECT 45.745 166.380 46.245 166.410 ;
        RECT 46.960 166.380 47.130 166.550 ;
        RECT 47.855 166.480 48.375 167.020 ;
        RECT 49.240 166.970 49.575 167.940 ;
        RECT 49.745 166.970 49.915 168.110 ;
        RECT 50.085 167.770 52.115 167.940 ;
        RECT 35.440 165.560 40.785 166.105 ;
        RECT 40.955 165.560 41.245 166.285 ;
        RECT 41.415 165.560 44.925 166.330 ;
        RECT 45.245 165.560 45.575 166.360 ;
        RECT 45.745 166.210 46.755 166.380 ;
        RECT 46.960 166.210 47.595 166.380 ;
        RECT 48.545 166.310 49.065 166.850 ;
        RECT 45.745 165.730 45.915 166.210 ;
        RECT 46.085 165.560 46.415 166.040 ;
        RECT 46.585 165.730 46.755 166.210 ;
        RECT 47.005 165.560 47.245 166.040 ;
        RECT 47.425 165.730 47.595 166.210 ;
        RECT 47.855 165.560 49.065 166.310 ;
        RECT 49.240 166.300 49.410 166.970 ;
        RECT 50.085 166.800 50.255 167.770 ;
        RECT 49.580 166.470 49.835 166.800 ;
        RECT 50.060 166.470 50.255 166.800 ;
        RECT 50.425 167.430 51.550 167.600 ;
        RECT 49.665 166.300 49.835 166.470 ;
        RECT 50.425 166.300 50.595 167.430 ;
        RECT 49.240 165.730 49.495 166.300 ;
        RECT 49.665 166.130 50.595 166.300 ;
        RECT 50.765 167.090 51.775 167.260 ;
        RECT 50.765 166.290 50.935 167.090 ;
        RECT 51.140 166.750 51.415 166.890 ;
        RECT 51.135 166.580 51.415 166.750 ;
        RECT 50.420 166.095 50.595 166.130 ;
        RECT 49.665 165.560 49.995 165.960 ;
        RECT 50.420 165.730 50.950 166.095 ;
        RECT 51.140 165.730 51.415 166.580 ;
        RECT 51.585 165.730 51.775 167.090 ;
        RECT 51.945 167.105 52.115 167.770 ;
        RECT 52.285 167.350 52.455 168.110 ;
        RECT 52.690 167.350 53.205 167.760 ;
        RECT 51.945 166.915 52.695 167.105 ;
        RECT 52.865 166.540 53.205 167.350 ;
        RECT 53.750 167.130 54.005 167.800 ;
        RECT 54.185 167.310 54.470 168.110 ;
        RECT 54.650 167.390 54.980 167.900 ;
        RECT 53.750 166.750 53.930 167.130 ;
        RECT 54.650 166.800 54.900 167.390 ;
        RECT 55.250 167.240 55.420 167.850 ;
        RECT 55.590 167.420 55.920 168.110 ;
        RECT 56.150 167.560 56.390 167.850 ;
        RECT 56.590 167.730 57.010 168.110 ;
        RECT 57.190 167.640 57.820 167.890 ;
        RECT 58.290 167.730 58.620 168.110 ;
        RECT 57.190 167.560 57.360 167.640 ;
        RECT 58.790 167.560 58.960 167.850 ;
        RECT 59.140 167.730 59.520 168.110 ;
        RECT 59.760 167.725 60.590 167.895 ;
        RECT 56.150 167.390 57.360 167.560 ;
        RECT 53.665 166.580 53.930 166.750 ;
        RECT 51.975 166.370 53.205 166.540 ;
        RECT 51.955 165.560 52.465 166.095 ;
        RECT 52.685 165.765 52.930 166.370 ;
        RECT 53.750 166.270 53.930 166.580 ;
        RECT 54.100 166.470 54.900 166.800 ;
        RECT 53.750 165.740 54.005 166.270 ;
        RECT 54.185 165.560 54.470 166.020 ;
        RECT 54.650 165.820 54.900 166.470 ;
        RECT 55.100 167.220 55.420 167.240 ;
        RECT 55.100 167.050 57.020 167.220 ;
        RECT 55.100 166.155 55.290 167.050 ;
        RECT 57.190 166.880 57.360 167.390 ;
        RECT 57.530 167.130 58.050 167.440 ;
        RECT 55.460 166.710 57.360 166.880 ;
        RECT 55.460 166.650 55.790 166.710 ;
        RECT 55.940 166.480 56.270 166.540 ;
        RECT 55.610 166.210 56.270 166.480 ;
        RECT 55.100 165.825 55.420 166.155 ;
        RECT 55.600 165.560 56.260 166.040 ;
        RECT 56.460 165.950 56.630 166.710 ;
        RECT 57.530 166.540 57.710 166.950 ;
        RECT 56.800 166.370 57.130 166.490 ;
        RECT 57.880 166.370 58.050 167.130 ;
        RECT 56.800 166.200 58.050 166.370 ;
        RECT 58.220 167.310 59.590 167.560 ;
        RECT 58.220 166.540 58.410 167.310 ;
        RECT 59.340 167.050 59.590 167.310 ;
        RECT 58.580 166.880 58.830 167.040 ;
        RECT 59.760 166.880 59.930 167.725 ;
        RECT 60.825 167.440 60.995 167.940 ;
        RECT 61.165 167.610 61.495 168.110 ;
        RECT 60.100 167.050 60.600 167.430 ;
        RECT 60.825 167.270 61.520 167.440 ;
        RECT 58.580 166.710 59.930 166.880 ;
        RECT 59.510 166.670 59.930 166.710 ;
        RECT 58.220 166.200 58.640 166.540 ;
        RECT 58.930 166.210 59.340 166.540 ;
        RECT 56.460 165.780 57.310 165.950 ;
        RECT 57.870 165.560 58.190 166.020 ;
        RECT 58.390 165.770 58.640 166.200 ;
        RECT 58.930 165.560 59.340 166.000 ;
        RECT 59.510 165.940 59.680 166.670 ;
        RECT 59.850 166.120 60.200 166.490 ;
        RECT 60.380 166.180 60.600 167.050 ;
        RECT 60.770 166.480 61.180 167.100 ;
        RECT 61.350 166.300 61.520 167.270 ;
        RECT 60.825 166.110 61.520 166.300 ;
        RECT 59.510 165.740 60.525 165.940 ;
        RECT 60.825 165.780 60.995 166.110 ;
        RECT 61.165 165.560 61.495 165.940 ;
        RECT 61.710 165.820 61.935 167.940 ;
        RECT 62.105 167.610 62.435 168.110 ;
        RECT 62.605 167.440 62.775 167.940 ;
        RECT 62.110 167.270 62.775 167.440 ;
        RECT 62.110 166.280 62.340 167.270 ;
        RECT 64.045 167.180 64.215 167.940 ;
        RECT 64.430 167.350 64.760 168.110 ;
        RECT 62.510 166.450 62.860 167.100 ;
        RECT 64.045 167.010 64.760 167.180 ;
        RECT 64.930 167.035 65.185 167.940 ;
        RECT 63.955 166.460 64.310 166.830 ;
        RECT 64.590 166.800 64.760 167.010 ;
        RECT 64.590 166.470 64.845 166.800 ;
        RECT 64.590 166.280 64.760 166.470 ;
        RECT 65.015 166.305 65.185 167.035 ;
        RECT 65.360 166.960 65.620 168.110 ;
        RECT 66.715 166.945 67.005 168.110 ;
        RECT 67.265 167.180 67.435 167.940 ;
        RECT 67.650 167.350 67.980 168.110 ;
        RECT 67.265 167.010 67.980 167.180 ;
        RECT 68.150 167.035 68.405 167.940 ;
        RECT 67.175 166.460 67.530 166.830 ;
        RECT 67.810 166.800 67.980 167.010 ;
        RECT 67.810 166.470 68.065 166.800 ;
        RECT 62.110 166.110 62.775 166.280 ;
        RECT 62.105 165.560 62.435 165.940 ;
        RECT 62.605 165.820 62.775 166.110 ;
        RECT 64.045 166.110 64.760 166.280 ;
        RECT 64.045 165.730 64.215 166.110 ;
        RECT 64.430 165.560 64.760 165.940 ;
        RECT 64.930 165.730 65.185 166.305 ;
        RECT 65.360 165.560 65.620 166.400 ;
        RECT 66.715 165.560 67.005 166.285 ;
        RECT 67.810 166.280 67.980 166.470 ;
        RECT 68.235 166.305 68.405 167.035 ;
        RECT 68.580 166.960 68.840 168.110 ;
        RECT 69.105 167.180 69.275 167.940 ;
        RECT 69.490 167.350 69.820 168.110 ;
        RECT 69.105 167.010 69.820 167.180 ;
        RECT 69.990 167.035 70.245 167.940 ;
        RECT 69.015 166.460 69.370 166.830 ;
        RECT 69.650 166.800 69.820 167.010 ;
        RECT 69.650 166.470 69.905 166.800 ;
        RECT 67.265 166.110 67.980 166.280 ;
        RECT 67.265 165.730 67.435 166.110 ;
        RECT 67.650 165.560 67.980 165.940 ;
        RECT 68.150 165.730 68.405 166.305 ;
        RECT 68.580 165.560 68.840 166.400 ;
        RECT 69.650 166.280 69.820 166.470 ;
        RECT 70.075 166.305 70.245 167.035 ;
        RECT 70.420 166.960 70.680 168.110 ;
        RECT 71.320 167.675 76.665 168.110 ;
        RECT 77.210 167.770 77.465 167.800 ;
        RECT 72.910 166.425 73.260 167.675 ;
        RECT 77.125 167.600 77.465 167.770 ;
        RECT 77.210 167.130 77.465 167.600 ;
        RECT 77.645 167.310 77.930 168.110 ;
        RECT 78.110 167.390 78.440 167.900 ;
        RECT 69.105 166.110 69.820 166.280 ;
        RECT 69.105 165.730 69.275 166.110 ;
        RECT 69.490 165.560 69.820 165.940 ;
        RECT 69.990 165.730 70.245 166.305 ;
        RECT 70.420 165.560 70.680 166.400 ;
        RECT 74.740 166.105 75.080 166.935 ;
        RECT 77.210 166.270 77.390 167.130 ;
        RECT 78.110 166.800 78.360 167.390 ;
        RECT 78.710 167.240 78.880 167.850 ;
        RECT 79.050 167.420 79.380 168.110 ;
        RECT 79.610 167.560 79.850 167.850 ;
        RECT 80.050 167.730 80.470 168.110 ;
        RECT 80.650 167.640 81.280 167.890 ;
        RECT 81.750 167.730 82.080 168.110 ;
        RECT 80.650 167.560 80.820 167.640 ;
        RECT 82.250 167.560 82.420 167.850 ;
        RECT 82.600 167.730 82.980 168.110 ;
        RECT 83.220 167.725 84.050 167.895 ;
        RECT 79.610 167.390 80.820 167.560 ;
        RECT 77.560 166.470 78.360 166.800 ;
        RECT 71.320 165.560 76.665 166.105 ;
        RECT 77.210 165.740 77.465 166.270 ;
        RECT 77.645 165.560 77.930 166.020 ;
        RECT 78.110 165.820 78.360 166.470 ;
        RECT 78.560 167.220 78.880 167.240 ;
        RECT 78.560 167.050 80.480 167.220 ;
        RECT 78.560 166.155 78.750 167.050 ;
        RECT 80.650 166.880 80.820 167.390 ;
        RECT 80.990 167.130 81.510 167.440 ;
        RECT 78.920 166.710 80.820 166.880 ;
        RECT 78.920 166.650 79.250 166.710 ;
        RECT 79.400 166.480 79.730 166.540 ;
        RECT 79.070 166.210 79.730 166.480 ;
        RECT 78.560 165.825 78.880 166.155 ;
        RECT 79.060 165.560 79.720 166.040 ;
        RECT 79.920 165.950 80.090 166.710 ;
        RECT 80.990 166.540 81.170 166.950 ;
        RECT 80.260 166.370 80.590 166.490 ;
        RECT 81.340 166.370 81.510 167.130 ;
        RECT 80.260 166.200 81.510 166.370 ;
        RECT 81.680 167.310 83.050 167.560 ;
        RECT 81.680 166.540 81.870 167.310 ;
        RECT 82.800 167.050 83.050 167.310 ;
        RECT 82.040 166.880 82.290 167.040 ;
        RECT 83.220 166.880 83.390 167.725 ;
        RECT 84.285 167.440 84.455 167.940 ;
        RECT 84.625 167.610 84.955 168.110 ;
        RECT 83.560 167.050 84.060 167.430 ;
        RECT 84.285 167.270 84.980 167.440 ;
        RECT 82.040 166.710 83.390 166.880 ;
        RECT 82.970 166.670 83.390 166.710 ;
        RECT 81.680 166.200 82.100 166.540 ;
        RECT 82.390 166.210 82.800 166.540 ;
        RECT 79.920 165.780 80.770 165.950 ;
        RECT 81.330 165.560 81.650 166.020 ;
        RECT 81.850 165.770 82.100 166.200 ;
        RECT 82.390 165.560 82.800 166.000 ;
        RECT 82.970 165.940 83.140 166.670 ;
        RECT 83.310 166.120 83.660 166.490 ;
        RECT 83.840 166.180 84.060 167.050 ;
        RECT 84.230 166.480 84.640 167.100 ;
        RECT 84.810 166.300 84.980 167.270 ;
        RECT 84.285 166.110 84.980 166.300 ;
        RECT 82.970 165.740 83.985 165.940 ;
        RECT 84.285 165.780 84.455 166.110 ;
        RECT 84.625 165.560 84.955 165.940 ;
        RECT 85.170 165.820 85.395 167.940 ;
        RECT 85.565 167.610 85.895 168.110 ;
        RECT 86.065 167.440 86.235 167.940 ;
        RECT 86.960 167.675 92.305 168.110 ;
        RECT 85.570 167.270 86.235 167.440 ;
        RECT 85.570 166.280 85.800 167.270 ;
        RECT 85.970 166.450 86.320 167.100 ;
        RECT 88.550 166.425 88.900 167.675 ;
        RECT 92.475 166.945 92.765 168.110 ;
        RECT 94.060 167.140 94.390 167.940 ;
        RECT 94.560 167.310 94.890 168.110 ;
        RECT 95.190 167.140 95.520 167.940 ;
        RECT 96.165 167.310 96.415 168.110 ;
        RECT 94.060 166.970 96.495 167.140 ;
        RECT 96.685 166.970 96.855 168.110 ;
        RECT 97.025 166.970 97.365 167.940 ;
        RECT 85.570 166.110 86.235 166.280 ;
        RECT 85.565 165.560 85.895 165.940 ;
        RECT 86.065 165.820 86.235 166.110 ;
        RECT 90.380 166.105 90.720 166.935 ;
        RECT 93.855 166.550 94.205 166.800 ;
        RECT 94.390 166.340 94.560 166.970 ;
        RECT 94.730 166.550 95.060 166.750 ;
        RECT 95.230 166.550 95.560 166.750 ;
        RECT 95.730 166.550 96.150 166.750 ;
        RECT 96.325 166.720 96.495 166.970 ;
        RECT 96.325 166.550 97.020 166.720 ;
        RECT 86.960 165.560 92.305 166.105 ;
        RECT 92.475 165.560 92.765 166.285 ;
        RECT 94.060 165.730 94.560 166.340 ;
        RECT 95.190 166.210 96.415 166.380 ;
        RECT 97.190 166.360 97.365 166.970 ;
        RECT 97.995 167.020 100.585 168.110 ;
        RECT 100.760 167.675 106.105 168.110 ;
        RECT 106.280 167.675 111.625 168.110 ;
        RECT 111.800 167.675 117.145 168.110 ;
        RECT 97.995 166.500 99.205 167.020 ;
        RECT 95.190 165.730 95.520 166.210 ;
        RECT 95.690 165.560 95.915 166.020 ;
        RECT 96.085 165.730 96.415 166.210 ;
        RECT 96.605 165.560 96.855 166.360 ;
        RECT 97.025 165.730 97.365 166.360 ;
        RECT 99.375 166.330 100.585 166.850 ;
        RECT 102.350 166.425 102.700 167.675 ;
        RECT 97.995 165.560 100.585 166.330 ;
        RECT 104.180 166.105 104.520 166.935 ;
        RECT 107.870 166.425 108.220 167.675 ;
        RECT 109.700 166.105 110.040 166.935 ;
        RECT 113.390 166.425 113.740 167.675 ;
        RECT 117.315 167.020 118.525 168.110 ;
        RECT 115.220 166.105 115.560 166.935 ;
        RECT 117.315 166.480 117.835 167.020 ;
        RECT 118.005 166.310 118.525 166.850 ;
        RECT 100.760 165.560 106.105 166.105 ;
        RECT 106.280 165.560 111.625 166.105 ;
        RECT 111.800 165.560 117.145 166.105 ;
        RECT 117.315 165.560 118.525 166.310 ;
        RECT 11.430 165.390 118.610 165.560 ;
        RECT 11.515 164.640 12.725 165.390 ;
        RECT 11.515 164.100 12.035 164.640 ;
        RECT 12.895 164.620 15.485 165.390 ;
        RECT 12.205 163.930 12.725 164.470 ;
        RECT 11.515 162.840 12.725 163.930 ;
        RECT 12.895 163.930 14.105 164.450 ;
        RECT 14.275 164.100 15.485 164.620 ;
        RECT 15.695 164.570 15.925 165.390 ;
        RECT 16.095 164.590 16.425 165.220 ;
        RECT 15.675 164.150 16.005 164.400 ;
        RECT 16.175 163.990 16.425 164.590 ;
        RECT 16.595 164.570 16.805 165.390 ;
        RECT 17.125 164.840 17.295 165.220 ;
        RECT 17.475 165.010 17.805 165.390 ;
        RECT 17.125 164.670 17.790 164.840 ;
        RECT 17.985 164.715 18.245 165.220 ;
        RECT 17.055 164.120 17.385 164.490 ;
        RECT 17.620 164.415 17.790 164.670 ;
        RECT 12.895 162.840 15.485 163.930 ;
        RECT 15.695 162.840 15.925 163.980 ;
        RECT 16.095 163.010 16.425 163.990 ;
        RECT 17.620 164.085 17.905 164.415 ;
        RECT 16.595 162.840 16.805 163.980 ;
        RECT 17.620 163.940 17.790 164.085 ;
        RECT 17.125 163.770 17.790 163.940 ;
        RECT 18.075 163.915 18.245 164.715 ;
        RECT 17.125 163.010 17.295 163.770 ;
        RECT 17.475 162.840 17.805 163.600 ;
        RECT 17.975 163.010 18.245 163.915 ;
        RECT 18.420 164.650 18.675 165.220 ;
        RECT 18.845 164.990 19.175 165.390 ;
        RECT 19.600 164.855 20.130 165.220 ;
        RECT 19.600 164.820 19.775 164.855 ;
        RECT 18.845 164.650 19.775 164.820 ;
        RECT 18.420 163.980 18.590 164.650 ;
        RECT 18.845 164.480 19.015 164.650 ;
        RECT 18.760 164.150 19.015 164.480 ;
        RECT 19.240 164.150 19.435 164.480 ;
        RECT 18.420 163.010 18.755 163.980 ;
        RECT 18.925 162.840 19.095 163.980 ;
        RECT 19.265 163.180 19.435 164.150 ;
        RECT 19.605 163.520 19.775 164.650 ;
        RECT 19.945 163.860 20.115 164.660 ;
        RECT 20.320 164.370 20.595 165.220 ;
        RECT 20.315 164.200 20.595 164.370 ;
        RECT 20.320 164.060 20.595 164.200 ;
        RECT 20.765 163.860 20.955 165.220 ;
        RECT 21.135 164.855 21.645 165.390 ;
        RECT 21.865 164.580 22.110 165.185 ;
        RECT 22.560 164.845 27.905 165.390 ;
        RECT 21.155 164.410 22.385 164.580 ;
        RECT 19.945 163.690 20.955 163.860 ;
        RECT 21.125 163.845 21.875 164.035 ;
        RECT 19.605 163.350 20.730 163.520 ;
        RECT 21.125 163.180 21.295 163.845 ;
        RECT 22.045 163.600 22.385 164.410 ;
        RECT 19.265 163.010 21.295 163.180 ;
        RECT 21.465 162.840 21.635 163.600 ;
        RECT 21.870 163.190 22.385 163.600 ;
        RECT 24.150 163.275 24.500 164.525 ;
        RECT 25.980 164.015 26.320 164.845 ;
        RECT 28.075 164.665 28.365 165.390 ;
        RECT 28.625 164.840 28.795 165.130 ;
        RECT 28.965 165.010 29.295 165.390 ;
        RECT 28.625 164.670 29.290 164.840 ;
        RECT 22.560 162.840 27.905 163.275 ;
        RECT 28.075 162.840 28.365 164.005 ;
        RECT 28.540 163.850 28.890 164.500 ;
        RECT 29.060 163.680 29.290 164.670 ;
        RECT 28.625 163.510 29.290 163.680 ;
        RECT 28.625 163.010 28.795 163.510 ;
        RECT 28.965 162.840 29.295 163.340 ;
        RECT 29.465 163.010 29.690 165.130 ;
        RECT 29.905 165.010 30.235 165.390 ;
        RECT 30.405 164.840 30.575 165.170 ;
        RECT 30.875 165.010 31.890 165.210 ;
        RECT 29.880 164.650 30.575 164.840 ;
        RECT 29.880 163.680 30.050 164.650 ;
        RECT 30.220 163.850 30.630 164.470 ;
        RECT 30.800 163.900 31.020 164.770 ;
        RECT 31.200 164.460 31.550 164.830 ;
        RECT 31.720 164.280 31.890 165.010 ;
        RECT 32.060 164.950 32.470 165.390 ;
        RECT 32.760 164.750 33.010 165.180 ;
        RECT 33.210 164.930 33.530 165.390 ;
        RECT 34.090 165.000 34.940 165.170 ;
        RECT 32.060 164.410 32.470 164.740 ;
        RECT 32.760 164.410 33.180 164.750 ;
        RECT 31.470 164.240 31.890 164.280 ;
        RECT 31.470 164.070 32.820 164.240 ;
        RECT 29.880 163.510 30.575 163.680 ;
        RECT 30.800 163.520 31.300 163.900 ;
        RECT 29.905 162.840 30.235 163.340 ;
        RECT 30.405 163.010 30.575 163.510 ;
        RECT 31.470 163.225 31.640 164.070 ;
        RECT 32.570 163.910 32.820 164.070 ;
        RECT 31.810 163.640 32.060 163.900 ;
        RECT 32.990 163.640 33.180 164.410 ;
        RECT 31.810 163.390 33.180 163.640 ;
        RECT 33.350 164.580 34.600 164.750 ;
        RECT 33.350 163.820 33.520 164.580 ;
        RECT 34.270 164.460 34.600 164.580 ;
        RECT 33.690 164.000 33.870 164.410 ;
        RECT 34.770 164.240 34.940 165.000 ;
        RECT 35.140 164.910 35.800 165.390 ;
        RECT 35.980 164.795 36.300 165.125 ;
        RECT 35.130 164.470 35.790 164.740 ;
        RECT 35.130 164.410 35.460 164.470 ;
        RECT 35.610 164.240 35.940 164.300 ;
        RECT 34.040 164.070 35.940 164.240 ;
        RECT 33.350 163.510 33.870 163.820 ;
        RECT 34.040 163.560 34.210 164.070 ;
        RECT 36.110 163.900 36.300 164.795 ;
        RECT 34.380 163.730 36.300 163.900 ;
        RECT 35.980 163.710 36.300 163.730 ;
        RECT 36.500 164.480 36.750 165.130 ;
        RECT 36.930 164.930 37.215 165.390 ;
        RECT 37.395 164.680 37.650 165.210 ;
        RECT 36.500 164.150 37.300 164.480 ;
        RECT 34.040 163.390 35.250 163.560 ;
        RECT 30.810 163.055 31.640 163.225 ;
        RECT 31.880 162.840 32.260 163.220 ;
        RECT 32.440 163.100 32.610 163.390 ;
        RECT 34.040 163.310 34.210 163.390 ;
        RECT 32.780 162.840 33.110 163.220 ;
        RECT 33.580 163.060 34.210 163.310 ;
        RECT 34.390 162.840 34.810 163.220 ;
        RECT 35.010 163.100 35.250 163.390 ;
        RECT 35.480 162.840 35.810 163.530 ;
        RECT 35.980 163.100 36.150 163.710 ;
        RECT 36.500 163.560 36.750 164.150 ;
        RECT 37.470 164.030 37.650 164.680 ;
        RECT 38.195 164.620 39.865 165.390 ;
        RECT 37.470 163.860 37.735 164.030 ;
        RECT 38.195 163.930 38.945 164.450 ;
        RECT 39.115 164.100 39.865 164.620 ;
        RECT 40.240 164.610 40.740 165.220 ;
        RECT 40.035 164.150 40.385 164.400 ;
        RECT 40.570 163.980 40.740 164.610 ;
        RECT 41.370 164.740 41.700 165.220 ;
        RECT 41.870 164.930 42.095 165.390 ;
        RECT 42.265 164.740 42.595 165.220 ;
        RECT 41.370 164.570 42.595 164.740 ;
        RECT 42.785 164.590 43.035 165.390 ;
        RECT 43.205 164.590 43.545 165.220 ;
        RECT 43.920 164.610 44.420 165.220 ;
        RECT 40.910 164.200 41.240 164.400 ;
        RECT 41.410 164.200 41.740 164.400 ;
        RECT 41.910 164.200 42.330 164.400 ;
        RECT 42.505 164.230 43.200 164.400 ;
        RECT 42.505 163.980 42.675 164.230 ;
        RECT 43.370 163.980 43.545 164.590 ;
        RECT 43.715 164.150 44.065 164.400 ;
        RECT 44.250 163.980 44.420 164.610 ;
        RECT 45.050 164.740 45.380 165.220 ;
        RECT 45.550 164.930 45.775 165.390 ;
        RECT 45.945 164.740 46.275 165.220 ;
        RECT 45.050 164.570 46.275 164.740 ;
        RECT 46.465 164.590 46.715 165.390 ;
        RECT 46.885 164.590 47.225 165.220 ;
        RECT 44.590 164.200 44.920 164.400 ;
        RECT 45.090 164.200 45.420 164.400 ;
        RECT 45.590 164.200 46.010 164.400 ;
        RECT 46.185 164.230 46.880 164.400 ;
        RECT 46.185 163.980 46.355 164.230 ;
        RECT 47.050 163.980 47.225 164.590 ;
        RECT 37.470 163.820 37.650 163.860 ;
        RECT 36.420 163.050 36.750 163.560 ;
        RECT 36.930 162.840 37.215 163.640 ;
        RECT 37.395 163.150 37.650 163.820 ;
        RECT 38.195 162.840 39.865 163.930 ;
        RECT 40.240 163.810 42.675 163.980 ;
        RECT 40.240 163.010 40.570 163.810 ;
        RECT 40.740 162.840 41.070 163.640 ;
        RECT 41.370 163.010 41.700 163.810 ;
        RECT 42.345 162.840 42.595 163.640 ;
        RECT 42.865 162.840 43.035 163.980 ;
        RECT 43.205 163.010 43.545 163.980 ;
        RECT 43.920 163.810 46.355 163.980 ;
        RECT 43.920 163.010 44.250 163.810 ;
        RECT 44.420 162.840 44.750 163.640 ;
        RECT 45.050 163.010 45.380 163.810 ;
        RECT 46.025 162.840 46.275 163.640 ;
        RECT 46.545 162.840 46.715 163.980 ;
        RECT 46.885 163.010 47.225 163.980 ;
        RECT 47.395 164.715 47.655 165.220 ;
        RECT 47.835 165.010 48.165 165.390 ;
        RECT 48.345 164.840 48.515 165.220 ;
        RECT 47.395 163.915 47.565 164.715 ;
        RECT 47.850 164.670 48.515 164.840 ;
        RECT 47.850 164.415 48.020 164.670 ;
        RECT 48.775 164.650 49.160 165.220 ;
        RECT 49.330 164.930 49.655 165.390 ;
        RECT 50.175 164.760 50.455 165.220 ;
        RECT 47.735 164.085 48.020 164.415 ;
        RECT 48.255 164.120 48.585 164.490 ;
        RECT 47.850 163.940 48.020 164.085 ;
        RECT 48.775 163.980 49.055 164.650 ;
        RECT 49.330 164.590 50.455 164.760 ;
        RECT 49.330 164.480 49.780 164.590 ;
        RECT 49.225 164.150 49.780 164.480 ;
        RECT 50.645 164.420 51.045 165.220 ;
        RECT 51.445 164.930 51.715 165.390 ;
        RECT 51.885 164.760 52.170 165.220 ;
        RECT 47.395 163.010 47.665 163.915 ;
        RECT 47.850 163.770 48.515 163.940 ;
        RECT 47.835 162.840 48.165 163.600 ;
        RECT 48.345 163.010 48.515 163.770 ;
        RECT 48.775 163.010 49.160 163.980 ;
        RECT 49.330 163.690 49.780 164.150 ;
        RECT 49.950 163.860 51.045 164.420 ;
        RECT 49.330 163.470 50.455 163.690 ;
        RECT 49.330 162.840 49.655 163.300 ;
        RECT 50.175 163.010 50.455 163.470 ;
        RECT 50.645 163.010 51.045 163.860 ;
        RECT 51.215 164.590 52.170 164.760 ;
        RECT 52.455 164.640 53.665 165.390 ;
        RECT 53.835 164.665 54.125 165.390 ;
        RECT 51.215 163.690 51.425 164.590 ;
        RECT 51.595 163.860 52.285 164.420 ;
        RECT 52.455 163.930 52.975 164.470 ;
        RECT 53.145 164.100 53.665 164.640 ;
        RECT 54.755 164.590 55.095 165.220 ;
        RECT 55.265 164.590 55.515 165.390 ;
        RECT 55.705 164.740 56.035 165.220 ;
        RECT 56.205 164.930 56.430 165.390 ;
        RECT 56.600 164.740 56.930 165.220 ;
        RECT 51.215 163.470 52.170 163.690 ;
        RECT 51.445 162.840 51.715 163.300 ;
        RECT 51.885 163.010 52.170 163.470 ;
        RECT 52.455 162.840 53.665 163.930 ;
        RECT 53.835 162.840 54.125 164.005 ;
        RECT 54.755 163.980 54.930 164.590 ;
        RECT 55.705 164.570 56.930 164.740 ;
        RECT 57.560 164.610 58.060 165.220 ;
        RECT 55.100 164.230 55.795 164.400 ;
        RECT 55.625 163.980 55.795 164.230 ;
        RECT 55.970 164.200 56.390 164.400 ;
        RECT 56.560 164.200 56.890 164.400 ;
        RECT 57.060 164.200 57.390 164.400 ;
        RECT 57.560 163.980 57.730 164.610 ;
        RECT 58.710 164.580 58.955 165.185 ;
        RECT 59.175 164.855 59.685 165.390 ;
        RECT 58.435 164.410 59.665 164.580 ;
        RECT 57.915 164.150 58.265 164.400 ;
        RECT 54.755 163.010 55.095 163.980 ;
        RECT 55.265 162.840 55.435 163.980 ;
        RECT 55.625 163.810 58.060 163.980 ;
        RECT 55.705 162.840 55.955 163.640 ;
        RECT 56.600 163.010 56.930 163.810 ;
        RECT 57.230 162.840 57.560 163.640 ;
        RECT 57.730 163.010 58.060 163.810 ;
        RECT 58.435 163.600 58.775 164.410 ;
        RECT 58.945 163.845 59.695 164.035 ;
        RECT 58.435 163.190 58.950 163.600 ;
        RECT 59.185 162.840 59.355 163.600 ;
        RECT 59.525 163.180 59.695 163.845 ;
        RECT 59.865 163.860 60.055 165.220 ;
        RECT 60.225 165.050 60.500 165.220 ;
        RECT 60.225 164.880 60.505 165.050 ;
        RECT 60.225 164.060 60.500 164.880 ;
        RECT 60.690 164.855 61.220 165.220 ;
        RECT 61.645 164.990 61.975 165.390 ;
        RECT 61.045 164.820 61.220 164.855 ;
        RECT 60.705 163.860 60.875 164.660 ;
        RECT 59.865 163.690 60.875 163.860 ;
        RECT 61.045 164.650 61.975 164.820 ;
        RECT 62.145 164.650 62.400 165.220 ;
        RECT 62.950 164.710 63.205 165.210 ;
        RECT 63.385 164.930 63.670 165.390 ;
        RECT 61.045 163.520 61.215 164.650 ;
        RECT 61.805 164.480 61.975 164.650 ;
        RECT 60.090 163.350 61.215 163.520 ;
        RECT 61.385 164.150 61.580 164.480 ;
        RECT 61.805 164.150 62.060 164.480 ;
        RECT 61.385 163.180 61.555 164.150 ;
        RECT 62.230 163.980 62.400 164.650 ;
        RECT 62.865 164.680 63.205 164.710 ;
        RECT 62.865 164.540 63.130 164.680 ;
        RECT 59.525 163.010 61.555 163.180 ;
        RECT 61.725 162.840 61.895 163.980 ;
        RECT 62.065 163.010 62.400 163.980 ;
        RECT 62.950 163.820 63.130 164.540 ;
        RECT 63.850 164.480 64.100 165.130 ;
        RECT 63.300 164.150 64.100 164.480 ;
        RECT 62.950 163.150 63.205 163.820 ;
        RECT 63.385 162.840 63.670 163.640 ;
        RECT 63.850 163.560 64.100 164.150 ;
        RECT 64.300 164.795 64.620 165.125 ;
        RECT 64.800 164.910 65.460 165.390 ;
        RECT 65.660 165.000 66.510 165.170 ;
        RECT 64.300 163.900 64.490 164.795 ;
        RECT 64.810 164.470 65.470 164.740 ;
        RECT 65.140 164.410 65.470 164.470 ;
        RECT 64.660 164.240 64.990 164.300 ;
        RECT 65.660 164.240 65.830 165.000 ;
        RECT 67.070 164.930 67.390 165.390 ;
        RECT 67.590 164.750 67.840 165.180 ;
        RECT 68.130 164.950 68.540 165.390 ;
        RECT 68.710 165.010 69.725 165.210 ;
        RECT 66.000 164.580 67.250 164.750 ;
        RECT 66.000 164.460 66.330 164.580 ;
        RECT 64.660 164.070 66.560 164.240 ;
        RECT 64.300 163.730 66.220 163.900 ;
        RECT 64.300 163.710 64.620 163.730 ;
        RECT 63.850 163.050 64.180 163.560 ;
        RECT 64.450 163.100 64.620 163.710 ;
        RECT 66.390 163.560 66.560 164.070 ;
        RECT 66.730 164.000 66.910 164.410 ;
        RECT 67.080 163.820 67.250 164.580 ;
        RECT 64.790 162.840 65.120 163.530 ;
        RECT 65.350 163.390 66.560 163.560 ;
        RECT 66.730 163.510 67.250 163.820 ;
        RECT 67.420 164.410 67.840 164.750 ;
        RECT 68.130 164.410 68.540 164.740 ;
        RECT 67.420 163.640 67.610 164.410 ;
        RECT 68.710 164.280 68.880 165.010 ;
        RECT 70.025 164.840 70.195 165.170 ;
        RECT 70.365 165.010 70.695 165.390 ;
        RECT 69.050 164.460 69.400 164.830 ;
        RECT 68.710 164.240 69.130 164.280 ;
        RECT 67.780 164.070 69.130 164.240 ;
        RECT 67.780 163.910 68.030 164.070 ;
        RECT 68.540 163.640 68.790 163.900 ;
        RECT 67.420 163.390 68.790 163.640 ;
        RECT 65.350 163.100 65.590 163.390 ;
        RECT 66.390 163.310 66.560 163.390 ;
        RECT 65.790 162.840 66.210 163.220 ;
        RECT 66.390 163.060 67.020 163.310 ;
        RECT 67.490 162.840 67.820 163.220 ;
        RECT 67.990 163.100 68.160 163.390 ;
        RECT 68.960 163.225 69.130 164.070 ;
        RECT 69.580 163.900 69.800 164.770 ;
        RECT 70.025 164.650 70.720 164.840 ;
        RECT 69.300 163.520 69.800 163.900 ;
        RECT 69.970 163.850 70.380 164.470 ;
        RECT 70.550 163.680 70.720 164.650 ;
        RECT 70.025 163.510 70.720 163.680 ;
        RECT 68.340 162.840 68.720 163.220 ;
        RECT 68.960 163.055 69.790 163.225 ;
        RECT 70.025 163.010 70.195 163.510 ;
        RECT 70.365 162.840 70.695 163.340 ;
        RECT 70.910 163.010 71.135 165.130 ;
        RECT 71.305 165.010 71.635 165.390 ;
        RECT 71.805 164.840 71.975 165.130 ;
        RECT 71.310 164.670 71.975 164.840 ;
        RECT 72.235 164.715 72.495 165.220 ;
        RECT 72.675 165.010 73.005 165.390 ;
        RECT 73.185 164.840 73.355 165.220 ;
        RECT 74.080 164.845 79.425 165.390 ;
        RECT 71.310 163.680 71.540 164.670 ;
        RECT 71.710 163.850 72.060 164.500 ;
        RECT 72.235 163.915 72.405 164.715 ;
        RECT 72.690 164.670 73.355 164.840 ;
        RECT 72.690 164.415 72.860 164.670 ;
        RECT 72.575 164.085 72.860 164.415 ;
        RECT 73.095 164.120 73.425 164.490 ;
        RECT 72.690 163.940 72.860 164.085 ;
        RECT 71.310 163.510 71.975 163.680 ;
        RECT 71.305 162.840 71.635 163.340 ;
        RECT 71.805 163.010 71.975 163.510 ;
        RECT 72.235 163.010 72.505 163.915 ;
        RECT 72.690 163.770 73.355 163.940 ;
        RECT 72.675 162.840 73.005 163.600 ;
        RECT 73.185 163.010 73.355 163.770 ;
        RECT 75.670 163.275 76.020 164.525 ;
        RECT 77.500 164.015 77.840 164.845 ;
        RECT 79.595 164.665 79.885 165.390 ;
        RECT 80.515 164.620 83.105 165.390 ;
        RECT 83.280 164.845 88.625 165.390 ;
        RECT 74.080 162.840 79.425 163.275 ;
        RECT 79.595 162.840 79.885 164.005 ;
        RECT 80.515 163.930 81.725 164.450 ;
        RECT 81.895 164.100 83.105 164.620 ;
        RECT 80.515 162.840 83.105 163.930 ;
        RECT 84.870 163.275 85.220 164.525 ;
        RECT 86.700 164.015 87.040 164.845 ;
        RECT 89.000 164.610 89.500 165.220 ;
        RECT 88.795 164.150 89.145 164.400 ;
        RECT 89.330 163.980 89.500 164.610 ;
        RECT 90.130 164.740 90.460 165.220 ;
        RECT 90.630 164.930 90.855 165.390 ;
        RECT 91.025 164.740 91.355 165.220 ;
        RECT 90.130 164.570 91.355 164.740 ;
        RECT 91.545 164.590 91.795 165.390 ;
        RECT 91.965 164.590 92.305 165.220 ;
        RECT 92.680 164.610 93.180 165.220 ;
        RECT 89.670 164.200 90.000 164.400 ;
        RECT 90.170 164.200 90.500 164.400 ;
        RECT 90.670 164.200 91.090 164.400 ;
        RECT 91.265 164.230 91.960 164.400 ;
        RECT 91.265 163.980 91.435 164.230 ;
        RECT 92.130 163.980 92.305 164.590 ;
        RECT 92.475 164.150 92.825 164.400 ;
        RECT 93.010 163.980 93.180 164.610 ;
        RECT 93.810 164.740 94.140 165.220 ;
        RECT 94.310 164.930 94.535 165.390 ;
        RECT 94.705 164.740 95.035 165.220 ;
        RECT 93.810 164.570 95.035 164.740 ;
        RECT 95.225 164.590 95.475 165.390 ;
        RECT 95.645 164.590 95.985 165.220 ;
        RECT 96.360 164.610 96.860 165.220 ;
        RECT 93.350 164.200 93.680 164.400 ;
        RECT 93.850 164.200 94.180 164.400 ;
        RECT 94.350 164.200 94.770 164.400 ;
        RECT 94.945 164.230 95.640 164.400 ;
        RECT 94.945 163.980 95.115 164.230 ;
        RECT 95.810 163.980 95.985 164.590 ;
        RECT 96.155 164.150 96.505 164.400 ;
        RECT 96.690 163.980 96.860 164.610 ;
        RECT 97.490 164.740 97.820 165.220 ;
        RECT 97.990 164.930 98.215 165.390 ;
        RECT 98.385 164.740 98.715 165.220 ;
        RECT 97.490 164.570 98.715 164.740 ;
        RECT 98.905 164.590 99.155 165.390 ;
        RECT 99.325 164.590 99.665 165.220 ;
        RECT 99.845 164.890 100.175 165.390 ;
        RECT 100.375 164.820 100.545 165.170 ;
        RECT 100.745 164.990 101.075 165.390 ;
        RECT 101.245 164.820 101.415 165.170 ;
        RECT 101.585 164.990 101.965 165.390 ;
        RECT 97.030 164.200 97.360 164.400 ;
        RECT 97.530 164.200 97.860 164.400 ;
        RECT 98.030 164.200 98.450 164.400 ;
        RECT 98.625 164.230 99.320 164.400 ;
        RECT 98.625 163.980 98.795 164.230 ;
        RECT 99.490 163.980 99.665 164.590 ;
        RECT 99.840 164.150 100.190 164.720 ;
        RECT 100.375 164.650 101.985 164.820 ;
        RECT 102.155 164.715 102.425 165.060 ;
        RECT 101.815 164.480 101.985 164.650 ;
        RECT 89.000 163.810 91.435 163.980 ;
        RECT 83.280 162.840 88.625 163.275 ;
        RECT 89.000 163.010 89.330 163.810 ;
        RECT 89.500 162.840 89.830 163.640 ;
        RECT 90.130 163.010 90.460 163.810 ;
        RECT 91.105 162.840 91.355 163.640 ;
        RECT 91.625 162.840 91.795 163.980 ;
        RECT 91.965 163.010 92.305 163.980 ;
        RECT 92.680 163.810 95.115 163.980 ;
        RECT 92.680 163.010 93.010 163.810 ;
        RECT 93.180 162.840 93.510 163.640 ;
        RECT 93.810 163.010 94.140 163.810 ;
        RECT 94.785 162.840 95.035 163.640 ;
        RECT 95.305 162.840 95.475 163.980 ;
        RECT 95.645 163.010 95.985 163.980 ;
        RECT 96.360 163.810 98.795 163.980 ;
        RECT 96.360 163.010 96.690 163.810 ;
        RECT 96.860 162.840 97.190 163.640 ;
        RECT 97.490 163.010 97.820 163.810 ;
        RECT 98.465 162.840 98.715 163.640 ;
        RECT 98.985 162.840 99.155 163.980 ;
        RECT 99.325 163.010 99.665 163.980 ;
        RECT 99.840 163.690 100.160 163.980 ;
        RECT 100.360 163.860 101.070 164.480 ;
        RECT 101.240 164.150 101.645 164.480 ;
        RECT 101.815 164.150 102.085 164.480 ;
        RECT 101.815 163.980 101.985 164.150 ;
        RECT 102.255 163.980 102.425 164.715 ;
        RECT 102.595 164.620 105.185 165.390 ;
        RECT 105.355 164.665 105.645 165.390 ;
        RECT 101.260 163.810 101.985 163.980 ;
        RECT 101.260 163.690 101.430 163.810 ;
        RECT 99.840 163.520 101.430 163.690 ;
        RECT 99.840 163.060 101.495 163.350 ;
        RECT 101.665 162.840 101.945 163.640 ;
        RECT 102.155 163.010 102.425 163.980 ;
        RECT 102.595 163.930 103.805 164.450 ;
        RECT 103.975 164.100 105.185 164.620 ;
        RECT 105.855 164.570 106.085 165.390 ;
        RECT 106.255 164.590 106.585 165.220 ;
        RECT 105.835 164.150 106.165 164.400 ;
        RECT 102.595 162.840 105.185 163.930 ;
        RECT 105.355 162.840 105.645 164.005 ;
        RECT 106.335 163.990 106.585 164.590 ;
        RECT 106.755 164.570 106.965 165.390 ;
        RECT 107.200 164.680 107.455 165.210 ;
        RECT 107.625 164.930 107.930 165.390 ;
        RECT 108.175 165.010 109.245 165.180 ;
        RECT 105.855 162.840 106.085 163.980 ;
        RECT 106.255 163.010 106.585 163.990 ;
        RECT 107.200 164.030 107.410 164.680 ;
        RECT 108.175 164.655 108.495 165.010 ;
        RECT 108.170 164.480 108.495 164.655 ;
        RECT 107.580 164.180 108.495 164.480 ;
        RECT 108.665 164.440 108.905 164.840 ;
        RECT 109.075 164.780 109.245 165.010 ;
        RECT 109.415 164.950 109.605 165.390 ;
        RECT 109.775 164.940 110.725 165.220 ;
        RECT 110.945 165.030 111.295 165.200 ;
        RECT 109.075 164.610 109.605 164.780 ;
        RECT 107.580 164.150 108.320 164.180 ;
        RECT 106.755 162.840 106.965 163.980 ;
        RECT 107.200 163.150 107.455 164.030 ;
        RECT 107.625 162.840 107.930 163.980 ;
        RECT 108.150 163.560 108.320 164.150 ;
        RECT 108.665 164.070 109.205 164.440 ;
        RECT 109.385 164.330 109.605 164.610 ;
        RECT 109.775 164.160 109.945 164.940 ;
        RECT 109.540 163.990 109.945 164.160 ;
        RECT 110.115 164.150 110.465 164.770 ;
        RECT 109.540 163.900 109.710 163.990 ;
        RECT 110.635 163.980 110.845 164.770 ;
        RECT 108.490 163.730 109.710 163.900 ;
        RECT 110.170 163.820 110.845 163.980 ;
        RECT 108.150 163.390 108.950 163.560 ;
        RECT 108.270 162.840 108.600 163.220 ;
        RECT 108.780 163.100 108.950 163.390 ;
        RECT 109.540 163.350 109.710 163.730 ;
        RECT 109.880 163.810 110.845 163.820 ;
        RECT 111.035 164.640 111.295 165.030 ;
        RECT 111.505 164.930 111.835 165.390 ;
        RECT 112.710 165.000 113.565 165.170 ;
        RECT 113.770 165.000 114.265 165.170 ;
        RECT 114.435 165.030 114.765 165.390 ;
        RECT 111.035 163.950 111.205 164.640 ;
        RECT 111.375 164.290 111.545 164.470 ;
        RECT 111.715 164.460 112.505 164.710 ;
        RECT 112.710 164.290 112.880 165.000 ;
        RECT 113.050 164.490 113.405 164.710 ;
        RECT 111.375 164.120 113.065 164.290 ;
        RECT 109.880 163.520 110.340 163.810 ;
        RECT 111.035 163.780 112.535 163.950 ;
        RECT 111.035 163.640 111.205 163.780 ;
        RECT 110.645 163.470 111.205 163.640 ;
        RECT 109.120 162.840 109.370 163.300 ;
        RECT 109.540 163.010 110.410 163.350 ;
        RECT 110.645 163.010 110.815 163.470 ;
        RECT 111.650 163.440 112.725 163.610 ;
        RECT 110.985 162.840 111.355 163.300 ;
        RECT 111.650 163.100 111.820 163.440 ;
        RECT 111.990 162.840 112.320 163.270 ;
        RECT 112.555 163.100 112.725 163.440 ;
        RECT 112.895 163.340 113.065 164.120 ;
        RECT 113.235 163.900 113.405 164.490 ;
        RECT 113.575 164.090 113.925 164.710 ;
        RECT 113.235 163.510 113.700 163.900 ;
        RECT 114.095 163.640 114.265 165.000 ;
        RECT 114.435 163.810 114.895 164.860 ;
        RECT 113.870 163.470 114.265 163.640 ;
        RECT 113.870 163.340 114.040 163.470 ;
        RECT 112.895 163.010 113.575 163.340 ;
        RECT 113.790 163.010 114.040 163.340 ;
        RECT 114.210 162.840 114.460 163.300 ;
        RECT 114.630 163.025 114.955 163.810 ;
        RECT 115.125 163.010 115.295 165.130 ;
        RECT 115.465 165.010 115.795 165.390 ;
        RECT 115.965 164.840 116.220 165.130 ;
        RECT 115.470 164.670 116.220 164.840 ;
        RECT 115.470 163.680 115.700 164.670 ;
        RECT 117.315 164.640 118.525 165.390 ;
        RECT 115.870 163.850 116.220 164.500 ;
        RECT 117.315 163.930 117.835 164.470 ;
        RECT 118.005 164.100 118.525 164.640 ;
        RECT 115.470 163.510 116.220 163.680 ;
        RECT 115.465 162.840 115.795 163.340 ;
        RECT 115.965 163.010 116.220 163.510 ;
        RECT 117.315 162.840 118.525 163.930 ;
        RECT 11.430 162.670 118.610 162.840 ;
        RECT 11.515 161.580 12.725 162.670 ;
        RECT 11.515 160.870 12.035 161.410 ;
        RECT 12.205 161.040 12.725 161.580 ;
        RECT 13.355 161.580 15.025 162.670 ;
        RECT 13.355 161.060 14.105 161.580 ;
        RECT 15.195 161.505 15.485 162.670 ;
        RECT 15.660 161.480 15.915 162.360 ;
        RECT 16.085 161.530 16.390 162.670 ;
        RECT 16.730 162.290 17.060 162.670 ;
        RECT 17.240 162.120 17.410 162.410 ;
        RECT 17.580 162.210 17.830 162.670 ;
        RECT 16.610 161.950 17.410 162.120 ;
        RECT 18.000 162.160 18.870 162.500 ;
        RECT 14.275 160.890 15.025 161.410 ;
        RECT 11.515 160.120 12.725 160.870 ;
        RECT 13.355 160.120 15.025 160.890 ;
        RECT 15.195 160.120 15.485 160.845 ;
        RECT 15.660 160.830 15.870 161.480 ;
        RECT 16.610 161.360 16.780 161.950 ;
        RECT 18.000 161.780 18.170 162.160 ;
        RECT 19.105 162.040 19.275 162.500 ;
        RECT 19.445 162.210 19.815 162.670 ;
        RECT 20.110 162.070 20.280 162.410 ;
        RECT 20.450 162.240 20.780 162.670 ;
        RECT 21.015 162.070 21.185 162.410 ;
        RECT 16.950 161.610 18.170 161.780 ;
        RECT 18.340 161.700 18.800 161.990 ;
        RECT 19.105 161.870 19.665 162.040 ;
        RECT 20.110 161.900 21.185 162.070 ;
        RECT 21.355 162.170 22.035 162.500 ;
        RECT 22.250 162.170 22.500 162.500 ;
        RECT 22.670 162.210 22.920 162.670 ;
        RECT 19.495 161.730 19.665 161.870 ;
        RECT 18.340 161.690 19.305 161.700 ;
        RECT 18.000 161.520 18.170 161.610 ;
        RECT 18.630 161.530 19.305 161.690 ;
        RECT 16.040 161.330 16.780 161.360 ;
        RECT 16.040 161.030 16.955 161.330 ;
        RECT 16.630 160.855 16.955 161.030 ;
        RECT 15.660 160.300 15.915 160.830 ;
        RECT 16.085 160.120 16.390 160.580 ;
        RECT 16.635 160.500 16.955 160.855 ;
        RECT 17.125 161.070 17.665 161.440 ;
        RECT 18.000 161.350 18.405 161.520 ;
        RECT 17.125 160.670 17.365 161.070 ;
        RECT 17.845 160.900 18.065 161.180 ;
        RECT 17.535 160.730 18.065 160.900 ;
        RECT 17.535 160.500 17.705 160.730 ;
        RECT 18.235 160.570 18.405 161.350 ;
        RECT 18.575 160.740 18.925 161.360 ;
        RECT 19.095 160.740 19.305 161.530 ;
        RECT 19.495 161.560 20.995 161.730 ;
        RECT 19.495 160.870 19.665 161.560 ;
        RECT 21.355 161.390 21.525 162.170 ;
        RECT 22.330 162.040 22.500 162.170 ;
        RECT 19.835 161.220 21.525 161.390 ;
        RECT 21.695 161.610 22.160 162.000 ;
        RECT 22.330 161.870 22.725 162.040 ;
        RECT 19.835 161.040 20.005 161.220 ;
        RECT 16.635 160.330 17.705 160.500 ;
        RECT 17.875 160.120 18.065 160.560 ;
        RECT 18.235 160.290 19.185 160.570 ;
        RECT 19.495 160.480 19.755 160.870 ;
        RECT 20.175 160.800 20.965 161.050 ;
        RECT 19.405 160.310 19.755 160.480 ;
        RECT 19.965 160.120 20.295 160.580 ;
        RECT 21.170 160.510 21.340 161.220 ;
        RECT 21.695 161.020 21.865 161.610 ;
        RECT 21.510 160.800 21.865 161.020 ;
        RECT 22.035 160.800 22.385 161.420 ;
        RECT 22.555 160.510 22.725 161.870 ;
        RECT 23.090 161.700 23.415 162.485 ;
        RECT 22.895 160.650 23.355 161.700 ;
        RECT 21.170 160.340 22.025 160.510 ;
        RECT 22.230 160.340 22.725 160.510 ;
        RECT 22.895 160.120 23.225 160.480 ;
        RECT 23.585 160.380 23.755 162.500 ;
        RECT 23.925 162.170 24.255 162.670 ;
        RECT 24.425 162.000 24.680 162.500 ;
        RECT 23.930 161.830 24.680 162.000 ;
        RECT 23.930 160.840 24.160 161.830 ;
        RECT 24.330 161.010 24.680 161.660 ;
        RECT 25.315 161.580 27.905 162.670 ;
        RECT 28.080 162.235 33.425 162.670 ;
        RECT 25.315 161.060 26.525 161.580 ;
        RECT 26.695 160.890 27.905 161.410 ;
        RECT 29.670 160.985 30.020 162.235 ;
        RECT 33.595 161.595 33.865 162.500 ;
        RECT 34.035 161.910 34.365 162.670 ;
        RECT 34.545 161.740 34.715 162.500 ;
        RECT 23.930 160.670 24.680 160.840 ;
        RECT 23.925 160.120 24.255 160.500 ;
        RECT 24.425 160.380 24.680 160.670 ;
        RECT 25.315 160.120 27.905 160.890 ;
        RECT 31.500 160.665 31.840 161.495 ;
        RECT 33.595 160.795 33.765 161.595 ;
        RECT 34.050 161.570 34.715 161.740 ;
        RECT 35.435 161.580 37.105 162.670 ;
        RECT 37.480 161.700 37.810 162.500 ;
        RECT 37.980 161.870 38.310 162.670 ;
        RECT 38.610 161.700 38.940 162.500 ;
        RECT 39.585 161.870 39.835 162.670 ;
        RECT 34.050 161.425 34.220 161.570 ;
        RECT 33.935 161.095 34.220 161.425 ;
        RECT 34.050 160.840 34.220 161.095 ;
        RECT 34.455 161.020 34.785 161.390 ;
        RECT 35.435 161.060 36.185 161.580 ;
        RECT 37.480 161.530 39.915 161.700 ;
        RECT 40.105 161.530 40.275 162.670 ;
        RECT 40.445 161.530 40.785 162.500 ;
        RECT 36.355 160.890 37.105 161.410 ;
        RECT 37.275 161.110 37.625 161.360 ;
        RECT 37.810 160.900 37.980 161.530 ;
        RECT 38.150 161.110 38.480 161.310 ;
        RECT 38.650 161.110 38.980 161.310 ;
        RECT 39.150 161.110 39.570 161.310 ;
        RECT 39.745 161.280 39.915 161.530 ;
        RECT 39.745 161.110 40.440 161.280 ;
        RECT 28.080 160.120 33.425 160.665 ;
        RECT 33.595 160.290 33.855 160.795 ;
        RECT 34.050 160.670 34.715 160.840 ;
        RECT 34.035 160.120 34.365 160.500 ;
        RECT 34.545 160.290 34.715 160.670 ;
        RECT 35.435 160.120 37.105 160.890 ;
        RECT 37.480 160.290 37.980 160.900 ;
        RECT 38.610 160.770 39.835 160.940 ;
        RECT 40.610 160.920 40.785 161.530 ;
        RECT 40.955 161.505 41.245 162.670 ;
        RECT 42.335 161.530 42.675 162.500 ;
        RECT 42.845 161.530 43.015 162.670 ;
        RECT 43.285 161.870 43.535 162.670 ;
        RECT 44.180 161.700 44.510 162.500 ;
        RECT 44.810 161.870 45.140 162.670 ;
        RECT 45.310 161.700 45.640 162.500 ;
        RECT 43.205 161.530 45.640 161.700 ;
        RECT 46.015 161.580 47.225 162.670 ;
        RECT 47.400 162.280 47.735 162.500 ;
        RECT 48.740 162.290 49.095 162.670 ;
        RECT 47.400 161.660 47.655 162.280 ;
        RECT 47.905 162.120 48.135 162.160 ;
        RECT 49.265 162.120 49.515 162.500 ;
        RECT 47.905 161.920 49.515 162.120 ;
        RECT 47.905 161.830 48.090 161.920 ;
        RECT 48.680 161.910 49.515 161.920 ;
        RECT 49.765 161.890 50.015 162.670 ;
        RECT 50.185 161.820 50.445 162.500 ;
        RECT 48.245 161.720 48.575 161.750 ;
        RECT 48.245 161.660 50.045 161.720 ;
        RECT 38.610 160.290 38.940 160.770 ;
        RECT 39.110 160.120 39.335 160.580 ;
        RECT 39.505 160.290 39.835 160.770 ;
        RECT 40.025 160.120 40.275 160.920 ;
        RECT 40.445 160.290 40.785 160.920 ;
        RECT 42.335 160.920 42.510 161.530 ;
        RECT 43.205 161.280 43.375 161.530 ;
        RECT 42.680 161.110 43.375 161.280 ;
        RECT 43.550 161.110 43.970 161.310 ;
        RECT 44.140 161.110 44.470 161.310 ;
        RECT 44.640 161.110 44.970 161.310 ;
        RECT 40.955 160.120 41.245 160.845 ;
        RECT 42.335 160.290 42.675 160.920 ;
        RECT 42.845 160.120 43.095 160.920 ;
        RECT 43.285 160.770 44.510 160.940 ;
        RECT 43.285 160.290 43.615 160.770 ;
        RECT 43.785 160.120 44.010 160.580 ;
        RECT 44.180 160.290 44.510 160.770 ;
        RECT 45.140 160.900 45.310 161.530 ;
        RECT 45.495 161.110 45.845 161.360 ;
        RECT 46.015 161.040 46.535 161.580 ;
        RECT 47.400 161.550 50.105 161.660 ;
        RECT 47.400 161.490 48.575 161.550 ;
        RECT 49.905 161.515 50.105 161.550 ;
        RECT 45.140 160.290 45.640 160.900 ;
        RECT 46.705 160.870 47.225 161.410 ;
        RECT 47.395 161.110 47.885 161.310 ;
        RECT 48.075 161.110 48.550 161.320 ;
        RECT 46.015 160.120 47.225 160.870 ;
        RECT 47.400 160.120 47.855 160.885 ;
        RECT 48.330 160.710 48.550 161.110 ;
        RECT 48.795 161.110 49.125 161.320 ;
        RECT 48.795 160.710 49.005 161.110 ;
        RECT 49.295 161.075 49.705 161.380 ;
        RECT 49.935 160.940 50.105 161.515 ;
        RECT 49.835 160.820 50.105 160.940 ;
        RECT 49.260 160.775 50.105 160.820 ;
        RECT 49.260 160.650 50.015 160.775 ;
        RECT 49.260 160.500 49.430 160.650 ;
        RECT 50.275 160.620 50.445 161.820 ;
        RECT 48.130 160.290 49.430 160.500 ;
        RECT 49.685 160.120 50.015 160.480 ;
        RECT 50.185 160.290 50.445 160.620 ;
        RECT 50.615 161.530 50.955 162.500 ;
        RECT 51.125 161.530 51.295 162.670 ;
        RECT 51.565 161.870 51.815 162.670 ;
        RECT 52.460 161.700 52.790 162.500 ;
        RECT 53.090 161.870 53.420 162.670 ;
        RECT 53.590 161.700 53.920 162.500 ;
        RECT 51.485 161.530 53.920 161.700 ;
        RECT 54.295 161.530 54.635 162.500 ;
        RECT 54.805 161.530 54.975 162.670 ;
        RECT 55.245 161.870 55.495 162.670 ;
        RECT 56.140 161.700 56.470 162.500 ;
        RECT 56.770 161.870 57.100 162.670 ;
        RECT 57.270 161.700 57.600 162.500 ;
        RECT 55.165 161.530 57.600 161.700 ;
        RECT 57.975 161.580 59.645 162.670 ;
        RECT 59.815 161.910 60.330 162.320 ;
        RECT 60.565 161.910 60.735 162.670 ;
        RECT 60.905 162.330 62.935 162.500 ;
        RECT 50.615 160.920 50.790 161.530 ;
        RECT 51.485 161.280 51.655 161.530 ;
        RECT 50.960 161.110 51.655 161.280 ;
        RECT 51.830 161.110 52.250 161.310 ;
        RECT 52.420 161.110 52.750 161.310 ;
        RECT 52.920 161.110 53.250 161.310 ;
        RECT 50.615 160.290 50.955 160.920 ;
        RECT 51.125 160.120 51.375 160.920 ;
        RECT 51.565 160.770 52.790 160.940 ;
        RECT 51.565 160.290 51.895 160.770 ;
        RECT 52.065 160.120 52.290 160.580 ;
        RECT 52.460 160.290 52.790 160.770 ;
        RECT 53.420 160.900 53.590 161.530 ;
        RECT 54.295 161.480 54.525 161.530 ;
        RECT 53.775 161.110 54.125 161.360 ;
        RECT 54.295 160.920 54.470 161.480 ;
        RECT 55.165 161.280 55.335 161.530 ;
        RECT 54.640 161.110 55.335 161.280 ;
        RECT 55.510 161.110 55.930 161.310 ;
        RECT 56.100 161.110 56.430 161.310 ;
        RECT 56.600 161.110 56.930 161.310 ;
        RECT 53.420 160.290 53.920 160.900 ;
        RECT 54.295 160.290 54.635 160.920 ;
        RECT 54.805 160.120 55.055 160.920 ;
        RECT 55.245 160.770 56.470 160.940 ;
        RECT 55.245 160.290 55.575 160.770 ;
        RECT 55.745 160.120 55.970 160.580 ;
        RECT 56.140 160.290 56.470 160.770 ;
        RECT 57.100 160.900 57.270 161.530 ;
        RECT 57.455 161.110 57.805 161.360 ;
        RECT 57.975 161.060 58.725 161.580 ;
        RECT 57.100 160.290 57.600 160.900 ;
        RECT 58.895 160.890 59.645 161.410 ;
        RECT 59.815 161.100 60.155 161.910 ;
        RECT 60.905 161.665 61.075 162.330 ;
        RECT 61.470 161.990 62.595 162.160 ;
        RECT 60.325 161.475 61.075 161.665 ;
        RECT 61.245 161.650 62.255 161.820 ;
        RECT 59.815 160.930 61.045 161.100 ;
        RECT 57.975 160.120 59.645 160.890 ;
        RECT 60.090 160.325 60.335 160.930 ;
        RECT 60.555 160.120 61.065 160.655 ;
        RECT 61.245 160.290 61.435 161.650 ;
        RECT 61.605 160.630 61.880 161.450 ;
        RECT 62.085 160.850 62.255 161.650 ;
        RECT 62.425 160.860 62.595 161.990 ;
        RECT 62.765 161.360 62.935 162.330 ;
        RECT 63.105 161.530 63.275 162.670 ;
        RECT 63.445 161.530 63.780 162.500 ;
        RECT 62.765 161.030 62.960 161.360 ;
        RECT 63.185 161.030 63.440 161.360 ;
        RECT 63.185 160.860 63.355 161.030 ;
        RECT 63.610 160.860 63.780 161.530 ;
        RECT 63.955 161.580 66.545 162.670 ;
        RECT 63.955 161.060 65.165 161.580 ;
        RECT 66.715 161.505 67.005 162.670 ;
        RECT 68.100 161.520 68.360 162.670 ;
        RECT 68.535 161.595 68.790 162.500 ;
        RECT 68.960 161.910 69.290 162.670 ;
        RECT 69.505 161.740 69.675 162.500 ;
        RECT 65.335 160.890 66.545 161.410 ;
        RECT 62.425 160.690 63.355 160.860 ;
        RECT 62.425 160.655 62.600 160.690 ;
        RECT 61.605 160.460 61.885 160.630 ;
        RECT 61.605 160.290 61.880 160.460 ;
        RECT 62.070 160.290 62.600 160.655 ;
        RECT 63.025 160.120 63.355 160.520 ;
        RECT 63.525 160.290 63.780 160.860 ;
        RECT 63.955 160.120 66.545 160.890 ;
        RECT 66.715 160.120 67.005 160.845 ;
        RECT 68.100 160.120 68.360 160.960 ;
        RECT 68.535 160.865 68.705 161.595 ;
        RECT 68.960 161.570 69.675 161.740 ;
        RECT 69.935 161.580 73.445 162.670 ;
        RECT 73.620 162.235 78.965 162.670 ;
        RECT 79.140 162.235 84.485 162.670 ;
        RECT 68.960 161.360 69.130 161.570 ;
        RECT 68.875 161.030 69.130 161.360 ;
        RECT 68.535 160.290 68.790 160.865 ;
        RECT 68.960 160.840 69.130 161.030 ;
        RECT 69.410 161.020 69.765 161.390 ;
        RECT 69.935 161.060 71.625 161.580 ;
        RECT 71.795 160.890 73.445 161.410 ;
        RECT 75.210 160.985 75.560 162.235 ;
        RECT 68.960 160.670 69.675 160.840 ;
        RECT 68.960 160.120 69.290 160.500 ;
        RECT 69.505 160.290 69.675 160.670 ;
        RECT 69.935 160.120 73.445 160.890 ;
        RECT 77.040 160.665 77.380 161.495 ;
        RECT 80.730 160.985 81.080 162.235 ;
        RECT 84.745 161.740 84.915 162.500 ;
        RECT 85.095 161.910 85.425 162.670 ;
        RECT 84.745 161.570 85.410 161.740 ;
        RECT 85.595 161.595 85.865 162.500 ;
        RECT 82.560 160.665 82.900 161.495 ;
        RECT 85.240 161.425 85.410 161.570 ;
        RECT 84.675 161.020 85.005 161.390 ;
        RECT 85.240 161.095 85.525 161.425 ;
        RECT 85.240 160.840 85.410 161.095 ;
        RECT 84.745 160.670 85.410 160.840 ;
        RECT 85.695 160.795 85.865 161.595 ;
        RECT 86.035 161.580 88.625 162.670 ;
        RECT 89.000 161.700 89.330 162.500 ;
        RECT 89.500 161.870 89.830 162.670 ;
        RECT 90.130 161.700 90.460 162.500 ;
        RECT 91.105 161.870 91.355 162.670 ;
        RECT 86.035 161.060 87.245 161.580 ;
        RECT 89.000 161.530 91.435 161.700 ;
        RECT 91.625 161.530 91.795 162.670 ;
        RECT 91.965 161.530 92.305 162.500 ;
        RECT 87.415 160.890 88.625 161.410 ;
        RECT 88.795 161.110 89.145 161.360 ;
        RECT 89.330 160.900 89.500 161.530 ;
        RECT 89.670 161.110 90.000 161.310 ;
        RECT 90.170 161.110 90.500 161.310 ;
        RECT 90.670 161.110 91.090 161.310 ;
        RECT 91.265 161.280 91.435 161.530 ;
        RECT 91.265 161.110 91.960 161.280 ;
        RECT 73.620 160.120 78.965 160.665 ;
        RECT 79.140 160.120 84.485 160.665 ;
        RECT 84.745 160.290 84.915 160.670 ;
        RECT 85.095 160.120 85.425 160.500 ;
        RECT 85.605 160.290 85.865 160.795 ;
        RECT 86.035 160.120 88.625 160.890 ;
        RECT 89.000 160.290 89.500 160.900 ;
        RECT 90.130 160.770 91.355 160.940 ;
        RECT 92.130 160.920 92.305 161.530 ;
        RECT 92.475 161.505 92.765 162.670 ;
        RECT 93.600 161.700 93.930 162.500 ;
        RECT 94.100 161.870 94.430 162.670 ;
        RECT 94.730 161.700 95.060 162.500 ;
        RECT 95.705 161.870 95.955 162.670 ;
        RECT 93.600 161.530 96.035 161.700 ;
        RECT 96.225 161.530 96.395 162.670 ;
        RECT 96.565 161.530 96.905 162.500 ;
        RECT 93.395 161.110 93.745 161.360 ;
        RECT 90.130 160.290 90.460 160.770 ;
        RECT 90.630 160.120 90.855 160.580 ;
        RECT 91.025 160.290 91.355 160.770 ;
        RECT 91.545 160.120 91.795 160.920 ;
        RECT 91.965 160.290 92.305 160.920 ;
        RECT 93.930 160.900 94.100 161.530 ;
        RECT 94.270 161.110 94.600 161.310 ;
        RECT 94.770 161.110 95.100 161.310 ;
        RECT 95.270 161.110 95.690 161.310 ;
        RECT 95.865 161.280 96.035 161.530 ;
        RECT 95.865 161.110 96.560 161.280 ;
        RECT 92.475 160.120 92.765 160.845 ;
        RECT 93.600 160.290 94.100 160.900 ;
        RECT 94.730 160.770 95.955 160.940 ;
        RECT 96.730 160.920 96.905 161.530 ;
        RECT 97.075 161.580 98.745 162.670 ;
        RECT 98.920 162.160 100.575 162.450 ;
        RECT 98.920 161.820 100.510 161.990 ;
        RECT 100.745 161.870 101.025 162.670 ;
        RECT 97.075 161.060 97.825 161.580 ;
        RECT 98.920 161.530 99.240 161.820 ;
        RECT 100.340 161.700 100.510 161.820 ;
        RECT 99.435 161.480 100.150 161.650 ;
        RECT 100.340 161.530 101.065 161.700 ;
        RECT 101.235 161.530 101.505 162.500 ;
        RECT 94.730 160.290 95.060 160.770 ;
        RECT 95.230 160.120 95.455 160.580 ;
        RECT 95.625 160.290 95.955 160.770 ;
        RECT 96.145 160.120 96.395 160.920 ;
        RECT 96.565 160.290 96.905 160.920 ;
        RECT 97.995 160.890 98.745 161.410 ;
        RECT 97.075 160.120 98.745 160.890 ;
        RECT 98.920 160.790 99.270 161.360 ;
        RECT 99.440 161.030 100.150 161.480 ;
        RECT 100.895 161.360 101.065 161.530 ;
        RECT 100.320 161.030 100.725 161.360 ;
        RECT 100.895 161.030 101.165 161.360 ;
        RECT 100.895 160.860 101.065 161.030 ;
        RECT 99.455 160.690 101.065 160.860 ;
        RECT 101.335 160.795 101.505 161.530 ;
        RECT 98.925 160.120 99.255 160.620 ;
        RECT 99.455 160.340 99.625 160.690 ;
        RECT 99.825 160.120 100.155 160.520 ;
        RECT 100.325 160.340 100.495 160.690 ;
        RECT 100.665 160.120 101.045 160.520 ;
        RECT 101.235 160.450 101.505 160.795 ;
        RECT 101.675 161.530 102.015 162.500 ;
        RECT 102.185 161.530 102.355 162.670 ;
        RECT 102.625 161.870 102.875 162.670 ;
        RECT 103.520 161.700 103.850 162.500 ;
        RECT 104.150 161.870 104.480 162.670 ;
        RECT 104.650 161.700 104.980 162.500 ;
        RECT 102.545 161.530 104.980 161.700 ;
        RECT 105.815 161.910 106.330 162.320 ;
        RECT 106.565 161.910 106.735 162.670 ;
        RECT 106.905 162.330 108.935 162.500 ;
        RECT 101.675 160.920 101.850 161.530 ;
        RECT 102.545 161.280 102.715 161.530 ;
        RECT 102.020 161.110 102.715 161.280 ;
        RECT 102.890 161.110 103.310 161.310 ;
        RECT 103.480 161.110 103.810 161.310 ;
        RECT 103.980 161.110 104.310 161.310 ;
        RECT 101.675 160.290 102.015 160.920 ;
        RECT 102.185 160.120 102.435 160.920 ;
        RECT 102.625 160.770 103.850 160.940 ;
        RECT 102.625 160.290 102.955 160.770 ;
        RECT 103.125 160.120 103.350 160.580 ;
        RECT 103.520 160.290 103.850 160.770 ;
        RECT 104.480 160.900 104.650 161.530 ;
        RECT 104.835 161.110 105.185 161.360 ;
        RECT 105.815 161.100 106.155 161.910 ;
        RECT 106.905 161.665 107.075 162.330 ;
        RECT 107.470 161.990 108.595 162.160 ;
        RECT 106.325 161.475 107.075 161.665 ;
        RECT 107.245 161.650 108.255 161.820 ;
        RECT 105.815 160.930 107.045 161.100 ;
        RECT 104.480 160.290 104.980 160.900 ;
        RECT 106.090 160.325 106.335 160.930 ;
        RECT 106.555 160.120 107.065 160.655 ;
        RECT 107.245 160.290 107.435 161.650 ;
        RECT 107.605 160.630 107.880 161.450 ;
        RECT 108.085 160.850 108.255 161.650 ;
        RECT 108.425 160.860 108.595 161.990 ;
        RECT 108.765 161.360 108.935 162.330 ;
        RECT 109.105 161.530 109.275 162.670 ;
        RECT 109.445 161.530 109.780 162.500 ;
        RECT 110.455 161.530 110.685 162.670 ;
        RECT 108.765 161.030 108.960 161.360 ;
        RECT 109.185 161.030 109.440 161.360 ;
        RECT 109.185 160.860 109.355 161.030 ;
        RECT 109.610 160.860 109.780 161.530 ;
        RECT 110.855 161.520 111.185 162.500 ;
        RECT 111.355 161.530 111.565 162.670 ;
        RECT 112.805 161.740 112.975 162.500 ;
        RECT 113.155 161.910 113.485 162.670 ;
        RECT 112.805 161.570 113.470 161.740 ;
        RECT 113.655 161.595 113.925 162.500 ;
        RECT 110.435 161.110 110.765 161.360 ;
        RECT 108.425 160.690 109.355 160.860 ;
        RECT 108.425 160.655 108.600 160.690 ;
        RECT 107.605 160.460 107.885 160.630 ;
        RECT 107.605 160.290 107.880 160.460 ;
        RECT 108.070 160.290 108.600 160.655 ;
        RECT 109.025 160.120 109.355 160.520 ;
        RECT 109.525 160.290 109.780 160.860 ;
        RECT 110.455 160.120 110.685 160.940 ;
        RECT 110.935 160.920 111.185 161.520 ;
        RECT 113.300 161.425 113.470 161.570 ;
        RECT 112.735 161.020 113.065 161.390 ;
        RECT 113.300 161.095 113.585 161.425 ;
        RECT 110.855 160.290 111.185 160.920 ;
        RECT 111.355 160.120 111.565 160.940 ;
        RECT 113.300 160.840 113.470 161.095 ;
        RECT 112.805 160.670 113.470 160.840 ;
        RECT 113.755 160.795 113.925 161.595 ;
        RECT 114.185 161.740 114.355 162.500 ;
        RECT 114.535 161.910 114.865 162.670 ;
        RECT 114.185 161.570 114.850 161.740 ;
        RECT 115.035 161.595 115.305 162.500 ;
        RECT 114.680 161.425 114.850 161.570 ;
        RECT 114.115 161.020 114.445 161.390 ;
        RECT 114.680 161.095 114.965 161.425 ;
        RECT 114.680 160.840 114.850 161.095 ;
        RECT 112.805 160.290 112.975 160.670 ;
        RECT 113.155 160.120 113.485 160.500 ;
        RECT 113.665 160.290 113.925 160.795 ;
        RECT 114.185 160.670 114.850 160.840 ;
        RECT 115.135 160.795 115.305 161.595 ;
        RECT 115.475 161.580 117.145 162.670 ;
        RECT 117.315 161.580 118.525 162.670 ;
        RECT 115.475 161.060 116.225 161.580 ;
        RECT 116.395 160.890 117.145 161.410 ;
        RECT 117.315 161.040 117.835 161.580 ;
        RECT 114.185 160.290 114.355 160.670 ;
        RECT 114.535 160.120 114.865 160.500 ;
        RECT 115.045 160.290 115.305 160.795 ;
        RECT 115.475 160.120 117.145 160.890 ;
        RECT 118.005 160.870 118.525 161.410 ;
        RECT 117.315 160.120 118.525 160.870 ;
        RECT 11.430 159.950 118.610 160.120 ;
        RECT 11.515 159.200 12.725 159.950 ;
        RECT 12.900 159.405 18.245 159.950 ;
        RECT 11.515 158.660 12.035 159.200 ;
        RECT 12.205 158.490 12.725 159.030 ;
        RECT 11.515 157.400 12.725 158.490 ;
        RECT 14.490 157.835 14.840 159.085 ;
        RECT 16.320 158.575 16.660 159.405 ;
        RECT 18.420 159.210 18.675 159.780 ;
        RECT 18.845 159.550 19.175 159.950 ;
        RECT 19.600 159.415 20.130 159.780 ;
        RECT 19.600 159.380 19.775 159.415 ;
        RECT 18.845 159.210 19.775 159.380 ;
        RECT 18.420 158.540 18.590 159.210 ;
        RECT 18.845 159.040 19.015 159.210 ;
        RECT 18.760 158.710 19.015 159.040 ;
        RECT 19.240 158.710 19.435 159.040 ;
        RECT 12.900 157.400 18.245 157.835 ;
        RECT 18.420 157.570 18.755 158.540 ;
        RECT 18.925 157.400 19.095 158.540 ;
        RECT 19.265 157.740 19.435 158.710 ;
        RECT 19.605 158.080 19.775 159.210 ;
        RECT 19.945 158.420 20.115 159.220 ;
        RECT 20.320 158.930 20.595 159.780 ;
        RECT 20.315 158.760 20.595 158.930 ;
        RECT 20.320 158.620 20.595 158.760 ;
        RECT 20.765 158.420 20.955 159.780 ;
        RECT 21.135 159.415 21.645 159.950 ;
        RECT 21.865 159.140 22.110 159.745 ;
        RECT 22.560 159.405 27.905 159.950 ;
        RECT 21.155 158.970 22.385 159.140 ;
        RECT 19.945 158.250 20.955 158.420 ;
        RECT 21.125 158.405 21.875 158.595 ;
        RECT 19.605 157.910 20.730 158.080 ;
        RECT 21.125 157.740 21.295 158.405 ;
        RECT 22.045 158.160 22.385 158.970 ;
        RECT 19.265 157.570 21.295 157.740 ;
        RECT 21.465 157.400 21.635 158.160 ;
        RECT 21.870 157.750 22.385 158.160 ;
        RECT 24.150 157.835 24.500 159.085 ;
        RECT 25.980 158.575 26.320 159.405 ;
        RECT 28.075 159.225 28.365 159.950 ;
        RECT 28.535 159.180 30.205 159.950 ;
        RECT 22.560 157.400 27.905 157.835 ;
        RECT 28.075 157.400 28.365 158.565 ;
        RECT 28.535 158.490 29.285 159.010 ;
        RECT 29.455 158.660 30.205 159.180 ;
        RECT 30.650 159.140 30.895 159.745 ;
        RECT 31.115 159.415 31.625 159.950 ;
        RECT 30.375 158.970 31.605 159.140 ;
        RECT 28.535 157.400 30.205 158.490 ;
        RECT 30.375 158.160 30.715 158.970 ;
        RECT 30.885 158.405 31.635 158.595 ;
        RECT 30.375 157.750 30.890 158.160 ;
        RECT 31.125 157.400 31.295 158.160 ;
        RECT 31.465 157.740 31.635 158.405 ;
        RECT 31.805 158.420 31.995 159.780 ;
        RECT 32.165 159.610 32.440 159.780 ;
        RECT 32.165 159.440 32.445 159.610 ;
        RECT 32.165 158.620 32.440 159.440 ;
        RECT 32.630 159.415 33.160 159.780 ;
        RECT 33.585 159.550 33.915 159.950 ;
        RECT 32.985 159.380 33.160 159.415 ;
        RECT 32.645 158.420 32.815 159.220 ;
        RECT 31.805 158.250 32.815 158.420 ;
        RECT 32.985 159.210 33.915 159.380 ;
        RECT 34.085 159.210 34.340 159.780 ;
        RECT 32.985 158.080 33.155 159.210 ;
        RECT 33.745 159.040 33.915 159.210 ;
        RECT 32.030 157.910 33.155 158.080 ;
        RECT 33.325 158.710 33.520 159.040 ;
        RECT 33.745 158.710 34.000 159.040 ;
        RECT 33.325 157.740 33.495 158.710 ;
        RECT 34.170 158.540 34.340 159.210 ;
        RECT 31.465 157.570 33.495 157.740 ;
        RECT 33.665 157.400 33.835 158.540 ;
        RECT 34.005 157.570 34.340 158.540 ;
        RECT 34.515 159.275 34.775 159.780 ;
        RECT 34.955 159.570 35.285 159.950 ;
        RECT 35.465 159.400 35.635 159.780 ;
        RECT 34.515 158.475 34.685 159.275 ;
        RECT 34.970 159.230 35.635 159.400 ;
        RECT 34.970 158.975 35.140 159.230 ;
        RECT 35.895 159.180 37.565 159.950 ;
        RECT 34.855 158.645 35.140 158.975 ;
        RECT 35.375 158.680 35.705 159.050 ;
        RECT 34.970 158.500 35.140 158.645 ;
        RECT 34.515 157.570 34.785 158.475 ;
        RECT 34.970 158.330 35.635 158.500 ;
        RECT 34.955 157.400 35.285 158.160 ;
        RECT 35.465 157.570 35.635 158.330 ;
        RECT 35.895 158.490 36.645 159.010 ;
        RECT 36.815 158.660 37.565 159.180 ;
        RECT 37.735 159.275 38.005 159.620 ;
        RECT 38.195 159.550 38.575 159.950 ;
        RECT 38.745 159.380 38.915 159.730 ;
        RECT 39.085 159.550 39.415 159.950 ;
        RECT 39.615 159.380 39.785 159.730 ;
        RECT 39.985 159.450 40.315 159.950 ;
        RECT 37.735 158.540 37.905 159.275 ;
        RECT 38.175 159.210 39.785 159.380 ;
        RECT 38.175 159.040 38.345 159.210 ;
        RECT 38.075 158.710 38.345 159.040 ;
        RECT 38.515 158.710 38.920 159.040 ;
        RECT 38.175 158.540 38.345 158.710 ;
        RECT 39.090 158.590 39.800 159.040 ;
        RECT 39.970 158.710 40.320 159.280 ;
        RECT 40.495 159.275 40.765 159.620 ;
        RECT 40.955 159.550 41.335 159.950 ;
        RECT 41.505 159.380 41.675 159.730 ;
        RECT 41.845 159.550 42.175 159.950 ;
        RECT 42.375 159.380 42.545 159.730 ;
        RECT 42.745 159.450 43.075 159.950 ;
        RECT 35.895 157.400 37.565 158.490 ;
        RECT 37.735 157.570 38.005 158.540 ;
        RECT 38.175 158.370 38.900 158.540 ;
        RECT 39.090 158.420 39.805 158.590 ;
        RECT 40.495 158.540 40.665 159.275 ;
        RECT 40.935 159.210 42.545 159.380 ;
        RECT 40.935 159.040 41.105 159.210 ;
        RECT 40.835 158.710 41.105 159.040 ;
        RECT 41.275 158.710 41.680 159.040 ;
        RECT 40.935 158.540 41.105 158.710 ;
        RECT 38.730 158.250 38.900 158.370 ;
        RECT 40.000 158.250 40.320 158.540 ;
        RECT 38.215 157.400 38.495 158.200 ;
        RECT 38.730 158.080 40.320 158.250 ;
        RECT 38.665 157.620 40.320 157.910 ;
        RECT 40.495 157.570 40.765 158.540 ;
        RECT 40.935 158.370 41.660 158.540 ;
        RECT 41.850 158.420 42.560 159.040 ;
        RECT 42.730 158.710 43.080 159.280 ;
        RECT 43.460 159.170 43.960 159.780 ;
        RECT 43.255 158.710 43.605 158.960 ;
        RECT 43.790 158.540 43.960 159.170 ;
        RECT 44.590 159.300 44.920 159.780 ;
        RECT 45.090 159.490 45.315 159.950 ;
        RECT 45.485 159.300 45.815 159.780 ;
        RECT 44.590 159.130 45.815 159.300 ;
        RECT 46.005 159.150 46.255 159.950 ;
        RECT 46.425 159.150 46.765 159.780 ;
        RECT 44.130 158.760 44.460 158.960 ;
        RECT 44.630 158.760 44.960 158.960 ;
        RECT 45.130 158.760 45.550 158.960 ;
        RECT 45.725 158.790 46.420 158.960 ;
        RECT 45.725 158.540 45.895 158.790 ;
        RECT 46.590 158.590 46.765 159.150 ;
        RECT 46.535 158.540 46.765 158.590 ;
        RECT 41.490 158.250 41.660 158.370 ;
        RECT 42.760 158.250 43.080 158.540 ;
        RECT 40.975 157.400 41.255 158.200 ;
        RECT 41.490 158.080 43.080 158.250 ;
        RECT 43.460 158.370 45.895 158.540 ;
        RECT 41.425 157.620 43.080 157.910 ;
        RECT 43.460 157.570 43.790 158.370 ;
        RECT 43.960 157.400 44.290 158.200 ;
        RECT 44.590 157.570 44.920 158.370 ;
        RECT 45.565 157.400 45.815 158.200 ;
        RECT 46.085 157.400 46.255 158.540 ;
        RECT 46.425 157.570 46.765 158.540 ;
        RECT 46.935 159.275 47.205 159.620 ;
        RECT 47.395 159.550 47.775 159.950 ;
        RECT 47.945 159.380 48.115 159.730 ;
        RECT 48.285 159.550 48.615 159.950 ;
        RECT 48.815 159.380 48.985 159.730 ;
        RECT 49.185 159.450 49.515 159.950 ;
        RECT 46.935 158.540 47.105 159.275 ;
        RECT 47.375 159.210 48.985 159.380 ;
        RECT 47.375 159.040 47.545 159.210 ;
        RECT 47.275 158.710 47.545 159.040 ;
        RECT 47.715 158.710 48.120 159.040 ;
        RECT 47.375 158.540 47.545 158.710 ;
        RECT 46.935 157.570 47.205 158.540 ;
        RECT 47.375 158.370 48.100 158.540 ;
        RECT 48.290 158.420 49.000 159.040 ;
        RECT 49.170 158.710 49.520 159.280 ;
        RECT 50.155 159.180 53.665 159.950 ;
        RECT 53.835 159.225 54.125 159.950 ;
        RECT 54.295 159.180 55.965 159.950 ;
        RECT 56.225 159.470 56.525 159.950 ;
        RECT 56.695 159.300 56.955 159.755 ;
        RECT 57.125 159.470 57.385 159.950 ;
        RECT 57.565 159.300 57.825 159.755 ;
        RECT 57.995 159.470 58.245 159.950 ;
        RECT 58.425 159.300 58.685 159.755 ;
        RECT 58.855 159.470 59.105 159.950 ;
        RECT 59.285 159.300 59.545 159.755 ;
        RECT 59.715 159.470 59.960 159.950 ;
        RECT 60.130 159.300 60.405 159.755 ;
        RECT 60.575 159.470 60.820 159.950 ;
        RECT 60.990 159.300 61.250 159.755 ;
        RECT 61.420 159.470 61.680 159.950 ;
        RECT 61.850 159.300 62.110 159.755 ;
        RECT 62.280 159.470 62.540 159.950 ;
        RECT 62.710 159.300 62.970 159.755 ;
        RECT 63.140 159.390 63.400 159.950 ;
        RECT 47.930 158.250 48.100 158.370 ;
        RECT 49.200 158.250 49.520 158.540 ;
        RECT 47.415 157.400 47.695 158.200 ;
        RECT 47.930 158.080 49.520 158.250 ;
        RECT 50.155 158.490 51.845 159.010 ;
        RECT 52.015 158.660 53.665 159.180 ;
        RECT 47.865 157.620 49.520 157.910 ;
        RECT 50.155 157.400 53.665 158.490 ;
        RECT 53.835 157.400 54.125 158.565 ;
        RECT 54.295 158.490 55.045 159.010 ;
        RECT 55.215 158.660 55.965 159.180 ;
        RECT 56.225 159.130 62.970 159.300 ;
        RECT 56.225 158.540 57.390 159.130 ;
        RECT 63.570 158.960 63.820 159.770 ;
        RECT 64.000 159.425 64.260 159.950 ;
        RECT 64.430 158.960 64.680 159.770 ;
        RECT 64.860 159.440 65.165 159.950 ;
        RECT 57.560 158.710 64.680 158.960 ;
        RECT 64.850 158.710 65.165 159.270 ;
        RECT 65.340 159.110 65.600 159.950 ;
        RECT 65.775 159.205 66.030 159.780 ;
        RECT 66.200 159.570 66.530 159.950 ;
        RECT 66.745 159.400 66.915 159.780 ;
        RECT 66.200 159.230 66.915 159.400 ;
        RECT 54.295 157.400 55.965 158.490 ;
        RECT 56.225 158.315 62.970 158.540 ;
        RECT 56.225 157.400 56.495 158.145 ;
        RECT 56.665 157.575 56.955 158.315 ;
        RECT 57.565 158.300 62.970 158.315 ;
        RECT 57.125 157.405 57.380 158.130 ;
        RECT 57.565 157.575 57.825 158.300 ;
        RECT 57.995 157.405 58.240 158.130 ;
        RECT 58.425 157.575 58.685 158.300 ;
        RECT 58.855 157.405 59.100 158.130 ;
        RECT 59.285 157.575 59.545 158.300 ;
        RECT 59.715 157.405 59.960 158.130 ;
        RECT 60.130 157.575 60.390 158.300 ;
        RECT 60.560 157.405 60.820 158.130 ;
        RECT 60.990 157.575 61.250 158.300 ;
        RECT 61.420 157.405 61.680 158.130 ;
        RECT 61.850 157.575 62.110 158.300 ;
        RECT 62.280 157.405 62.540 158.130 ;
        RECT 62.710 157.575 62.970 158.300 ;
        RECT 63.140 157.405 63.400 158.200 ;
        RECT 63.570 157.575 63.820 158.710 ;
        RECT 57.125 157.400 63.400 157.405 ;
        RECT 64.000 157.400 64.260 158.210 ;
        RECT 64.435 157.570 64.680 158.710 ;
        RECT 64.860 157.400 65.155 158.210 ;
        RECT 65.340 157.400 65.600 158.550 ;
        RECT 65.775 158.475 65.945 159.205 ;
        RECT 66.200 159.040 66.370 159.230 ;
        RECT 68.100 159.110 68.360 159.950 ;
        RECT 68.535 159.205 68.790 159.780 ;
        RECT 68.960 159.570 69.290 159.950 ;
        RECT 69.505 159.400 69.675 159.780 ;
        RECT 68.960 159.230 69.675 159.400 ;
        RECT 69.935 159.275 70.195 159.780 ;
        RECT 70.375 159.570 70.705 159.950 ;
        RECT 70.885 159.400 71.055 159.780 ;
        RECT 66.115 158.710 66.370 159.040 ;
        RECT 66.200 158.500 66.370 158.710 ;
        RECT 66.650 158.680 67.005 159.050 ;
        RECT 65.775 157.570 66.030 158.475 ;
        RECT 66.200 158.330 66.915 158.500 ;
        RECT 66.200 157.400 66.530 158.160 ;
        RECT 66.745 157.570 66.915 158.330 ;
        RECT 68.100 157.400 68.360 158.550 ;
        RECT 68.535 158.475 68.705 159.205 ;
        RECT 68.960 159.040 69.130 159.230 ;
        RECT 68.875 158.710 69.130 159.040 ;
        RECT 68.960 158.500 69.130 158.710 ;
        RECT 69.410 158.680 69.765 159.050 ;
        RECT 68.535 157.570 68.790 158.475 ;
        RECT 68.960 158.330 69.675 158.500 ;
        RECT 68.960 157.400 69.290 158.160 ;
        RECT 69.505 157.570 69.675 158.330 ;
        RECT 69.935 158.475 70.105 159.275 ;
        RECT 70.390 159.230 71.055 159.400 ;
        RECT 70.390 158.975 70.560 159.230 ;
        RECT 71.315 159.200 72.525 159.950 ;
        RECT 70.275 158.645 70.560 158.975 ;
        RECT 70.795 158.680 71.125 159.050 ;
        RECT 70.390 158.500 70.560 158.645 ;
        RECT 69.935 157.570 70.205 158.475 ;
        RECT 70.390 158.330 71.055 158.500 ;
        RECT 70.375 157.400 70.705 158.160 ;
        RECT 70.885 157.570 71.055 158.330 ;
        RECT 71.315 158.490 71.835 159.030 ;
        RECT 72.005 158.660 72.525 159.200 ;
        RECT 72.900 159.170 73.400 159.780 ;
        RECT 72.695 158.710 73.045 158.960 ;
        RECT 73.230 158.540 73.400 159.170 ;
        RECT 74.030 159.300 74.360 159.780 ;
        RECT 74.530 159.490 74.755 159.950 ;
        RECT 74.925 159.300 75.255 159.780 ;
        RECT 74.030 159.130 75.255 159.300 ;
        RECT 75.445 159.150 75.695 159.950 ;
        RECT 75.865 159.150 76.205 159.780 ;
        RECT 76.375 159.180 78.045 159.950 ;
        RECT 73.570 158.760 73.900 158.960 ;
        RECT 74.070 158.760 74.400 158.960 ;
        RECT 74.570 158.760 74.990 158.960 ;
        RECT 75.165 158.790 75.860 158.960 ;
        RECT 75.165 158.540 75.335 158.790 ;
        RECT 76.030 158.540 76.205 159.150 ;
        RECT 71.315 157.400 72.525 158.490 ;
        RECT 72.900 158.370 75.335 158.540 ;
        RECT 72.900 157.570 73.230 158.370 ;
        RECT 73.400 157.400 73.730 158.200 ;
        RECT 74.030 157.570 74.360 158.370 ;
        RECT 75.005 157.400 75.255 158.200 ;
        RECT 75.525 157.400 75.695 158.540 ;
        RECT 75.865 157.570 76.205 158.540 ;
        RECT 76.375 158.490 77.125 159.010 ;
        RECT 77.295 158.660 78.045 159.180 ;
        RECT 78.275 159.130 78.485 159.950 ;
        RECT 78.655 159.150 78.985 159.780 ;
        RECT 78.655 158.550 78.905 159.150 ;
        RECT 79.155 159.130 79.385 159.950 ;
        RECT 79.595 159.225 79.885 159.950 ;
        RECT 80.060 159.240 80.315 159.770 ;
        RECT 80.485 159.490 80.790 159.950 ;
        RECT 81.035 159.570 82.105 159.740 ;
        RECT 79.075 158.710 79.405 158.960 ;
        RECT 80.060 158.590 80.270 159.240 ;
        RECT 81.035 159.215 81.355 159.570 ;
        RECT 81.030 159.040 81.355 159.215 ;
        RECT 80.440 158.740 81.355 159.040 ;
        RECT 81.525 159.000 81.765 159.400 ;
        RECT 81.935 159.340 82.105 159.570 ;
        RECT 82.275 159.510 82.465 159.950 ;
        RECT 82.635 159.500 83.585 159.780 ;
        RECT 83.805 159.590 84.155 159.760 ;
        RECT 81.935 159.170 82.465 159.340 ;
        RECT 80.440 158.710 81.180 158.740 ;
        RECT 76.375 157.400 78.045 158.490 ;
        RECT 78.275 157.400 78.485 158.540 ;
        RECT 78.655 157.570 78.985 158.550 ;
        RECT 79.155 157.400 79.385 158.540 ;
        RECT 79.595 157.400 79.885 158.565 ;
        RECT 80.060 157.710 80.315 158.590 ;
        RECT 80.485 157.400 80.790 158.540 ;
        RECT 81.010 158.120 81.180 158.710 ;
        RECT 81.525 158.630 82.065 159.000 ;
        RECT 82.245 158.890 82.465 159.170 ;
        RECT 82.635 158.720 82.805 159.500 ;
        RECT 82.400 158.550 82.805 158.720 ;
        RECT 82.975 158.710 83.325 159.330 ;
        RECT 82.400 158.460 82.570 158.550 ;
        RECT 83.495 158.540 83.705 159.330 ;
        RECT 81.350 158.290 82.570 158.460 ;
        RECT 83.030 158.380 83.705 158.540 ;
        RECT 81.010 157.950 81.810 158.120 ;
        RECT 81.130 157.400 81.460 157.780 ;
        RECT 81.640 157.660 81.810 157.950 ;
        RECT 82.400 157.910 82.570 158.290 ;
        RECT 82.740 158.370 83.705 158.380 ;
        RECT 83.895 159.200 84.155 159.590 ;
        RECT 84.365 159.490 84.695 159.950 ;
        RECT 85.570 159.560 86.425 159.730 ;
        RECT 86.630 159.560 87.125 159.730 ;
        RECT 87.295 159.590 87.625 159.950 ;
        RECT 83.895 158.510 84.065 159.200 ;
        RECT 84.235 158.850 84.405 159.030 ;
        RECT 84.575 159.020 85.365 159.270 ;
        RECT 85.570 158.850 85.740 159.560 ;
        RECT 85.910 159.050 86.265 159.270 ;
        RECT 84.235 158.680 85.925 158.850 ;
        RECT 82.740 158.080 83.200 158.370 ;
        RECT 83.895 158.340 85.395 158.510 ;
        RECT 83.895 158.200 84.065 158.340 ;
        RECT 83.505 158.030 84.065 158.200 ;
        RECT 81.980 157.400 82.230 157.860 ;
        RECT 82.400 157.570 83.270 157.910 ;
        RECT 83.505 157.570 83.675 158.030 ;
        RECT 84.510 158.000 85.585 158.170 ;
        RECT 83.845 157.400 84.215 157.860 ;
        RECT 84.510 157.660 84.680 158.000 ;
        RECT 84.850 157.400 85.180 157.830 ;
        RECT 85.415 157.660 85.585 158.000 ;
        RECT 85.755 157.900 85.925 158.680 ;
        RECT 86.095 158.460 86.265 159.050 ;
        RECT 86.435 158.650 86.785 159.270 ;
        RECT 86.095 158.070 86.560 158.460 ;
        RECT 86.955 158.200 87.125 159.560 ;
        RECT 87.295 158.370 87.755 159.420 ;
        RECT 86.730 158.030 87.125 158.200 ;
        RECT 86.730 157.900 86.900 158.030 ;
        RECT 85.755 157.570 86.435 157.900 ;
        RECT 86.650 157.570 86.900 157.900 ;
        RECT 87.070 157.400 87.320 157.860 ;
        RECT 87.490 157.585 87.815 158.370 ;
        RECT 87.985 157.570 88.155 159.690 ;
        RECT 88.325 159.570 88.655 159.950 ;
        RECT 88.825 159.400 89.080 159.690 ;
        RECT 88.330 159.230 89.080 159.400 ;
        RECT 88.330 158.240 88.560 159.230 ;
        RECT 89.255 159.200 90.465 159.950 ;
        RECT 88.730 158.410 89.080 159.060 ;
        RECT 89.255 158.490 89.775 159.030 ;
        RECT 89.945 158.660 90.465 159.200 ;
        RECT 90.635 159.180 94.145 159.950 ;
        RECT 90.635 158.490 92.325 159.010 ;
        RECT 92.495 158.660 94.145 159.180 ;
        RECT 94.315 159.275 94.585 159.620 ;
        RECT 94.775 159.550 95.155 159.950 ;
        RECT 95.325 159.380 95.495 159.730 ;
        RECT 95.665 159.550 95.995 159.950 ;
        RECT 96.195 159.380 96.365 159.730 ;
        RECT 96.565 159.450 96.895 159.950 ;
        RECT 94.315 158.540 94.485 159.275 ;
        RECT 94.755 159.210 96.365 159.380 ;
        RECT 94.755 159.040 94.925 159.210 ;
        RECT 94.655 158.710 94.925 159.040 ;
        RECT 95.095 158.710 95.500 159.040 ;
        RECT 94.755 158.540 94.925 158.710 ;
        RECT 88.330 158.070 89.080 158.240 ;
        RECT 88.325 157.400 88.655 157.900 ;
        RECT 88.825 157.570 89.080 158.070 ;
        RECT 89.255 157.400 90.465 158.490 ;
        RECT 90.635 157.400 94.145 158.490 ;
        RECT 94.315 157.570 94.585 158.540 ;
        RECT 94.755 158.370 95.480 158.540 ;
        RECT 95.670 158.420 96.380 159.040 ;
        RECT 96.550 158.710 96.900 159.280 ;
        RECT 97.075 159.150 97.415 159.780 ;
        RECT 97.585 159.150 97.835 159.950 ;
        RECT 98.025 159.300 98.355 159.780 ;
        RECT 98.525 159.490 98.750 159.950 ;
        RECT 98.920 159.300 99.250 159.780 ;
        RECT 97.075 159.100 97.305 159.150 ;
        RECT 98.025 159.130 99.250 159.300 ;
        RECT 99.880 159.170 100.380 159.780 ;
        RECT 97.075 158.540 97.250 159.100 ;
        RECT 97.420 158.790 98.115 158.960 ;
        RECT 97.945 158.540 98.115 158.790 ;
        RECT 98.290 158.760 98.710 158.960 ;
        RECT 98.880 158.760 99.210 158.960 ;
        RECT 99.380 158.760 99.710 158.960 ;
        RECT 99.880 158.540 100.050 159.170 ;
        RECT 101.675 159.150 102.015 159.780 ;
        RECT 102.185 159.150 102.435 159.950 ;
        RECT 102.625 159.300 102.955 159.780 ;
        RECT 103.125 159.490 103.350 159.950 ;
        RECT 103.520 159.300 103.850 159.780 ;
        RECT 100.235 158.710 100.585 158.960 ;
        RECT 101.675 158.540 101.850 159.150 ;
        RECT 102.625 159.130 103.850 159.300 ;
        RECT 104.480 159.170 104.980 159.780 ;
        RECT 105.355 159.225 105.645 159.950 ;
        RECT 105.815 159.200 107.025 159.950 ;
        RECT 102.020 158.790 102.715 158.960 ;
        RECT 102.545 158.540 102.715 158.790 ;
        RECT 102.890 158.760 103.310 158.960 ;
        RECT 103.480 158.760 103.810 158.960 ;
        RECT 103.980 158.760 104.310 158.960 ;
        RECT 104.480 158.540 104.650 159.170 ;
        RECT 104.835 158.710 105.185 158.960 ;
        RECT 95.310 158.250 95.480 158.370 ;
        RECT 96.580 158.250 96.900 158.540 ;
        RECT 94.795 157.400 95.075 158.200 ;
        RECT 95.310 158.080 96.900 158.250 ;
        RECT 95.245 157.620 96.900 157.910 ;
        RECT 97.075 157.570 97.415 158.540 ;
        RECT 97.585 157.400 97.755 158.540 ;
        RECT 97.945 158.370 100.380 158.540 ;
        RECT 98.025 157.400 98.275 158.200 ;
        RECT 98.920 157.570 99.250 158.370 ;
        RECT 99.550 157.400 99.880 158.200 ;
        RECT 100.050 157.570 100.380 158.370 ;
        RECT 101.675 157.570 102.015 158.540 ;
        RECT 102.185 157.400 102.355 158.540 ;
        RECT 102.545 158.370 104.980 158.540 ;
        RECT 102.625 157.400 102.875 158.200 ;
        RECT 103.520 157.570 103.850 158.370 ;
        RECT 104.150 157.400 104.480 158.200 ;
        RECT 104.650 157.570 104.980 158.370 ;
        RECT 105.355 157.400 105.645 158.565 ;
        RECT 105.815 158.490 106.335 159.030 ;
        RECT 106.505 158.660 107.025 159.200 ;
        RECT 107.570 159.240 107.825 159.770 ;
        RECT 108.005 159.490 108.290 159.950 ;
        RECT 105.815 157.400 107.025 158.490 ;
        RECT 107.570 158.380 107.750 159.240 ;
        RECT 108.470 159.040 108.720 159.690 ;
        RECT 107.920 158.710 108.720 159.040 ;
        RECT 107.570 157.910 107.825 158.380 ;
        RECT 107.485 157.740 107.825 157.910 ;
        RECT 107.570 157.710 107.825 157.740 ;
        RECT 108.005 157.400 108.290 158.200 ;
        RECT 108.470 158.120 108.720 158.710 ;
        RECT 108.920 159.355 109.240 159.685 ;
        RECT 109.420 159.470 110.080 159.950 ;
        RECT 110.280 159.560 111.130 159.730 ;
        RECT 108.920 158.460 109.110 159.355 ;
        RECT 109.430 159.030 110.090 159.300 ;
        RECT 109.760 158.970 110.090 159.030 ;
        RECT 109.280 158.800 109.610 158.860 ;
        RECT 110.280 158.800 110.450 159.560 ;
        RECT 111.690 159.490 112.010 159.950 ;
        RECT 112.210 159.310 112.460 159.740 ;
        RECT 112.750 159.510 113.160 159.950 ;
        RECT 113.330 159.570 114.345 159.770 ;
        RECT 110.620 159.140 111.870 159.310 ;
        RECT 110.620 159.020 110.950 159.140 ;
        RECT 109.280 158.630 111.180 158.800 ;
        RECT 108.920 158.290 110.840 158.460 ;
        RECT 108.920 158.270 109.240 158.290 ;
        RECT 108.470 157.610 108.800 158.120 ;
        RECT 109.070 157.660 109.240 158.270 ;
        RECT 111.010 158.120 111.180 158.630 ;
        RECT 111.350 158.560 111.530 158.970 ;
        RECT 111.700 158.380 111.870 159.140 ;
        RECT 109.410 157.400 109.740 158.090 ;
        RECT 109.970 157.950 111.180 158.120 ;
        RECT 111.350 158.070 111.870 158.380 ;
        RECT 112.040 158.970 112.460 159.310 ;
        RECT 112.750 158.970 113.160 159.300 ;
        RECT 112.040 158.200 112.230 158.970 ;
        RECT 113.330 158.840 113.500 159.570 ;
        RECT 114.645 159.400 114.815 159.730 ;
        RECT 114.985 159.570 115.315 159.950 ;
        RECT 113.670 159.020 114.020 159.390 ;
        RECT 113.330 158.800 113.750 158.840 ;
        RECT 112.400 158.630 113.750 158.800 ;
        RECT 112.400 158.470 112.650 158.630 ;
        RECT 113.160 158.200 113.410 158.460 ;
        RECT 112.040 157.950 113.410 158.200 ;
        RECT 109.970 157.660 110.210 157.950 ;
        RECT 111.010 157.870 111.180 157.950 ;
        RECT 110.410 157.400 110.830 157.780 ;
        RECT 111.010 157.620 111.640 157.870 ;
        RECT 112.110 157.400 112.440 157.780 ;
        RECT 112.610 157.660 112.780 157.950 ;
        RECT 113.580 157.785 113.750 158.630 ;
        RECT 114.200 158.460 114.420 159.330 ;
        RECT 114.645 159.210 115.340 159.400 ;
        RECT 113.920 158.080 114.420 158.460 ;
        RECT 114.590 158.410 115.000 159.030 ;
        RECT 115.170 158.240 115.340 159.210 ;
        RECT 114.645 158.070 115.340 158.240 ;
        RECT 112.960 157.400 113.340 157.780 ;
        RECT 113.580 157.615 114.410 157.785 ;
        RECT 114.645 157.570 114.815 158.070 ;
        RECT 114.985 157.400 115.315 157.900 ;
        RECT 115.530 157.570 115.755 159.690 ;
        RECT 115.925 159.570 116.255 159.950 ;
        RECT 116.425 159.400 116.595 159.690 ;
        RECT 115.930 159.230 116.595 159.400 ;
        RECT 115.930 158.240 116.160 159.230 ;
        RECT 117.315 159.200 118.525 159.950 ;
        RECT 116.330 158.410 116.680 159.060 ;
        RECT 117.315 158.490 117.835 159.030 ;
        RECT 118.005 158.660 118.525 159.200 ;
        RECT 115.930 158.070 116.595 158.240 ;
        RECT 115.925 157.400 116.255 157.900 ;
        RECT 116.425 157.570 116.595 158.070 ;
        RECT 117.315 157.400 118.525 158.490 ;
        RECT 11.430 157.230 118.610 157.400 ;
        RECT 11.515 156.140 12.725 157.230 ;
        RECT 11.515 155.430 12.035 155.970 ;
        RECT 12.205 155.600 12.725 156.140 ;
        RECT 13.355 156.140 15.025 157.230 ;
        RECT 13.355 155.620 14.105 156.140 ;
        RECT 15.195 156.065 15.485 157.230 ;
        RECT 15.655 156.140 17.325 157.230 ;
        RECT 14.275 155.450 15.025 155.970 ;
        RECT 15.655 155.620 16.405 156.140 ;
        RECT 17.555 156.090 17.765 157.230 ;
        RECT 17.935 156.080 18.265 157.060 ;
        RECT 18.435 156.090 18.665 157.230 ;
        RECT 18.875 156.140 22.385 157.230 ;
        RECT 22.555 156.155 22.825 157.060 ;
        RECT 22.995 156.470 23.325 157.230 ;
        RECT 23.505 156.300 23.675 157.060 ;
        RECT 16.575 155.450 17.325 155.970 ;
        RECT 11.515 154.680 12.725 155.430 ;
        RECT 13.355 154.680 15.025 155.450 ;
        RECT 15.195 154.680 15.485 155.405 ;
        RECT 15.655 154.680 17.325 155.450 ;
        RECT 17.555 154.680 17.765 155.500 ;
        RECT 17.935 155.480 18.185 156.080 ;
        RECT 18.355 155.670 18.685 155.920 ;
        RECT 18.875 155.620 20.565 156.140 ;
        RECT 17.935 154.850 18.265 155.480 ;
        RECT 18.435 154.680 18.665 155.500 ;
        RECT 20.735 155.450 22.385 155.970 ;
        RECT 18.875 154.680 22.385 155.450 ;
        RECT 22.555 155.355 22.725 156.155 ;
        RECT 23.010 156.130 23.675 156.300 ;
        RECT 23.935 156.140 25.145 157.230 ;
        RECT 23.010 155.985 23.180 156.130 ;
        RECT 22.895 155.655 23.180 155.985 ;
        RECT 23.010 155.400 23.180 155.655 ;
        RECT 23.415 155.580 23.745 155.950 ;
        RECT 23.935 155.600 24.455 156.140 ;
        RECT 25.355 156.090 25.585 157.230 ;
        RECT 25.755 156.080 26.085 157.060 ;
        RECT 26.255 156.090 26.465 157.230 ;
        RECT 24.625 155.430 25.145 155.970 ;
        RECT 25.335 155.670 25.665 155.920 ;
        RECT 22.555 154.850 22.815 155.355 ;
        RECT 23.010 155.230 23.675 155.400 ;
        RECT 22.995 154.680 23.325 155.060 ;
        RECT 23.505 154.850 23.675 155.230 ;
        RECT 23.935 154.680 25.145 155.430 ;
        RECT 25.355 154.680 25.585 155.500 ;
        RECT 25.835 155.480 26.085 156.080 ;
        RECT 26.700 156.040 26.955 156.920 ;
        RECT 27.125 156.090 27.430 157.230 ;
        RECT 27.770 156.850 28.100 157.230 ;
        RECT 28.280 156.680 28.450 156.970 ;
        RECT 28.620 156.770 28.870 157.230 ;
        RECT 27.650 156.510 28.450 156.680 ;
        RECT 29.040 156.720 29.910 157.060 ;
        RECT 25.755 154.850 26.085 155.480 ;
        RECT 26.255 154.680 26.465 155.500 ;
        RECT 26.700 155.390 26.910 156.040 ;
        RECT 27.650 155.920 27.820 156.510 ;
        RECT 29.040 156.340 29.210 156.720 ;
        RECT 30.145 156.600 30.315 157.060 ;
        RECT 30.485 156.770 30.855 157.230 ;
        RECT 31.150 156.630 31.320 156.970 ;
        RECT 31.490 156.800 31.820 157.230 ;
        RECT 32.055 156.630 32.225 156.970 ;
        RECT 27.990 156.170 29.210 156.340 ;
        RECT 29.380 156.260 29.840 156.550 ;
        RECT 30.145 156.430 30.705 156.600 ;
        RECT 31.150 156.460 32.225 156.630 ;
        RECT 32.395 156.730 33.075 157.060 ;
        RECT 33.290 156.730 33.540 157.060 ;
        RECT 33.710 156.770 33.960 157.230 ;
        RECT 30.535 156.290 30.705 156.430 ;
        RECT 29.380 156.250 30.345 156.260 ;
        RECT 29.040 156.080 29.210 156.170 ;
        RECT 29.670 156.090 30.345 156.250 ;
        RECT 27.080 155.890 27.820 155.920 ;
        RECT 27.080 155.590 27.995 155.890 ;
        RECT 27.670 155.415 27.995 155.590 ;
        RECT 26.700 154.860 26.955 155.390 ;
        RECT 27.125 154.680 27.430 155.140 ;
        RECT 27.675 155.060 27.995 155.415 ;
        RECT 28.165 155.630 28.705 156.000 ;
        RECT 29.040 155.910 29.445 156.080 ;
        RECT 28.165 155.230 28.405 155.630 ;
        RECT 28.885 155.460 29.105 155.740 ;
        RECT 28.575 155.290 29.105 155.460 ;
        RECT 28.575 155.060 28.745 155.290 ;
        RECT 29.275 155.130 29.445 155.910 ;
        RECT 29.615 155.300 29.965 155.920 ;
        RECT 30.135 155.300 30.345 156.090 ;
        RECT 30.535 156.120 32.035 156.290 ;
        RECT 30.535 155.430 30.705 156.120 ;
        RECT 32.395 155.950 32.565 156.730 ;
        RECT 33.370 156.600 33.540 156.730 ;
        RECT 30.875 155.780 32.565 155.950 ;
        RECT 32.735 156.170 33.200 156.560 ;
        RECT 33.370 156.430 33.765 156.600 ;
        RECT 30.875 155.600 31.045 155.780 ;
        RECT 27.675 154.890 28.745 155.060 ;
        RECT 28.915 154.680 29.105 155.120 ;
        RECT 29.275 154.850 30.225 155.130 ;
        RECT 30.535 155.040 30.795 155.430 ;
        RECT 31.215 155.360 32.005 155.610 ;
        RECT 30.445 154.870 30.795 155.040 ;
        RECT 31.005 154.680 31.335 155.140 ;
        RECT 32.210 155.070 32.380 155.780 ;
        RECT 32.735 155.580 32.905 156.170 ;
        RECT 32.550 155.360 32.905 155.580 ;
        RECT 33.075 155.360 33.425 155.980 ;
        RECT 33.595 155.070 33.765 156.430 ;
        RECT 34.130 156.260 34.455 157.045 ;
        RECT 33.935 155.210 34.395 156.260 ;
        RECT 32.210 154.900 33.065 155.070 ;
        RECT 33.270 154.900 33.765 155.070 ;
        RECT 33.935 154.680 34.265 155.040 ;
        RECT 34.625 154.940 34.795 157.060 ;
        RECT 34.965 156.730 35.295 157.230 ;
        RECT 35.465 156.560 35.720 157.060 ;
        RECT 34.970 156.390 35.720 156.560 ;
        RECT 34.970 155.400 35.200 156.390 ;
        RECT 35.370 155.570 35.720 156.220 ;
        RECT 35.895 156.140 37.105 157.230 ;
        RECT 37.275 156.140 40.785 157.230 ;
        RECT 35.895 155.600 36.415 156.140 ;
        RECT 36.585 155.430 37.105 155.970 ;
        RECT 37.275 155.620 38.965 156.140 ;
        RECT 40.955 156.065 41.245 157.230 ;
        RECT 41.875 156.140 44.465 157.230 ;
        RECT 39.135 155.450 40.785 155.970 ;
        RECT 41.875 155.620 43.085 156.140 ;
        RECT 44.635 156.090 44.905 157.060 ;
        RECT 45.115 156.430 45.395 157.230 ;
        RECT 45.565 156.720 47.220 157.010 ;
        RECT 45.630 156.380 47.220 156.550 ;
        RECT 45.630 156.260 45.800 156.380 ;
        RECT 45.075 156.090 45.800 156.260 ;
        RECT 43.255 155.450 44.465 155.970 ;
        RECT 34.970 155.230 35.720 155.400 ;
        RECT 34.965 154.680 35.295 155.060 ;
        RECT 35.465 154.940 35.720 155.230 ;
        RECT 35.895 154.680 37.105 155.430 ;
        RECT 37.275 154.680 40.785 155.450 ;
        RECT 40.955 154.680 41.245 155.405 ;
        RECT 41.875 154.680 44.465 155.450 ;
        RECT 44.635 155.355 44.805 156.090 ;
        RECT 45.075 155.920 45.245 156.090 ;
        RECT 45.990 156.040 46.705 156.210 ;
        RECT 46.900 156.090 47.220 156.380 ;
        RECT 47.915 156.090 48.125 157.230 ;
        RECT 48.295 156.080 48.625 157.060 ;
        RECT 48.795 156.090 49.025 157.230 ;
        RECT 49.235 156.470 49.750 156.880 ;
        RECT 49.985 156.470 50.155 157.230 ;
        RECT 50.325 156.890 52.355 157.060 ;
        RECT 44.975 155.590 45.245 155.920 ;
        RECT 45.415 155.590 45.820 155.920 ;
        RECT 45.990 155.590 46.700 156.040 ;
        RECT 45.075 155.420 45.245 155.590 ;
        RECT 44.635 155.010 44.905 155.355 ;
        RECT 45.075 155.250 46.685 155.420 ;
        RECT 46.870 155.350 47.220 155.920 ;
        RECT 45.095 154.680 45.475 155.080 ;
        RECT 45.645 154.900 45.815 155.250 ;
        RECT 45.985 154.680 46.315 155.080 ;
        RECT 46.515 154.900 46.685 155.250 ;
        RECT 46.885 154.680 47.215 155.180 ;
        RECT 47.915 154.680 48.125 155.500 ;
        RECT 48.295 155.480 48.545 156.080 ;
        RECT 48.715 155.670 49.045 155.920 ;
        RECT 49.235 155.660 49.575 156.470 ;
        RECT 50.325 156.225 50.495 156.890 ;
        RECT 50.890 156.550 52.015 156.720 ;
        RECT 49.745 156.035 50.495 156.225 ;
        RECT 50.665 156.210 51.675 156.380 ;
        RECT 48.295 154.850 48.625 155.480 ;
        RECT 48.795 154.680 49.025 155.500 ;
        RECT 49.235 155.490 50.465 155.660 ;
        RECT 49.510 154.885 49.755 155.490 ;
        RECT 49.975 154.680 50.485 155.215 ;
        RECT 50.665 154.850 50.855 156.210 ;
        RECT 51.025 155.870 51.300 156.010 ;
        RECT 51.025 155.700 51.305 155.870 ;
        RECT 51.025 154.850 51.300 155.700 ;
        RECT 51.505 155.410 51.675 156.210 ;
        RECT 51.845 155.420 52.015 156.550 ;
        RECT 52.185 155.920 52.355 156.890 ;
        RECT 52.525 156.090 52.695 157.230 ;
        RECT 52.865 156.090 53.200 157.060 ;
        RECT 52.185 155.590 52.380 155.920 ;
        RECT 52.605 155.590 52.860 155.920 ;
        RECT 52.605 155.420 52.775 155.590 ;
        RECT 53.030 155.420 53.200 156.090 ;
        RECT 51.845 155.250 52.775 155.420 ;
        RECT 51.845 155.215 52.020 155.250 ;
        RECT 51.490 154.850 52.020 155.215 ;
        RECT 52.445 154.680 52.775 155.080 ;
        RECT 52.945 154.850 53.200 155.420 ;
        RECT 53.375 156.090 53.715 157.060 ;
        RECT 53.885 156.090 54.055 157.230 ;
        RECT 54.325 156.430 54.575 157.230 ;
        RECT 55.220 156.260 55.550 157.060 ;
        RECT 55.850 156.430 56.180 157.230 ;
        RECT 56.350 156.260 56.680 157.060 ;
        RECT 57.430 156.890 57.685 156.920 ;
        RECT 57.345 156.720 57.685 156.890 ;
        RECT 54.245 156.090 56.680 156.260 ;
        RECT 57.430 156.250 57.685 156.720 ;
        RECT 57.865 156.430 58.150 157.230 ;
        RECT 58.330 156.510 58.660 157.020 ;
        RECT 53.375 155.530 53.550 156.090 ;
        RECT 54.245 155.840 54.415 156.090 ;
        RECT 53.720 155.670 54.415 155.840 ;
        RECT 54.590 155.670 55.010 155.870 ;
        RECT 55.180 155.670 55.510 155.870 ;
        RECT 55.680 155.670 56.010 155.870 ;
        RECT 53.375 155.480 53.605 155.530 ;
        RECT 53.375 154.850 53.715 155.480 ;
        RECT 53.885 154.680 54.135 155.480 ;
        RECT 54.325 155.330 55.550 155.500 ;
        RECT 54.325 154.850 54.655 155.330 ;
        RECT 54.825 154.680 55.050 155.140 ;
        RECT 55.220 154.850 55.550 155.330 ;
        RECT 56.180 155.460 56.350 156.090 ;
        RECT 56.535 155.670 56.885 155.920 ;
        RECT 56.180 154.850 56.680 155.460 ;
        RECT 57.430 155.390 57.610 156.250 ;
        RECT 58.330 155.920 58.580 156.510 ;
        RECT 58.930 156.360 59.100 156.970 ;
        RECT 59.270 156.540 59.600 157.230 ;
        RECT 59.830 156.680 60.070 156.970 ;
        RECT 60.270 156.850 60.690 157.230 ;
        RECT 60.870 156.760 61.500 157.010 ;
        RECT 61.970 156.850 62.300 157.230 ;
        RECT 60.870 156.680 61.040 156.760 ;
        RECT 62.470 156.680 62.640 156.970 ;
        RECT 62.820 156.850 63.200 157.230 ;
        RECT 63.440 156.845 64.270 157.015 ;
        RECT 59.830 156.510 61.040 156.680 ;
        RECT 57.780 155.590 58.580 155.920 ;
        RECT 57.430 154.860 57.685 155.390 ;
        RECT 57.865 154.680 58.150 155.140 ;
        RECT 58.330 154.940 58.580 155.590 ;
        RECT 58.780 156.340 59.100 156.360 ;
        RECT 58.780 156.170 60.700 156.340 ;
        RECT 58.780 155.275 58.970 156.170 ;
        RECT 60.870 156.000 61.040 156.510 ;
        RECT 61.210 156.250 61.730 156.560 ;
        RECT 59.140 155.830 61.040 156.000 ;
        RECT 59.140 155.770 59.470 155.830 ;
        RECT 59.620 155.600 59.950 155.660 ;
        RECT 59.290 155.330 59.950 155.600 ;
        RECT 58.780 154.945 59.100 155.275 ;
        RECT 59.280 154.680 59.940 155.160 ;
        RECT 60.140 155.070 60.310 155.830 ;
        RECT 61.210 155.660 61.390 156.070 ;
        RECT 60.480 155.490 60.810 155.610 ;
        RECT 61.560 155.490 61.730 156.250 ;
        RECT 60.480 155.320 61.730 155.490 ;
        RECT 61.900 156.430 63.270 156.680 ;
        RECT 61.900 155.660 62.090 156.430 ;
        RECT 63.020 156.170 63.270 156.430 ;
        RECT 62.260 156.000 62.510 156.160 ;
        RECT 63.440 156.000 63.610 156.845 ;
        RECT 64.505 156.560 64.675 157.060 ;
        RECT 64.845 156.730 65.175 157.230 ;
        RECT 63.780 156.170 64.280 156.550 ;
        RECT 64.505 156.390 65.200 156.560 ;
        RECT 62.260 155.830 63.610 156.000 ;
        RECT 63.190 155.790 63.610 155.830 ;
        RECT 61.900 155.320 62.320 155.660 ;
        RECT 62.610 155.330 63.020 155.660 ;
        RECT 60.140 154.900 60.990 155.070 ;
        RECT 61.550 154.680 61.870 155.140 ;
        RECT 62.070 154.890 62.320 155.320 ;
        RECT 62.610 154.680 63.020 155.120 ;
        RECT 63.190 155.060 63.360 155.790 ;
        RECT 63.530 155.240 63.880 155.610 ;
        RECT 64.060 155.300 64.280 156.170 ;
        RECT 64.450 155.600 64.860 156.220 ;
        RECT 65.030 155.420 65.200 156.390 ;
        RECT 64.505 155.230 65.200 155.420 ;
        RECT 63.190 154.860 64.205 155.060 ;
        RECT 64.505 154.900 64.675 155.230 ;
        RECT 64.845 154.680 65.175 155.060 ;
        RECT 65.390 154.940 65.615 157.060 ;
        RECT 65.785 156.730 66.115 157.230 ;
        RECT 66.285 156.560 66.455 157.060 ;
        RECT 65.790 156.390 66.455 156.560 ;
        RECT 65.790 155.400 66.020 156.390 ;
        RECT 66.190 155.570 66.540 156.220 ;
        RECT 66.715 156.065 67.005 157.230 ;
        RECT 67.185 156.170 67.515 157.230 ;
        RECT 67.695 155.920 67.865 156.890 ;
        RECT 68.035 156.640 68.365 157.040 ;
        RECT 68.535 156.870 68.865 157.230 ;
        RECT 69.065 156.640 69.765 157.060 ;
        RECT 68.035 156.410 69.765 156.640 ;
        RECT 68.035 156.190 68.365 156.410 ;
        RECT 68.560 155.920 68.885 156.210 ;
        RECT 67.175 155.590 67.485 155.920 ;
        RECT 67.695 155.590 68.070 155.920 ;
        RECT 68.390 155.590 68.885 155.920 ;
        RECT 69.060 155.670 69.390 156.210 ;
        RECT 69.560 155.440 69.765 156.410 ;
        RECT 65.790 155.230 66.455 155.400 ;
        RECT 65.785 154.680 66.115 155.060 ;
        RECT 66.285 154.940 66.455 155.230 ;
        RECT 66.715 154.680 67.005 155.405 ;
        RECT 67.185 155.210 68.545 155.420 ;
        RECT 67.185 154.850 67.515 155.210 ;
        RECT 67.685 154.680 68.015 155.040 ;
        RECT 68.215 154.850 68.545 155.210 ;
        RECT 69.055 154.850 69.765 155.440 ;
        RECT 69.935 156.260 70.245 157.060 ;
        RECT 70.415 156.430 70.725 157.230 ;
        RECT 70.895 156.600 71.155 157.060 ;
        RECT 71.325 156.770 71.580 157.230 ;
        RECT 71.755 156.600 72.015 157.060 ;
        RECT 70.895 156.430 72.015 156.600 ;
        RECT 69.935 156.090 70.965 156.260 ;
        RECT 69.935 155.180 70.105 156.090 ;
        RECT 70.275 155.350 70.625 155.920 ;
        RECT 70.795 155.840 70.965 156.090 ;
        RECT 71.755 156.180 72.015 156.430 ;
        RECT 72.185 156.360 72.470 157.230 ;
        RECT 72.900 156.260 73.230 157.060 ;
        RECT 73.400 156.430 73.730 157.230 ;
        RECT 74.030 156.260 74.360 157.060 ;
        RECT 75.005 156.430 75.255 157.230 ;
        RECT 71.755 156.010 72.510 156.180 ;
        RECT 72.900 156.090 75.335 156.260 ;
        RECT 75.525 156.090 75.695 157.230 ;
        RECT 75.865 156.090 76.205 157.060 ;
        RECT 70.795 155.670 71.935 155.840 ;
        RECT 72.105 155.500 72.510 156.010 ;
        RECT 72.695 155.670 73.045 155.920 ;
        RECT 70.860 155.330 72.510 155.500 ;
        RECT 73.230 155.460 73.400 156.090 ;
        RECT 73.570 155.670 73.900 155.870 ;
        RECT 74.070 155.670 74.400 155.870 ;
        RECT 74.570 155.700 74.995 155.870 ;
        RECT 75.165 155.840 75.335 156.090 ;
        RECT 74.570 155.670 74.990 155.700 ;
        RECT 75.165 155.670 75.860 155.840 ;
        RECT 69.935 154.850 70.235 155.180 ;
        RECT 70.405 154.680 70.680 155.160 ;
        RECT 70.860 154.940 71.155 155.330 ;
        RECT 71.325 154.680 71.580 155.160 ;
        RECT 71.755 154.940 72.015 155.330 ;
        RECT 72.185 154.680 72.465 155.160 ;
        RECT 72.900 154.850 73.400 155.460 ;
        RECT 74.030 155.330 75.255 155.500 ;
        RECT 76.030 155.480 76.205 156.090 ;
        RECT 76.835 156.140 80.345 157.230 ;
        RECT 80.515 156.470 81.030 156.880 ;
        RECT 81.265 156.470 81.435 157.230 ;
        RECT 81.605 156.890 83.635 157.060 ;
        RECT 76.835 155.620 78.525 156.140 ;
        RECT 74.030 154.850 74.360 155.330 ;
        RECT 74.530 154.680 74.755 155.140 ;
        RECT 74.925 154.850 75.255 155.330 ;
        RECT 75.445 154.680 75.695 155.480 ;
        RECT 75.865 154.850 76.205 155.480 ;
        RECT 78.695 155.450 80.345 155.970 ;
        RECT 80.515 155.660 80.855 156.470 ;
        RECT 81.605 156.225 81.775 156.890 ;
        RECT 82.170 156.550 83.295 156.720 ;
        RECT 81.025 156.035 81.775 156.225 ;
        RECT 81.945 156.210 82.955 156.380 ;
        RECT 80.515 155.490 81.745 155.660 ;
        RECT 76.835 154.680 80.345 155.450 ;
        RECT 80.790 154.885 81.035 155.490 ;
        RECT 81.255 154.680 81.765 155.215 ;
        RECT 81.945 154.850 82.135 156.210 ;
        RECT 82.305 155.190 82.580 156.010 ;
        RECT 82.785 155.410 82.955 156.210 ;
        RECT 83.125 155.420 83.295 156.550 ;
        RECT 83.465 155.920 83.635 156.890 ;
        RECT 83.805 156.090 83.975 157.230 ;
        RECT 84.145 156.090 84.480 157.060 ;
        RECT 83.465 155.590 83.660 155.920 ;
        RECT 83.885 155.590 84.140 155.920 ;
        RECT 83.885 155.420 84.055 155.590 ;
        RECT 84.310 155.420 84.480 156.090 ;
        RECT 85.115 156.140 86.785 157.230 ;
        RECT 86.960 156.795 92.305 157.230 ;
        RECT 85.115 155.620 85.865 156.140 ;
        RECT 86.035 155.450 86.785 155.970 ;
        RECT 88.550 155.545 88.900 156.795 ;
        RECT 92.475 156.065 92.765 157.230 ;
        RECT 92.935 156.140 96.445 157.230 ;
        RECT 83.125 155.250 84.055 155.420 ;
        RECT 83.125 155.215 83.300 155.250 ;
        RECT 82.305 155.020 82.585 155.190 ;
        RECT 82.305 154.850 82.580 155.020 ;
        RECT 82.770 154.850 83.300 155.215 ;
        RECT 83.725 154.680 84.055 155.080 ;
        RECT 84.225 154.850 84.480 155.420 ;
        RECT 85.115 154.680 86.785 155.450 ;
        RECT 90.380 155.225 90.720 156.055 ;
        RECT 92.935 155.620 94.625 156.140 ;
        RECT 96.615 156.090 96.885 157.060 ;
        RECT 97.095 156.430 97.375 157.230 ;
        RECT 97.545 156.720 99.200 157.010 ;
        RECT 97.610 156.380 99.200 156.550 ;
        RECT 97.610 156.260 97.780 156.380 ;
        RECT 97.055 156.090 97.780 156.260 ;
        RECT 94.795 155.450 96.445 155.970 ;
        RECT 86.960 154.680 92.305 155.225 ;
        RECT 92.475 154.680 92.765 155.405 ;
        RECT 92.935 154.680 96.445 155.450 ;
        RECT 96.615 155.355 96.785 156.090 ;
        RECT 97.055 155.920 97.225 156.090 ;
        RECT 96.955 155.590 97.225 155.920 ;
        RECT 97.395 155.590 97.800 155.920 ;
        RECT 97.970 155.590 98.680 156.210 ;
        RECT 98.880 156.090 99.200 156.380 ;
        RECT 99.375 156.140 101.045 157.230 ;
        RECT 97.055 155.420 97.225 155.590 ;
        RECT 96.615 155.010 96.885 155.355 ;
        RECT 97.055 155.250 98.665 155.420 ;
        RECT 98.850 155.350 99.200 155.920 ;
        RECT 99.375 155.620 100.125 156.140 ;
        RECT 101.215 156.090 101.555 157.060 ;
        RECT 101.725 156.090 101.895 157.230 ;
        RECT 102.165 156.430 102.415 157.230 ;
        RECT 103.060 156.260 103.390 157.060 ;
        RECT 103.690 156.430 104.020 157.230 ;
        RECT 104.190 156.260 104.520 157.060 ;
        RECT 102.085 156.090 104.520 156.260 ;
        RECT 105.355 156.140 107.025 157.230 ;
        RECT 107.195 156.470 107.710 156.880 ;
        RECT 107.945 156.470 108.115 157.230 ;
        RECT 108.285 156.890 110.315 157.060 ;
        RECT 100.295 155.450 101.045 155.970 ;
        RECT 97.075 154.680 97.455 155.080 ;
        RECT 97.625 154.900 97.795 155.250 ;
        RECT 97.965 154.680 98.295 155.080 ;
        RECT 98.495 154.900 98.665 155.250 ;
        RECT 98.865 154.680 99.195 155.180 ;
        RECT 99.375 154.680 101.045 155.450 ;
        RECT 101.215 155.480 101.390 156.090 ;
        RECT 102.085 155.840 102.255 156.090 ;
        RECT 101.560 155.670 102.255 155.840 ;
        RECT 102.430 155.670 102.850 155.870 ;
        RECT 103.020 155.670 103.350 155.870 ;
        RECT 103.520 155.670 103.850 155.870 ;
        RECT 101.215 154.850 101.555 155.480 ;
        RECT 101.725 154.680 101.975 155.480 ;
        RECT 102.165 155.330 103.390 155.500 ;
        RECT 102.165 154.850 102.495 155.330 ;
        RECT 102.665 154.680 102.890 155.140 ;
        RECT 103.060 154.850 103.390 155.330 ;
        RECT 104.020 155.460 104.190 156.090 ;
        RECT 104.375 155.670 104.725 155.920 ;
        RECT 105.355 155.620 106.105 156.140 ;
        RECT 104.020 154.850 104.520 155.460 ;
        RECT 106.275 155.450 107.025 155.970 ;
        RECT 107.195 155.660 107.535 156.470 ;
        RECT 108.285 156.225 108.455 156.890 ;
        RECT 108.850 156.550 109.975 156.720 ;
        RECT 107.705 156.035 108.455 156.225 ;
        RECT 108.625 156.210 109.635 156.380 ;
        RECT 107.195 155.490 108.425 155.660 ;
        RECT 105.355 154.680 107.025 155.450 ;
        RECT 107.470 154.885 107.715 155.490 ;
        RECT 107.935 154.680 108.445 155.215 ;
        RECT 108.625 154.850 108.815 156.210 ;
        RECT 108.985 155.870 109.260 156.010 ;
        RECT 108.985 155.700 109.265 155.870 ;
        RECT 108.985 154.850 109.260 155.700 ;
        RECT 109.465 155.410 109.635 156.210 ;
        RECT 109.805 155.420 109.975 156.550 ;
        RECT 110.145 155.920 110.315 156.890 ;
        RECT 110.485 156.090 110.655 157.230 ;
        RECT 110.825 156.090 111.160 157.060 ;
        RECT 111.800 156.795 117.145 157.230 ;
        RECT 110.145 155.590 110.340 155.920 ;
        RECT 110.565 155.590 110.820 155.920 ;
        RECT 110.565 155.420 110.735 155.590 ;
        RECT 110.990 155.420 111.160 156.090 ;
        RECT 113.390 155.545 113.740 156.795 ;
        RECT 117.315 156.140 118.525 157.230 ;
        RECT 109.805 155.250 110.735 155.420 ;
        RECT 109.805 155.215 109.980 155.250 ;
        RECT 109.450 154.850 109.980 155.215 ;
        RECT 110.405 154.680 110.735 155.080 ;
        RECT 110.905 154.850 111.160 155.420 ;
        RECT 115.220 155.225 115.560 156.055 ;
        RECT 117.315 155.600 117.835 156.140 ;
        RECT 118.005 155.430 118.525 155.970 ;
        RECT 111.800 154.680 117.145 155.225 ;
        RECT 117.315 154.680 118.525 155.430 ;
        RECT 11.430 154.510 118.610 154.680 ;
        RECT 11.515 153.760 12.725 154.510 ;
        RECT 13.360 153.800 13.615 154.330 ;
        RECT 13.785 154.050 14.090 154.510 ;
        RECT 14.335 154.130 15.405 154.300 ;
        RECT 11.515 153.220 12.035 153.760 ;
        RECT 12.205 153.050 12.725 153.590 ;
        RECT 11.515 151.960 12.725 153.050 ;
        RECT 13.360 153.150 13.570 153.800 ;
        RECT 14.335 153.775 14.655 154.130 ;
        RECT 14.330 153.600 14.655 153.775 ;
        RECT 13.740 153.300 14.655 153.600 ;
        RECT 14.825 153.560 15.065 153.960 ;
        RECT 15.235 153.900 15.405 154.130 ;
        RECT 15.575 154.070 15.765 154.510 ;
        RECT 15.935 154.060 16.885 154.340 ;
        RECT 17.105 154.150 17.455 154.320 ;
        RECT 15.235 153.730 15.765 153.900 ;
        RECT 13.740 153.270 14.480 153.300 ;
        RECT 13.360 152.270 13.615 153.150 ;
        RECT 13.785 151.960 14.090 153.100 ;
        RECT 14.310 152.680 14.480 153.270 ;
        RECT 14.825 153.190 15.365 153.560 ;
        RECT 15.545 153.450 15.765 153.730 ;
        RECT 15.935 153.280 16.105 154.060 ;
        RECT 15.700 153.110 16.105 153.280 ;
        RECT 16.275 153.270 16.625 153.890 ;
        RECT 15.700 153.020 15.870 153.110 ;
        RECT 16.795 153.100 17.005 153.890 ;
        RECT 14.650 152.850 15.870 153.020 ;
        RECT 16.330 152.940 17.005 153.100 ;
        RECT 14.310 152.510 15.110 152.680 ;
        RECT 14.430 151.960 14.760 152.340 ;
        RECT 14.940 152.220 15.110 152.510 ;
        RECT 15.700 152.470 15.870 152.850 ;
        RECT 16.040 152.930 17.005 152.940 ;
        RECT 17.195 153.760 17.455 154.150 ;
        RECT 17.665 154.050 17.995 154.510 ;
        RECT 18.870 154.120 19.725 154.290 ;
        RECT 19.930 154.120 20.425 154.290 ;
        RECT 20.595 154.150 20.925 154.510 ;
        RECT 17.195 153.070 17.365 153.760 ;
        RECT 17.535 153.410 17.705 153.590 ;
        RECT 17.875 153.580 18.665 153.830 ;
        RECT 18.870 153.410 19.040 154.120 ;
        RECT 19.210 153.610 19.565 153.830 ;
        RECT 17.535 153.240 19.225 153.410 ;
        RECT 16.040 152.640 16.500 152.930 ;
        RECT 17.195 152.900 18.695 153.070 ;
        RECT 17.195 152.760 17.365 152.900 ;
        RECT 16.805 152.590 17.365 152.760 ;
        RECT 15.280 151.960 15.530 152.420 ;
        RECT 15.700 152.130 16.570 152.470 ;
        RECT 16.805 152.130 16.975 152.590 ;
        RECT 17.810 152.560 18.885 152.730 ;
        RECT 17.145 151.960 17.515 152.420 ;
        RECT 17.810 152.220 17.980 152.560 ;
        RECT 18.150 151.960 18.480 152.390 ;
        RECT 18.715 152.220 18.885 152.560 ;
        RECT 19.055 152.460 19.225 153.240 ;
        RECT 19.395 153.020 19.565 153.610 ;
        RECT 19.735 153.210 20.085 153.830 ;
        RECT 19.395 152.630 19.860 153.020 ;
        RECT 20.255 152.760 20.425 154.120 ;
        RECT 20.595 152.930 21.055 153.980 ;
        RECT 20.030 152.590 20.425 152.760 ;
        RECT 20.030 152.460 20.200 152.590 ;
        RECT 19.055 152.130 19.735 152.460 ;
        RECT 19.950 152.130 20.200 152.460 ;
        RECT 20.370 151.960 20.620 152.420 ;
        RECT 20.790 152.145 21.115 152.930 ;
        RECT 21.285 152.130 21.455 154.250 ;
        RECT 21.625 154.130 21.955 154.510 ;
        RECT 22.125 153.960 22.380 154.250 ;
        RECT 21.630 153.790 22.380 153.960 ;
        RECT 22.670 153.880 22.955 154.340 ;
        RECT 23.125 154.050 23.395 154.510 ;
        RECT 21.630 152.800 21.860 153.790 ;
        RECT 22.670 153.710 23.625 153.880 ;
        RECT 22.030 152.970 22.380 153.620 ;
        RECT 22.555 152.980 23.245 153.540 ;
        RECT 23.415 152.810 23.625 153.710 ;
        RECT 21.630 152.630 22.380 152.800 ;
        RECT 21.625 151.960 21.955 152.460 ;
        RECT 22.125 152.130 22.380 152.630 ;
        RECT 22.670 152.590 23.625 152.810 ;
        RECT 23.795 153.540 24.195 154.340 ;
        RECT 24.385 153.880 24.665 154.340 ;
        RECT 25.185 154.050 25.510 154.510 ;
        RECT 24.385 153.710 25.510 153.880 ;
        RECT 25.680 153.770 26.065 154.340 ;
        RECT 25.060 153.600 25.510 153.710 ;
        RECT 23.795 152.980 24.890 153.540 ;
        RECT 25.060 153.270 25.615 153.600 ;
        RECT 22.670 152.130 22.955 152.590 ;
        RECT 23.125 151.960 23.395 152.420 ;
        RECT 23.795 152.130 24.195 152.980 ;
        RECT 25.060 152.810 25.510 153.270 ;
        RECT 25.785 153.100 26.065 153.770 ;
        RECT 26.235 153.740 27.905 154.510 ;
        RECT 28.075 153.785 28.365 154.510 ;
        RECT 24.385 152.590 25.510 152.810 ;
        RECT 24.385 152.130 24.665 152.590 ;
        RECT 25.185 151.960 25.510 152.420 ;
        RECT 25.680 152.130 26.065 153.100 ;
        RECT 26.235 153.050 26.985 153.570 ;
        RECT 27.155 153.220 27.905 153.740 ;
        RECT 28.540 153.770 28.795 154.340 ;
        RECT 28.965 154.110 29.295 154.510 ;
        RECT 29.720 153.975 30.250 154.340 ;
        RECT 29.720 153.940 29.895 153.975 ;
        RECT 28.965 153.770 29.895 153.940 ;
        RECT 26.235 151.960 27.905 153.050 ;
        RECT 28.075 151.960 28.365 153.125 ;
        RECT 28.540 153.100 28.710 153.770 ;
        RECT 28.965 153.600 29.135 153.770 ;
        RECT 28.880 153.270 29.135 153.600 ;
        RECT 29.360 153.270 29.555 153.600 ;
        RECT 28.540 152.130 28.875 153.100 ;
        RECT 29.045 151.960 29.215 153.100 ;
        RECT 29.385 152.300 29.555 153.270 ;
        RECT 29.725 152.640 29.895 153.770 ;
        RECT 30.065 152.980 30.235 153.780 ;
        RECT 30.440 153.490 30.715 154.340 ;
        RECT 30.435 153.320 30.715 153.490 ;
        RECT 30.440 153.180 30.715 153.320 ;
        RECT 30.885 152.980 31.075 154.340 ;
        RECT 31.255 153.975 31.765 154.510 ;
        RECT 31.985 153.700 32.230 154.305 ;
        RECT 33.135 153.740 35.725 154.510 ;
        RECT 31.275 153.530 32.505 153.700 ;
        RECT 30.065 152.810 31.075 152.980 ;
        RECT 31.245 152.965 31.995 153.155 ;
        RECT 29.725 152.470 30.850 152.640 ;
        RECT 31.245 152.300 31.415 152.965 ;
        RECT 32.165 152.720 32.505 153.530 ;
        RECT 29.385 152.130 31.415 152.300 ;
        RECT 31.585 151.960 31.755 152.720 ;
        RECT 31.990 152.310 32.505 152.720 ;
        RECT 33.135 153.050 34.345 153.570 ;
        RECT 34.515 153.220 35.725 153.740 ;
        RECT 35.895 153.710 36.235 154.340 ;
        RECT 36.405 153.710 36.655 154.510 ;
        RECT 36.845 153.860 37.175 154.340 ;
        RECT 37.345 154.050 37.570 154.510 ;
        RECT 37.740 153.860 38.070 154.340 ;
        RECT 35.895 153.100 36.070 153.710 ;
        RECT 36.845 153.690 38.070 153.860 ;
        RECT 38.700 153.730 39.200 154.340 ;
        RECT 39.665 153.860 39.835 154.340 ;
        RECT 40.015 154.030 40.255 154.510 ;
        RECT 40.505 153.860 40.675 154.340 ;
        RECT 40.845 154.030 41.175 154.510 ;
        RECT 41.345 153.860 41.515 154.340 ;
        RECT 36.240 153.350 36.935 153.520 ;
        RECT 36.765 153.100 36.935 153.350 ;
        RECT 37.110 153.320 37.530 153.520 ;
        RECT 37.700 153.320 38.030 153.520 ;
        RECT 38.200 153.320 38.530 153.520 ;
        RECT 38.700 153.100 38.870 153.730 ;
        RECT 39.665 153.690 40.300 153.860 ;
        RECT 40.505 153.690 41.515 153.860 ;
        RECT 41.685 153.710 42.015 154.510 ;
        RECT 42.335 153.740 44.005 154.510 ;
        RECT 40.130 153.520 40.300 153.690 ;
        RECT 39.055 153.270 39.405 153.520 ;
        RECT 39.580 153.280 39.960 153.520 ;
        RECT 40.130 153.350 40.630 153.520 ;
        RECT 40.130 153.110 40.300 153.350 ;
        RECT 41.020 153.150 41.515 153.690 ;
        RECT 33.135 151.960 35.725 153.050 ;
        RECT 35.895 152.130 36.235 153.100 ;
        RECT 36.405 151.960 36.575 153.100 ;
        RECT 36.765 152.930 39.200 153.100 ;
        RECT 36.845 151.960 37.095 152.760 ;
        RECT 37.740 152.130 38.070 152.930 ;
        RECT 38.370 151.960 38.700 152.760 ;
        RECT 38.870 152.130 39.200 152.930 ;
        RECT 39.585 152.940 40.300 153.110 ;
        RECT 40.505 152.980 41.515 153.150 ;
        RECT 39.585 152.130 39.915 152.940 ;
        RECT 40.085 151.960 40.325 152.760 ;
        RECT 40.505 152.130 40.675 152.980 ;
        RECT 40.845 151.960 41.175 152.760 ;
        RECT 41.345 152.130 41.515 152.980 ;
        RECT 41.685 151.960 42.015 153.110 ;
        RECT 42.335 153.050 43.085 153.570 ;
        RECT 43.255 153.220 44.005 153.740 ;
        RECT 44.550 153.800 44.805 154.330 ;
        RECT 44.985 154.050 45.270 154.510 ;
        RECT 42.335 151.960 44.005 153.050 ;
        RECT 44.550 152.940 44.730 153.800 ;
        RECT 45.450 153.600 45.700 154.250 ;
        RECT 44.900 153.270 45.700 153.600 ;
        RECT 44.550 152.470 44.805 152.940 ;
        RECT 44.465 152.300 44.805 152.470 ;
        RECT 44.550 152.270 44.805 152.300 ;
        RECT 44.985 151.960 45.270 152.760 ;
        RECT 45.450 152.680 45.700 153.270 ;
        RECT 45.900 153.915 46.220 154.245 ;
        RECT 46.400 154.030 47.060 154.510 ;
        RECT 47.260 154.120 48.110 154.290 ;
        RECT 45.900 153.020 46.090 153.915 ;
        RECT 46.410 153.590 47.070 153.860 ;
        RECT 46.740 153.530 47.070 153.590 ;
        RECT 46.260 153.360 46.590 153.420 ;
        RECT 47.260 153.360 47.430 154.120 ;
        RECT 48.670 154.050 48.990 154.510 ;
        RECT 49.190 153.870 49.440 154.300 ;
        RECT 49.730 154.070 50.140 154.510 ;
        RECT 50.310 154.130 51.325 154.330 ;
        RECT 47.600 153.700 48.850 153.870 ;
        RECT 47.600 153.580 47.930 153.700 ;
        RECT 46.260 153.190 48.160 153.360 ;
        RECT 45.900 152.850 47.820 153.020 ;
        RECT 45.900 152.830 46.220 152.850 ;
        RECT 45.450 152.170 45.780 152.680 ;
        RECT 46.050 152.220 46.220 152.830 ;
        RECT 47.990 152.680 48.160 153.190 ;
        RECT 48.330 153.120 48.510 153.530 ;
        RECT 48.680 152.940 48.850 153.700 ;
        RECT 46.390 151.960 46.720 152.650 ;
        RECT 46.950 152.510 48.160 152.680 ;
        RECT 48.330 152.630 48.850 152.940 ;
        RECT 49.020 153.530 49.440 153.870 ;
        RECT 49.730 153.530 50.140 153.860 ;
        RECT 49.020 152.760 49.210 153.530 ;
        RECT 50.310 153.400 50.480 154.130 ;
        RECT 51.625 153.960 51.795 154.290 ;
        RECT 51.965 154.130 52.295 154.510 ;
        RECT 50.650 153.580 51.000 153.950 ;
        RECT 50.310 153.360 50.730 153.400 ;
        RECT 49.380 153.190 50.730 153.360 ;
        RECT 49.380 153.030 49.630 153.190 ;
        RECT 50.140 152.760 50.390 153.020 ;
        RECT 49.020 152.510 50.390 152.760 ;
        RECT 46.950 152.220 47.190 152.510 ;
        RECT 47.990 152.430 48.160 152.510 ;
        RECT 47.390 151.960 47.810 152.340 ;
        RECT 47.990 152.180 48.620 152.430 ;
        RECT 49.090 151.960 49.420 152.340 ;
        RECT 49.590 152.220 49.760 152.510 ;
        RECT 50.560 152.345 50.730 153.190 ;
        RECT 51.180 153.020 51.400 153.890 ;
        RECT 51.625 153.770 52.320 153.960 ;
        RECT 50.900 152.640 51.400 153.020 ;
        RECT 51.570 152.970 51.980 153.590 ;
        RECT 52.150 152.800 52.320 153.770 ;
        RECT 51.625 152.630 52.320 152.800 ;
        RECT 49.940 151.960 50.320 152.340 ;
        RECT 50.560 152.175 51.390 152.345 ;
        RECT 51.625 152.130 51.795 152.630 ;
        RECT 51.965 151.960 52.295 152.460 ;
        RECT 52.510 152.130 52.735 154.250 ;
        RECT 52.905 154.130 53.235 154.510 ;
        RECT 53.405 153.960 53.575 154.250 ;
        RECT 52.910 153.790 53.575 153.960 ;
        RECT 52.910 152.800 53.140 153.790 ;
        RECT 53.835 153.785 54.125 154.510 ;
        RECT 54.295 153.835 54.555 154.340 ;
        RECT 54.735 154.130 55.065 154.510 ;
        RECT 55.245 153.960 55.415 154.340 ;
        RECT 53.310 152.970 53.660 153.620 ;
        RECT 52.910 152.630 53.575 152.800 ;
        RECT 52.905 151.960 53.235 152.460 ;
        RECT 53.405 152.130 53.575 152.630 ;
        RECT 53.835 151.960 54.125 153.125 ;
        RECT 54.295 153.035 54.465 153.835 ;
        RECT 54.750 153.790 55.415 153.960 ;
        RECT 54.750 153.535 54.920 153.790 ;
        RECT 55.675 153.740 59.185 154.510 ;
        RECT 59.445 153.960 59.615 154.340 ;
        RECT 59.830 154.130 60.160 154.510 ;
        RECT 59.445 153.790 60.160 153.960 ;
        RECT 54.635 153.205 54.920 153.535 ;
        RECT 55.155 153.240 55.485 153.610 ;
        RECT 54.750 153.060 54.920 153.205 ;
        RECT 54.295 152.130 54.565 153.035 ;
        RECT 54.750 152.890 55.415 153.060 ;
        RECT 54.735 151.960 55.065 152.720 ;
        RECT 55.245 152.130 55.415 152.890 ;
        RECT 55.675 153.050 57.365 153.570 ;
        RECT 57.535 153.220 59.185 153.740 ;
        RECT 59.355 153.240 59.710 153.610 ;
        RECT 59.990 153.600 60.160 153.790 ;
        RECT 60.330 153.765 60.585 154.340 ;
        RECT 59.990 153.270 60.245 153.600 ;
        RECT 59.990 153.060 60.160 153.270 ;
        RECT 55.675 151.960 59.185 153.050 ;
        RECT 59.445 152.890 60.160 153.060 ;
        RECT 60.415 153.035 60.585 153.765 ;
        RECT 60.760 153.670 61.020 154.510 ;
        RECT 61.285 153.960 61.455 154.340 ;
        RECT 61.670 154.130 62.000 154.510 ;
        RECT 61.285 153.790 62.000 153.960 ;
        RECT 61.195 153.240 61.550 153.610 ;
        RECT 61.830 153.600 62.000 153.790 ;
        RECT 62.170 153.765 62.425 154.340 ;
        RECT 61.830 153.270 62.085 153.600 ;
        RECT 59.445 152.130 59.615 152.890 ;
        RECT 59.830 151.960 60.160 152.720 ;
        RECT 60.330 152.130 60.585 153.035 ;
        RECT 60.760 151.960 61.020 153.110 ;
        RECT 61.830 153.060 62.000 153.270 ;
        RECT 61.285 152.890 62.000 153.060 ;
        RECT 62.255 153.035 62.425 153.765 ;
        RECT 62.600 153.670 62.860 154.510 ;
        RECT 63.555 154.030 63.835 154.510 ;
        RECT 64.005 153.860 64.265 154.250 ;
        RECT 64.440 154.030 64.695 154.510 ;
        RECT 64.865 153.860 65.160 154.250 ;
        RECT 65.340 154.030 65.615 154.510 ;
        RECT 65.785 154.010 66.085 154.340 ;
        RECT 63.510 153.690 65.160 153.860 ;
        RECT 63.510 153.180 63.915 153.690 ;
        RECT 64.085 153.350 65.225 153.520 ;
        RECT 61.285 152.130 61.455 152.890 ;
        RECT 61.670 151.960 62.000 152.720 ;
        RECT 62.170 152.130 62.425 153.035 ;
        RECT 62.600 151.960 62.860 153.110 ;
        RECT 63.510 153.010 64.265 153.180 ;
        RECT 63.550 151.960 63.835 152.830 ;
        RECT 64.005 152.760 64.265 153.010 ;
        RECT 65.055 153.100 65.225 153.350 ;
        RECT 65.395 153.270 65.745 153.840 ;
        RECT 65.915 153.100 66.085 154.010 ;
        RECT 66.345 153.960 66.515 154.340 ;
        RECT 66.730 154.130 67.060 154.510 ;
        RECT 66.345 153.790 67.060 153.960 ;
        RECT 66.255 153.240 66.610 153.610 ;
        RECT 66.890 153.600 67.060 153.790 ;
        RECT 67.230 153.765 67.485 154.340 ;
        RECT 66.890 153.270 67.145 153.600 ;
        RECT 65.055 152.930 66.085 153.100 ;
        RECT 66.890 153.060 67.060 153.270 ;
        RECT 64.005 152.590 65.125 152.760 ;
        RECT 64.005 152.130 64.265 152.590 ;
        RECT 64.440 151.960 64.695 152.420 ;
        RECT 64.865 152.130 65.125 152.590 ;
        RECT 65.295 151.960 65.605 152.760 ;
        RECT 65.775 152.130 66.085 152.930 ;
        RECT 66.345 152.890 67.060 153.060 ;
        RECT 67.315 153.035 67.485 153.765 ;
        RECT 67.660 153.670 67.920 154.510 ;
        RECT 68.185 153.960 68.355 154.340 ;
        RECT 68.570 154.130 68.900 154.510 ;
        RECT 68.185 153.790 68.900 153.960 ;
        RECT 68.095 153.240 68.450 153.610 ;
        RECT 68.730 153.600 68.900 153.790 ;
        RECT 69.070 153.765 69.325 154.340 ;
        RECT 68.730 153.270 68.985 153.600 ;
        RECT 66.345 152.130 66.515 152.890 ;
        RECT 66.730 151.960 67.060 152.720 ;
        RECT 67.230 152.130 67.485 153.035 ;
        RECT 67.660 151.960 67.920 153.110 ;
        RECT 68.730 153.060 68.900 153.270 ;
        RECT 68.185 152.890 68.900 153.060 ;
        RECT 69.155 153.035 69.325 153.765 ;
        RECT 69.500 153.670 69.760 154.510 ;
        RECT 70.025 153.960 70.195 154.340 ;
        RECT 70.410 154.130 70.740 154.510 ;
        RECT 70.025 153.790 70.740 153.960 ;
        RECT 69.935 153.240 70.290 153.610 ;
        RECT 70.570 153.600 70.740 153.790 ;
        RECT 70.910 153.765 71.165 154.340 ;
        RECT 70.570 153.270 70.825 153.600 ;
        RECT 68.185 152.130 68.355 152.890 ;
        RECT 68.570 151.960 68.900 152.720 ;
        RECT 69.070 152.130 69.325 153.035 ;
        RECT 69.500 151.960 69.760 153.110 ;
        RECT 70.570 153.060 70.740 153.270 ;
        RECT 70.025 152.890 70.740 153.060 ;
        RECT 70.995 153.035 71.165 153.765 ;
        RECT 71.340 153.670 71.600 154.510 ;
        RECT 71.980 153.730 72.480 154.340 ;
        RECT 71.775 153.270 72.125 153.520 ;
        RECT 70.025 152.130 70.195 152.890 ;
        RECT 70.410 151.960 70.740 152.720 ;
        RECT 70.910 152.130 71.165 153.035 ;
        RECT 71.340 151.960 71.600 153.110 ;
        RECT 72.310 153.100 72.480 153.730 ;
        RECT 73.110 153.860 73.440 154.340 ;
        RECT 73.610 154.050 73.835 154.510 ;
        RECT 74.005 153.860 74.335 154.340 ;
        RECT 73.110 153.690 74.335 153.860 ;
        RECT 74.525 153.710 74.775 154.510 ;
        RECT 74.945 153.710 75.285 154.340 ;
        RECT 75.915 153.740 79.425 154.510 ;
        RECT 79.595 153.785 79.885 154.510 ;
        RECT 80.430 154.170 80.685 154.330 ;
        RECT 80.345 154.000 80.685 154.170 ;
        RECT 80.865 154.050 81.150 154.510 ;
        RECT 80.430 153.800 80.685 154.000 ;
        RECT 72.650 153.320 72.980 153.520 ;
        RECT 73.150 153.320 73.480 153.520 ;
        RECT 73.650 153.320 74.070 153.520 ;
        RECT 74.245 153.350 74.940 153.520 ;
        RECT 74.245 153.100 74.415 153.350 ;
        RECT 75.110 153.100 75.285 153.710 ;
        RECT 71.980 152.930 74.415 153.100 ;
        RECT 71.980 152.130 72.310 152.930 ;
        RECT 72.480 151.960 72.810 152.760 ;
        RECT 73.110 152.130 73.440 152.930 ;
        RECT 74.085 151.960 74.335 152.760 ;
        RECT 74.605 151.960 74.775 153.100 ;
        RECT 74.945 152.130 75.285 153.100 ;
        RECT 75.915 153.050 77.605 153.570 ;
        RECT 77.775 153.220 79.425 153.740 ;
        RECT 75.915 151.960 79.425 153.050 ;
        RECT 79.595 151.960 79.885 153.125 ;
        RECT 80.430 152.940 80.610 153.800 ;
        RECT 81.330 153.600 81.580 154.250 ;
        RECT 80.780 153.270 81.580 153.600 ;
        RECT 80.430 152.270 80.685 152.940 ;
        RECT 80.865 151.960 81.150 152.760 ;
        RECT 81.330 152.680 81.580 153.270 ;
        RECT 81.780 153.915 82.100 154.245 ;
        RECT 82.280 154.030 82.940 154.510 ;
        RECT 83.140 154.120 83.990 154.290 ;
        RECT 81.780 153.020 81.970 153.915 ;
        RECT 82.290 153.590 82.950 153.860 ;
        RECT 82.620 153.530 82.950 153.590 ;
        RECT 82.140 153.360 82.470 153.420 ;
        RECT 83.140 153.360 83.310 154.120 ;
        RECT 84.550 154.050 84.870 154.510 ;
        RECT 85.070 153.870 85.320 154.300 ;
        RECT 85.610 154.070 86.020 154.510 ;
        RECT 86.190 154.130 87.205 154.330 ;
        RECT 83.480 153.700 84.730 153.870 ;
        RECT 83.480 153.580 83.810 153.700 ;
        RECT 82.140 153.190 84.040 153.360 ;
        RECT 81.780 152.850 83.700 153.020 ;
        RECT 81.780 152.830 82.100 152.850 ;
        RECT 81.330 152.170 81.660 152.680 ;
        RECT 81.930 152.220 82.100 152.830 ;
        RECT 83.870 152.680 84.040 153.190 ;
        RECT 84.210 153.120 84.390 153.530 ;
        RECT 84.560 152.940 84.730 153.700 ;
        RECT 82.270 151.960 82.600 152.650 ;
        RECT 82.830 152.510 84.040 152.680 ;
        RECT 84.210 152.630 84.730 152.940 ;
        RECT 84.900 153.530 85.320 153.870 ;
        RECT 85.610 153.530 86.020 153.860 ;
        RECT 84.900 152.760 85.090 153.530 ;
        RECT 86.190 153.400 86.360 154.130 ;
        RECT 87.505 153.960 87.675 154.290 ;
        RECT 87.845 154.130 88.175 154.510 ;
        RECT 86.530 153.580 86.880 153.950 ;
        RECT 86.190 153.360 86.610 153.400 ;
        RECT 85.260 153.190 86.610 153.360 ;
        RECT 85.260 153.030 85.510 153.190 ;
        RECT 86.020 152.760 86.270 153.020 ;
        RECT 84.900 152.510 86.270 152.760 ;
        RECT 82.830 152.220 83.070 152.510 ;
        RECT 83.870 152.430 84.040 152.510 ;
        RECT 83.270 151.960 83.690 152.340 ;
        RECT 83.870 152.180 84.500 152.430 ;
        RECT 84.970 151.960 85.300 152.340 ;
        RECT 85.470 152.220 85.640 152.510 ;
        RECT 86.440 152.345 86.610 153.190 ;
        RECT 87.060 153.020 87.280 153.890 ;
        RECT 87.505 153.770 88.200 153.960 ;
        RECT 86.780 152.640 87.280 153.020 ;
        RECT 87.450 152.970 87.860 153.590 ;
        RECT 88.030 152.800 88.200 153.770 ;
        RECT 87.505 152.630 88.200 152.800 ;
        RECT 85.820 151.960 86.200 152.340 ;
        RECT 86.440 152.175 87.270 152.345 ;
        RECT 87.505 152.130 87.675 152.630 ;
        RECT 87.845 151.960 88.175 152.460 ;
        RECT 88.390 152.130 88.615 154.250 ;
        RECT 88.785 154.130 89.115 154.510 ;
        RECT 89.285 153.960 89.455 154.250 ;
        RECT 88.790 153.790 89.455 153.960 ;
        RECT 90.175 153.835 90.445 154.180 ;
        RECT 90.635 154.110 91.015 154.510 ;
        RECT 91.185 153.940 91.355 154.290 ;
        RECT 91.525 154.110 91.855 154.510 ;
        RECT 92.055 153.940 92.225 154.290 ;
        RECT 92.425 154.010 92.755 154.510 ;
        RECT 88.790 152.800 89.020 153.790 ;
        RECT 89.190 152.970 89.540 153.620 ;
        RECT 90.175 153.100 90.345 153.835 ;
        RECT 90.615 153.770 92.225 153.940 ;
        RECT 90.615 153.600 90.785 153.770 ;
        RECT 90.515 153.270 90.785 153.600 ;
        RECT 90.955 153.270 91.360 153.600 ;
        RECT 90.615 153.100 90.785 153.270 ;
        RECT 91.530 153.150 92.240 153.600 ;
        RECT 92.410 153.270 92.760 153.840 ;
        RECT 92.935 153.710 93.275 154.340 ;
        RECT 93.445 153.710 93.695 154.510 ;
        RECT 93.885 153.860 94.215 154.340 ;
        RECT 94.385 154.050 94.610 154.510 ;
        RECT 94.780 153.860 95.110 154.340 ;
        RECT 92.935 153.660 93.165 153.710 ;
        RECT 93.885 153.690 95.110 153.860 ;
        RECT 95.740 153.730 96.240 154.340 ;
        RECT 97.075 153.740 98.745 154.510 ;
        RECT 88.790 152.630 89.455 152.800 ;
        RECT 88.785 151.960 89.115 152.460 ;
        RECT 89.285 152.130 89.455 152.630 ;
        RECT 90.175 152.130 90.445 153.100 ;
        RECT 90.615 152.930 91.340 153.100 ;
        RECT 91.530 152.980 92.245 153.150 ;
        RECT 92.935 153.100 93.110 153.660 ;
        RECT 93.280 153.350 93.975 153.520 ;
        RECT 93.805 153.100 93.975 153.350 ;
        RECT 94.150 153.320 94.570 153.520 ;
        RECT 94.740 153.320 95.070 153.520 ;
        RECT 95.240 153.320 95.570 153.520 ;
        RECT 95.740 153.100 95.910 153.730 ;
        RECT 96.095 153.270 96.445 153.520 ;
        RECT 91.170 152.810 91.340 152.930 ;
        RECT 92.440 152.810 92.760 153.100 ;
        RECT 90.655 151.960 90.935 152.760 ;
        RECT 91.170 152.640 92.760 152.810 ;
        RECT 91.105 152.180 92.760 152.470 ;
        RECT 92.935 152.130 93.275 153.100 ;
        RECT 93.445 151.960 93.615 153.100 ;
        RECT 93.805 152.930 96.240 153.100 ;
        RECT 93.885 151.960 94.135 152.760 ;
        RECT 94.780 152.130 95.110 152.930 ;
        RECT 95.410 151.960 95.740 152.760 ;
        RECT 95.910 152.130 96.240 152.930 ;
        RECT 97.075 153.050 97.825 153.570 ;
        RECT 97.995 153.220 98.745 153.740 ;
        RECT 98.915 153.710 99.255 154.340 ;
        RECT 99.425 153.710 99.675 154.510 ;
        RECT 99.865 153.860 100.195 154.340 ;
        RECT 100.365 154.050 100.590 154.510 ;
        RECT 100.760 153.860 101.090 154.340 ;
        RECT 98.915 153.100 99.090 153.710 ;
        RECT 99.865 153.690 101.090 153.860 ;
        RECT 101.720 153.730 102.220 154.340 ;
        RECT 102.595 153.740 105.185 154.510 ;
        RECT 105.355 153.785 105.645 154.510 ;
        RECT 105.815 153.760 107.025 154.510 ;
        RECT 99.260 153.350 99.955 153.520 ;
        RECT 99.785 153.100 99.955 153.350 ;
        RECT 100.130 153.320 100.550 153.520 ;
        RECT 100.720 153.320 101.050 153.520 ;
        RECT 101.220 153.320 101.550 153.520 ;
        RECT 101.720 153.100 101.890 153.730 ;
        RECT 102.075 153.270 102.425 153.520 ;
        RECT 97.075 151.960 98.745 153.050 ;
        RECT 98.915 152.130 99.255 153.100 ;
        RECT 99.425 151.960 99.595 153.100 ;
        RECT 99.785 152.930 102.220 153.100 ;
        RECT 99.865 151.960 100.115 152.760 ;
        RECT 100.760 152.130 101.090 152.930 ;
        RECT 101.390 151.960 101.720 152.760 ;
        RECT 101.890 152.130 102.220 152.930 ;
        RECT 102.595 153.050 103.805 153.570 ;
        RECT 103.975 153.220 105.185 153.740 ;
        RECT 102.595 151.960 105.185 153.050 ;
        RECT 105.355 151.960 105.645 153.125 ;
        RECT 105.815 153.050 106.335 153.590 ;
        RECT 106.505 153.220 107.025 153.760 ;
        RECT 107.470 153.700 107.715 154.305 ;
        RECT 107.935 153.975 108.445 154.510 ;
        RECT 107.195 153.530 108.425 153.700 ;
        RECT 105.815 151.960 107.025 153.050 ;
        RECT 107.195 152.720 107.535 153.530 ;
        RECT 107.705 152.965 108.455 153.155 ;
        RECT 107.195 152.310 107.710 152.720 ;
        RECT 107.945 151.960 108.115 152.720 ;
        RECT 108.285 152.300 108.455 152.965 ;
        RECT 108.625 152.980 108.815 154.340 ;
        RECT 108.985 154.170 109.260 154.340 ;
        RECT 108.985 154.000 109.265 154.170 ;
        RECT 108.985 153.180 109.260 154.000 ;
        RECT 109.450 153.975 109.980 154.340 ;
        RECT 110.405 154.110 110.735 154.510 ;
        RECT 109.805 153.940 109.980 153.975 ;
        RECT 109.465 152.980 109.635 153.780 ;
        RECT 108.625 152.810 109.635 152.980 ;
        RECT 109.805 153.770 110.735 153.940 ;
        RECT 110.905 153.770 111.160 154.340 ;
        RECT 109.805 152.640 109.975 153.770 ;
        RECT 110.565 153.600 110.735 153.770 ;
        RECT 108.850 152.470 109.975 152.640 ;
        RECT 110.145 153.270 110.340 153.600 ;
        RECT 110.565 153.270 110.820 153.600 ;
        RECT 110.145 152.300 110.315 153.270 ;
        RECT 110.990 153.100 111.160 153.770 ;
        RECT 111.485 153.710 111.815 154.510 ;
        RECT 111.985 153.860 112.155 154.340 ;
        RECT 112.325 154.030 112.655 154.510 ;
        RECT 112.825 153.860 112.995 154.340 ;
        RECT 113.245 154.030 113.485 154.510 ;
        RECT 113.665 153.860 113.835 154.340 ;
        RECT 111.985 153.690 112.995 153.860 ;
        RECT 113.200 153.690 113.835 153.860 ;
        RECT 114.555 153.740 117.145 154.510 ;
        RECT 117.315 153.760 118.525 154.510 ;
        RECT 111.985 153.150 112.480 153.690 ;
        RECT 113.200 153.520 113.370 153.690 ;
        RECT 112.870 153.350 113.370 153.520 ;
        RECT 108.285 152.130 110.315 152.300 ;
        RECT 110.485 151.960 110.655 153.100 ;
        RECT 110.825 152.130 111.160 153.100 ;
        RECT 111.485 151.960 111.815 153.110 ;
        RECT 111.985 152.980 112.995 153.150 ;
        RECT 111.985 152.130 112.155 152.980 ;
        RECT 112.325 151.960 112.655 152.760 ;
        RECT 112.825 152.130 112.995 152.980 ;
        RECT 113.200 153.110 113.370 153.350 ;
        RECT 113.540 153.280 113.920 153.520 ;
        RECT 113.200 152.940 113.915 153.110 ;
        RECT 113.175 151.960 113.415 152.760 ;
        RECT 113.585 152.130 113.915 152.940 ;
        RECT 114.555 153.050 115.765 153.570 ;
        RECT 115.935 153.220 117.145 153.740 ;
        RECT 117.315 153.050 117.835 153.590 ;
        RECT 118.005 153.220 118.525 153.760 ;
        RECT 114.555 151.960 117.145 153.050 ;
        RECT 117.315 151.960 118.525 153.050 ;
        RECT 11.430 151.790 118.610 151.960 ;
        RECT 11.515 150.700 12.725 151.790 ;
        RECT 11.515 149.990 12.035 150.530 ;
        RECT 12.205 150.160 12.725 150.700 ;
        RECT 13.355 150.700 15.025 151.790 ;
        RECT 13.355 150.180 14.105 150.700 ;
        RECT 15.195 150.625 15.485 151.790 ;
        RECT 16.115 150.700 17.785 151.790 ;
        RECT 17.955 151.030 18.470 151.440 ;
        RECT 18.705 151.030 18.875 151.790 ;
        RECT 19.045 151.450 21.075 151.620 ;
        RECT 14.275 150.010 15.025 150.530 ;
        RECT 16.115 150.180 16.865 150.700 ;
        RECT 17.035 150.010 17.785 150.530 ;
        RECT 17.955 150.220 18.295 151.030 ;
        RECT 19.045 150.785 19.215 151.450 ;
        RECT 19.610 151.110 20.735 151.280 ;
        RECT 18.465 150.595 19.215 150.785 ;
        RECT 19.385 150.770 20.395 150.940 ;
        RECT 17.955 150.050 19.185 150.220 ;
        RECT 11.515 149.240 12.725 149.990 ;
        RECT 13.355 149.240 15.025 150.010 ;
        RECT 15.195 149.240 15.485 149.965 ;
        RECT 16.115 149.240 17.785 150.010 ;
        RECT 18.230 149.445 18.475 150.050 ;
        RECT 18.695 149.240 19.205 149.775 ;
        RECT 19.385 149.410 19.575 150.770 ;
        RECT 19.745 149.750 20.020 150.570 ;
        RECT 20.225 149.970 20.395 150.770 ;
        RECT 20.565 149.980 20.735 151.110 ;
        RECT 20.905 150.480 21.075 151.450 ;
        RECT 21.245 150.650 21.415 151.790 ;
        RECT 21.585 150.650 21.920 151.620 ;
        RECT 22.135 150.650 22.365 151.790 ;
        RECT 20.905 150.150 21.100 150.480 ;
        RECT 21.325 150.150 21.580 150.480 ;
        RECT 21.325 149.980 21.495 150.150 ;
        RECT 21.750 149.980 21.920 150.650 ;
        RECT 22.535 150.640 22.865 151.620 ;
        RECT 23.035 150.650 23.245 151.790 ;
        RECT 22.115 150.230 22.445 150.480 ;
        RECT 20.565 149.810 21.495 149.980 ;
        RECT 20.565 149.775 20.740 149.810 ;
        RECT 19.745 149.580 20.025 149.750 ;
        RECT 19.745 149.410 20.020 149.580 ;
        RECT 20.210 149.410 20.740 149.775 ;
        RECT 21.165 149.240 21.495 149.640 ;
        RECT 21.665 149.410 21.920 149.980 ;
        RECT 22.135 149.240 22.365 150.060 ;
        RECT 22.615 150.040 22.865 150.640 ;
        RECT 23.480 150.600 23.735 151.480 ;
        RECT 23.905 150.650 24.210 151.790 ;
        RECT 24.550 151.410 24.880 151.790 ;
        RECT 25.060 151.240 25.230 151.530 ;
        RECT 25.400 151.330 25.650 151.790 ;
        RECT 24.430 151.070 25.230 151.240 ;
        RECT 25.820 151.280 26.690 151.620 ;
        RECT 22.535 149.410 22.865 150.040 ;
        RECT 23.035 149.240 23.245 150.060 ;
        RECT 23.480 149.950 23.690 150.600 ;
        RECT 24.430 150.480 24.600 151.070 ;
        RECT 25.820 150.900 25.990 151.280 ;
        RECT 26.925 151.160 27.095 151.620 ;
        RECT 27.265 151.330 27.635 151.790 ;
        RECT 27.930 151.190 28.100 151.530 ;
        RECT 28.270 151.360 28.600 151.790 ;
        RECT 28.835 151.190 29.005 151.530 ;
        RECT 24.770 150.730 25.990 150.900 ;
        RECT 26.160 150.820 26.620 151.110 ;
        RECT 26.925 150.990 27.485 151.160 ;
        RECT 27.930 151.020 29.005 151.190 ;
        RECT 29.175 151.290 29.855 151.620 ;
        RECT 30.070 151.290 30.320 151.620 ;
        RECT 30.490 151.330 30.740 151.790 ;
        RECT 27.315 150.850 27.485 150.990 ;
        RECT 26.160 150.810 27.125 150.820 ;
        RECT 25.820 150.640 25.990 150.730 ;
        RECT 26.450 150.650 27.125 150.810 ;
        RECT 23.860 150.450 24.600 150.480 ;
        RECT 23.860 150.150 24.775 150.450 ;
        RECT 24.450 149.975 24.775 150.150 ;
        RECT 23.480 149.420 23.735 149.950 ;
        RECT 23.905 149.240 24.210 149.700 ;
        RECT 24.455 149.620 24.775 149.975 ;
        RECT 24.945 150.190 25.485 150.560 ;
        RECT 25.820 150.470 26.225 150.640 ;
        RECT 24.945 149.790 25.185 150.190 ;
        RECT 25.665 150.020 25.885 150.300 ;
        RECT 25.355 149.850 25.885 150.020 ;
        RECT 25.355 149.620 25.525 149.850 ;
        RECT 26.055 149.690 26.225 150.470 ;
        RECT 26.395 149.860 26.745 150.480 ;
        RECT 26.915 149.860 27.125 150.650 ;
        RECT 27.315 150.680 28.815 150.850 ;
        RECT 27.315 149.990 27.485 150.680 ;
        RECT 29.175 150.510 29.345 151.290 ;
        RECT 30.150 151.160 30.320 151.290 ;
        RECT 27.655 150.340 29.345 150.510 ;
        RECT 29.515 150.730 29.980 151.120 ;
        RECT 30.150 150.990 30.545 151.160 ;
        RECT 27.655 150.160 27.825 150.340 ;
        RECT 24.455 149.450 25.525 149.620 ;
        RECT 25.695 149.240 25.885 149.680 ;
        RECT 26.055 149.410 27.005 149.690 ;
        RECT 27.315 149.600 27.575 149.990 ;
        RECT 27.995 149.920 28.785 150.170 ;
        RECT 27.225 149.430 27.575 149.600 ;
        RECT 27.785 149.240 28.115 149.700 ;
        RECT 28.990 149.630 29.160 150.340 ;
        RECT 29.515 150.140 29.685 150.730 ;
        RECT 29.330 149.920 29.685 150.140 ;
        RECT 29.855 149.920 30.205 150.540 ;
        RECT 30.375 149.630 30.545 150.990 ;
        RECT 30.910 150.820 31.235 151.605 ;
        RECT 30.715 149.770 31.175 150.820 ;
        RECT 28.990 149.460 29.845 149.630 ;
        RECT 30.050 149.460 30.545 149.630 ;
        RECT 30.715 149.240 31.045 149.600 ;
        RECT 31.405 149.500 31.575 151.620 ;
        RECT 31.745 151.290 32.075 151.790 ;
        RECT 32.245 151.120 32.500 151.620 ;
        RECT 31.750 150.950 32.500 151.120 ;
        RECT 31.750 149.960 31.980 150.950 ;
        RECT 32.150 150.130 32.500 150.780 ;
        RECT 33.135 150.700 34.805 151.790 ;
        RECT 33.135 150.180 33.885 150.700 ;
        RECT 34.975 150.650 35.315 151.620 ;
        RECT 35.485 150.650 35.655 151.790 ;
        RECT 35.925 150.990 36.175 151.790 ;
        RECT 36.820 150.820 37.150 151.620 ;
        RECT 37.450 150.990 37.780 151.790 ;
        RECT 37.950 150.820 38.280 151.620 ;
        RECT 35.845 150.650 38.280 150.820 ;
        RECT 39.115 150.700 40.785 151.790 ;
        RECT 34.055 150.010 34.805 150.530 ;
        RECT 31.750 149.790 32.500 149.960 ;
        RECT 31.745 149.240 32.075 149.620 ;
        RECT 32.245 149.500 32.500 149.790 ;
        RECT 33.135 149.240 34.805 150.010 ;
        RECT 34.975 150.040 35.150 150.650 ;
        RECT 35.845 150.400 36.015 150.650 ;
        RECT 35.320 150.230 36.015 150.400 ;
        RECT 36.190 150.230 36.610 150.430 ;
        RECT 36.780 150.230 37.110 150.430 ;
        RECT 37.280 150.230 37.610 150.430 ;
        RECT 34.975 149.410 35.315 150.040 ;
        RECT 35.485 149.240 35.735 150.040 ;
        RECT 35.925 149.890 37.150 150.060 ;
        RECT 35.925 149.410 36.255 149.890 ;
        RECT 36.425 149.240 36.650 149.700 ;
        RECT 36.820 149.410 37.150 149.890 ;
        RECT 37.780 150.020 37.950 150.650 ;
        RECT 38.135 150.230 38.485 150.480 ;
        RECT 39.115 150.180 39.865 150.700 ;
        RECT 40.955 150.625 41.245 151.790 ;
        RECT 41.415 150.700 44.005 151.790 ;
        RECT 37.780 149.410 38.280 150.020 ;
        RECT 40.035 150.010 40.785 150.530 ;
        RECT 41.415 150.180 42.625 150.700 ;
        RECT 44.175 150.650 44.515 151.620 ;
        RECT 44.685 150.650 44.855 151.790 ;
        RECT 45.125 150.990 45.375 151.790 ;
        RECT 46.020 150.820 46.350 151.620 ;
        RECT 46.650 150.990 46.980 151.790 ;
        RECT 47.150 150.820 47.480 151.620 ;
        RECT 45.045 150.650 47.480 150.820 ;
        RECT 47.855 150.700 49.525 151.790 ;
        RECT 49.695 151.030 50.210 151.440 ;
        RECT 50.445 151.030 50.615 151.790 ;
        RECT 50.785 151.450 52.815 151.620 ;
        RECT 42.795 150.010 44.005 150.530 ;
        RECT 39.115 149.240 40.785 150.010 ;
        RECT 40.955 149.240 41.245 149.965 ;
        RECT 41.415 149.240 44.005 150.010 ;
        RECT 44.175 150.040 44.350 150.650 ;
        RECT 45.045 150.400 45.215 150.650 ;
        RECT 44.520 150.230 45.215 150.400 ;
        RECT 45.390 150.230 45.810 150.430 ;
        RECT 45.980 150.230 46.310 150.430 ;
        RECT 46.480 150.230 46.810 150.430 ;
        RECT 44.175 149.410 44.515 150.040 ;
        RECT 44.685 149.240 44.935 150.040 ;
        RECT 45.125 149.890 46.350 150.060 ;
        RECT 45.125 149.410 45.455 149.890 ;
        RECT 45.625 149.240 45.850 149.700 ;
        RECT 46.020 149.410 46.350 149.890 ;
        RECT 46.980 150.020 47.150 150.650 ;
        RECT 47.335 150.230 47.685 150.480 ;
        RECT 47.855 150.180 48.605 150.700 ;
        RECT 46.980 149.410 47.480 150.020 ;
        RECT 48.775 150.010 49.525 150.530 ;
        RECT 49.695 150.220 50.035 151.030 ;
        RECT 50.785 150.785 50.955 151.450 ;
        RECT 51.350 151.110 52.475 151.280 ;
        RECT 50.205 150.595 50.955 150.785 ;
        RECT 51.125 150.770 52.135 150.940 ;
        RECT 49.695 150.050 50.925 150.220 ;
        RECT 47.855 149.240 49.525 150.010 ;
        RECT 49.970 149.445 50.215 150.050 ;
        RECT 50.435 149.240 50.945 149.775 ;
        RECT 51.125 149.410 51.315 150.770 ;
        RECT 51.485 150.090 51.760 150.570 ;
        RECT 51.485 149.920 51.765 150.090 ;
        RECT 51.965 149.970 52.135 150.770 ;
        RECT 52.305 149.980 52.475 151.110 ;
        RECT 52.645 150.480 52.815 151.450 ;
        RECT 52.985 150.650 53.155 151.790 ;
        RECT 53.325 150.650 53.660 151.620 ;
        RECT 52.645 150.150 52.840 150.480 ;
        RECT 53.065 150.150 53.320 150.480 ;
        RECT 53.065 149.980 53.235 150.150 ;
        RECT 53.490 149.980 53.660 150.650 ;
        RECT 53.835 150.700 57.345 151.790 ;
        RECT 57.520 151.355 62.865 151.790 ;
        RECT 53.835 150.180 55.525 150.700 ;
        RECT 55.695 150.010 57.345 150.530 ;
        RECT 59.110 150.105 59.460 151.355 ;
        RECT 63.095 150.650 63.305 151.790 ;
        RECT 63.475 150.640 63.805 151.620 ;
        RECT 63.975 150.650 64.205 151.790 ;
        RECT 64.875 150.700 66.545 151.790 ;
        RECT 51.485 149.410 51.760 149.920 ;
        RECT 52.305 149.810 53.235 149.980 ;
        RECT 52.305 149.775 52.480 149.810 ;
        RECT 51.950 149.410 52.480 149.775 ;
        RECT 52.905 149.240 53.235 149.640 ;
        RECT 53.405 149.410 53.660 149.980 ;
        RECT 53.835 149.240 57.345 150.010 ;
        RECT 60.940 149.785 61.280 150.615 ;
        RECT 57.520 149.240 62.865 149.785 ;
        RECT 63.095 149.240 63.305 150.060 ;
        RECT 63.475 150.040 63.725 150.640 ;
        RECT 63.895 150.230 64.225 150.480 ;
        RECT 64.875 150.180 65.625 150.700 ;
        RECT 66.715 150.625 67.005 151.790 ;
        RECT 67.635 150.700 71.145 151.790 ;
        RECT 71.520 150.820 71.850 151.620 ;
        RECT 72.020 150.990 72.350 151.790 ;
        RECT 72.650 150.820 72.980 151.620 ;
        RECT 73.625 150.990 73.875 151.790 ;
        RECT 63.475 149.410 63.805 150.040 ;
        RECT 63.975 149.240 64.205 150.060 ;
        RECT 65.795 150.010 66.545 150.530 ;
        RECT 67.635 150.180 69.325 150.700 ;
        RECT 71.520 150.650 73.955 150.820 ;
        RECT 74.145 150.650 74.315 151.790 ;
        RECT 74.485 150.650 74.825 151.620 ;
        RECT 69.495 150.010 71.145 150.530 ;
        RECT 71.315 150.230 71.665 150.480 ;
        RECT 71.850 150.020 72.020 150.650 ;
        RECT 72.190 150.230 72.520 150.430 ;
        RECT 72.690 150.230 73.020 150.430 ;
        RECT 73.190 150.230 73.610 150.430 ;
        RECT 73.785 150.400 73.955 150.650 ;
        RECT 73.785 150.230 74.480 150.400 ;
        RECT 64.875 149.240 66.545 150.010 ;
        RECT 66.715 149.240 67.005 149.965 ;
        RECT 67.635 149.240 71.145 150.010 ;
        RECT 71.520 149.410 72.020 150.020 ;
        RECT 72.650 149.890 73.875 150.060 ;
        RECT 74.650 150.040 74.825 150.650 ;
        RECT 72.650 149.410 72.980 149.890 ;
        RECT 73.150 149.240 73.375 149.700 ;
        RECT 73.545 149.410 73.875 149.890 ;
        RECT 74.065 149.240 74.315 150.040 ;
        RECT 74.485 149.410 74.825 150.040 ;
        RECT 74.995 150.650 75.335 151.620 ;
        RECT 75.505 150.650 75.675 151.790 ;
        RECT 75.945 150.990 76.195 151.790 ;
        RECT 76.840 150.820 77.170 151.620 ;
        RECT 77.470 150.990 77.800 151.790 ;
        RECT 77.970 150.820 78.300 151.620 ;
        RECT 75.865 150.650 78.300 150.820 ;
        RECT 78.675 150.700 80.345 151.790 ;
        RECT 80.515 151.030 81.030 151.440 ;
        RECT 81.265 151.030 81.435 151.790 ;
        RECT 81.605 151.450 83.635 151.620 ;
        RECT 74.995 150.040 75.170 150.650 ;
        RECT 75.865 150.400 76.035 150.650 ;
        RECT 75.340 150.230 76.035 150.400 ;
        RECT 76.210 150.230 76.630 150.430 ;
        RECT 76.800 150.230 77.130 150.430 ;
        RECT 77.300 150.230 77.630 150.430 ;
        RECT 74.995 149.410 75.335 150.040 ;
        RECT 75.505 149.240 75.755 150.040 ;
        RECT 75.945 149.890 77.170 150.060 ;
        RECT 75.945 149.410 76.275 149.890 ;
        RECT 76.445 149.240 76.670 149.700 ;
        RECT 76.840 149.410 77.170 149.890 ;
        RECT 77.800 150.020 77.970 150.650 ;
        RECT 78.155 150.230 78.505 150.480 ;
        RECT 78.675 150.180 79.425 150.700 ;
        RECT 77.800 149.410 78.300 150.020 ;
        RECT 79.595 150.010 80.345 150.530 ;
        RECT 80.515 150.220 80.855 151.030 ;
        RECT 81.605 150.785 81.775 151.450 ;
        RECT 82.170 151.110 83.295 151.280 ;
        RECT 81.025 150.595 81.775 150.785 ;
        RECT 81.945 150.770 82.955 150.940 ;
        RECT 80.515 150.050 81.745 150.220 ;
        RECT 78.675 149.240 80.345 150.010 ;
        RECT 80.790 149.445 81.035 150.050 ;
        RECT 81.255 149.240 81.765 149.775 ;
        RECT 81.945 149.410 82.135 150.770 ;
        RECT 82.305 149.750 82.580 150.570 ;
        RECT 82.785 149.970 82.955 150.770 ;
        RECT 83.125 149.980 83.295 151.110 ;
        RECT 83.465 150.480 83.635 151.450 ;
        RECT 83.805 150.650 83.975 151.790 ;
        RECT 84.145 150.650 84.480 151.620 ;
        RECT 85.175 150.650 85.385 151.790 ;
        RECT 83.465 150.150 83.660 150.480 ;
        RECT 83.885 150.150 84.140 150.480 ;
        RECT 83.885 149.980 84.055 150.150 ;
        RECT 84.310 149.980 84.480 150.650 ;
        RECT 85.555 150.640 85.885 151.620 ;
        RECT 86.055 150.650 86.285 151.790 ;
        RECT 86.585 150.860 86.755 151.620 ;
        RECT 86.935 151.030 87.265 151.790 ;
        RECT 86.585 150.690 87.250 150.860 ;
        RECT 87.435 150.715 87.705 151.620 ;
        RECT 83.125 149.810 84.055 149.980 ;
        RECT 83.125 149.775 83.300 149.810 ;
        RECT 82.305 149.580 82.585 149.750 ;
        RECT 82.305 149.410 82.580 149.580 ;
        RECT 82.770 149.410 83.300 149.775 ;
        RECT 83.725 149.240 84.055 149.640 ;
        RECT 84.225 149.410 84.480 149.980 ;
        RECT 85.175 149.240 85.385 150.060 ;
        RECT 85.555 150.040 85.805 150.640 ;
        RECT 87.080 150.545 87.250 150.690 ;
        RECT 85.975 150.230 86.305 150.480 ;
        RECT 86.515 150.140 86.845 150.510 ;
        RECT 87.080 150.215 87.365 150.545 ;
        RECT 85.555 149.410 85.885 150.040 ;
        RECT 86.055 149.240 86.285 150.060 ;
        RECT 87.080 149.960 87.250 150.215 ;
        RECT 86.585 149.790 87.250 149.960 ;
        RECT 87.535 149.915 87.705 150.715 ;
        RECT 88.795 150.700 92.305 151.790 ;
        RECT 88.795 150.180 90.485 150.700 ;
        RECT 92.475 150.625 92.765 151.790 ;
        RECT 93.860 151.355 99.205 151.790 ;
        RECT 90.655 150.010 92.305 150.530 ;
        RECT 95.450 150.105 95.800 151.355 ;
        RECT 99.380 151.280 101.035 151.570 ;
        RECT 99.380 150.940 100.970 151.110 ;
        RECT 101.205 150.990 101.485 151.790 ;
        RECT 99.380 150.650 99.700 150.940 ;
        RECT 100.800 150.820 100.970 150.940 ;
        RECT 86.585 149.410 86.755 149.790 ;
        RECT 86.935 149.240 87.265 149.620 ;
        RECT 87.445 149.410 87.705 149.915 ;
        RECT 88.795 149.240 92.305 150.010 ;
        RECT 92.475 149.240 92.765 149.965 ;
        RECT 97.280 149.785 97.620 150.615 ;
        RECT 99.895 150.600 100.610 150.770 ;
        RECT 100.800 150.650 101.525 150.820 ;
        RECT 101.695 150.650 101.965 151.620 ;
        RECT 99.380 149.910 99.730 150.480 ;
        RECT 99.900 150.150 100.610 150.600 ;
        RECT 101.355 150.480 101.525 150.650 ;
        RECT 100.780 150.150 101.185 150.480 ;
        RECT 101.355 150.150 101.625 150.480 ;
        RECT 101.355 149.980 101.525 150.150 ;
        RECT 99.915 149.810 101.525 149.980 ;
        RECT 101.795 149.915 101.965 150.650 ;
        RECT 102.135 150.700 104.725 151.790 ;
        RECT 102.135 150.180 103.345 150.700 ;
        RECT 104.935 150.650 105.165 151.790 ;
        RECT 105.335 150.640 105.665 151.620 ;
        RECT 105.835 150.650 106.045 151.790 ;
        RECT 106.650 151.110 106.905 151.480 ;
        RECT 106.565 150.940 106.905 151.110 ;
        RECT 107.085 150.990 107.370 151.790 ;
        RECT 107.550 151.070 107.880 151.580 ;
        RECT 106.650 150.810 106.905 150.940 ;
        RECT 103.515 150.010 104.725 150.530 ;
        RECT 104.915 150.230 105.245 150.480 ;
        RECT 93.860 149.240 99.205 149.785 ;
        RECT 99.385 149.240 99.715 149.740 ;
        RECT 99.915 149.460 100.085 149.810 ;
        RECT 100.285 149.240 100.615 149.640 ;
        RECT 100.785 149.460 100.955 149.810 ;
        RECT 101.125 149.240 101.505 149.640 ;
        RECT 101.695 149.570 101.965 149.915 ;
        RECT 102.135 149.240 104.725 150.010 ;
        RECT 104.935 149.240 105.165 150.060 ;
        RECT 105.415 150.040 105.665 150.640 ;
        RECT 105.335 149.410 105.665 150.040 ;
        RECT 105.835 149.240 106.045 150.060 ;
        RECT 106.650 149.950 106.830 150.810 ;
        RECT 107.550 150.480 107.800 151.070 ;
        RECT 108.150 150.920 108.320 151.530 ;
        RECT 108.490 151.100 108.820 151.790 ;
        RECT 109.050 151.240 109.290 151.530 ;
        RECT 109.490 151.410 109.910 151.790 ;
        RECT 110.090 151.320 110.720 151.570 ;
        RECT 111.190 151.410 111.520 151.790 ;
        RECT 110.090 151.240 110.260 151.320 ;
        RECT 111.690 151.240 111.860 151.530 ;
        RECT 112.040 151.410 112.420 151.790 ;
        RECT 112.660 151.405 113.490 151.575 ;
        RECT 109.050 151.070 110.260 151.240 ;
        RECT 107.000 150.150 107.800 150.480 ;
        RECT 106.650 149.420 106.905 149.950 ;
        RECT 107.085 149.240 107.370 149.700 ;
        RECT 107.550 149.500 107.800 150.150 ;
        RECT 108.000 150.900 108.320 150.920 ;
        RECT 108.000 150.730 109.920 150.900 ;
        RECT 108.000 149.835 108.190 150.730 ;
        RECT 110.090 150.560 110.260 151.070 ;
        RECT 110.430 150.810 110.950 151.120 ;
        RECT 108.360 150.390 110.260 150.560 ;
        RECT 108.360 150.330 108.690 150.390 ;
        RECT 108.840 150.160 109.170 150.220 ;
        RECT 108.510 149.890 109.170 150.160 ;
        RECT 108.000 149.505 108.320 149.835 ;
        RECT 108.500 149.240 109.160 149.720 ;
        RECT 109.360 149.630 109.530 150.390 ;
        RECT 110.430 150.220 110.610 150.630 ;
        RECT 109.700 150.050 110.030 150.170 ;
        RECT 110.780 150.050 110.950 150.810 ;
        RECT 109.700 149.880 110.950 150.050 ;
        RECT 111.120 150.990 112.490 151.240 ;
        RECT 111.120 150.220 111.310 150.990 ;
        RECT 112.240 150.730 112.490 150.990 ;
        RECT 111.480 150.560 111.730 150.720 ;
        RECT 112.660 150.560 112.830 151.405 ;
        RECT 113.725 151.120 113.895 151.620 ;
        RECT 114.065 151.290 114.395 151.790 ;
        RECT 113.000 150.730 113.500 151.110 ;
        RECT 113.725 150.950 114.420 151.120 ;
        RECT 111.480 150.390 112.830 150.560 ;
        RECT 112.410 150.350 112.830 150.390 ;
        RECT 111.120 149.880 111.540 150.220 ;
        RECT 111.830 149.890 112.240 150.220 ;
        RECT 109.360 149.460 110.210 149.630 ;
        RECT 110.770 149.240 111.090 149.700 ;
        RECT 111.290 149.450 111.540 149.880 ;
        RECT 111.830 149.240 112.240 149.680 ;
        RECT 112.410 149.620 112.580 150.350 ;
        RECT 112.750 149.800 113.100 150.170 ;
        RECT 113.280 149.860 113.500 150.730 ;
        RECT 113.670 150.160 114.080 150.780 ;
        RECT 114.250 149.980 114.420 150.950 ;
        RECT 113.725 149.790 114.420 149.980 ;
        RECT 112.410 149.420 113.425 149.620 ;
        RECT 113.725 149.460 113.895 149.790 ;
        RECT 114.065 149.240 114.395 149.620 ;
        RECT 114.610 149.500 114.835 151.620 ;
        RECT 115.005 151.290 115.335 151.790 ;
        RECT 115.505 151.120 115.675 151.620 ;
        RECT 115.010 150.950 115.675 151.120 ;
        RECT 115.010 149.960 115.240 150.950 ;
        RECT 115.410 150.130 115.760 150.780 ;
        RECT 115.935 150.715 116.205 151.620 ;
        RECT 116.375 151.030 116.705 151.790 ;
        RECT 116.885 150.860 117.055 151.620 ;
        RECT 115.010 149.790 115.675 149.960 ;
        RECT 115.005 149.240 115.335 149.620 ;
        RECT 115.505 149.500 115.675 149.790 ;
        RECT 115.935 149.915 116.105 150.715 ;
        RECT 116.390 150.690 117.055 150.860 ;
        RECT 117.315 150.700 118.525 151.790 ;
        RECT 116.390 150.545 116.560 150.690 ;
        RECT 116.275 150.215 116.560 150.545 ;
        RECT 116.390 149.960 116.560 150.215 ;
        RECT 116.795 150.140 117.125 150.510 ;
        RECT 117.315 150.160 117.835 150.700 ;
        RECT 118.005 149.990 118.525 150.530 ;
        RECT 115.935 149.410 116.195 149.915 ;
        RECT 116.390 149.790 117.055 149.960 ;
        RECT 116.375 149.240 116.705 149.620 ;
        RECT 116.885 149.410 117.055 149.790 ;
        RECT 117.315 149.240 118.525 149.990 ;
        RECT 11.430 149.070 118.610 149.240 ;
        RECT 11.515 148.320 12.725 149.070 ;
        RECT 13.820 148.360 14.075 148.890 ;
        RECT 14.245 148.610 14.550 149.070 ;
        RECT 14.795 148.690 15.865 148.860 ;
        RECT 11.515 147.780 12.035 148.320 ;
        RECT 12.205 147.610 12.725 148.150 ;
        RECT 11.515 146.520 12.725 147.610 ;
        RECT 13.820 147.710 14.030 148.360 ;
        RECT 14.795 148.335 15.115 148.690 ;
        RECT 14.790 148.160 15.115 148.335 ;
        RECT 14.200 147.860 15.115 148.160 ;
        RECT 15.285 148.120 15.525 148.520 ;
        RECT 15.695 148.460 15.865 148.690 ;
        RECT 16.035 148.630 16.225 149.070 ;
        RECT 16.395 148.620 17.345 148.900 ;
        RECT 17.565 148.710 17.915 148.880 ;
        RECT 15.695 148.290 16.225 148.460 ;
        RECT 14.200 147.830 14.940 147.860 ;
        RECT 13.820 146.830 14.075 147.710 ;
        RECT 14.245 146.520 14.550 147.660 ;
        RECT 14.770 147.240 14.940 147.830 ;
        RECT 15.285 147.750 15.825 148.120 ;
        RECT 16.005 148.010 16.225 148.290 ;
        RECT 16.395 147.840 16.565 148.620 ;
        RECT 16.160 147.670 16.565 147.840 ;
        RECT 16.735 147.830 17.085 148.450 ;
        RECT 16.160 147.580 16.330 147.670 ;
        RECT 17.255 147.660 17.465 148.450 ;
        RECT 15.110 147.410 16.330 147.580 ;
        RECT 16.790 147.500 17.465 147.660 ;
        RECT 14.770 147.070 15.570 147.240 ;
        RECT 14.890 146.520 15.220 146.900 ;
        RECT 15.400 146.780 15.570 147.070 ;
        RECT 16.160 147.030 16.330 147.410 ;
        RECT 16.500 147.490 17.465 147.500 ;
        RECT 17.655 148.320 17.915 148.710 ;
        RECT 18.125 148.610 18.455 149.070 ;
        RECT 19.330 148.680 20.185 148.850 ;
        RECT 20.390 148.680 20.885 148.850 ;
        RECT 21.055 148.710 21.385 149.070 ;
        RECT 17.655 147.630 17.825 148.320 ;
        RECT 17.995 147.970 18.165 148.150 ;
        RECT 18.335 148.140 19.125 148.390 ;
        RECT 19.330 147.970 19.500 148.680 ;
        RECT 19.670 148.170 20.025 148.390 ;
        RECT 17.995 147.800 19.685 147.970 ;
        RECT 16.500 147.200 16.960 147.490 ;
        RECT 17.655 147.460 19.155 147.630 ;
        RECT 17.655 147.320 17.825 147.460 ;
        RECT 17.265 147.150 17.825 147.320 ;
        RECT 15.740 146.520 15.990 146.980 ;
        RECT 16.160 146.690 17.030 147.030 ;
        RECT 17.265 146.690 17.435 147.150 ;
        RECT 18.270 147.120 19.345 147.290 ;
        RECT 17.605 146.520 17.975 146.980 ;
        RECT 18.270 146.780 18.440 147.120 ;
        RECT 18.610 146.520 18.940 146.950 ;
        RECT 19.175 146.780 19.345 147.120 ;
        RECT 19.515 147.020 19.685 147.800 ;
        RECT 19.855 147.580 20.025 148.170 ;
        RECT 20.195 147.770 20.545 148.390 ;
        RECT 19.855 147.190 20.320 147.580 ;
        RECT 20.715 147.320 20.885 148.680 ;
        RECT 21.055 147.490 21.515 148.540 ;
        RECT 20.490 147.150 20.885 147.320 ;
        RECT 20.490 147.020 20.660 147.150 ;
        RECT 19.515 146.690 20.195 147.020 ;
        RECT 20.410 146.690 20.660 147.020 ;
        RECT 20.830 146.520 21.080 146.980 ;
        RECT 21.250 146.705 21.575 147.490 ;
        RECT 21.745 146.690 21.915 148.810 ;
        RECT 22.085 148.690 22.415 149.070 ;
        RECT 22.585 148.520 22.840 148.810 ;
        RECT 22.090 148.350 22.840 148.520 ;
        RECT 22.090 147.360 22.320 148.350 ;
        RECT 23.480 148.330 23.735 148.900 ;
        RECT 23.905 148.670 24.235 149.070 ;
        RECT 24.660 148.535 25.190 148.900 ;
        RECT 25.380 148.730 25.655 148.900 ;
        RECT 25.375 148.560 25.655 148.730 ;
        RECT 24.660 148.500 24.835 148.535 ;
        RECT 23.905 148.330 24.835 148.500 ;
        RECT 22.490 147.530 22.840 148.180 ;
        RECT 23.480 147.660 23.650 148.330 ;
        RECT 23.905 148.160 24.075 148.330 ;
        RECT 23.820 147.830 24.075 148.160 ;
        RECT 24.300 147.830 24.495 148.160 ;
        RECT 22.090 147.190 22.840 147.360 ;
        RECT 22.085 146.520 22.415 147.020 ;
        RECT 22.585 146.690 22.840 147.190 ;
        RECT 23.480 146.690 23.815 147.660 ;
        RECT 23.985 146.520 24.155 147.660 ;
        RECT 24.325 146.860 24.495 147.830 ;
        RECT 24.665 147.200 24.835 148.330 ;
        RECT 25.005 147.540 25.175 148.340 ;
        RECT 25.380 147.740 25.655 148.560 ;
        RECT 25.825 147.540 26.015 148.900 ;
        RECT 26.195 148.535 26.705 149.070 ;
        RECT 26.925 148.260 27.170 148.865 ;
        RECT 28.075 148.345 28.365 149.070 ;
        RECT 28.535 148.320 29.745 149.070 ;
        RECT 30.005 148.520 30.175 148.900 ;
        RECT 30.355 148.690 30.685 149.070 ;
        RECT 30.005 148.350 30.670 148.520 ;
        RECT 30.865 148.395 31.125 148.900 ;
        RECT 26.215 148.090 27.445 148.260 ;
        RECT 25.005 147.370 26.015 147.540 ;
        RECT 26.185 147.525 26.935 147.715 ;
        RECT 24.665 147.030 25.790 147.200 ;
        RECT 26.185 146.860 26.355 147.525 ;
        RECT 27.105 147.280 27.445 148.090 ;
        RECT 24.325 146.690 26.355 146.860 ;
        RECT 26.525 146.520 26.695 147.280 ;
        RECT 26.930 146.870 27.445 147.280 ;
        RECT 28.075 146.520 28.365 147.685 ;
        RECT 28.535 147.610 29.055 148.150 ;
        RECT 29.225 147.780 29.745 148.320 ;
        RECT 29.935 147.800 30.265 148.170 ;
        RECT 30.500 148.095 30.670 148.350 ;
        RECT 30.500 147.765 30.785 148.095 ;
        RECT 30.500 147.620 30.670 147.765 ;
        RECT 28.535 146.520 29.745 147.610 ;
        RECT 30.005 147.450 30.670 147.620 ;
        RECT 30.955 147.595 31.125 148.395 ;
        RECT 31.500 148.290 32.000 148.900 ;
        RECT 31.295 147.830 31.645 148.080 ;
        RECT 31.830 147.660 32.000 148.290 ;
        RECT 32.630 148.420 32.960 148.900 ;
        RECT 33.130 148.610 33.355 149.070 ;
        RECT 33.525 148.420 33.855 148.900 ;
        RECT 32.630 148.250 33.855 148.420 ;
        RECT 34.045 148.270 34.295 149.070 ;
        RECT 34.465 148.270 34.805 148.900 ;
        RECT 35.180 148.290 35.680 148.900 ;
        RECT 32.170 147.880 32.500 148.080 ;
        RECT 32.670 147.880 33.000 148.080 ;
        RECT 33.170 147.880 33.590 148.080 ;
        RECT 33.765 147.910 34.460 148.080 ;
        RECT 33.765 147.660 33.935 147.910 ;
        RECT 34.630 147.660 34.805 148.270 ;
        RECT 34.975 147.830 35.325 148.080 ;
        RECT 35.510 147.660 35.680 148.290 ;
        RECT 36.310 148.420 36.640 148.900 ;
        RECT 36.810 148.610 37.035 149.070 ;
        RECT 37.205 148.420 37.535 148.900 ;
        RECT 36.310 148.250 37.535 148.420 ;
        RECT 37.725 148.270 37.975 149.070 ;
        RECT 38.145 148.270 38.485 148.900 ;
        RECT 38.655 148.300 40.325 149.070 ;
        RECT 35.850 147.880 36.180 148.080 ;
        RECT 36.350 147.880 36.680 148.080 ;
        RECT 36.850 147.880 37.270 148.080 ;
        RECT 37.445 147.910 38.140 148.080 ;
        RECT 37.445 147.660 37.615 147.910 ;
        RECT 38.310 147.660 38.485 148.270 ;
        RECT 30.005 146.690 30.175 147.450 ;
        RECT 30.355 146.520 30.685 147.280 ;
        RECT 30.855 146.690 31.125 147.595 ;
        RECT 31.500 147.490 33.935 147.660 ;
        RECT 31.500 146.690 31.830 147.490 ;
        RECT 32.000 146.520 32.330 147.320 ;
        RECT 32.630 146.690 32.960 147.490 ;
        RECT 33.605 146.520 33.855 147.320 ;
        RECT 34.125 146.520 34.295 147.660 ;
        RECT 34.465 146.690 34.805 147.660 ;
        RECT 35.180 147.490 37.615 147.660 ;
        RECT 35.180 146.690 35.510 147.490 ;
        RECT 35.680 146.520 36.010 147.320 ;
        RECT 36.310 146.690 36.640 147.490 ;
        RECT 37.285 146.520 37.535 147.320 ;
        RECT 37.805 146.520 37.975 147.660 ;
        RECT 38.145 146.690 38.485 147.660 ;
        RECT 38.655 147.610 39.405 148.130 ;
        RECT 39.575 147.780 40.325 148.300 ;
        RECT 40.495 148.270 40.835 148.900 ;
        RECT 41.005 148.270 41.255 149.070 ;
        RECT 41.445 148.420 41.775 148.900 ;
        RECT 41.945 148.610 42.170 149.070 ;
        RECT 42.340 148.420 42.670 148.900 ;
        RECT 40.495 147.660 40.670 148.270 ;
        RECT 41.445 148.250 42.670 148.420 ;
        RECT 43.300 148.290 43.800 148.900 ;
        RECT 44.550 148.360 44.805 148.890 ;
        RECT 44.985 148.610 45.270 149.070 ;
        RECT 40.840 147.910 41.535 148.080 ;
        RECT 41.365 147.660 41.535 147.910 ;
        RECT 41.710 147.880 42.130 148.080 ;
        RECT 42.300 147.880 42.630 148.080 ;
        RECT 42.800 147.880 43.130 148.080 ;
        RECT 43.300 147.660 43.470 148.290 ;
        RECT 43.655 147.830 44.005 148.080 ;
        RECT 38.655 146.520 40.325 147.610 ;
        RECT 40.495 146.690 40.835 147.660 ;
        RECT 41.005 146.520 41.175 147.660 ;
        RECT 41.365 147.490 43.800 147.660 ;
        RECT 41.445 146.520 41.695 147.320 ;
        RECT 42.340 146.690 42.670 147.490 ;
        RECT 42.970 146.520 43.300 147.320 ;
        RECT 43.470 146.690 43.800 147.490 ;
        RECT 44.550 147.500 44.730 148.360 ;
        RECT 45.450 148.160 45.700 148.810 ;
        RECT 44.900 147.830 45.700 148.160 ;
        RECT 44.550 147.030 44.805 147.500 ;
        RECT 44.465 146.860 44.805 147.030 ;
        RECT 44.550 146.830 44.805 146.860 ;
        RECT 44.985 146.520 45.270 147.320 ;
        RECT 45.450 147.240 45.700 147.830 ;
        RECT 45.900 148.475 46.220 148.805 ;
        RECT 46.400 148.590 47.060 149.070 ;
        RECT 47.260 148.680 48.110 148.850 ;
        RECT 45.900 147.580 46.090 148.475 ;
        RECT 46.410 148.150 47.070 148.420 ;
        RECT 46.740 148.090 47.070 148.150 ;
        RECT 46.260 147.920 46.590 147.980 ;
        RECT 47.260 147.920 47.430 148.680 ;
        RECT 48.670 148.610 48.990 149.070 ;
        RECT 49.190 148.430 49.440 148.860 ;
        RECT 49.730 148.630 50.140 149.070 ;
        RECT 50.310 148.690 51.325 148.890 ;
        RECT 47.600 148.260 48.850 148.430 ;
        RECT 47.600 148.140 47.930 148.260 ;
        RECT 46.260 147.750 48.160 147.920 ;
        RECT 45.900 147.410 47.820 147.580 ;
        RECT 45.900 147.390 46.220 147.410 ;
        RECT 45.450 146.730 45.780 147.240 ;
        RECT 46.050 146.780 46.220 147.390 ;
        RECT 47.990 147.240 48.160 147.750 ;
        RECT 48.330 147.680 48.510 148.090 ;
        RECT 48.680 147.500 48.850 148.260 ;
        RECT 46.390 146.520 46.720 147.210 ;
        RECT 46.950 147.070 48.160 147.240 ;
        RECT 48.330 147.190 48.850 147.500 ;
        RECT 49.020 148.090 49.440 148.430 ;
        RECT 49.730 148.090 50.140 148.420 ;
        RECT 49.020 147.320 49.210 148.090 ;
        RECT 50.310 147.960 50.480 148.690 ;
        RECT 51.625 148.520 51.795 148.850 ;
        RECT 51.965 148.690 52.295 149.070 ;
        RECT 50.650 148.140 51.000 148.510 ;
        RECT 50.310 147.920 50.730 147.960 ;
        RECT 49.380 147.750 50.730 147.920 ;
        RECT 49.380 147.590 49.630 147.750 ;
        RECT 50.140 147.320 50.390 147.580 ;
        RECT 49.020 147.070 50.390 147.320 ;
        RECT 46.950 146.780 47.190 147.070 ;
        RECT 47.990 146.990 48.160 147.070 ;
        RECT 47.390 146.520 47.810 146.900 ;
        RECT 47.990 146.740 48.620 146.990 ;
        RECT 49.090 146.520 49.420 146.900 ;
        RECT 49.590 146.780 49.760 147.070 ;
        RECT 50.560 146.905 50.730 147.750 ;
        RECT 51.180 147.580 51.400 148.450 ;
        RECT 51.625 148.330 52.320 148.520 ;
        RECT 50.900 147.200 51.400 147.580 ;
        RECT 51.570 147.530 51.980 148.150 ;
        RECT 52.150 147.360 52.320 148.330 ;
        RECT 51.625 147.190 52.320 147.360 ;
        RECT 49.940 146.520 50.320 146.900 ;
        RECT 50.560 146.735 51.390 146.905 ;
        RECT 51.625 146.690 51.795 147.190 ;
        RECT 51.965 146.520 52.295 147.020 ;
        RECT 52.510 146.690 52.735 148.810 ;
        RECT 52.905 148.690 53.235 149.070 ;
        RECT 53.405 148.520 53.575 148.810 ;
        RECT 52.910 148.350 53.575 148.520 ;
        RECT 52.910 147.360 53.140 148.350 ;
        RECT 53.835 148.345 54.125 149.070 ;
        RECT 54.295 148.395 54.555 148.900 ;
        RECT 54.735 148.690 55.065 149.070 ;
        RECT 55.245 148.520 55.415 148.900 ;
        RECT 53.310 147.530 53.660 148.180 ;
        RECT 52.910 147.190 53.575 147.360 ;
        RECT 52.905 146.520 53.235 147.020 ;
        RECT 53.405 146.690 53.575 147.190 ;
        RECT 53.835 146.520 54.125 147.685 ;
        RECT 54.295 147.595 54.465 148.395 ;
        RECT 54.750 148.350 55.415 148.520 ;
        RECT 54.750 148.095 54.920 148.350 ;
        RECT 55.675 148.300 57.345 149.070 ;
        RECT 54.635 147.765 54.920 148.095 ;
        RECT 55.155 147.800 55.485 148.170 ;
        RECT 54.750 147.620 54.920 147.765 ;
        RECT 54.295 146.690 54.565 147.595 ;
        RECT 54.750 147.450 55.415 147.620 ;
        RECT 54.735 146.520 55.065 147.280 ;
        RECT 55.245 146.690 55.415 147.450 ;
        RECT 55.675 147.610 56.425 148.130 ;
        RECT 56.595 147.780 57.345 148.300 ;
        RECT 57.555 148.250 57.785 149.070 ;
        RECT 57.955 148.270 58.285 148.900 ;
        RECT 57.535 147.830 57.865 148.080 ;
        RECT 58.035 147.670 58.285 148.270 ;
        RECT 58.455 148.250 58.665 149.070 ;
        RECT 59.820 148.525 65.165 149.070 ;
        RECT 55.675 146.520 57.345 147.610 ;
        RECT 57.555 146.520 57.785 147.660 ;
        RECT 57.955 146.690 58.285 147.670 ;
        RECT 58.455 146.520 58.665 147.660 ;
        RECT 61.410 146.955 61.760 148.205 ;
        RECT 63.240 147.695 63.580 148.525 ;
        RECT 65.335 148.395 65.595 148.900 ;
        RECT 65.775 148.690 66.105 149.070 ;
        RECT 66.285 148.520 66.455 148.900 ;
        RECT 66.720 148.525 72.065 149.070 ;
        RECT 65.335 147.595 65.515 148.395 ;
        RECT 65.790 148.350 66.455 148.520 ;
        RECT 65.790 148.095 65.960 148.350 ;
        RECT 65.685 147.765 65.960 148.095 ;
        RECT 66.185 147.800 66.525 148.170 ;
        RECT 65.790 147.620 65.960 147.765 ;
        RECT 59.820 146.520 65.165 146.955 ;
        RECT 65.335 146.690 65.605 147.595 ;
        RECT 65.790 147.450 66.465 147.620 ;
        RECT 65.775 146.520 66.105 147.280 ;
        RECT 66.285 146.690 66.465 147.450 ;
        RECT 68.310 146.955 68.660 148.205 ;
        RECT 70.140 147.695 70.480 148.525 ;
        RECT 72.235 148.395 72.505 148.740 ;
        RECT 72.695 148.670 73.075 149.070 ;
        RECT 73.245 148.500 73.415 148.850 ;
        RECT 73.585 148.670 73.915 149.070 ;
        RECT 74.115 148.500 74.285 148.850 ;
        RECT 74.485 148.570 74.815 149.070 ;
        RECT 72.235 147.660 72.405 148.395 ;
        RECT 72.675 148.330 74.285 148.500 ;
        RECT 72.675 148.160 72.845 148.330 ;
        RECT 72.575 147.830 72.845 148.160 ;
        RECT 73.015 147.830 73.420 148.160 ;
        RECT 72.675 147.660 72.845 147.830 ;
        RECT 73.590 147.710 74.300 148.160 ;
        RECT 74.470 147.830 74.820 148.400 ;
        RECT 75.915 148.300 79.425 149.070 ;
        RECT 79.595 148.345 79.885 149.070 ;
        RECT 81.350 148.360 81.605 148.890 ;
        RECT 81.785 148.610 82.070 149.070 ;
        RECT 66.720 146.520 72.065 146.955 ;
        RECT 72.235 146.690 72.505 147.660 ;
        RECT 72.675 147.490 73.400 147.660 ;
        RECT 73.590 147.540 74.305 147.710 ;
        RECT 73.230 147.370 73.400 147.490 ;
        RECT 74.500 147.370 74.820 147.660 ;
        RECT 72.715 146.520 72.995 147.320 ;
        RECT 73.230 147.200 74.820 147.370 ;
        RECT 75.915 147.610 77.605 148.130 ;
        RECT 77.775 147.780 79.425 148.300 ;
        RECT 73.165 146.740 74.820 147.030 ;
        RECT 75.915 146.520 79.425 147.610 ;
        RECT 79.595 146.520 79.885 147.685 ;
        RECT 81.350 147.500 81.530 148.360 ;
        RECT 82.250 148.160 82.500 148.810 ;
        RECT 81.700 147.830 82.500 148.160 ;
        RECT 81.350 147.370 81.605 147.500 ;
        RECT 81.265 147.200 81.605 147.370 ;
        RECT 81.350 146.830 81.605 147.200 ;
        RECT 81.785 146.520 82.070 147.320 ;
        RECT 82.250 147.240 82.500 147.830 ;
        RECT 82.700 148.475 83.020 148.805 ;
        RECT 83.200 148.590 83.860 149.070 ;
        RECT 84.060 148.680 84.910 148.850 ;
        RECT 82.700 147.580 82.890 148.475 ;
        RECT 83.210 148.150 83.870 148.420 ;
        RECT 83.540 148.090 83.870 148.150 ;
        RECT 83.060 147.920 83.390 147.980 ;
        RECT 84.060 147.920 84.230 148.680 ;
        RECT 85.470 148.610 85.790 149.070 ;
        RECT 85.990 148.430 86.240 148.860 ;
        RECT 86.530 148.630 86.940 149.070 ;
        RECT 87.110 148.690 88.125 148.890 ;
        RECT 84.400 148.260 85.650 148.430 ;
        RECT 84.400 148.140 84.730 148.260 ;
        RECT 83.060 147.750 84.960 147.920 ;
        RECT 82.700 147.410 84.620 147.580 ;
        RECT 82.700 147.390 83.020 147.410 ;
        RECT 82.250 146.730 82.580 147.240 ;
        RECT 82.850 146.780 83.020 147.390 ;
        RECT 84.790 147.240 84.960 147.750 ;
        RECT 85.130 147.680 85.310 148.090 ;
        RECT 85.480 147.500 85.650 148.260 ;
        RECT 83.190 146.520 83.520 147.210 ;
        RECT 83.750 147.070 84.960 147.240 ;
        RECT 85.130 147.190 85.650 147.500 ;
        RECT 85.820 148.090 86.240 148.430 ;
        RECT 86.530 148.090 86.940 148.420 ;
        RECT 85.820 147.320 86.010 148.090 ;
        RECT 87.110 147.960 87.280 148.690 ;
        RECT 88.425 148.520 88.595 148.850 ;
        RECT 88.765 148.690 89.095 149.070 ;
        RECT 87.450 148.140 87.800 148.510 ;
        RECT 87.110 147.920 87.530 147.960 ;
        RECT 86.180 147.750 87.530 147.920 ;
        RECT 86.180 147.590 86.430 147.750 ;
        RECT 86.940 147.320 87.190 147.580 ;
        RECT 85.820 147.070 87.190 147.320 ;
        RECT 83.750 146.780 83.990 147.070 ;
        RECT 84.790 146.990 84.960 147.070 ;
        RECT 84.190 146.520 84.610 146.900 ;
        RECT 84.790 146.740 85.420 146.990 ;
        RECT 85.890 146.520 86.220 146.900 ;
        RECT 86.390 146.780 86.560 147.070 ;
        RECT 87.360 146.905 87.530 147.750 ;
        RECT 87.980 147.580 88.200 148.450 ;
        RECT 88.425 148.330 89.120 148.520 ;
        RECT 87.700 147.200 88.200 147.580 ;
        RECT 88.370 147.530 88.780 148.150 ;
        RECT 88.950 147.360 89.120 148.330 ;
        RECT 88.425 147.190 89.120 147.360 ;
        RECT 86.740 146.520 87.120 146.900 ;
        RECT 87.360 146.735 88.190 146.905 ;
        RECT 88.425 146.690 88.595 147.190 ;
        RECT 88.765 146.520 89.095 147.020 ;
        RECT 89.310 146.690 89.535 148.810 ;
        RECT 89.705 148.690 90.035 149.070 ;
        RECT 90.205 148.520 90.375 148.810 ;
        RECT 89.710 148.350 90.375 148.520 ;
        RECT 89.710 147.360 89.940 148.350 ;
        RECT 90.635 148.300 94.145 149.070 ;
        RECT 90.110 147.530 90.460 148.180 ;
        RECT 90.635 147.610 92.325 148.130 ;
        RECT 92.495 147.780 94.145 148.300 ;
        RECT 94.590 148.260 94.835 148.865 ;
        RECT 95.055 148.535 95.565 149.070 ;
        RECT 94.315 148.090 95.545 148.260 ;
        RECT 89.710 147.190 90.375 147.360 ;
        RECT 89.705 146.520 90.035 147.020 ;
        RECT 90.205 146.690 90.375 147.190 ;
        RECT 90.635 146.520 94.145 147.610 ;
        RECT 94.315 147.280 94.655 148.090 ;
        RECT 94.825 147.525 95.575 147.715 ;
        RECT 94.315 146.870 94.830 147.280 ;
        RECT 95.065 146.520 95.235 147.280 ;
        RECT 95.405 146.860 95.575 147.525 ;
        RECT 95.745 147.540 95.935 148.900 ;
        RECT 96.105 148.730 96.380 148.900 ;
        RECT 96.105 148.560 96.385 148.730 ;
        RECT 96.105 147.740 96.380 148.560 ;
        RECT 96.570 148.535 97.100 148.900 ;
        RECT 97.525 148.670 97.855 149.070 ;
        RECT 96.925 148.500 97.100 148.535 ;
        RECT 96.585 147.540 96.755 148.340 ;
        RECT 95.745 147.370 96.755 147.540 ;
        RECT 96.925 148.330 97.855 148.500 ;
        RECT 98.025 148.330 98.280 148.900 ;
        RECT 96.925 147.200 97.095 148.330 ;
        RECT 97.685 148.160 97.855 148.330 ;
        RECT 95.970 147.030 97.095 147.200 ;
        RECT 97.265 147.830 97.460 148.160 ;
        RECT 97.685 147.830 97.940 148.160 ;
        RECT 97.265 146.860 97.435 147.830 ;
        RECT 98.110 147.660 98.280 148.330 ;
        RECT 98.730 148.260 98.975 148.865 ;
        RECT 99.195 148.535 99.705 149.070 ;
        RECT 95.405 146.690 97.435 146.860 ;
        RECT 97.605 146.520 97.775 147.660 ;
        RECT 97.945 146.690 98.280 147.660 ;
        RECT 98.455 148.090 99.685 148.260 ;
        RECT 98.455 147.280 98.795 148.090 ;
        RECT 98.965 147.525 99.715 147.715 ;
        RECT 98.455 146.870 98.970 147.280 ;
        RECT 99.205 146.520 99.375 147.280 ;
        RECT 99.545 146.860 99.715 147.525 ;
        RECT 99.885 147.540 100.075 148.900 ;
        RECT 100.245 148.390 100.520 148.900 ;
        RECT 100.710 148.535 101.240 148.900 ;
        RECT 101.665 148.670 101.995 149.070 ;
        RECT 101.065 148.500 101.240 148.535 ;
        RECT 100.245 148.220 100.525 148.390 ;
        RECT 100.245 147.740 100.520 148.220 ;
        RECT 100.725 147.540 100.895 148.340 ;
        RECT 99.885 147.370 100.895 147.540 ;
        RECT 101.065 148.330 101.995 148.500 ;
        RECT 102.165 148.330 102.420 148.900 ;
        RECT 101.065 147.200 101.235 148.330 ;
        RECT 101.825 148.160 101.995 148.330 ;
        RECT 100.110 147.030 101.235 147.200 ;
        RECT 101.405 147.830 101.600 148.160 ;
        RECT 101.825 147.830 102.080 148.160 ;
        RECT 101.405 146.860 101.575 147.830 ;
        RECT 102.250 147.660 102.420 148.330 ;
        RECT 102.595 148.300 105.185 149.070 ;
        RECT 105.355 148.345 105.645 149.070 ;
        RECT 99.545 146.690 101.575 146.860 ;
        RECT 101.745 146.520 101.915 147.660 ;
        RECT 102.085 146.690 102.420 147.660 ;
        RECT 102.595 147.610 103.805 148.130 ;
        RECT 103.975 147.780 105.185 148.300 ;
        RECT 106.315 148.250 106.545 149.070 ;
        RECT 106.715 148.270 107.045 148.900 ;
        RECT 106.295 147.830 106.625 148.080 ;
        RECT 102.595 146.520 105.185 147.610 ;
        RECT 105.355 146.520 105.645 147.685 ;
        RECT 106.795 147.670 107.045 148.270 ;
        RECT 107.215 148.250 107.425 149.070 ;
        RECT 108.030 148.730 108.285 148.890 ;
        RECT 107.945 148.560 108.285 148.730 ;
        RECT 108.465 148.610 108.750 149.070 ;
        RECT 108.030 148.360 108.285 148.560 ;
        RECT 106.315 146.520 106.545 147.660 ;
        RECT 106.715 146.690 107.045 147.670 ;
        RECT 107.215 146.520 107.425 147.660 ;
        RECT 108.030 147.500 108.210 148.360 ;
        RECT 108.930 148.160 109.180 148.810 ;
        RECT 108.380 147.830 109.180 148.160 ;
        RECT 108.030 146.830 108.285 147.500 ;
        RECT 108.465 146.520 108.750 147.320 ;
        RECT 108.930 147.240 109.180 147.830 ;
        RECT 109.380 148.475 109.700 148.805 ;
        RECT 109.880 148.590 110.540 149.070 ;
        RECT 110.740 148.680 111.590 148.850 ;
        RECT 109.380 147.580 109.570 148.475 ;
        RECT 109.890 148.150 110.550 148.420 ;
        RECT 110.220 148.090 110.550 148.150 ;
        RECT 109.740 147.920 110.070 147.980 ;
        RECT 110.740 147.920 110.910 148.680 ;
        RECT 112.150 148.610 112.470 149.070 ;
        RECT 112.670 148.430 112.920 148.860 ;
        RECT 113.210 148.630 113.620 149.070 ;
        RECT 113.790 148.690 114.805 148.890 ;
        RECT 111.080 148.260 112.330 148.430 ;
        RECT 111.080 148.140 111.410 148.260 ;
        RECT 109.740 147.750 111.640 147.920 ;
        RECT 109.380 147.410 111.300 147.580 ;
        RECT 109.380 147.390 109.700 147.410 ;
        RECT 108.930 146.730 109.260 147.240 ;
        RECT 109.530 146.780 109.700 147.390 ;
        RECT 111.470 147.240 111.640 147.750 ;
        RECT 111.810 147.680 111.990 148.090 ;
        RECT 112.160 147.500 112.330 148.260 ;
        RECT 109.870 146.520 110.200 147.210 ;
        RECT 110.430 147.070 111.640 147.240 ;
        RECT 111.810 147.190 112.330 147.500 ;
        RECT 112.500 148.090 112.920 148.430 ;
        RECT 113.210 148.090 113.620 148.420 ;
        RECT 112.500 147.320 112.690 148.090 ;
        RECT 113.790 147.960 113.960 148.690 ;
        RECT 115.105 148.520 115.275 148.850 ;
        RECT 115.445 148.690 115.775 149.070 ;
        RECT 114.130 148.140 114.480 148.510 ;
        RECT 113.790 147.920 114.210 147.960 ;
        RECT 112.860 147.750 114.210 147.920 ;
        RECT 112.860 147.590 113.110 147.750 ;
        RECT 113.620 147.320 113.870 147.580 ;
        RECT 112.500 147.070 113.870 147.320 ;
        RECT 110.430 146.780 110.670 147.070 ;
        RECT 111.470 146.990 111.640 147.070 ;
        RECT 110.870 146.520 111.290 146.900 ;
        RECT 111.470 146.740 112.100 146.990 ;
        RECT 112.570 146.520 112.900 146.900 ;
        RECT 113.070 146.780 113.240 147.070 ;
        RECT 114.040 146.905 114.210 147.750 ;
        RECT 114.660 147.580 114.880 148.450 ;
        RECT 115.105 148.330 115.800 148.520 ;
        RECT 114.380 147.200 114.880 147.580 ;
        RECT 115.050 147.530 115.460 148.150 ;
        RECT 115.630 147.360 115.800 148.330 ;
        RECT 115.105 147.190 115.800 147.360 ;
        RECT 113.420 146.520 113.800 146.900 ;
        RECT 114.040 146.735 114.870 146.905 ;
        RECT 115.105 146.690 115.275 147.190 ;
        RECT 115.445 146.520 115.775 147.020 ;
        RECT 115.990 146.690 116.215 148.810 ;
        RECT 116.385 148.690 116.715 149.070 ;
        RECT 116.885 148.520 117.055 148.810 ;
        RECT 116.390 148.350 117.055 148.520 ;
        RECT 116.390 147.360 116.620 148.350 ;
        RECT 117.315 148.320 118.525 149.070 ;
        RECT 116.790 147.530 117.140 148.180 ;
        RECT 117.315 147.610 117.835 148.150 ;
        RECT 118.005 147.780 118.525 148.320 ;
        RECT 116.390 147.190 117.055 147.360 ;
        RECT 116.385 146.520 116.715 147.020 ;
        RECT 116.885 146.690 117.055 147.190 ;
        RECT 117.315 146.520 118.525 147.610 ;
        RECT 11.430 146.350 118.610 146.520 ;
        RECT 11.515 145.260 12.725 146.350 ;
        RECT 11.515 144.550 12.035 145.090 ;
        RECT 12.205 144.720 12.725 145.260 ;
        RECT 13.875 145.210 14.085 146.350 ;
        RECT 14.255 145.200 14.585 146.180 ;
        RECT 14.755 145.210 14.985 146.350 ;
        RECT 11.515 143.800 12.725 144.550 ;
        RECT 13.875 143.800 14.085 144.620 ;
        RECT 14.255 144.600 14.505 145.200 ;
        RECT 15.195 145.185 15.485 146.350 ;
        RECT 15.695 145.210 15.925 146.350 ;
        RECT 16.095 145.200 16.425 146.180 ;
        RECT 16.595 145.210 16.805 146.350 ;
        RECT 17.125 145.420 17.295 146.180 ;
        RECT 17.475 145.590 17.805 146.350 ;
        RECT 17.125 145.250 17.790 145.420 ;
        RECT 17.975 145.275 18.245 146.180 ;
        RECT 14.675 144.790 15.005 145.040 ;
        RECT 15.675 144.790 16.005 145.040 ;
        RECT 14.255 143.970 14.585 144.600 ;
        RECT 14.755 143.800 14.985 144.620 ;
        RECT 15.195 143.800 15.485 144.525 ;
        RECT 15.695 143.800 15.925 144.620 ;
        RECT 16.175 144.600 16.425 145.200 ;
        RECT 17.620 145.105 17.790 145.250 ;
        RECT 17.055 144.700 17.385 145.070 ;
        RECT 17.620 144.775 17.905 145.105 ;
        RECT 16.095 143.970 16.425 144.600 ;
        RECT 16.595 143.800 16.805 144.620 ;
        RECT 17.620 144.520 17.790 144.775 ;
        RECT 17.125 144.350 17.790 144.520 ;
        RECT 18.075 144.475 18.245 145.275 ;
        RECT 17.125 143.970 17.295 144.350 ;
        RECT 17.475 143.800 17.805 144.180 ;
        RECT 17.985 143.970 18.245 144.475 ;
        RECT 18.420 145.160 18.675 146.040 ;
        RECT 18.845 145.210 19.150 146.350 ;
        RECT 19.490 145.970 19.820 146.350 ;
        RECT 20.000 145.800 20.170 146.090 ;
        RECT 20.340 145.890 20.590 146.350 ;
        RECT 19.370 145.630 20.170 145.800 ;
        RECT 20.760 145.840 21.630 146.180 ;
        RECT 18.420 144.510 18.630 145.160 ;
        RECT 19.370 145.040 19.540 145.630 ;
        RECT 20.760 145.460 20.930 145.840 ;
        RECT 21.865 145.720 22.035 146.180 ;
        RECT 22.205 145.890 22.575 146.350 ;
        RECT 22.870 145.750 23.040 146.090 ;
        RECT 23.210 145.920 23.540 146.350 ;
        RECT 23.775 145.750 23.945 146.090 ;
        RECT 19.710 145.290 20.930 145.460 ;
        RECT 21.100 145.380 21.560 145.670 ;
        RECT 21.865 145.550 22.425 145.720 ;
        RECT 22.870 145.580 23.945 145.750 ;
        RECT 24.115 145.850 24.795 146.180 ;
        RECT 25.010 145.850 25.260 146.180 ;
        RECT 25.430 145.890 25.680 146.350 ;
        RECT 22.255 145.410 22.425 145.550 ;
        RECT 21.100 145.370 22.065 145.380 ;
        RECT 20.760 145.200 20.930 145.290 ;
        RECT 21.390 145.210 22.065 145.370 ;
        RECT 18.800 145.010 19.540 145.040 ;
        RECT 18.800 144.710 19.715 145.010 ;
        RECT 19.390 144.535 19.715 144.710 ;
        RECT 18.420 143.980 18.675 144.510 ;
        RECT 18.845 143.800 19.150 144.260 ;
        RECT 19.395 144.180 19.715 144.535 ;
        RECT 19.885 144.750 20.425 145.120 ;
        RECT 20.760 145.030 21.165 145.200 ;
        RECT 19.885 144.350 20.125 144.750 ;
        RECT 20.605 144.580 20.825 144.860 ;
        RECT 20.295 144.410 20.825 144.580 ;
        RECT 20.295 144.180 20.465 144.410 ;
        RECT 20.995 144.250 21.165 145.030 ;
        RECT 21.335 144.420 21.685 145.040 ;
        RECT 21.855 144.420 22.065 145.210 ;
        RECT 22.255 145.240 23.755 145.410 ;
        RECT 22.255 144.550 22.425 145.240 ;
        RECT 24.115 145.070 24.285 145.850 ;
        RECT 25.090 145.720 25.260 145.850 ;
        RECT 22.595 144.900 24.285 145.070 ;
        RECT 24.455 145.290 24.920 145.680 ;
        RECT 25.090 145.550 25.485 145.720 ;
        RECT 22.595 144.720 22.765 144.900 ;
        RECT 19.395 144.010 20.465 144.180 ;
        RECT 20.635 143.800 20.825 144.240 ;
        RECT 20.995 143.970 21.945 144.250 ;
        RECT 22.255 144.160 22.515 144.550 ;
        RECT 22.935 144.480 23.725 144.730 ;
        RECT 22.165 143.990 22.515 144.160 ;
        RECT 22.725 143.800 23.055 144.260 ;
        RECT 23.930 144.190 24.100 144.900 ;
        RECT 24.455 144.700 24.625 145.290 ;
        RECT 24.270 144.480 24.625 144.700 ;
        RECT 24.795 144.480 25.145 145.100 ;
        RECT 25.315 144.190 25.485 145.550 ;
        RECT 25.850 145.380 26.175 146.165 ;
        RECT 25.655 144.330 26.115 145.380 ;
        RECT 23.930 144.020 24.785 144.190 ;
        RECT 24.990 144.020 25.485 144.190 ;
        RECT 25.655 143.800 25.985 144.160 ;
        RECT 26.345 144.060 26.515 146.180 ;
        RECT 26.685 145.850 27.015 146.350 ;
        RECT 27.185 145.680 27.440 146.180 ;
        RECT 26.690 145.510 27.440 145.680 ;
        RECT 26.690 144.520 26.920 145.510 ;
        RECT 27.090 144.690 27.440 145.340 ;
        RECT 28.535 145.260 32.045 146.350 ;
        RECT 28.535 144.740 30.225 145.260 ;
        RECT 32.215 145.210 32.485 146.180 ;
        RECT 32.695 145.550 32.975 146.350 ;
        RECT 33.145 145.840 34.800 146.130 ;
        RECT 33.210 145.500 34.800 145.670 ;
        RECT 33.210 145.380 33.380 145.500 ;
        RECT 32.655 145.210 33.380 145.380 ;
        RECT 30.395 144.570 32.045 145.090 ;
        RECT 26.690 144.350 27.440 144.520 ;
        RECT 26.685 143.800 27.015 144.180 ;
        RECT 27.185 144.060 27.440 144.350 ;
        RECT 28.535 143.800 32.045 144.570 ;
        RECT 32.215 144.475 32.385 145.210 ;
        RECT 32.655 145.040 32.825 145.210 ;
        RECT 32.555 144.710 32.825 145.040 ;
        RECT 32.995 144.710 33.400 145.040 ;
        RECT 33.570 144.710 34.280 145.330 ;
        RECT 34.480 145.210 34.800 145.500 ;
        RECT 34.975 145.210 35.315 146.180 ;
        RECT 35.485 145.210 35.655 146.350 ;
        RECT 35.925 145.550 36.175 146.350 ;
        RECT 36.820 145.380 37.150 146.180 ;
        RECT 37.450 145.550 37.780 146.350 ;
        RECT 37.950 145.380 38.280 146.180 ;
        RECT 35.845 145.210 38.280 145.380 ;
        RECT 39.115 145.260 40.785 146.350 ;
        RECT 32.655 144.540 32.825 144.710 ;
        RECT 32.215 144.130 32.485 144.475 ;
        RECT 32.655 144.370 34.265 144.540 ;
        RECT 34.450 144.470 34.800 145.040 ;
        RECT 34.975 144.600 35.150 145.210 ;
        RECT 35.845 144.960 36.015 145.210 ;
        RECT 35.320 144.790 36.015 144.960 ;
        RECT 36.190 144.790 36.610 144.990 ;
        RECT 36.780 144.790 37.110 144.990 ;
        RECT 37.280 144.790 37.610 144.990 ;
        RECT 32.675 143.800 33.055 144.200 ;
        RECT 33.225 144.020 33.395 144.370 ;
        RECT 33.565 143.800 33.895 144.200 ;
        RECT 34.095 144.020 34.265 144.370 ;
        RECT 34.465 143.800 34.795 144.300 ;
        RECT 34.975 143.970 35.315 144.600 ;
        RECT 35.485 143.800 35.735 144.600 ;
        RECT 35.925 144.450 37.150 144.620 ;
        RECT 35.925 143.970 36.255 144.450 ;
        RECT 36.425 143.800 36.650 144.260 ;
        RECT 36.820 143.970 37.150 144.450 ;
        RECT 37.780 144.580 37.950 145.210 ;
        RECT 38.135 144.790 38.485 145.040 ;
        RECT 39.115 144.740 39.865 145.260 ;
        RECT 40.955 145.185 41.245 146.350 ;
        RECT 41.875 145.260 44.465 146.350 ;
        RECT 37.780 143.970 38.280 144.580 ;
        RECT 40.035 144.570 40.785 145.090 ;
        RECT 41.875 144.740 43.085 145.260 ;
        RECT 44.635 145.210 44.975 146.180 ;
        RECT 45.145 145.210 45.315 146.350 ;
        RECT 45.585 145.550 45.835 146.350 ;
        RECT 46.480 145.380 46.810 146.180 ;
        RECT 47.110 145.550 47.440 146.350 ;
        RECT 47.610 145.380 47.940 146.180 ;
        RECT 45.505 145.210 47.940 145.380 ;
        RECT 48.775 145.260 50.445 146.350 ;
        RECT 43.255 144.570 44.465 145.090 ;
        RECT 39.115 143.800 40.785 144.570 ;
        RECT 40.955 143.800 41.245 144.525 ;
        RECT 41.875 143.800 44.465 144.570 ;
        RECT 44.635 144.600 44.810 145.210 ;
        RECT 45.505 144.960 45.675 145.210 ;
        RECT 44.980 144.790 45.675 144.960 ;
        RECT 45.850 144.790 46.270 144.990 ;
        RECT 46.440 144.790 46.770 144.990 ;
        RECT 46.940 144.790 47.270 144.990 ;
        RECT 44.635 143.970 44.975 144.600 ;
        RECT 45.145 143.800 45.395 144.600 ;
        RECT 45.585 144.450 46.810 144.620 ;
        RECT 45.585 143.970 45.915 144.450 ;
        RECT 46.085 143.800 46.310 144.260 ;
        RECT 46.480 143.970 46.810 144.450 ;
        RECT 47.440 144.580 47.610 145.210 ;
        RECT 47.795 144.790 48.145 145.040 ;
        RECT 48.775 144.740 49.525 145.260 ;
        RECT 50.675 145.210 50.885 146.350 ;
        RECT 51.055 145.200 51.385 146.180 ;
        RECT 51.555 145.210 51.785 146.350 ;
        RECT 52.455 145.260 54.125 146.350 ;
        RECT 47.440 143.970 47.940 144.580 ;
        RECT 49.695 144.570 50.445 145.090 ;
        RECT 48.775 143.800 50.445 144.570 ;
        RECT 50.675 143.800 50.885 144.620 ;
        RECT 51.055 144.600 51.305 145.200 ;
        RECT 51.475 144.790 51.805 145.040 ;
        RECT 52.455 144.740 53.205 145.260 ;
        RECT 54.335 145.210 54.565 146.350 ;
        RECT 54.735 145.200 55.065 146.180 ;
        RECT 55.235 145.210 55.445 146.350 ;
        RECT 56.050 146.010 56.305 146.040 ;
        RECT 55.965 145.840 56.305 146.010 ;
        RECT 56.050 145.370 56.305 145.840 ;
        RECT 56.485 145.550 56.770 146.350 ;
        RECT 56.950 145.630 57.280 146.140 ;
        RECT 51.055 143.970 51.385 144.600 ;
        RECT 51.555 143.800 51.785 144.620 ;
        RECT 53.375 144.570 54.125 145.090 ;
        RECT 54.315 144.790 54.645 145.040 ;
        RECT 52.455 143.800 54.125 144.570 ;
        RECT 54.335 143.800 54.565 144.620 ;
        RECT 54.815 144.600 55.065 145.200 ;
        RECT 54.735 143.970 55.065 144.600 ;
        RECT 55.235 143.800 55.445 144.620 ;
        RECT 56.050 144.510 56.230 145.370 ;
        RECT 56.950 145.040 57.200 145.630 ;
        RECT 57.550 145.480 57.720 146.090 ;
        RECT 57.890 145.660 58.220 146.350 ;
        RECT 58.450 145.800 58.690 146.090 ;
        RECT 58.890 145.970 59.310 146.350 ;
        RECT 59.490 145.880 60.120 146.130 ;
        RECT 60.590 145.970 60.920 146.350 ;
        RECT 59.490 145.800 59.660 145.880 ;
        RECT 61.090 145.800 61.260 146.090 ;
        RECT 61.440 145.970 61.820 146.350 ;
        RECT 62.060 145.965 62.890 146.135 ;
        RECT 58.450 145.630 59.660 145.800 ;
        RECT 56.400 144.710 57.200 145.040 ;
        RECT 56.050 143.980 56.305 144.510 ;
        RECT 56.485 143.800 56.770 144.260 ;
        RECT 56.950 144.060 57.200 144.710 ;
        RECT 57.400 145.460 57.720 145.480 ;
        RECT 57.400 145.290 59.320 145.460 ;
        RECT 57.400 144.395 57.590 145.290 ;
        RECT 59.490 145.120 59.660 145.630 ;
        RECT 59.830 145.370 60.350 145.680 ;
        RECT 57.760 144.950 59.660 145.120 ;
        RECT 57.760 144.890 58.090 144.950 ;
        RECT 58.240 144.720 58.570 144.780 ;
        RECT 57.910 144.450 58.570 144.720 ;
        RECT 57.400 144.065 57.720 144.395 ;
        RECT 57.900 143.800 58.560 144.280 ;
        RECT 58.760 144.190 58.930 144.950 ;
        RECT 59.830 144.780 60.010 145.190 ;
        RECT 59.100 144.610 59.430 144.730 ;
        RECT 60.180 144.610 60.350 145.370 ;
        RECT 59.100 144.440 60.350 144.610 ;
        RECT 60.520 145.550 61.890 145.800 ;
        RECT 60.520 144.780 60.710 145.550 ;
        RECT 61.640 145.290 61.890 145.550 ;
        RECT 60.880 145.120 61.130 145.280 ;
        RECT 62.060 145.120 62.230 145.965 ;
        RECT 63.125 145.680 63.295 146.180 ;
        RECT 63.465 145.850 63.795 146.350 ;
        RECT 62.400 145.290 62.900 145.670 ;
        RECT 63.125 145.510 63.820 145.680 ;
        RECT 60.880 144.950 62.230 145.120 ;
        RECT 61.810 144.910 62.230 144.950 ;
        RECT 60.520 144.440 60.940 144.780 ;
        RECT 61.230 144.450 61.640 144.780 ;
        RECT 58.760 144.020 59.610 144.190 ;
        RECT 60.170 143.800 60.490 144.260 ;
        RECT 60.690 144.010 60.940 144.440 ;
        RECT 61.230 143.800 61.640 144.240 ;
        RECT 61.810 144.180 61.980 144.910 ;
        RECT 62.150 144.360 62.500 144.730 ;
        RECT 62.680 144.420 62.900 145.290 ;
        RECT 63.070 144.720 63.480 145.340 ;
        RECT 63.650 144.540 63.820 145.510 ;
        RECT 63.125 144.350 63.820 144.540 ;
        RECT 61.810 143.980 62.825 144.180 ;
        RECT 63.125 144.020 63.295 144.350 ;
        RECT 63.465 143.800 63.795 144.180 ;
        RECT 64.010 144.060 64.235 146.180 ;
        RECT 64.405 145.850 64.735 146.350 ;
        RECT 64.905 145.680 65.075 146.180 ;
        RECT 64.410 145.510 65.075 145.680 ;
        RECT 64.410 144.520 64.640 145.510 ;
        RECT 64.810 144.690 65.160 145.340 ;
        RECT 65.335 145.260 66.545 146.350 ;
        RECT 65.335 144.720 65.855 145.260 ;
        RECT 66.715 145.185 67.005 146.350 ;
        RECT 67.635 145.260 71.145 146.350 ;
        RECT 66.025 144.550 66.545 145.090 ;
        RECT 67.635 144.740 69.325 145.260 ;
        RECT 71.315 145.210 71.585 146.180 ;
        RECT 71.795 145.550 72.075 146.350 ;
        RECT 72.245 145.840 73.900 146.130 ;
        RECT 72.310 145.500 73.900 145.670 ;
        RECT 72.310 145.380 72.480 145.500 ;
        RECT 71.755 145.210 72.480 145.380 ;
        RECT 69.495 144.570 71.145 145.090 ;
        RECT 64.410 144.350 65.075 144.520 ;
        RECT 64.405 143.800 64.735 144.180 ;
        RECT 64.905 144.060 65.075 144.350 ;
        RECT 65.335 143.800 66.545 144.550 ;
        RECT 66.715 143.800 67.005 144.525 ;
        RECT 67.635 143.800 71.145 144.570 ;
        RECT 71.315 144.475 71.485 145.210 ;
        RECT 71.755 145.040 71.925 145.210 ;
        RECT 71.655 144.710 71.925 145.040 ;
        RECT 72.095 144.710 72.500 145.040 ;
        RECT 72.670 144.710 73.380 145.330 ;
        RECT 73.580 145.210 73.900 145.500 ;
        RECT 74.075 145.210 74.415 146.180 ;
        RECT 74.585 145.210 74.755 146.350 ;
        RECT 75.025 145.550 75.275 146.350 ;
        RECT 75.920 145.380 76.250 146.180 ;
        RECT 76.550 145.550 76.880 146.350 ;
        RECT 77.050 145.380 77.380 146.180 ;
        RECT 74.945 145.210 77.380 145.380 ;
        RECT 77.755 145.260 81.265 146.350 ;
        RECT 81.435 145.590 81.950 146.000 ;
        RECT 82.185 145.590 82.355 146.350 ;
        RECT 82.525 146.010 84.555 146.180 ;
        RECT 71.755 144.540 71.925 144.710 ;
        RECT 71.315 144.130 71.585 144.475 ;
        RECT 71.755 144.370 73.365 144.540 ;
        RECT 73.550 144.470 73.900 145.040 ;
        RECT 74.075 144.650 74.250 145.210 ;
        RECT 74.945 144.960 75.115 145.210 ;
        RECT 74.420 144.790 75.115 144.960 ;
        RECT 75.290 144.790 75.710 144.990 ;
        RECT 75.880 144.790 76.210 144.990 ;
        RECT 76.380 144.790 76.710 144.990 ;
        RECT 74.075 144.600 74.305 144.650 ;
        RECT 71.775 143.800 72.155 144.200 ;
        RECT 72.325 144.020 72.495 144.370 ;
        RECT 72.665 143.800 72.995 144.200 ;
        RECT 73.195 144.020 73.365 144.370 ;
        RECT 73.565 143.800 73.895 144.300 ;
        RECT 74.075 143.970 74.415 144.600 ;
        RECT 74.585 143.800 74.835 144.600 ;
        RECT 75.025 144.450 76.250 144.620 ;
        RECT 75.025 143.970 75.355 144.450 ;
        RECT 75.525 143.800 75.750 144.260 ;
        RECT 75.920 143.970 76.250 144.450 ;
        RECT 76.880 144.580 77.050 145.210 ;
        RECT 77.235 144.790 77.585 145.040 ;
        RECT 77.755 144.740 79.445 145.260 ;
        RECT 76.880 143.970 77.380 144.580 ;
        RECT 79.615 144.570 81.265 145.090 ;
        RECT 81.435 144.780 81.775 145.590 ;
        RECT 82.525 145.345 82.695 146.010 ;
        RECT 83.090 145.670 84.215 145.840 ;
        RECT 81.945 145.155 82.695 145.345 ;
        RECT 82.865 145.330 83.875 145.500 ;
        RECT 81.435 144.610 82.665 144.780 ;
        RECT 77.755 143.800 81.265 144.570 ;
        RECT 81.710 144.005 81.955 144.610 ;
        RECT 82.175 143.800 82.685 144.335 ;
        RECT 82.865 143.970 83.055 145.330 ;
        RECT 83.225 144.310 83.500 145.130 ;
        RECT 83.705 144.530 83.875 145.330 ;
        RECT 84.045 144.540 84.215 145.670 ;
        RECT 84.385 145.040 84.555 146.010 ;
        RECT 84.725 145.210 84.895 146.350 ;
        RECT 85.065 145.210 85.400 146.180 ;
        RECT 85.635 145.210 85.845 146.350 ;
        RECT 84.385 144.710 84.580 145.040 ;
        RECT 84.805 144.710 85.060 145.040 ;
        RECT 84.805 144.540 84.975 144.710 ;
        RECT 85.230 144.540 85.400 145.210 ;
        RECT 86.015 145.200 86.345 146.180 ;
        RECT 86.515 145.210 86.745 146.350 ;
        RECT 87.045 145.420 87.215 146.180 ;
        RECT 87.395 145.590 87.725 146.350 ;
        RECT 87.045 145.250 87.710 145.420 ;
        RECT 87.895 145.275 88.165 146.180 ;
        RECT 84.045 144.370 84.975 144.540 ;
        RECT 84.045 144.335 84.220 144.370 ;
        RECT 83.225 144.140 83.505 144.310 ;
        RECT 83.225 143.970 83.500 144.140 ;
        RECT 83.690 143.970 84.220 144.335 ;
        RECT 84.645 143.800 84.975 144.200 ;
        RECT 85.145 143.970 85.400 144.540 ;
        RECT 85.635 143.800 85.845 144.620 ;
        RECT 86.015 144.600 86.265 145.200 ;
        RECT 87.540 145.105 87.710 145.250 ;
        RECT 86.435 144.790 86.765 145.040 ;
        RECT 86.975 144.700 87.305 145.070 ;
        RECT 87.540 144.775 87.825 145.105 ;
        RECT 86.015 143.970 86.345 144.600 ;
        RECT 86.515 143.800 86.745 144.620 ;
        RECT 87.540 144.520 87.710 144.775 ;
        RECT 87.045 144.350 87.710 144.520 ;
        RECT 87.995 144.475 88.165 145.275 ;
        RECT 88.795 145.260 92.305 146.350 ;
        RECT 88.795 144.740 90.485 145.260 ;
        RECT 92.475 145.185 92.765 146.350 ;
        RECT 93.895 145.210 94.125 146.350 ;
        RECT 94.295 145.200 94.625 146.180 ;
        RECT 94.795 145.210 95.005 146.350 ;
        RECT 95.610 146.010 95.865 146.040 ;
        RECT 95.525 145.840 95.865 146.010 ;
        RECT 95.610 145.370 95.865 145.840 ;
        RECT 96.045 145.550 96.330 146.350 ;
        RECT 96.510 145.630 96.840 146.140 ;
        RECT 90.655 144.570 92.305 145.090 ;
        RECT 93.875 144.790 94.205 145.040 ;
        RECT 87.045 143.970 87.215 144.350 ;
        RECT 87.395 143.800 87.725 144.180 ;
        RECT 87.905 143.970 88.165 144.475 ;
        RECT 88.795 143.800 92.305 144.570 ;
        RECT 92.475 143.800 92.765 144.525 ;
        RECT 93.895 143.800 94.125 144.620 ;
        RECT 94.375 144.600 94.625 145.200 ;
        RECT 94.295 143.970 94.625 144.600 ;
        RECT 94.795 143.800 95.005 144.620 ;
        RECT 95.610 144.510 95.790 145.370 ;
        RECT 96.510 145.040 96.760 145.630 ;
        RECT 97.110 145.480 97.280 146.090 ;
        RECT 97.450 145.660 97.780 146.350 ;
        RECT 98.010 145.800 98.250 146.090 ;
        RECT 98.450 145.970 98.870 146.350 ;
        RECT 99.050 145.880 99.680 146.130 ;
        RECT 100.150 145.970 100.480 146.350 ;
        RECT 99.050 145.800 99.220 145.880 ;
        RECT 100.650 145.800 100.820 146.090 ;
        RECT 101.000 145.970 101.380 146.350 ;
        RECT 101.620 145.965 102.450 146.135 ;
        RECT 98.010 145.630 99.220 145.800 ;
        RECT 95.960 144.710 96.760 145.040 ;
        RECT 95.610 143.980 95.865 144.510 ;
        RECT 96.045 143.800 96.330 144.260 ;
        RECT 96.510 144.060 96.760 144.710 ;
        RECT 96.960 145.460 97.280 145.480 ;
        RECT 96.960 145.290 98.880 145.460 ;
        RECT 96.960 144.395 97.150 145.290 ;
        RECT 99.050 145.120 99.220 145.630 ;
        RECT 99.390 145.370 99.910 145.680 ;
        RECT 97.320 144.950 99.220 145.120 ;
        RECT 97.320 144.890 97.650 144.950 ;
        RECT 97.800 144.720 98.130 144.780 ;
        RECT 97.470 144.450 98.130 144.720 ;
        RECT 96.960 144.065 97.280 144.395 ;
        RECT 97.460 143.800 98.120 144.280 ;
        RECT 98.320 144.190 98.490 144.950 ;
        RECT 99.390 144.780 99.570 145.190 ;
        RECT 98.660 144.610 98.990 144.730 ;
        RECT 99.740 144.610 99.910 145.370 ;
        RECT 98.660 144.440 99.910 144.610 ;
        RECT 100.080 145.550 101.450 145.800 ;
        RECT 100.080 144.780 100.270 145.550 ;
        RECT 101.200 145.290 101.450 145.550 ;
        RECT 100.440 145.120 100.690 145.280 ;
        RECT 101.620 145.120 101.790 145.965 ;
        RECT 102.685 145.680 102.855 146.180 ;
        RECT 103.025 145.850 103.355 146.350 ;
        RECT 101.960 145.290 102.460 145.670 ;
        RECT 102.685 145.510 103.380 145.680 ;
        RECT 100.440 144.950 101.790 145.120 ;
        RECT 101.370 144.910 101.790 144.950 ;
        RECT 100.080 144.440 100.500 144.780 ;
        RECT 100.790 144.450 101.200 144.780 ;
        RECT 98.320 144.020 99.170 144.190 ;
        RECT 99.730 143.800 100.050 144.260 ;
        RECT 100.250 144.010 100.500 144.440 ;
        RECT 100.790 143.800 101.200 144.240 ;
        RECT 101.370 144.180 101.540 144.910 ;
        RECT 101.710 144.360 102.060 144.730 ;
        RECT 102.240 144.420 102.460 145.290 ;
        RECT 102.630 144.720 103.040 145.340 ;
        RECT 103.210 144.540 103.380 145.510 ;
        RECT 102.685 144.350 103.380 144.540 ;
        RECT 101.370 143.980 102.385 144.180 ;
        RECT 102.685 144.020 102.855 144.350 ;
        RECT 103.025 143.800 103.355 144.180 ;
        RECT 103.570 144.060 103.795 146.180 ;
        RECT 103.965 145.850 104.295 146.350 ;
        RECT 104.465 145.680 104.635 146.180 ;
        RECT 103.970 145.510 104.635 145.680 ;
        RECT 103.970 144.520 104.200 145.510 ;
        RECT 104.370 144.690 104.720 145.340 ;
        RECT 104.895 145.260 106.105 146.350 ;
        RECT 106.275 145.590 106.790 146.000 ;
        RECT 107.025 145.590 107.195 146.350 ;
        RECT 107.365 146.010 109.395 146.180 ;
        RECT 104.895 144.720 105.415 145.260 ;
        RECT 105.585 144.550 106.105 145.090 ;
        RECT 106.275 144.780 106.615 145.590 ;
        RECT 107.365 145.345 107.535 146.010 ;
        RECT 107.930 145.670 109.055 145.840 ;
        RECT 106.785 145.155 107.535 145.345 ;
        RECT 107.705 145.330 108.715 145.500 ;
        RECT 106.275 144.610 107.505 144.780 ;
        RECT 103.970 144.350 104.635 144.520 ;
        RECT 103.965 143.800 104.295 144.180 ;
        RECT 104.465 144.060 104.635 144.350 ;
        RECT 104.895 143.800 106.105 144.550 ;
        RECT 106.550 144.005 106.795 144.610 ;
        RECT 107.015 143.800 107.525 144.335 ;
        RECT 107.705 143.970 107.895 145.330 ;
        RECT 108.065 144.990 108.340 145.130 ;
        RECT 108.065 144.820 108.345 144.990 ;
        RECT 108.065 143.970 108.340 144.820 ;
        RECT 108.545 144.530 108.715 145.330 ;
        RECT 108.885 144.540 109.055 145.670 ;
        RECT 109.225 145.040 109.395 146.010 ;
        RECT 109.565 145.210 109.735 146.350 ;
        RECT 109.905 145.210 110.240 146.180 ;
        RECT 111.425 145.420 111.595 146.180 ;
        RECT 111.775 145.590 112.105 146.350 ;
        RECT 111.425 145.250 112.090 145.420 ;
        RECT 112.275 145.275 112.545 146.180 ;
        RECT 109.225 144.710 109.420 145.040 ;
        RECT 109.645 144.710 109.900 145.040 ;
        RECT 109.645 144.540 109.815 144.710 ;
        RECT 110.070 144.540 110.240 145.210 ;
        RECT 111.920 145.105 112.090 145.250 ;
        RECT 111.355 144.700 111.685 145.070 ;
        RECT 111.920 144.775 112.205 145.105 ;
        RECT 108.885 144.370 109.815 144.540 ;
        RECT 108.885 144.335 109.060 144.370 ;
        RECT 108.530 143.970 109.060 144.335 ;
        RECT 109.485 143.800 109.815 144.200 ;
        RECT 109.985 143.970 110.240 144.540 ;
        RECT 111.920 144.520 112.090 144.775 ;
        RECT 111.425 144.350 112.090 144.520 ;
        RECT 112.375 144.475 112.545 145.275 ;
        RECT 113.635 145.260 117.145 146.350 ;
        RECT 117.315 145.260 118.525 146.350 ;
        RECT 113.635 144.740 115.325 145.260 ;
        RECT 115.495 144.570 117.145 145.090 ;
        RECT 117.315 144.720 117.835 145.260 ;
        RECT 111.425 143.970 111.595 144.350 ;
        RECT 111.775 143.800 112.105 144.180 ;
        RECT 112.285 143.970 112.545 144.475 ;
        RECT 113.635 143.800 117.145 144.570 ;
        RECT 118.005 144.550 118.525 145.090 ;
        RECT 117.315 143.800 118.525 144.550 ;
        RECT 11.430 143.630 118.610 143.800 ;
        RECT 11.515 142.880 12.725 143.630 ;
        RECT 13.470 143.000 13.755 143.460 ;
        RECT 13.925 143.170 14.195 143.630 ;
        RECT 11.515 142.340 12.035 142.880 ;
        RECT 13.470 142.830 14.425 143.000 ;
        RECT 12.205 142.170 12.725 142.710 ;
        RECT 11.515 141.080 12.725 142.170 ;
        RECT 13.355 142.100 14.045 142.660 ;
        RECT 14.215 141.930 14.425 142.830 ;
        RECT 13.470 141.710 14.425 141.930 ;
        RECT 14.595 142.660 14.995 143.460 ;
        RECT 15.185 143.000 15.465 143.460 ;
        RECT 15.985 143.170 16.310 143.630 ;
        RECT 15.185 142.830 16.310 143.000 ;
        RECT 16.480 142.890 16.865 143.460 ;
        RECT 15.860 142.720 16.310 142.830 ;
        RECT 14.595 142.100 15.690 142.660 ;
        RECT 15.860 142.390 16.415 142.720 ;
        RECT 13.470 141.250 13.755 141.710 ;
        RECT 13.925 141.080 14.195 141.540 ;
        RECT 14.595 141.250 14.995 142.100 ;
        RECT 15.860 141.930 16.310 142.390 ;
        RECT 16.585 142.220 16.865 142.890 ;
        RECT 17.035 142.860 18.705 143.630 ;
        RECT 15.185 141.710 16.310 141.930 ;
        RECT 15.185 141.250 15.465 141.710 ;
        RECT 15.985 141.080 16.310 141.540 ;
        RECT 16.480 141.250 16.865 142.220 ;
        RECT 17.035 142.170 17.785 142.690 ;
        RECT 17.955 142.340 18.705 142.860 ;
        RECT 18.880 142.890 19.135 143.460 ;
        RECT 19.305 143.230 19.635 143.630 ;
        RECT 20.060 143.095 20.590 143.460 ;
        RECT 20.780 143.290 21.055 143.460 ;
        RECT 20.775 143.120 21.055 143.290 ;
        RECT 20.060 143.060 20.235 143.095 ;
        RECT 19.305 142.890 20.235 143.060 ;
        RECT 18.880 142.220 19.050 142.890 ;
        RECT 19.305 142.720 19.475 142.890 ;
        RECT 19.220 142.390 19.475 142.720 ;
        RECT 19.700 142.390 19.895 142.720 ;
        RECT 17.035 141.080 18.705 142.170 ;
        RECT 18.880 141.250 19.215 142.220 ;
        RECT 19.385 141.080 19.555 142.220 ;
        RECT 19.725 141.420 19.895 142.390 ;
        RECT 20.065 141.760 20.235 142.890 ;
        RECT 20.405 142.100 20.575 142.900 ;
        RECT 20.780 142.300 21.055 143.120 ;
        RECT 21.225 142.100 21.415 143.460 ;
        RECT 21.595 143.095 22.105 143.630 ;
        RECT 22.325 142.820 22.570 143.425 ;
        RECT 23.015 142.880 24.225 143.630 ;
        RECT 24.485 143.080 24.655 143.460 ;
        RECT 24.835 143.250 25.165 143.630 ;
        RECT 24.485 142.910 25.150 143.080 ;
        RECT 25.345 142.955 25.605 143.460 ;
        RECT 21.615 142.650 22.845 142.820 ;
        RECT 20.405 141.930 21.415 142.100 ;
        RECT 21.585 142.085 22.335 142.275 ;
        RECT 20.065 141.590 21.190 141.760 ;
        RECT 21.585 141.420 21.755 142.085 ;
        RECT 22.505 141.840 22.845 142.650 ;
        RECT 19.725 141.250 21.755 141.420 ;
        RECT 21.925 141.080 22.095 141.840 ;
        RECT 22.330 141.430 22.845 141.840 ;
        RECT 23.015 142.170 23.535 142.710 ;
        RECT 23.705 142.340 24.225 142.880 ;
        RECT 24.415 142.360 24.745 142.730 ;
        RECT 24.980 142.655 25.150 142.910 ;
        RECT 24.980 142.325 25.265 142.655 ;
        RECT 24.980 142.180 25.150 142.325 ;
        RECT 23.015 141.080 24.225 142.170 ;
        RECT 24.485 142.010 25.150 142.180 ;
        RECT 25.435 142.155 25.605 142.955 ;
        RECT 26.235 142.860 27.905 143.630 ;
        RECT 28.075 142.905 28.365 143.630 ;
        RECT 28.995 142.860 32.505 143.630 ;
        RECT 32.685 143.130 33.015 143.630 ;
        RECT 33.215 143.060 33.385 143.410 ;
        RECT 33.585 143.230 33.915 143.630 ;
        RECT 34.085 143.060 34.255 143.410 ;
        RECT 34.425 143.230 34.805 143.630 ;
        RECT 24.485 141.250 24.655 142.010 ;
        RECT 24.835 141.080 25.165 141.840 ;
        RECT 25.335 141.250 25.605 142.155 ;
        RECT 26.235 142.170 26.985 142.690 ;
        RECT 27.155 142.340 27.905 142.860 ;
        RECT 26.235 141.080 27.905 142.170 ;
        RECT 28.075 141.080 28.365 142.245 ;
        RECT 28.995 142.170 30.685 142.690 ;
        RECT 30.855 142.340 32.505 142.860 ;
        RECT 32.680 142.390 33.030 142.960 ;
        RECT 33.215 142.890 34.825 143.060 ;
        RECT 34.995 142.955 35.265 143.300 ;
        RECT 34.655 142.720 34.825 142.890 ;
        RECT 28.995 141.080 32.505 142.170 ;
        RECT 32.680 141.930 33.000 142.220 ;
        RECT 33.200 142.100 33.910 142.720 ;
        RECT 34.080 142.390 34.485 142.720 ;
        RECT 34.655 142.390 34.925 142.720 ;
        RECT 34.655 142.220 34.825 142.390 ;
        RECT 35.095 142.220 35.265 142.955 ;
        RECT 34.100 142.050 34.825 142.220 ;
        RECT 34.100 141.930 34.270 142.050 ;
        RECT 32.680 141.760 34.270 141.930 ;
        RECT 32.680 141.300 34.335 141.590 ;
        RECT 34.505 141.080 34.785 141.880 ;
        RECT 34.995 141.250 35.265 142.220 ;
        RECT 35.435 142.955 35.705 143.300 ;
        RECT 35.895 143.230 36.275 143.630 ;
        RECT 36.445 143.060 36.615 143.410 ;
        RECT 36.785 143.230 37.115 143.630 ;
        RECT 37.315 143.060 37.485 143.410 ;
        RECT 37.685 143.130 38.015 143.630 ;
        RECT 35.435 142.220 35.605 142.955 ;
        RECT 35.875 142.890 37.485 143.060 ;
        RECT 35.875 142.720 36.045 142.890 ;
        RECT 35.775 142.390 36.045 142.720 ;
        RECT 36.215 142.390 36.620 142.720 ;
        RECT 35.875 142.220 36.045 142.390 ;
        RECT 35.435 141.250 35.705 142.220 ;
        RECT 35.875 142.050 36.600 142.220 ;
        RECT 36.790 142.100 37.500 142.720 ;
        RECT 37.670 142.390 38.020 142.960 ;
        RECT 38.655 142.860 40.325 143.630 ;
        RECT 40.500 143.085 45.845 143.630 ;
        RECT 36.430 141.930 36.600 142.050 ;
        RECT 37.700 141.930 38.020 142.220 ;
        RECT 35.915 141.080 36.195 141.880 ;
        RECT 36.430 141.760 38.020 141.930 ;
        RECT 38.655 142.170 39.405 142.690 ;
        RECT 39.575 142.340 40.325 142.860 ;
        RECT 36.365 141.300 38.020 141.590 ;
        RECT 38.655 141.080 40.325 142.170 ;
        RECT 42.090 141.515 42.440 142.765 ;
        RECT 43.920 142.255 44.260 143.085 ;
        RECT 46.015 142.830 46.355 143.460 ;
        RECT 46.525 142.830 46.775 143.630 ;
        RECT 46.965 142.980 47.295 143.460 ;
        RECT 47.465 143.170 47.690 143.630 ;
        RECT 47.860 142.980 48.190 143.460 ;
        RECT 46.015 142.220 46.190 142.830 ;
        RECT 46.965 142.810 48.190 142.980 ;
        RECT 48.820 142.850 49.320 143.460 ;
        RECT 46.360 142.470 47.055 142.640 ;
        RECT 46.885 142.220 47.055 142.470 ;
        RECT 47.230 142.440 47.650 142.640 ;
        RECT 47.820 142.440 48.150 142.640 ;
        RECT 48.320 142.440 48.650 142.640 ;
        RECT 48.820 142.220 48.990 142.850 ;
        RECT 49.970 142.820 50.215 143.425 ;
        RECT 50.435 143.095 50.945 143.630 ;
        RECT 49.695 142.650 50.925 142.820 ;
        RECT 49.175 142.390 49.525 142.640 ;
        RECT 40.500 141.080 45.845 141.515 ;
        RECT 46.015 141.250 46.355 142.220 ;
        RECT 46.525 141.080 46.695 142.220 ;
        RECT 46.885 142.050 49.320 142.220 ;
        RECT 46.965 141.080 47.215 141.880 ;
        RECT 47.860 141.250 48.190 142.050 ;
        RECT 48.490 141.080 48.820 141.880 ;
        RECT 48.990 141.250 49.320 142.050 ;
        RECT 49.695 141.840 50.035 142.650 ;
        RECT 50.205 142.085 50.955 142.275 ;
        RECT 49.695 141.430 50.210 141.840 ;
        RECT 50.445 141.080 50.615 141.840 ;
        RECT 50.785 141.420 50.955 142.085 ;
        RECT 51.125 142.100 51.315 143.460 ;
        RECT 51.485 143.290 51.760 143.460 ;
        RECT 51.485 143.120 51.765 143.290 ;
        RECT 51.485 142.300 51.760 143.120 ;
        RECT 51.950 143.095 52.480 143.460 ;
        RECT 52.905 143.230 53.235 143.630 ;
        RECT 52.305 143.060 52.480 143.095 ;
        RECT 51.965 142.100 52.135 142.900 ;
        RECT 51.125 141.930 52.135 142.100 ;
        RECT 52.305 142.890 53.235 143.060 ;
        RECT 53.405 142.890 53.660 143.460 ;
        RECT 53.835 142.905 54.125 143.630 ;
        RECT 52.305 141.760 52.475 142.890 ;
        RECT 53.065 142.720 53.235 142.890 ;
        RECT 51.350 141.590 52.475 141.760 ;
        RECT 52.645 142.390 52.840 142.720 ;
        RECT 53.065 142.390 53.320 142.720 ;
        RECT 52.645 141.420 52.815 142.390 ;
        RECT 53.490 142.220 53.660 142.890 ;
        RECT 54.295 142.880 55.505 143.630 ;
        RECT 50.785 141.250 52.815 141.420 ;
        RECT 52.985 141.080 53.155 142.220 ;
        RECT 53.325 141.250 53.660 142.220 ;
        RECT 53.835 141.080 54.125 142.245 ;
        RECT 54.295 142.170 54.815 142.710 ;
        RECT 54.985 142.340 55.505 142.880 ;
        RECT 56.050 142.920 56.305 143.450 ;
        RECT 56.485 143.170 56.770 143.630 ;
        RECT 54.295 141.080 55.505 142.170 ;
        RECT 56.050 142.060 56.230 142.920 ;
        RECT 56.950 142.720 57.200 143.370 ;
        RECT 56.400 142.390 57.200 142.720 ;
        RECT 56.050 141.930 56.305 142.060 ;
        RECT 55.965 141.760 56.305 141.930 ;
        RECT 56.050 141.390 56.305 141.760 ;
        RECT 56.485 141.080 56.770 141.880 ;
        RECT 56.950 141.800 57.200 142.390 ;
        RECT 57.400 143.035 57.720 143.365 ;
        RECT 57.900 143.150 58.560 143.630 ;
        RECT 58.760 143.240 59.610 143.410 ;
        RECT 57.400 142.140 57.590 143.035 ;
        RECT 57.910 142.710 58.570 142.980 ;
        RECT 58.240 142.650 58.570 142.710 ;
        RECT 57.760 142.480 58.090 142.540 ;
        RECT 58.760 142.480 58.930 143.240 ;
        RECT 60.170 143.170 60.490 143.630 ;
        RECT 60.690 142.990 60.940 143.420 ;
        RECT 61.230 143.190 61.640 143.630 ;
        RECT 61.810 143.250 62.825 143.450 ;
        RECT 59.100 142.820 60.350 142.990 ;
        RECT 59.100 142.700 59.430 142.820 ;
        RECT 57.760 142.310 59.660 142.480 ;
        RECT 57.400 141.970 59.320 142.140 ;
        RECT 57.400 141.950 57.720 141.970 ;
        RECT 56.950 141.290 57.280 141.800 ;
        RECT 57.550 141.340 57.720 141.950 ;
        RECT 59.490 141.800 59.660 142.310 ;
        RECT 59.830 142.240 60.010 142.650 ;
        RECT 60.180 142.060 60.350 142.820 ;
        RECT 57.890 141.080 58.220 141.770 ;
        RECT 58.450 141.630 59.660 141.800 ;
        RECT 59.830 141.750 60.350 142.060 ;
        RECT 60.520 142.650 60.940 142.990 ;
        RECT 61.230 142.650 61.640 142.980 ;
        RECT 60.520 141.880 60.710 142.650 ;
        RECT 61.810 142.520 61.980 143.250 ;
        RECT 63.125 143.080 63.295 143.410 ;
        RECT 63.465 143.250 63.795 143.630 ;
        RECT 62.150 142.700 62.500 143.070 ;
        RECT 61.810 142.480 62.230 142.520 ;
        RECT 60.880 142.310 62.230 142.480 ;
        RECT 60.880 142.150 61.130 142.310 ;
        RECT 61.640 141.880 61.890 142.140 ;
        RECT 60.520 141.630 61.890 141.880 ;
        RECT 58.450 141.340 58.690 141.630 ;
        RECT 59.490 141.550 59.660 141.630 ;
        RECT 58.890 141.080 59.310 141.460 ;
        RECT 59.490 141.300 60.120 141.550 ;
        RECT 60.590 141.080 60.920 141.460 ;
        RECT 61.090 141.340 61.260 141.630 ;
        RECT 62.060 141.465 62.230 142.310 ;
        RECT 62.680 142.140 62.900 143.010 ;
        RECT 63.125 142.890 63.820 143.080 ;
        RECT 62.400 141.760 62.900 142.140 ;
        RECT 63.070 142.090 63.480 142.710 ;
        RECT 63.650 141.920 63.820 142.890 ;
        RECT 63.125 141.750 63.820 141.920 ;
        RECT 61.440 141.080 61.820 141.460 ;
        RECT 62.060 141.295 62.890 141.465 ;
        RECT 63.125 141.250 63.295 141.750 ;
        RECT 63.465 141.080 63.795 141.580 ;
        RECT 64.010 141.250 64.235 143.370 ;
        RECT 64.405 143.250 64.735 143.630 ;
        RECT 64.905 143.080 65.075 143.370 ;
        RECT 65.340 143.085 70.685 143.630 ;
        RECT 64.410 142.910 65.075 143.080 ;
        RECT 64.410 141.920 64.640 142.910 ;
        RECT 64.810 142.090 65.160 142.740 ;
        RECT 64.410 141.750 65.075 141.920 ;
        RECT 64.405 141.080 64.735 141.580 ;
        RECT 64.905 141.250 65.075 141.750 ;
        RECT 66.930 141.515 67.280 142.765 ;
        RECT 68.760 142.255 69.100 143.085 ;
        RECT 71.060 142.850 71.560 143.460 ;
        RECT 70.855 142.390 71.205 142.640 ;
        RECT 71.390 142.220 71.560 142.850 ;
        RECT 72.190 142.980 72.520 143.460 ;
        RECT 72.690 143.170 72.915 143.630 ;
        RECT 73.085 142.980 73.415 143.460 ;
        RECT 72.190 142.810 73.415 142.980 ;
        RECT 73.605 142.830 73.855 143.630 ;
        RECT 74.025 142.830 74.365 143.460 ;
        RECT 71.730 142.440 72.060 142.640 ;
        RECT 72.230 142.440 72.560 142.640 ;
        RECT 72.730 142.440 73.150 142.640 ;
        RECT 73.325 142.470 74.020 142.640 ;
        RECT 73.325 142.220 73.495 142.470 ;
        RECT 74.190 142.220 74.365 142.830 ;
        RECT 71.060 142.050 73.495 142.220 ;
        RECT 65.340 141.080 70.685 141.515 ;
        RECT 71.060 141.250 71.390 142.050 ;
        RECT 71.560 141.080 71.890 141.880 ;
        RECT 72.190 141.250 72.520 142.050 ;
        RECT 73.165 141.080 73.415 141.880 ;
        RECT 73.685 141.080 73.855 142.220 ;
        RECT 74.025 141.250 74.365 142.220 ;
        RECT 74.535 142.830 74.875 143.460 ;
        RECT 75.045 142.830 75.295 143.630 ;
        RECT 75.485 142.980 75.815 143.460 ;
        RECT 75.985 143.170 76.210 143.630 ;
        RECT 76.380 142.980 76.710 143.460 ;
        RECT 74.535 142.270 74.710 142.830 ;
        RECT 75.485 142.810 76.710 142.980 ;
        RECT 77.340 142.850 77.840 143.460 ;
        RECT 78.215 142.880 79.425 143.630 ;
        RECT 79.595 142.905 79.885 143.630 ;
        RECT 74.880 142.470 75.575 142.640 ;
        RECT 74.535 142.220 74.765 142.270 ;
        RECT 75.405 142.220 75.575 142.470 ;
        RECT 75.750 142.440 76.170 142.640 ;
        RECT 76.340 142.440 76.670 142.640 ;
        RECT 76.840 142.440 77.170 142.640 ;
        RECT 77.340 142.220 77.510 142.850 ;
        RECT 77.695 142.390 78.045 142.640 ;
        RECT 74.535 141.250 74.875 142.220 ;
        RECT 75.045 141.080 75.215 142.220 ;
        RECT 75.405 142.050 77.840 142.220 ;
        RECT 75.485 141.080 75.735 141.880 ;
        RECT 76.380 141.250 76.710 142.050 ;
        RECT 77.010 141.080 77.340 141.880 ;
        RECT 77.510 141.250 77.840 142.050 ;
        RECT 78.215 142.170 78.735 142.710 ;
        RECT 78.905 142.340 79.425 142.880 ;
        RECT 80.055 142.860 82.645 143.630 ;
        RECT 78.215 141.080 79.425 142.170 ;
        RECT 79.595 141.080 79.885 142.245 ;
        RECT 80.055 142.170 81.265 142.690 ;
        RECT 81.435 142.340 82.645 142.860 ;
        RECT 83.090 142.820 83.335 143.425 ;
        RECT 83.555 143.095 84.065 143.630 ;
        RECT 82.815 142.650 84.045 142.820 ;
        RECT 80.055 141.080 82.645 142.170 ;
        RECT 82.815 141.840 83.155 142.650 ;
        RECT 83.325 142.085 84.075 142.275 ;
        RECT 82.815 141.430 83.330 141.840 ;
        RECT 83.565 141.080 83.735 141.840 ;
        RECT 83.905 141.420 84.075 142.085 ;
        RECT 84.245 142.100 84.435 143.460 ;
        RECT 84.605 142.610 84.880 143.460 ;
        RECT 85.070 143.095 85.600 143.460 ;
        RECT 86.025 143.230 86.355 143.630 ;
        RECT 85.425 143.060 85.600 143.095 ;
        RECT 84.605 142.440 84.885 142.610 ;
        RECT 84.605 142.300 84.880 142.440 ;
        RECT 85.085 142.100 85.255 142.900 ;
        RECT 84.245 141.930 85.255 142.100 ;
        RECT 85.425 142.890 86.355 143.060 ;
        RECT 86.525 142.890 86.780 143.460 ;
        RECT 87.045 143.080 87.215 143.460 ;
        RECT 87.395 143.250 87.725 143.630 ;
        RECT 87.045 142.910 87.710 143.080 ;
        RECT 87.905 142.955 88.165 143.460 ;
        RECT 85.425 141.760 85.595 142.890 ;
        RECT 86.185 142.720 86.355 142.890 ;
        RECT 84.470 141.590 85.595 141.760 ;
        RECT 85.765 142.390 85.960 142.720 ;
        RECT 86.185 142.390 86.440 142.720 ;
        RECT 85.765 141.420 85.935 142.390 ;
        RECT 86.610 142.220 86.780 142.890 ;
        RECT 86.975 142.360 87.305 142.730 ;
        RECT 87.540 142.655 87.710 142.910 ;
        RECT 83.905 141.250 85.935 141.420 ;
        RECT 86.105 141.080 86.275 142.220 ;
        RECT 86.445 141.250 86.780 142.220 ;
        RECT 87.540 142.325 87.825 142.655 ;
        RECT 87.540 142.180 87.710 142.325 ;
        RECT 87.045 142.010 87.710 142.180 ;
        RECT 87.995 142.155 88.165 142.955 ;
        RECT 88.335 142.860 91.845 143.630 ;
        RECT 92.390 143.290 92.645 143.450 ;
        RECT 92.305 143.120 92.645 143.290 ;
        RECT 92.825 143.170 93.110 143.630 ;
        RECT 87.045 141.250 87.215 142.010 ;
        RECT 87.395 141.080 87.725 141.840 ;
        RECT 87.895 141.250 88.165 142.155 ;
        RECT 88.335 142.170 90.025 142.690 ;
        RECT 90.195 142.340 91.845 142.860 ;
        RECT 92.390 142.920 92.645 143.120 ;
        RECT 88.335 141.080 91.845 142.170 ;
        RECT 92.390 142.060 92.570 142.920 ;
        RECT 93.290 142.720 93.540 143.370 ;
        RECT 92.740 142.390 93.540 142.720 ;
        RECT 92.390 141.390 92.645 142.060 ;
        RECT 92.825 141.080 93.110 141.880 ;
        RECT 93.290 141.800 93.540 142.390 ;
        RECT 93.740 143.035 94.060 143.365 ;
        RECT 94.240 143.150 94.900 143.630 ;
        RECT 95.100 143.240 95.950 143.410 ;
        RECT 93.740 142.140 93.930 143.035 ;
        RECT 94.250 142.710 94.910 142.980 ;
        RECT 94.580 142.650 94.910 142.710 ;
        RECT 94.100 142.480 94.430 142.540 ;
        RECT 95.100 142.480 95.270 143.240 ;
        RECT 96.510 143.170 96.830 143.630 ;
        RECT 97.030 142.990 97.280 143.420 ;
        RECT 97.570 143.190 97.980 143.630 ;
        RECT 98.150 143.250 99.165 143.450 ;
        RECT 95.440 142.820 96.690 142.990 ;
        RECT 95.440 142.700 95.770 142.820 ;
        RECT 94.100 142.310 96.000 142.480 ;
        RECT 93.740 141.970 95.660 142.140 ;
        RECT 93.740 141.950 94.060 141.970 ;
        RECT 93.290 141.290 93.620 141.800 ;
        RECT 93.890 141.340 94.060 141.950 ;
        RECT 95.830 141.800 96.000 142.310 ;
        RECT 96.170 142.240 96.350 142.650 ;
        RECT 96.520 142.060 96.690 142.820 ;
        RECT 94.230 141.080 94.560 141.770 ;
        RECT 94.790 141.630 96.000 141.800 ;
        RECT 96.170 141.750 96.690 142.060 ;
        RECT 96.860 142.650 97.280 142.990 ;
        RECT 97.570 142.650 97.980 142.980 ;
        RECT 96.860 141.880 97.050 142.650 ;
        RECT 98.150 142.520 98.320 143.250 ;
        RECT 99.465 143.080 99.635 143.410 ;
        RECT 99.805 143.250 100.135 143.630 ;
        RECT 98.490 142.700 98.840 143.070 ;
        RECT 98.150 142.480 98.570 142.520 ;
        RECT 97.220 142.310 98.570 142.480 ;
        RECT 97.220 142.150 97.470 142.310 ;
        RECT 97.980 141.880 98.230 142.140 ;
        RECT 96.860 141.630 98.230 141.880 ;
        RECT 94.790 141.340 95.030 141.630 ;
        RECT 95.830 141.550 96.000 141.630 ;
        RECT 95.230 141.080 95.650 141.460 ;
        RECT 95.830 141.300 96.460 141.550 ;
        RECT 96.930 141.080 97.260 141.460 ;
        RECT 97.430 141.340 97.600 141.630 ;
        RECT 98.400 141.465 98.570 142.310 ;
        RECT 99.020 142.140 99.240 143.010 ;
        RECT 99.465 142.890 100.160 143.080 ;
        RECT 98.740 141.760 99.240 142.140 ;
        RECT 99.410 142.090 99.820 142.710 ;
        RECT 99.990 141.920 100.160 142.890 ;
        RECT 99.465 141.750 100.160 141.920 ;
        RECT 97.780 141.080 98.160 141.460 ;
        RECT 98.400 141.295 99.230 141.465 ;
        RECT 99.465 141.250 99.635 141.750 ;
        RECT 99.805 141.080 100.135 141.580 ;
        RECT 100.350 141.250 100.575 143.370 ;
        RECT 100.745 143.250 101.075 143.630 ;
        RECT 101.245 143.080 101.415 143.370 ;
        RECT 100.750 142.910 101.415 143.080 ;
        RECT 101.765 143.080 101.935 143.460 ;
        RECT 102.115 143.250 102.445 143.630 ;
        RECT 101.765 142.910 102.430 143.080 ;
        RECT 102.625 142.955 102.885 143.460 ;
        RECT 100.750 141.920 100.980 142.910 ;
        RECT 101.150 142.090 101.500 142.740 ;
        RECT 101.695 142.360 102.025 142.730 ;
        RECT 102.260 142.655 102.430 142.910 ;
        RECT 102.260 142.325 102.545 142.655 ;
        RECT 102.260 142.180 102.430 142.325 ;
        RECT 101.765 142.010 102.430 142.180 ;
        RECT 102.715 142.155 102.885 142.955 ;
        RECT 103.515 142.860 105.185 143.630 ;
        RECT 105.355 142.905 105.645 143.630 ;
        RECT 106.280 143.085 111.625 143.630 ;
        RECT 111.800 143.085 117.145 143.630 ;
        RECT 100.750 141.750 101.415 141.920 ;
        RECT 100.745 141.080 101.075 141.580 ;
        RECT 101.245 141.250 101.415 141.750 ;
        RECT 101.765 141.250 101.935 142.010 ;
        RECT 102.115 141.080 102.445 141.840 ;
        RECT 102.615 141.250 102.885 142.155 ;
        RECT 103.515 142.170 104.265 142.690 ;
        RECT 104.435 142.340 105.185 142.860 ;
        RECT 103.515 141.080 105.185 142.170 ;
        RECT 105.355 141.080 105.645 142.245 ;
        RECT 107.870 141.515 108.220 142.765 ;
        RECT 109.700 142.255 110.040 143.085 ;
        RECT 113.390 141.515 113.740 142.765 ;
        RECT 115.220 142.255 115.560 143.085 ;
        RECT 117.315 142.880 118.525 143.630 ;
        RECT 117.315 142.170 117.835 142.710 ;
        RECT 118.005 142.340 118.525 142.880 ;
        RECT 106.280 141.080 111.625 141.515 ;
        RECT 111.800 141.080 117.145 141.515 ;
        RECT 117.315 141.080 118.525 142.170 ;
        RECT 11.430 140.910 118.610 141.080 ;
        RECT 11.515 139.820 12.725 140.910 ;
        RECT 11.515 139.110 12.035 139.650 ;
        RECT 12.205 139.280 12.725 139.820 ;
        RECT 13.355 139.820 15.025 140.910 ;
        RECT 13.355 139.300 14.105 139.820 ;
        RECT 15.195 139.745 15.485 140.910 ;
        RECT 16.120 140.475 21.465 140.910 ;
        RECT 21.640 140.475 26.985 140.910 ;
        RECT 27.160 140.475 32.505 140.910 ;
        RECT 14.275 139.130 15.025 139.650 ;
        RECT 17.710 139.225 18.060 140.475 ;
        RECT 11.515 138.360 12.725 139.110 ;
        RECT 13.355 138.360 15.025 139.130 ;
        RECT 15.195 138.360 15.485 139.085 ;
        RECT 19.540 138.905 19.880 139.735 ;
        RECT 23.230 139.225 23.580 140.475 ;
        RECT 25.060 138.905 25.400 139.735 ;
        RECT 28.750 139.225 29.100 140.475 ;
        RECT 32.675 139.770 32.945 140.740 ;
        RECT 33.155 140.110 33.435 140.910 ;
        RECT 33.605 140.400 35.260 140.690 ;
        RECT 33.670 140.060 35.260 140.230 ;
        RECT 33.670 139.940 33.840 140.060 ;
        RECT 33.115 139.770 33.840 139.940 ;
        RECT 30.580 138.905 30.920 139.735 ;
        RECT 32.675 139.035 32.845 139.770 ;
        RECT 33.115 139.600 33.285 139.770 ;
        RECT 34.030 139.720 34.745 139.890 ;
        RECT 34.940 139.770 35.260 140.060 ;
        RECT 35.435 139.770 35.705 140.740 ;
        RECT 35.915 140.110 36.195 140.910 ;
        RECT 36.365 140.400 38.020 140.690 ;
        RECT 36.430 140.060 38.020 140.230 ;
        RECT 36.430 139.940 36.600 140.060 ;
        RECT 35.875 139.770 36.600 139.940 ;
        RECT 33.015 139.270 33.285 139.600 ;
        RECT 33.455 139.270 33.860 139.600 ;
        RECT 34.030 139.270 34.740 139.720 ;
        RECT 33.115 139.100 33.285 139.270 ;
        RECT 16.120 138.360 21.465 138.905 ;
        RECT 21.640 138.360 26.985 138.905 ;
        RECT 27.160 138.360 32.505 138.905 ;
        RECT 32.675 138.690 32.945 139.035 ;
        RECT 33.115 138.930 34.725 139.100 ;
        RECT 34.910 139.030 35.260 139.600 ;
        RECT 35.435 139.035 35.605 139.770 ;
        RECT 35.875 139.600 36.045 139.770 ;
        RECT 35.775 139.270 36.045 139.600 ;
        RECT 36.215 139.270 36.620 139.600 ;
        RECT 36.790 139.270 37.500 139.890 ;
        RECT 37.700 139.770 38.020 140.060 ;
        RECT 38.195 139.820 40.785 140.910 ;
        RECT 35.875 139.100 36.045 139.270 ;
        RECT 33.135 138.360 33.515 138.760 ;
        RECT 33.685 138.580 33.855 138.930 ;
        RECT 34.025 138.360 34.355 138.760 ;
        RECT 34.555 138.580 34.725 138.930 ;
        RECT 34.925 138.360 35.255 138.860 ;
        RECT 35.435 138.690 35.705 139.035 ;
        RECT 35.875 138.930 37.485 139.100 ;
        RECT 37.670 139.030 38.020 139.600 ;
        RECT 38.195 139.300 39.405 139.820 ;
        RECT 40.955 139.745 41.245 140.910 ;
        RECT 41.415 139.820 43.085 140.910 ;
        RECT 39.575 139.130 40.785 139.650 ;
        RECT 41.415 139.300 42.165 139.820 ;
        RECT 43.255 139.770 43.525 140.740 ;
        RECT 43.735 140.110 44.015 140.910 ;
        RECT 44.185 140.400 45.840 140.690 ;
        RECT 44.250 140.060 45.840 140.230 ;
        RECT 44.250 139.940 44.420 140.060 ;
        RECT 43.695 139.770 44.420 139.940 ;
        RECT 42.335 139.130 43.085 139.650 ;
        RECT 35.895 138.360 36.275 138.760 ;
        RECT 36.445 138.580 36.615 138.930 ;
        RECT 36.785 138.360 37.115 138.760 ;
        RECT 37.315 138.580 37.485 138.930 ;
        RECT 37.685 138.360 38.015 138.860 ;
        RECT 38.195 138.360 40.785 139.130 ;
        RECT 40.955 138.360 41.245 139.085 ;
        RECT 41.415 138.360 43.085 139.130 ;
        RECT 43.255 139.035 43.425 139.770 ;
        RECT 43.695 139.600 43.865 139.770 ;
        RECT 44.610 139.720 45.325 139.890 ;
        RECT 45.520 139.770 45.840 140.060 ;
        RECT 46.015 139.770 46.355 140.740 ;
        RECT 46.525 139.770 46.695 140.910 ;
        RECT 46.965 140.110 47.215 140.910 ;
        RECT 47.860 139.940 48.190 140.740 ;
        RECT 48.490 140.110 48.820 140.910 ;
        RECT 48.990 139.940 49.320 140.740 ;
        RECT 46.885 139.770 49.320 139.940 ;
        RECT 49.695 139.770 50.035 140.740 ;
        RECT 50.205 139.770 50.375 140.910 ;
        RECT 50.645 140.110 50.895 140.910 ;
        RECT 51.540 139.940 51.870 140.740 ;
        RECT 52.170 140.110 52.500 140.910 ;
        RECT 52.670 139.940 53.000 140.740 ;
        RECT 50.565 139.770 53.000 139.940 ;
        RECT 53.375 139.820 55.965 140.910 ;
        RECT 56.135 140.150 56.650 140.560 ;
        RECT 56.885 140.150 57.055 140.910 ;
        RECT 57.225 140.570 59.255 140.740 ;
        RECT 43.595 139.270 43.865 139.600 ;
        RECT 44.035 139.270 44.440 139.600 ;
        RECT 44.610 139.270 45.320 139.720 ;
        RECT 43.695 139.100 43.865 139.270 ;
        RECT 43.255 138.690 43.525 139.035 ;
        RECT 43.695 138.930 45.305 139.100 ;
        RECT 45.490 139.030 45.840 139.600 ;
        RECT 46.015 139.160 46.190 139.770 ;
        RECT 46.885 139.520 47.055 139.770 ;
        RECT 46.360 139.350 47.055 139.520 ;
        RECT 47.230 139.350 47.650 139.550 ;
        RECT 47.820 139.350 48.150 139.550 ;
        RECT 48.320 139.350 48.650 139.550 ;
        RECT 43.715 138.360 44.095 138.760 ;
        RECT 44.265 138.580 44.435 138.930 ;
        RECT 44.605 138.360 44.935 138.760 ;
        RECT 45.135 138.580 45.305 138.930 ;
        RECT 45.505 138.360 45.835 138.860 ;
        RECT 46.015 138.530 46.355 139.160 ;
        RECT 46.525 138.360 46.775 139.160 ;
        RECT 46.965 139.010 48.190 139.180 ;
        RECT 46.965 138.530 47.295 139.010 ;
        RECT 47.465 138.360 47.690 138.820 ;
        RECT 47.860 138.530 48.190 139.010 ;
        RECT 48.820 139.140 48.990 139.770 ;
        RECT 49.175 139.350 49.525 139.600 ;
        RECT 49.695 139.210 49.870 139.770 ;
        RECT 50.565 139.520 50.735 139.770 ;
        RECT 50.040 139.350 50.735 139.520 ;
        RECT 50.910 139.350 51.330 139.550 ;
        RECT 51.500 139.350 51.830 139.550 ;
        RECT 52.000 139.350 52.330 139.550 ;
        RECT 49.695 139.160 49.925 139.210 ;
        RECT 48.820 138.530 49.320 139.140 ;
        RECT 49.695 138.530 50.035 139.160 ;
        RECT 50.205 138.360 50.455 139.160 ;
        RECT 50.645 139.010 51.870 139.180 ;
        RECT 50.645 138.530 50.975 139.010 ;
        RECT 51.145 138.360 51.370 138.820 ;
        RECT 51.540 138.530 51.870 139.010 ;
        RECT 52.500 139.140 52.670 139.770 ;
        RECT 52.855 139.350 53.205 139.600 ;
        RECT 53.375 139.300 54.585 139.820 ;
        RECT 52.500 138.530 53.000 139.140 ;
        RECT 54.755 139.130 55.965 139.650 ;
        RECT 56.135 139.340 56.475 140.150 ;
        RECT 57.225 139.905 57.395 140.570 ;
        RECT 57.790 140.230 58.915 140.400 ;
        RECT 56.645 139.715 57.395 139.905 ;
        RECT 57.565 139.890 58.575 140.060 ;
        RECT 56.135 139.170 57.365 139.340 ;
        RECT 53.375 138.360 55.965 139.130 ;
        RECT 56.410 138.565 56.655 139.170 ;
        RECT 56.875 138.360 57.385 138.895 ;
        RECT 57.565 138.530 57.755 139.890 ;
        RECT 57.925 139.550 58.200 139.690 ;
        RECT 57.925 139.380 58.205 139.550 ;
        RECT 57.925 138.530 58.200 139.380 ;
        RECT 58.405 139.090 58.575 139.890 ;
        RECT 58.745 139.100 58.915 140.230 ;
        RECT 59.085 139.600 59.255 140.570 ;
        RECT 59.425 139.770 59.595 140.910 ;
        RECT 59.765 139.770 60.100 140.740 ;
        RECT 60.365 139.980 60.535 140.740 ;
        RECT 60.715 140.150 61.045 140.910 ;
        RECT 60.365 139.810 61.030 139.980 ;
        RECT 61.215 139.835 61.485 140.740 ;
        RECT 59.085 139.270 59.280 139.600 ;
        RECT 59.505 139.270 59.760 139.600 ;
        RECT 59.505 139.100 59.675 139.270 ;
        RECT 59.930 139.100 60.100 139.770 ;
        RECT 60.860 139.665 61.030 139.810 ;
        RECT 60.295 139.260 60.625 139.630 ;
        RECT 60.860 139.335 61.145 139.665 ;
        RECT 58.745 138.930 59.675 139.100 ;
        RECT 58.745 138.895 58.920 138.930 ;
        RECT 58.390 138.530 58.920 138.895 ;
        RECT 59.345 138.360 59.675 138.760 ;
        RECT 59.845 138.530 60.100 139.100 ;
        RECT 60.860 139.080 61.030 139.335 ;
        RECT 60.365 138.910 61.030 139.080 ;
        RECT 61.315 139.035 61.485 139.835 ;
        RECT 61.745 139.980 61.915 140.740 ;
        RECT 62.095 140.150 62.425 140.910 ;
        RECT 61.745 139.810 62.410 139.980 ;
        RECT 62.595 139.835 62.865 140.740 ;
        RECT 62.240 139.665 62.410 139.810 ;
        RECT 61.675 139.260 62.005 139.630 ;
        RECT 62.240 139.335 62.525 139.665 ;
        RECT 62.240 139.080 62.410 139.335 ;
        RECT 60.365 138.530 60.535 138.910 ;
        RECT 60.715 138.360 61.045 138.740 ;
        RECT 61.225 138.530 61.485 139.035 ;
        RECT 61.745 138.910 62.410 139.080 ;
        RECT 62.695 139.035 62.865 139.835 ;
        RECT 63.035 139.820 66.545 140.910 ;
        RECT 63.035 139.300 64.725 139.820 ;
        RECT 66.715 139.745 67.005 140.910 ;
        RECT 67.635 139.820 69.305 140.910 ;
        RECT 64.895 139.130 66.545 139.650 ;
        RECT 67.635 139.300 68.385 139.820 ;
        RECT 69.475 139.770 69.745 140.740 ;
        RECT 69.955 140.110 70.235 140.910 ;
        RECT 70.405 140.400 72.060 140.690 ;
        RECT 70.470 140.060 72.060 140.230 ;
        RECT 70.470 139.940 70.640 140.060 ;
        RECT 69.915 139.770 70.640 139.940 ;
        RECT 68.555 139.130 69.305 139.650 ;
        RECT 61.745 138.530 61.915 138.910 ;
        RECT 62.095 138.360 62.425 138.740 ;
        RECT 62.605 138.530 62.865 139.035 ;
        RECT 63.035 138.360 66.545 139.130 ;
        RECT 66.715 138.360 67.005 139.085 ;
        RECT 67.635 138.360 69.305 139.130 ;
        RECT 69.475 139.035 69.645 139.770 ;
        RECT 69.915 139.600 70.085 139.770 ;
        RECT 69.815 139.270 70.085 139.600 ;
        RECT 70.255 139.270 70.660 139.600 ;
        RECT 70.830 139.270 71.540 139.890 ;
        RECT 71.740 139.770 72.060 140.060 ;
        RECT 72.235 139.770 72.505 140.740 ;
        RECT 72.715 140.110 72.995 140.910 ;
        RECT 73.165 140.400 74.820 140.690 ;
        RECT 75.460 140.475 80.805 140.910 ;
        RECT 81.350 140.570 81.605 140.600 ;
        RECT 73.230 140.060 74.820 140.230 ;
        RECT 73.230 139.940 73.400 140.060 ;
        RECT 72.675 139.770 73.400 139.940 ;
        RECT 69.915 139.100 70.085 139.270 ;
        RECT 69.475 138.690 69.745 139.035 ;
        RECT 69.915 138.930 71.525 139.100 ;
        RECT 71.710 139.030 72.060 139.600 ;
        RECT 72.235 139.035 72.405 139.770 ;
        RECT 72.675 139.600 72.845 139.770 ;
        RECT 73.590 139.720 74.305 139.890 ;
        RECT 74.500 139.770 74.820 140.060 ;
        RECT 72.575 139.270 72.845 139.600 ;
        RECT 73.015 139.270 73.420 139.600 ;
        RECT 73.590 139.270 74.300 139.720 ;
        RECT 72.675 139.100 72.845 139.270 ;
        RECT 69.935 138.360 70.315 138.760 ;
        RECT 70.485 138.580 70.655 138.930 ;
        RECT 70.825 138.360 71.155 138.760 ;
        RECT 71.355 138.580 71.525 138.930 ;
        RECT 71.725 138.360 72.055 138.860 ;
        RECT 72.235 138.690 72.505 139.035 ;
        RECT 72.675 138.930 74.285 139.100 ;
        RECT 74.470 139.030 74.820 139.600 ;
        RECT 77.050 139.225 77.400 140.475 ;
        RECT 81.265 140.400 81.605 140.570 ;
        RECT 81.350 139.930 81.605 140.400 ;
        RECT 81.785 140.110 82.070 140.910 ;
        RECT 82.250 140.190 82.580 140.700 ;
        RECT 72.695 138.360 73.075 138.760 ;
        RECT 73.245 138.580 73.415 138.930 ;
        RECT 73.585 138.360 73.915 138.760 ;
        RECT 74.115 138.580 74.285 138.930 ;
        RECT 78.880 138.905 79.220 139.735 ;
        RECT 81.350 139.070 81.530 139.930 ;
        RECT 82.250 139.600 82.500 140.190 ;
        RECT 82.850 140.040 83.020 140.650 ;
        RECT 83.190 140.220 83.520 140.910 ;
        RECT 83.750 140.360 83.990 140.650 ;
        RECT 84.190 140.530 84.610 140.910 ;
        RECT 84.790 140.440 85.420 140.690 ;
        RECT 85.890 140.530 86.220 140.910 ;
        RECT 84.790 140.360 84.960 140.440 ;
        RECT 86.390 140.360 86.560 140.650 ;
        RECT 86.740 140.530 87.120 140.910 ;
        RECT 87.360 140.525 88.190 140.695 ;
        RECT 83.750 140.190 84.960 140.360 ;
        RECT 81.700 139.270 82.500 139.600 ;
        RECT 74.485 138.360 74.815 138.860 ;
        RECT 75.460 138.360 80.805 138.905 ;
        RECT 81.350 138.540 81.605 139.070 ;
        RECT 81.785 138.360 82.070 138.820 ;
        RECT 82.250 138.620 82.500 139.270 ;
        RECT 82.700 140.020 83.020 140.040 ;
        RECT 82.700 139.850 84.620 140.020 ;
        RECT 82.700 138.955 82.890 139.850 ;
        RECT 84.790 139.680 84.960 140.190 ;
        RECT 85.130 139.930 85.650 140.240 ;
        RECT 83.060 139.510 84.960 139.680 ;
        RECT 83.060 139.450 83.390 139.510 ;
        RECT 83.540 139.280 83.870 139.340 ;
        RECT 83.210 139.010 83.870 139.280 ;
        RECT 82.700 138.625 83.020 138.955 ;
        RECT 83.200 138.360 83.860 138.840 ;
        RECT 84.060 138.750 84.230 139.510 ;
        RECT 85.130 139.340 85.310 139.750 ;
        RECT 84.400 139.170 84.730 139.290 ;
        RECT 85.480 139.170 85.650 139.930 ;
        RECT 84.400 139.000 85.650 139.170 ;
        RECT 85.820 140.110 87.190 140.360 ;
        RECT 85.820 139.340 86.010 140.110 ;
        RECT 86.940 139.850 87.190 140.110 ;
        RECT 86.180 139.680 86.430 139.840 ;
        RECT 87.360 139.680 87.530 140.525 ;
        RECT 88.425 140.240 88.595 140.740 ;
        RECT 88.765 140.410 89.095 140.910 ;
        RECT 87.700 139.850 88.200 140.230 ;
        RECT 88.425 140.070 89.120 140.240 ;
        RECT 86.180 139.510 87.530 139.680 ;
        RECT 87.110 139.470 87.530 139.510 ;
        RECT 85.820 139.000 86.240 139.340 ;
        RECT 86.530 139.010 86.940 139.340 ;
        RECT 84.060 138.580 84.910 138.750 ;
        RECT 85.470 138.360 85.790 138.820 ;
        RECT 85.990 138.570 86.240 139.000 ;
        RECT 86.530 138.360 86.940 138.800 ;
        RECT 87.110 138.740 87.280 139.470 ;
        RECT 87.450 138.920 87.800 139.290 ;
        RECT 87.980 138.980 88.200 139.850 ;
        RECT 88.370 139.280 88.780 139.900 ;
        RECT 88.950 139.100 89.120 140.070 ;
        RECT 88.425 138.910 89.120 139.100 ;
        RECT 87.110 138.540 88.125 138.740 ;
        RECT 88.425 138.580 88.595 138.910 ;
        RECT 88.765 138.360 89.095 138.740 ;
        RECT 89.310 138.620 89.535 140.740 ;
        RECT 89.705 140.410 90.035 140.910 ;
        RECT 90.205 140.240 90.375 140.740 ;
        RECT 89.710 140.070 90.375 140.240 ;
        RECT 89.710 139.080 89.940 140.070 ;
        RECT 90.110 139.250 90.460 139.900 ;
        RECT 90.635 139.820 92.305 140.910 ;
        RECT 90.635 139.300 91.385 139.820 ;
        RECT 92.475 139.745 92.765 140.910 ;
        RECT 92.935 139.820 95.525 140.910 ;
        RECT 91.555 139.130 92.305 139.650 ;
        RECT 92.935 139.300 94.145 139.820 ;
        RECT 95.755 139.770 95.965 140.910 ;
        RECT 96.135 139.760 96.465 140.740 ;
        RECT 96.635 139.770 96.865 140.910 ;
        RECT 98.085 139.980 98.255 140.740 ;
        RECT 98.435 140.150 98.765 140.910 ;
        RECT 98.085 139.810 98.750 139.980 ;
        RECT 98.935 139.835 99.205 140.740 ;
        RECT 94.315 139.130 95.525 139.650 ;
        RECT 89.710 138.910 90.375 139.080 ;
        RECT 89.705 138.360 90.035 138.740 ;
        RECT 90.205 138.620 90.375 138.910 ;
        RECT 90.635 138.360 92.305 139.130 ;
        RECT 92.475 138.360 92.765 139.085 ;
        RECT 92.935 138.360 95.525 139.130 ;
        RECT 95.755 138.360 95.965 139.180 ;
        RECT 96.135 139.160 96.385 139.760 ;
        RECT 98.580 139.665 98.750 139.810 ;
        RECT 96.555 139.350 96.885 139.600 ;
        RECT 98.015 139.260 98.345 139.630 ;
        RECT 98.580 139.335 98.865 139.665 ;
        RECT 96.135 138.530 96.465 139.160 ;
        RECT 96.635 138.360 96.865 139.180 ;
        RECT 98.580 139.080 98.750 139.335 ;
        RECT 98.085 138.910 98.750 139.080 ;
        RECT 99.035 139.035 99.205 139.835 ;
        RECT 100.295 139.820 103.805 140.910 ;
        RECT 103.980 140.475 109.325 140.910 ;
        RECT 100.295 139.300 101.985 139.820 ;
        RECT 102.155 139.130 103.805 139.650 ;
        RECT 105.570 139.225 105.920 140.475 ;
        RECT 109.535 139.770 109.765 140.910 ;
        RECT 109.935 139.760 110.265 140.740 ;
        RECT 110.435 139.770 110.645 140.910 ;
        RECT 110.965 139.980 111.135 140.740 ;
        RECT 111.315 140.150 111.645 140.910 ;
        RECT 110.965 139.810 111.630 139.980 ;
        RECT 111.815 139.835 112.085 140.740 ;
        RECT 98.085 138.530 98.255 138.910 ;
        RECT 98.435 138.360 98.765 138.740 ;
        RECT 98.945 138.530 99.205 139.035 ;
        RECT 100.295 138.360 103.805 139.130 ;
        RECT 107.400 138.905 107.740 139.735 ;
        RECT 109.515 139.350 109.845 139.600 ;
        RECT 103.980 138.360 109.325 138.905 ;
        RECT 109.535 138.360 109.765 139.180 ;
        RECT 110.015 139.160 110.265 139.760 ;
        RECT 111.460 139.665 111.630 139.810 ;
        RECT 110.895 139.260 111.225 139.630 ;
        RECT 111.460 139.335 111.745 139.665 ;
        RECT 109.935 138.530 110.265 139.160 ;
        RECT 110.435 138.360 110.645 139.180 ;
        RECT 111.460 139.080 111.630 139.335 ;
        RECT 110.965 138.910 111.630 139.080 ;
        RECT 111.915 139.035 112.085 139.835 ;
        RECT 112.255 139.820 113.465 140.910 ;
        RECT 113.635 139.820 117.145 140.910 ;
        RECT 117.315 139.820 118.525 140.910 ;
        RECT 112.255 139.280 112.775 139.820 ;
        RECT 112.945 139.110 113.465 139.650 ;
        RECT 113.635 139.300 115.325 139.820 ;
        RECT 115.495 139.130 117.145 139.650 ;
        RECT 117.315 139.280 117.835 139.820 ;
        RECT 110.965 138.530 111.135 138.910 ;
        RECT 111.315 138.360 111.645 138.740 ;
        RECT 111.825 138.530 112.085 139.035 ;
        RECT 112.255 138.360 113.465 139.110 ;
        RECT 113.635 138.360 117.145 139.130 ;
        RECT 118.005 139.110 118.525 139.650 ;
        RECT 117.315 138.360 118.525 139.110 ;
        RECT 11.430 138.190 118.610 138.360 ;
        RECT 11.515 137.440 12.725 138.190 ;
        RECT 13.730 137.480 13.985 138.010 ;
        RECT 14.165 137.730 14.450 138.190 ;
        RECT 11.515 136.900 12.035 137.440 ;
        RECT 12.205 136.730 12.725 137.270 ;
        RECT 11.515 135.640 12.725 136.730 ;
        RECT 13.730 136.620 13.910 137.480 ;
        RECT 14.630 137.280 14.880 137.930 ;
        RECT 14.080 136.950 14.880 137.280 ;
        RECT 13.730 136.150 13.985 136.620 ;
        RECT 13.645 135.980 13.985 136.150 ;
        RECT 13.730 135.950 13.985 135.980 ;
        RECT 14.165 135.640 14.450 136.440 ;
        RECT 14.630 136.360 14.880 136.950 ;
        RECT 15.080 137.595 15.400 137.925 ;
        RECT 15.580 137.710 16.240 138.190 ;
        RECT 16.440 137.800 17.290 137.970 ;
        RECT 15.080 136.700 15.270 137.595 ;
        RECT 15.590 137.270 16.250 137.540 ;
        RECT 15.920 137.210 16.250 137.270 ;
        RECT 15.440 137.040 15.770 137.100 ;
        RECT 16.440 137.040 16.610 137.800 ;
        RECT 17.850 137.730 18.170 138.190 ;
        RECT 18.370 137.550 18.620 137.980 ;
        RECT 18.910 137.750 19.320 138.190 ;
        RECT 19.490 137.810 20.505 138.010 ;
        RECT 16.780 137.380 18.030 137.550 ;
        RECT 16.780 137.260 17.110 137.380 ;
        RECT 15.440 136.870 17.340 137.040 ;
        RECT 15.080 136.530 17.000 136.700 ;
        RECT 15.080 136.510 15.400 136.530 ;
        RECT 14.630 135.850 14.960 136.360 ;
        RECT 15.230 135.900 15.400 136.510 ;
        RECT 17.170 136.360 17.340 136.870 ;
        RECT 17.510 136.800 17.690 137.210 ;
        RECT 17.860 136.620 18.030 137.380 ;
        RECT 15.570 135.640 15.900 136.330 ;
        RECT 16.130 136.190 17.340 136.360 ;
        RECT 17.510 136.310 18.030 136.620 ;
        RECT 18.200 137.210 18.620 137.550 ;
        RECT 18.910 137.210 19.320 137.540 ;
        RECT 18.200 136.440 18.390 137.210 ;
        RECT 19.490 137.080 19.660 137.810 ;
        RECT 20.805 137.640 20.975 137.970 ;
        RECT 21.145 137.810 21.475 138.190 ;
        RECT 19.830 137.260 20.180 137.630 ;
        RECT 19.490 137.040 19.910 137.080 ;
        RECT 18.560 136.870 19.910 137.040 ;
        RECT 18.560 136.710 18.810 136.870 ;
        RECT 19.320 136.440 19.570 136.700 ;
        RECT 18.200 136.190 19.570 136.440 ;
        RECT 16.130 135.900 16.370 136.190 ;
        RECT 17.170 136.110 17.340 136.190 ;
        RECT 16.570 135.640 16.990 136.020 ;
        RECT 17.170 135.860 17.800 136.110 ;
        RECT 18.270 135.640 18.600 136.020 ;
        RECT 18.770 135.900 18.940 136.190 ;
        RECT 19.740 136.025 19.910 136.870 ;
        RECT 20.360 136.700 20.580 137.570 ;
        RECT 20.805 137.450 21.500 137.640 ;
        RECT 20.080 136.320 20.580 136.700 ;
        RECT 20.750 136.650 21.160 137.270 ;
        RECT 21.330 136.480 21.500 137.450 ;
        RECT 20.805 136.310 21.500 136.480 ;
        RECT 19.120 135.640 19.500 136.020 ;
        RECT 19.740 135.855 20.570 136.025 ;
        RECT 20.805 135.810 20.975 136.310 ;
        RECT 21.145 135.640 21.475 136.140 ;
        RECT 21.690 135.810 21.915 137.930 ;
        RECT 22.085 137.810 22.415 138.190 ;
        RECT 22.585 137.640 22.755 137.930 ;
        RECT 22.090 137.470 22.755 137.640 ;
        RECT 22.090 136.480 22.320 137.470 ;
        RECT 23.475 137.420 26.065 138.190 ;
        RECT 22.490 136.650 22.840 137.300 ;
        RECT 23.475 136.730 24.685 137.250 ;
        RECT 24.855 136.900 26.065 137.420 ;
        RECT 26.235 137.515 26.495 138.020 ;
        RECT 26.675 137.810 27.005 138.190 ;
        RECT 27.185 137.640 27.355 138.020 ;
        RECT 22.090 136.310 22.755 136.480 ;
        RECT 22.085 135.640 22.415 136.140 ;
        RECT 22.585 135.810 22.755 136.310 ;
        RECT 23.475 135.640 26.065 136.730 ;
        RECT 26.235 136.715 26.405 137.515 ;
        RECT 26.690 137.470 27.355 137.640 ;
        RECT 26.690 137.215 26.860 137.470 ;
        RECT 28.075 137.465 28.365 138.190 ;
        RECT 28.535 137.440 29.745 138.190 ;
        RECT 26.575 136.885 26.860 137.215 ;
        RECT 27.095 136.920 27.425 137.290 ;
        RECT 26.690 136.740 26.860 136.885 ;
        RECT 26.235 135.810 26.505 136.715 ;
        RECT 26.690 136.570 27.355 136.740 ;
        RECT 26.675 135.640 27.005 136.400 ;
        RECT 27.185 135.810 27.355 136.570 ;
        RECT 28.075 135.640 28.365 136.805 ;
        RECT 28.535 136.730 29.055 137.270 ;
        RECT 29.225 136.900 29.745 137.440 ;
        RECT 30.115 137.560 30.445 137.920 ;
        RECT 31.065 137.730 31.315 138.190 ;
        RECT 31.485 137.730 32.045 138.020 ;
        RECT 30.115 137.370 31.505 137.560 ;
        RECT 31.335 137.280 31.505 137.370 ;
        RECT 29.930 136.950 30.605 137.200 ;
        RECT 30.825 136.950 31.165 137.200 ;
        RECT 31.335 136.950 31.625 137.280 ;
        RECT 28.535 135.640 29.745 136.730 ;
        RECT 29.930 136.590 30.195 136.950 ;
        RECT 31.335 136.700 31.505 136.950 ;
        RECT 30.565 136.530 31.505 136.700 ;
        RECT 30.115 135.640 30.395 136.310 ;
        RECT 30.565 135.980 30.865 136.530 ;
        RECT 31.795 136.360 32.045 137.730 ;
        RECT 32.415 137.560 32.745 137.920 ;
        RECT 33.365 137.730 33.615 138.190 ;
        RECT 33.785 137.730 34.345 138.020 ;
        RECT 32.415 137.370 33.805 137.560 ;
        RECT 33.635 137.280 33.805 137.370 ;
        RECT 32.230 136.950 32.905 137.200 ;
        RECT 33.125 136.950 33.465 137.200 ;
        RECT 33.635 136.950 33.925 137.280 ;
        RECT 32.230 136.590 32.495 136.950 ;
        RECT 33.635 136.700 33.805 136.950 ;
        RECT 31.065 135.640 31.395 136.360 ;
        RECT 31.585 135.810 32.045 136.360 ;
        RECT 32.865 136.530 33.805 136.700 ;
        RECT 32.415 135.640 32.695 136.310 ;
        RECT 32.865 135.980 33.165 136.530 ;
        RECT 34.095 136.360 34.345 137.730 ;
        RECT 33.365 135.640 33.695 136.360 ;
        RECT 33.885 135.810 34.345 136.360 ;
        RECT 34.515 137.730 35.075 138.020 ;
        RECT 35.245 137.730 35.495 138.190 ;
        RECT 34.515 136.360 34.765 137.730 ;
        RECT 36.115 137.560 36.445 137.920 ;
        RECT 35.055 137.370 36.445 137.560 ;
        RECT 37.015 137.560 37.345 137.920 ;
        RECT 37.965 137.730 38.215 138.190 ;
        RECT 38.385 137.730 38.945 138.020 ;
        RECT 37.015 137.370 38.405 137.560 ;
        RECT 35.055 137.280 35.225 137.370 ;
        RECT 34.935 136.950 35.225 137.280 ;
        RECT 38.235 137.280 38.405 137.370 ;
        RECT 35.395 136.950 35.735 137.200 ;
        RECT 35.955 136.950 36.630 137.200 ;
        RECT 35.055 136.700 35.225 136.950 ;
        RECT 35.055 136.530 35.995 136.700 ;
        RECT 36.365 136.590 36.630 136.950 ;
        RECT 36.830 136.950 37.505 137.200 ;
        RECT 37.725 136.950 38.065 137.200 ;
        RECT 38.235 136.950 38.525 137.280 ;
        RECT 36.830 136.590 37.095 136.950 ;
        RECT 38.235 136.700 38.405 136.950 ;
        RECT 34.515 135.810 34.975 136.360 ;
        RECT 35.165 135.640 35.495 136.360 ;
        RECT 35.695 135.980 35.995 136.530 ;
        RECT 37.465 136.530 38.405 136.700 ;
        RECT 36.165 135.640 36.445 136.310 ;
        RECT 37.015 135.640 37.295 136.310 ;
        RECT 37.465 135.980 37.765 136.530 ;
        RECT 38.695 136.360 38.945 137.730 ;
        RECT 39.115 137.420 42.625 138.190 ;
        RECT 42.800 137.645 48.145 138.190 ;
        RECT 48.320 137.645 53.665 138.190 ;
        RECT 37.965 135.640 38.295 136.360 ;
        RECT 38.485 135.810 38.945 136.360 ;
        RECT 39.115 136.730 40.805 137.250 ;
        RECT 40.975 136.900 42.625 137.420 ;
        RECT 39.115 135.640 42.625 136.730 ;
        RECT 44.390 136.075 44.740 137.325 ;
        RECT 46.220 136.815 46.560 137.645 ;
        RECT 49.910 136.075 50.260 137.325 ;
        RECT 51.740 136.815 52.080 137.645 ;
        RECT 53.835 137.465 54.125 138.190 ;
        RECT 54.755 137.420 57.345 138.190 ;
        RECT 42.800 135.640 48.145 136.075 ;
        RECT 48.320 135.640 53.665 136.075 ;
        RECT 53.835 135.640 54.125 136.805 ;
        RECT 54.755 136.730 55.965 137.250 ;
        RECT 56.135 136.900 57.345 137.420 ;
        RECT 57.790 137.380 58.035 137.985 ;
        RECT 58.255 137.655 58.765 138.190 ;
        RECT 57.515 137.210 58.745 137.380 ;
        RECT 54.755 135.640 57.345 136.730 ;
        RECT 57.515 136.400 57.855 137.210 ;
        RECT 58.025 136.645 58.775 136.835 ;
        RECT 57.515 135.990 58.030 136.400 ;
        RECT 58.265 135.640 58.435 136.400 ;
        RECT 58.605 135.980 58.775 136.645 ;
        RECT 58.945 136.660 59.135 138.020 ;
        RECT 59.305 137.850 59.580 138.020 ;
        RECT 59.305 137.680 59.585 137.850 ;
        RECT 59.305 136.860 59.580 137.680 ;
        RECT 59.770 137.655 60.300 138.020 ;
        RECT 60.725 137.790 61.055 138.190 ;
        RECT 60.125 137.620 60.300 137.655 ;
        RECT 59.785 136.660 59.955 137.460 ;
        RECT 58.945 136.490 59.955 136.660 ;
        RECT 60.125 137.450 61.055 137.620 ;
        RECT 61.225 137.450 61.480 138.020 ;
        RECT 62.665 137.640 62.835 138.020 ;
        RECT 63.015 137.810 63.345 138.190 ;
        RECT 62.665 137.470 63.330 137.640 ;
        RECT 63.525 137.515 63.785 138.020 ;
        RECT 60.125 136.320 60.295 137.450 ;
        RECT 60.885 137.280 61.055 137.450 ;
        RECT 59.170 136.150 60.295 136.320 ;
        RECT 60.465 136.950 60.660 137.280 ;
        RECT 60.885 136.950 61.140 137.280 ;
        RECT 60.465 135.980 60.635 136.950 ;
        RECT 61.310 136.780 61.480 137.450 ;
        RECT 62.595 136.920 62.925 137.290 ;
        RECT 63.160 137.215 63.330 137.470 ;
        RECT 58.605 135.810 60.635 135.980 ;
        RECT 60.805 135.640 60.975 136.780 ;
        RECT 61.145 135.810 61.480 136.780 ;
        RECT 63.160 136.885 63.445 137.215 ;
        RECT 63.160 136.740 63.330 136.885 ;
        RECT 62.665 136.570 63.330 136.740 ;
        RECT 63.615 136.715 63.785 137.515 ;
        RECT 64.505 137.640 64.675 138.020 ;
        RECT 64.855 137.810 65.185 138.190 ;
        RECT 64.505 137.470 65.170 137.640 ;
        RECT 65.365 137.515 65.625 138.020 ;
        RECT 64.435 136.920 64.765 137.290 ;
        RECT 65.000 137.215 65.170 137.470 ;
        RECT 65.000 136.885 65.285 137.215 ;
        RECT 65.000 136.740 65.170 136.885 ;
        RECT 62.665 135.810 62.835 136.570 ;
        RECT 63.015 135.640 63.345 136.400 ;
        RECT 63.515 135.810 63.785 136.715 ;
        RECT 64.505 136.570 65.170 136.740 ;
        RECT 65.455 136.715 65.625 137.515 ;
        RECT 64.505 135.810 64.675 136.570 ;
        RECT 64.855 135.640 65.185 136.400 ;
        RECT 65.355 135.810 65.625 136.715 ;
        RECT 65.795 137.690 66.055 138.020 ;
        RECT 66.265 137.710 66.540 138.190 ;
        RECT 65.795 136.780 65.965 137.690 ;
        RECT 66.750 137.620 66.955 138.020 ;
        RECT 67.125 137.790 67.460 138.190 ;
        RECT 66.135 136.950 66.495 137.530 ;
        RECT 66.750 137.450 67.435 137.620 ;
        RECT 66.675 136.780 66.925 137.280 ;
        RECT 65.795 136.610 66.925 136.780 ;
        RECT 65.795 135.840 66.065 136.610 ;
        RECT 67.095 136.420 67.435 137.450 ;
        RECT 67.635 137.420 70.225 138.190 ;
        RECT 66.235 135.640 66.565 136.420 ;
        RECT 66.770 136.245 67.435 136.420 ;
        RECT 67.635 136.730 68.845 137.250 ;
        RECT 69.015 136.900 70.225 137.420 ;
        RECT 70.595 137.560 70.925 137.920 ;
        RECT 71.545 137.730 71.795 138.190 ;
        RECT 71.965 137.730 72.525 138.020 ;
        RECT 70.595 137.370 71.985 137.560 ;
        RECT 71.815 137.280 71.985 137.370 ;
        RECT 70.410 136.950 71.085 137.200 ;
        RECT 71.305 136.950 71.645 137.200 ;
        RECT 71.815 136.950 72.105 137.280 ;
        RECT 66.770 135.840 66.955 136.245 ;
        RECT 67.125 135.640 67.460 136.065 ;
        RECT 67.635 135.640 70.225 136.730 ;
        RECT 70.410 136.590 70.675 136.950 ;
        RECT 71.815 136.700 71.985 136.950 ;
        RECT 71.045 136.530 71.985 136.700 ;
        RECT 70.595 135.640 70.875 136.310 ;
        RECT 71.045 135.980 71.345 136.530 ;
        RECT 72.275 136.360 72.525 137.730 ;
        RECT 71.545 135.640 71.875 136.360 ;
        RECT 72.065 135.810 72.525 136.360 ;
        RECT 72.695 137.730 73.255 138.020 ;
        RECT 73.425 137.730 73.675 138.190 ;
        RECT 72.695 136.360 72.945 137.730 ;
        RECT 74.295 137.560 74.625 137.920 ;
        RECT 73.235 137.370 74.625 137.560 ;
        RECT 75.915 137.420 79.425 138.190 ;
        RECT 79.595 137.465 79.885 138.190 ;
        RECT 80.515 137.420 83.105 138.190 ;
        RECT 73.235 137.280 73.405 137.370 ;
        RECT 73.115 136.950 73.405 137.280 ;
        RECT 73.575 136.950 73.915 137.200 ;
        RECT 74.135 136.950 74.810 137.200 ;
        RECT 73.235 136.700 73.405 136.950 ;
        RECT 73.235 136.530 74.175 136.700 ;
        RECT 74.545 136.590 74.810 136.950 ;
        RECT 75.915 136.730 77.605 137.250 ;
        RECT 77.775 136.900 79.425 137.420 ;
        RECT 72.695 135.810 73.155 136.360 ;
        RECT 73.345 135.640 73.675 136.360 ;
        RECT 73.875 135.980 74.175 136.530 ;
        RECT 74.345 135.640 74.625 136.310 ;
        RECT 75.915 135.640 79.425 136.730 ;
        RECT 79.595 135.640 79.885 136.805 ;
        RECT 80.515 136.730 81.725 137.250 ;
        RECT 81.895 136.900 83.105 137.420 ;
        RECT 83.335 137.370 83.545 138.190 ;
        RECT 83.715 137.390 84.045 138.020 ;
        RECT 83.715 136.790 83.965 137.390 ;
        RECT 84.215 137.370 84.445 138.190 ;
        RECT 85.635 137.370 85.845 138.190 ;
        RECT 86.015 137.390 86.345 138.020 ;
        RECT 84.135 136.950 84.465 137.200 ;
        RECT 86.015 136.790 86.265 137.390 ;
        RECT 86.515 137.370 86.745 138.190 ;
        RECT 86.955 137.420 90.465 138.190 ;
        RECT 86.435 136.950 86.765 137.200 ;
        RECT 80.515 135.640 83.105 136.730 ;
        RECT 83.335 135.640 83.545 136.780 ;
        RECT 83.715 135.810 84.045 136.790 ;
        RECT 84.215 135.640 84.445 136.780 ;
        RECT 85.635 135.640 85.845 136.780 ;
        RECT 86.015 135.810 86.345 136.790 ;
        RECT 86.515 135.640 86.745 136.780 ;
        RECT 86.955 136.730 88.645 137.250 ;
        RECT 88.815 136.900 90.465 137.420 ;
        RECT 90.910 137.380 91.155 137.985 ;
        RECT 91.375 137.655 91.885 138.190 ;
        RECT 90.635 137.210 91.865 137.380 ;
        RECT 86.955 135.640 90.465 136.730 ;
        RECT 90.635 136.400 90.975 137.210 ;
        RECT 91.145 136.645 91.895 136.835 ;
        RECT 90.635 135.990 91.150 136.400 ;
        RECT 91.385 135.640 91.555 136.400 ;
        RECT 91.725 135.980 91.895 136.645 ;
        RECT 92.065 136.660 92.255 138.020 ;
        RECT 92.425 137.510 92.700 138.020 ;
        RECT 92.890 137.655 93.420 138.020 ;
        RECT 93.845 137.790 94.175 138.190 ;
        RECT 93.245 137.620 93.420 137.655 ;
        RECT 92.425 137.340 92.705 137.510 ;
        RECT 92.425 136.860 92.700 137.340 ;
        RECT 92.905 136.660 93.075 137.460 ;
        RECT 92.065 136.490 93.075 136.660 ;
        RECT 93.245 137.450 94.175 137.620 ;
        RECT 94.345 137.450 94.600 138.020 ;
        RECT 93.245 136.320 93.415 137.450 ;
        RECT 94.005 137.280 94.175 137.450 ;
        RECT 92.290 136.150 93.415 136.320 ;
        RECT 93.585 136.950 93.780 137.280 ;
        RECT 94.005 136.950 94.260 137.280 ;
        RECT 93.585 135.980 93.755 136.950 ;
        RECT 94.430 136.780 94.600 137.450 ;
        RECT 91.725 135.810 93.755 135.980 ;
        RECT 93.925 135.640 94.095 136.780 ;
        RECT 94.265 135.810 94.600 136.780 ;
        RECT 95.695 137.515 95.955 138.020 ;
        RECT 96.135 137.810 96.465 138.190 ;
        RECT 96.645 137.640 96.815 138.020 ;
        RECT 95.695 136.715 95.865 137.515 ;
        RECT 96.150 137.470 96.815 137.640 ;
        RECT 97.075 137.730 97.635 138.020 ;
        RECT 97.805 137.730 98.055 138.190 ;
        RECT 96.150 137.215 96.320 137.470 ;
        RECT 96.035 136.885 96.320 137.215 ;
        RECT 96.555 136.920 96.885 137.290 ;
        RECT 96.150 136.740 96.320 136.885 ;
        RECT 95.695 135.810 95.965 136.715 ;
        RECT 96.150 136.570 96.815 136.740 ;
        RECT 96.135 135.640 96.465 136.400 ;
        RECT 96.645 135.810 96.815 136.570 ;
        RECT 97.075 136.360 97.325 137.730 ;
        RECT 98.675 137.560 99.005 137.920 ;
        RECT 97.615 137.370 99.005 137.560 ;
        RECT 99.375 137.420 101.965 138.190 ;
        RECT 97.615 137.280 97.785 137.370 ;
        RECT 97.495 136.950 97.785 137.280 ;
        RECT 97.955 136.950 98.295 137.200 ;
        RECT 98.515 136.950 99.190 137.200 ;
        RECT 97.615 136.700 97.785 136.950 ;
        RECT 97.615 136.530 98.555 136.700 ;
        RECT 98.925 136.590 99.190 136.950 ;
        RECT 99.375 136.730 100.585 137.250 ;
        RECT 100.755 136.900 101.965 137.420 ;
        RECT 102.135 137.730 102.695 138.020 ;
        RECT 102.865 137.730 103.115 138.190 ;
        RECT 97.075 135.810 97.535 136.360 ;
        RECT 97.725 135.640 98.055 136.360 ;
        RECT 98.255 135.980 98.555 136.530 ;
        RECT 98.725 135.640 99.005 136.310 ;
        RECT 99.375 135.640 101.965 136.730 ;
        RECT 102.135 136.360 102.385 137.730 ;
        RECT 103.735 137.560 104.065 137.920 ;
        RECT 102.675 137.370 104.065 137.560 ;
        RECT 105.355 137.465 105.645 138.190 ;
        RECT 106.650 137.480 106.905 138.010 ;
        RECT 107.085 137.730 107.370 138.190 ;
        RECT 102.675 137.280 102.845 137.370 ;
        RECT 102.555 136.950 102.845 137.280 ;
        RECT 103.015 136.950 103.355 137.200 ;
        RECT 103.575 136.950 104.250 137.200 ;
        RECT 102.675 136.700 102.845 136.950 ;
        RECT 102.675 136.530 103.615 136.700 ;
        RECT 103.985 136.590 104.250 136.950 ;
        RECT 106.650 136.830 106.830 137.480 ;
        RECT 107.550 137.280 107.800 137.930 ;
        RECT 107.000 136.950 107.800 137.280 ;
        RECT 102.135 135.810 102.595 136.360 ;
        RECT 102.785 135.640 103.115 136.360 ;
        RECT 103.315 135.980 103.615 136.530 ;
        RECT 103.785 135.640 104.065 136.310 ;
        RECT 105.355 135.640 105.645 136.805 ;
        RECT 106.565 136.660 106.830 136.830 ;
        RECT 106.650 136.620 106.830 136.660 ;
        RECT 106.650 135.950 106.905 136.620 ;
        RECT 107.085 135.640 107.370 136.440 ;
        RECT 107.550 136.360 107.800 136.950 ;
        RECT 108.000 137.595 108.320 137.925 ;
        RECT 108.500 137.710 109.160 138.190 ;
        RECT 109.360 137.800 110.210 137.970 ;
        RECT 108.000 136.700 108.190 137.595 ;
        RECT 108.510 137.270 109.170 137.540 ;
        RECT 108.840 137.210 109.170 137.270 ;
        RECT 108.360 137.040 108.690 137.100 ;
        RECT 109.360 137.040 109.530 137.800 ;
        RECT 110.770 137.730 111.090 138.190 ;
        RECT 111.290 137.550 111.540 137.980 ;
        RECT 111.830 137.750 112.240 138.190 ;
        RECT 112.410 137.810 113.425 138.010 ;
        RECT 109.700 137.380 110.950 137.550 ;
        RECT 109.700 137.260 110.030 137.380 ;
        RECT 108.360 136.870 110.260 137.040 ;
        RECT 108.000 136.530 109.920 136.700 ;
        RECT 108.000 136.510 108.320 136.530 ;
        RECT 107.550 135.850 107.880 136.360 ;
        RECT 108.150 135.900 108.320 136.510 ;
        RECT 110.090 136.360 110.260 136.870 ;
        RECT 110.430 136.800 110.610 137.210 ;
        RECT 110.780 136.620 110.950 137.380 ;
        RECT 108.490 135.640 108.820 136.330 ;
        RECT 109.050 136.190 110.260 136.360 ;
        RECT 110.430 136.310 110.950 136.620 ;
        RECT 111.120 137.210 111.540 137.550 ;
        RECT 111.830 137.210 112.240 137.540 ;
        RECT 111.120 136.440 111.310 137.210 ;
        RECT 112.410 137.080 112.580 137.810 ;
        RECT 113.725 137.640 113.895 137.970 ;
        RECT 114.065 137.810 114.395 138.190 ;
        RECT 112.750 137.260 113.100 137.630 ;
        RECT 112.410 137.040 112.830 137.080 ;
        RECT 111.480 136.870 112.830 137.040 ;
        RECT 111.480 136.710 111.730 136.870 ;
        RECT 112.240 136.440 112.490 136.700 ;
        RECT 111.120 136.190 112.490 136.440 ;
        RECT 109.050 135.900 109.290 136.190 ;
        RECT 110.090 136.110 110.260 136.190 ;
        RECT 109.490 135.640 109.910 136.020 ;
        RECT 110.090 135.860 110.720 136.110 ;
        RECT 111.190 135.640 111.520 136.020 ;
        RECT 111.690 135.900 111.860 136.190 ;
        RECT 112.660 136.025 112.830 136.870 ;
        RECT 113.280 136.700 113.500 137.570 ;
        RECT 113.725 137.450 114.420 137.640 ;
        RECT 113.000 136.320 113.500 136.700 ;
        RECT 113.670 136.650 114.080 137.270 ;
        RECT 114.250 136.480 114.420 137.450 ;
        RECT 113.725 136.310 114.420 136.480 ;
        RECT 112.040 135.640 112.420 136.020 ;
        RECT 112.660 135.855 113.490 136.025 ;
        RECT 113.725 135.810 113.895 136.310 ;
        RECT 114.065 135.640 114.395 136.140 ;
        RECT 114.610 135.810 114.835 137.930 ;
        RECT 115.005 137.810 115.335 138.190 ;
        RECT 115.505 137.640 115.675 137.930 ;
        RECT 115.010 137.470 115.675 137.640 ;
        RECT 115.010 136.480 115.240 137.470 ;
        RECT 115.935 137.440 117.145 138.190 ;
        RECT 117.315 137.440 118.525 138.190 ;
        RECT 115.410 136.650 115.760 137.300 ;
        RECT 115.935 136.730 116.455 137.270 ;
        RECT 116.625 136.900 117.145 137.440 ;
        RECT 117.315 136.730 117.835 137.270 ;
        RECT 118.005 136.900 118.525 137.440 ;
        RECT 115.010 136.310 115.675 136.480 ;
        RECT 115.005 135.640 115.335 136.140 ;
        RECT 115.505 135.810 115.675 136.310 ;
        RECT 115.935 135.640 117.145 136.730 ;
        RECT 117.315 135.640 118.525 136.730 ;
        RECT 11.430 135.470 118.610 135.640 ;
        RECT 11.515 134.380 12.725 135.470 ;
        RECT 11.515 133.670 12.035 134.210 ;
        RECT 12.205 133.840 12.725 134.380 ;
        RECT 13.875 134.330 14.085 135.470 ;
        RECT 14.255 134.320 14.585 135.300 ;
        RECT 14.755 134.330 14.985 135.470 ;
        RECT 11.515 132.920 12.725 133.670 ;
        RECT 13.875 132.920 14.085 133.740 ;
        RECT 14.255 133.720 14.505 134.320 ;
        RECT 15.195 134.305 15.485 135.470 ;
        RECT 15.695 134.330 15.925 135.470 ;
        RECT 16.095 134.320 16.425 135.300 ;
        RECT 16.595 134.330 16.805 135.470 ;
        RECT 17.125 134.540 17.295 135.300 ;
        RECT 17.475 134.710 17.805 135.470 ;
        RECT 17.125 134.370 17.790 134.540 ;
        RECT 17.975 134.395 18.245 135.300 ;
        RECT 14.675 133.910 15.005 134.160 ;
        RECT 15.675 133.910 16.005 134.160 ;
        RECT 14.255 133.090 14.585 133.720 ;
        RECT 14.755 132.920 14.985 133.740 ;
        RECT 15.195 132.920 15.485 133.645 ;
        RECT 15.695 132.920 15.925 133.740 ;
        RECT 16.175 133.720 16.425 134.320 ;
        RECT 17.620 134.225 17.790 134.370 ;
        RECT 17.055 133.820 17.385 134.190 ;
        RECT 17.620 133.895 17.905 134.225 ;
        RECT 16.095 133.090 16.425 133.720 ;
        RECT 16.595 132.920 16.805 133.740 ;
        RECT 17.620 133.640 17.790 133.895 ;
        RECT 17.125 133.470 17.790 133.640 ;
        RECT 18.075 133.595 18.245 134.395 ;
        RECT 17.125 133.090 17.295 133.470 ;
        RECT 17.475 132.920 17.805 133.300 ;
        RECT 17.985 133.090 18.245 133.595 ;
        RECT 18.790 134.490 19.045 135.160 ;
        RECT 19.225 134.670 19.510 135.470 ;
        RECT 19.690 134.750 20.020 135.260 ;
        RECT 18.790 133.630 18.970 134.490 ;
        RECT 19.690 134.160 19.940 134.750 ;
        RECT 20.290 134.600 20.460 135.210 ;
        RECT 20.630 134.780 20.960 135.470 ;
        RECT 21.190 134.920 21.430 135.210 ;
        RECT 21.630 135.090 22.050 135.470 ;
        RECT 22.230 135.000 22.860 135.250 ;
        RECT 23.330 135.090 23.660 135.470 ;
        RECT 22.230 134.920 22.400 135.000 ;
        RECT 23.830 134.920 24.000 135.210 ;
        RECT 24.180 135.090 24.560 135.470 ;
        RECT 24.800 135.085 25.630 135.255 ;
        RECT 21.190 134.750 22.400 134.920 ;
        RECT 19.140 133.830 19.940 134.160 ;
        RECT 18.790 133.430 19.045 133.630 ;
        RECT 18.705 133.260 19.045 133.430 ;
        RECT 18.790 133.100 19.045 133.260 ;
        RECT 19.225 132.920 19.510 133.380 ;
        RECT 19.690 133.180 19.940 133.830 ;
        RECT 20.140 134.580 20.460 134.600 ;
        RECT 20.140 134.410 22.060 134.580 ;
        RECT 20.140 133.515 20.330 134.410 ;
        RECT 22.230 134.240 22.400 134.750 ;
        RECT 22.570 134.490 23.090 134.800 ;
        RECT 20.500 134.070 22.400 134.240 ;
        RECT 20.500 134.010 20.830 134.070 ;
        RECT 20.980 133.840 21.310 133.900 ;
        RECT 20.650 133.570 21.310 133.840 ;
        RECT 20.140 133.185 20.460 133.515 ;
        RECT 20.640 132.920 21.300 133.400 ;
        RECT 21.500 133.310 21.670 134.070 ;
        RECT 22.570 133.900 22.750 134.310 ;
        RECT 21.840 133.730 22.170 133.850 ;
        RECT 22.920 133.730 23.090 134.490 ;
        RECT 21.840 133.560 23.090 133.730 ;
        RECT 23.260 134.670 24.630 134.920 ;
        RECT 23.260 133.900 23.450 134.670 ;
        RECT 24.380 134.410 24.630 134.670 ;
        RECT 23.620 134.240 23.870 134.400 ;
        RECT 24.800 134.240 24.970 135.085 ;
        RECT 25.865 134.800 26.035 135.300 ;
        RECT 26.205 134.970 26.535 135.470 ;
        RECT 25.140 134.410 25.640 134.790 ;
        RECT 25.865 134.630 26.560 134.800 ;
        RECT 23.620 134.070 24.970 134.240 ;
        RECT 24.550 134.030 24.970 134.070 ;
        RECT 23.260 133.560 23.680 133.900 ;
        RECT 23.970 133.570 24.380 133.900 ;
        RECT 21.500 133.140 22.350 133.310 ;
        RECT 22.910 132.920 23.230 133.380 ;
        RECT 23.430 133.130 23.680 133.560 ;
        RECT 23.970 132.920 24.380 133.360 ;
        RECT 24.550 133.300 24.720 134.030 ;
        RECT 24.890 133.480 25.240 133.850 ;
        RECT 25.420 133.540 25.640 134.410 ;
        RECT 25.810 133.840 26.220 134.460 ;
        RECT 26.390 133.660 26.560 134.630 ;
        RECT 25.865 133.470 26.560 133.660 ;
        RECT 24.550 133.100 25.565 133.300 ;
        RECT 25.865 133.140 26.035 133.470 ;
        RECT 26.205 132.920 26.535 133.300 ;
        RECT 26.750 133.180 26.975 135.300 ;
        RECT 27.145 134.970 27.475 135.470 ;
        RECT 27.645 134.800 27.815 135.300 ;
        RECT 27.150 134.630 27.815 134.800 ;
        RECT 27.150 133.640 27.380 134.630 ;
        RECT 27.550 133.810 27.900 134.460 ;
        RECT 28.080 134.330 28.415 135.300 ;
        RECT 28.585 134.330 28.755 135.470 ;
        RECT 28.925 135.130 30.955 135.300 ;
        RECT 28.080 133.660 28.250 134.330 ;
        RECT 28.925 134.160 29.095 135.130 ;
        RECT 28.420 133.830 28.675 134.160 ;
        RECT 28.900 133.830 29.095 134.160 ;
        RECT 29.265 134.790 30.390 134.960 ;
        RECT 28.505 133.660 28.675 133.830 ;
        RECT 29.265 133.660 29.435 134.790 ;
        RECT 27.150 133.470 27.815 133.640 ;
        RECT 27.145 132.920 27.475 133.300 ;
        RECT 27.645 133.180 27.815 133.470 ;
        RECT 28.080 133.090 28.335 133.660 ;
        RECT 28.505 133.490 29.435 133.660 ;
        RECT 29.605 134.450 30.615 134.620 ;
        RECT 29.605 133.650 29.775 134.450 ;
        RECT 29.980 134.110 30.255 134.250 ;
        RECT 29.975 133.940 30.255 134.110 ;
        RECT 29.260 133.455 29.435 133.490 ;
        RECT 28.505 132.920 28.835 133.320 ;
        RECT 29.260 133.090 29.790 133.455 ;
        RECT 29.980 133.090 30.255 133.940 ;
        RECT 30.425 133.090 30.615 134.450 ;
        RECT 30.785 134.465 30.955 135.130 ;
        RECT 31.125 134.710 31.295 135.470 ;
        RECT 31.530 134.710 32.045 135.120 ;
        RECT 30.785 134.275 31.535 134.465 ;
        RECT 31.705 133.900 32.045 134.710 ;
        RECT 30.815 133.730 32.045 133.900 ;
        RECT 32.675 134.710 33.190 135.120 ;
        RECT 33.425 134.710 33.595 135.470 ;
        RECT 33.765 135.130 35.795 135.300 ;
        RECT 32.675 133.900 33.015 134.710 ;
        RECT 33.765 134.465 33.935 135.130 ;
        RECT 34.330 134.790 35.455 134.960 ;
        RECT 33.185 134.275 33.935 134.465 ;
        RECT 34.105 134.450 35.115 134.620 ;
        RECT 32.675 133.730 33.905 133.900 ;
        RECT 30.795 132.920 31.305 133.455 ;
        RECT 31.525 133.125 31.770 133.730 ;
        RECT 32.950 133.125 33.195 133.730 ;
        RECT 33.415 132.920 33.925 133.455 ;
        RECT 34.105 133.090 34.295 134.450 ;
        RECT 34.465 133.430 34.740 134.250 ;
        RECT 34.945 133.650 35.115 134.450 ;
        RECT 35.285 133.660 35.455 134.790 ;
        RECT 35.625 134.160 35.795 135.130 ;
        RECT 35.965 134.330 36.135 135.470 ;
        RECT 36.305 134.330 36.640 135.300 ;
        RECT 35.625 133.830 35.820 134.160 ;
        RECT 36.045 133.830 36.300 134.160 ;
        RECT 36.045 133.660 36.215 133.830 ;
        RECT 36.470 133.660 36.640 134.330 ;
        RECT 36.815 134.380 38.485 135.470 ;
        RECT 38.655 134.750 39.115 135.300 ;
        RECT 39.305 134.750 39.635 135.470 ;
        RECT 36.815 133.860 37.565 134.380 ;
        RECT 37.735 133.690 38.485 134.210 ;
        RECT 35.285 133.490 36.215 133.660 ;
        RECT 35.285 133.455 35.460 133.490 ;
        RECT 34.465 133.260 34.745 133.430 ;
        RECT 34.465 133.090 34.740 133.260 ;
        RECT 34.930 133.090 35.460 133.455 ;
        RECT 35.885 132.920 36.215 133.320 ;
        RECT 36.385 133.090 36.640 133.660 ;
        RECT 36.815 132.920 38.485 133.690 ;
        RECT 38.655 133.380 38.905 134.750 ;
        RECT 39.835 134.580 40.135 135.130 ;
        RECT 40.305 134.800 40.585 135.470 ;
        RECT 39.195 134.410 40.135 134.580 ;
        RECT 39.195 134.160 39.365 134.410 ;
        RECT 40.505 134.160 40.770 134.520 ;
        RECT 40.955 134.305 41.245 135.470 ;
        RECT 41.615 134.800 41.895 135.470 ;
        RECT 42.065 134.580 42.365 135.130 ;
        RECT 42.565 134.750 42.895 135.470 ;
        RECT 43.085 134.750 43.545 135.300 ;
        RECT 43.915 134.800 44.195 135.470 ;
        RECT 39.075 133.830 39.365 134.160 ;
        RECT 39.535 133.910 39.875 134.160 ;
        RECT 40.095 133.910 40.770 134.160 ;
        RECT 41.430 134.160 41.695 134.520 ;
        RECT 42.065 134.410 43.005 134.580 ;
        RECT 42.835 134.160 43.005 134.410 ;
        RECT 41.430 133.910 42.105 134.160 ;
        RECT 42.325 133.910 42.665 134.160 ;
        RECT 39.195 133.740 39.365 133.830 ;
        RECT 42.835 133.830 43.125 134.160 ;
        RECT 42.835 133.740 43.005 133.830 ;
        RECT 39.195 133.550 40.585 133.740 ;
        RECT 38.655 133.090 39.215 133.380 ;
        RECT 39.385 132.920 39.635 133.380 ;
        RECT 40.255 133.190 40.585 133.550 ;
        RECT 40.955 132.920 41.245 133.645 ;
        RECT 41.615 133.550 43.005 133.740 ;
        RECT 41.615 133.190 41.945 133.550 ;
        RECT 43.295 133.380 43.545 134.750 ;
        RECT 44.365 134.580 44.665 135.130 ;
        RECT 44.865 134.750 45.195 135.470 ;
        RECT 45.385 134.750 45.845 135.300 ;
        RECT 43.730 134.160 43.995 134.520 ;
        RECT 44.365 134.410 45.305 134.580 ;
        RECT 45.135 134.160 45.305 134.410 ;
        RECT 43.730 133.910 44.405 134.160 ;
        RECT 44.625 133.910 44.965 134.160 ;
        RECT 45.135 133.830 45.425 134.160 ;
        RECT 45.135 133.740 45.305 133.830 ;
        RECT 42.565 132.920 42.815 133.380 ;
        RECT 42.985 133.090 43.545 133.380 ;
        RECT 43.915 133.550 45.305 133.740 ;
        RECT 43.915 133.190 44.245 133.550 ;
        RECT 45.595 133.380 45.845 134.750 ;
        RECT 44.865 132.920 45.115 133.380 ;
        RECT 45.285 133.090 45.845 133.380 ;
        RECT 46.015 134.750 46.475 135.300 ;
        RECT 46.665 134.750 46.995 135.470 ;
        RECT 46.015 133.380 46.265 134.750 ;
        RECT 47.195 134.580 47.495 135.130 ;
        RECT 47.665 134.800 47.945 135.470 ;
        RECT 46.555 134.410 47.495 134.580 ;
        RECT 46.555 134.160 46.725 134.410 ;
        RECT 47.865 134.160 48.130 134.520 ;
        RECT 46.435 133.830 46.725 134.160 ;
        RECT 46.895 133.910 47.235 134.160 ;
        RECT 47.455 133.910 48.130 134.160 ;
        RECT 48.315 134.380 49.985 135.470 ;
        RECT 50.160 135.035 55.505 135.470 ;
        RECT 48.315 133.860 49.065 134.380 ;
        RECT 46.555 133.740 46.725 133.830 ;
        RECT 46.555 133.550 47.945 133.740 ;
        RECT 49.235 133.690 49.985 134.210 ;
        RECT 51.750 133.785 52.100 135.035 ;
        RECT 55.735 134.330 55.945 135.470 ;
        RECT 56.115 134.320 56.445 135.300 ;
        RECT 56.615 134.330 56.845 135.470 ;
        RECT 57.430 135.130 57.685 135.160 ;
        RECT 57.345 134.960 57.685 135.130 ;
        RECT 57.430 134.490 57.685 134.960 ;
        RECT 57.865 134.670 58.150 135.470 ;
        RECT 58.330 134.750 58.660 135.260 ;
        RECT 46.015 133.090 46.575 133.380 ;
        RECT 46.745 132.920 46.995 133.380 ;
        RECT 47.615 133.190 47.945 133.550 ;
        RECT 48.315 132.920 49.985 133.690 ;
        RECT 53.580 133.465 53.920 134.295 ;
        RECT 50.160 132.920 55.505 133.465 ;
        RECT 55.735 132.920 55.945 133.740 ;
        RECT 56.115 133.720 56.365 134.320 ;
        RECT 56.535 133.910 56.865 134.160 ;
        RECT 56.115 133.090 56.445 133.720 ;
        RECT 56.615 132.920 56.845 133.740 ;
        RECT 57.430 133.630 57.610 134.490 ;
        RECT 58.330 134.160 58.580 134.750 ;
        RECT 58.930 134.600 59.100 135.210 ;
        RECT 59.270 134.780 59.600 135.470 ;
        RECT 59.830 134.920 60.070 135.210 ;
        RECT 60.270 135.090 60.690 135.470 ;
        RECT 60.870 135.000 61.500 135.250 ;
        RECT 61.970 135.090 62.300 135.470 ;
        RECT 60.870 134.920 61.040 135.000 ;
        RECT 62.470 134.920 62.640 135.210 ;
        RECT 62.820 135.090 63.200 135.470 ;
        RECT 63.440 135.085 64.270 135.255 ;
        RECT 59.830 134.750 61.040 134.920 ;
        RECT 57.780 133.830 58.580 134.160 ;
        RECT 57.430 133.100 57.685 133.630 ;
        RECT 57.865 132.920 58.150 133.380 ;
        RECT 58.330 133.180 58.580 133.830 ;
        RECT 58.780 134.580 59.100 134.600 ;
        RECT 58.780 134.410 60.700 134.580 ;
        RECT 58.780 133.515 58.970 134.410 ;
        RECT 60.870 134.240 61.040 134.750 ;
        RECT 61.210 134.490 61.730 134.800 ;
        RECT 59.140 134.070 61.040 134.240 ;
        RECT 59.140 134.010 59.470 134.070 ;
        RECT 59.620 133.840 59.950 133.900 ;
        RECT 59.290 133.570 59.950 133.840 ;
        RECT 58.780 133.185 59.100 133.515 ;
        RECT 59.280 132.920 59.940 133.400 ;
        RECT 60.140 133.310 60.310 134.070 ;
        RECT 61.210 133.900 61.390 134.310 ;
        RECT 60.480 133.730 60.810 133.850 ;
        RECT 61.560 133.730 61.730 134.490 ;
        RECT 60.480 133.560 61.730 133.730 ;
        RECT 61.900 134.670 63.270 134.920 ;
        RECT 61.900 133.900 62.090 134.670 ;
        RECT 63.020 134.410 63.270 134.670 ;
        RECT 62.260 134.240 62.510 134.400 ;
        RECT 63.440 134.240 63.610 135.085 ;
        RECT 64.505 134.800 64.675 135.300 ;
        RECT 64.845 134.970 65.175 135.470 ;
        RECT 63.780 134.410 64.280 134.790 ;
        RECT 64.505 134.630 65.200 134.800 ;
        RECT 62.260 134.070 63.610 134.240 ;
        RECT 63.190 134.030 63.610 134.070 ;
        RECT 61.900 133.560 62.320 133.900 ;
        RECT 62.610 133.570 63.020 133.900 ;
        RECT 60.140 133.140 60.990 133.310 ;
        RECT 61.550 132.920 61.870 133.380 ;
        RECT 62.070 133.130 62.320 133.560 ;
        RECT 62.610 132.920 63.020 133.360 ;
        RECT 63.190 133.300 63.360 134.030 ;
        RECT 63.530 133.480 63.880 133.850 ;
        RECT 64.060 133.540 64.280 134.410 ;
        RECT 64.450 133.840 64.860 134.460 ;
        RECT 65.030 133.660 65.200 134.630 ;
        RECT 64.505 133.470 65.200 133.660 ;
        RECT 63.190 133.100 64.205 133.300 ;
        RECT 64.505 133.140 64.675 133.470 ;
        RECT 64.845 132.920 65.175 133.300 ;
        RECT 65.390 133.180 65.615 135.300 ;
        RECT 65.785 134.970 66.115 135.470 ;
        RECT 66.285 134.800 66.455 135.300 ;
        RECT 65.790 134.630 66.455 134.800 ;
        RECT 65.790 133.640 66.020 134.630 ;
        RECT 66.190 133.810 66.540 134.460 ;
        RECT 66.715 134.305 67.005 135.470 ;
        RECT 67.175 134.500 67.445 135.270 ;
        RECT 67.615 134.690 67.945 135.470 ;
        RECT 68.150 134.865 68.335 135.270 ;
        RECT 68.505 135.045 68.840 135.470 ;
        RECT 68.150 134.690 68.815 134.865 ;
        RECT 67.175 134.330 68.305 134.500 ;
        RECT 65.790 133.470 66.455 133.640 ;
        RECT 65.785 132.920 66.115 133.300 ;
        RECT 66.285 133.180 66.455 133.470 ;
        RECT 66.715 132.920 67.005 133.645 ;
        RECT 67.175 133.420 67.345 134.330 ;
        RECT 67.515 133.580 67.875 134.160 ;
        RECT 68.055 133.830 68.305 134.330 ;
        RECT 68.475 133.660 68.815 134.690 ;
        RECT 69.015 134.380 70.685 135.470 ;
        RECT 70.855 134.750 71.315 135.300 ;
        RECT 71.505 134.750 71.835 135.470 ;
        RECT 69.015 133.860 69.765 134.380 ;
        RECT 69.935 133.690 70.685 134.210 ;
        RECT 68.130 133.490 68.815 133.660 ;
        RECT 67.175 133.090 67.435 133.420 ;
        RECT 67.645 132.920 67.920 133.400 ;
        RECT 68.130 133.090 68.335 133.490 ;
        RECT 68.505 132.920 68.840 133.320 ;
        RECT 69.015 132.920 70.685 133.690 ;
        RECT 70.855 133.380 71.105 134.750 ;
        RECT 72.035 134.580 72.335 135.130 ;
        RECT 72.505 134.800 72.785 135.470 ;
        RECT 71.395 134.410 72.335 134.580 ;
        RECT 73.155 134.750 73.615 135.300 ;
        RECT 73.805 134.750 74.135 135.470 ;
        RECT 71.395 134.160 71.565 134.410 ;
        RECT 72.705 134.160 72.970 134.520 ;
        RECT 71.275 133.830 71.565 134.160 ;
        RECT 71.735 133.910 72.075 134.160 ;
        RECT 72.295 133.910 72.970 134.160 ;
        RECT 71.395 133.740 71.565 133.830 ;
        RECT 71.395 133.550 72.785 133.740 ;
        RECT 70.855 133.090 71.415 133.380 ;
        RECT 71.585 132.920 71.835 133.380 ;
        RECT 72.455 133.190 72.785 133.550 ;
        RECT 73.155 133.380 73.405 134.750 ;
        RECT 74.335 134.580 74.635 135.130 ;
        RECT 74.805 134.800 75.085 135.470 ;
        RECT 73.695 134.410 74.635 134.580 ;
        RECT 75.455 134.710 75.970 135.120 ;
        RECT 76.205 134.710 76.375 135.470 ;
        RECT 76.545 135.130 78.575 135.300 ;
        RECT 73.695 134.160 73.865 134.410 ;
        RECT 75.005 134.160 75.270 134.520 ;
        RECT 73.575 133.830 73.865 134.160 ;
        RECT 74.035 133.910 74.375 134.160 ;
        RECT 74.595 133.910 75.270 134.160 ;
        RECT 73.695 133.740 73.865 133.830 ;
        RECT 75.455 133.900 75.795 134.710 ;
        RECT 76.545 134.465 76.715 135.130 ;
        RECT 77.110 134.790 78.235 134.960 ;
        RECT 75.965 134.275 76.715 134.465 ;
        RECT 76.885 134.450 77.895 134.620 ;
        RECT 73.695 133.550 75.085 133.740 ;
        RECT 75.455 133.730 76.685 133.900 ;
        RECT 73.155 133.090 73.715 133.380 ;
        RECT 73.885 132.920 74.135 133.380 ;
        RECT 74.755 133.190 75.085 133.550 ;
        RECT 75.730 133.125 75.975 133.730 ;
        RECT 76.195 132.920 76.705 133.455 ;
        RECT 76.885 133.090 77.075 134.450 ;
        RECT 77.245 134.110 77.520 134.250 ;
        RECT 77.245 133.940 77.525 134.110 ;
        RECT 77.245 133.090 77.520 133.940 ;
        RECT 77.725 133.650 77.895 134.450 ;
        RECT 78.065 133.660 78.235 134.790 ;
        RECT 78.405 134.160 78.575 135.130 ;
        RECT 78.745 134.330 78.915 135.470 ;
        RECT 79.085 134.330 79.420 135.300 ;
        RECT 78.405 133.830 78.600 134.160 ;
        RECT 78.825 133.830 79.080 134.160 ;
        RECT 78.825 133.660 78.995 133.830 ;
        RECT 79.250 133.660 79.420 134.330 ;
        RECT 79.970 134.490 80.225 135.160 ;
        RECT 80.405 134.670 80.690 135.470 ;
        RECT 80.870 134.750 81.200 135.260 ;
        RECT 79.970 134.110 80.150 134.490 ;
        RECT 80.870 134.160 81.120 134.750 ;
        RECT 81.470 134.600 81.640 135.210 ;
        RECT 81.810 134.780 82.140 135.470 ;
        RECT 82.370 134.920 82.610 135.210 ;
        RECT 82.810 135.090 83.230 135.470 ;
        RECT 83.410 135.000 84.040 135.250 ;
        RECT 84.510 135.090 84.840 135.470 ;
        RECT 83.410 134.920 83.580 135.000 ;
        RECT 85.010 134.920 85.180 135.210 ;
        RECT 85.360 135.090 85.740 135.470 ;
        RECT 85.980 135.085 86.810 135.255 ;
        RECT 82.370 134.750 83.580 134.920 ;
        RECT 79.885 133.940 80.150 134.110 ;
        RECT 78.065 133.490 78.995 133.660 ;
        RECT 78.065 133.455 78.240 133.490 ;
        RECT 77.710 133.090 78.240 133.455 ;
        RECT 78.665 132.920 78.995 133.320 ;
        RECT 79.165 133.090 79.420 133.660 ;
        RECT 79.970 133.630 80.150 133.940 ;
        RECT 80.320 133.830 81.120 134.160 ;
        RECT 79.970 133.100 80.225 133.630 ;
        RECT 80.405 132.920 80.690 133.380 ;
        RECT 80.870 133.180 81.120 133.830 ;
        RECT 81.320 134.580 81.640 134.600 ;
        RECT 81.320 134.410 83.240 134.580 ;
        RECT 81.320 133.515 81.510 134.410 ;
        RECT 83.410 134.240 83.580 134.750 ;
        RECT 83.750 134.490 84.270 134.800 ;
        RECT 81.680 134.070 83.580 134.240 ;
        RECT 81.680 134.010 82.010 134.070 ;
        RECT 82.160 133.840 82.490 133.900 ;
        RECT 81.830 133.570 82.490 133.840 ;
        RECT 81.320 133.185 81.640 133.515 ;
        RECT 81.820 132.920 82.480 133.400 ;
        RECT 82.680 133.310 82.850 134.070 ;
        RECT 83.750 133.900 83.930 134.310 ;
        RECT 83.020 133.730 83.350 133.850 ;
        RECT 84.100 133.730 84.270 134.490 ;
        RECT 83.020 133.560 84.270 133.730 ;
        RECT 84.440 134.670 85.810 134.920 ;
        RECT 84.440 133.900 84.630 134.670 ;
        RECT 85.560 134.410 85.810 134.670 ;
        RECT 84.800 134.240 85.050 134.400 ;
        RECT 85.980 134.240 86.150 135.085 ;
        RECT 87.045 134.800 87.215 135.300 ;
        RECT 87.385 134.970 87.715 135.470 ;
        RECT 86.320 134.410 86.820 134.790 ;
        RECT 87.045 134.630 87.740 134.800 ;
        RECT 84.800 134.070 86.150 134.240 ;
        RECT 85.730 134.030 86.150 134.070 ;
        RECT 84.440 133.560 84.860 133.900 ;
        RECT 85.150 133.570 85.560 133.900 ;
        RECT 82.680 133.140 83.530 133.310 ;
        RECT 84.090 132.920 84.410 133.380 ;
        RECT 84.610 133.130 84.860 133.560 ;
        RECT 85.150 132.920 85.560 133.360 ;
        RECT 85.730 133.300 85.900 134.030 ;
        RECT 86.070 133.480 86.420 133.850 ;
        RECT 86.600 133.540 86.820 134.410 ;
        RECT 86.990 133.840 87.400 134.460 ;
        RECT 87.570 133.660 87.740 134.630 ;
        RECT 87.045 133.470 87.740 133.660 ;
        RECT 85.730 133.100 86.745 133.300 ;
        RECT 87.045 133.140 87.215 133.470 ;
        RECT 87.385 132.920 87.715 133.300 ;
        RECT 87.930 133.180 88.155 135.300 ;
        RECT 88.325 134.970 88.655 135.470 ;
        RECT 88.825 134.800 88.995 135.300 ;
        RECT 88.330 134.630 88.995 134.800 ;
        RECT 88.330 133.640 88.560 134.630 ;
        RECT 88.730 133.810 89.080 134.460 ;
        RECT 89.255 134.380 90.925 135.470 ;
        RECT 89.255 133.860 90.005 134.380 ;
        RECT 91.135 134.330 91.365 135.470 ;
        RECT 91.535 134.320 91.865 135.300 ;
        RECT 92.035 134.330 92.245 135.470 ;
        RECT 90.175 133.690 90.925 134.210 ;
        RECT 91.115 133.910 91.445 134.160 ;
        RECT 88.330 133.470 88.995 133.640 ;
        RECT 88.325 132.920 88.655 133.300 ;
        RECT 88.825 133.180 88.995 133.470 ;
        RECT 89.255 132.920 90.925 133.690 ;
        RECT 91.135 132.920 91.365 133.740 ;
        RECT 91.615 133.720 91.865 134.320 ;
        RECT 92.475 134.305 92.765 135.470 ;
        RECT 93.025 134.800 93.195 135.300 ;
        RECT 93.365 134.970 93.695 135.470 ;
        RECT 93.025 134.630 93.690 134.800 ;
        RECT 92.940 133.810 93.290 134.460 ;
        RECT 91.535 133.090 91.865 133.720 ;
        RECT 92.035 132.920 92.245 133.740 ;
        RECT 92.475 132.920 92.765 133.645 ;
        RECT 93.460 133.640 93.690 134.630 ;
        RECT 93.025 133.470 93.690 133.640 ;
        RECT 93.025 133.180 93.195 133.470 ;
        RECT 93.365 132.920 93.695 133.300 ;
        RECT 93.865 133.180 94.090 135.300 ;
        RECT 94.305 134.970 94.635 135.470 ;
        RECT 94.805 134.800 94.975 135.300 ;
        RECT 95.210 135.085 96.040 135.255 ;
        RECT 96.280 135.090 96.660 135.470 ;
        RECT 94.280 134.630 94.975 134.800 ;
        RECT 94.280 133.660 94.450 134.630 ;
        RECT 94.620 133.840 95.030 134.460 ;
        RECT 95.200 134.410 95.700 134.790 ;
        RECT 94.280 133.470 94.975 133.660 ;
        RECT 95.200 133.540 95.420 134.410 ;
        RECT 95.870 134.240 96.040 135.085 ;
        RECT 96.840 134.920 97.010 135.210 ;
        RECT 97.180 135.090 97.510 135.470 ;
        RECT 97.980 135.000 98.610 135.250 ;
        RECT 98.790 135.090 99.210 135.470 ;
        RECT 98.440 134.920 98.610 135.000 ;
        RECT 99.410 134.920 99.650 135.210 ;
        RECT 96.210 134.670 97.580 134.920 ;
        RECT 96.210 134.410 96.460 134.670 ;
        RECT 96.970 134.240 97.220 134.400 ;
        RECT 95.870 134.070 97.220 134.240 ;
        RECT 95.870 134.030 96.290 134.070 ;
        RECT 95.600 133.480 95.950 133.850 ;
        RECT 94.305 132.920 94.635 133.300 ;
        RECT 94.805 133.140 94.975 133.470 ;
        RECT 96.120 133.300 96.290 134.030 ;
        RECT 97.390 133.900 97.580 134.670 ;
        RECT 96.460 133.570 96.870 133.900 ;
        RECT 97.160 133.560 97.580 133.900 ;
        RECT 97.750 134.490 98.270 134.800 ;
        RECT 98.440 134.750 99.650 134.920 ;
        RECT 99.880 134.780 100.210 135.470 ;
        RECT 97.750 133.730 97.920 134.490 ;
        RECT 98.090 133.900 98.270 134.310 ;
        RECT 98.440 134.240 98.610 134.750 ;
        RECT 100.380 134.600 100.550 135.210 ;
        RECT 100.820 134.750 101.150 135.260 ;
        RECT 100.380 134.580 100.700 134.600 ;
        RECT 98.780 134.410 100.700 134.580 ;
        RECT 98.440 134.070 100.340 134.240 ;
        RECT 98.670 133.730 99.000 133.850 ;
        RECT 97.750 133.560 99.000 133.730 ;
        RECT 95.275 133.100 96.290 133.300 ;
        RECT 96.460 132.920 96.870 133.360 ;
        RECT 97.160 133.130 97.410 133.560 ;
        RECT 97.610 132.920 97.930 133.380 ;
        RECT 99.170 133.310 99.340 134.070 ;
        RECT 100.010 134.010 100.340 134.070 ;
        RECT 99.530 133.840 99.860 133.900 ;
        RECT 99.530 133.570 100.190 133.840 ;
        RECT 100.510 133.515 100.700 134.410 ;
        RECT 98.490 133.140 99.340 133.310 ;
        RECT 99.540 132.920 100.200 133.400 ;
        RECT 100.380 133.185 100.700 133.515 ;
        RECT 100.900 134.160 101.150 134.750 ;
        RECT 101.330 134.670 101.615 135.470 ;
        RECT 101.795 134.490 102.050 135.160 ;
        RECT 100.900 133.830 101.700 134.160 ;
        RECT 101.870 134.110 102.050 134.490 ;
        RECT 102.595 134.380 104.265 135.470 ;
        RECT 104.435 134.710 104.950 135.120 ;
        RECT 105.185 134.710 105.355 135.470 ;
        RECT 105.525 135.130 107.555 135.300 ;
        RECT 101.870 133.940 102.135 134.110 ;
        RECT 100.900 133.180 101.150 133.830 ;
        RECT 101.870 133.630 102.050 133.940 ;
        RECT 102.595 133.860 103.345 134.380 ;
        RECT 103.515 133.690 104.265 134.210 ;
        RECT 104.435 133.900 104.775 134.710 ;
        RECT 105.525 134.465 105.695 135.130 ;
        RECT 106.090 134.790 107.215 134.960 ;
        RECT 104.945 134.275 105.695 134.465 ;
        RECT 105.865 134.450 106.875 134.620 ;
        RECT 104.435 133.730 105.665 133.900 ;
        RECT 101.330 132.920 101.615 133.380 ;
        RECT 101.795 133.100 102.050 133.630 ;
        RECT 102.595 132.920 104.265 133.690 ;
        RECT 104.710 133.125 104.955 133.730 ;
        RECT 105.175 132.920 105.685 133.455 ;
        RECT 105.865 133.090 106.055 134.450 ;
        RECT 106.225 134.110 106.500 134.250 ;
        RECT 106.225 133.940 106.505 134.110 ;
        RECT 106.225 133.090 106.500 133.940 ;
        RECT 106.705 133.650 106.875 134.450 ;
        RECT 107.045 133.660 107.215 134.790 ;
        RECT 107.385 134.160 107.555 135.130 ;
        RECT 107.725 134.330 107.895 135.470 ;
        RECT 108.065 134.330 108.400 135.300 ;
        RECT 107.385 133.830 107.580 134.160 ;
        RECT 107.805 133.830 108.060 134.160 ;
        RECT 107.805 133.660 107.975 133.830 ;
        RECT 108.230 133.660 108.400 134.330 ;
        RECT 108.575 134.710 109.090 135.120 ;
        RECT 109.325 134.710 109.495 135.470 ;
        RECT 109.665 135.130 111.695 135.300 ;
        RECT 108.575 133.900 108.915 134.710 ;
        RECT 109.665 134.465 109.835 135.130 ;
        RECT 110.230 134.790 111.355 134.960 ;
        RECT 109.085 134.275 109.835 134.465 ;
        RECT 110.005 134.450 111.015 134.620 ;
        RECT 108.575 133.730 109.805 133.900 ;
        RECT 107.045 133.490 107.975 133.660 ;
        RECT 107.045 133.455 107.220 133.490 ;
        RECT 106.690 133.090 107.220 133.455 ;
        RECT 107.645 132.920 107.975 133.320 ;
        RECT 108.145 133.090 108.400 133.660 ;
        RECT 108.850 133.125 109.095 133.730 ;
        RECT 109.315 132.920 109.825 133.455 ;
        RECT 110.005 133.090 110.195 134.450 ;
        RECT 110.365 133.430 110.640 134.250 ;
        RECT 110.845 133.650 111.015 134.450 ;
        RECT 111.185 133.660 111.355 134.790 ;
        RECT 111.525 134.160 111.695 135.130 ;
        RECT 111.865 134.330 112.035 135.470 ;
        RECT 112.205 134.330 112.540 135.300 ;
        RECT 111.525 133.830 111.720 134.160 ;
        RECT 111.945 133.830 112.200 134.160 ;
        RECT 111.945 133.660 112.115 133.830 ;
        RECT 112.370 133.660 112.540 134.330 ;
        RECT 113.635 134.380 117.145 135.470 ;
        RECT 117.315 134.380 118.525 135.470 ;
        RECT 113.635 133.860 115.325 134.380 ;
        RECT 115.495 133.690 117.145 134.210 ;
        RECT 117.315 133.840 117.835 134.380 ;
        RECT 111.185 133.490 112.115 133.660 ;
        RECT 111.185 133.455 111.360 133.490 ;
        RECT 110.365 133.260 110.645 133.430 ;
        RECT 110.365 133.090 110.640 133.260 ;
        RECT 110.830 133.090 111.360 133.455 ;
        RECT 111.785 132.920 112.115 133.320 ;
        RECT 112.285 133.090 112.540 133.660 ;
        RECT 113.635 132.920 117.145 133.690 ;
        RECT 118.005 133.670 118.525 134.210 ;
        RECT 117.315 132.920 118.525 133.670 ;
        RECT 11.430 132.750 118.610 132.920 ;
        RECT 11.515 132.000 12.725 132.750 ;
        RECT 12.895 132.000 14.105 132.750 ;
        RECT 11.515 131.460 12.035 132.000 ;
        RECT 12.205 131.290 12.725 131.830 ;
        RECT 11.515 130.200 12.725 131.290 ;
        RECT 12.895 131.290 13.415 131.830 ;
        RECT 13.585 131.460 14.105 132.000 ;
        RECT 14.550 131.940 14.795 132.545 ;
        RECT 15.015 132.215 15.525 132.750 ;
        RECT 14.275 131.770 15.505 131.940 ;
        RECT 12.895 130.200 14.105 131.290 ;
        RECT 14.275 130.960 14.615 131.770 ;
        RECT 14.785 131.205 15.535 131.395 ;
        RECT 14.275 130.550 14.790 130.960 ;
        RECT 15.025 130.200 15.195 130.960 ;
        RECT 15.365 130.540 15.535 131.205 ;
        RECT 15.705 131.220 15.895 132.580 ;
        RECT 16.065 131.730 16.340 132.580 ;
        RECT 16.530 132.215 17.060 132.580 ;
        RECT 17.485 132.350 17.815 132.750 ;
        RECT 16.885 132.180 17.060 132.215 ;
        RECT 16.065 131.560 16.345 131.730 ;
        RECT 16.065 131.420 16.340 131.560 ;
        RECT 16.545 131.220 16.715 132.020 ;
        RECT 15.705 131.050 16.715 131.220 ;
        RECT 16.885 132.010 17.815 132.180 ;
        RECT 17.985 132.010 18.240 132.580 ;
        RECT 16.885 130.880 17.055 132.010 ;
        RECT 17.645 131.840 17.815 132.010 ;
        RECT 15.930 130.710 17.055 130.880 ;
        RECT 17.225 131.510 17.420 131.840 ;
        RECT 17.645 131.510 17.900 131.840 ;
        RECT 17.225 130.540 17.395 131.510 ;
        RECT 18.070 131.340 18.240 132.010 ;
        RECT 15.365 130.370 17.395 130.540 ;
        RECT 17.565 130.200 17.735 131.340 ;
        RECT 17.905 130.370 18.240 131.340 ;
        RECT 18.420 132.010 18.675 132.580 ;
        RECT 18.845 132.350 19.175 132.750 ;
        RECT 19.600 132.215 20.130 132.580 ;
        RECT 20.320 132.410 20.595 132.580 ;
        RECT 20.315 132.240 20.595 132.410 ;
        RECT 19.600 132.180 19.775 132.215 ;
        RECT 18.845 132.010 19.775 132.180 ;
        RECT 18.420 131.340 18.590 132.010 ;
        RECT 18.845 131.840 19.015 132.010 ;
        RECT 18.760 131.510 19.015 131.840 ;
        RECT 19.240 131.510 19.435 131.840 ;
        RECT 18.420 130.370 18.755 131.340 ;
        RECT 18.925 130.200 19.095 131.340 ;
        RECT 19.265 130.540 19.435 131.510 ;
        RECT 19.605 130.880 19.775 132.010 ;
        RECT 19.945 131.220 20.115 132.020 ;
        RECT 20.320 131.420 20.595 132.240 ;
        RECT 20.765 131.220 20.955 132.580 ;
        RECT 21.135 132.215 21.645 132.750 ;
        RECT 21.865 131.940 22.110 132.545 ;
        RECT 23.015 131.980 26.525 132.750 ;
        RECT 21.155 131.770 22.385 131.940 ;
        RECT 19.945 131.050 20.955 131.220 ;
        RECT 21.125 131.205 21.875 131.395 ;
        RECT 19.605 130.710 20.730 130.880 ;
        RECT 21.125 130.540 21.295 131.205 ;
        RECT 22.045 130.960 22.385 131.770 ;
        RECT 19.265 130.370 21.295 130.540 ;
        RECT 21.465 130.200 21.635 130.960 ;
        RECT 21.870 130.550 22.385 130.960 ;
        RECT 23.015 131.290 24.705 131.810 ;
        RECT 24.875 131.460 26.525 131.980 ;
        RECT 26.735 131.930 26.965 132.750 ;
        RECT 27.135 131.950 27.465 132.580 ;
        RECT 26.715 131.510 27.045 131.760 ;
        RECT 27.215 131.350 27.465 131.950 ;
        RECT 27.635 131.930 27.845 132.750 ;
        RECT 28.075 132.025 28.365 132.750 ;
        RECT 28.910 132.410 29.165 132.570 ;
        RECT 28.825 132.240 29.165 132.410 ;
        RECT 29.345 132.290 29.630 132.750 ;
        RECT 28.910 132.040 29.165 132.240 ;
        RECT 23.015 130.200 26.525 131.290 ;
        RECT 26.735 130.200 26.965 131.340 ;
        RECT 27.135 130.370 27.465 131.350 ;
        RECT 27.635 130.200 27.845 131.340 ;
        RECT 28.075 130.200 28.365 131.365 ;
        RECT 28.910 131.180 29.090 132.040 ;
        RECT 29.810 131.840 30.060 132.490 ;
        RECT 29.260 131.510 30.060 131.840 ;
        RECT 28.910 130.510 29.165 131.180 ;
        RECT 29.345 130.200 29.630 131.000 ;
        RECT 29.810 130.920 30.060 131.510 ;
        RECT 30.260 132.155 30.580 132.485 ;
        RECT 30.760 132.270 31.420 132.750 ;
        RECT 31.620 132.360 32.470 132.530 ;
        RECT 30.260 131.260 30.450 132.155 ;
        RECT 30.770 131.830 31.430 132.100 ;
        RECT 31.100 131.770 31.430 131.830 ;
        RECT 30.620 131.600 30.950 131.660 ;
        RECT 31.620 131.600 31.790 132.360 ;
        RECT 33.030 132.290 33.350 132.750 ;
        RECT 33.550 132.110 33.800 132.540 ;
        RECT 34.090 132.310 34.500 132.750 ;
        RECT 34.670 132.370 35.685 132.570 ;
        RECT 31.960 131.940 33.210 132.110 ;
        RECT 31.960 131.820 32.290 131.940 ;
        RECT 30.620 131.430 32.520 131.600 ;
        RECT 30.260 131.090 32.180 131.260 ;
        RECT 30.260 131.070 30.580 131.090 ;
        RECT 29.810 130.410 30.140 130.920 ;
        RECT 30.410 130.460 30.580 131.070 ;
        RECT 32.350 130.920 32.520 131.430 ;
        RECT 32.690 131.360 32.870 131.770 ;
        RECT 33.040 131.180 33.210 131.940 ;
        RECT 30.750 130.200 31.080 130.890 ;
        RECT 31.310 130.750 32.520 130.920 ;
        RECT 32.690 130.870 33.210 131.180 ;
        RECT 33.380 131.770 33.800 132.110 ;
        RECT 34.090 131.770 34.500 132.100 ;
        RECT 33.380 131.000 33.570 131.770 ;
        RECT 34.670 131.640 34.840 132.370 ;
        RECT 35.985 132.200 36.155 132.530 ;
        RECT 36.325 132.370 36.655 132.750 ;
        RECT 35.010 131.820 35.360 132.190 ;
        RECT 34.670 131.600 35.090 131.640 ;
        RECT 33.740 131.430 35.090 131.600 ;
        RECT 33.740 131.270 33.990 131.430 ;
        RECT 34.500 131.000 34.750 131.260 ;
        RECT 33.380 130.750 34.750 131.000 ;
        RECT 31.310 130.460 31.550 130.750 ;
        RECT 32.350 130.670 32.520 130.750 ;
        RECT 31.750 130.200 32.170 130.580 ;
        RECT 32.350 130.420 32.980 130.670 ;
        RECT 33.450 130.200 33.780 130.580 ;
        RECT 33.950 130.460 34.120 130.750 ;
        RECT 34.920 130.585 35.090 131.430 ;
        RECT 35.540 131.260 35.760 132.130 ;
        RECT 35.985 132.010 36.680 132.200 ;
        RECT 35.260 130.880 35.760 131.260 ;
        RECT 35.930 131.210 36.340 131.830 ;
        RECT 36.510 131.040 36.680 132.010 ;
        RECT 35.985 130.870 36.680 131.040 ;
        RECT 34.300 130.200 34.680 130.580 ;
        RECT 34.920 130.415 35.750 130.585 ;
        RECT 35.985 130.370 36.155 130.870 ;
        RECT 36.325 130.200 36.655 130.700 ;
        RECT 36.870 130.370 37.095 132.490 ;
        RECT 37.265 132.370 37.595 132.750 ;
        RECT 37.765 132.200 37.935 132.490 ;
        RECT 37.270 132.030 37.935 132.200 ;
        RECT 38.195 132.075 38.455 132.580 ;
        RECT 38.635 132.370 38.965 132.750 ;
        RECT 39.145 132.200 39.315 132.580 ;
        RECT 37.270 131.040 37.500 132.030 ;
        RECT 37.670 131.210 38.020 131.860 ;
        RECT 38.195 131.275 38.365 132.075 ;
        RECT 38.650 132.030 39.315 132.200 ;
        RECT 38.650 131.775 38.820 132.030 ;
        RECT 40.035 131.980 42.625 132.750 ;
        RECT 42.800 132.205 48.145 132.750 ;
        RECT 48.315 132.290 48.875 132.580 ;
        RECT 49.045 132.290 49.295 132.750 ;
        RECT 38.535 131.445 38.820 131.775 ;
        RECT 39.055 131.480 39.385 131.850 ;
        RECT 38.650 131.300 38.820 131.445 ;
        RECT 37.270 130.870 37.935 131.040 ;
        RECT 37.265 130.200 37.595 130.700 ;
        RECT 37.765 130.370 37.935 130.870 ;
        RECT 38.195 130.370 38.465 131.275 ;
        RECT 38.650 131.130 39.315 131.300 ;
        RECT 38.635 130.200 38.965 130.960 ;
        RECT 39.145 130.370 39.315 131.130 ;
        RECT 40.035 131.290 41.245 131.810 ;
        RECT 41.415 131.460 42.625 131.980 ;
        RECT 40.035 130.200 42.625 131.290 ;
        RECT 44.390 130.635 44.740 131.885 ;
        RECT 46.220 131.375 46.560 132.205 ;
        RECT 48.315 130.920 48.565 132.290 ;
        RECT 49.915 132.120 50.245 132.480 ;
        RECT 48.855 131.930 50.245 132.120 ;
        RECT 51.075 131.980 53.665 132.750 ;
        RECT 53.835 132.025 54.125 132.750 ;
        RECT 54.755 131.980 56.425 132.750 ;
        RECT 56.655 132.270 56.935 132.750 ;
        RECT 57.105 132.100 57.365 132.490 ;
        RECT 57.540 132.270 57.795 132.750 ;
        RECT 57.965 132.100 58.260 132.490 ;
        RECT 58.440 132.270 58.715 132.750 ;
        RECT 58.885 132.250 59.185 132.580 ;
        RECT 48.855 131.840 49.025 131.930 ;
        RECT 48.735 131.510 49.025 131.840 ;
        RECT 49.195 131.510 49.535 131.760 ;
        RECT 49.755 131.510 50.430 131.760 ;
        RECT 48.855 131.260 49.025 131.510 ;
        RECT 48.855 131.090 49.795 131.260 ;
        RECT 50.165 131.150 50.430 131.510 ;
        RECT 51.075 131.290 52.285 131.810 ;
        RECT 52.455 131.460 53.665 131.980 ;
        RECT 42.800 130.200 48.145 130.635 ;
        RECT 48.315 130.370 48.775 130.920 ;
        RECT 48.965 130.200 49.295 130.920 ;
        RECT 49.495 130.540 49.795 131.090 ;
        RECT 49.965 130.200 50.245 130.870 ;
        RECT 51.075 130.200 53.665 131.290 ;
        RECT 53.835 130.200 54.125 131.365 ;
        RECT 54.755 131.290 55.505 131.810 ;
        RECT 55.675 131.460 56.425 131.980 ;
        RECT 56.610 131.930 58.260 132.100 ;
        RECT 56.610 131.420 57.015 131.930 ;
        RECT 57.185 131.590 58.325 131.760 ;
        RECT 54.755 130.200 56.425 131.290 ;
        RECT 56.610 131.250 57.365 131.420 ;
        RECT 56.650 130.200 56.935 131.070 ;
        RECT 57.105 131.000 57.365 131.250 ;
        RECT 58.155 131.340 58.325 131.590 ;
        RECT 58.495 131.510 58.845 132.080 ;
        RECT 59.015 131.340 59.185 132.250 ;
        RECT 59.630 131.940 59.875 132.545 ;
        RECT 60.095 132.215 60.605 132.750 ;
        RECT 58.155 131.170 59.185 131.340 ;
        RECT 57.105 130.830 58.225 131.000 ;
        RECT 57.105 130.370 57.365 130.830 ;
        RECT 57.540 130.200 57.795 130.660 ;
        RECT 57.965 130.370 58.225 130.830 ;
        RECT 58.395 130.200 58.705 131.000 ;
        RECT 58.875 130.370 59.185 131.170 ;
        RECT 59.355 131.770 60.585 131.940 ;
        RECT 59.355 130.960 59.695 131.770 ;
        RECT 59.865 131.205 60.615 131.395 ;
        RECT 59.355 130.550 59.870 130.960 ;
        RECT 60.105 130.200 60.275 130.960 ;
        RECT 60.445 130.540 60.615 131.205 ;
        RECT 60.785 131.220 60.975 132.580 ;
        RECT 61.145 132.410 61.420 132.580 ;
        RECT 61.145 132.240 61.425 132.410 ;
        RECT 61.145 131.420 61.420 132.240 ;
        RECT 61.610 132.215 62.140 132.580 ;
        RECT 62.565 132.350 62.895 132.750 ;
        RECT 61.965 132.180 62.140 132.215 ;
        RECT 61.625 131.220 61.795 132.020 ;
        RECT 60.785 131.050 61.795 131.220 ;
        RECT 61.965 132.010 62.895 132.180 ;
        RECT 63.065 132.010 63.320 132.580 ;
        RECT 64.505 132.200 64.675 132.580 ;
        RECT 64.855 132.370 65.185 132.750 ;
        RECT 64.505 132.030 65.170 132.200 ;
        RECT 65.365 132.075 65.625 132.580 ;
        RECT 61.965 130.880 62.135 132.010 ;
        RECT 62.725 131.840 62.895 132.010 ;
        RECT 61.010 130.710 62.135 130.880 ;
        RECT 62.305 131.510 62.500 131.840 ;
        RECT 62.725 131.510 62.980 131.840 ;
        RECT 62.305 130.540 62.475 131.510 ;
        RECT 63.150 131.340 63.320 132.010 ;
        RECT 64.435 131.480 64.765 131.850 ;
        RECT 65.000 131.775 65.170 132.030 ;
        RECT 60.445 130.370 62.475 130.540 ;
        RECT 62.645 130.200 62.815 131.340 ;
        RECT 62.985 130.370 63.320 131.340 ;
        RECT 65.000 131.445 65.285 131.775 ;
        RECT 65.000 131.300 65.170 131.445 ;
        RECT 64.505 131.130 65.170 131.300 ;
        RECT 65.455 131.275 65.625 132.075 ;
        RECT 65.995 132.120 66.325 132.480 ;
        RECT 66.945 132.290 67.195 132.750 ;
        RECT 67.365 132.290 67.925 132.580 ;
        RECT 65.995 131.930 67.385 132.120 ;
        RECT 67.215 131.840 67.385 131.930 ;
        RECT 64.505 130.370 64.675 131.130 ;
        RECT 64.855 130.200 65.185 130.960 ;
        RECT 65.355 130.370 65.625 131.275 ;
        RECT 65.810 131.510 66.485 131.760 ;
        RECT 66.705 131.510 67.045 131.760 ;
        RECT 67.215 131.510 67.505 131.840 ;
        RECT 65.810 131.150 66.075 131.510 ;
        RECT 67.215 131.260 67.385 131.510 ;
        RECT 66.445 131.090 67.385 131.260 ;
        RECT 65.995 130.200 66.275 130.870 ;
        RECT 66.445 130.540 66.745 131.090 ;
        RECT 67.675 130.920 67.925 132.290 ;
        RECT 66.945 130.200 67.275 130.920 ;
        RECT 67.465 130.370 67.925 130.920 ;
        RECT 68.555 132.250 68.855 132.580 ;
        RECT 69.025 132.270 69.300 132.750 ;
        RECT 68.555 131.340 68.725 132.250 ;
        RECT 69.480 132.100 69.775 132.490 ;
        RECT 69.945 132.270 70.200 132.750 ;
        RECT 70.375 132.100 70.635 132.490 ;
        RECT 70.805 132.270 71.085 132.750 ;
        RECT 68.895 131.510 69.245 132.080 ;
        RECT 69.480 131.930 71.130 132.100 ;
        RECT 71.775 131.980 73.445 132.750 ;
        RECT 69.415 131.590 70.555 131.760 ;
        RECT 69.415 131.340 69.585 131.590 ;
        RECT 70.725 131.420 71.130 131.930 ;
        RECT 68.555 131.170 69.585 131.340 ;
        RECT 70.375 131.250 71.130 131.420 ;
        RECT 71.775 131.290 72.525 131.810 ;
        RECT 72.695 131.460 73.445 131.980 ;
        RECT 73.890 131.940 74.135 132.545 ;
        RECT 74.355 132.215 74.865 132.750 ;
        RECT 73.615 131.770 74.845 131.940 ;
        RECT 68.555 130.370 68.865 131.170 ;
        RECT 70.375 131.000 70.635 131.250 ;
        RECT 69.035 130.200 69.345 131.000 ;
        RECT 69.515 130.830 70.635 131.000 ;
        RECT 69.515 130.370 69.775 130.830 ;
        RECT 69.945 130.200 70.200 130.660 ;
        RECT 70.375 130.370 70.635 130.830 ;
        RECT 70.805 130.200 71.090 131.070 ;
        RECT 71.775 130.200 73.445 131.290 ;
        RECT 73.615 130.960 73.955 131.770 ;
        RECT 74.125 131.205 74.875 131.395 ;
        RECT 73.615 130.550 74.130 130.960 ;
        RECT 74.365 130.200 74.535 130.960 ;
        RECT 74.705 130.540 74.875 131.205 ;
        RECT 75.045 131.220 75.235 132.580 ;
        RECT 75.405 131.730 75.680 132.580 ;
        RECT 75.870 132.215 76.400 132.580 ;
        RECT 76.825 132.350 77.155 132.750 ;
        RECT 76.225 132.180 76.400 132.215 ;
        RECT 75.405 131.560 75.685 131.730 ;
        RECT 75.405 131.420 75.680 131.560 ;
        RECT 75.885 131.220 76.055 132.020 ;
        RECT 75.045 131.050 76.055 131.220 ;
        RECT 76.225 132.010 77.155 132.180 ;
        RECT 77.325 132.010 77.580 132.580 ;
        RECT 76.225 130.880 76.395 132.010 ;
        RECT 76.985 131.840 77.155 132.010 ;
        RECT 75.270 130.710 76.395 130.880 ;
        RECT 76.565 131.510 76.760 131.840 ;
        RECT 76.985 131.510 77.240 131.840 ;
        RECT 76.565 130.540 76.735 131.510 ;
        RECT 77.410 131.340 77.580 132.010 ;
        RECT 77.755 131.980 79.425 132.750 ;
        RECT 79.595 132.025 79.885 132.750 ;
        RECT 80.055 132.075 80.315 132.580 ;
        RECT 80.495 132.370 80.825 132.750 ;
        RECT 81.005 132.200 81.175 132.580 ;
        RECT 74.705 130.370 76.735 130.540 ;
        RECT 76.905 130.200 77.075 131.340 ;
        RECT 77.245 130.370 77.580 131.340 ;
        RECT 77.755 131.290 78.505 131.810 ;
        RECT 78.675 131.460 79.425 131.980 ;
        RECT 77.755 130.200 79.425 131.290 ;
        RECT 79.595 130.200 79.885 131.365 ;
        RECT 80.055 131.275 80.225 132.075 ;
        RECT 80.510 132.030 81.175 132.200 ;
        RECT 80.510 131.775 80.680 132.030 ;
        RECT 81.435 131.980 84.025 132.750 ;
        RECT 84.285 132.200 84.455 132.580 ;
        RECT 84.635 132.370 84.965 132.750 ;
        RECT 84.285 132.030 84.950 132.200 ;
        RECT 85.145 132.075 85.405 132.580 ;
        RECT 85.580 132.205 90.925 132.750 ;
        RECT 91.095 132.290 91.655 132.580 ;
        RECT 91.825 132.290 92.075 132.750 ;
        RECT 80.395 131.445 80.680 131.775 ;
        RECT 80.915 131.480 81.245 131.850 ;
        RECT 80.510 131.300 80.680 131.445 ;
        RECT 80.055 130.370 80.325 131.275 ;
        RECT 80.510 131.130 81.175 131.300 ;
        RECT 80.495 130.200 80.825 130.960 ;
        RECT 81.005 130.370 81.175 131.130 ;
        RECT 81.435 131.290 82.645 131.810 ;
        RECT 82.815 131.460 84.025 131.980 ;
        RECT 84.215 131.480 84.545 131.850 ;
        RECT 84.780 131.775 84.950 132.030 ;
        RECT 84.780 131.445 85.065 131.775 ;
        RECT 84.780 131.300 84.950 131.445 ;
        RECT 81.435 130.200 84.025 131.290 ;
        RECT 84.285 131.130 84.950 131.300 ;
        RECT 85.235 131.275 85.405 132.075 ;
        RECT 84.285 130.370 84.455 131.130 ;
        RECT 84.635 130.200 84.965 130.960 ;
        RECT 85.135 130.370 85.405 131.275 ;
        RECT 87.170 130.635 87.520 131.885 ;
        RECT 89.000 131.375 89.340 132.205 ;
        RECT 91.095 130.920 91.345 132.290 ;
        RECT 92.695 132.120 93.025 132.480 ;
        RECT 91.635 131.930 93.025 132.120 ;
        RECT 93.670 131.940 93.915 132.545 ;
        RECT 94.135 132.215 94.645 132.750 ;
        RECT 91.635 131.840 91.805 131.930 ;
        RECT 91.515 131.510 91.805 131.840 ;
        RECT 93.395 131.770 94.625 131.940 ;
        RECT 91.975 131.510 92.315 131.760 ;
        RECT 92.535 131.510 93.210 131.760 ;
        RECT 91.635 131.260 91.805 131.510 ;
        RECT 91.635 131.090 92.575 131.260 ;
        RECT 92.945 131.150 93.210 131.510 ;
        RECT 85.580 130.200 90.925 130.635 ;
        RECT 91.095 130.370 91.555 130.920 ;
        RECT 91.745 130.200 92.075 130.920 ;
        RECT 92.275 130.540 92.575 131.090 ;
        RECT 93.395 130.960 93.735 131.770 ;
        RECT 93.905 131.205 94.655 131.395 ;
        RECT 92.745 130.200 93.025 130.870 ;
        RECT 93.395 130.550 93.910 130.960 ;
        RECT 94.145 130.200 94.315 130.960 ;
        RECT 94.485 130.540 94.655 131.205 ;
        RECT 94.825 131.220 95.015 132.580 ;
        RECT 95.185 131.730 95.460 132.580 ;
        RECT 95.650 132.215 96.180 132.580 ;
        RECT 96.605 132.350 96.935 132.750 ;
        RECT 96.005 132.180 96.180 132.215 ;
        RECT 95.185 131.560 95.465 131.730 ;
        RECT 95.185 131.420 95.460 131.560 ;
        RECT 95.665 131.220 95.835 132.020 ;
        RECT 94.825 131.050 95.835 131.220 ;
        RECT 96.005 132.010 96.935 132.180 ;
        RECT 97.105 132.010 97.360 132.580 ;
        RECT 96.005 130.880 96.175 132.010 ;
        RECT 96.765 131.840 96.935 132.010 ;
        RECT 95.050 130.710 96.175 130.880 ;
        RECT 96.345 131.510 96.540 131.840 ;
        RECT 96.765 131.510 97.020 131.840 ;
        RECT 96.345 130.540 96.515 131.510 ;
        RECT 97.190 131.340 97.360 132.010 ;
        RECT 94.485 130.370 96.515 130.540 ;
        RECT 96.685 130.200 96.855 131.340 ;
        RECT 97.025 130.370 97.360 131.340 ;
        RECT 97.995 132.290 98.555 132.580 ;
        RECT 98.725 132.290 98.975 132.750 ;
        RECT 97.995 130.920 98.245 132.290 ;
        RECT 99.595 132.120 99.925 132.480 ;
        RECT 98.535 131.930 99.925 132.120 ;
        RECT 100.295 132.290 100.855 132.580 ;
        RECT 101.025 132.290 101.275 132.750 ;
        RECT 98.535 131.840 98.705 131.930 ;
        RECT 98.415 131.510 98.705 131.840 ;
        RECT 98.875 131.510 99.215 131.760 ;
        RECT 99.435 131.510 100.110 131.760 ;
        RECT 98.535 131.260 98.705 131.510 ;
        RECT 98.535 131.090 99.475 131.260 ;
        RECT 99.845 131.150 100.110 131.510 ;
        RECT 97.995 130.370 98.455 130.920 ;
        RECT 98.645 130.200 98.975 130.920 ;
        RECT 99.175 130.540 99.475 131.090 ;
        RECT 100.295 130.920 100.545 132.290 ;
        RECT 101.895 132.120 102.225 132.480 ;
        RECT 100.835 131.930 102.225 132.120 ;
        RECT 102.595 132.290 103.155 132.580 ;
        RECT 103.325 132.290 103.575 132.750 ;
        RECT 100.835 131.840 101.005 131.930 ;
        RECT 100.715 131.510 101.005 131.840 ;
        RECT 101.175 131.510 101.515 131.760 ;
        RECT 101.735 131.510 102.410 131.760 ;
        RECT 100.835 131.260 101.005 131.510 ;
        RECT 100.835 131.090 101.775 131.260 ;
        RECT 102.145 131.150 102.410 131.510 ;
        RECT 99.645 130.200 99.925 130.870 ;
        RECT 100.295 130.370 100.755 130.920 ;
        RECT 100.945 130.200 101.275 130.920 ;
        RECT 101.475 130.540 101.775 131.090 ;
        RECT 102.595 130.920 102.845 132.290 ;
        RECT 104.195 132.120 104.525 132.480 ;
        RECT 103.135 131.930 104.525 132.120 ;
        RECT 105.355 132.025 105.645 132.750 ;
        RECT 107.110 132.040 107.365 132.570 ;
        RECT 107.545 132.290 107.830 132.750 ;
        RECT 103.135 131.840 103.305 131.930 ;
        RECT 103.015 131.510 103.305 131.840 ;
        RECT 103.475 131.510 103.815 131.760 ;
        RECT 104.035 131.510 104.710 131.760 ;
        RECT 103.135 131.260 103.305 131.510 ;
        RECT 103.135 131.090 104.075 131.260 ;
        RECT 104.445 131.150 104.710 131.510 ;
        RECT 107.110 131.390 107.290 132.040 ;
        RECT 108.010 131.840 108.260 132.490 ;
        RECT 107.460 131.510 108.260 131.840 ;
        RECT 101.945 130.200 102.225 130.870 ;
        RECT 102.595 130.370 103.055 130.920 ;
        RECT 103.245 130.200 103.575 130.920 ;
        RECT 103.775 130.540 104.075 131.090 ;
        RECT 104.245 130.200 104.525 130.870 ;
        RECT 105.355 130.200 105.645 131.365 ;
        RECT 107.025 131.220 107.290 131.390 ;
        RECT 107.110 131.180 107.290 131.220 ;
        RECT 107.110 130.510 107.365 131.180 ;
        RECT 107.545 130.200 107.830 131.000 ;
        RECT 108.010 130.920 108.260 131.510 ;
        RECT 108.460 132.155 108.780 132.485 ;
        RECT 108.960 132.270 109.620 132.750 ;
        RECT 109.820 132.360 110.670 132.530 ;
        RECT 108.460 131.260 108.650 132.155 ;
        RECT 108.970 131.830 109.630 132.100 ;
        RECT 109.300 131.770 109.630 131.830 ;
        RECT 108.820 131.600 109.150 131.660 ;
        RECT 109.820 131.600 109.990 132.360 ;
        RECT 111.230 132.290 111.550 132.750 ;
        RECT 111.750 132.110 112.000 132.540 ;
        RECT 112.290 132.310 112.700 132.750 ;
        RECT 112.870 132.370 113.885 132.570 ;
        RECT 110.160 131.940 111.410 132.110 ;
        RECT 110.160 131.820 110.490 131.940 ;
        RECT 108.820 131.430 110.720 131.600 ;
        RECT 108.460 131.090 110.380 131.260 ;
        RECT 108.460 131.070 108.780 131.090 ;
        RECT 108.010 130.410 108.340 130.920 ;
        RECT 108.610 130.460 108.780 131.070 ;
        RECT 110.550 130.920 110.720 131.430 ;
        RECT 110.890 131.360 111.070 131.770 ;
        RECT 111.240 131.180 111.410 131.940 ;
        RECT 108.950 130.200 109.280 130.890 ;
        RECT 109.510 130.750 110.720 130.920 ;
        RECT 110.890 130.870 111.410 131.180 ;
        RECT 111.580 131.770 112.000 132.110 ;
        RECT 112.290 131.770 112.700 132.100 ;
        RECT 111.580 131.000 111.770 131.770 ;
        RECT 112.870 131.640 113.040 132.370 ;
        RECT 114.185 132.200 114.355 132.530 ;
        RECT 114.525 132.370 114.855 132.750 ;
        RECT 113.210 131.820 113.560 132.190 ;
        RECT 112.870 131.600 113.290 131.640 ;
        RECT 111.940 131.430 113.290 131.600 ;
        RECT 111.940 131.270 112.190 131.430 ;
        RECT 112.700 131.000 112.950 131.260 ;
        RECT 111.580 130.750 112.950 131.000 ;
        RECT 109.510 130.460 109.750 130.750 ;
        RECT 110.550 130.670 110.720 130.750 ;
        RECT 109.950 130.200 110.370 130.580 ;
        RECT 110.550 130.420 111.180 130.670 ;
        RECT 111.650 130.200 111.980 130.580 ;
        RECT 112.150 130.460 112.320 130.750 ;
        RECT 113.120 130.585 113.290 131.430 ;
        RECT 113.740 131.260 113.960 132.130 ;
        RECT 114.185 132.010 114.880 132.200 ;
        RECT 113.460 130.880 113.960 131.260 ;
        RECT 114.130 131.210 114.540 131.830 ;
        RECT 114.710 131.040 114.880 132.010 ;
        RECT 114.185 130.870 114.880 131.040 ;
        RECT 112.500 130.200 112.880 130.580 ;
        RECT 113.120 130.415 113.950 130.585 ;
        RECT 114.185 130.370 114.355 130.870 ;
        RECT 114.525 130.200 114.855 130.700 ;
        RECT 115.070 130.370 115.295 132.490 ;
        RECT 115.465 132.370 115.795 132.750 ;
        RECT 115.965 132.200 116.135 132.490 ;
        RECT 115.470 132.030 116.135 132.200 ;
        RECT 115.470 131.040 115.700 132.030 ;
        RECT 117.315 132.000 118.525 132.750 ;
        RECT 115.870 131.210 116.220 131.860 ;
        RECT 117.315 131.290 117.835 131.830 ;
        RECT 118.005 131.460 118.525 132.000 ;
        RECT 115.470 130.870 116.135 131.040 ;
        RECT 115.465 130.200 115.795 130.700 ;
        RECT 115.965 130.370 116.135 130.870 ;
        RECT 117.315 130.200 118.525 131.290 ;
        RECT 11.430 130.030 118.610 130.200 ;
        RECT 11.515 128.940 12.725 130.030 ;
        RECT 11.515 128.230 12.035 128.770 ;
        RECT 12.205 128.400 12.725 128.940 ;
        RECT 13.875 128.890 14.085 130.030 ;
        RECT 14.255 128.880 14.585 129.860 ;
        RECT 14.755 128.890 14.985 130.030 ;
        RECT 11.515 127.480 12.725 128.230 ;
        RECT 13.875 127.480 14.085 128.300 ;
        RECT 14.255 128.280 14.505 128.880 ;
        RECT 15.195 128.865 15.485 130.030 ;
        RECT 16.665 129.100 16.835 129.860 ;
        RECT 17.015 129.270 17.345 130.030 ;
        RECT 16.665 128.930 17.330 129.100 ;
        RECT 17.515 128.955 17.785 129.860 ;
        RECT 17.160 128.785 17.330 128.930 ;
        RECT 14.675 128.470 15.005 128.720 ;
        RECT 16.595 128.380 16.925 128.750 ;
        RECT 17.160 128.455 17.445 128.785 ;
        RECT 14.255 127.650 14.585 128.280 ;
        RECT 14.755 127.480 14.985 128.300 ;
        RECT 15.195 127.480 15.485 128.205 ;
        RECT 17.160 128.200 17.330 128.455 ;
        RECT 16.665 128.030 17.330 128.200 ;
        RECT 17.615 128.155 17.785 128.955 ;
        RECT 16.665 127.650 16.835 128.030 ;
        RECT 17.015 127.480 17.345 127.860 ;
        RECT 17.525 127.650 17.785 128.155 ;
        RECT 17.960 128.890 18.295 129.860 ;
        RECT 18.465 128.890 18.635 130.030 ;
        RECT 18.805 129.690 20.835 129.860 ;
        RECT 17.960 128.220 18.130 128.890 ;
        RECT 18.805 128.720 18.975 129.690 ;
        RECT 18.300 128.390 18.555 128.720 ;
        RECT 18.780 128.390 18.975 128.720 ;
        RECT 19.145 129.350 20.270 129.520 ;
        RECT 18.385 128.220 18.555 128.390 ;
        RECT 19.145 128.220 19.315 129.350 ;
        RECT 17.960 127.650 18.215 128.220 ;
        RECT 18.385 128.050 19.315 128.220 ;
        RECT 19.485 129.010 20.495 129.180 ;
        RECT 19.485 128.210 19.655 129.010 ;
        RECT 19.140 128.015 19.315 128.050 ;
        RECT 18.385 127.480 18.715 127.880 ;
        RECT 19.140 127.650 19.670 128.015 ;
        RECT 19.860 127.990 20.135 128.810 ;
        RECT 19.855 127.820 20.135 127.990 ;
        RECT 19.860 127.650 20.135 127.820 ;
        RECT 20.305 127.650 20.495 129.010 ;
        RECT 20.665 129.025 20.835 129.690 ;
        RECT 21.005 129.270 21.175 130.030 ;
        RECT 21.410 129.270 21.925 129.680 ;
        RECT 23.020 129.595 28.365 130.030 ;
        RECT 28.540 129.595 33.885 130.030 ;
        RECT 20.665 128.835 21.415 129.025 ;
        RECT 21.585 128.460 21.925 129.270 ;
        RECT 20.695 128.290 21.925 128.460 ;
        RECT 24.610 128.345 24.960 129.595 ;
        RECT 20.675 127.480 21.185 128.015 ;
        RECT 21.405 127.685 21.650 128.290 ;
        RECT 26.440 128.025 26.780 128.855 ;
        RECT 30.130 128.345 30.480 129.595 ;
        RECT 34.255 129.360 34.535 130.030 ;
        RECT 34.705 129.140 35.005 129.690 ;
        RECT 35.205 129.310 35.535 130.030 ;
        RECT 35.725 129.310 36.185 129.860 ;
        RECT 31.960 128.025 32.300 128.855 ;
        RECT 34.070 128.720 34.335 129.080 ;
        RECT 34.705 128.970 35.645 129.140 ;
        RECT 35.475 128.720 35.645 128.970 ;
        RECT 34.070 128.470 34.745 128.720 ;
        RECT 34.965 128.470 35.305 128.720 ;
        RECT 35.475 128.390 35.765 128.720 ;
        RECT 35.475 128.300 35.645 128.390 ;
        RECT 34.255 128.110 35.645 128.300 ;
        RECT 23.020 127.480 28.365 128.025 ;
        RECT 28.540 127.480 33.885 128.025 ;
        RECT 34.255 127.750 34.585 128.110 ;
        RECT 35.935 127.940 36.185 129.310 ;
        RECT 36.815 129.270 37.330 129.680 ;
        RECT 37.565 129.270 37.735 130.030 ;
        RECT 37.905 129.690 39.935 129.860 ;
        RECT 36.815 128.460 37.155 129.270 ;
        RECT 37.905 129.025 38.075 129.690 ;
        RECT 38.470 129.350 39.595 129.520 ;
        RECT 37.325 128.835 38.075 129.025 ;
        RECT 38.245 129.010 39.255 129.180 ;
        RECT 36.815 128.290 38.045 128.460 ;
        RECT 35.205 127.480 35.455 127.940 ;
        RECT 35.625 127.650 36.185 127.940 ;
        RECT 37.090 127.685 37.335 128.290 ;
        RECT 37.555 127.480 38.065 128.015 ;
        RECT 38.245 127.650 38.435 129.010 ;
        RECT 38.605 127.990 38.880 128.810 ;
        RECT 39.085 128.210 39.255 129.010 ;
        RECT 39.425 128.220 39.595 129.350 ;
        RECT 39.765 128.720 39.935 129.690 ;
        RECT 40.105 128.890 40.275 130.030 ;
        RECT 40.445 128.890 40.780 129.860 ;
        RECT 39.765 128.390 39.960 128.720 ;
        RECT 40.185 128.390 40.440 128.720 ;
        RECT 40.185 128.220 40.355 128.390 ;
        RECT 40.610 128.220 40.780 128.890 ;
        RECT 40.955 128.865 41.245 130.030 ;
        RECT 42.250 129.050 42.505 129.720 ;
        RECT 42.685 129.230 42.970 130.030 ;
        RECT 43.150 129.310 43.480 129.820 ;
        RECT 42.250 128.330 42.430 129.050 ;
        RECT 43.150 128.720 43.400 129.310 ;
        RECT 43.750 129.160 43.920 129.770 ;
        RECT 44.090 129.340 44.420 130.030 ;
        RECT 44.650 129.480 44.890 129.770 ;
        RECT 45.090 129.650 45.510 130.030 ;
        RECT 45.690 129.560 46.320 129.810 ;
        RECT 46.790 129.650 47.120 130.030 ;
        RECT 45.690 129.480 45.860 129.560 ;
        RECT 47.290 129.480 47.460 129.770 ;
        RECT 47.640 129.650 48.020 130.030 ;
        RECT 48.260 129.645 49.090 129.815 ;
        RECT 44.650 129.310 45.860 129.480 ;
        RECT 42.600 128.390 43.400 128.720 ;
        RECT 39.425 128.050 40.355 128.220 ;
        RECT 39.425 128.015 39.600 128.050 ;
        RECT 38.605 127.820 38.885 127.990 ;
        RECT 38.605 127.650 38.880 127.820 ;
        RECT 39.070 127.650 39.600 128.015 ;
        RECT 40.025 127.480 40.355 127.880 ;
        RECT 40.525 127.650 40.780 128.220 ;
        RECT 40.955 127.480 41.245 128.205 ;
        RECT 42.165 128.190 42.430 128.330 ;
        RECT 42.165 128.160 42.505 128.190 ;
        RECT 42.250 127.660 42.505 128.160 ;
        RECT 42.685 127.480 42.970 127.940 ;
        RECT 43.150 127.740 43.400 128.390 ;
        RECT 43.600 129.140 43.920 129.160 ;
        RECT 43.600 128.970 45.520 129.140 ;
        RECT 43.600 128.075 43.790 128.970 ;
        RECT 45.690 128.800 45.860 129.310 ;
        RECT 46.030 129.050 46.550 129.360 ;
        RECT 43.960 128.630 45.860 128.800 ;
        RECT 43.960 128.570 44.290 128.630 ;
        RECT 44.440 128.400 44.770 128.460 ;
        RECT 44.110 128.130 44.770 128.400 ;
        RECT 43.600 127.745 43.920 128.075 ;
        RECT 44.100 127.480 44.760 127.960 ;
        RECT 44.960 127.870 45.130 128.630 ;
        RECT 46.030 128.460 46.210 128.870 ;
        RECT 45.300 128.290 45.630 128.410 ;
        RECT 46.380 128.290 46.550 129.050 ;
        RECT 45.300 128.120 46.550 128.290 ;
        RECT 46.720 129.230 48.090 129.480 ;
        RECT 46.720 128.460 46.910 129.230 ;
        RECT 47.840 128.970 48.090 129.230 ;
        RECT 47.080 128.800 47.330 128.960 ;
        RECT 48.260 128.800 48.430 129.645 ;
        RECT 49.325 129.360 49.495 129.860 ;
        RECT 49.665 129.530 49.995 130.030 ;
        RECT 48.600 128.970 49.100 129.350 ;
        RECT 49.325 129.190 50.020 129.360 ;
        RECT 47.080 128.630 48.430 128.800 ;
        RECT 48.010 128.590 48.430 128.630 ;
        RECT 46.720 128.120 47.140 128.460 ;
        RECT 47.430 128.130 47.840 128.460 ;
        RECT 44.960 127.700 45.810 127.870 ;
        RECT 46.370 127.480 46.690 127.940 ;
        RECT 46.890 127.690 47.140 128.120 ;
        RECT 47.430 127.480 47.840 127.920 ;
        RECT 48.010 127.860 48.180 128.590 ;
        RECT 48.350 128.040 48.700 128.410 ;
        RECT 48.880 128.100 49.100 128.970 ;
        RECT 49.270 128.400 49.680 129.020 ;
        RECT 49.850 128.220 50.020 129.190 ;
        RECT 49.325 128.030 50.020 128.220 ;
        RECT 48.010 127.660 49.025 127.860 ;
        RECT 49.325 127.700 49.495 128.030 ;
        RECT 49.665 127.480 49.995 127.860 ;
        RECT 50.210 127.740 50.435 129.860 ;
        RECT 50.605 129.530 50.935 130.030 ;
        RECT 51.105 129.360 51.275 129.860 ;
        RECT 50.610 129.190 51.275 129.360 ;
        RECT 50.610 128.200 50.840 129.190 ;
        RECT 51.010 128.370 51.360 129.020 ;
        RECT 51.595 128.890 51.805 130.030 ;
        RECT 51.975 128.880 52.305 129.860 ;
        RECT 52.475 128.890 52.705 130.030 ;
        RECT 53.375 128.955 53.645 129.860 ;
        RECT 53.815 129.270 54.145 130.030 ;
        RECT 54.325 129.100 54.495 129.860 ;
        RECT 50.610 128.030 51.275 128.200 ;
        RECT 50.605 127.480 50.935 127.860 ;
        RECT 51.105 127.740 51.275 128.030 ;
        RECT 51.595 127.480 51.805 128.300 ;
        RECT 51.975 128.280 52.225 128.880 ;
        RECT 52.395 128.470 52.725 128.720 ;
        RECT 51.975 127.650 52.305 128.280 ;
        RECT 52.475 127.480 52.705 128.300 ;
        RECT 53.375 128.155 53.545 128.955 ;
        RECT 53.830 128.930 54.495 129.100 ;
        RECT 55.215 129.060 55.495 130.030 ;
        RECT 53.830 128.785 54.000 128.930 ;
        RECT 53.715 128.455 54.000 128.785 ;
        RECT 53.830 128.200 54.000 128.455 ;
        RECT 54.235 128.380 54.565 128.750 ;
        RECT 55.665 128.685 55.995 129.860 ;
        RECT 56.165 129.060 56.425 130.030 ;
        RECT 57.430 129.690 57.685 129.720 ;
        RECT 57.345 129.520 57.685 129.690 ;
        RECT 57.430 129.050 57.685 129.520 ;
        RECT 57.865 129.230 58.150 130.030 ;
        RECT 58.330 129.310 58.660 129.820 ;
        RECT 53.375 127.650 53.635 128.155 ;
        RECT 53.830 128.030 54.495 128.200 ;
        RECT 55.215 128.155 55.995 128.685 ;
        RECT 53.815 127.480 54.145 127.860 ;
        RECT 54.325 127.650 54.495 128.030 ;
        RECT 55.215 127.480 55.500 127.985 ;
        RECT 55.670 127.650 55.995 128.155 ;
        RECT 56.185 127.770 56.425 128.720 ;
        RECT 57.430 128.190 57.610 129.050 ;
        RECT 58.330 128.720 58.580 129.310 ;
        RECT 58.930 129.160 59.100 129.770 ;
        RECT 59.270 129.340 59.600 130.030 ;
        RECT 59.830 129.480 60.070 129.770 ;
        RECT 60.270 129.650 60.690 130.030 ;
        RECT 60.870 129.560 61.500 129.810 ;
        RECT 61.970 129.650 62.300 130.030 ;
        RECT 60.870 129.480 61.040 129.560 ;
        RECT 62.470 129.480 62.640 129.770 ;
        RECT 62.820 129.650 63.200 130.030 ;
        RECT 63.440 129.645 64.270 129.815 ;
        RECT 59.830 129.310 61.040 129.480 ;
        RECT 57.780 128.390 58.580 128.720 ;
        RECT 57.430 127.660 57.685 128.190 ;
        RECT 57.865 127.480 58.150 127.940 ;
        RECT 58.330 127.740 58.580 128.390 ;
        RECT 58.780 129.140 59.100 129.160 ;
        RECT 58.780 128.970 60.700 129.140 ;
        RECT 58.780 128.075 58.970 128.970 ;
        RECT 60.870 128.800 61.040 129.310 ;
        RECT 61.210 129.050 61.730 129.360 ;
        RECT 59.140 128.630 61.040 128.800 ;
        RECT 59.140 128.570 59.470 128.630 ;
        RECT 59.620 128.400 59.950 128.460 ;
        RECT 59.290 128.130 59.950 128.400 ;
        RECT 58.780 127.745 59.100 128.075 ;
        RECT 59.280 127.480 59.940 127.960 ;
        RECT 60.140 127.870 60.310 128.630 ;
        RECT 61.210 128.460 61.390 128.870 ;
        RECT 60.480 128.290 60.810 128.410 ;
        RECT 61.560 128.290 61.730 129.050 ;
        RECT 60.480 128.120 61.730 128.290 ;
        RECT 61.900 129.230 63.270 129.480 ;
        RECT 61.900 128.460 62.090 129.230 ;
        RECT 63.020 128.970 63.270 129.230 ;
        RECT 62.260 128.800 62.510 128.960 ;
        RECT 63.440 128.800 63.610 129.645 ;
        RECT 64.505 129.360 64.675 129.860 ;
        RECT 64.845 129.530 65.175 130.030 ;
        RECT 63.780 128.970 64.280 129.350 ;
        RECT 64.505 129.190 65.200 129.360 ;
        RECT 62.260 128.630 63.610 128.800 ;
        RECT 63.190 128.590 63.610 128.630 ;
        RECT 61.900 128.120 62.320 128.460 ;
        RECT 62.610 128.130 63.020 128.460 ;
        RECT 60.140 127.700 60.990 127.870 ;
        RECT 61.550 127.480 61.870 127.940 ;
        RECT 62.070 127.690 62.320 128.120 ;
        RECT 62.610 127.480 63.020 127.920 ;
        RECT 63.190 127.860 63.360 128.590 ;
        RECT 63.530 128.040 63.880 128.410 ;
        RECT 64.060 128.100 64.280 128.970 ;
        RECT 64.450 128.400 64.860 129.020 ;
        RECT 65.030 128.220 65.200 129.190 ;
        RECT 64.505 128.030 65.200 128.220 ;
        RECT 63.190 127.660 64.205 127.860 ;
        RECT 64.505 127.700 64.675 128.030 ;
        RECT 64.845 127.480 65.175 127.860 ;
        RECT 65.390 127.740 65.615 129.860 ;
        RECT 65.785 129.530 66.115 130.030 ;
        RECT 66.285 129.360 66.455 129.860 ;
        RECT 65.790 129.190 66.455 129.360 ;
        RECT 65.790 128.200 66.020 129.190 ;
        RECT 66.190 128.370 66.540 129.020 ;
        RECT 66.715 128.865 67.005 130.030 ;
        RECT 67.635 128.940 70.225 130.030 ;
        RECT 70.770 129.690 71.025 129.720 ;
        RECT 70.685 129.520 71.025 129.690 ;
        RECT 70.770 129.050 71.025 129.520 ;
        RECT 71.205 129.230 71.490 130.030 ;
        RECT 71.670 129.310 72.000 129.820 ;
        RECT 67.635 128.420 68.845 128.940 ;
        RECT 69.015 128.250 70.225 128.770 ;
        RECT 65.790 128.030 66.455 128.200 ;
        RECT 65.785 127.480 66.115 127.860 ;
        RECT 66.285 127.740 66.455 128.030 ;
        RECT 66.715 127.480 67.005 128.205 ;
        RECT 67.635 127.480 70.225 128.250 ;
        RECT 70.770 128.190 70.950 129.050 ;
        RECT 71.670 128.720 71.920 129.310 ;
        RECT 72.270 129.160 72.440 129.770 ;
        RECT 72.610 129.340 72.940 130.030 ;
        RECT 73.170 129.480 73.410 129.770 ;
        RECT 73.610 129.650 74.030 130.030 ;
        RECT 74.210 129.560 74.840 129.810 ;
        RECT 75.310 129.650 75.640 130.030 ;
        RECT 74.210 129.480 74.380 129.560 ;
        RECT 75.810 129.480 75.980 129.770 ;
        RECT 76.160 129.650 76.540 130.030 ;
        RECT 76.780 129.645 77.610 129.815 ;
        RECT 73.170 129.310 74.380 129.480 ;
        RECT 71.120 128.390 71.920 128.720 ;
        RECT 70.770 127.660 71.025 128.190 ;
        RECT 71.205 127.480 71.490 127.940 ;
        RECT 71.670 127.740 71.920 128.390 ;
        RECT 72.120 129.140 72.440 129.160 ;
        RECT 72.120 128.970 74.040 129.140 ;
        RECT 72.120 128.075 72.310 128.970 ;
        RECT 74.210 128.800 74.380 129.310 ;
        RECT 74.550 129.050 75.070 129.360 ;
        RECT 72.480 128.630 74.380 128.800 ;
        RECT 72.480 128.570 72.810 128.630 ;
        RECT 72.960 128.400 73.290 128.460 ;
        RECT 72.630 128.130 73.290 128.400 ;
        RECT 72.120 127.745 72.440 128.075 ;
        RECT 72.620 127.480 73.280 127.960 ;
        RECT 73.480 127.870 73.650 128.630 ;
        RECT 74.550 128.460 74.730 128.870 ;
        RECT 73.820 128.290 74.150 128.410 ;
        RECT 74.900 128.290 75.070 129.050 ;
        RECT 73.820 128.120 75.070 128.290 ;
        RECT 75.240 129.230 76.610 129.480 ;
        RECT 75.240 128.460 75.430 129.230 ;
        RECT 76.360 128.970 76.610 129.230 ;
        RECT 75.600 128.800 75.850 128.960 ;
        RECT 76.780 128.800 76.950 129.645 ;
        RECT 77.845 129.360 78.015 129.860 ;
        RECT 78.185 129.530 78.515 130.030 ;
        RECT 77.120 128.970 77.620 129.350 ;
        RECT 77.845 129.190 78.540 129.360 ;
        RECT 75.600 128.630 76.950 128.800 ;
        RECT 76.530 128.590 76.950 128.630 ;
        RECT 75.240 128.120 75.660 128.460 ;
        RECT 75.950 128.130 76.360 128.460 ;
        RECT 73.480 127.700 74.330 127.870 ;
        RECT 74.890 127.480 75.210 127.940 ;
        RECT 75.410 127.690 75.660 128.120 ;
        RECT 75.950 127.480 76.360 127.920 ;
        RECT 76.530 127.860 76.700 128.590 ;
        RECT 76.870 128.040 77.220 128.410 ;
        RECT 77.400 128.100 77.620 128.970 ;
        RECT 77.790 128.400 78.200 129.020 ;
        RECT 78.370 128.220 78.540 129.190 ;
        RECT 77.845 128.030 78.540 128.220 ;
        RECT 76.530 127.660 77.545 127.860 ;
        RECT 77.845 127.700 78.015 128.030 ;
        RECT 78.185 127.480 78.515 127.860 ;
        RECT 78.730 127.740 78.955 129.860 ;
        RECT 79.125 129.530 79.455 130.030 ;
        RECT 79.625 129.360 79.795 129.860 ;
        RECT 79.130 129.190 79.795 129.360 ;
        RECT 80.145 129.285 80.415 130.030 ;
        RECT 81.045 130.025 87.320 130.030 ;
        RECT 79.130 128.200 79.360 129.190 ;
        RECT 80.585 129.115 80.875 129.855 ;
        RECT 81.045 129.300 81.300 130.025 ;
        RECT 81.485 129.130 81.745 129.855 ;
        RECT 81.915 129.300 82.160 130.025 ;
        RECT 82.345 129.130 82.605 129.855 ;
        RECT 82.775 129.300 83.020 130.025 ;
        RECT 83.205 129.130 83.465 129.855 ;
        RECT 83.635 129.300 83.880 130.025 ;
        RECT 84.050 129.130 84.310 129.855 ;
        RECT 84.480 129.300 84.740 130.025 ;
        RECT 84.910 129.130 85.170 129.855 ;
        RECT 85.340 129.300 85.600 130.025 ;
        RECT 85.770 129.130 86.030 129.855 ;
        RECT 86.200 129.300 86.460 130.025 ;
        RECT 86.630 129.130 86.890 129.855 ;
        RECT 87.060 129.230 87.320 130.025 ;
        RECT 81.485 129.115 86.890 129.130 ;
        RECT 79.530 128.370 79.880 129.020 ;
        RECT 80.145 128.890 86.890 129.115 ;
        RECT 80.145 128.300 81.310 128.890 ;
        RECT 87.490 128.720 87.740 129.855 ;
        RECT 87.920 129.220 88.180 130.030 ;
        RECT 88.355 128.720 88.600 129.860 ;
        RECT 88.780 129.220 89.075 130.030 ;
        RECT 89.295 128.890 89.525 130.030 ;
        RECT 89.695 128.880 90.025 129.860 ;
        RECT 90.195 128.890 90.405 130.030 ;
        RECT 90.635 128.940 92.305 130.030 ;
        RECT 81.480 128.470 88.600 128.720 ;
        RECT 79.130 128.030 79.795 128.200 ;
        RECT 80.145 128.130 86.890 128.300 ;
        RECT 79.125 127.480 79.455 127.860 ;
        RECT 79.625 127.740 79.795 128.030 ;
        RECT 80.145 127.480 80.445 127.960 ;
        RECT 80.615 127.675 80.875 128.130 ;
        RECT 81.045 127.480 81.305 127.960 ;
        RECT 81.485 127.675 81.745 128.130 ;
        RECT 81.915 127.480 82.165 127.960 ;
        RECT 82.345 127.675 82.605 128.130 ;
        RECT 82.775 127.480 83.025 127.960 ;
        RECT 83.205 127.675 83.465 128.130 ;
        RECT 83.635 127.480 83.880 127.960 ;
        RECT 84.050 127.675 84.325 128.130 ;
        RECT 84.495 127.480 84.740 127.960 ;
        RECT 84.910 127.675 85.170 128.130 ;
        RECT 85.340 127.480 85.600 127.960 ;
        RECT 85.770 127.675 86.030 128.130 ;
        RECT 86.200 127.480 86.460 127.960 ;
        RECT 86.630 127.675 86.890 128.130 ;
        RECT 87.060 127.480 87.320 128.040 ;
        RECT 87.490 127.660 87.740 128.470 ;
        RECT 87.920 127.480 88.180 128.005 ;
        RECT 88.350 127.660 88.600 128.470 ;
        RECT 88.770 128.160 89.085 128.720 ;
        RECT 89.275 128.470 89.605 128.720 ;
        RECT 88.780 127.480 89.085 127.990 ;
        RECT 89.295 127.480 89.525 128.300 ;
        RECT 89.775 128.280 90.025 128.880 ;
        RECT 90.635 128.420 91.385 128.940 ;
        RECT 92.475 128.865 92.765 130.030 ;
        RECT 93.395 128.940 95.065 130.030 ;
        RECT 95.325 129.100 95.495 129.860 ;
        RECT 95.675 129.270 96.005 130.030 ;
        RECT 89.695 127.650 90.025 128.280 ;
        RECT 90.195 127.480 90.405 128.300 ;
        RECT 91.555 128.250 92.305 128.770 ;
        RECT 93.395 128.420 94.145 128.940 ;
        RECT 95.325 128.930 95.990 129.100 ;
        RECT 96.175 128.955 96.445 129.860 ;
        RECT 96.625 129.220 96.920 130.030 ;
        RECT 95.820 128.785 95.990 128.930 ;
        RECT 94.315 128.250 95.065 128.770 ;
        RECT 95.255 128.380 95.585 128.750 ;
        RECT 95.820 128.455 96.105 128.785 ;
        RECT 90.635 127.480 92.305 128.250 ;
        RECT 92.475 127.480 92.765 128.205 ;
        RECT 93.395 127.480 95.065 128.250 ;
        RECT 95.820 128.200 95.990 128.455 ;
        RECT 95.325 128.030 95.990 128.200 ;
        RECT 96.275 128.155 96.445 128.955 ;
        RECT 97.100 128.720 97.345 129.860 ;
        RECT 97.520 129.220 97.780 130.030 ;
        RECT 98.380 130.025 104.655 130.030 ;
        RECT 97.960 128.720 98.210 129.855 ;
        RECT 98.380 129.230 98.640 130.025 ;
        RECT 98.810 129.130 99.070 129.855 ;
        RECT 99.240 129.300 99.500 130.025 ;
        RECT 99.670 129.130 99.930 129.855 ;
        RECT 100.100 129.300 100.360 130.025 ;
        RECT 100.530 129.130 100.790 129.855 ;
        RECT 100.960 129.300 101.220 130.025 ;
        RECT 101.390 129.130 101.650 129.855 ;
        RECT 101.820 129.300 102.065 130.025 ;
        RECT 102.235 129.130 102.495 129.855 ;
        RECT 102.680 129.300 102.925 130.025 ;
        RECT 103.095 129.130 103.355 129.855 ;
        RECT 103.540 129.300 103.785 130.025 ;
        RECT 103.955 129.130 104.215 129.855 ;
        RECT 104.400 129.300 104.655 130.025 ;
        RECT 98.810 129.115 104.215 129.130 ;
        RECT 104.825 129.115 105.115 129.855 ;
        RECT 105.285 129.285 105.555 130.030 ;
        RECT 105.815 129.270 106.330 129.680 ;
        RECT 106.565 129.270 106.735 130.030 ;
        RECT 106.905 129.690 108.935 129.860 ;
        RECT 98.810 128.890 105.555 129.115 ;
        RECT 96.615 128.160 96.930 128.720 ;
        RECT 97.100 128.470 104.220 128.720 ;
        RECT 95.325 127.650 95.495 128.030 ;
        RECT 95.675 127.480 96.005 127.860 ;
        RECT 96.185 127.650 96.445 128.155 ;
        RECT 96.615 127.480 96.920 127.990 ;
        RECT 97.100 127.660 97.350 128.470 ;
        RECT 97.520 127.480 97.780 128.005 ;
        RECT 97.960 127.660 98.210 128.470 ;
        RECT 104.390 128.330 105.555 128.890 ;
        RECT 105.815 128.460 106.155 129.270 ;
        RECT 106.905 129.025 107.075 129.690 ;
        RECT 107.470 129.350 108.595 129.520 ;
        RECT 106.325 128.835 107.075 129.025 ;
        RECT 107.245 129.010 108.255 129.180 ;
        RECT 104.390 128.300 105.585 128.330 ;
        RECT 98.810 128.160 105.585 128.300 ;
        RECT 105.815 128.290 107.045 128.460 ;
        RECT 98.810 128.130 105.555 128.160 ;
        RECT 98.380 127.480 98.640 128.040 ;
        RECT 98.810 127.675 99.070 128.130 ;
        RECT 99.240 127.480 99.500 127.960 ;
        RECT 99.670 127.675 99.930 128.130 ;
        RECT 100.100 127.480 100.360 127.960 ;
        RECT 100.530 127.675 100.790 128.130 ;
        RECT 100.960 127.480 101.205 127.960 ;
        RECT 101.375 127.675 101.650 128.130 ;
        RECT 101.820 127.480 102.065 127.960 ;
        RECT 102.235 127.675 102.495 128.130 ;
        RECT 102.675 127.480 102.925 127.960 ;
        RECT 103.095 127.675 103.355 128.130 ;
        RECT 103.535 127.480 103.785 127.960 ;
        RECT 103.955 127.675 104.215 128.130 ;
        RECT 104.395 127.480 104.655 127.960 ;
        RECT 104.825 127.675 105.085 128.130 ;
        RECT 105.255 127.480 105.555 127.960 ;
        RECT 106.090 127.685 106.335 128.290 ;
        RECT 106.555 127.480 107.065 128.015 ;
        RECT 107.245 127.650 107.435 129.010 ;
        RECT 107.605 128.670 107.880 128.810 ;
        RECT 107.605 128.500 107.885 128.670 ;
        RECT 107.605 127.650 107.880 128.500 ;
        RECT 108.085 128.210 108.255 129.010 ;
        RECT 108.425 128.220 108.595 129.350 ;
        RECT 108.765 128.720 108.935 129.690 ;
        RECT 109.105 128.890 109.275 130.030 ;
        RECT 109.445 128.890 109.780 129.860 ;
        RECT 109.955 129.060 110.235 130.030 ;
        RECT 108.765 128.390 108.960 128.720 ;
        RECT 109.185 128.390 109.440 128.720 ;
        RECT 109.185 128.220 109.355 128.390 ;
        RECT 109.610 128.220 109.780 128.890 ;
        RECT 110.405 128.685 110.735 129.860 ;
        RECT 110.905 129.060 111.165 130.030 ;
        RECT 111.395 128.890 111.605 130.030 ;
        RECT 111.775 128.880 112.105 129.860 ;
        RECT 112.275 128.890 112.505 130.030 ;
        RECT 112.805 129.100 112.975 129.860 ;
        RECT 113.155 129.270 113.485 130.030 ;
        RECT 112.805 128.930 113.470 129.100 ;
        RECT 113.655 128.955 113.925 129.860 ;
        RECT 108.425 128.050 109.355 128.220 ;
        RECT 108.425 128.015 108.600 128.050 ;
        RECT 108.070 127.650 108.600 128.015 ;
        RECT 109.025 127.480 109.355 127.880 ;
        RECT 109.525 127.650 109.780 128.220 ;
        RECT 109.955 128.155 110.735 128.685 ;
        RECT 109.955 127.480 110.240 127.985 ;
        RECT 110.410 127.650 110.735 128.155 ;
        RECT 110.925 127.770 111.165 128.720 ;
        RECT 111.395 127.480 111.605 128.300 ;
        RECT 111.775 128.280 112.025 128.880 ;
        RECT 113.300 128.785 113.470 128.930 ;
        RECT 112.195 128.470 112.525 128.720 ;
        RECT 112.735 128.380 113.065 128.750 ;
        RECT 113.300 128.455 113.585 128.785 ;
        RECT 111.775 127.650 112.105 128.280 ;
        RECT 112.275 127.480 112.505 128.300 ;
        RECT 113.300 128.200 113.470 128.455 ;
        RECT 112.805 128.030 113.470 128.200 ;
        RECT 113.755 128.155 113.925 128.955 ;
        RECT 114.555 128.940 117.145 130.030 ;
        RECT 117.315 128.940 118.525 130.030 ;
        RECT 114.555 128.420 115.765 128.940 ;
        RECT 115.935 128.250 117.145 128.770 ;
        RECT 117.315 128.400 117.835 128.940 ;
        RECT 112.805 127.650 112.975 128.030 ;
        RECT 113.155 127.480 113.485 127.860 ;
        RECT 113.665 127.650 113.925 128.155 ;
        RECT 114.555 127.480 117.145 128.250 ;
        RECT 118.005 128.230 118.525 128.770 ;
        RECT 117.315 127.480 118.525 128.230 ;
        RECT 11.430 127.310 118.610 127.480 ;
        RECT 11.515 126.560 12.725 127.310 ;
        RECT 14.190 126.600 14.445 127.130 ;
        RECT 14.625 126.850 14.910 127.310 ;
        RECT 11.515 126.020 12.035 126.560 ;
        RECT 12.205 125.850 12.725 126.390 ;
        RECT 14.190 125.950 14.370 126.600 ;
        RECT 15.090 126.400 15.340 127.050 ;
        RECT 14.540 126.070 15.340 126.400 ;
        RECT 11.515 124.760 12.725 125.850 ;
        RECT 14.105 125.780 14.370 125.950 ;
        RECT 14.190 125.740 14.370 125.780 ;
        RECT 14.190 125.070 14.445 125.740 ;
        RECT 14.625 124.760 14.910 125.560 ;
        RECT 15.090 125.480 15.340 126.070 ;
        RECT 15.540 126.715 15.860 127.045 ;
        RECT 16.040 126.830 16.700 127.310 ;
        RECT 16.900 126.920 17.750 127.090 ;
        RECT 15.540 125.820 15.730 126.715 ;
        RECT 16.050 126.390 16.710 126.660 ;
        RECT 16.380 126.330 16.710 126.390 ;
        RECT 15.900 126.160 16.230 126.220 ;
        RECT 16.900 126.160 17.070 126.920 ;
        RECT 18.310 126.850 18.630 127.310 ;
        RECT 18.830 126.670 19.080 127.100 ;
        RECT 19.370 126.870 19.780 127.310 ;
        RECT 19.950 126.930 20.965 127.130 ;
        RECT 17.240 126.500 18.490 126.670 ;
        RECT 17.240 126.380 17.570 126.500 ;
        RECT 15.900 125.990 17.800 126.160 ;
        RECT 15.540 125.650 17.460 125.820 ;
        RECT 15.540 125.630 15.860 125.650 ;
        RECT 15.090 124.970 15.420 125.480 ;
        RECT 15.690 125.020 15.860 125.630 ;
        RECT 17.630 125.480 17.800 125.990 ;
        RECT 17.970 125.920 18.150 126.330 ;
        RECT 18.320 125.740 18.490 126.500 ;
        RECT 16.030 124.760 16.360 125.450 ;
        RECT 16.590 125.310 17.800 125.480 ;
        RECT 17.970 125.430 18.490 125.740 ;
        RECT 18.660 126.330 19.080 126.670 ;
        RECT 19.370 126.330 19.780 126.660 ;
        RECT 18.660 125.560 18.850 126.330 ;
        RECT 19.950 126.200 20.120 126.930 ;
        RECT 21.265 126.760 21.435 127.090 ;
        RECT 21.605 126.930 21.935 127.310 ;
        RECT 20.290 126.380 20.640 126.750 ;
        RECT 19.950 126.160 20.370 126.200 ;
        RECT 19.020 125.990 20.370 126.160 ;
        RECT 19.020 125.830 19.270 125.990 ;
        RECT 19.780 125.560 20.030 125.820 ;
        RECT 18.660 125.310 20.030 125.560 ;
        RECT 16.590 125.020 16.830 125.310 ;
        RECT 17.630 125.230 17.800 125.310 ;
        RECT 17.030 124.760 17.450 125.140 ;
        RECT 17.630 124.980 18.260 125.230 ;
        RECT 18.730 124.760 19.060 125.140 ;
        RECT 19.230 125.020 19.400 125.310 ;
        RECT 20.200 125.145 20.370 125.990 ;
        RECT 20.820 125.820 21.040 126.690 ;
        RECT 21.265 126.570 21.960 126.760 ;
        RECT 20.540 125.440 21.040 125.820 ;
        RECT 21.210 125.770 21.620 126.390 ;
        RECT 21.790 125.600 21.960 126.570 ;
        RECT 21.265 125.430 21.960 125.600 ;
        RECT 19.580 124.760 19.960 125.140 ;
        RECT 20.200 124.975 21.030 125.145 ;
        RECT 21.265 124.930 21.435 125.430 ;
        RECT 21.605 124.760 21.935 125.260 ;
        RECT 22.150 124.930 22.375 127.050 ;
        RECT 22.545 126.930 22.875 127.310 ;
        RECT 23.045 126.760 23.215 127.050 ;
        RECT 22.550 126.590 23.215 126.760 ;
        RECT 22.550 125.600 22.780 126.590 ;
        RECT 23.975 126.490 24.205 127.310 ;
        RECT 24.375 126.510 24.705 127.140 ;
        RECT 22.950 125.770 23.300 126.420 ;
        RECT 23.955 126.070 24.285 126.320 ;
        RECT 24.455 125.910 24.705 126.510 ;
        RECT 24.875 126.490 25.085 127.310 ;
        RECT 25.375 126.830 25.655 127.310 ;
        RECT 25.825 126.660 26.085 127.050 ;
        RECT 26.260 126.830 26.515 127.310 ;
        RECT 26.685 126.660 26.980 127.050 ;
        RECT 27.160 126.830 27.435 127.310 ;
        RECT 27.605 126.810 27.905 127.140 ;
        RECT 25.330 126.490 26.980 126.660 ;
        RECT 22.550 125.430 23.215 125.600 ;
        RECT 22.545 124.760 22.875 125.260 ;
        RECT 23.045 124.930 23.215 125.430 ;
        RECT 23.975 124.760 24.205 125.900 ;
        RECT 24.375 124.930 24.705 125.910 ;
        RECT 25.330 125.980 25.735 126.490 ;
        RECT 25.905 126.150 27.045 126.320 ;
        RECT 24.875 124.760 25.085 125.900 ;
        RECT 25.330 125.810 26.085 125.980 ;
        RECT 25.370 124.760 25.655 125.630 ;
        RECT 25.825 125.560 26.085 125.810 ;
        RECT 26.875 125.900 27.045 126.150 ;
        RECT 27.215 126.070 27.565 126.640 ;
        RECT 27.735 125.900 27.905 126.810 ;
        RECT 28.075 126.585 28.365 127.310 ;
        RECT 28.810 126.500 29.055 127.105 ;
        RECT 29.275 126.775 29.785 127.310 ;
        RECT 28.535 126.330 29.765 126.500 ;
        RECT 26.875 125.730 27.905 125.900 ;
        RECT 25.825 125.390 26.945 125.560 ;
        RECT 25.825 124.930 26.085 125.390 ;
        RECT 26.260 124.760 26.515 125.220 ;
        RECT 26.685 124.930 26.945 125.390 ;
        RECT 27.115 124.760 27.425 125.560 ;
        RECT 27.595 124.930 27.905 125.730 ;
        RECT 28.075 124.760 28.365 125.925 ;
        RECT 28.535 125.520 28.875 126.330 ;
        RECT 29.045 125.765 29.795 125.955 ;
        RECT 28.535 125.110 29.050 125.520 ;
        RECT 29.285 124.760 29.455 125.520 ;
        RECT 29.625 125.100 29.795 125.765 ;
        RECT 29.965 125.780 30.155 127.140 ;
        RECT 30.325 126.290 30.600 127.140 ;
        RECT 30.790 126.775 31.320 127.140 ;
        RECT 31.745 126.910 32.075 127.310 ;
        RECT 31.145 126.740 31.320 126.775 ;
        RECT 30.325 126.120 30.605 126.290 ;
        RECT 30.325 125.980 30.600 126.120 ;
        RECT 30.805 125.780 30.975 126.580 ;
        RECT 29.965 125.610 30.975 125.780 ;
        RECT 31.145 126.570 32.075 126.740 ;
        RECT 32.245 126.570 32.500 127.140 ;
        RECT 31.145 125.440 31.315 126.570 ;
        RECT 31.905 126.400 32.075 126.570 ;
        RECT 30.190 125.270 31.315 125.440 ;
        RECT 31.485 126.070 31.680 126.400 ;
        RECT 31.905 126.070 32.160 126.400 ;
        RECT 31.485 125.100 31.655 126.070 ;
        RECT 32.330 125.900 32.500 126.570 ;
        RECT 32.675 126.560 33.885 127.310 ;
        RECT 34.430 126.970 34.685 127.130 ;
        RECT 34.345 126.800 34.685 126.970 ;
        RECT 34.865 126.850 35.150 127.310 ;
        RECT 29.625 124.930 31.655 125.100 ;
        RECT 31.825 124.760 31.995 125.900 ;
        RECT 32.165 124.930 32.500 125.900 ;
        RECT 32.675 125.850 33.195 126.390 ;
        RECT 33.365 126.020 33.885 126.560 ;
        RECT 34.430 126.600 34.685 126.800 ;
        RECT 32.675 124.760 33.885 125.850 ;
        RECT 34.430 125.740 34.610 126.600 ;
        RECT 35.330 126.400 35.580 127.050 ;
        RECT 34.780 126.070 35.580 126.400 ;
        RECT 34.430 125.070 34.685 125.740 ;
        RECT 34.865 124.760 35.150 125.560 ;
        RECT 35.330 125.480 35.580 126.070 ;
        RECT 35.780 126.715 36.100 127.045 ;
        RECT 36.280 126.830 36.940 127.310 ;
        RECT 37.140 126.920 37.990 127.090 ;
        RECT 35.780 125.820 35.970 126.715 ;
        RECT 36.290 126.390 36.950 126.660 ;
        RECT 36.620 126.330 36.950 126.390 ;
        RECT 36.140 126.160 36.470 126.220 ;
        RECT 37.140 126.160 37.310 126.920 ;
        RECT 38.550 126.850 38.870 127.310 ;
        RECT 39.070 126.670 39.320 127.100 ;
        RECT 39.610 126.870 40.020 127.310 ;
        RECT 40.190 126.930 41.205 127.130 ;
        RECT 37.480 126.500 38.730 126.670 ;
        RECT 37.480 126.380 37.810 126.500 ;
        RECT 36.140 125.990 38.040 126.160 ;
        RECT 35.780 125.650 37.700 125.820 ;
        RECT 35.780 125.630 36.100 125.650 ;
        RECT 35.330 124.970 35.660 125.480 ;
        RECT 35.930 125.020 36.100 125.630 ;
        RECT 37.870 125.480 38.040 125.990 ;
        RECT 38.210 125.920 38.390 126.330 ;
        RECT 38.560 125.740 38.730 126.500 ;
        RECT 36.270 124.760 36.600 125.450 ;
        RECT 36.830 125.310 38.040 125.480 ;
        RECT 38.210 125.430 38.730 125.740 ;
        RECT 38.900 126.330 39.320 126.670 ;
        RECT 39.610 126.330 40.020 126.660 ;
        RECT 38.900 125.560 39.090 126.330 ;
        RECT 40.190 126.200 40.360 126.930 ;
        RECT 41.505 126.760 41.675 127.090 ;
        RECT 41.845 126.930 42.175 127.310 ;
        RECT 40.530 126.380 40.880 126.750 ;
        RECT 40.190 126.160 40.610 126.200 ;
        RECT 39.260 125.990 40.610 126.160 ;
        RECT 39.260 125.830 39.510 125.990 ;
        RECT 40.020 125.560 40.270 125.820 ;
        RECT 38.900 125.310 40.270 125.560 ;
        RECT 36.830 125.020 37.070 125.310 ;
        RECT 37.870 125.230 38.040 125.310 ;
        RECT 37.270 124.760 37.690 125.140 ;
        RECT 37.870 124.980 38.500 125.230 ;
        RECT 38.970 124.760 39.300 125.140 ;
        RECT 39.470 125.020 39.640 125.310 ;
        RECT 40.440 125.145 40.610 125.990 ;
        RECT 41.060 125.820 41.280 126.690 ;
        RECT 41.505 126.570 42.200 126.760 ;
        RECT 40.780 125.440 41.280 125.820 ;
        RECT 41.450 125.770 41.860 126.390 ;
        RECT 42.030 125.600 42.200 126.570 ;
        RECT 41.505 125.430 42.200 125.600 ;
        RECT 39.820 124.760 40.200 125.140 ;
        RECT 40.440 124.975 41.270 125.145 ;
        RECT 41.505 124.930 41.675 125.430 ;
        RECT 41.845 124.760 42.175 125.260 ;
        RECT 42.390 124.930 42.615 127.050 ;
        RECT 42.785 126.930 43.115 127.310 ;
        RECT 43.285 126.760 43.455 127.050 ;
        RECT 42.790 126.590 43.455 126.760 ;
        RECT 44.550 126.600 44.805 127.130 ;
        RECT 44.985 126.850 45.270 127.310 ;
        RECT 42.790 125.600 43.020 126.590 ;
        RECT 43.190 125.770 43.540 126.420 ;
        RECT 44.550 126.290 44.730 126.600 ;
        RECT 45.450 126.400 45.700 127.050 ;
        RECT 44.465 126.120 44.730 126.290 ;
        RECT 44.550 125.740 44.730 126.120 ;
        RECT 44.900 126.070 45.700 126.400 ;
        RECT 42.790 125.430 43.455 125.600 ;
        RECT 42.785 124.760 43.115 125.260 ;
        RECT 43.285 124.930 43.455 125.430 ;
        RECT 44.550 125.070 44.805 125.740 ;
        RECT 44.985 124.760 45.270 125.560 ;
        RECT 45.450 125.480 45.700 126.070 ;
        RECT 45.900 126.715 46.220 127.045 ;
        RECT 46.400 126.830 47.060 127.310 ;
        RECT 47.260 126.920 48.110 127.090 ;
        RECT 45.900 125.820 46.090 126.715 ;
        RECT 46.410 126.390 47.070 126.660 ;
        RECT 46.740 126.330 47.070 126.390 ;
        RECT 46.260 126.160 46.590 126.220 ;
        RECT 47.260 126.160 47.430 126.920 ;
        RECT 48.670 126.850 48.990 127.310 ;
        RECT 49.190 126.670 49.440 127.100 ;
        RECT 49.730 126.870 50.140 127.310 ;
        RECT 50.310 126.930 51.325 127.130 ;
        RECT 47.600 126.500 48.850 126.670 ;
        RECT 47.600 126.380 47.930 126.500 ;
        RECT 46.260 125.990 48.160 126.160 ;
        RECT 45.900 125.650 47.820 125.820 ;
        RECT 45.900 125.630 46.220 125.650 ;
        RECT 45.450 124.970 45.780 125.480 ;
        RECT 46.050 125.020 46.220 125.630 ;
        RECT 47.990 125.480 48.160 125.990 ;
        RECT 48.330 125.920 48.510 126.330 ;
        RECT 48.680 125.740 48.850 126.500 ;
        RECT 46.390 124.760 46.720 125.450 ;
        RECT 46.950 125.310 48.160 125.480 ;
        RECT 48.330 125.430 48.850 125.740 ;
        RECT 49.020 126.330 49.440 126.670 ;
        RECT 49.730 126.330 50.140 126.660 ;
        RECT 49.020 125.560 49.210 126.330 ;
        RECT 50.310 126.200 50.480 126.930 ;
        RECT 51.625 126.760 51.795 127.090 ;
        RECT 51.965 126.930 52.295 127.310 ;
        RECT 50.650 126.380 51.000 126.750 ;
        RECT 50.310 126.160 50.730 126.200 ;
        RECT 49.380 125.990 50.730 126.160 ;
        RECT 49.380 125.830 49.630 125.990 ;
        RECT 50.140 125.560 50.390 125.820 ;
        RECT 49.020 125.310 50.390 125.560 ;
        RECT 46.950 125.020 47.190 125.310 ;
        RECT 47.990 125.230 48.160 125.310 ;
        RECT 47.390 124.760 47.810 125.140 ;
        RECT 47.990 124.980 48.620 125.230 ;
        RECT 49.090 124.760 49.420 125.140 ;
        RECT 49.590 125.020 49.760 125.310 ;
        RECT 50.560 125.145 50.730 125.990 ;
        RECT 51.180 125.820 51.400 126.690 ;
        RECT 51.625 126.570 52.320 126.760 ;
        RECT 50.900 125.440 51.400 125.820 ;
        RECT 51.570 125.770 51.980 126.390 ;
        RECT 52.150 125.600 52.320 126.570 ;
        RECT 51.625 125.430 52.320 125.600 ;
        RECT 49.940 124.760 50.320 125.140 ;
        RECT 50.560 124.975 51.390 125.145 ;
        RECT 51.625 124.930 51.795 125.430 ;
        RECT 51.965 124.760 52.295 125.260 ;
        RECT 52.510 124.930 52.735 127.050 ;
        RECT 52.905 126.930 53.235 127.310 ;
        RECT 53.405 126.760 53.575 127.050 ;
        RECT 52.910 126.590 53.575 126.760 ;
        RECT 52.910 125.600 53.140 126.590 ;
        RECT 53.835 126.585 54.125 127.310 ;
        RECT 54.300 126.570 54.555 127.140 ;
        RECT 54.725 126.910 55.055 127.310 ;
        RECT 55.480 126.775 56.010 127.140 ;
        RECT 56.200 126.970 56.475 127.140 ;
        RECT 56.195 126.800 56.475 126.970 ;
        RECT 55.480 126.740 55.655 126.775 ;
        RECT 54.725 126.570 55.655 126.740 ;
        RECT 53.310 125.770 53.660 126.420 ;
        RECT 52.910 125.430 53.575 125.600 ;
        RECT 52.905 124.760 53.235 125.260 ;
        RECT 53.405 124.930 53.575 125.430 ;
        RECT 53.835 124.760 54.125 125.925 ;
        RECT 54.300 125.900 54.470 126.570 ;
        RECT 54.725 126.400 54.895 126.570 ;
        RECT 54.640 126.070 54.895 126.400 ;
        RECT 55.120 126.070 55.315 126.400 ;
        RECT 54.300 124.930 54.635 125.900 ;
        RECT 54.805 124.760 54.975 125.900 ;
        RECT 55.145 125.100 55.315 126.070 ;
        RECT 55.485 125.440 55.655 126.570 ;
        RECT 55.825 125.780 55.995 126.580 ;
        RECT 56.200 125.980 56.475 126.800 ;
        RECT 56.645 125.780 56.835 127.140 ;
        RECT 57.015 126.775 57.525 127.310 ;
        RECT 57.745 126.500 57.990 127.105 ;
        RECT 59.355 126.540 62.865 127.310 ;
        RECT 57.035 126.330 58.265 126.500 ;
        RECT 55.825 125.610 56.835 125.780 ;
        RECT 57.005 125.765 57.755 125.955 ;
        RECT 55.485 125.270 56.610 125.440 ;
        RECT 57.005 125.100 57.175 125.765 ;
        RECT 57.925 125.520 58.265 126.330 ;
        RECT 55.145 124.930 57.175 125.100 ;
        RECT 57.345 124.760 57.515 125.520 ;
        RECT 57.750 125.110 58.265 125.520 ;
        RECT 59.355 125.850 61.045 126.370 ;
        RECT 61.215 126.020 62.865 126.540 ;
        RECT 63.095 126.490 63.305 127.310 ;
        RECT 63.475 126.510 63.805 127.140 ;
        RECT 63.475 125.910 63.725 126.510 ;
        RECT 63.975 126.490 64.205 127.310 ;
        RECT 64.875 126.540 66.545 127.310 ;
        RECT 66.720 126.765 72.065 127.310 ;
        RECT 63.895 126.070 64.225 126.320 ;
        RECT 59.355 124.760 62.865 125.850 ;
        RECT 63.095 124.760 63.305 125.900 ;
        RECT 63.475 124.930 63.805 125.910 ;
        RECT 63.975 124.760 64.205 125.900 ;
        RECT 64.875 125.850 65.625 126.370 ;
        RECT 65.795 126.020 66.545 126.540 ;
        RECT 64.875 124.760 66.545 125.850 ;
        RECT 68.310 125.195 68.660 126.445 ;
        RECT 70.140 125.935 70.480 126.765 ;
        RECT 72.275 126.490 72.505 127.310 ;
        RECT 72.675 126.510 73.005 127.140 ;
        RECT 72.255 126.070 72.585 126.320 ;
        RECT 72.755 125.910 73.005 126.510 ;
        RECT 73.175 126.490 73.385 127.310 ;
        RECT 73.655 126.490 73.885 127.310 ;
        RECT 74.055 126.510 74.385 127.140 ;
        RECT 73.635 126.070 73.965 126.320 ;
        RECT 74.135 125.910 74.385 126.510 ;
        RECT 74.555 126.490 74.765 127.310 ;
        RECT 75.730 126.500 75.975 127.105 ;
        RECT 76.195 126.775 76.705 127.310 ;
        RECT 66.720 124.760 72.065 125.195 ;
        RECT 72.275 124.760 72.505 125.900 ;
        RECT 72.675 124.930 73.005 125.910 ;
        RECT 73.175 124.760 73.385 125.900 ;
        RECT 73.655 124.760 73.885 125.900 ;
        RECT 74.055 124.930 74.385 125.910 ;
        RECT 75.455 126.330 76.685 126.500 ;
        RECT 74.555 124.760 74.765 125.900 ;
        RECT 75.455 125.520 75.795 126.330 ;
        RECT 75.965 125.765 76.715 125.955 ;
        RECT 75.455 125.110 75.970 125.520 ;
        RECT 76.205 124.760 76.375 125.520 ;
        RECT 76.545 125.100 76.715 125.765 ;
        RECT 76.885 125.780 77.075 127.140 ;
        RECT 77.245 126.290 77.520 127.140 ;
        RECT 77.710 126.775 78.240 127.140 ;
        RECT 78.665 126.910 78.995 127.310 ;
        RECT 78.065 126.740 78.240 126.775 ;
        RECT 77.245 126.120 77.525 126.290 ;
        RECT 77.245 125.980 77.520 126.120 ;
        RECT 77.725 125.780 77.895 126.580 ;
        RECT 76.885 125.610 77.895 125.780 ;
        RECT 78.065 126.570 78.995 126.740 ;
        RECT 79.165 126.570 79.420 127.140 ;
        RECT 79.595 126.585 79.885 127.310 ;
        RECT 78.065 125.440 78.235 126.570 ;
        RECT 78.825 126.400 78.995 126.570 ;
        RECT 77.110 125.270 78.235 125.440 ;
        RECT 78.405 126.070 78.600 126.400 ;
        RECT 78.825 126.070 79.080 126.400 ;
        RECT 78.405 125.100 78.575 126.070 ;
        RECT 79.250 125.900 79.420 126.570 ;
        RECT 80.055 126.540 81.725 127.310 ;
        RECT 76.545 124.930 78.575 125.100 ;
        RECT 78.745 124.760 78.915 125.900 ;
        RECT 79.085 124.930 79.420 125.900 ;
        RECT 79.595 124.760 79.885 125.925 ;
        RECT 80.055 125.850 80.805 126.370 ;
        RECT 80.975 126.020 81.725 126.540 ;
        RECT 81.935 126.490 82.165 127.310 ;
        RECT 82.335 126.510 82.665 127.140 ;
        RECT 81.915 126.070 82.245 126.320 ;
        RECT 82.415 125.910 82.665 126.510 ;
        RECT 82.835 126.490 83.045 127.310 ;
        RECT 83.550 126.500 83.795 127.105 ;
        RECT 84.015 126.775 84.525 127.310 ;
        RECT 80.055 124.760 81.725 125.850 ;
        RECT 81.935 124.760 82.165 125.900 ;
        RECT 82.335 124.930 82.665 125.910 ;
        RECT 83.275 126.330 84.505 126.500 ;
        RECT 82.835 124.760 83.045 125.900 ;
        RECT 83.275 125.520 83.615 126.330 ;
        RECT 83.785 125.765 84.535 125.955 ;
        RECT 83.275 125.110 83.790 125.520 ;
        RECT 84.025 124.760 84.195 125.520 ;
        RECT 84.365 125.100 84.535 125.765 ;
        RECT 84.705 125.780 84.895 127.140 ;
        RECT 85.065 126.970 85.340 127.140 ;
        RECT 85.065 126.800 85.345 126.970 ;
        RECT 85.065 125.980 85.340 126.800 ;
        RECT 85.530 126.775 86.060 127.140 ;
        RECT 86.485 126.910 86.815 127.310 ;
        RECT 85.885 126.740 86.060 126.775 ;
        RECT 85.545 125.780 85.715 126.580 ;
        RECT 84.705 125.610 85.715 125.780 ;
        RECT 85.885 126.570 86.815 126.740 ;
        RECT 86.985 126.570 87.240 127.140 ;
        RECT 87.790 126.630 88.045 127.130 ;
        RECT 88.225 126.850 88.510 127.310 ;
        RECT 85.885 125.440 86.055 126.570 ;
        RECT 86.645 126.400 86.815 126.570 ;
        RECT 84.930 125.270 86.055 125.440 ;
        RECT 86.225 126.070 86.420 126.400 ;
        RECT 86.645 126.070 86.900 126.400 ;
        RECT 86.225 125.100 86.395 126.070 ;
        RECT 87.070 125.900 87.240 126.570 ;
        RECT 87.705 126.600 88.045 126.630 ;
        RECT 87.705 126.460 87.970 126.600 ;
        RECT 84.365 124.930 86.395 125.100 ;
        RECT 86.565 124.760 86.735 125.900 ;
        RECT 86.905 124.930 87.240 125.900 ;
        RECT 87.790 125.740 87.970 126.460 ;
        RECT 88.690 126.400 88.940 127.050 ;
        RECT 88.140 126.070 88.940 126.400 ;
        RECT 87.790 125.070 88.045 125.740 ;
        RECT 88.225 124.760 88.510 125.560 ;
        RECT 88.690 125.480 88.940 126.070 ;
        RECT 89.140 126.715 89.460 127.045 ;
        RECT 89.640 126.830 90.300 127.310 ;
        RECT 90.500 126.920 91.350 127.090 ;
        RECT 89.140 125.820 89.330 126.715 ;
        RECT 89.650 126.390 90.310 126.660 ;
        RECT 89.980 126.330 90.310 126.390 ;
        RECT 89.500 126.160 89.830 126.220 ;
        RECT 90.500 126.160 90.670 126.920 ;
        RECT 91.910 126.850 92.230 127.310 ;
        RECT 92.430 126.670 92.680 127.100 ;
        RECT 92.970 126.870 93.380 127.310 ;
        RECT 93.550 126.930 94.565 127.130 ;
        RECT 90.840 126.500 92.090 126.670 ;
        RECT 90.840 126.380 91.170 126.500 ;
        RECT 89.500 125.990 91.400 126.160 ;
        RECT 89.140 125.650 91.060 125.820 ;
        RECT 89.140 125.630 89.460 125.650 ;
        RECT 88.690 124.970 89.020 125.480 ;
        RECT 89.290 125.020 89.460 125.630 ;
        RECT 91.230 125.480 91.400 125.990 ;
        RECT 91.570 125.920 91.750 126.330 ;
        RECT 91.920 125.740 92.090 126.500 ;
        RECT 89.630 124.760 89.960 125.450 ;
        RECT 90.190 125.310 91.400 125.480 ;
        RECT 91.570 125.430 92.090 125.740 ;
        RECT 92.260 126.330 92.680 126.670 ;
        RECT 92.970 126.330 93.380 126.660 ;
        RECT 92.260 125.560 92.450 126.330 ;
        RECT 93.550 126.200 93.720 126.930 ;
        RECT 94.865 126.760 95.035 127.090 ;
        RECT 95.205 126.930 95.535 127.310 ;
        RECT 93.890 126.380 94.240 126.750 ;
        RECT 93.550 126.160 93.970 126.200 ;
        RECT 92.620 125.990 93.970 126.160 ;
        RECT 92.620 125.830 92.870 125.990 ;
        RECT 93.380 125.560 93.630 125.820 ;
        RECT 92.260 125.310 93.630 125.560 ;
        RECT 90.190 125.020 90.430 125.310 ;
        RECT 91.230 125.230 91.400 125.310 ;
        RECT 90.630 124.760 91.050 125.140 ;
        RECT 91.230 124.980 91.860 125.230 ;
        RECT 92.330 124.760 92.660 125.140 ;
        RECT 92.830 125.020 93.000 125.310 ;
        RECT 93.800 125.145 93.970 125.990 ;
        RECT 94.420 125.820 94.640 126.690 ;
        RECT 94.865 126.570 95.560 126.760 ;
        RECT 94.140 125.440 94.640 125.820 ;
        RECT 94.810 125.770 95.220 126.390 ;
        RECT 95.390 125.600 95.560 126.570 ;
        RECT 94.865 125.430 95.560 125.600 ;
        RECT 93.180 124.760 93.560 125.140 ;
        RECT 93.800 124.975 94.630 125.145 ;
        RECT 94.865 124.930 95.035 125.430 ;
        RECT 95.205 124.760 95.535 125.260 ;
        RECT 95.750 124.930 95.975 127.050 ;
        RECT 96.145 126.930 96.475 127.310 ;
        RECT 96.645 126.760 96.815 127.050 ;
        RECT 96.150 126.590 96.815 126.760 ;
        RECT 96.150 125.600 96.380 126.590 ;
        RECT 97.535 126.540 99.205 127.310 ;
        RECT 96.550 125.770 96.900 126.420 ;
        RECT 97.535 125.850 98.285 126.370 ;
        RECT 98.455 126.020 99.205 126.540 ;
        RECT 99.415 126.490 99.645 127.310 ;
        RECT 99.815 126.510 100.145 127.140 ;
        RECT 99.395 126.070 99.725 126.320 ;
        RECT 99.895 125.910 100.145 126.510 ;
        RECT 100.315 126.490 100.525 127.310 ;
        RECT 100.760 126.570 101.015 127.140 ;
        RECT 101.185 126.910 101.515 127.310 ;
        RECT 101.940 126.775 102.470 127.140 ;
        RECT 101.940 126.740 102.115 126.775 ;
        RECT 101.185 126.570 102.115 126.740 ;
        RECT 102.660 126.630 102.935 127.140 ;
        RECT 96.150 125.430 96.815 125.600 ;
        RECT 96.145 124.760 96.475 125.260 ;
        RECT 96.645 124.930 96.815 125.430 ;
        RECT 97.535 124.760 99.205 125.850 ;
        RECT 99.415 124.760 99.645 125.900 ;
        RECT 99.815 124.930 100.145 125.910 ;
        RECT 100.760 125.900 100.930 126.570 ;
        RECT 101.185 126.400 101.355 126.570 ;
        RECT 101.100 126.070 101.355 126.400 ;
        RECT 101.580 126.070 101.775 126.400 ;
        RECT 100.315 124.760 100.525 125.900 ;
        RECT 100.760 124.930 101.095 125.900 ;
        RECT 101.265 124.760 101.435 125.900 ;
        RECT 101.605 125.100 101.775 126.070 ;
        RECT 101.945 125.440 102.115 126.570 ;
        RECT 102.285 125.780 102.455 126.580 ;
        RECT 102.655 126.460 102.935 126.630 ;
        RECT 102.660 125.980 102.935 126.460 ;
        RECT 103.105 125.780 103.295 127.140 ;
        RECT 103.475 126.775 103.985 127.310 ;
        RECT 104.205 126.500 104.450 127.105 ;
        RECT 105.355 126.585 105.645 127.310 ;
        RECT 106.190 126.970 106.445 127.130 ;
        RECT 106.105 126.800 106.445 126.970 ;
        RECT 106.625 126.850 106.910 127.310 ;
        RECT 106.190 126.600 106.445 126.800 ;
        RECT 103.495 126.330 104.725 126.500 ;
        RECT 102.285 125.610 103.295 125.780 ;
        RECT 103.465 125.765 104.215 125.955 ;
        RECT 101.945 125.270 103.070 125.440 ;
        RECT 103.465 125.100 103.635 125.765 ;
        RECT 104.385 125.520 104.725 126.330 ;
        RECT 101.605 124.930 103.635 125.100 ;
        RECT 103.805 124.760 103.975 125.520 ;
        RECT 104.210 125.110 104.725 125.520 ;
        RECT 105.355 124.760 105.645 125.925 ;
        RECT 106.190 125.740 106.370 126.600 ;
        RECT 107.090 126.400 107.340 127.050 ;
        RECT 106.540 126.070 107.340 126.400 ;
        RECT 106.190 125.070 106.445 125.740 ;
        RECT 106.625 124.760 106.910 125.560 ;
        RECT 107.090 125.480 107.340 126.070 ;
        RECT 107.540 126.715 107.860 127.045 ;
        RECT 108.040 126.830 108.700 127.310 ;
        RECT 108.900 126.920 109.750 127.090 ;
        RECT 107.540 125.820 107.730 126.715 ;
        RECT 108.050 126.390 108.710 126.660 ;
        RECT 108.380 126.330 108.710 126.390 ;
        RECT 107.900 126.160 108.230 126.220 ;
        RECT 108.900 126.160 109.070 126.920 ;
        RECT 110.310 126.850 110.630 127.310 ;
        RECT 110.830 126.670 111.080 127.100 ;
        RECT 111.370 126.870 111.780 127.310 ;
        RECT 111.950 126.930 112.965 127.130 ;
        RECT 109.240 126.500 110.490 126.670 ;
        RECT 109.240 126.380 109.570 126.500 ;
        RECT 107.900 125.990 109.800 126.160 ;
        RECT 107.540 125.650 109.460 125.820 ;
        RECT 107.540 125.630 107.860 125.650 ;
        RECT 107.090 124.970 107.420 125.480 ;
        RECT 107.690 125.020 107.860 125.630 ;
        RECT 109.630 125.480 109.800 125.990 ;
        RECT 109.970 125.920 110.150 126.330 ;
        RECT 110.320 125.740 110.490 126.500 ;
        RECT 108.030 124.760 108.360 125.450 ;
        RECT 108.590 125.310 109.800 125.480 ;
        RECT 109.970 125.430 110.490 125.740 ;
        RECT 110.660 126.330 111.080 126.670 ;
        RECT 111.370 126.330 111.780 126.660 ;
        RECT 110.660 125.560 110.850 126.330 ;
        RECT 111.950 126.200 112.120 126.930 ;
        RECT 113.265 126.760 113.435 127.090 ;
        RECT 113.605 126.930 113.935 127.310 ;
        RECT 112.290 126.380 112.640 126.750 ;
        RECT 111.950 126.160 112.370 126.200 ;
        RECT 111.020 125.990 112.370 126.160 ;
        RECT 111.020 125.830 111.270 125.990 ;
        RECT 111.780 125.560 112.030 125.820 ;
        RECT 110.660 125.310 112.030 125.560 ;
        RECT 108.590 125.020 108.830 125.310 ;
        RECT 109.630 125.230 109.800 125.310 ;
        RECT 109.030 124.760 109.450 125.140 ;
        RECT 109.630 124.980 110.260 125.230 ;
        RECT 110.730 124.760 111.060 125.140 ;
        RECT 111.230 125.020 111.400 125.310 ;
        RECT 112.200 125.145 112.370 125.990 ;
        RECT 112.820 125.820 113.040 126.690 ;
        RECT 113.265 126.570 113.960 126.760 ;
        RECT 112.540 125.440 113.040 125.820 ;
        RECT 113.210 125.770 113.620 126.390 ;
        RECT 113.790 125.600 113.960 126.570 ;
        RECT 113.265 125.430 113.960 125.600 ;
        RECT 111.580 124.760 111.960 125.140 ;
        RECT 112.200 124.975 113.030 125.145 ;
        RECT 113.265 124.930 113.435 125.430 ;
        RECT 113.605 124.760 113.935 125.260 ;
        RECT 114.150 124.930 114.375 127.050 ;
        RECT 114.545 126.930 114.875 127.310 ;
        RECT 115.045 126.760 115.215 127.050 ;
        RECT 114.550 126.590 115.215 126.760 ;
        RECT 114.550 125.600 114.780 126.590 ;
        RECT 115.475 126.540 117.145 127.310 ;
        RECT 117.315 126.560 118.525 127.310 ;
        RECT 114.950 125.770 115.300 126.420 ;
        RECT 115.475 125.850 116.225 126.370 ;
        RECT 116.395 126.020 117.145 126.540 ;
        RECT 117.315 125.850 117.835 126.390 ;
        RECT 118.005 126.020 118.525 126.560 ;
        RECT 114.550 125.430 115.215 125.600 ;
        RECT 114.545 124.760 114.875 125.260 ;
        RECT 115.045 124.930 115.215 125.430 ;
        RECT 115.475 124.760 117.145 125.850 ;
        RECT 117.315 124.760 118.525 125.850 ;
        RECT 11.430 124.590 118.610 124.760 ;
        RECT 11.515 123.500 12.725 124.590 ;
        RECT 11.515 122.790 12.035 123.330 ;
        RECT 12.205 122.960 12.725 123.500 ;
        RECT 13.875 123.450 14.085 124.590 ;
        RECT 14.255 123.440 14.585 124.420 ;
        RECT 14.755 123.450 14.985 124.590 ;
        RECT 11.515 122.040 12.725 122.790 ;
        RECT 13.875 122.040 14.085 122.860 ;
        RECT 14.255 122.840 14.505 123.440 ;
        RECT 15.195 123.425 15.485 124.590 ;
        RECT 16.030 124.250 16.285 124.280 ;
        RECT 15.945 124.080 16.285 124.250 ;
        RECT 16.030 123.610 16.285 124.080 ;
        RECT 16.465 123.790 16.750 124.590 ;
        RECT 16.930 123.870 17.260 124.380 ;
        RECT 14.675 123.030 15.005 123.280 ;
        RECT 14.255 122.210 14.585 122.840 ;
        RECT 14.755 122.040 14.985 122.860 ;
        RECT 15.195 122.040 15.485 122.765 ;
        RECT 16.030 122.750 16.210 123.610 ;
        RECT 16.930 123.280 17.180 123.870 ;
        RECT 17.530 123.720 17.700 124.330 ;
        RECT 17.870 123.900 18.200 124.590 ;
        RECT 18.430 124.040 18.670 124.330 ;
        RECT 18.870 124.210 19.290 124.590 ;
        RECT 19.470 124.120 20.100 124.370 ;
        RECT 20.570 124.210 20.900 124.590 ;
        RECT 19.470 124.040 19.640 124.120 ;
        RECT 21.070 124.040 21.240 124.330 ;
        RECT 21.420 124.210 21.800 124.590 ;
        RECT 22.040 124.205 22.870 124.375 ;
        RECT 18.430 123.870 19.640 124.040 ;
        RECT 16.380 122.950 17.180 123.280 ;
        RECT 16.030 122.220 16.285 122.750 ;
        RECT 16.465 122.040 16.750 122.500 ;
        RECT 16.930 122.300 17.180 122.950 ;
        RECT 17.380 123.700 17.700 123.720 ;
        RECT 17.380 123.530 19.300 123.700 ;
        RECT 17.380 122.635 17.570 123.530 ;
        RECT 19.470 123.360 19.640 123.870 ;
        RECT 19.810 123.610 20.330 123.920 ;
        RECT 17.740 123.190 19.640 123.360 ;
        RECT 17.740 123.130 18.070 123.190 ;
        RECT 18.220 122.960 18.550 123.020 ;
        RECT 17.890 122.690 18.550 122.960 ;
        RECT 17.380 122.305 17.700 122.635 ;
        RECT 17.880 122.040 18.540 122.520 ;
        RECT 18.740 122.430 18.910 123.190 ;
        RECT 19.810 123.020 19.990 123.430 ;
        RECT 19.080 122.850 19.410 122.970 ;
        RECT 20.160 122.850 20.330 123.610 ;
        RECT 19.080 122.680 20.330 122.850 ;
        RECT 20.500 123.790 21.870 124.040 ;
        RECT 20.500 123.020 20.690 123.790 ;
        RECT 21.620 123.530 21.870 123.790 ;
        RECT 20.860 123.360 21.110 123.520 ;
        RECT 22.040 123.360 22.210 124.205 ;
        RECT 23.105 123.920 23.275 124.420 ;
        RECT 23.445 124.090 23.775 124.590 ;
        RECT 22.380 123.530 22.880 123.910 ;
        RECT 23.105 123.750 23.800 123.920 ;
        RECT 20.860 123.190 22.210 123.360 ;
        RECT 21.790 123.150 22.210 123.190 ;
        RECT 20.500 122.680 20.920 123.020 ;
        RECT 21.210 122.690 21.620 123.020 ;
        RECT 18.740 122.260 19.590 122.430 ;
        RECT 20.150 122.040 20.470 122.500 ;
        RECT 20.670 122.250 20.920 122.680 ;
        RECT 21.210 122.040 21.620 122.480 ;
        RECT 21.790 122.420 21.960 123.150 ;
        RECT 22.130 122.600 22.480 122.970 ;
        RECT 22.660 122.660 22.880 123.530 ;
        RECT 23.050 122.960 23.460 123.580 ;
        RECT 23.630 122.780 23.800 123.750 ;
        RECT 23.105 122.590 23.800 122.780 ;
        RECT 21.790 122.220 22.805 122.420 ;
        RECT 23.105 122.260 23.275 122.590 ;
        RECT 23.445 122.040 23.775 122.420 ;
        RECT 23.990 122.300 24.215 124.420 ;
        RECT 24.385 124.090 24.715 124.590 ;
        RECT 24.885 123.920 25.055 124.420 ;
        RECT 25.690 124.250 25.945 124.280 ;
        RECT 25.605 124.080 25.945 124.250 ;
        RECT 24.390 123.750 25.055 123.920 ;
        RECT 24.390 122.760 24.620 123.750 ;
        RECT 25.690 123.610 25.945 124.080 ;
        RECT 26.125 123.790 26.410 124.590 ;
        RECT 26.590 123.870 26.920 124.380 ;
        RECT 24.790 122.930 25.140 123.580 ;
        RECT 24.390 122.590 25.055 122.760 ;
        RECT 24.385 122.040 24.715 122.420 ;
        RECT 24.885 122.300 25.055 122.590 ;
        RECT 25.690 122.750 25.870 123.610 ;
        RECT 26.590 123.280 26.840 123.870 ;
        RECT 27.190 123.720 27.360 124.330 ;
        RECT 27.530 123.900 27.860 124.590 ;
        RECT 28.090 124.040 28.330 124.330 ;
        RECT 28.530 124.210 28.950 124.590 ;
        RECT 29.130 124.120 29.760 124.370 ;
        RECT 30.230 124.210 30.560 124.590 ;
        RECT 29.130 124.040 29.300 124.120 ;
        RECT 30.730 124.040 30.900 124.330 ;
        RECT 31.080 124.210 31.460 124.590 ;
        RECT 31.700 124.205 32.530 124.375 ;
        RECT 28.090 123.870 29.300 124.040 ;
        RECT 26.040 122.950 26.840 123.280 ;
        RECT 25.690 122.220 25.945 122.750 ;
        RECT 26.125 122.040 26.410 122.500 ;
        RECT 26.590 122.300 26.840 122.950 ;
        RECT 27.040 123.700 27.360 123.720 ;
        RECT 27.040 123.530 28.960 123.700 ;
        RECT 27.040 122.635 27.230 123.530 ;
        RECT 29.130 123.360 29.300 123.870 ;
        RECT 29.470 123.610 29.990 123.920 ;
        RECT 27.400 123.190 29.300 123.360 ;
        RECT 27.400 123.130 27.730 123.190 ;
        RECT 27.880 122.960 28.210 123.020 ;
        RECT 27.550 122.690 28.210 122.960 ;
        RECT 27.040 122.305 27.360 122.635 ;
        RECT 27.540 122.040 28.200 122.520 ;
        RECT 28.400 122.430 28.570 123.190 ;
        RECT 29.470 123.020 29.650 123.430 ;
        RECT 28.740 122.850 29.070 122.970 ;
        RECT 29.820 122.850 29.990 123.610 ;
        RECT 28.740 122.680 29.990 122.850 ;
        RECT 30.160 123.790 31.530 124.040 ;
        RECT 30.160 123.020 30.350 123.790 ;
        RECT 31.280 123.530 31.530 123.790 ;
        RECT 30.520 123.360 30.770 123.520 ;
        RECT 31.700 123.360 31.870 124.205 ;
        RECT 32.765 123.920 32.935 124.420 ;
        RECT 33.105 124.090 33.435 124.590 ;
        RECT 32.040 123.530 32.540 123.910 ;
        RECT 32.765 123.750 33.460 123.920 ;
        RECT 30.520 123.190 31.870 123.360 ;
        RECT 31.450 123.150 31.870 123.190 ;
        RECT 30.160 122.680 30.580 123.020 ;
        RECT 30.870 122.690 31.280 123.020 ;
        RECT 28.400 122.260 29.250 122.430 ;
        RECT 29.810 122.040 30.130 122.500 ;
        RECT 30.330 122.250 30.580 122.680 ;
        RECT 30.870 122.040 31.280 122.480 ;
        RECT 31.450 122.420 31.620 123.150 ;
        RECT 31.790 122.600 32.140 122.970 ;
        RECT 32.320 122.660 32.540 123.530 ;
        RECT 32.710 122.960 33.120 123.580 ;
        RECT 33.290 122.780 33.460 123.750 ;
        RECT 32.765 122.590 33.460 122.780 ;
        RECT 31.450 122.220 32.465 122.420 ;
        RECT 32.765 122.260 32.935 122.590 ;
        RECT 33.105 122.040 33.435 122.420 ;
        RECT 33.650 122.300 33.875 124.420 ;
        RECT 34.045 124.090 34.375 124.590 ;
        RECT 34.545 123.920 34.715 124.420 ;
        RECT 34.050 123.750 34.715 123.920 ;
        RECT 34.050 122.760 34.280 123.750 ;
        RECT 34.450 122.930 34.800 123.580 ;
        RECT 35.435 123.500 37.105 124.590 ;
        RECT 35.435 122.980 36.185 123.500 ;
        RECT 37.315 123.450 37.545 124.590 ;
        RECT 37.715 123.440 38.045 124.420 ;
        RECT 38.215 123.450 38.425 124.590 ;
        RECT 39.115 123.500 40.785 124.590 ;
        RECT 36.355 122.810 37.105 123.330 ;
        RECT 37.295 123.030 37.625 123.280 ;
        RECT 34.050 122.590 34.715 122.760 ;
        RECT 34.045 122.040 34.375 122.420 ;
        RECT 34.545 122.300 34.715 122.590 ;
        RECT 35.435 122.040 37.105 122.810 ;
        RECT 37.315 122.040 37.545 122.860 ;
        RECT 37.795 122.840 38.045 123.440 ;
        RECT 39.115 122.980 39.865 123.500 ;
        RECT 40.955 123.425 41.245 124.590 ;
        RECT 41.505 123.660 41.675 124.420 ;
        RECT 41.855 123.830 42.185 124.590 ;
        RECT 41.505 123.490 42.170 123.660 ;
        RECT 42.355 123.515 42.625 124.420 ;
        RECT 42.000 123.345 42.170 123.490 ;
        RECT 37.715 122.210 38.045 122.840 ;
        RECT 38.215 122.040 38.425 122.860 ;
        RECT 40.035 122.810 40.785 123.330 ;
        RECT 41.435 122.940 41.765 123.310 ;
        RECT 42.000 123.015 42.285 123.345 ;
        RECT 39.115 122.040 40.785 122.810 ;
        RECT 40.955 122.040 41.245 122.765 ;
        RECT 42.000 122.760 42.170 123.015 ;
        RECT 41.505 122.590 42.170 122.760 ;
        RECT 42.455 122.715 42.625 123.515 ;
        RECT 42.835 123.450 43.065 124.590 ;
        RECT 43.235 123.440 43.565 124.420 ;
        RECT 43.735 123.450 43.945 124.590 ;
        RECT 44.265 123.845 44.535 124.590 ;
        RECT 45.165 124.585 51.440 124.590 ;
        RECT 44.705 123.675 44.995 124.415 ;
        RECT 45.165 123.860 45.420 124.585 ;
        RECT 45.605 123.690 45.865 124.415 ;
        RECT 46.035 123.860 46.280 124.585 ;
        RECT 46.465 123.690 46.725 124.415 ;
        RECT 46.895 123.860 47.140 124.585 ;
        RECT 47.325 123.690 47.585 124.415 ;
        RECT 47.755 123.860 48.000 124.585 ;
        RECT 48.170 123.690 48.430 124.415 ;
        RECT 48.600 123.860 48.860 124.585 ;
        RECT 49.030 123.690 49.290 124.415 ;
        RECT 49.460 123.860 49.720 124.585 ;
        RECT 49.890 123.690 50.150 124.415 ;
        RECT 50.320 123.860 50.580 124.585 ;
        RECT 50.750 123.690 51.010 124.415 ;
        RECT 51.180 123.790 51.440 124.585 ;
        RECT 45.605 123.675 51.010 123.690 ;
        RECT 44.265 123.450 51.010 123.675 ;
        RECT 42.815 123.030 43.145 123.280 ;
        RECT 41.505 122.210 41.675 122.590 ;
        RECT 41.855 122.040 42.185 122.420 ;
        RECT 42.365 122.210 42.625 122.715 ;
        RECT 42.835 122.040 43.065 122.860 ;
        RECT 43.315 122.840 43.565 123.440 ;
        RECT 44.265 122.860 45.430 123.450 ;
        RECT 51.610 123.280 51.860 124.415 ;
        RECT 52.040 123.780 52.300 124.590 ;
        RECT 52.475 123.280 52.720 124.420 ;
        RECT 52.900 123.780 53.195 124.590 ;
        RECT 53.750 124.250 54.005 124.280 ;
        RECT 53.665 124.080 54.005 124.250 ;
        RECT 53.750 123.610 54.005 124.080 ;
        RECT 54.185 123.790 54.470 124.590 ;
        RECT 54.650 123.870 54.980 124.380 ;
        RECT 45.600 123.030 52.720 123.280 ;
        RECT 43.235 122.210 43.565 122.840 ;
        RECT 43.735 122.040 43.945 122.860 ;
        RECT 44.265 122.690 51.010 122.860 ;
        RECT 44.265 122.040 44.565 122.520 ;
        RECT 44.735 122.235 44.995 122.690 ;
        RECT 45.165 122.040 45.425 122.520 ;
        RECT 45.605 122.235 45.865 122.690 ;
        RECT 46.035 122.040 46.285 122.520 ;
        RECT 46.465 122.235 46.725 122.690 ;
        RECT 46.895 122.040 47.145 122.520 ;
        RECT 47.325 122.235 47.585 122.690 ;
        RECT 47.755 122.040 48.000 122.520 ;
        RECT 48.170 122.235 48.445 122.690 ;
        RECT 48.615 122.040 48.860 122.520 ;
        RECT 49.030 122.235 49.290 122.690 ;
        RECT 49.460 122.040 49.720 122.520 ;
        RECT 49.890 122.235 50.150 122.690 ;
        RECT 50.320 122.040 50.580 122.520 ;
        RECT 50.750 122.235 51.010 122.690 ;
        RECT 51.180 122.040 51.440 122.600 ;
        RECT 51.610 122.220 51.860 123.030 ;
        RECT 52.040 122.040 52.300 122.565 ;
        RECT 52.470 122.220 52.720 123.030 ;
        RECT 52.890 122.720 53.205 123.280 ;
        RECT 53.750 122.750 53.930 123.610 ;
        RECT 54.650 123.280 54.900 123.870 ;
        RECT 55.250 123.720 55.420 124.330 ;
        RECT 55.590 123.900 55.920 124.590 ;
        RECT 56.150 124.040 56.390 124.330 ;
        RECT 56.590 124.210 57.010 124.590 ;
        RECT 57.190 124.120 57.820 124.370 ;
        RECT 58.290 124.210 58.620 124.590 ;
        RECT 57.190 124.040 57.360 124.120 ;
        RECT 58.790 124.040 58.960 124.330 ;
        RECT 59.140 124.210 59.520 124.590 ;
        RECT 59.760 124.205 60.590 124.375 ;
        RECT 56.150 123.870 57.360 124.040 ;
        RECT 54.100 122.950 54.900 123.280 ;
        RECT 52.900 122.040 53.205 122.550 ;
        RECT 53.750 122.220 54.005 122.750 ;
        RECT 54.185 122.040 54.470 122.500 ;
        RECT 54.650 122.300 54.900 122.950 ;
        RECT 55.100 123.700 55.420 123.720 ;
        RECT 55.100 123.530 57.020 123.700 ;
        RECT 55.100 122.635 55.290 123.530 ;
        RECT 57.190 123.360 57.360 123.870 ;
        RECT 57.530 123.610 58.050 123.920 ;
        RECT 55.460 123.190 57.360 123.360 ;
        RECT 55.460 123.130 55.790 123.190 ;
        RECT 55.940 122.960 56.270 123.020 ;
        RECT 55.610 122.690 56.270 122.960 ;
        RECT 55.100 122.305 55.420 122.635 ;
        RECT 55.600 122.040 56.260 122.520 ;
        RECT 56.460 122.430 56.630 123.190 ;
        RECT 57.530 123.020 57.710 123.430 ;
        RECT 56.800 122.850 57.130 122.970 ;
        RECT 57.880 122.850 58.050 123.610 ;
        RECT 56.800 122.680 58.050 122.850 ;
        RECT 58.220 123.790 59.590 124.040 ;
        RECT 58.220 123.020 58.410 123.790 ;
        RECT 59.340 123.530 59.590 123.790 ;
        RECT 58.580 123.360 58.830 123.520 ;
        RECT 59.760 123.360 59.930 124.205 ;
        RECT 60.825 123.920 60.995 124.420 ;
        RECT 61.165 124.090 61.495 124.590 ;
        RECT 60.100 123.530 60.600 123.910 ;
        RECT 60.825 123.750 61.520 123.920 ;
        RECT 58.580 123.190 59.930 123.360 ;
        RECT 59.510 123.150 59.930 123.190 ;
        RECT 58.220 122.680 58.640 123.020 ;
        RECT 58.930 122.690 59.340 123.020 ;
        RECT 56.460 122.260 57.310 122.430 ;
        RECT 57.870 122.040 58.190 122.500 ;
        RECT 58.390 122.250 58.640 122.680 ;
        RECT 58.930 122.040 59.340 122.480 ;
        RECT 59.510 122.420 59.680 123.150 ;
        RECT 59.850 122.600 60.200 122.970 ;
        RECT 60.380 122.660 60.600 123.530 ;
        RECT 60.770 122.960 61.180 123.580 ;
        RECT 61.350 122.780 61.520 123.750 ;
        RECT 60.825 122.590 61.520 122.780 ;
        RECT 59.510 122.220 60.525 122.420 ;
        RECT 60.825 122.260 60.995 122.590 ;
        RECT 61.165 122.040 61.495 122.420 ;
        RECT 61.710 122.300 61.935 124.420 ;
        RECT 62.105 124.090 62.435 124.590 ;
        RECT 62.605 123.920 62.775 124.420 ;
        RECT 62.110 123.750 62.775 123.920 ;
        RECT 62.110 122.760 62.340 123.750 ;
        RECT 62.510 122.930 62.860 123.580 ;
        RECT 63.035 123.500 66.545 124.590 ;
        RECT 63.035 122.980 64.725 123.500 ;
        RECT 66.715 123.425 67.005 124.590 ;
        RECT 67.635 123.500 70.225 124.590 ;
        RECT 64.895 122.810 66.545 123.330 ;
        RECT 67.635 122.980 68.845 123.500 ;
        RECT 70.455 123.450 70.665 124.590 ;
        RECT 70.835 123.440 71.165 124.420 ;
        RECT 71.335 123.450 71.565 124.590 ;
        RECT 72.610 124.250 72.865 124.280 ;
        RECT 72.525 124.080 72.865 124.250 ;
        RECT 72.610 123.610 72.865 124.080 ;
        RECT 73.045 123.790 73.330 124.590 ;
        RECT 73.510 123.870 73.840 124.380 ;
        RECT 69.015 122.810 70.225 123.330 ;
        RECT 62.110 122.590 62.775 122.760 ;
        RECT 62.105 122.040 62.435 122.420 ;
        RECT 62.605 122.300 62.775 122.590 ;
        RECT 63.035 122.040 66.545 122.810 ;
        RECT 66.715 122.040 67.005 122.765 ;
        RECT 67.635 122.040 70.225 122.810 ;
        RECT 70.455 122.040 70.665 122.860 ;
        RECT 70.835 122.840 71.085 123.440 ;
        RECT 71.255 123.030 71.585 123.280 ;
        RECT 70.835 122.210 71.165 122.840 ;
        RECT 71.335 122.040 71.565 122.860 ;
        RECT 72.610 122.750 72.790 123.610 ;
        RECT 73.510 123.280 73.760 123.870 ;
        RECT 74.110 123.720 74.280 124.330 ;
        RECT 74.450 123.900 74.780 124.590 ;
        RECT 75.010 124.040 75.250 124.330 ;
        RECT 75.450 124.210 75.870 124.590 ;
        RECT 76.050 124.120 76.680 124.370 ;
        RECT 77.150 124.210 77.480 124.590 ;
        RECT 76.050 124.040 76.220 124.120 ;
        RECT 77.650 124.040 77.820 124.330 ;
        RECT 78.000 124.210 78.380 124.590 ;
        RECT 78.620 124.205 79.450 124.375 ;
        RECT 75.010 123.870 76.220 124.040 ;
        RECT 72.960 122.950 73.760 123.280 ;
        RECT 72.610 122.220 72.865 122.750 ;
        RECT 73.045 122.040 73.330 122.500 ;
        RECT 73.510 122.300 73.760 122.950 ;
        RECT 73.960 123.700 74.280 123.720 ;
        RECT 73.960 123.530 75.880 123.700 ;
        RECT 73.960 122.635 74.150 123.530 ;
        RECT 76.050 123.360 76.220 123.870 ;
        RECT 76.390 123.610 76.910 123.920 ;
        RECT 74.320 123.190 76.220 123.360 ;
        RECT 74.320 123.130 74.650 123.190 ;
        RECT 74.800 122.960 75.130 123.020 ;
        RECT 74.470 122.690 75.130 122.960 ;
        RECT 73.960 122.305 74.280 122.635 ;
        RECT 74.460 122.040 75.120 122.520 ;
        RECT 75.320 122.430 75.490 123.190 ;
        RECT 76.390 123.020 76.570 123.430 ;
        RECT 75.660 122.850 75.990 122.970 ;
        RECT 76.740 122.850 76.910 123.610 ;
        RECT 75.660 122.680 76.910 122.850 ;
        RECT 77.080 123.790 78.450 124.040 ;
        RECT 77.080 123.020 77.270 123.790 ;
        RECT 78.200 123.530 78.450 123.790 ;
        RECT 77.440 123.360 77.690 123.520 ;
        RECT 78.620 123.360 78.790 124.205 ;
        RECT 79.685 123.920 79.855 124.420 ;
        RECT 80.025 124.090 80.355 124.590 ;
        RECT 78.960 123.530 79.460 123.910 ;
        RECT 79.685 123.750 80.380 123.920 ;
        RECT 77.440 123.190 78.790 123.360 ;
        RECT 78.370 123.150 78.790 123.190 ;
        RECT 77.080 122.680 77.500 123.020 ;
        RECT 77.790 122.690 78.200 123.020 ;
        RECT 75.320 122.260 76.170 122.430 ;
        RECT 76.730 122.040 77.050 122.500 ;
        RECT 77.250 122.250 77.500 122.680 ;
        RECT 77.790 122.040 78.200 122.480 ;
        RECT 78.370 122.420 78.540 123.150 ;
        RECT 78.710 122.600 79.060 122.970 ;
        RECT 79.240 122.660 79.460 123.530 ;
        RECT 79.630 122.960 80.040 123.580 ;
        RECT 80.210 122.780 80.380 123.750 ;
        RECT 79.685 122.590 80.380 122.780 ;
        RECT 78.370 122.220 79.385 122.420 ;
        RECT 79.685 122.260 79.855 122.590 ;
        RECT 80.025 122.040 80.355 122.420 ;
        RECT 80.570 122.300 80.795 124.420 ;
        RECT 80.965 124.090 81.295 124.590 ;
        RECT 81.465 123.920 81.635 124.420 ;
        RECT 82.270 124.250 82.525 124.280 ;
        RECT 82.185 124.080 82.525 124.250 ;
        RECT 80.970 123.750 81.635 123.920 ;
        RECT 80.970 122.760 81.200 123.750 ;
        RECT 82.270 123.610 82.525 124.080 ;
        RECT 82.705 123.790 82.990 124.590 ;
        RECT 83.170 123.870 83.500 124.380 ;
        RECT 81.370 122.930 81.720 123.580 ;
        RECT 80.970 122.590 81.635 122.760 ;
        RECT 80.965 122.040 81.295 122.420 ;
        RECT 81.465 122.300 81.635 122.590 ;
        RECT 82.270 122.750 82.450 123.610 ;
        RECT 83.170 123.280 83.420 123.870 ;
        RECT 83.770 123.720 83.940 124.330 ;
        RECT 84.110 123.900 84.440 124.590 ;
        RECT 84.670 124.040 84.910 124.330 ;
        RECT 85.110 124.210 85.530 124.590 ;
        RECT 85.710 124.120 86.340 124.370 ;
        RECT 86.810 124.210 87.140 124.590 ;
        RECT 85.710 124.040 85.880 124.120 ;
        RECT 87.310 124.040 87.480 124.330 ;
        RECT 87.660 124.210 88.040 124.590 ;
        RECT 88.280 124.205 89.110 124.375 ;
        RECT 84.670 123.870 85.880 124.040 ;
        RECT 82.620 122.950 83.420 123.280 ;
        RECT 82.270 122.220 82.525 122.750 ;
        RECT 82.705 122.040 82.990 122.500 ;
        RECT 83.170 122.300 83.420 122.950 ;
        RECT 83.620 123.700 83.940 123.720 ;
        RECT 83.620 123.530 85.540 123.700 ;
        RECT 83.620 122.635 83.810 123.530 ;
        RECT 85.710 123.360 85.880 123.870 ;
        RECT 86.050 123.610 86.570 123.920 ;
        RECT 83.980 123.190 85.880 123.360 ;
        RECT 83.980 123.130 84.310 123.190 ;
        RECT 84.460 122.960 84.790 123.020 ;
        RECT 84.130 122.690 84.790 122.960 ;
        RECT 83.620 122.305 83.940 122.635 ;
        RECT 84.120 122.040 84.780 122.520 ;
        RECT 84.980 122.430 85.150 123.190 ;
        RECT 86.050 123.020 86.230 123.430 ;
        RECT 85.320 122.850 85.650 122.970 ;
        RECT 86.400 122.850 86.570 123.610 ;
        RECT 85.320 122.680 86.570 122.850 ;
        RECT 86.740 123.790 88.110 124.040 ;
        RECT 86.740 123.020 86.930 123.790 ;
        RECT 87.860 123.530 88.110 123.790 ;
        RECT 87.100 123.360 87.350 123.520 ;
        RECT 88.280 123.360 88.450 124.205 ;
        RECT 89.345 123.920 89.515 124.420 ;
        RECT 89.685 124.090 90.015 124.590 ;
        RECT 88.620 123.530 89.120 123.910 ;
        RECT 89.345 123.750 90.040 123.920 ;
        RECT 87.100 123.190 88.450 123.360 ;
        RECT 88.030 123.150 88.450 123.190 ;
        RECT 86.740 122.680 87.160 123.020 ;
        RECT 87.450 122.690 87.860 123.020 ;
        RECT 84.980 122.260 85.830 122.430 ;
        RECT 86.390 122.040 86.710 122.500 ;
        RECT 86.910 122.250 87.160 122.680 ;
        RECT 87.450 122.040 87.860 122.480 ;
        RECT 88.030 122.420 88.200 123.150 ;
        RECT 88.370 122.600 88.720 122.970 ;
        RECT 88.900 122.660 89.120 123.530 ;
        RECT 89.290 122.960 89.700 123.580 ;
        RECT 89.870 122.780 90.040 123.750 ;
        RECT 89.345 122.590 90.040 122.780 ;
        RECT 88.030 122.220 89.045 122.420 ;
        RECT 89.345 122.260 89.515 122.590 ;
        RECT 89.685 122.040 90.015 122.420 ;
        RECT 90.230 122.300 90.455 124.420 ;
        RECT 90.625 124.090 90.955 124.590 ;
        RECT 91.125 123.920 91.295 124.420 ;
        RECT 90.630 123.750 91.295 123.920 ;
        RECT 90.630 122.760 90.860 123.750 ;
        RECT 91.030 122.930 91.380 123.580 ;
        RECT 92.475 123.425 92.765 124.590 ;
        RECT 93.395 123.500 95.065 124.590 ;
        RECT 95.235 123.515 95.505 124.420 ;
        RECT 95.675 123.830 96.005 124.590 ;
        RECT 96.185 123.660 96.355 124.420 ;
        RECT 96.990 124.250 97.245 124.280 ;
        RECT 96.905 124.080 97.245 124.250 ;
        RECT 93.395 122.980 94.145 123.500 ;
        RECT 94.315 122.810 95.065 123.330 ;
        RECT 90.630 122.590 91.295 122.760 ;
        RECT 90.625 122.040 90.955 122.420 ;
        RECT 91.125 122.300 91.295 122.590 ;
        RECT 92.475 122.040 92.765 122.765 ;
        RECT 93.395 122.040 95.065 122.810 ;
        RECT 95.235 122.715 95.405 123.515 ;
        RECT 95.690 123.490 96.355 123.660 ;
        RECT 96.990 123.610 97.245 124.080 ;
        RECT 97.425 123.790 97.710 124.590 ;
        RECT 97.890 123.870 98.220 124.380 ;
        RECT 95.690 123.345 95.860 123.490 ;
        RECT 95.575 123.015 95.860 123.345 ;
        RECT 95.690 122.760 95.860 123.015 ;
        RECT 96.095 122.940 96.425 123.310 ;
        RECT 95.235 122.210 95.495 122.715 ;
        RECT 95.690 122.590 96.355 122.760 ;
        RECT 95.675 122.040 96.005 122.420 ;
        RECT 96.185 122.210 96.355 122.590 ;
        RECT 96.990 122.750 97.170 123.610 ;
        RECT 97.890 123.280 98.140 123.870 ;
        RECT 98.490 123.720 98.660 124.330 ;
        RECT 98.830 123.900 99.160 124.590 ;
        RECT 99.390 124.040 99.630 124.330 ;
        RECT 99.830 124.210 100.250 124.590 ;
        RECT 100.430 124.120 101.060 124.370 ;
        RECT 101.530 124.210 101.860 124.590 ;
        RECT 100.430 124.040 100.600 124.120 ;
        RECT 102.030 124.040 102.200 124.330 ;
        RECT 102.380 124.210 102.760 124.590 ;
        RECT 103.000 124.205 103.830 124.375 ;
        RECT 99.390 123.870 100.600 124.040 ;
        RECT 97.340 122.950 98.140 123.280 ;
        RECT 96.990 122.220 97.245 122.750 ;
        RECT 97.425 122.040 97.710 122.500 ;
        RECT 97.890 122.300 98.140 122.950 ;
        RECT 98.340 123.700 98.660 123.720 ;
        RECT 98.340 123.530 100.260 123.700 ;
        RECT 98.340 122.635 98.530 123.530 ;
        RECT 100.430 123.360 100.600 123.870 ;
        RECT 100.770 123.610 101.290 123.920 ;
        RECT 98.700 123.190 100.600 123.360 ;
        RECT 98.700 123.130 99.030 123.190 ;
        RECT 99.180 122.960 99.510 123.020 ;
        RECT 98.850 122.690 99.510 122.960 ;
        RECT 98.340 122.305 98.660 122.635 ;
        RECT 98.840 122.040 99.500 122.520 ;
        RECT 99.700 122.430 99.870 123.190 ;
        RECT 100.770 123.020 100.950 123.430 ;
        RECT 100.040 122.850 100.370 122.970 ;
        RECT 101.120 122.850 101.290 123.610 ;
        RECT 100.040 122.680 101.290 122.850 ;
        RECT 101.460 123.790 102.830 124.040 ;
        RECT 101.460 123.020 101.650 123.790 ;
        RECT 102.580 123.530 102.830 123.790 ;
        RECT 101.820 123.360 102.070 123.520 ;
        RECT 103.000 123.360 103.170 124.205 ;
        RECT 104.065 123.920 104.235 124.420 ;
        RECT 104.405 124.090 104.735 124.590 ;
        RECT 103.340 123.530 103.840 123.910 ;
        RECT 104.065 123.750 104.760 123.920 ;
        RECT 101.820 123.190 103.170 123.360 ;
        RECT 102.750 123.150 103.170 123.190 ;
        RECT 101.460 122.680 101.880 123.020 ;
        RECT 102.170 122.690 102.580 123.020 ;
        RECT 99.700 122.260 100.550 122.430 ;
        RECT 101.110 122.040 101.430 122.500 ;
        RECT 101.630 122.250 101.880 122.680 ;
        RECT 102.170 122.040 102.580 122.480 ;
        RECT 102.750 122.420 102.920 123.150 ;
        RECT 103.090 122.600 103.440 122.970 ;
        RECT 103.620 122.660 103.840 123.530 ;
        RECT 104.010 122.960 104.420 123.580 ;
        RECT 104.590 122.780 104.760 123.750 ;
        RECT 104.065 122.590 104.760 122.780 ;
        RECT 102.750 122.220 103.765 122.420 ;
        RECT 104.065 122.260 104.235 122.590 ;
        RECT 104.405 122.040 104.735 122.420 ;
        RECT 104.950 122.300 105.175 124.420 ;
        RECT 105.345 124.090 105.675 124.590 ;
        RECT 105.845 123.920 106.015 124.420 ;
        RECT 105.350 123.750 106.015 123.920 ;
        RECT 105.350 122.760 105.580 123.750 ;
        RECT 105.750 122.930 106.100 123.580 ;
        RECT 106.275 123.500 108.865 124.590 ;
        RECT 106.275 122.980 107.485 123.500 ;
        RECT 109.075 123.450 109.305 124.590 ;
        RECT 109.475 123.440 109.805 124.420 ;
        RECT 109.975 123.450 110.185 124.590 ;
        RECT 110.965 123.660 111.135 124.420 ;
        RECT 111.315 123.830 111.645 124.590 ;
        RECT 110.965 123.490 111.630 123.660 ;
        RECT 111.815 123.515 112.085 124.420 ;
        RECT 107.655 122.810 108.865 123.330 ;
        RECT 109.055 123.030 109.385 123.280 ;
        RECT 105.350 122.590 106.015 122.760 ;
        RECT 105.345 122.040 105.675 122.420 ;
        RECT 105.845 122.300 106.015 122.590 ;
        RECT 106.275 122.040 108.865 122.810 ;
        RECT 109.075 122.040 109.305 122.860 ;
        RECT 109.555 122.840 109.805 123.440 ;
        RECT 111.460 123.345 111.630 123.490 ;
        RECT 110.895 122.940 111.225 123.310 ;
        RECT 111.460 123.015 111.745 123.345 ;
        RECT 109.475 122.210 109.805 122.840 ;
        RECT 109.975 122.040 110.185 122.860 ;
        RECT 111.460 122.760 111.630 123.015 ;
        RECT 110.965 122.590 111.630 122.760 ;
        RECT 111.915 122.715 112.085 123.515 ;
        RECT 112.255 123.500 113.465 124.590 ;
        RECT 113.635 123.500 117.145 124.590 ;
        RECT 117.315 123.500 118.525 124.590 ;
        RECT 112.255 122.960 112.775 123.500 ;
        RECT 112.945 122.790 113.465 123.330 ;
        RECT 113.635 122.980 115.325 123.500 ;
        RECT 115.495 122.810 117.145 123.330 ;
        RECT 117.315 122.960 117.835 123.500 ;
        RECT 110.965 122.210 111.135 122.590 ;
        RECT 111.315 122.040 111.645 122.420 ;
        RECT 111.825 122.210 112.085 122.715 ;
        RECT 112.255 122.040 113.465 122.790 ;
        RECT 113.635 122.040 117.145 122.810 ;
        RECT 118.005 122.790 118.525 123.330 ;
        RECT 117.315 122.040 118.525 122.790 ;
        RECT 11.430 121.870 118.610 122.040 ;
        RECT 11.515 121.120 12.725 121.870 ;
        RECT 11.515 120.580 12.035 121.120 ;
        RECT 13.815 121.100 17.325 121.870 ;
        RECT 17.585 121.320 17.755 121.700 ;
        RECT 17.935 121.490 18.265 121.870 ;
        RECT 17.585 121.150 18.250 121.320 ;
        RECT 18.445 121.195 18.705 121.700 ;
        RECT 18.965 121.390 19.265 121.870 ;
        RECT 19.435 121.220 19.695 121.675 ;
        RECT 19.865 121.390 20.125 121.870 ;
        RECT 20.305 121.220 20.565 121.675 ;
        RECT 20.735 121.390 20.985 121.870 ;
        RECT 21.165 121.220 21.425 121.675 ;
        RECT 21.595 121.390 21.845 121.870 ;
        RECT 22.025 121.220 22.285 121.675 ;
        RECT 22.455 121.390 22.700 121.870 ;
        RECT 22.870 121.220 23.145 121.675 ;
        RECT 23.315 121.390 23.560 121.870 ;
        RECT 23.730 121.220 23.990 121.675 ;
        RECT 24.160 121.390 24.420 121.870 ;
        RECT 24.590 121.220 24.850 121.675 ;
        RECT 25.020 121.390 25.280 121.870 ;
        RECT 25.450 121.220 25.710 121.675 ;
        RECT 25.880 121.310 26.140 121.870 ;
        RECT 12.205 120.410 12.725 120.950 ;
        RECT 11.515 119.320 12.725 120.410 ;
        RECT 13.815 120.410 15.505 120.930 ;
        RECT 15.675 120.580 17.325 121.100 ;
        RECT 17.515 120.600 17.845 120.970 ;
        RECT 18.080 120.895 18.250 121.150 ;
        RECT 18.080 120.565 18.365 120.895 ;
        RECT 18.080 120.420 18.250 120.565 ;
        RECT 13.815 119.320 17.325 120.410 ;
        RECT 17.585 120.250 18.250 120.420 ;
        RECT 18.535 120.395 18.705 121.195 ;
        RECT 17.585 119.490 17.755 120.250 ;
        RECT 17.935 119.320 18.265 120.080 ;
        RECT 18.435 119.490 18.705 120.395 ;
        RECT 18.965 121.050 25.710 121.220 ;
        RECT 18.965 120.460 20.130 121.050 ;
        RECT 26.310 120.880 26.560 121.690 ;
        RECT 26.740 121.345 27.000 121.870 ;
        RECT 27.170 120.880 27.420 121.690 ;
        RECT 27.600 121.360 27.905 121.870 ;
        RECT 20.300 120.630 27.420 120.880 ;
        RECT 27.590 120.630 27.905 121.190 ;
        RECT 28.075 121.145 28.365 121.870 ;
        RECT 28.995 121.100 31.585 121.870 ;
        RECT 31.845 121.320 32.015 121.700 ;
        RECT 32.195 121.490 32.525 121.870 ;
        RECT 31.845 121.150 32.510 121.320 ;
        RECT 32.705 121.195 32.965 121.700 ;
        RECT 33.600 121.325 38.945 121.870 ;
        RECT 39.120 121.325 44.465 121.870 ;
        RECT 18.965 120.235 25.710 120.460 ;
        RECT 18.965 119.320 19.235 120.065 ;
        RECT 19.405 119.495 19.695 120.235 ;
        RECT 20.305 120.220 25.710 120.235 ;
        RECT 19.865 119.325 20.120 120.050 ;
        RECT 20.305 119.495 20.565 120.220 ;
        RECT 20.735 119.325 20.980 120.050 ;
        RECT 21.165 119.495 21.425 120.220 ;
        RECT 21.595 119.325 21.840 120.050 ;
        RECT 22.025 119.495 22.285 120.220 ;
        RECT 22.455 119.325 22.700 120.050 ;
        RECT 22.870 119.495 23.130 120.220 ;
        RECT 23.300 119.325 23.560 120.050 ;
        RECT 23.730 119.495 23.990 120.220 ;
        RECT 24.160 119.325 24.420 120.050 ;
        RECT 24.590 119.495 24.850 120.220 ;
        RECT 25.020 119.325 25.280 120.050 ;
        RECT 25.450 119.495 25.710 120.220 ;
        RECT 25.880 119.325 26.140 120.120 ;
        RECT 26.310 119.495 26.560 120.630 ;
        RECT 19.865 119.320 26.140 119.325 ;
        RECT 26.740 119.320 27.000 120.130 ;
        RECT 27.175 119.490 27.420 120.630 ;
        RECT 27.600 119.320 27.895 120.130 ;
        RECT 28.075 119.320 28.365 120.485 ;
        RECT 28.995 120.410 30.205 120.930 ;
        RECT 30.375 120.580 31.585 121.100 ;
        RECT 31.775 120.600 32.105 120.970 ;
        RECT 32.340 120.895 32.510 121.150 ;
        RECT 32.340 120.565 32.625 120.895 ;
        RECT 32.340 120.420 32.510 120.565 ;
        RECT 28.995 119.320 31.585 120.410 ;
        RECT 31.845 120.250 32.510 120.420 ;
        RECT 32.795 120.395 32.965 121.195 ;
        RECT 31.845 119.490 32.015 120.250 ;
        RECT 32.195 119.320 32.525 120.080 ;
        RECT 32.695 119.490 32.965 120.395 ;
        RECT 35.190 119.755 35.540 121.005 ;
        RECT 37.020 120.495 37.360 121.325 ;
        RECT 40.710 119.755 41.060 121.005 ;
        RECT 42.540 120.495 42.880 121.325 ;
        RECT 44.910 121.060 45.155 121.665 ;
        RECT 45.375 121.335 45.885 121.870 ;
        RECT 44.635 120.890 45.865 121.060 ;
        RECT 44.635 120.080 44.975 120.890 ;
        RECT 45.145 120.325 45.895 120.515 ;
        RECT 33.600 119.320 38.945 119.755 ;
        RECT 39.120 119.320 44.465 119.755 ;
        RECT 44.635 119.670 45.150 120.080 ;
        RECT 45.385 119.320 45.555 120.080 ;
        RECT 45.725 119.660 45.895 120.325 ;
        RECT 46.065 120.340 46.255 121.700 ;
        RECT 46.425 120.850 46.700 121.700 ;
        RECT 46.890 121.335 47.420 121.700 ;
        RECT 47.845 121.470 48.175 121.870 ;
        RECT 47.245 121.300 47.420 121.335 ;
        RECT 46.425 120.680 46.705 120.850 ;
        RECT 46.425 120.540 46.700 120.680 ;
        RECT 46.905 120.340 47.075 121.140 ;
        RECT 46.065 120.170 47.075 120.340 ;
        RECT 47.245 121.130 48.175 121.300 ;
        RECT 48.345 121.130 48.600 121.700 ;
        RECT 47.245 120.000 47.415 121.130 ;
        RECT 48.005 120.960 48.175 121.130 ;
        RECT 46.290 119.830 47.415 120.000 ;
        RECT 47.585 120.630 47.780 120.960 ;
        RECT 48.005 120.630 48.260 120.960 ;
        RECT 47.585 119.660 47.755 120.630 ;
        RECT 48.430 120.460 48.600 121.130 ;
        RECT 49.510 121.060 49.755 121.665 ;
        RECT 49.975 121.335 50.485 121.870 ;
        RECT 45.725 119.490 47.755 119.660 ;
        RECT 47.925 119.320 48.095 120.460 ;
        RECT 48.265 119.490 48.600 120.460 ;
        RECT 49.235 120.890 50.465 121.060 ;
        RECT 49.235 120.080 49.575 120.890 ;
        RECT 49.745 120.325 50.495 120.515 ;
        RECT 49.235 119.670 49.750 120.080 ;
        RECT 49.985 119.320 50.155 120.080 ;
        RECT 50.325 119.660 50.495 120.325 ;
        RECT 50.665 120.340 50.855 121.700 ;
        RECT 51.025 121.190 51.300 121.700 ;
        RECT 51.490 121.335 52.020 121.700 ;
        RECT 52.445 121.470 52.775 121.870 ;
        RECT 51.845 121.300 52.020 121.335 ;
        RECT 51.025 121.020 51.305 121.190 ;
        RECT 51.025 120.540 51.300 121.020 ;
        RECT 51.505 120.340 51.675 121.140 ;
        RECT 50.665 120.170 51.675 120.340 ;
        RECT 51.845 121.130 52.775 121.300 ;
        RECT 52.945 121.130 53.200 121.700 ;
        RECT 53.835 121.145 54.125 121.870 ;
        RECT 51.845 120.000 52.015 121.130 ;
        RECT 52.605 120.960 52.775 121.130 ;
        RECT 50.890 119.830 52.015 120.000 ;
        RECT 52.185 120.630 52.380 120.960 ;
        RECT 52.605 120.630 52.860 120.960 ;
        RECT 52.185 119.660 52.355 120.630 ;
        RECT 53.030 120.460 53.200 121.130 ;
        RECT 54.335 121.050 54.565 121.870 ;
        RECT 54.735 121.070 55.065 121.700 ;
        RECT 54.315 120.630 54.645 120.880 ;
        RECT 50.325 119.490 52.355 119.660 ;
        RECT 52.525 119.320 52.695 120.460 ;
        RECT 52.865 119.490 53.200 120.460 ;
        RECT 53.835 119.320 54.125 120.485 ;
        RECT 54.815 120.470 55.065 121.070 ;
        RECT 55.235 121.050 55.445 121.870 ;
        RECT 55.765 121.320 55.935 121.700 ;
        RECT 56.115 121.490 56.445 121.870 ;
        RECT 55.765 121.150 56.430 121.320 ;
        RECT 56.625 121.195 56.885 121.700 ;
        RECT 55.695 120.600 56.025 120.970 ;
        RECT 56.260 120.895 56.430 121.150 ;
        RECT 54.335 119.320 54.565 120.460 ;
        RECT 54.735 119.490 55.065 120.470 ;
        RECT 56.260 120.565 56.545 120.895 ;
        RECT 55.235 119.320 55.445 120.460 ;
        RECT 56.260 120.420 56.430 120.565 ;
        RECT 55.765 120.250 56.430 120.420 ;
        RECT 56.715 120.395 56.885 121.195 ;
        RECT 57.205 121.070 57.535 121.870 ;
        RECT 57.705 121.220 57.875 121.700 ;
        RECT 58.045 121.390 58.375 121.870 ;
        RECT 58.545 121.220 58.715 121.700 ;
        RECT 58.965 121.390 59.205 121.870 ;
        RECT 59.385 121.220 59.555 121.700 ;
        RECT 57.705 121.050 58.715 121.220 ;
        RECT 58.920 121.050 59.555 121.220 ;
        RECT 59.815 121.120 61.025 121.870 ;
        RECT 61.200 121.325 66.545 121.870 ;
        RECT 66.720 121.325 72.065 121.870 ;
        RECT 57.705 121.020 58.205 121.050 ;
        RECT 57.705 120.510 58.200 121.020 ;
        RECT 58.920 120.880 59.090 121.050 ;
        RECT 58.590 120.710 59.090 120.880 ;
        RECT 55.765 119.490 55.935 120.250 ;
        RECT 56.115 119.320 56.445 120.080 ;
        RECT 56.615 119.490 56.885 120.395 ;
        RECT 57.205 119.320 57.535 120.470 ;
        RECT 57.705 120.340 58.715 120.510 ;
        RECT 57.705 119.490 57.875 120.340 ;
        RECT 58.045 119.320 58.375 120.120 ;
        RECT 58.545 119.490 58.715 120.340 ;
        RECT 58.920 120.470 59.090 120.710 ;
        RECT 59.260 120.640 59.640 120.880 ;
        RECT 58.920 120.300 59.635 120.470 ;
        RECT 58.895 119.320 59.135 120.120 ;
        RECT 59.305 119.490 59.635 120.300 ;
        RECT 59.815 120.410 60.335 120.950 ;
        RECT 60.505 120.580 61.025 121.120 ;
        RECT 59.815 119.320 61.025 120.410 ;
        RECT 62.790 119.755 63.140 121.005 ;
        RECT 64.620 120.495 64.960 121.325 ;
        RECT 68.310 119.755 68.660 121.005 ;
        RECT 70.140 120.495 70.480 121.325 ;
        RECT 72.295 121.050 72.505 121.870 ;
        RECT 72.675 121.070 73.005 121.700 ;
        RECT 72.675 120.470 72.925 121.070 ;
        RECT 73.175 121.050 73.405 121.870 ;
        RECT 74.535 121.100 78.045 121.870 ;
        RECT 78.305 121.320 78.475 121.700 ;
        RECT 78.655 121.490 78.985 121.870 ;
        RECT 78.305 121.150 78.970 121.320 ;
        RECT 79.165 121.195 79.425 121.700 ;
        RECT 73.095 120.630 73.425 120.880 ;
        RECT 61.200 119.320 66.545 119.755 ;
        RECT 66.720 119.320 72.065 119.755 ;
        RECT 72.295 119.320 72.505 120.460 ;
        RECT 72.675 119.490 73.005 120.470 ;
        RECT 73.175 119.320 73.405 120.460 ;
        RECT 74.535 120.410 76.225 120.930 ;
        RECT 76.395 120.580 78.045 121.100 ;
        RECT 78.235 120.600 78.565 120.970 ;
        RECT 78.800 120.895 78.970 121.150 ;
        RECT 78.800 120.565 79.085 120.895 ;
        RECT 78.800 120.420 78.970 120.565 ;
        RECT 74.535 119.320 78.045 120.410 ;
        RECT 78.305 120.250 78.970 120.420 ;
        RECT 79.255 120.395 79.425 121.195 ;
        RECT 79.595 121.145 79.885 121.870 ;
        RECT 80.055 121.100 82.645 121.870 ;
        RECT 82.820 121.325 88.165 121.870 ;
        RECT 78.305 119.490 78.475 120.250 ;
        RECT 78.655 119.320 78.985 120.080 ;
        RECT 79.155 119.490 79.425 120.395 ;
        RECT 79.595 119.320 79.885 120.485 ;
        RECT 80.055 120.410 81.265 120.930 ;
        RECT 81.435 120.580 82.645 121.100 ;
        RECT 80.055 119.320 82.645 120.410 ;
        RECT 84.410 119.755 84.760 121.005 ;
        RECT 86.240 120.495 86.580 121.325 ;
        RECT 88.425 121.320 88.595 121.700 ;
        RECT 88.775 121.490 89.105 121.870 ;
        RECT 88.425 121.150 89.090 121.320 ;
        RECT 89.285 121.195 89.545 121.700 ;
        RECT 88.355 120.600 88.685 120.970 ;
        RECT 88.920 120.895 89.090 121.150 ;
        RECT 88.920 120.565 89.205 120.895 ;
        RECT 88.920 120.420 89.090 120.565 ;
        RECT 88.425 120.250 89.090 120.420 ;
        RECT 89.375 120.395 89.545 121.195 ;
        RECT 90.635 121.100 94.145 121.870 ;
        RECT 94.320 121.325 99.665 121.870 ;
        RECT 99.840 121.325 105.185 121.870 ;
        RECT 82.820 119.320 88.165 119.755 ;
        RECT 88.425 119.490 88.595 120.250 ;
        RECT 88.775 119.320 89.105 120.080 ;
        RECT 89.275 119.490 89.545 120.395 ;
        RECT 90.635 120.410 92.325 120.930 ;
        RECT 92.495 120.580 94.145 121.100 ;
        RECT 90.635 119.320 94.145 120.410 ;
        RECT 95.910 119.755 96.260 121.005 ;
        RECT 97.740 120.495 98.080 121.325 ;
        RECT 101.430 119.755 101.780 121.005 ;
        RECT 103.260 120.495 103.600 121.325 ;
        RECT 105.355 121.145 105.645 121.870 ;
        RECT 105.815 121.120 107.025 121.870 ;
        RECT 94.320 119.320 99.665 119.755 ;
        RECT 99.840 119.320 105.185 119.755 ;
        RECT 105.355 119.320 105.645 120.485 ;
        RECT 105.815 120.410 106.335 120.950 ;
        RECT 106.505 120.580 107.025 121.120 ;
        RECT 107.195 121.100 110.705 121.870 ;
        RECT 107.195 120.410 108.885 120.930 ;
        RECT 109.055 120.580 110.705 121.100 ;
        RECT 110.915 121.050 111.145 121.870 ;
        RECT 111.315 121.070 111.645 121.700 ;
        RECT 110.895 120.630 111.225 120.880 ;
        RECT 111.395 120.470 111.645 121.070 ;
        RECT 111.815 121.050 112.025 121.870 ;
        RECT 113.265 121.320 113.435 121.700 ;
        RECT 113.615 121.490 113.945 121.870 ;
        RECT 113.265 121.150 113.930 121.320 ;
        RECT 114.125 121.195 114.385 121.700 ;
        RECT 113.195 120.600 113.525 120.970 ;
        RECT 113.760 120.895 113.930 121.150 ;
        RECT 105.815 119.320 107.025 120.410 ;
        RECT 107.195 119.320 110.705 120.410 ;
        RECT 110.915 119.320 111.145 120.460 ;
        RECT 111.315 119.490 111.645 120.470 ;
        RECT 113.760 120.565 114.045 120.895 ;
        RECT 111.815 119.320 112.025 120.460 ;
        RECT 113.760 120.420 113.930 120.565 ;
        RECT 113.265 120.250 113.930 120.420 ;
        RECT 114.215 120.395 114.385 121.195 ;
        RECT 114.555 121.120 115.765 121.870 ;
        RECT 113.265 119.490 113.435 120.250 ;
        RECT 113.615 119.320 113.945 120.080 ;
        RECT 114.115 119.490 114.385 120.395 ;
        RECT 114.555 120.410 115.075 120.950 ;
        RECT 115.245 120.580 115.765 121.120 ;
        RECT 115.935 121.195 116.195 121.700 ;
        RECT 116.375 121.490 116.705 121.870 ;
        RECT 116.885 121.320 117.055 121.700 ;
        RECT 114.555 119.320 115.765 120.410 ;
        RECT 115.935 120.395 116.115 121.195 ;
        RECT 116.390 121.150 117.055 121.320 ;
        RECT 116.390 120.895 116.560 121.150 ;
        RECT 117.315 121.120 118.525 121.870 ;
        RECT 116.285 120.565 116.560 120.895 ;
        RECT 116.785 120.600 117.125 120.970 ;
        RECT 116.390 120.420 116.560 120.565 ;
        RECT 115.935 119.490 116.205 120.395 ;
        RECT 116.390 120.250 117.065 120.420 ;
        RECT 116.375 119.320 116.705 120.080 ;
        RECT 116.885 119.490 117.065 120.250 ;
        RECT 117.315 120.410 117.835 120.950 ;
        RECT 118.005 120.580 118.525 121.120 ;
        RECT 117.315 119.320 118.525 120.410 ;
        RECT 11.430 119.150 118.610 119.320 ;
        RECT 11.515 118.060 12.725 119.150 ;
        RECT 11.515 117.350 12.035 117.890 ;
        RECT 12.205 117.520 12.725 118.060 ;
        RECT 13.355 118.060 15.025 119.150 ;
        RECT 13.355 117.540 14.105 118.060 ;
        RECT 15.195 117.985 15.485 119.150 ;
        RECT 15.655 118.060 18.245 119.150 ;
        RECT 18.420 118.715 23.765 119.150 ;
        RECT 14.275 117.370 15.025 117.890 ;
        RECT 15.655 117.540 16.865 118.060 ;
        RECT 17.035 117.370 18.245 117.890 ;
        RECT 20.010 117.465 20.360 118.715 ;
        RECT 23.935 118.075 24.205 118.980 ;
        RECT 24.375 118.390 24.705 119.150 ;
        RECT 24.885 118.220 25.055 118.980 ;
        RECT 11.515 116.600 12.725 117.350 ;
        RECT 13.355 116.600 15.025 117.370 ;
        RECT 15.195 116.600 15.485 117.325 ;
        RECT 15.655 116.600 18.245 117.370 ;
        RECT 21.840 117.145 22.180 117.975 ;
        RECT 23.935 117.275 24.105 118.075 ;
        RECT 24.390 118.050 25.055 118.220 ;
        RECT 25.315 118.060 26.525 119.150 ;
        RECT 26.695 118.060 30.205 119.150 ;
        RECT 30.685 118.310 30.855 119.150 ;
        RECT 31.065 118.140 31.315 118.980 ;
        RECT 31.525 118.310 31.695 119.150 ;
        RECT 31.865 118.140 32.155 118.980 ;
        RECT 24.390 117.905 24.560 118.050 ;
        RECT 24.275 117.575 24.560 117.905 ;
        RECT 24.390 117.320 24.560 117.575 ;
        RECT 24.795 117.500 25.125 117.870 ;
        RECT 25.315 117.520 25.835 118.060 ;
        RECT 26.005 117.350 26.525 117.890 ;
        RECT 26.695 117.540 28.385 118.060 ;
        RECT 30.430 117.970 32.155 118.140 ;
        RECT 32.365 118.090 32.535 119.150 ;
        RECT 32.830 118.770 33.160 119.150 ;
        RECT 33.340 118.600 33.510 118.890 ;
        RECT 33.680 118.690 33.930 119.150 ;
        RECT 32.710 118.430 33.510 118.600 ;
        RECT 34.100 118.640 34.970 118.980 ;
        RECT 28.555 117.370 30.205 117.890 ;
        RECT 18.420 116.600 23.765 117.145 ;
        RECT 23.935 116.770 24.195 117.275 ;
        RECT 24.390 117.150 25.055 117.320 ;
        RECT 24.375 116.600 24.705 116.980 ;
        RECT 24.885 116.770 25.055 117.150 ;
        RECT 25.315 116.600 26.525 117.350 ;
        RECT 26.695 116.600 30.205 117.370 ;
        RECT 30.430 117.420 30.840 117.970 ;
        RECT 32.710 117.810 32.880 118.430 ;
        RECT 34.100 118.260 34.270 118.640 ;
        RECT 35.205 118.520 35.375 118.980 ;
        RECT 35.545 118.690 35.915 119.150 ;
        RECT 36.210 118.550 36.380 118.890 ;
        RECT 36.550 118.720 36.880 119.150 ;
        RECT 37.115 118.550 37.285 118.890 ;
        RECT 33.050 118.090 34.270 118.260 ;
        RECT 34.440 118.180 34.900 118.470 ;
        RECT 35.205 118.350 35.765 118.520 ;
        RECT 36.210 118.380 37.285 118.550 ;
        RECT 37.455 118.650 38.135 118.980 ;
        RECT 38.350 118.650 38.600 118.980 ;
        RECT 38.770 118.690 39.020 119.150 ;
        RECT 35.595 118.210 35.765 118.350 ;
        RECT 34.440 118.170 35.405 118.180 ;
        RECT 34.100 118.000 34.270 118.090 ;
        RECT 34.730 118.010 35.405 118.170 ;
        RECT 32.710 117.800 33.055 117.810 ;
        RECT 31.025 117.590 33.055 117.800 ;
        RECT 30.430 117.250 32.195 117.420 ;
        RECT 30.685 116.600 30.855 117.070 ;
        RECT 31.025 116.770 31.355 117.250 ;
        RECT 31.525 116.600 31.695 117.070 ;
        RECT 31.865 116.770 32.195 117.250 ;
        RECT 32.365 116.600 32.535 117.410 ;
        RECT 32.730 117.335 33.055 117.590 ;
        RECT 32.735 116.980 33.055 117.335 ;
        RECT 33.225 117.550 33.765 117.920 ;
        RECT 34.100 117.830 34.505 118.000 ;
        RECT 33.225 117.150 33.465 117.550 ;
        RECT 33.945 117.380 34.165 117.660 ;
        RECT 33.635 117.210 34.165 117.380 ;
        RECT 33.635 116.980 33.805 117.210 ;
        RECT 34.335 117.050 34.505 117.830 ;
        RECT 34.675 117.220 35.025 117.840 ;
        RECT 35.195 117.220 35.405 118.010 ;
        RECT 35.595 118.040 37.095 118.210 ;
        RECT 35.595 117.350 35.765 118.040 ;
        RECT 37.455 117.870 37.625 118.650 ;
        RECT 38.430 118.520 38.600 118.650 ;
        RECT 35.935 117.700 37.625 117.870 ;
        RECT 37.795 118.090 38.260 118.480 ;
        RECT 38.430 118.350 38.825 118.520 ;
        RECT 35.935 117.520 36.105 117.700 ;
        RECT 32.735 116.810 33.805 116.980 ;
        RECT 33.975 116.600 34.165 117.040 ;
        RECT 34.335 116.770 35.285 117.050 ;
        RECT 35.595 116.960 35.855 117.350 ;
        RECT 36.275 117.280 37.065 117.530 ;
        RECT 35.505 116.790 35.855 116.960 ;
        RECT 36.065 116.600 36.395 117.060 ;
        RECT 37.270 116.990 37.440 117.700 ;
        RECT 37.795 117.500 37.965 118.090 ;
        RECT 37.610 117.280 37.965 117.500 ;
        RECT 38.135 117.280 38.485 117.900 ;
        RECT 38.655 116.990 38.825 118.350 ;
        RECT 39.190 118.180 39.515 118.965 ;
        RECT 38.995 117.130 39.455 118.180 ;
        RECT 37.270 116.820 38.125 116.990 ;
        RECT 38.330 116.820 38.825 116.990 ;
        RECT 38.995 116.600 39.325 116.960 ;
        RECT 39.685 116.860 39.855 118.980 ;
        RECT 40.025 118.650 40.355 119.150 ;
        RECT 40.525 118.480 40.780 118.980 ;
        RECT 40.030 118.310 40.780 118.480 ;
        RECT 40.030 117.320 40.260 118.310 ;
        RECT 40.430 117.490 40.780 118.140 ;
        RECT 40.955 117.985 41.245 119.150 ;
        RECT 41.415 118.075 41.685 118.980 ;
        RECT 41.855 118.390 42.185 119.150 ;
        RECT 42.365 118.220 42.535 118.980 ;
        RECT 40.030 117.150 40.780 117.320 ;
        RECT 40.025 116.600 40.355 116.980 ;
        RECT 40.525 116.860 40.780 117.150 ;
        RECT 40.955 116.600 41.245 117.325 ;
        RECT 41.415 117.275 41.585 118.075 ;
        RECT 41.870 118.050 42.535 118.220 ;
        RECT 42.795 118.075 43.065 118.980 ;
        RECT 43.235 118.390 43.565 119.150 ;
        RECT 43.745 118.220 43.915 118.980 ;
        RECT 41.870 117.905 42.040 118.050 ;
        RECT 41.755 117.575 42.040 117.905 ;
        RECT 41.870 117.320 42.040 117.575 ;
        RECT 42.275 117.500 42.605 117.870 ;
        RECT 41.415 116.770 41.675 117.275 ;
        RECT 41.870 117.150 42.535 117.320 ;
        RECT 41.855 116.600 42.185 116.980 ;
        RECT 42.365 116.770 42.535 117.150 ;
        RECT 42.795 117.275 42.965 118.075 ;
        RECT 43.250 118.050 43.915 118.220 ;
        RECT 44.175 118.060 46.765 119.150 ;
        RECT 47.025 118.220 47.195 118.980 ;
        RECT 47.375 118.390 47.705 119.150 ;
        RECT 43.250 117.905 43.420 118.050 ;
        RECT 43.135 117.575 43.420 117.905 ;
        RECT 43.250 117.320 43.420 117.575 ;
        RECT 43.655 117.500 43.985 117.870 ;
        RECT 44.175 117.540 45.385 118.060 ;
        RECT 47.025 118.050 47.690 118.220 ;
        RECT 47.875 118.075 48.145 118.980 ;
        RECT 47.520 117.905 47.690 118.050 ;
        RECT 45.555 117.370 46.765 117.890 ;
        RECT 46.955 117.500 47.285 117.870 ;
        RECT 47.520 117.575 47.805 117.905 ;
        RECT 42.795 116.770 43.055 117.275 ;
        RECT 43.250 117.150 43.915 117.320 ;
        RECT 43.235 116.600 43.565 116.980 ;
        RECT 43.745 116.770 43.915 117.150 ;
        RECT 44.175 116.600 46.765 117.370 ;
        RECT 47.520 117.320 47.690 117.575 ;
        RECT 47.025 117.150 47.690 117.320 ;
        RECT 47.975 117.275 48.145 118.075 ;
        RECT 48.405 118.220 48.575 118.980 ;
        RECT 48.755 118.390 49.085 119.150 ;
        RECT 48.405 118.050 49.070 118.220 ;
        RECT 49.255 118.075 49.525 118.980 ;
        RECT 48.900 117.905 49.070 118.050 ;
        RECT 48.335 117.500 48.665 117.870 ;
        RECT 48.900 117.575 49.185 117.905 ;
        RECT 48.900 117.320 49.070 117.575 ;
        RECT 47.025 116.770 47.195 117.150 ;
        RECT 47.375 116.600 47.705 116.980 ;
        RECT 47.885 116.770 48.145 117.275 ;
        RECT 48.405 117.150 49.070 117.320 ;
        RECT 49.355 117.275 49.525 118.075 ;
        RECT 50.155 118.060 51.825 119.150 ;
        RECT 52.000 118.715 57.345 119.150 ;
        RECT 50.155 117.540 50.905 118.060 ;
        RECT 51.075 117.370 51.825 117.890 ;
        RECT 53.590 117.465 53.940 118.715 ;
        RECT 57.555 118.010 57.785 119.150 ;
        RECT 57.955 118.000 58.285 118.980 ;
        RECT 58.455 118.010 58.665 119.150 ;
        RECT 59.045 118.000 59.375 119.150 ;
        RECT 59.545 118.130 59.715 118.980 ;
        RECT 59.885 118.350 60.215 119.150 ;
        RECT 60.385 118.130 60.555 118.980 ;
        RECT 60.735 118.350 60.975 119.150 ;
        RECT 61.145 118.170 61.475 118.980 ;
        RECT 48.405 116.770 48.575 117.150 ;
        RECT 48.755 116.600 49.085 116.980 ;
        RECT 49.265 116.770 49.525 117.275 ;
        RECT 50.155 116.600 51.825 117.370 ;
        RECT 55.420 117.145 55.760 117.975 ;
        RECT 57.535 117.590 57.865 117.840 ;
        RECT 52.000 116.600 57.345 117.145 ;
        RECT 57.555 116.600 57.785 117.420 ;
        RECT 58.035 117.400 58.285 118.000 ;
        RECT 59.545 117.960 60.555 118.130 ;
        RECT 60.760 118.000 61.475 118.170 ;
        RECT 61.655 118.060 63.325 119.150 ;
        RECT 63.585 118.220 63.755 118.980 ;
        RECT 63.935 118.390 64.265 119.150 ;
        RECT 59.545 117.790 60.040 117.960 ;
        RECT 59.545 117.620 60.045 117.790 ;
        RECT 60.760 117.760 60.930 118.000 ;
        RECT 59.545 117.420 60.040 117.620 ;
        RECT 60.430 117.590 60.930 117.760 ;
        RECT 61.100 117.590 61.480 117.830 ;
        RECT 60.760 117.420 60.930 117.590 ;
        RECT 61.655 117.540 62.405 118.060 ;
        RECT 63.585 118.050 64.250 118.220 ;
        RECT 64.435 118.075 64.705 118.980 ;
        RECT 64.080 117.905 64.250 118.050 ;
        RECT 57.955 116.770 58.285 117.400 ;
        RECT 58.455 116.600 58.665 117.420 ;
        RECT 59.045 116.600 59.375 117.400 ;
        RECT 59.545 117.250 60.555 117.420 ;
        RECT 60.760 117.250 61.395 117.420 ;
        RECT 62.575 117.370 63.325 117.890 ;
        RECT 63.515 117.500 63.845 117.870 ;
        RECT 64.080 117.575 64.365 117.905 ;
        RECT 59.545 116.770 59.715 117.250 ;
        RECT 59.885 116.600 60.215 117.080 ;
        RECT 60.385 116.770 60.555 117.250 ;
        RECT 60.805 116.600 61.045 117.080 ;
        RECT 61.225 116.770 61.395 117.250 ;
        RECT 61.655 116.600 63.325 117.370 ;
        RECT 64.080 117.320 64.250 117.575 ;
        RECT 63.585 117.150 64.250 117.320 ;
        RECT 64.535 117.275 64.705 118.075 ;
        RECT 64.875 118.060 66.545 119.150 ;
        RECT 64.875 117.540 65.625 118.060 ;
        RECT 66.715 117.985 67.005 119.150 ;
        RECT 67.175 118.060 68.385 119.150 ;
        RECT 65.795 117.370 66.545 117.890 ;
        RECT 67.175 117.520 67.695 118.060 ;
        RECT 68.615 118.010 68.825 119.150 ;
        RECT 68.995 118.000 69.325 118.980 ;
        RECT 69.495 118.010 69.725 119.150 ;
        RECT 69.945 118.170 70.275 118.980 ;
        RECT 70.445 118.350 70.685 119.150 ;
        RECT 69.945 118.000 70.660 118.170 ;
        RECT 63.585 116.770 63.755 117.150 ;
        RECT 63.935 116.600 64.265 116.980 ;
        RECT 64.445 116.770 64.705 117.275 ;
        RECT 64.875 116.600 66.545 117.370 ;
        RECT 67.865 117.350 68.385 117.890 ;
        RECT 66.715 116.600 67.005 117.325 ;
        RECT 67.175 116.600 68.385 117.350 ;
        RECT 68.615 116.600 68.825 117.420 ;
        RECT 68.995 117.400 69.245 118.000 ;
        RECT 69.415 117.590 69.745 117.840 ;
        RECT 69.940 117.590 70.320 117.830 ;
        RECT 70.490 117.760 70.660 118.000 ;
        RECT 70.865 118.130 71.035 118.980 ;
        RECT 71.205 118.350 71.535 119.150 ;
        RECT 71.705 118.130 71.875 118.980 ;
        RECT 70.865 117.960 71.875 118.130 ;
        RECT 72.045 118.000 72.375 119.150 ;
        RECT 72.785 118.220 72.955 118.980 ;
        RECT 73.135 118.390 73.465 119.150 ;
        RECT 72.785 118.050 73.450 118.220 ;
        RECT 73.635 118.075 73.905 118.980 ;
        RECT 70.490 117.590 70.990 117.760 ;
        RECT 70.490 117.420 70.660 117.590 ;
        RECT 71.380 117.420 71.875 117.960 ;
        RECT 73.280 117.905 73.450 118.050 ;
        RECT 72.715 117.500 73.045 117.870 ;
        RECT 73.280 117.575 73.565 117.905 ;
        RECT 68.995 116.770 69.325 117.400 ;
        RECT 69.495 116.600 69.725 117.420 ;
        RECT 70.025 117.250 70.660 117.420 ;
        RECT 70.865 117.250 71.875 117.420 ;
        RECT 70.025 116.770 70.195 117.250 ;
        RECT 70.375 116.600 70.615 117.080 ;
        RECT 70.865 116.770 71.035 117.250 ;
        RECT 71.205 116.600 71.535 117.080 ;
        RECT 71.705 116.770 71.875 117.250 ;
        RECT 72.045 116.600 72.375 117.400 ;
        RECT 73.280 117.320 73.450 117.575 ;
        RECT 72.785 117.150 73.450 117.320 ;
        RECT 73.735 117.275 73.905 118.075 ;
        RECT 74.165 118.220 74.335 118.980 ;
        RECT 74.515 118.390 74.845 119.150 ;
        RECT 74.165 118.050 74.830 118.220 ;
        RECT 75.015 118.075 75.285 118.980 ;
        RECT 74.660 117.905 74.830 118.050 ;
        RECT 74.095 117.500 74.425 117.870 ;
        RECT 74.660 117.575 74.945 117.905 ;
        RECT 74.660 117.320 74.830 117.575 ;
        RECT 72.785 116.770 72.955 117.150 ;
        RECT 73.135 116.600 73.465 116.980 ;
        RECT 73.645 116.770 73.905 117.275 ;
        RECT 74.165 117.150 74.830 117.320 ;
        RECT 75.115 117.275 75.285 118.075 ;
        RECT 75.915 118.060 77.585 119.150 ;
        RECT 77.845 118.220 78.015 118.980 ;
        RECT 78.195 118.390 78.525 119.150 ;
        RECT 75.915 117.540 76.665 118.060 ;
        RECT 77.845 118.050 78.510 118.220 ;
        RECT 78.695 118.075 78.965 118.980 ;
        RECT 79.600 118.715 84.945 119.150 ;
        RECT 78.340 117.905 78.510 118.050 ;
        RECT 76.835 117.370 77.585 117.890 ;
        RECT 77.775 117.500 78.105 117.870 ;
        RECT 78.340 117.575 78.625 117.905 ;
        RECT 74.165 116.770 74.335 117.150 ;
        RECT 74.515 116.600 74.845 116.980 ;
        RECT 75.025 116.770 75.285 117.275 ;
        RECT 75.915 116.600 77.585 117.370 ;
        RECT 78.340 117.320 78.510 117.575 ;
        RECT 77.845 117.150 78.510 117.320 ;
        RECT 78.795 117.275 78.965 118.075 ;
        RECT 81.190 117.465 81.540 118.715 ;
        RECT 85.205 118.220 85.375 118.980 ;
        RECT 85.555 118.390 85.885 119.150 ;
        RECT 85.205 118.050 85.870 118.220 ;
        RECT 86.055 118.075 86.325 118.980 ;
        RECT 86.960 118.715 92.305 119.150 ;
        RECT 77.845 116.770 78.015 117.150 ;
        RECT 78.195 116.600 78.525 116.980 ;
        RECT 78.705 116.770 78.965 117.275 ;
        RECT 83.020 117.145 83.360 117.975 ;
        RECT 85.700 117.905 85.870 118.050 ;
        RECT 85.135 117.500 85.465 117.870 ;
        RECT 85.700 117.575 85.985 117.905 ;
        RECT 85.700 117.320 85.870 117.575 ;
        RECT 85.205 117.150 85.870 117.320 ;
        RECT 86.155 117.275 86.325 118.075 ;
        RECT 88.550 117.465 88.900 118.715 ;
        RECT 92.475 117.985 92.765 119.150 ;
        RECT 92.935 118.060 94.145 119.150 ;
        RECT 94.315 118.060 97.825 119.150 ;
        RECT 98.085 118.220 98.255 118.980 ;
        RECT 98.435 118.390 98.765 119.150 ;
        RECT 79.600 116.600 84.945 117.145 ;
        RECT 85.205 116.770 85.375 117.150 ;
        RECT 85.555 116.600 85.885 116.980 ;
        RECT 86.065 116.770 86.325 117.275 ;
        RECT 90.380 117.145 90.720 117.975 ;
        RECT 92.935 117.520 93.455 118.060 ;
        RECT 93.625 117.350 94.145 117.890 ;
        RECT 94.315 117.540 96.005 118.060 ;
        RECT 98.085 118.050 98.750 118.220 ;
        RECT 98.935 118.075 99.205 118.980 ;
        RECT 98.580 117.905 98.750 118.050 ;
        RECT 96.175 117.370 97.825 117.890 ;
        RECT 98.015 117.500 98.345 117.870 ;
        RECT 98.580 117.575 98.865 117.905 ;
        RECT 86.960 116.600 92.305 117.145 ;
        RECT 92.475 116.600 92.765 117.325 ;
        RECT 92.935 116.600 94.145 117.350 ;
        RECT 94.315 116.600 97.825 117.370 ;
        RECT 98.580 117.320 98.750 117.575 ;
        RECT 98.085 117.150 98.750 117.320 ;
        RECT 99.035 117.275 99.205 118.075 ;
        RECT 99.895 118.010 100.105 119.150 ;
        RECT 100.275 118.000 100.605 118.980 ;
        RECT 100.775 118.010 101.005 119.150 ;
        RECT 101.305 118.220 101.475 118.980 ;
        RECT 101.655 118.390 101.985 119.150 ;
        RECT 101.305 118.050 101.970 118.220 ;
        RECT 102.155 118.075 102.425 118.980 ;
        RECT 98.085 116.770 98.255 117.150 ;
        RECT 98.435 116.600 98.765 116.980 ;
        RECT 98.945 116.770 99.205 117.275 ;
        RECT 99.895 116.600 100.105 117.420 ;
        RECT 100.275 117.400 100.525 118.000 ;
        RECT 101.800 117.905 101.970 118.050 ;
        RECT 100.695 117.590 101.025 117.840 ;
        RECT 101.235 117.500 101.565 117.870 ;
        RECT 101.800 117.575 102.085 117.905 ;
        RECT 100.275 116.770 100.605 117.400 ;
        RECT 100.775 116.600 101.005 117.420 ;
        RECT 101.800 117.320 101.970 117.575 ;
        RECT 101.305 117.150 101.970 117.320 ;
        RECT 102.255 117.275 102.425 118.075 ;
        RECT 102.595 118.060 103.805 119.150 ;
        RECT 102.595 117.520 103.115 118.060 ;
        RECT 104.015 118.010 104.245 119.150 ;
        RECT 104.415 118.000 104.745 118.980 ;
        RECT 104.915 118.010 105.125 119.150 ;
        RECT 105.445 118.220 105.615 118.980 ;
        RECT 105.795 118.390 106.125 119.150 ;
        RECT 105.445 118.050 106.110 118.220 ;
        RECT 106.295 118.075 106.565 118.980 ;
        RECT 106.740 118.480 106.995 118.980 ;
        RECT 107.165 118.650 107.495 119.150 ;
        RECT 106.740 118.310 107.490 118.480 ;
        RECT 103.285 117.350 103.805 117.890 ;
        RECT 103.995 117.590 104.325 117.840 ;
        RECT 101.305 116.770 101.475 117.150 ;
        RECT 101.655 116.600 101.985 116.980 ;
        RECT 102.165 116.770 102.425 117.275 ;
        RECT 102.595 116.600 103.805 117.350 ;
        RECT 104.015 116.600 104.245 117.420 ;
        RECT 104.495 117.400 104.745 118.000 ;
        RECT 105.940 117.905 106.110 118.050 ;
        RECT 105.375 117.500 105.705 117.870 ;
        RECT 105.940 117.575 106.225 117.905 ;
        RECT 104.415 116.770 104.745 117.400 ;
        RECT 104.915 116.600 105.125 117.420 ;
        RECT 105.940 117.320 106.110 117.575 ;
        RECT 105.445 117.150 106.110 117.320 ;
        RECT 106.395 117.275 106.565 118.075 ;
        RECT 106.740 117.490 107.090 118.140 ;
        RECT 107.260 117.320 107.490 118.310 ;
        RECT 105.445 116.770 105.615 117.150 ;
        RECT 105.795 116.600 106.125 116.980 ;
        RECT 106.305 116.770 106.565 117.275 ;
        RECT 106.740 117.150 107.490 117.320 ;
        RECT 106.740 116.860 106.995 117.150 ;
        RECT 107.165 116.600 107.495 116.980 ;
        RECT 107.665 116.860 107.835 118.980 ;
        RECT 108.005 118.180 108.330 118.965 ;
        RECT 108.500 118.690 108.750 119.150 ;
        RECT 108.920 118.650 109.170 118.980 ;
        RECT 109.385 118.650 110.065 118.980 ;
        RECT 108.920 118.520 109.090 118.650 ;
        RECT 108.695 118.350 109.090 118.520 ;
        RECT 108.065 117.130 108.525 118.180 ;
        RECT 108.695 116.990 108.865 118.350 ;
        RECT 109.260 118.090 109.725 118.480 ;
        RECT 109.035 117.280 109.385 117.900 ;
        RECT 109.555 117.500 109.725 118.090 ;
        RECT 109.895 117.870 110.065 118.650 ;
        RECT 110.235 118.550 110.405 118.890 ;
        RECT 110.640 118.720 110.970 119.150 ;
        RECT 111.140 118.550 111.310 118.890 ;
        RECT 111.605 118.690 111.975 119.150 ;
        RECT 110.235 118.380 111.310 118.550 ;
        RECT 112.145 118.520 112.315 118.980 ;
        RECT 112.550 118.640 113.420 118.980 ;
        RECT 113.590 118.690 113.840 119.150 ;
        RECT 111.755 118.350 112.315 118.520 ;
        RECT 111.755 118.210 111.925 118.350 ;
        RECT 110.425 118.040 111.925 118.210 ;
        RECT 112.620 118.180 113.080 118.470 ;
        RECT 109.895 117.700 111.585 117.870 ;
        RECT 109.555 117.280 109.910 117.500 ;
        RECT 110.080 116.990 110.250 117.700 ;
        RECT 110.455 117.280 111.245 117.530 ;
        RECT 111.415 117.520 111.585 117.700 ;
        RECT 111.755 117.350 111.925 118.040 ;
        RECT 108.195 116.600 108.525 116.960 ;
        RECT 108.695 116.820 109.190 116.990 ;
        RECT 109.395 116.820 110.250 116.990 ;
        RECT 111.125 116.600 111.455 117.060 ;
        RECT 111.665 116.960 111.925 117.350 ;
        RECT 112.115 118.170 113.080 118.180 ;
        RECT 113.250 118.260 113.420 118.640 ;
        RECT 114.010 118.600 114.180 118.890 ;
        RECT 114.360 118.770 114.690 119.150 ;
        RECT 114.010 118.430 114.810 118.600 ;
        RECT 112.115 118.010 112.790 118.170 ;
        RECT 113.250 118.090 114.470 118.260 ;
        RECT 112.115 117.220 112.325 118.010 ;
        RECT 113.250 118.000 113.420 118.090 ;
        RECT 112.495 117.220 112.845 117.840 ;
        RECT 113.015 117.830 113.420 118.000 ;
        RECT 113.015 117.050 113.185 117.830 ;
        RECT 113.355 117.380 113.575 117.660 ;
        RECT 113.755 117.550 114.295 117.920 ;
        RECT 114.640 117.810 114.810 118.430 ;
        RECT 114.985 118.090 115.155 119.150 ;
        RECT 115.365 118.140 115.655 118.980 ;
        RECT 115.825 118.310 115.995 119.150 ;
        RECT 116.205 118.140 116.455 118.980 ;
        RECT 116.665 118.310 116.835 119.150 ;
        RECT 115.365 117.970 117.090 118.140 ;
        RECT 113.355 117.210 113.885 117.380 ;
        RECT 111.665 116.790 112.015 116.960 ;
        RECT 112.235 116.770 113.185 117.050 ;
        RECT 113.355 116.600 113.545 117.040 ;
        RECT 113.715 116.980 113.885 117.210 ;
        RECT 114.055 117.150 114.295 117.550 ;
        RECT 114.465 117.800 114.810 117.810 ;
        RECT 114.465 117.590 116.495 117.800 ;
        RECT 114.465 117.335 114.790 117.590 ;
        RECT 116.680 117.420 117.090 117.970 ;
        RECT 117.315 118.060 118.525 119.150 ;
        RECT 117.315 117.520 117.835 118.060 ;
        RECT 114.465 116.980 114.785 117.335 ;
        RECT 113.715 116.810 114.785 116.980 ;
        RECT 114.985 116.600 115.155 117.410 ;
        RECT 115.325 117.250 117.090 117.420 ;
        RECT 118.005 117.350 118.525 117.890 ;
        RECT 115.325 116.770 115.655 117.250 ;
        RECT 115.825 116.600 115.995 117.070 ;
        RECT 116.165 116.770 116.495 117.250 ;
        RECT 116.665 116.600 116.835 117.070 ;
        RECT 117.315 116.600 118.525 117.350 ;
        RECT 11.430 116.430 118.610 116.600 ;
        RECT 11.515 115.680 12.725 116.430 ;
        RECT 11.515 115.140 12.035 115.680 ;
        RECT 13.355 115.660 15.945 116.430 ;
        RECT 16.425 115.960 16.595 116.430 ;
        RECT 16.765 115.780 17.095 116.260 ;
        RECT 17.265 115.960 17.435 116.430 ;
        RECT 17.605 115.780 17.935 116.260 ;
        RECT 12.205 114.970 12.725 115.510 ;
        RECT 11.515 113.880 12.725 114.970 ;
        RECT 13.355 114.970 14.565 115.490 ;
        RECT 14.735 115.140 15.945 115.660 ;
        RECT 16.170 115.610 17.935 115.780 ;
        RECT 18.105 115.620 18.275 116.430 ;
        RECT 18.475 116.050 19.545 116.220 ;
        RECT 18.475 115.695 18.795 116.050 ;
        RECT 16.170 115.060 16.580 115.610 ;
        RECT 18.470 115.440 18.795 115.695 ;
        RECT 16.765 115.230 18.795 115.440 ;
        RECT 18.450 115.220 18.795 115.230 ;
        RECT 18.965 115.480 19.205 115.880 ;
        RECT 19.375 115.820 19.545 116.050 ;
        RECT 19.715 115.990 19.905 116.430 ;
        RECT 20.075 115.980 21.025 116.260 ;
        RECT 21.245 116.070 21.595 116.240 ;
        RECT 19.375 115.650 19.905 115.820 ;
        RECT 13.355 113.880 15.945 114.970 ;
        RECT 16.170 114.890 17.895 115.060 ;
        RECT 16.425 113.880 16.595 114.720 ;
        RECT 16.805 114.050 17.055 114.890 ;
        RECT 17.265 113.880 17.435 114.720 ;
        RECT 17.605 114.050 17.895 114.890 ;
        RECT 18.105 113.880 18.275 114.940 ;
        RECT 18.450 114.600 18.620 115.220 ;
        RECT 18.965 115.110 19.505 115.480 ;
        RECT 19.685 115.370 19.905 115.650 ;
        RECT 20.075 115.200 20.245 115.980 ;
        RECT 19.840 115.030 20.245 115.200 ;
        RECT 20.415 115.190 20.765 115.810 ;
        RECT 19.840 114.940 20.010 115.030 ;
        RECT 20.935 115.020 21.145 115.810 ;
        RECT 18.790 114.770 20.010 114.940 ;
        RECT 20.470 114.860 21.145 115.020 ;
        RECT 18.450 114.430 19.250 114.600 ;
        RECT 18.570 113.880 18.900 114.260 ;
        RECT 19.080 114.140 19.250 114.430 ;
        RECT 19.840 114.390 20.010 114.770 ;
        RECT 20.180 114.850 21.145 114.860 ;
        RECT 21.335 115.680 21.595 116.070 ;
        RECT 21.805 115.970 22.135 116.430 ;
        RECT 23.010 116.040 23.865 116.210 ;
        RECT 24.070 116.040 24.565 116.210 ;
        RECT 24.735 116.070 25.065 116.430 ;
        RECT 21.335 114.990 21.505 115.680 ;
        RECT 21.675 115.330 21.845 115.510 ;
        RECT 22.015 115.500 22.805 115.750 ;
        RECT 23.010 115.330 23.180 116.040 ;
        RECT 23.350 115.530 23.705 115.750 ;
        RECT 21.675 115.160 23.365 115.330 ;
        RECT 20.180 114.560 20.640 114.850 ;
        RECT 21.335 114.820 22.835 114.990 ;
        RECT 21.335 114.680 21.505 114.820 ;
        RECT 20.945 114.510 21.505 114.680 ;
        RECT 19.420 113.880 19.670 114.340 ;
        RECT 19.840 114.050 20.710 114.390 ;
        RECT 20.945 114.050 21.115 114.510 ;
        RECT 21.950 114.480 23.025 114.650 ;
        RECT 21.285 113.880 21.655 114.340 ;
        RECT 21.950 114.140 22.120 114.480 ;
        RECT 22.290 113.880 22.620 114.310 ;
        RECT 22.855 114.140 23.025 114.480 ;
        RECT 23.195 114.380 23.365 115.160 ;
        RECT 23.535 114.940 23.705 115.530 ;
        RECT 23.875 115.130 24.225 115.750 ;
        RECT 23.535 114.550 24.000 114.940 ;
        RECT 24.395 114.680 24.565 116.040 ;
        RECT 24.735 114.850 25.195 115.900 ;
        RECT 24.170 114.510 24.565 114.680 ;
        RECT 24.170 114.380 24.340 114.510 ;
        RECT 23.195 114.050 23.875 114.380 ;
        RECT 24.090 114.050 24.340 114.380 ;
        RECT 24.510 113.880 24.760 114.340 ;
        RECT 24.930 114.065 25.255 114.850 ;
        RECT 25.425 114.050 25.595 116.170 ;
        RECT 25.765 116.050 26.095 116.430 ;
        RECT 26.265 115.880 26.520 116.170 ;
        RECT 25.770 115.710 26.520 115.880 ;
        RECT 26.695 115.755 26.955 116.260 ;
        RECT 27.135 116.050 27.465 116.430 ;
        RECT 27.645 115.880 27.815 116.260 ;
        RECT 25.770 114.720 26.000 115.710 ;
        RECT 26.170 114.890 26.520 115.540 ;
        RECT 26.695 114.955 26.865 115.755 ;
        RECT 27.150 115.710 27.815 115.880 ;
        RECT 27.150 115.455 27.320 115.710 ;
        RECT 28.075 115.705 28.365 116.430 ;
        RECT 28.575 115.610 28.805 116.430 ;
        RECT 28.975 115.630 29.305 116.260 ;
        RECT 27.035 115.125 27.320 115.455 ;
        RECT 27.555 115.160 27.885 115.530 ;
        RECT 28.555 115.190 28.885 115.440 ;
        RECT 27.150 114.980 27.320 115.125 ;
        RECT 25.770 114.550 26.520 114.720 ;
        RECT 25.765 113.880 26.095 114.380 ;
        RECT 26.265 114.050 26.520 114.550 ;
        RECT 26.695 114.050 26.965 114.955 ;
        RECT 27.150 114.810 27.815 114.980 ;
        RECT 27.135 113.880 27.465 114.640 ;
        RECT 27.645 114.050 27.815 114.810 ;
        RECT 28.075 113.880 28.365 115.045 ;
        RECT 29.055 115.030 29.305 115.630 ;
        RECT 29.475 115.610 29.685 116.430 ;
        RECT 29.955 115.610 30.185 116.430 ;
        RECT 30.355 115.630 30.685 116.260 ;
        RECT 29.935 115.190 30.265 115.440 ;
        RECT 30.435 115.030 30.685 115.630 ;
        RECT 30.855 115.610 31.065 116.430 ;
        RECT 31.295 115.755 31.555 116.260 ;
        RECT 31.735 116.050 32.065 116.430 ;
        RECT 32.245 115.880 32.415 116.260 ;
        RECT 32.985 115.960 33.155 116.430 ;
        RECT 28.575 113.880 28.805 115.020 ;
        RECT 28.975 114.050 29.305 115.030 ;
        RECT 29.475 113.880 29.685 115.020 ;
        RECT 29.955 113.880 30.185 115.020 ;
        RECT 30.355 114.050 30.685 115.030 ;
        RECT 30.855 113.880 31.065 115.020 ;
        RECT 31.295 114.955 31.465 115.755 ;
        RECT 31.750 115.710 32.415 115.880 ;
        RECT 33.325 115.780 33.655 116.260 ;
        RECT 33.825 115.960 33.995 116.430 ;
        RECT 34.165 115.780 34.495 116.260 ;
        RECT 31.750 115.455 31.920 115.710 ;
        RECT 32.730 115.610 34.495 115.780 ;
        RECT 34.665 115.620 34.835 116.430 ;
        RECT 35.035 116.050 36.105 116.220 ;
        RECT 35.035 115.695 35.355 116.050 ;
        RECT 31.635 115.125 31.920 115.455 ;
        RECT 32.155 115.160 32.485 115.530 ;
        RECT 31.750 114.980 31.920 115.125 ;
        RECT 32.730 115.060 33.140 115.610 ;
        RECT 35.030 115.440 35.355 115.695 ;
        RECT 33.325 115.230 35.355 115.440 ;
        RECT 35.010 115.220 35.355 115.230 ;
        RECT 35.525 115.480 35.765 115.880 ;
        RECT 35.935 115.820 36.105 116.050 ;
        RECT 36.275 115.990 36.465 116.430 ;
        RECT 36.635 115.980 37.585 116.260 ;
        RECT 37.805 116.070 38.155 116.240 ;
        RECT 35.935 115.650 36.465 115.820 ;
        RECT 31.295 114.050 31.565 114.955 ;
        RECT 31.750 114.810 32.415 114.980 ;
        RECT 32.730 114.890 34.455 115.060 ;
        RECT 31.735 113.880 32.065 114.640 ;
        RECT 32.245 114.050 32.415 114.810 ;
        RECT 32.985 113.880 33.155 114.720 ;
        RECT 33.365 114.050 33.615 114.890 ;
        RECT 33.825 113.880 33.995 114.720 ;
        RECT 34.165 114.050 34.455 114.890 ;
        RECT 34.665 113.880 34.835 114.940 ;
        RECT 35.010 114.600 35.180 115.220 ;
        RECT 35.525 115.110 36.065 115.480 ;
        RECT 36.245 115.370 36.465 115.650 ;
        RECT 36.635 115.200 36.805 115.980 ;
        RECT 36.400 115.030 36.805 115.200 ;
        RECT 36.975 115.190 37.325 115.810 ;
        RECT 36.400 114.940 36.570 115.030 ;
        RECT 37.495 115.020 37.705 115.810 ;
        RECT 35.350 114.770 36.570 114.940 ;
        RECT 37.030 114.860 37.705 115.020 ;
        RECT 35.010 114.430 35.810 114.600 ;
        RECT 35.130 113.880 35.460 114.260 ;
        RECT 35.640 114.140 35.810 114.430 ;
        RECT 36.400 114.390 36.570 114.770 ;
        RECT 36.740 114.850 37.705 114.860 ;
        RECT 37.895 115.680 38.155 116.070 ;
        RECT 38.365 115.970 38.695 116.430 ;
        RECT 39.570 116.040 40.425 116.210 ;
        RECT 40.630 116.040 41.125 116.210 ;
        RECT 41.295 116.070 41.625 116.430 ;
        RECT 37.895 114.990 38.065 115.680 ;
        RECT 38.235 115.330 38.405 115.510 ;
        RECT 38.575 115.500 39.365 115.750 ;
        RECT 39.570 115.330 39.740 116.040 ;
        RECT 39.910 115.530 40.265 115.750 ;
        RECT 38.235 115.160 39.925 115.330 ;
        RECT 36.740 114.560 37.200 114.850 ;
        RECT 37.895 114.820 39.395 114.990 ;
        RECT 37.895 114.680 38.065 114.820 ;
        RECT 37.505 114.510 38.065 114.680 ;
        RECT 35.980 113.880 36.230 114.340 ;
        RECT 36.400 114.050 37.270 114.390 ;
        RECT 37.505 114.050 37.675 114.510 ;
        RECT 38.510 114.480 39.585 114.650 ;
        RECT 37.845 113.880 38.215 114.340 ;
        RECT 38.510 114.140 38.680 114.480 ;
        RECT 38.850 113.880 39.180 114.310 ;
        RECT 39.415 114.140 39.585 114.480 ;
        RECT 39.755 114.380 39.925 115.160 ;
        RECT 40.095 114.940 40.265 115.530 ;
        RECT 40.435 115.130 40.785 115.750 ;
        RECT 40.095 114.550 40.560 114.940 ;
        RECT 40.955 114.680 41.125 116.040 ;
        RECT 41.295 114.850 41.755 115.900 ;
        RECT 40.730 114.510 41.125 114.680 ;
        RECT 40.730 114.380 40.900 114.510 ;
        RECT 39.755 114.050 40.435 114.380 ;
        RECT 40.650 114.050 40.900 114.380 ;
        RECT 41.070 113.880 41.320 114.340 ;
        RECT 41.490 114.065 41.815 114.850 ;
        RECT 41.985 114.050 42.155 116.170 ;
        RECT 42.325 116.050 42.655 116.430 ;
        RECT 42.825 115.880 43.080 116.170 ;
        RECT 43.565 115.960 43.735 116.430 ;
        RECT 42.330 115.710 43.080 115.880 ;
        RECT 43.905 115.780 44.235 116.260 ;
        RECT 44.405 115.960 44.575 116.430 ;
        RECT 44.745 115.780 45.075 116.260 ;
        RECT 42.330 114.720 42.560 115.710 ;
        RECT 43.310 115.610 45.075 115.780 ;
        RECT 45.245 115.620 45.415 116.430 ;
        RECT 45.615 116.050 46.685 116.220 ;
        RECT 45.615 115.695 45.935 116.050 ;
        RECT 42.730 114.890 43.080 115.540 ;
        RECT 43.310 115.060 43.720 115.610 ;
        RECT 45.610 115.440 45.935 115.695 ;
        RECT 43.905 115.230 45.935 115.440 ;
        RECT 45.590 115.220 45.935 115.230 ;
        RECT 46.105 115.480 46.345 115.880 ;
        RECT 46.515 115.820 46.685 116.050 ;
        RECT 46.855 115.990 47.045 116.430 ;
        RECT 47.215 115.980 48.165 116.260 ;
        RECT 48.385 116.070 48.735 116.240 ;
        RECT 46.515 115.650 47.045 115.820 ;
        RECT 43.310 114.890 45.035 115.060 ;
        RECT 42.330 114.550 43.080 114.720 ;
        RECT 42.325 113.880 42.655 114.380 ;
        RECT 42.825 114.050 43.080 114.550 ;
        RECT 43.565 113.880 43.735 114.720 ;
        RECT 43.945 114.050 44.195 114.890 ;
        RECT 44.405 113.880 44.575 114.720 ;
        RECT 44.745 114.050 45.035 114.890 ;
        RECT 45.245 113.880 45.415 114.940 ;
        RECT 45.590 114.600 45.760 115.220 ;
        RECT 46.105 115.110 46.645 115.480 ;
        RECT 46.825 115.370 47.045 115.650 ;
        RECT 47.215 115.200 47.385 115.980 ;
        RECT 46.980 115.030 47.385 115.200 ;
        RECT 47.555 115.190 47.905 115.810 ;
        RECT 46.980 114.940 47.150 115.030 ;
        RECT 48.075 115.020 48.285 115.810 ;
        RECT 45.930 114.770 47.150 114.940 ;
        RECT 47.610 114.860 48.285 115.020 ;
        RECT 45.590 114.430 46.390 114.600 ;
        RECT 45.710 113.880 46.040 114.260 ;
        RECT 46.220 114.140 46.390 114.430 ;
        RECT 46.980 114.390 47.150 114.770 ;
        RECT 47.320 114.850 48.285 114.860 ;
        RECT 48.475 115.680 48.735 116.070 ;
        RECT 48.945 115.970 49.275 116.430 ;
        RECT 50.150 116.040 51.005 116.210 ;
        RECT 51.210 116.040 51.705 116.210 ;
        RECT 51.875 116.070 52.205 116.430 ;
        RECT 48.475 114.990 48.645 115.680 ;
        RECT 48.815 115.330 48.985 115.510 ;
        RECT 49.155 115.500 49.945 115.750 ;
        RECT 50.150 115.330 50.320 116.040 ;
        RECT 50.490 115.530 50.845 115.750 ;
        RECT 48.815 115.160 50.505 115.330 ;
        RECT 47.320 114.560 47.780 114.850 ;
        RECT 48.475 114.820 49.975 114.990 ;
        RECT 48.475 114.680 48.645 114.820 ;
        RECT 48.085 114.510 48.645 114.680 ;
        RECT 46.560 113.880 46.810 114.340 ;
        RECT 46.980 114.050 47.850 114.390 ;
        RECT 48.085 114.050 48.255 114.510 ;
        RECT 49.090 114.480 50.165 114.650 ;
        RECT 48.425 113.880 48.795 114.340 ;
        RECT 49.090 114.140 49.260 114.480 ;
        RECT 49.430 113.880 49.760 114.310 ;
        RECT 49.995 114.140 50.165 114.480 ;
        RECT 50.335 114.380 50.505 115.160 ;
        RECT 50.675 114.940 50.845 115.530 ;
        RECT 51.015 115.130 51.365 115.750 ;
        RECT 50.675 114.550 51.140 114.940 ;
        RECT 51.535 114.680 51.705 116.040 ;
        RECT 51.875 114.850 52.335 115.900 ;
        RECT 51.310 114.510 51.705 114.680 ;
        RECT 51.310 114.380 51.480 114.510 ;
        RECT 50.335 114.050 51.015 114.380 ;
        RECT 51.230 114.050 51.480 114.380 ;
        RECT 51.650 113.880 51.900 114.340 ;
        RECT 52.070 114.065 52.395 114.850 ;
        RECT 52.565 114.050 52.735 116.170 ;
        RECT 52.905 116.050 53.235 116.430 ;
        RECT 53.405 115.880 53.660 116.170 ;
        RECT 52.910 115.710 53.660 115.880 ;
        RECT 52.910 114.720 53.140 115.710 ;
        RECT 53.835 115.705 54.125 116.430 ;
        RECT 54.295 115.755 54.555 116.260 ;
        RECT 54.735 116.050 55.065 116.430 ;
        RECT 55.245 115.880 55.415 116.260 ;
        RECT 53.310 114.890 53.660 115.540 ;
        RECT 52.910 114.550 53.660 114.720 ;
        RECT 52.905 113.880 53.235 114.380 ;
        RECT 53.405 114.050 53.660 114.550 ;
        RECT 53.835 113.880 54.125 115.045 ;
        RECT 54.295 114.955 54.465 115.755 ;
        RECT 54.750 115.710 55.415 115.880 ;
        RECT 56.225 115.880 56.395 116.260 ;
        RECT 56.575 116.050 56.905 116.430 ;
        RECT 56.225 115.710 56.890 115.880 ;
        RECT 57.085 115.755 57.345 116.260 ;
        RECT 57.825 115.960 57.995 116.430 ;
        RECT 58.165 115.780 58.495 116.260 ;
        RECT 58.665 115.960 58.835 116.430 ;
        RECT 59.005 115.780 59.335 116.260 ;
        RECT 54.750 115.455 54.920 115.710 ;
        RECT 54.635 115.125 54.920 115.455 ;
        RECT 55.155 115.160 55.485 115.530 ;
        RECT 56.155 115.160 56.485 115.530 ;
        RECT 56.720 115.455 56.890 115.710 ;
        RECT 54.750 114.980 54.920 115.125 ;
        RECT 56.720 115.125 57.005 115.455 ;
        RECT 56.720 114.980 56.890 115.125 ;
        RECT 54.295 114.050 54.565 114.955 ;
        RECT 54.750 114.810 55.415 114.980 ;
        RECT 54.735 113.880 55.065 114.640 ;
        RECT 55.245 114.050 55.415 114.810 ;
        RECT 56.225 114.810 56.890 114.980 ;
        RECT 57.175 114.955 57.345 115.755 ;
        RECT 56.225 114.050 56.395 114.810 ;
        RECT 56.575 113.880 56.905 114.640 ;
        RECT 57.075 114.050 57.345 114.955 ;
        RECT 57.570 115.610 59.335 115.780 ;
        RECT 59.505 115.620 59.675 116.430 ;
        RECT 59.875 116.050 60.945 116.220 ;
        RECT 59.875 115.695 60.195 116.050 ;
        RECT 57.570 115.060 57.980 115.610 ;
        RECT 59.870 115.440 60.195 115.695 ;
        RECT 58.165 115.230 60.195 115.440 ;
        RECT 59.850 115.220 60.195 115.230 ;
        RECT 60.365 115.480 60.605 115.880 ;
        RECT 60.775 115.820 60.945 116.050 ;
        RECT 61.115 115.990 61.305 116.430 ;
        RECT 61.475 115.980 62.425 116.260 ;
        RECT 62.645 116.070 62.995 116.240 ;
        RECT 60.775 115.650 61.305 115.820 ;
        RECT 57.570 114.890 59.295 115.060 ;
        RECT 57.825 113.880 57.995 114.720 ;
        RECT 58.205 114.050 58.455 114.890 ;
        RECT 58.665 113.880 58.835 114.720 ;
        RECT 59.005 114.050 59.295 114.890 ;
        RECT 59.505 113.880 59.675 114.940 ;
        RECT 59.850 114.600 60.020 115.220 ;
        RECT 60.365 115.110 60.905 115.480 ;
        RECT 61.085 115.370 61.305 115.650 ;
        RECT 61.475 115.200 61.645 115.980 ;
        RECT 61.240 115.030 61.645 115.200 ;
        RECT 61.815 115.190 62.165 115.810 ;
        RECT 61.240 114.940 61.410 115.030 ;
        RECT 62.335 115.020 62.545 115.810 ;
        RECT 60.190 114.770 61.410 114.940 ;
        RECT 61.870 114.860 62.545 115.020 ;
        RECT 59.850 114.430 60.650 114.600 ;
        RECT 59.970 113.880 60.300 114.260 ;
        RECT 60.480 114.140 60.650 114.430 ;
        RECT 61.240 114.390 61.410 114.770 ;
        RECT 61.580 114.850 62.545 114.860 ;
        RECT 62.735 115.680 62.995 116.070 ;
        RECT 63.205 115.970 63.535 116.430 ;
        RECT 64.410 116.040 65.265 116.210 ;
        RECT 65.470 116.040 65.965 116.210 ;
        RECT 66.135 116.070 66.465 116.430 ;
        RECT 62.735 114.990 62.905 115.680 ;
        RECT 63.075 115.330 63.245 115.510 ;
        RECT 63.415 115.500 64.205 115.750 ;
        RECT 64.410 115.330 64.580 116.040 ;
        RECT 64.750 115.530 65.105 115.750 ;
        RECT 63.075 115.160 64.765 115.330 ;
        RECT 61.580 114.560 62.040 114.850 ;
        RECT 62.735 114.820 64.235 114.990 ;
        RECT 62.735 114.680 62.905 114.820 ;
        RECT 62.345 114.510 62.905 114.680 ;
        RECT 60.820 113.880 61.070 114.340 ;
        RECT 61.240 114.050 62.110 114.390 ;
        RECT 62.345 114.050 62.515 114.510 ;
        RECT 63.350 114.480 64.425 114.650 ;
        RECT 62.685 113.880 63.055 114.340 ;
        RECT 63.350 114.140 63.520 114.480 ;
        RECT 63.690 113.880 64.020 114.310 ;
        RECT 64.255 114.140 64.425 114.480 ;
        RECT 64.595 114.380 64.765 115.160 ;
        RECT 64.935 114.940 65.105 115.530 ;
        RECT 65.275 115.130 65.625 115.750 ;
        RECT 64.935 114.550 65.400 114.940 ;
        RECT 65.795 114.680 65.965 116.040 ;
        RECT 66.135 114.850 66.595 115.900 ;
        RECT 65.570 114.510 65.965 114.680 ;
        RECT 65.570 114.380 65.740 114.510 ;
        RECT 64.595 114.050 65.275 114.380 ;
        RECT 65.490 114.050 65.740 114.380 ;
        RECT 65.910 113.880 66.160 114.340 ;
        RECT 66.330 114.065 66.655 114.850 ;
        RECT 66.825 114.050 66.995 116.170 ;
        RECT 67.165 116.050 67.495 116.430 ;
        RECT 67.665 115.880 67.920 116.170 ;
        RECT 68.405 115.960 68.575 116.430 ;
        RECT 67.170 115.710 67.920 115.880 ;
        RECT 68.745 115.780 69.075 116.260 ;
        RECT 69.245 115.960 69.415 116.430 ;
        RECT 69.585 115.780 69.915 116.260 ;
        RECT 67.170 114.720 67.400 115.710 ;
        RECT 68.150 115.610 69.915 115.780 ;
        RECT 70.085 115.620 70.255 116.430 ;
        RECT 70.455 116.050 71.525 116.220 ;
        RECT 70.455 115.695 70.775 116.050 ;
        RECT 67.570 114.890 67.920 115.540 ;
        RECT 68.150 115.060 68.560 115.610 ;
        RECT 70.450 115.440 70.775 115.695 ;
        RECT 68.745 115.230 70.775 115.440 ;
        RECT 70.430 115.220 70.775 115.230 ;
        RECT 70.945 115.480 71.185 115.880 ;
        RECT 71.355 115.820 71.525 116.050 ;
        RECT 71.695 115.990 71.885 116.430 ;
        RECT 72.055 115.980 73.005 116.260 ;
        RECT 73.225 116.070 73.575 116.240 ;
        RECT 71.355 115.650 71.885 115.820 ;
        RECT 68.150 114.890 69.875 115.060 ;
        RECT 67.170 114.550 67.920 114.720 ;
        RECT 67.165 113.880 67.495 114.380 ;
        RECT 67.665 114.050 67.920 114.550 ;
        RECT 68.405 113.880 68.575 114.720 ;
        RECT 68.785 114.050 69.035 114.890 ;
        RECT 69.245 113.880 69.415 114.720 ;
        RECT 69.585 114.050 69.875 114.890 ;
        RECT 70.085 113.880 70.255 114.940 ;
        RECT 70.430 114.600 70.600 115.220 ;
        RECT 70.945 115.110 71.485 115.480 ;
        RECT 71.665 115.370 71.885 115.650 ;
        RECT 72.055 115.200 72.225 115.980 ;
        RECT 71.820 115.030 72.225 115.200 ;
        RECT 72.395 115.190 72.745 115.810 ;
        RECT 71.820 114.940 71.990 115.030 ;
        RECT 72.915 115.020 73.125 115.810 ;
        RECT 70.770 114.770 71.990 114.940 ;
        RECT 72.450 114.860 73.125 115.020 ;
        RECT 70.430 114.430 71.230 114.600 ;
        RECT 70.550 113.880 70.880 114.260 ;
        RECT 71.060 114.140 71.230 114.430 ;
        RECT 71.820 114.390 71.990 114.770 ;
        RECT 72.160 114.850 73.125 114.860 ;
        RECT 73.315 115.680 73.575 116.070 ;
        RECT 73.785 115.970 74.115 116.430 ;
        RECT 74.990 116.040 75.845 116.210 ;
        RECT 76.050 116.040 76.545 116.210 ;
        RECT 76.715 116.070 77.045 116.430 ;
        RECT 73.315 114.990 73.485 115.680 ;
        RECT 73.655 115.330 73.825 115.510 ;
        RECT 73.995 115.500 74.785 115.750 ;
        RECT 74.990 115.330 75.160 116.040 ;
        RECT 75.330 115.530 75.685 115.750 ;
        RECT 73.655 115.160 75.345 115.330 ;
        RECT 72.160 114.560 72.620 114.850 ;
        RECT 73.315 114.820 74.815 114.990 ;
        RECT 73.315 114.680 73.485 114.820 ;
        RECT 72.925 114.510 73.485 114.680 ;
        RECT 71.400 113.880 71.650 114.340 ;
        RECT 71.820 114.050 72.690 114.390 ;
        RECT 72.925 114.050 73.095 114.510 ;
        RECT 73.930 114.480 75.005 114.650 ;
        RECT 73.265 113.880 73.635 114.340 ;
        RECT 73.930 114.140 74.100 114.480 ;
        RECT 74.270 113.880 74.600 114.310 ;
        RECT 74.835 114.140 75.005 114.480 ;
        RECT 75.175 114.380 75.345 115.160 ;
        RECT 75.515 114.940 75.685 115.530 ;
        RECT 75.855 115.130 76.205 115.750 ;
        RECT 75.515 114.550 75.980 114.940 ;
        RECT 76.375 114.680 76.545 116.040 ;
        RECT 76.715 114.850 77.175 115.900 ;
        RECT 76.150 114.510 76.545 114.680 ;
        RECT 76.150 114.380 76.320 114.510 ;
        RECT 75.175 114.050 75.855 114.380 ;
        RECT 76.070 114.050 76.320 114.380 ;
        RECT 76.490 113.880 76.740 114.340 ;
        RECT 76.910 114.065 77.235 114.850 ;
        RECT 77.405 114.050 77.575 116.170 ;
        RECT 77.745 116.050 78.075 116.430 ;
        RECT 78.245 115.880 78.500 116.170 ;
        RECT 77.750 115.710 78.500 115.880 ;
        RECT 77.750 114.720 77.980 115.710 ;
        RECT 79.595 115.705 79.885 116.430 ;
        RECT 80.365 115.960 80.535 116.430 ;
        RECT 80.705 115.780 81.035 116.260 ;
        RECT 81.205 115.960 81.375 116.430 ;
        RECT 81.545 115.780 81.875 116.260 ;
        RECT 80.110 115.610 81.875 115.780 ;
        RECT 82.045 115.620 82.215 116.430 ;
        RECT 82.415 116.050 83.485 116.220 ;
        RECT 82.415 115.695 82.735 116.050 ;
        RECT 78.150 114.890 78.500 115.540 ;
        RECT 80.110 115.060 80.520 115.610 ;
        RECT 82.410 115.440 82.735 115.695 ;
        RECT 80.705 115.230 82.735 115.440 ;
        RECT 82.390 115.220 82.735 115.230 ;
        RECT 82.905 115.480 83.145 115.880 ;
        RECT 83.315 115.820 83.485 116.050 ;
        RECT 83.655 115.990 83.845 116.430 ;
        RECT 84.015 115.980 84.965 116.260 ;
        RECT 85.185 116.070 85.535 116.240 ;
        RECT 83.315 115.650 83.845 115.820 ;
        RECT 77.750 114.550 78.500 114.720 ;
        RECT 77.745 113.880 78.075 114.380 ;
        RECT 78.245 114.050 78.500 114.550 ;
        RECT 79.595 113.880 79.885 115.045 ;
        RECT 80.110 114.890 81.835 115.060 ;
        RECT 80.365 113.880 80.535 114.720 ;
        RECT 80.745 114.050 80.995 114.890 ;
        RECT 81.205 113.880 81.375 114.720 ;
        RECT 81.545 114.050 81.835 114.890 ;
        RECT 82.045 113.880 82.215 114.940 ;
        RECT 82.390 114.600 82.560 115.220 ;
        RECT 82.905 115.110 83.445 115.480 ;
        RECT 83.625 115.370 83.845 115.650 ;
        RECT 84.015 115.200 84.185 115.980 ;
        RECT 83.780 115.030 84.185 115.200 ;
        RECT 84.355 115.190 84.705 115.810 ;
        RECT 83.780 114.940 83.950 115.030 ;
        RECT 84.875 115.020 85.085 115.810 ;
        RECT 82.730 114.770 83.950 114.940 ;
        RECT 84.410 114.860 85.085 115.020 ;
        RECT 82.390 114.430 83.190 114.600 ;
        RECT 82.510 113.880 82.840 114.260 ;
        RECT 83.020 114.140 83.190 114.430 ;
        RECT 83.780 114.390 83.950 114.770 ;
        RECT 84.120 114.850 85.085 114.860 ;
        RECT 85.275 115.680 85.535 116.070 ;
        RECT 85.745 115.970 86.075 116.430 ;
        RECT 86.950 116.040 87.805 116.210 ;
        RECT 88.010 116.040 88.505 116.210 ;
        RECT 88.675 116.070 89.005 116.430 ;
        RECT 85.275 114.990 85.445 115.680 ;
        RECT 85.615 115.330 85.785 115.510 ;
        RECT 85.955 115.500 86.745 115.750 ;
        RECT 86.950 115.330 87.120 116.040 ;
        RECT 87.290 115.530 87.645 115.750 ;
        RECT 85.615 115.160 87.305 115.330 ;
        RECT 84.120 114.560 84.580 114.850 ;
        RECT 85.275 114.820 86.775 114.990 ;
        RECT 85.275 114.680 85.445 114.820 ;
        RECT 84.885 114.510 85.445 114.680 ;
        RECT 83.360 113.880 83.610 114.340 ;
        RECT 83.780 114.050 84.650 114.390 ;
        RECT 84.885 114.050 85.055 114.510 ;
        RECT 85.890 114.480 86.965 114.650 ;
        RECT 85.225 113.880 85.595 114.340 ;
        RECT 85.890 114.140 86.060 114.480 ;
        RECT 86.230 113.880 86.560 114.310 ;
        RECT 86.795 114.140 86.965 114.480 ;
        RECT 87.135 114.380 87.305 115.160 ;
        RECT 87.475 114.940 87.645 115.530 ;
        RECT 87.815 115.130 88.165 115.750 ;
        RECT 87.475 114.550 87.940 114.940 ;
        RECT 88.335 114.680 88.505 116.040 ;
        RECT 88.675 114.850 89.135 115.900 ;
        RECT 88.110 114.510 88.505 114.680 ;
        RECT 88.110 114.380 88.280 114.510 ;
        RECT 87.135 114.050 87.815 114.380 ;
        RECT 88.030 114.050 88.280 114.380 ;
        RECT 88.450 113.880 88.700 114.340 ;
        RECT 88.870 114.065 89.195 114.850 ;
        RECT 89.365 114.050 89.535 116.170 ;
        RECT 89.705 116.050 90.035 116.430 ;
        RECT 90.205 115.880 90.460 116.170 ;
        RECT 89.710 115.710 90.460 115.880 ;
        RECT 89.710 114.720 89.940 115.710 ;
        RECT 90.635 115.680 91.845 116.430 ;
        RECT 90.110 114.890 90.460 115.540 ;
        RECT 90.635 114.970 91.155 115.510 ;
        RECT 91.325 115.140 91.845 115.680 ;
        RECT 92.015 115.755 92.275 116.260 ;
        RECT 92.455 116.050 92.785 116.430 ;
        RECT 92.965 115.880 93.135 116.260 ;
        RECT 89.710 114.550 90.460 114.720 ;
        RECT 89.705 113.880 90.035 114.380 ;
        RECT 90.205 114.050 90.460 114.550 ;
        RECT 90.635 113.880 91.845 114.970 ;
        RECT 92.015 114.955 92.185 115.755 ;
        RECT 92.470 115.710 93.135 115.880 ;
        RECT 92.470 115.455 92.640 115.710 ;
        RECT 93.435 115.610 93.665 116.430 ;
        RECT 93.835 115.630 94.165 116.260 ;
        RECT 92.355 115.125 92.640 115.455 ;
        RECT 92.875 115.160 93.205 115.530 ;
        RECT 93.415 115.190 93.745 115.440 ;
        RECT 92.470 114.980 92.640 115.125 ;
        RECT 93.915 115.030 94.165 115.630 ;
        RECT 94.335 115.610 94.545 116.430 ;
        RECT 95.085 115.960 95.255 116.430 ;
        RECT 95.425 115.780 95.755 116.260 ;
        RECT 95.925 115.960 96.095 116.430 ;
        RECT 96.265 115.780 96.595 116.260 ;
        RECT 94.830 115.610 96.595 115.780 ;
        RECT 96.765 115.620 96.935 116.430 ;
        RECT 97.135 116.050 98.205 116.220 ;
        RECT 97.135 115.695 97.455 116.050 ;
        RECT 92.015 114.050 92.285 114.955 ;
        RECT 92.470 114.810 93.135 114.980 ;
        RECT 92.455 113.880 92.785 114.640 ;
        RECT 92.965 114.050 93.135 114.810 ;
        RECT 93.435 113.880 93.665 115.020 ;
        RECT 93.835 114.050 94.165 115.030 ;
        RECT 94.830 115.060 95.240 115.610 ;
        RECT 97.130 115.440 97.455 115.695 ;
        RECT 95.425 115.230 97.455 115.440 ;
        RECT 97.110 115.220 97.455 115.230 ;
        RECT 97.625 115.480 97.865 115.880 ;
        RECT 98.035 115.820 98.205 116.050 ;
        RECT 98.375 115.990 98.565 116.430 ;
        RECT 98.735 115.980 99.685 116.260 ;
        RECT 99.905 116.070 100.255 116.240 ;
        RECT 98.035 115.650 98.565 115.820 ;
        RECT 94.335 113.880 94.545 115.020 ;
        RECT 94.830 114.890 96.555 115.060 ;
        RECT 95.085 113.880 95.255 114.720 ;
        RECT 95.465 114.050 95.715 114.890 ;
        RECT 95.925 113.880 96.095 114.720 ;
        RECT 96.265 114.050 96.555 114.890 ;
        RECT 96.765 113.880 96.935 114.940 ;
        RECT 97.110 114.600 97.280 115.220 ;
        RECT 97.625 115.110 98.165 115.480 ;
        RECT 98.345 115.370 98.565 115.650 ;
        RECT 98.735 115.200 98.905 115.980 ;
        RECT 98.500 115.030 98.905 115.200 ;
        RECT 99.075 115.190 99.425 115.810 ;
        RECT 98.500 114.940 98.670 115.030 ;
        RECT 99.595 115.020 99.805 115.810 ;
        RECT 97.450 114.770 98.670 114.940 ;
        RECT 99.130 114.860 99.805 115.020 ;
        RECT 97.110 114.430 97.910 114.600 ;
        RECT 97.230 113.880 97.560 114.260 ;
        RECT 97.740 114.140 97.910 114.430 ;
        RECT 98.500 114.390 98.670 114.770 ;
        RECT 98.840 114.850 99.805 114.860 ;
        RECT 99.995 115.680 100.255 116.070 ;
        RECT 100.465 115.970 100.795 116.430 ;
        RECT 101.670 116.040 102.525 116.210 ;
        RECT 102.730 116.040 103.225 116.210 ;
        RECT 103.395 116.070 103.725 116.430 ;
        RECT 99.995 114.990 100.165 115.680 ;
        RECT 100.335 115.330 100.505 115.510 ;
        RECT 100.675 115.500 101.465 115.750 ;
        RECT 101.670 115.330 101.840 116.040 ;
        RECT 102.010 115.530 102.365 115.750 ;
        RECT 100.335 115.160 102.025 115.330 ;
        RECT 98.840 114.560 99.300 114.850 ;
        RECT 99.995 114.820 101.495 114.990 ;
        RECT 99.995 114.680 100.165 114.820 ;
        RECT 99.605 114.510 100.165 114.680 ;
        RECT 98.080 113.880 98.330 114.340 ;
        RECT 98.500 114.050 99.370 114.390 ;
        RECT 99.605 114.050 99.775 114.510 ;
        RECT 100.610 114.480 101.685 114.650 ;
        RECT 99.945 113.880 100.315 114.340 ;
        RECT 100.610 114.140 100.780 114.480 ;
        RECT 100.950 113.880 101.280 114.310 ;
        RECT 101.515 114.140 101.685 114.480 ;
        RECT 101.855 114.380 102.025 115.160 ;
        RECT 102.195 114.940 102.365 115.530 ;
        RECT 102.535 115.130 102.885 115.750 ;
        RECT 102.195 114.550 102.660 114.940 ;
        RECT 103.055 114.680 103.225 116.040 ;
        RECT 103.395 114.850 103.855 115.900 ;
        RECT 102.830 114.510 103.225 114.680 ;
        RECT 102.830 114.380 103.000 114.510 ;
        RECT 101.855 114.050 102.535 114.380 ;
        RECT 102.750 114.050 103.000 114.380 ;
        RECT 103.170 113.880 103.420 114.340 ;
        RECT 103.590 114.065 103.915 114.850 ;
        RECT 104.085 114.050 104.255 116.170 ;
        RECT 104.425 116.050 104.755 116.430 ;
        RECT 104.925 115.880 105.180 116.170 ;
        RECT 104.430 115.710 105.180 115.880 ;
        RECT 104.430 114.720 104.660 115.710 ;
        RECT 105.355 115.705 105.645 116.430 ;
        RECT 107.045 115.960 107.215 116.430 ;
        RECT 107.385 115.780 107.715 116.260 ;
        RECT 107.885 115.960 108.055 116.430 ;
        RECT 108.225 115.780 108.555 116.260 ;
        RECT 106.790 115.610 108.555 115.780 ;
        RECT 108.725 115.620 108.895 116.430 ;
        RECT 109.095 116.050 110.165 116.220 ;
        RECT 109.095 115.695 109.415 116.050 ;
        RECT 104.830 114.890 105.180 115.540 ;
        RECT 106.790 115.060 107.200 115.610 ;
        RECT 109.090 115.440 109.415 115.695 ;
        RECT 107.385 115.230 109.415 115.440 ;
        RECT 109.070 115.220 109.415 115.230 ;
        RECT 109.585 115.480 109.825 115.880 ;
        RECT 109.995 115.820 110.165 116.050 ;
        RECT 110.335 115.990 110.525 116.430 ;
        RECT 110.695 115.980 111.645 116.260 ;
        RECT 111.865 116.070 112.215 116.240 ;
        RECT 109.995 115.650 110.525 115.820 ;
        RECT 104.430 114.550 105.180 114.720 ;
        RECT 104.425 113.880 104.755 114.380 ;
        RECT 104.925 114.050 105.180 114.550 ;
        RECT 105.355 113.880 105.645 115.045 ;
        RECT 106.790 114.890 108.515 115.060 ;
        RECT 107.045 113.880 107.215 114.720 ;
        RECT 107.425 114.050 107.675 114.890 ;
        RECT 107.885 113.880 108.055 114.720 ;
        RECT 108.225 114.050 108.515 114.890 ;
        RECT 108.725 113.880 108.895 114.940 ;
        RECT 109.070 114.600 109.240 115.220 ;
        RECT 109.585 115.110 110.125 115.480 ;
        RECT 110.305 115.370 110.525 115.650 ;
        RECT 110.695 115.200 110.865 115.980 ;
        RECT 110.460 115.030 110.865 115.200 ;
        RECT 111.035 115.190 111.385 115.810 ;
        RECT 110.460 114.940 110.630 115.030 ;
        RECT 111.555 115.020 111.765 115.810 ;
        RECT 109.410 114.770 110.630 114.940 ;
        RECT 111.090 114.860 111.765 115.020 ;
        RECT 109.070 114.430 109.870 114.600 ;
        RECT 109.190 113.880 109.520 114.260 ;
        RECT 109.700 114.140 109.870 114.430 ;
        RECT 110.460 114.390 110.630 114.770 ;
        RECT 110.800 114.850 111.765 114.860 ;
        RECT 111.955 115.680 112.215 116.070 ;
        RECT 112.425 115.970 112.755 116.430 ;
        RECT 113.630 116.040 114.485 116.210 ;
        RECT 114.690 116.040 115.185 116.210 ;
        RECT 115.355 116.070 115.685 116.430 ;
        RECT 111.955 114.990 112.125 115.680 ;
        RECT 112.295 115.330 112.465 115.510 ;
        RECT 112.635 115.500 113.425 115.750 ;
        RECT 113.630 115.330 113.800 116.040 ;
        RECT 113.970 115.530 114.325 115.750 ;
        RECT 112.295 115.160 113.985 115.330 ;
        RECT 110.800 114.560 111.260 114.850 ;
        RECT 111.955 114.820 113.455 114.990 ;
        RECT 111.955 114.680 112.125 114.820 ;
        RECT 111.565 114.510 112.125 114.680 ;
        RECT 110.040 113.880 110.290 114.340 ;
        RECT 110.460 114.050 111.330 114.390 ;
        RECT 111.565 114.050 111.735 114.510 ;
        RECT 112.570 114.480 113.645 114.650 ;
        RECT 111.905 113.880 112.275 114.340 ;
        RECT 112.570 114.140 112.740 114.480 ;
        RECT 112.910 113.880 113.240 114.310 ;
        RECT 113.475 114.140 113.645 114.480 ;
        RECT 113.815 114.380 113.985 115.160 ;
        RECT 114.155 114.940 114.325 115.530 ;
        RECT 114.495 115.130 114.845 115.750 ;
        RECT 114.155 114.550 114.620 114.940 ;
        RECT 115.015 114.680 115.185 116.040 ;
        RECT 115.355 114.850 115.815 115.900 ;
        RECT 114.790 114.510 115.185 114.680 ;
        RECT 114.790 114.380 114.960 114.510 ;
        RECT 113.815 114.050 114.495 114.380 ;
        RECT 114.710 114.050 114.960 114.380 ;
        RECT 115.130 113.880 115.380 114.340 ;
        RECT 115.550 114.065 115.875 114.850 ;
        RECT 116.045 114.050 116.215 116.170 ;
        RECT 116.385 116.050 116.715 116.430 ;
        RECT 116.885 115.880 117.140 116.170 ;
        RECT 116.390 115.710 117.140 115.880 ;
        RECT 116.390 114.720 116.620 115.710 ;
        RECT 117.315 115.680 118.525 116.430 ;
        RECT 116.790 114.890 117.140 115.540 ;
        RECT 117.315 114.970 117.835 115.510 ;
        RECT 118.005 115.140 118.525 115.680 ;
        RECT 116.390 114.550 117.140 114.720 ;
        RECT 116.385 113.880 116.715 114.380 ;
        RECT 116.885 114.050 117.140 114.550 ;
        RECT 117.315 113.880 118.525 114.970 ;
        RECT 11.430 113.710 118.610 113.880 ;
        RECT 11.515 112.620 12.725 113.710 ;
        RECT 11.515 111.910 12.035 112.450 ;
        RECT 12.205 112.080 12.725 112.620 ;
        RECT 13.875 112.570 14.085 113.710 ;
        RECT 14.255 112.560 14.585 113.540 ;
        RECT 14.755 112.570 14.985 113.710 ;
        RECT 11.515 111.160 12.725 111.910 ;
        RECT 13.875 111.160 14.085 111.980 ;
        RECT 14.255 111.960 14.505 112.560 ;
        RECT 15.195 112.545 15.485 113.710 ;
        RECT 15.695 112.570 15.925 113.710 ;
        RECT 16.095 112.560 16.425 113.540 ;
        RECT 16.595 112.570 16.805 113.710 ;
        RECT 17.345 112.870 17.515 113.710 ;
        RECT 17.725 112.700 17.975 113.540 ;
        RECT 18.185 112.870 18.355 113.710 ;
        RECT 18.525 112.700 18.815 113.540 ;
        RECT 14.675 112.150 15.005 112.400 ;
        RECT 15.675 112.150 16.005 112.400 ;
        RECT 14.255 111.330 14.585 111.960 ;
        RECT 14.755 111.160 14.985 111.980 ;
        RECT 15.195 111.160 15.485 111.885 ;
        RECT 15.695 111.160 15.925 111.980 ;
        RECT 16.175 111.960 16.425 112.560 ;
        RECT 17.090 112.530 18.815 112.700 ;
        RECT 19.025 112.650 19.195 113.710 ;
        RECT 19.490 113.330 19.820 113.710 ;
        RECT 20.000 113.160 20.170 113.450 ;
        RECT 20.340 113.250 20.590 113.710 ;
        RECT 19.370 112.990 20.170 113.160 ;
        RECT 20.760 113.200 21.630 113.540 ;
        RECT 17.090 111.980 17.500 112.530 ;
        RECT 19.370 112.370 19.540 112.990 ;
        RECT 20.760 112.820 20.930 113.200 ;
        RECT 21.865 113.080 22.035 113.540 ;
        RECT 22.205 113.250 22.575 113.710 ;
        RECT 22.870 113.110 23.040 113.450 ;
        RECT 23.210 113.280 23.540 113.710 ;
        RECT 23.775 113.110 23.945 113.450 ;
        RECT 19.710 112.650 20.930 112.820 ;
        RECT 21.100 112.740 21.560 113.030 ;
        RECT 21.865 112.910 22.425 113.080 ;
        RECT 22.870 112.940 23.945 113.110 ;
        RECT 24.115 113.210 24.795 113.540 ;
        RECT 25.010 113.210 25.260 113.540 ;
        RECT 25.430 113.250 25.680 113.710 ;
        RECT 22.255 112.770 22.425 112.910 ;
        RECT 21.100 112.730 22.065 112.740 ;
        RECT 20.760 112.560 20.930 112.650 ;
        RECT 21.390 112.570 22.065 112.730 ;
        RECT 19.370 112.360 19.715 112.370 ;
        RECT 17.685 112.150 19.715 112.360 ;
        RECT 16.095 111.330 16.425 111.960 ;
        RECT 16.595 111.160 16.805 111.980 ;
        RECT 17.090 111.810 18.855 111.980 ;
        RECT 17.345 111.160 17.515 111.630 ;
        RECT 17.685 111.330 18.015 111.810 ;
        RECT 18.185 111.160 18.355 111.630 ;
        RECT 18.525 111.330 18.855 111.810 ;
        RECT 19.025 111.160 19.195 111.970 ;
        RECT 19.390 111.895 19.715 112.150 ;
        RECT 19.395 111.540 19.715 111.895 ;
        RECT 19.885 112.110 20.425 112.480 ;
        RECT 20.760 112.390 21.165 112.560 ;
        RECT 19.885 111.710 20.125 112.110 ;
        RECT 20.605 111.940 20.825 112.220 ;
        RECT 20.295 111.770 20.825 111.940 ;
        RECT 20.295 111.540 20.465 111.770 ;
        RECT 20.995 111.610 21.165 112.390 ;
        RECT 21.335 111.780 21.685 112.400 ;
        RECT 21.855 111.780 22.065 112.570 ;
        RECT 22.255 112.600 23.755 112.770 ;
        RECT 22.255 111.910 22.425 112.600 ;
        RECT 24.115 112.430 24.285 113.210 ;
        RECT 25.090 113.080 25.260 113.210 ;
        RECT 22.595 112.260 24.285 112.430 ;
        RECT 24.455 112.650 24.920 113.040 ;
        RECT 25.090 112.910 25.485 113.080 ;
        RECT 22.595 112.080 22.765 112.260 ;
        RECT 19.395 111.370 20.465 111.540 ;
        RECT 20.635 111.160 20.825 111.600 ;
        RECT 20.995 111.330 21.945 111.610 ;
        RECT 22.255 111.520 22.515 111.910 ;
        RECT 22.935 111.840 23.725 112.090 ;
        RECT 22.165 111.350 22.515 111.520 ;
        RECT 22.725 111.160 23.055 111.620 ;
        RECT 23.930 111.550 24.100 112.260 ;
        RECT 24.455 112.060 24.625 112.650 ;
        RECT 24.270 111.840 24.625 112.060 ;
        RECT 24.795 111.840 25.145 112.460 ;
        RECT 25.315 111.550 25.485 112.910 ;
        RECT 25.850 112.740 26.175 113.525 ;
        RECT 25.655 111.690 26.115 112.740 ;
        RECT 23.930 111.380 24.785 111.550 ;
        RECT 24.990 111.380 25.485 111.550 ;
        RECT 25.655 111.160 25.985 111.520 ;
        RECT 26.345 111.420 26.515 113.540 ;
        RECT 26.685 113.210 27.015 113.710 ;
        RECT 27.185 113.040 27.440 113.540 ;
        RECT 26.690 112.870 27.440 113.040 ;
        RECT 27.925 112.870 28.095 113.710 ;
        RECT 26.690 111.880 26.920 112.870 ;
        RECT 28.305 112.700 28.555 113.540 ;
        RECT 28.765 112.870 28.935 113.710 ;
        RECT 29.105 112.700 29.395 113.540 ;
        RECT 27.090 112.050 27.440 112.700 ;
        RECT 27.670 112.530 29.395 112.700 ;
        RECT 29.605 112.650 29.775 113.710 ;
        RECT 30.070 113.330 30.400 113.710 ;
        RECT 30.580 113.160 30.750 113.450 ;
        RECT 30.920 113.250 31.170 113.710 ;
        RECT 29.950 112.990 30.750 113.160 ;
        RECT 31.340 113.200 32.210 113.540 ;
        RECT 27.670 111.980 28.080 112.530 ;
        RECT 29.950 112.370 30.120 112.990 ;
        RECT 31.340 112.820 31.510 113.200 ;
        RECT 32.445 113.080 32.615 113.540 ;
        RECT 32.785 113.250 33.155 113.710 ;
        RECT 33.450 113.110 33.620 113.450 ;
        RECT 33.790 113.280 34.120 113.710 ;
        RECT 34.355 113.110 34.525 113.450 ;
        RECT 30.290 112.650 31.510 112.820 ;
        RECT 31.680 112.740 32.140 113.030 ;
        RECT 32.445 112.910 33.005 113.080 ;
        RECT 33.450 112.940 34.525 113.110 ;
        RECT 34.695 113.210 35.375 113.540 ;
        RECT 35.590 113.210 35.840 113.540 ;
        RECT 36.010 113.250 36.260 113.710 ;
        RECT 32.835 112.770 33.005 112.910 ;
        RECT 31.680 112.730 32.645 112.740 ;
        RECT 31.340 112.560 31.510 112.650 ;
        RECT 31.970 112.570 32.645 112.730 ;
        RECT 29.950 112.360 30.295 112.370 ;
        RECT 28.265 112.150 30.295 112.360 ;
        RECT 26.690 111.710 27.440 111.880 ;
        RECT 27.670 111.810 29.435 111.980 ;
        RECT 26.685 111.160 27.015 111.540 ;
        RECT 27.185 111.420 27.440 111.710 ;
        RECT 27.925 111.160 28.095 111.630 ;
        RECT 28.265 111.330 28.595 111.810 ;
        RECT 28.765 111.160 28.935 111.630 ;
        RECT 29.105 111.330 29.435 111.810 ;
        RECT 29.605 111.160 29.775 111.970 ;
        RECT 29.970 111.895 30.295 112.150 ;
        RECT 29.975 111.540 30.295 111.895 ;
        RECT 30.465 112.110 31.005 112.480 ;
        RECT 31.340 112.390 31.745 112.560 ;
        RECT 30.465 111.710 30.705 112.110 ;
        RECT 31.185 111.940 31.405 112.220 ;
        RECT 30.875 111.770 31.405 111.940 ;
        RECT 30.875 111.540 31.045 111.770 ;
        RECT 31.575 111.610 31.745 112.390 ;
        RECT 31.915 111.780 32.265 112.400 ;
        RECT 32.435 111.780 32.645 112.570 ;
        RECT 32.835 112.600 34.335 112.770 ;
        RECT 32.835 111.910 33.005 112.600 ;
        RECT 34.695 112.430 34.865 113.210 ;
        RECT 35.670 113.080 35.840 113.210 ;
        RECT 33.175 112.260 34.865 112.430 ;
        RECT 35.035 112.650 35.500 113.040 ;
        RECT 35.670 112.910 36.065 113.080 ;
        RECT 33.175 112.080 33.345 112.260 ;
        RECT 29.975 111.370 31.045 111.540 ;
        RECT 31.215 111.160 31.405 111.600 ;
        RECT 31.575 111.330 32.525 111.610 ;
        RECT 32.835 111.520 33.095 111.910 ;
        RECT 33.515 111.840 34.305 112.090 ;
        RECT 32.745 111.350 33.095 111.520 ;
        RECT 33.305 111.160 33.635 111.620 ;
        RECT 34.510 111.550 34.680 112.260 ;
        RECT 35.035 112.060 35.205 112.650 ;
        RECT 34.850 111.840 35.205 112.060 ;
        RECT 35.375 111.840 35.725 112.460 ;
        RECT 35.895 111.550 36.065 112.910 ;
        RECT 36.430 112.740 36.755 113.525 ;
        RECT 36.235 111.690 36.695 112.740 ;
        RECT 34.510 111.380 35.365 111.550 ;
        RECT 35.570 111.380 36.065 111.550 ;
        RECT 36.235 111.160 36.565 111.520 ;
        RECT 36.925 111.420 37.095 113.540 ;
        RECT 37.265 113.210 37.595 113.710 ;
        RECT 37.765 113.040 38.020 113.540 ;
        RECT 37.270 112.870 38.020 113.040 ;
        RECT 37.270 111.880 37.500 112.870 ;
        RECT 37.670 112.050 38.020 112.700 ;
        RECT 38.255 112.570 38.465 113.710 ;
        RECT 38.635 112.560 38.965 113.540 ;
        RECT 39.135 112.570 39.365 113.710 ;
        RECT 39.575 112.635 39.845 113.540 ;
        RECT 40.015 112.950 40.345 113.710 ;
        RECT 40.525 112.780 40.695 113.540 ;
        RECT 37.270 111.710 38.020 111.880 ;
        RECT 37.265 111.160 37.595 111.540 ;
        RECT 37.765 111.420 38.020 111.710 ;
        RECT 38.255 111.160 38.465 111.980 ;
        RECT 38.635 111.960 38.885 112.560 ;
        RECT 39.055 112.150 39.385 112.400 ;
        RECT 38.635 111.330 38.965 111.960 ;
        RECT 39.135 111.160 39.365 111.980 ;
        RECT 39.575 111.835 39.745 112.635 ;
        RECT 40.030 112.610 40.695 112.780 ;
        RECT 40.030 112.465 40.200 112.610 ;
        RECT 40.955 112.545 41.245 113.710 ;
        RECT 41.875 112.620 43.545 113.710 ;
        RECT 44.025 112.870 44.195 113.710 ;
        RECT 44.405 112.700 44.655 113.540 ;
        RECT 44.865 112.870 45.035 113.710 ;
        RECT 45.205 112.700 45.495 113.540 ;
        RECT 39.915 112.135 40.200 112.465 ;
        RECT 40.030 111.880 40.200 112.135 ;
        RECT 40.435 112.060 40.765 112.430 ;
        RECT 41.875 112.100 42.625 112.620 ;
        RECT 43.770 112.530 45.495 112.700 ;
        RECT 45.705 112.650 45.875 113.710 ;
        RECT 46.170 113.330 46.500 113.710 ;
        RECT 46.680 113.160 46.850 113.450 ;
        RECT 47.020 113.250 47.270 113.710 ;
        RECT 46.050 112.990 46.850 113.160 ;
        RECT 47.440 113.200 48.310 113.540 ;
        RECT 42.795 111.930 43.545 112.450 ;
        RECT 39.575 111.330 39.835 111.835 ;
        RECT 40.030 111.710 40.695 111.880 ;
        RECT 40.015 111.160 40.345 111.540 ;
        RECT 40.525 111.330 40.695 111.710 ;
        RECT 40.955 111.160 41.245 111.885 ;
        RECT 41.875 111.160 43.545 111.930 ;
        RECT 43.770 111.980 44.180 112.530 ;
        RECT 46.050 112.370 46.220 112.990 ;
        RECT 47.440 112.820 47.610 113.200 ;
        RECT 48.545 113.080 48.715 113.540 ;
        RECT 48.885 113.250 49.255 113.710 ;
        RECT 49.550 113.110 49.720 113.450 ;
        RECT 49.890 113.280 50.220 113.710 ;
        RECT 50.455 113.110 50.625 113.450 ;
        RECT 46.390 112.650 47.610 112.820 ;
        RECT 47.780 112.740 48.240 113.030 ;
        RECT 48.545 112.910 49.105 113.080 ;
        RECT 49.550 112.940 50.625 113.110 ;
        RECT 50.795 113.210 51.475 113.540 ;
        RECT 51.690 113.210 51.940 113.540 ;
        RECT 52.110 113.250 52.360 113.710 ;
        RECT 48.935 112.770 49.105 112.910 ;
        RECT 47.780 112.730 48.745 112.740 ;
        RECT 47.440 112.560 47.610 112.650 ;
        RECT 48.070 112.570 48.745 112.730 ;
        RECT 46.050 112.360 46.395 112.370 ;
        RECT 44.365 112.150 46.395 112.360 ;
        RECT 43.770 111.810 45.535 111.980 ;
        RECT 44.025 111.160 44.195 111.630 ;
        RECT 44.365 111.330 44.695 111.810 ;
        RECT 44.865 111.160 45.035 111.630 ;
        RECT 45.205 111.330 45.535 111.810 ;
        RECT 45.705 111.160 45.875 111.970 ;
        RECT 46.070 111.895 46.395 112.150 ;
        RECT 46.075 111.540 46.395 111.895 ;
        RECT 46.565 112.110 47.105 112.480 ;
        RECT 47.440 112.390 47.845 112.560 ;
        RECT 46.565 111.710 46.805 112.110 ;
        RECT 47.285 111.940 47.505 112.220 ;
        RECT 46.975 111.770 47.505 111.940 ;
        RECT 46.975 111.540 47.145 111.770 ;
        RECT 47.675 111.610 47.845 112.390 ;
        RECT 48.015 111.780 48.365 112.400 ;
        RECT 48.535 111.780 48.745 112.570 ;
        RECT 48.935 112.600 50.435 112.770 ;
        RECT 48.935 111.910 49.105 112.600 ;
        RECT 50.795 112.430 50.965 113.210 ;
        RECT 51.770 113.080 51.940 113.210 ;
        RECT 49.275 112.260 50.965 112.430 ;
        RECT 51.135 112.650 51.600 113.040 ;
        RECT 51.770 112.910 52.165 113.080 ;
        RECT 49.275 112.080 49.445 112.260 ;
        RECT 46.075 111.370 47.145 111.540 ;
        RECT 47.315 111.160 47.505 111.600 ;
        RECT 47.675 111.330 48.625 111.610 ;
        RECT 48.935 111.520 49.195 111.910 ;
        RECT 49.615 111.840 50.405 112.090 ;
        RECT 48.845 111.350 49.195 111.520 ;
        RECT 49.405 111.160 49.735 111.620 ;
        RECT 50.610 111.550 50.780 112.260 ;
        RECT 51.135 112.060 51.305 112.650 ;
        RECT 50.950 111.840 51.305 112.060 ;
        RECT 51.475 111.840 51.825 112.460 ;
        RECT 51.995 111.550 52.165 112.910 ;
        RECT 52.530 112.740 52.855 113.525 ;
        RECT 52.335 111.690 52.795 112.740 ;
        RECT 50.610 111.380 51.465 111.550 ;
        RECT 51.670 111.380 52.165 111.550 ;
        RECT 52.335 111.160 52.665 111.520 ;
        RECT 53.025 111.420 53.195 113.540 ;
        RECT 53.365 113.210 53.695 113.710 ;
        RECT 53.865 113.040 54.120 113.540 ;
        RECT 53.370 112.870 54.120 113.040 ;
        RECT 54.605 112.870 54.775 113.710 ;
        RECT 53.370 111.880 53.600 112.870 ;
        RECT 54.985 112.700 55.235 113.540 ;
        RECT 55.445 112.870 55.615 113.710 ;
        RECT 55.785 112.700 56.075 113.540 ;
        RECT 53.770 112.050 54.120 112.700 ;
        RECT 54.350 112.530 56.075 112.700 ;
        RECT 56.285 112.650 56.455 113.710 ;
        RECT 56.750 113.330 57.080 113.710 ;
        RECT 57.260 113.160 57.430 113.450 ;
        RECT 57.600 113.250 57.850 113.710 ;
        RECT 56.630 112.990 57.430 113.160 ;
        RECT 58.020 113.200 58.890 113.540 ;
        RECT 54.350 111.980 54.760 112.530 ;
        RECT 56.630 112.370 56.800 112.990 ;
        RECT 58.020 112.820 58.190 113.200 ;
        RECT 59.125 113.080 59.295 113.540 ;
        RECT 59.465 113.250 59.835 113.710 ;
        RECT 60.130 113.110 60.300 113.450 ;
        RECT 60.470 113.280 60.800 113.710 ;
        RECT 61.035 113.110 61.205 113.450 ;
        RECT 56.970 112.650 58.190 112.820 ;
        RECT 58.360 112.740 58.820 113.030 ;
        RECT 59.125 112.910 59.685 113.080 ;
        RECT 60.130 112.940 61.205 113.110 ;
        RECT 61.375 113.210 62.055 113.540 ;
        RECT 62.270 113.210 62.520 113.540 ;
        RECT 62.690 113.250 62.940 113.710 ;
        RECT 59.515 112.770 59.685 112.910 ;
        RECT 58.360 112.730 59.325 112.740 ;
        RECT 58.020 112.560 58.190 112.650 ;
        RECT 58.650 112.570 59.325 112.730 ;
        RECT 56.630 112.360 56.975 112.370 ;
        RECT 54.945 112.150 56.975 112.360 ;
        RECT 53.370 111.710 54.120 111.880 ;
        RECT 54.350 111.810 56.115 111.980 ;
        RECT 53.365 111.160 53.695 111.540 ;
        RECT 53.865 111.420 54.120 111.710 ;
        RECT 54.605 111.160 54.775 111.630 ;
        RECT 54.945 111.330 55.275 111.810 ;
        RECT 55.445 111.160 55.615 111.630 ;
        RECT 55.785 111.330 56.115 111.810 ;
        RECT 56.285 111.160 56.455 111.970 ;
        RECT 56.650 111.895 56.975 112.150 ;
        RECT 56.655 111.540 56.975 111.895 ;
        RECT 57.145 112.110 57.685 112.480 ;
        RECT 58.020 112.390 58.425 112.560 ;
        RECT 57.145 111.710 57.385 112.110 ;
        RECT 57.865 111.940 58.085 112.220 ;
        RECT 57.555 111.770 58.085 111.940 ;
        RECT 57.555 111.540 57.725 111.770 ;
        RECT 58.255 111.610 58.425 112.390 ;
        RECT 58.595 111.780 58.945 112.400 ;
        RECT 59.115 111.780 59.325 112.570 ;
        RECT 59.515 112.600 61.015 112.770 ;
        RECT 59.515 111.910 59.685 112.600 ;
        RECT 61.375 112.430 61.545 113.210 ;
        RECT 62.350 113.080 62.520 113.210 ;
        RECT 59.855 112.260 61.545 112.430 ;
        RECT 61.715 112.650 62.180 113.040 ;
        RECT 62.350 112.910 62.745 113.080 ;
        RECT 59.855 112.080 60.025 112.260 ;
        RECT 56.655 111.370 57.725 111.540 ;
        RECT 57.895 111.160 58.085 111.600 ;
        RECT 58.255 111.330 59.205 111.610 ;
        RECT 59.515 111.520 59.775 111.910 ;
        RECT 60.195 111.840 60.985 112.090 ;
        RECT 59.425 111.350 59.775 111.520 ;
        RECT 59.985 111.160 60.315 111.620 ;
        RECT 61.190 111.550 61.360 112.260 ;
        RECT 61.715 112.060 61.885 112.650 ;
        RECT 61.530 111.840 61.885 112.060 ;
        RECT 62.055 111.840 62.405 112.460 ;
        RECT 62.575 111.550 62.745 112.910 ;
        RECT 63.110 112.740 63.435 113.525 ;
        RECT 62.915 111.690 63.375 112.740 ;
        RECT 61.190 111.380 62.045 111.550 ;
        RECT 62.250 111.380 62.745 111.550 ;
        RECT 62.915 111.160 63.245 111.520 ;
        RECT 63.605 111.420 63.775 113.540 ;
        RECT 63.945 113.210 64.275 113.710 ;
        RECT 64.445 113.040 64.700 113.540 ;
        RECT 63.950 112.870 64.700 113.040 ;
        RECT 63.950 111.880 64.180 112.870 ;
        RECT 64.350 112.050 64.700 112.700 ;
        RECT 64.875 112.620 66.545 113.710 ;
        RECT 64.875 112.100 65.625 112.620 ;
        RECT 66.715 112.545 67.005 113.710 ;
        RECT 67.945 112.870 68.115 113.710 ;
        RECT 68.325 112.700 68.575 113.540 ;
        RECT 68.785 112.870 68.955 113.710 ;
        RECT 69.125 112.700 69.415 113.540 ;
        RECT 67.690 112.530 69.415 112.700 ;
        RECT 69.625 112.650 69.795 113.710 ;
        RECT 70.090 113.330 70.420 113.710 ;
        RECT 70.600 113.160 70.770 113.450 ;
        RECT 70.940 113.250 71.190 113.710 ;
        RECT 69.970 112.990 70.770 113.160 ;
        RECT 71.360 113.200 72.230 113.540 ;
        RECT 65.795 111.930 66.545 112.450 ;
        RECT 63.950 111.710 64.700 111.880 ;
        RECT 63.945 111.160 64.275 111.540 ;
        RECT 64.445 111.420 64.700 111.710 ;
        RECT 64.875 111.160 66.545 111.930 ;
        RECT 67.690 111.980 68.100 112.530 ;
        RECT 69.970 112.370 70.140 112.990 ;
        RECT 71.360 112.820 71.530 113.200 ;
        RECT 72.465 113.080 72.635 113.540 ;
        RECT 72.805 113.250 73.175 113.710 ;
        RECT 73.470 113.110 73.640 113.450 ;
        RECT 73.810 113.280 74.140 113.710 ;
        RECT 74.375 113.110 74.545 113.450 ;
        RECT 70.310 112.650 71.530 112.820 ;
        RECT 71.700 112.740 72.160 113.030 ;
        RECT 72.465 112.910 73.025 113.080 ;
        RECT 73.470 112.940 74.545 113.110 ;
        RECT 74.715 113.210 75.395 113.540 ;
        RECT 75.610 113.210 75.860 113.540 ;
        RECT 76.030 113.250 76.280 113.710 ;
        RECT 72.855 112.770 73.025 112.910 ;
        RECT 71.700 112.730 72.665 112.740 ;
        RECT 71.360 112.560 71.530 112.650 ;
        RECT 71.990 112.570 72.665 112.730 ;
        RECT 69.970 112.360 70.315 112.370 ;
        RECT 68.285 112.150 70.315 112.360 ;
        RECT 66.715 111.160 67.005 111.885 ;
        RECT 67.690 111.810 69.455 111.980 ;
        RECT 67.945 111.160 68.115 111.630 ;
        RECT 68.285 111.330 68.615 111.810 ;
        RECT 68.785 111.160 68.955 111.630 ;
        RECT 69.125 111.330 69.455 111.810 ;
        RECT 69.625 111.160 69.795 111.970 ;
        RECT 69.990 111.895 70.315 112.150 ;
        RECT 69.995 111.540 70.315 111.895 ;
        RECT 70.485 112.110 71.025 112.480 ;
        RECT 71.360 112.390 71.765 112.560 ;
        RECT 70.485 111.710 70.725 112.110 ;
        RECT 71.205 111.940 71.425 112.220 ;
        RECT 70.895 111.770 71.425 111.940 ;
        RECT 70.895 111.540 71.065 111.770 ;
        RECT 71.595 111.610 71.765 112.390 ;
        RECT 71.935 111.780 72.285 112.400 ;
        RECT 72.455 111.780 72.665 112.570 ;
        RECT 72.855 112.600 74.355 112.770 ;
        RECT 72.855 111.910 73.025 112.600 ;
        RECT 74.715 112.430 74.885 113.210 ;
        RECT 75.690 113.080 75.860 113.210 ;
        RECT 73.195 112.260 74.885 112.430 ;
        RECT 75.055 112.650 75.520 113.040 ;
        RECT 75.690 112.910 76.085 113.080 ;
        RECT 73.195 112.080 73.365 112.260 ;
        RECT 69.995 111.370 71.065 111.540 ;
        RECT 71.235 111.160 71.425 111.600 ;
        RECT 71.595 111.330 72.545 111.610 ;
        RECT 72.855 111.520 73.115 111.910 ;
        RECT 73.535 111.840 74.325 112.090 ;
        RECT 72.765 111.350 73.115 111.520 ;
        RECT 73.325 111.160 73.655 111.620 ;
        RECT 74.530 111.550 74.700 112.260 ;
        RECT 75.055 112.060 75.225 112.650 ;
        RECT 74.870 111.840 75.225 112.060 ;
        RECT 75.395 111.840 75.745 112.460 ;
        RECT 75.915 111.550 76.085 112.910 ;
        RECT 76.450 112.740 76.775 113.525 ;
        RECT 76.255 111.690 76.715 112.740 ;
        RECT 74.530 111.380 75.385 111.550 ;
        RECT 75.590 111.380 76.085 111.550 ;
        RECT 76.255 111.160 76.585 111.520 ;
        RECT 76.945 111.420 77.115 113.540 ;
        RECT 77.285 113.210 77.615 113.710 ;
        RECT 77.785 113.040 78.040 113.540 ;
        RECT 77.290 112.870 78.040 113.040 ;
        RECT 78.525 112.870 78.695 113.710 ;
        RECT 77.290 111.880 77.520 112.870 ;
        RECT 78.905 112.700 79.155 113.540 ;
        RECT 79.365 112.870 79.535 113.710 ;
        RECT 79.705 112.700 79.995 113.540 ;
        RECT 77.690 112.050 78.040 112.700 ;
        RECT 78.270 112.530 79.995 112.700 ;
        RECT 80.205 112.650 80.375 113.710 ;
        RECT 80.670 113.330 81.000 113.710 ;
        RECT 81.180 113.160 81.350 113.450 ;
        RECT 81.520 113.250 81.770 113.710 ;
        RECT 80.550 112.990 81.350 113.160 ;
        RECT 81.940 113.200 82.810 113.540 ;
        RECT 78.270 111.980 78.680 112.530 ;
        RECT 80.550 112.370 80.720 112.990 ;
        RECT 81.940 112.820 82.110 113.200 ;
        RECT 83.045 113.080 83.215 113.540 ;
        RECT 83.385 113.250 83.755 113.710 ;
        RECT 84.050 113.110 84.220 113.450 ;
        RECT 84.390 113.280 84.720 113.710 ;
        RECT 84.955 113.110 85.125 113.450 ;
        RECT 80.890 112.650 82.110 112.820 ;
        RECT 82.280 112.740 82.740 113.030 ;
        RECT 83.045 112.910 83.605 113.080 ;
        RECT 84.050 112.940 85.125 113.110 ;
        RECT 85.295 113.210 85.975 113.540 ;
        RECT 86.190 113.210 86.440 113.540 ;
        RECT 86.610 113.250 86.860 113.710 ;
        RECT 83.435 112.770 83.605 112.910 ;
        RECT 82.280 112.730 83.245 112.740 ;
        RECT 81.940 112.560 82.110 112.650 ;
        RECT 82.570 112.570 83.245 112.730 ;
        RECT 80.550 112.360 80.895 112.370 ;
        RECT 78.865 112.150 80.895 112.360 ;
        RECT 77.290 111.710 78.040 111.880 ;
        RECT 78.270 111.810 80.035 111.980 ;
        RECT 77.285 111.160 77.615 111.540 ;
        RECT 77.785 111.420 78.040 111.710 ;
        RECT 78.525 111.160 78.695 111.630 ;
        RECT 78.865 111.330 79.195 111.810 ;
        RECT 79.365 111.160 79.535 111.630 ;
        RECT 79.705 111.330 80.035 111.810 ;
        RECT 80.205 111.160 80.375 111.970 ;
        RECT 80.570 111.895 80.895 112.150 ;
        RECT 80.575 111.540 80.895 111.895 ;
        RECT 81.065 112.110 81.605 112.480 ;
        RECT 81.940 112.390 82.345 112.560 ;
        RECT 81.065 111.710 81.305 112.110 ;
        RECT 81.785 111.940 82.005 112.220 ;
        RECT 81.475 111.770 82.005 111.940 ;
        RECT 81.475 111.540 81.645 111.770 ;
        RECT 82.175 111.610 82.345 112.390 ;
        RECT 82.515 111.780 82.865 112.400 ;
        RECT 83.035 111.780 83.245 112.570 ;
        RECT 83.435 112.600 84.935 112.770 ;
        RECT 83.435 111.910 83.605 112.600 ;
        RECT 85.295 112.430 85.465 113.210 ;
        RECT 86.270 113.080 86.440 113.210 ;
        RECT 83.775 112.260 85.465 112.430 ;
        RECT 85.635 112.650 86.100 113.040 ;
        RECT 86.270 112.910 86.665 113.080 ;
        RECT 83.775 112.080 83.945 112.260 ;
        RECT 80.575 111.370 81.645 111.540 ;
        RECT 81.815 111.160 82.005 111.600 ;
        RECT 82.175 111.330 83.125 111.610 ;
        RECT 83.435 111.520 83.695 111.910 ;
        RECT 84.115 111.840 84.905 112.090 ;
        RECT 83.345 111.350 83.695 111.520 ;
        RECT 83.905 111.160 84.235 111.620 ;
        RECT 85.110 111.550 85.280 112.260 ;
        RECT 85.635 112.060 85.805 112.650 ;
        RECT 85.450 111.840 85.805 112.060 ;
        RECT 85.975 111.840 86.325 112.460 ;
        RECT 86.495 111.550 86.665 112.910 ;
        RECT 87.030 112.740 87.355 113.525 ;
        RECT 86.835 111.690 87.295 112.740 ;
        RECT 85.110 111.380 85.965 111.550 ;
        RECT 86.170 111.380 86.665 111.550 ;
        RECT 86.835 111.160 87.165 111.520 ;
        RECT 87.525 111.420 87.695 113.540 ;
        RECT 87.865 113.210 88.195 113.710 ;
        RECT 88.365 113.040 88.620 113.540 ;
        RECT 87.870 112.870 88.620 113.040 ;
        RECT 87.870 111.880 88.100 112.870 ;
        RECT 88.270 112.050 88.620 112.700 ;
        RECT 88.855 112.570 89.065 113.710 ;
        RECT 89.235 112.560 89.565 113.540 ;
        RECT 89.735 112.570 89.965 113.710 ;
        RECT 90.235 112.570 90.445 113.710 ;
        RECT 90.615 112.560 90.945 113.540 ;
        RECT 91.115 112.570 91.345 113.710 ;
        RECT 87.870 111.710 88.620 111.880 ;
        RECT 87.865 111.160 88.195 111.540 ;
        RECT 88.365 111.420 88.620 111.710 ;
        RECT 88.855 111.160 89.065 111.980 ;
        RECT 89.235 111.960 89.485 112.560 ;
        RECT 89.655 112.150 89.985 112.400 ;
        RECT 89.235 111.330 89.565 111.960 ;
        RECT 89.735 111.160 89.965 111.980 ;
        RECT 90.235 111.160 90.445 111.980 ;
        RECT 90.615 111.960 90.865 112.560 ;
        RECT 92.475 112.545 92.765 113.710 ;
        RECT 93.245 112.870 93.415 113.710 ;
        RECT 93.625 112.700 93.875 113.540 ;
        RECT 94.085 112.870 94.255 113.710 ;
        RECT 94.425 112.700 94.715 113.540 ;
        RECT 92.990 112.530 94.715 112.700 ;
        RECT 94.925 112.650 95.095 113.710 ;
        RECT 95.390 113.330 95.720 113.710 ;
        RECT 95.900 113.160 96.070 113.450 ;
        RECT 96.240 113.250 96.490 113.710 ;
        RECT 95.270 112.990 96.070 113.160 ;
        RECT 96.660 113.200 97.530 113.540 ;
        RECT 91.035 112.150 91.365 112.400 ;
        RECT 92.990 111.980 93.400 112.530 ;
        RECT 95.270 112.370 95.440 112.990 ;
        RECT 96.660 112.820 96.830 113.200 ;
        RECT 97.765 113.080 97.935 113.540 ;
        RECT 98.105 113.250 98.475 113.710 ;
        RECT 98.770 113.110 98.940 113.450 ;
        RECT 99.110 113.280 99.440 113.710 ;
        RECT 99.675 113.110 99.845 113.450 ;
        RECT 95.610 112.650 96.830 112.820 ;
        RECT 97.000 112.740 97.460 113.030 ;
        RECT 97.765 112.910 98.325 113.080 ;
        RECT 98.770 112.940 99.845 113.110 ;
        RECT 100.015 113.210 100.695 113.540 ;
        RECT 100.910 113.210 101.160 113.540 ;
        RECT 101.330 113.250 101.580 113.710 ;
        RECT 98.155 112.770 98.325 112.910 ;
        RECT 97.000 112.730 97.965 112.740 ;
        RECT 96.660 112.560 96.830 112.650 ;
        RECT 97.290 112.570 97.965 112.730 ;
        RECT 95.270 112.360 95.615 112.370 ;
        RECT 93.585 112.150 95.615 112.360 ;
        RECT 90.615 111.330 90.945 111.960 ;
        RECT 91.115 111.160 91.345 111.980 ;
        RECT 92.475 111.160 92.765 111.885 ;
        RECT 92.990 111.810 94.755 111.980 ;
        RECT 93.245 111.160 93.415 111.630 ;
        RECT 93.585 111.330 93.915 111.810 ;
        RECT 94.085 111.160 94.255 111.630 ;
        RECT 94.425 111.330 94.755 111.810 ;
        RECT 94.925 111.160 95.095 111.970 ;
        RECT 95.290 111.895 95.615 112.150 ;
        RECT 95.295 111.540 95.615 111.895 ;
        RECT 95.785 112.110 96.325 112.480 ;
        RECT 96.660 112.390 97.065 112.560 ;
        RECT 95.785 111.710 96.025 112.110 ;
        RECT 96.505 111.940 96.725 112.220 ;
        RECT 96.195 111.770 96.725 111.940 ;
        RECT 96.195 111.540 96.365 111.770 ;
        RECT 96.895 111.610 97.065 112.390 ;
        RECT 97.235 111.780 97.585 112.400 ;
        RECT 97.755 111.780 97.965 112.570 ;
        RECT 98.155 112.600 99.655 112.770 ;
        RECT 98.155 111.910 98.325 112.600 ;
        RECT 100.015 112.430 100.185 113.210 ;
        RECT 100.990 113.080 101.160 113.210 ;
        RECT 98.495 112.260 100.185 112.430 ;
        RECT 100.355 112.650 100.820 113.040 ;
        RECT 100.990 112.910 101.385 113.080 ;
        RECT 98.495 112.080 98.665 112.260 ;
        RECT 95.295 111.370 96.365 111.540 ;
        RECT 96.535 111.160 96.725 111.600 ;
        RECT 96.895 111.330 97.845 111.610 ;
        RECT 98.155 111.520 98.415 111.910 ;
        RECT 98.835 111.840 99.625 112.090 ;
        RECT 98.065 111.350 98.415 111.520 ;
        RECT 98.625 111.160 98.955 111.620 ;
        RECT 99.830 111.550 100.000 112.260 ;
        RECT 100.355 112.060 100.525 112.650 ;
        RECT 100.170 111.840 100.525 112.060 ;
        RECT 100.695 111.840 101.045 112.460 ;
        RECT 101.215 111.550 101.385 112.910 ;
        RECT 101.750 112.740 102.075 113.525 ;
        RECT 101.555 111.690 102.015 112.740 ;
        RECT 99.830 111.380 100.685 111.550 ;
        RECT 100.890 111.380 101.385 111.550 ;
        RECT 101.555 111.160 101.885 111.520 ;
        RECT 102.245 111.420 102.415 113.540 ;
        RECT 102.585 113.210 102.915 113.710 ;
        RECT 103.085 113.040 103.340 113.540 ;
        RECT 102.590 112.870 103.340 113.040 ;
        RECT 103.825 112.870 103.995 113.710 ;
        RECT 102.590 111.880 102.820 112.870 ;
        RECT 104.205 112.700 104.455 113.540 ;
        RECT 104.665 112.870 104.835 113.710 ;
        RECT 105.005 112.700 105.295 113.540 ;
        RECT 102.990 112.050 103.340 112.700 ;
        RECT 103.570 112.530 105.295 112.700 ;
        RECT 105.505 112.650 105.675 113.710 ;
        RECT 105.970 113.330 106.300 113.710 ;
        RECT 106.480 113.160 106.650 113.450 ;
        RECT 106.820 113.250 107.070 113.710 ;
        RECT 105.850 112.990 106.650 113.160 ;
        RECT 107.240 113.200 108.110 113.540 ;
        RECT 103.570 111.980 103.980 112.530 ;
        RECT 105.850 112.370 106.020 112.990 ;
        RECT 107.240 112.820 107.410 113.200 ;
        RECT 108.345 113.080 108.515 113.540 ;
        RECT 108.685 113.250 109.055 113.710 ;
        RECT 109.350 113.110 109.520 113.450 ;
        RECT 109.690 113.280 110.020 113.710 ;
        RECT 110.255 113.110 110.425 113.450 ;
        RECT 106.190 112.650 107.410 112.820 ;
        RECT 107.580 112.740 108.040 113.030 ;
        RECT 108.345 112.910 108.905 113.080 ;
        RECT 109.350 112.940 110.425 113.110 ;
        RECT 110.595 113.210 111.275 113.540 ;
        RECT 111.490 113.210 111.740 113.540 ;
        RECT 111.910 113.250 112.160 113.710 ;
        RECT 108.735 112.770 108.905 112.910 ;
        RECT 107.580 112.730 108.545 112.740 ;
        RECT 107.240 112.560 107.410 112.650 ;
        RECT 107.870 112.570 108.545 112.730 ;
        RECT 105.850 112.360 106.195 112.370 ;
        RECT 104.165 112.150 106.195 112.360 ;
        RECT 102.590 111.710 103.340 111.880 ;
        RECT 103.570 111.810 105.335 111.980 ;
        RECT 102.585 111.160 102.915 111.540 ;
        RECT 103.085 111.420 103.340 111.710 ;
        RECT 103.825 111.160 103.995 111.630 ;
        RECT 104.165 111.330 104.495 111.810 ;
        RECT 104.665 111.160 104.835 111.630 ;
        RECT 105.005 111.330 105.335 111.810 ;
        RECT 105.505 111.160 105.675 111.970 ;
        RECT 105.870 111.895 106.195 112.150 ;
        RECT 105.875 111.540 106.195 111.895 ;
        RECT 106.365 112.110 106.905 112.480 ;
        RECT 107.240 112.390 107.645 112.560 ;
        RECT 106.365 111.710 106.605 112.110 ;
        RECT 107.085 111.940 107.305 112.220 ;
        RECT 106.775 111.770 107.305 111.940 ;
        RECT 106.775 111.540 106.945 111.770 ;
        RECT 107.475 111.610 107.645 112.390 ;
        RECT 107.815 111.780 108.165 112.400 ;
        RECT 108.335 111.780 108.545 112.570 ;
        RECT 108.735 112.600 110.235 112.770 ;
        RECT 108.735 111.910 108.905 112.600 ;
        RECT 110.595 112.430 110.765 113.210 ;
        RECT 111.570 113.080 111.740 113.210 ;
        RECT 109.075 112.260 110.765 112.430 ;
        RECT 110.935 112.650 111.400 113.040 ;
        RECT 111.570 112.910 111.965 113.080 ;
        RECT 109.075 112.080 109.245 112.260 ;
        RECT 105.875 111.370 106.945 111.540 ;
        RECT 107.115 111.160 107.305 111.600 ;
        RECT 107.475 111.330 108.425 111.610 ;
        RECT 108.735 111.520 108.995 111.910 ;
        RECT 109.415 111.840 110.205 112.090 ;
        RECT 108.645 111.350 108.995 111.520 ;
        RECT 109.205 111.160 109.535 111.620 ;
        RECT 110.410 111.550 110.580 112.260 ;
        RECT 110.935 112.060 111.105 112.650 ;
        RECT 110.750 111.840 111.105 112.060 ;
        RECT 111.275 111.840 111.625 112.460 ;
        RECT 111.795 111.550 111.965 112.910 ;
        RECT 112.330 112.740 112.655 113.525 ;
        RECT 112.135 111.690 112.595 112.740 ;
        RECT 110.410 111.380 111.265 111.550 ;
        RECT 111.470 111.380 111.965 111.550 ;
        RECT 112.135 111.160 112.465 111.520 ;
        RECT 112.825 111.420 112.995 113.540 ;
        RECT 113.165 113.210 113.495 113.710 ;
        RECT 113.665 113.040 113.920 113.540 ;
        RECT 113.170 112.870 113.920 113.040 ;
        RECT 113.170 111.880 113.400 112.870 ;
        RECT 114.185 112.780 114.355 113.540 ;
        RECT 114.535 112.950 114.865 113.710 ;
        RECT 113.570 112.050 113.920 112.700 ;
        RECT 114.185 112.610 114.850 112.780 ;
        RECT 115.035 112.635 115.305 113.540 ;
        RECT 114.680 112.465 114.850 112.610 ;
        RECT 114.115 112.060 114.445 112.430 ;
        RECT 114.680 112.135 114.965 112.465 ;
        RECT 114.680 111.880 114.850 112.135 ;
        RECT 113.170 111.710 113.920 111.880 ;
        RECT 113.165 111.160 113.495 111.540 ;
        RECT 113.665 111.420 113.920 111.710 ;
        RECT 114.185 111.710 114.850 111.880 ;
        RECT 115.135 111.835 115.305 112.635 ;
        RECT 115.475 112.620 117.145 113.710 ;
        RECT 117.315 112.620 118.525 113.710 ;
        RECT 115.475 112.100 116.225 112.620 ;
        RECT 116.395 111.930 117.145 112.450 ;
        RECT 117.315 112.080 117.835 112.620 ;
        RECT 114.185 111.330 114.355 111.710 ;
        RECT 114.535 111.160 114.865 111.540 ;
        RECT 115.045 111.330 115.305 111.835 ;
        RECT 115.475 111.160 117.145 111.930 ;
        RECT 118.005 111.910 118.525 112.450 ;
        RECT 117.315 111.160 118.525 111.910 ;
        RECT 11.430 110.990 118.610 111.160 ;
        RECT 11.515 110.240 12.725 110.990 ;
        RECT 11.515 109.700 12.035 110.240 ;
        RECT 13.355 110.220 15.025 110.990 ;
        RECT 15.195 110.265 15.485 110.990 ;
        RECT 15.965 110.520 16.135 110.990 ;
        RECT 16.305 110.340 16.635 110.820 ;
        RECT 16.805 110.520 16.975 110.990 ;
        RECT 17.145 110.340 17.475 110.820 ;
        RECT 12.205 109.530 12.725 110.070 ;
        RECT 11.515 108.440 12.725 109.530 ;
        RECT 13.355 109.530 14.105 110.050 ;
        RECT 14.275 109.700 15.025 110.220 ;
        RECT 15.710 110.170 17.475 110.340 ;
        RECT 17.645 110.180 17.815 110.990 ;
        RECT 18.015 110.610 19.085 110.780 ;
        RECT 18.015 110.255 18.335 110.610 ;
        RECT 15.710 109.620 16.120 110.170 ;
        RECT 18.010 110.000 18.335 110.255 ;
        RECT 16.305 109.790 18.335 110.000 ;
        RECT 17.990 109.780 18.335 109.790 ;
        RECT 18.505 110.040 18.745 110.440 ;
        RECT 18.915 110.380 19.085 110.610 ;
        RECT 19.255 110.550 19.445 110.990 ;
        RECT 19.615 110.540 20.565 110.820 ;
        RECT 20.785 110.630 21.135 110.800 ;
        RECT 18.915 110.210 19.445 110.380 ;
        RECT 13.355 108.440 15.025 109.530 ;
        RECT 15.195 108.440 15.485 109.605 ;
        RECT 15.710 109.450 17.435 109.620 ;
        RECT 15.965 108.440 16.135 109.280 ;
        RECT 16.345 108.610 16.595 109.450 ;
        RECT 16.805 108.440 16.975 109.280 ;
        RECT 17.145 108.610 17.435 109.450 ;
        RECT 17.645 108.440 17.815 109.500 ;
        RECT 17.990 109.160 18.160 109.780 ;
        RECT 18.505 109.670 19.045 110.040 ;
        RECT 19.225 109.930 19.445 110.210 ;
        RECT 19.615 109.760 19.785 110.540 ;
        RECT 19.380 109.590 19.785 109.760 ;
        RECT 19.955 109.750 20.305 110.370 ;
        RECT 19.380 109.500 19.550 109.590 ;
        RECT 20.475 109.580 20.685 110.370 ;
        RECT 18.330 109.330 19.550 109.500 ;
        RECT 20.010 109.420 20.685 109.580 ;
        RECT 17.990 108.990 18.790 109.160 ;
        RECT 18.110 108.440 18.440 108.820 ;
        RECT 18.620 108.700 18.790 108.990 ;
        RECT 19.380 108.950 19.550 109.330 ;
        RECT 19.720 109.410 20.685 109.420 ;
        RECT 20.875 110.240 21.135 110.630 ;
        RECT 21.345 110.530 21.675 110.990 ;
        RECT 22.550 110.600 23.405 110.770 ;
        RECT 23.610 110.600 24.105 110.770 ;
        RECT 24.275 110.630 24.605 110.990 ;
        RECT 20.875 109.550 21.045 110.240 ;
        RECT 21.215 109.890 21.385 110.070 ;
        RECT 21.555 110.060 22.345 110.310 ;
        RECT 22.550 109.890 22.720 110.600 ;
        RECT 22.890 110.090 23.245 110.310 ;
        RECT 21.215 109.720 22.905 109.890 ;
        RECT 19.720 109.120 20.180 109.410 ;
        RECT 20.875 109.380 22.375 109.550 ;
        RECT 20.875 109.240 21.045 109.380 ;
        RECT 20.485 109.070 21.045 109.240 ;
        RECT 18.960 108.440 19.210 108.900 ;
        RECT 19.380 108.610 20.250 108.950 ;
        RECT 20.485 108.610 20.655 109.070 ;
        RECT 21.490 109.040 22.565 109.210 ;
        RECT 20.825 108.440 21.195 108.900 ;
        RECT 21.490 108.700 21.660 109.040 ;
        RECT 21.830 108.440 22.160 108.870 ;
        RECT 22.395 108.700 22.565 109.040 ;
        RECT 22.735 108.940 22.905 109.720 ;
        RECT 23.075 109.500 23.245 110.090 ;
        RECT 23.415 109.690 23.765 110.310 ;
        RECT 23.075 109.110 23.540 109.500 ;
        RECT 23.935 109.240 24.105 110.600 ;
        RECT 24.275 109.410 24.735 110.460 ;
        RECT 23.710 109.070 24.105 109.240 ;
        RECT 23.710 108.940 23.880 109.070 ;
        RECT 22.735 108.610 23.415 108.940 ;
        RECT 23.630 108.610 23.880 108.940 ;
        RECT 24.050 108.440 24.300 108.900 ;
        RECT 24.470 108.625 24.795 109.410 ;
        RECT 24.965 108.610 25.135 110.730 ;
        RECT 25.305 110.610 25.635 110.990 ;
        RECT 25.805 110.440 26.060 110.730 ;
        RECT 25.310 110.270 26.060 110.440 ;
        RECT 25.310 109.280 25.540 110.270 ;
        RECT 26.295 110.170 26.505 110.990 ;
        RECT 26.675 110.190 27.005 110.820 ;
        RECT 25.710 109.450 26.060 110.100 ;
        RECT 26.675 109.590 26.925 110.190 ;
        RECT 27.175 110.170 27.405 110.990 ;
        RECT 28.075 110.265 28.365 110.990 ;
        RECT 28.535 110.240 29.745 110.990 ;
        RECT 29.920 110.445 35.265 110.990 ;
        RECT 35.440 110.445 40.785 110.990 ;
        RECT 27.095 109.750 27.425 110.000 ;
        RECT 25.310 109.110 26.060 109.280 ;
        RECT 25.305 108.440 25.635 108.940 ;
        RECT 25.805 108.610 26.060 109.110 ;
        RECT 26.295 108.440 26.505 109.580 ;
        RECT 26.675 108.610 27.005 109.590 ;
        RECT 27.175 108.440 27.405 109.580 ;
        RECT 28.075 108.440 28.365 109.605 ;
        RECT 28.535 109.530 29.055 110.070 ;
        RECT 29.225 109.700 29.745 110.240 ;
        RECT 28.535 108.440 29.745 109.530 ;
        RECT 31.510 108.875 31.860 110.125 ;
        RECT 33.340 109.615 33.680 110.445 ;
        RECT 37.030 108.875 37.380 110.125 ;
        RECT 38.860 109.615 39.200 110.445 ;
        RECT 40.955 110.265 41.245 110.990 ;
        RECT 41.880 110.445 47.225 110.990 ;
        RECT 29.920 108.440 35.265 108.875 ;
        RECT 35.440 108.440 40.785 108.875 ;
        RECT 40.955 108.440 41.245 109.605 ;
        RECT 43.470 108.875 43.820 110.125 ;
        RECT 45.300 109.615 45.640 110.445 ;
        RECT 47.455 110.170 47.665 110.990 ;
        RECT 47.835 110.190 48.165 110.820 ;
        RECT 47.835 109.590 48.085 110.190 ;
        RECT 48.335 110.170 48.565 110.990 ;
        RECT 48.775 110.220 51.365 110.990 ;
        RECT 48.255 109.750 48.585 110.000 ;
        RECT 41.880 108.440 47.225 108.875 ;
        RECT 47.455 108.440 47.665 109.580 ;
        RECT 47.835 108.610 48.165 109.590 ;
        RECT 48.335 108.440 48.565 109.580 ;
        RECT 48.775 109.530 49.985 110.050 ;
        RECT 50.155 109.700 51.365 110.220 ;
        RECT 51.595 110.170 51.805 110.990 ;
        RECT 51.975 110.190 52.305 110.820 ;
        RECT 51.975 109.590 52.225 110.190 ;
        RECT 52.475 110.170 52.705 110.990 ;
        RECT 53.835 110.265 54.125 110.990 ;
        RECT 54.755 110.220 58.265 110.990 ;
        RECT 52.395 109.750 52.725 110.000 ;
        RECT 48.775 108.440 51.365 109.530 ;
        RECT 51.595 108.440 51.805 109.580 ;
        RECT 51.975 108.610 52.305 109.590 ;
        RECT 52.475 108.440 52.705 109.580 ;
        RECT 53.835 108.440 54.125 109.605 ;
        RECT 54.755 109.530 56.445 110.050 ;
        RECT 56.615 109.700 58.265 110.220 ;
        RECT 58.495 110.170 58.705 110.990 ;
        RECT 58.875 110.190 59.205 110.820 ;
        RECT 58.875 109.590 59.125 110.190 ;
        RECT 59.375 110.170 59.605 110.990 ;
        RECT 59.815 110.240 61.025 110.990 ;
        RECT 61.200 110.445 66.545 110.990 ;
        RECT 59.295 109.750 59.625 110.000 ;
        RECT 54.755 108.440 58.265 109.530 ;
        RECT 58.495 108.440 58.705 109.580 ;
        RECT 58.875 108.610 59.205 109.590 ;
        RECT 59.375 108.440 59.605 109.580 ;
        RECT 59.815 109.530 60.335 110.070 ;
        RECT 60.505 109.700 61.025 110.240 ;
        RECT 59.815 108.440 61.025 109.530 ;
        RECT 62.790 108.875 63.140 110.125 ;
        RECT 64.620 109.615 64.960 110.445 ;
        RECT 66.715 110.265 67.005 110.990 ;
        RECT 67.180 110.445 72.525 110.990 ;
        RECT 72.700 110.445 78.045 110.990 ;
        RECT 61.200 108.440 66.545 108.875 ;
        RECT 66.715 108.440 67.005 109.605 ;
        RECT 68.770 108.875 69.120 110.125 ;
        RECT 70.600 109.615 70.940 110.445 ;
        RECT 74.290 108.875 74.640 110.125 ;
        RECT 76.120 109.615 76.460 110.445 ;
        RECT 78.255 110.170 78.485 110.990 ;
        RECT 78.655 110.190 78.985 110.820 ;
        RECT 78.235 109.750 78.565 110.000 ;
        RECT 78.735 109.590 78.985 110.190 ;
        RECT 79.155 110.170 79.365 110.990 ;
        RECT 79.595 110.265 79.885 110.990 ;
        RECT 80.055 110.220 81.725 110.990 ;
        RECT 82.205 110.520 82.375 110.990 ;
        RECT 82.545 110.340 82.875 110.820 ;
        RECT 83.045 110.520 83.215 110.990 ;
        RECT 83.385 110.340 83.715 110.820 ;
        RECT 67.180 108.440 72.525 108.875 ;
        RECT 72.700 108.440 78.045 108.875 ;
        RECT 78.255 108.440 78.485 109.580 ;
        RECT 78.655 108.610 78.985 109.590 ;
        RECT 79.155 108.440 79.365 109.580 ;
        RECT 79.595 108.440 79.885 109.605 ;
        RECT 80.055 109.530 80.805 110.050 ;
        RECT 80.975 109.700 81.725 110.220 ;
        RECT 81.950 110.170 83.715 110.340 ;
        RECT 83.885 110.180 84.055 110.990 ;
        RECT 84.255 110.610 85.325 110.780 ;
        RECT 84.255 110.255 84.575 110.610 ;
        RECT 81.950 109.620 82.360 110.170 ;
        RECT 84.250 110.000 84.575 110.255 ;
        RECT 82.545 109.790 84.575 110.000 ;
        RECT 84.230 109.780 84.575 109.790 ;
        RECT 84.745 110.040 84.985 110.440 ;
        RECT 85.155 110.380 85.325 110.610 ;
        RECT 85.495 110.550 85.685 110.990 ;
        RECT 85.855 110.540 86.805 110.820 ;
        RECT 87.025 110.630 87.375 110.800 ;
        RECT 85.155 110.210 85.685 110.380 ;
        RECT 80.055 108.440 81.725 109.530 ;
        RECT 81.950 109.450 83.675 109.620 ;
        RECT 82.205 108.440 82.375 109.280 ;
        RECT 82.585 108.610 82.835 109.450 ;
        RECT 83.045 108.440 83.215 109.280 ;
        RECT 83.385 108.610 83.675 109.450 ;
        RECT 83.885 108.440 84.055 109.500 ;
        RECT 84.230 109.160 84.400 109.780 ;
        RECT 84.745 109.670 85.285 110.040 ;
        RECT 85.465 109.930 85.685 110.210 ;
        RECT 85.855 109.760 86.025 110.540 ;
        RECT 85.620 109.590 86.025 109.760 ;
        RECT 86.195 109.750 86.545 110.370 ;
        RECT 85.620 109.500 85.790 109.590 ;
        RECT 86.715 109.580 86.925 110.370 ;
        RECT 84.570 109.330 85.790 109.500 ;
        RECT 86.250 109.420 86.925 109.580 ;
        RECT 84.230 108.990 85.030 109.160 ;
        RECT 84.350 108.440 84.680 108.820 ;
        RECT 84.860 108.700 85.030 108.990 ;
        RECT 85.620 108.950 85.790 109.330 ;
        RECT 85.960 109.410 86.925 109.420 ;
        RECT 87.115 110.240 87.375 110.630 ;
        RECT 87.585 110.530 87.915 110.990 ;
        RECT 88.790 110.600 89.645 110.770 ;
        RECT 89.850 110.600 90.345 110.770 ;
        RECT 90.515 110.630 90.845 110.990 ;
        RECT 87.115 109.550 87.285 110.240 ;
        RECT 87.455 109.890 87.625 110.070 ;
        RECT 87.795 110.060 88.585 110.310 ;
        RECT 88.790 109.890 88.960 110.600 ;
        RECT 89.130 110.090 89.485 110.310 ;
        RECT 87.455 109.720 89.145 109.890 ;
        RECT 85.960 109.120 86.420 109.410 ;
        RECT 87.115 109.380 88.615 109.550 ;
        RECT 87.115 109.240 87.285 109.380 ;
        RECT 86.725 109.070 87.285 109.240 ;
        RECT 85.200 108.440 85.450 108.900 ;
        RECT 85.620 108.610 86.490 108.950 ;
        RECT 86.725 108.610 86.895 109.070 ;
        RECT 87.730 109.040 88.805 109.210 ;
        RECT 87.065 108.440 87.435 108.900 ;
        RECT 87.730 108.700 87.900 109.040 ;
        RECT 88.070 108.440 88.400 108.870 ;
        RECT 88.635 108.700 88.805 109.040 ;
        RECT 88.975 108.940 89.145 109.720 ;
        RECT 89.315 109.500 89.485 110.090 ;
        RECT 89.655 109.690 90.005 110.310 ;
        RECT 89.315 109.110 89.780 109.500 ;
        RECT 90.175 109.240 90.345 110.600 ;
        RECT 90.515 109.410 90.975 110.460 ;
        RECT 89.950 109.070 90.345 109.240 ;
        RECT 89.950 108.940 90.120 109.070 ;
        RECT 88.975 108.610 89.655 108.940 ;
        RECT 89.870 108.610 90.120 108.940 ;
        RECT 90.290 108.440 90.540 108.900 ;
        RECT 90.710 108.625 91.035 109.410 ;
        RECT 91.205 108.610 91.375 110.730 ;
        RECT 91.545 110.610 91.875 110.990 ;
        RECT 92.045 110.440 92.300 110.730 ;
        RECT 91.550 110.270 92.300 110.440 ;
        RECT 91.550 109.280 91.780 110.270 ;
        RECT 92.475 110.265 92.765 110.990 ;
        RECT 92.935 110.240 94.145 110.990 ;
        RECT 94.320 110.445 99.665 110.990 ;
        RECT 99.840 110.445 105.185 110.990 ;
        RECT 91.950 109.450 92.300 110.100 ;
        RECT 91.550 109.110 92.300 109.280 ;
        RECT 91.545 108.440 91.875 108.940 ;
        RECT 92.045 108.610 92.300 109.110 ;
        RECT 92.475 108.440 92.765 109.605 ;
        RECT 92.935 109.530 93.455 110.070 ;
        RECT 93.625 109.700 94.145 110.240 ;
        RECT 92.935 108.440 94.145 109.530 ;
        RECT 95.910 108.875 96.260 110.125 ;
        RECT 97.740 109.615 98.080 110.445 ;
        RECT 101.430 108.875 101.780 110.125 ;
        RECT 103.260 109.615 103.600 110.445 ;
        RECT 105.355 110.265 105.645 110.990 ;
        RECT 106.735 110.220 110.245 110.990 ;
        RECT 94.320 108.440 99.665 108.875 ;
        RECT 99.840 108.440 105.185 108.875 ;
        RECT 105.355 108.440 105.645 109.605 ;
        RECT 106.735 109.530 108.425 110.050 ;
        RECT 108.595 109.700 110.245 110.220 ;
        RECT 110.455 110.170 110.685 110.990 ;
        RECT 110.855 110.190 111.185 110.820 ;
        RECT 110.435 109.750 110.765 110.000 ;
        RECT 110.935 109.590 111.185 110.190 ;
        RECT 111.355 110.170 111.565 110.990 ;
        RECT 111.800 110.445 117.145 110.990 ;
        RECT 106.735 108.440 110.245 109.530 ;
        RECT 110.455 108.440 110.685 109.580 ;
        RECT 110.855 108.610 111.185 109.590 ;
        RECT 111.355 108.440 111.565 109.580 ;
        RECT 113.390 108.875 113.740 110.125 ;
        RECT 115.220 109.615 115.560 110.445 ;
        RECT 117.315 110.240 118.525 110.990 ;
        RECT 117.315 109.530 117.835 110.070 ;
        RECT 118.005 109.700 118.525 110.240 ;
        RECT 111.800 108.440 117.145 108.875 ;
        RECT 117.315 108.440 118.525 109.530 ;
        RECT 11.430 108.270 118.610 108.440 ;
        RECT 19.165 66.070 30.165 66.940 ;
        RECT 19.165 54.930 20.835 66.070 ;
        RECT 21.465 65.555 26.465 65.725 ;
        RECT 21.235 55.300 21.405 65.340 ;
        RECT 26.525 55.300 26.695 65.340 ;
        RECT 27.095 54.930 27.265 66.070 ;
        RECT 27.895 65.555 28.895 65.725 ;
        RECT 27.665 55.300 27.835 65.340 ;
        RECT 28.955 55.300 29.125 65.340 ;
        RECT 29.525 54.930 30.165 66.070 ;
        RECT 19.165 52.860 30.165 54.930 ;
        RECT 19.165 49.370 21.005 52.860 ;
        RECT 22.765 52.780 30.165 52.860 ;
        RECT 21.635 52.350 22.135 52.520 ;
        RECT 21.405 50.095 21.575 52.135 ;
        RECT 22.195 50.095 22.365 52.135 ;
        RECT 21.635 49.710 22.135 49.880 ;
        RECT 22.765 49.370 25.085 52.780 ;
        RECT 25.715 52.270 26.215 52.440 ;
        RECT 19.165 48.650 25.085 49.370 ;
        RECT 19.135 48.040 23.045 48.260 ;
        RECT 19.135 45.640 20.855 48.040 ;
        RECT 21.485 47.530 21.985 47.700 ;
        RECT 21.255 46.320 21.425 47.360 ;
        RECT 22.045 46.320 22.215 47.360 ;
        RECT 21.485 45.980 21.985 46.150 ;
        RECT 22.615 45.640 23.045 48.040 ;
        RECT 24.025 46.290 25.085 48.650 ;
        RECT 25.485 47.015 25.655 52.055 ;
        RECT 26.275 47.015 26.445 52.055 ;
        RECT 25.715 46.630 26.215 46.800 ;
        RECT 26.845 46.290 27.015 52.780 ;
        RECT 27.645 52.270 28.145 52.440 ;
        RECT 27.415 47.015 27.585 52.055 ;
        RECT 28.205 47.015 28.375 52.055 ;
        RECT 27.645 46.630 28.145 46.800 ;
        RECT 28.775 46.290 30.165 52.780 ;
        RECT 30.365 66.080 41.365 66.950 ;
        RECT 30.365 54.940 32.035 66.080 ;
        RECT 32.665 65.565 37.665 65.735 ;
        RECT 32.435 55.310 32.605 65.350 ;
        RECT 37.725 55.310 37.895 65.350 ;
        RECT 38.295 54.940 38.465 66.080 ;
        RECT 39.095 65.565 40.095 65.735 ;
        RECT 38.865 55.310 39.035 65.350 ;
        RECT 40.155 55.310 40.325 65.350 ;
        RECT 40.725 54.940 41.365 66.080 ;
        RECT 30.365 52.870 41.365 54.940 ;
        RECT 30.365 49.380 32.205 52.870 ;
        RECT 33.965 52.790 41.365 52.870 ;
        RECT 32.835 52.360 33.335 52.530 ;
        RECT 32.605 50.105 32.775 52.145 ;
        RECT 33.395 50.105 33.565 52.145 ;
        RECT 32.835 49.720 33.335 49.890 ;
        RECT 33.965 49.380 36.285 52.790 ;
        RECT 36.915 52.280 37.415 52.450 ;
        RECT 30.365 48.660 36.285 49.380 ;
        RECT 24.025 45.800 30.165 46.290 ;
        RECT 30.335 48.050 34.245 48.270 ;
        RECT 19.135 45.370 23.045 45.640 ;
        RECT 30.335 45.650 32.055 48.050 ;
        RECT 32.685 47.540 33.185 47.710 ;
        RECT 32.455 46.330 32.625 47.370 ;
        RECT 33.245 46.330 33.415 47.370 ;
        RECT 32.685 45.990 33.185 46.160 ;
        RECT 33.815 45.650 34.245 48.050 ;
        RECT 35.225 46.300 36.285 48.660 ;
        RECT 36.685 47.025 36.855 52.065 ;
        RECT 37.475 47.025 37.645 52.065 ;
        RECT 36.915 46.640 37.415 46.810 ;
        RECT 38.045 46.300 38.215 52.790 ;
        RECT 38.845 52.280 39.345 52.450 ;
        RECT 38.615 47.025 38.785 52.065 ;
        RECT 39.405 47.025 39.575 52.065 ;
        RECT 38.845 46.640 39.345 46.810 ;
        RECT 39.975 46.300 41.365 52.790 ;
        RECT 41.585 66.050 52.585 66.920 ;
        RECT 41.585 54.910 43.255 66.050 ;
        RECT 43.885 65.535 48.885 65.705 ;
        RECT 43.655 55.280 43.825 65.320 ;
        RECT 48.945 55.280 49.115 65.320 ;
        RECT 49.515 54.910 49.685 66.050 ;
        RECT 50.315 65.535 51.315 65.705 ;
        RECT 50.085 55.280 50.255 65.320 ;
        RECT 51.375 55.280 51.545 65.320 ;
        RECT 51.945 54.910 52.585 66.050 ;
        RECT 41.585 52.840 52.585 54.910 ;
        RECT 41.585 49.350 43.425 52.840 ;
        RECT 45.185 52.760 52.585 52.840 ;
        RECT 44.055 52.330 44.555 52.500 ;
        RECT 43.825 50.075 43.995 52.115 ;
        RECT 44.615 50.075 44.785 52.115 ;
        RECT 44.055 49.690 44.555 49.860 ;
        RECT 45.185 49.350 47.505 52.760 ;
        RECT 48.135 52.250 48.635 52.420 ;
        RECT 41.585 48.630 47.505 49.350 ;
        RECT 35.225 45.810 41.365 46.300 ;
        RECT 41.555 48.020 45.465 48.240 ;
        RECT 30.335 45.380 34.245 45.650 ;
        RECT 41.555 45.620 43.275 48.020 ;
        RECT 43.905 47.510 44.405 47.680 ;
        RECT 43.675 46.300 43.845 47.340 ;
        RECT 44.465 46.300 44.635 47.340 ;
        RECT 43.905 45.960 44.405 46.130 ;
        RECT 45.035 45.620 45.465 48.020 ;
        RECT 46.445 46.270 47.505 48.630 ;
        RECT 47.905 46.995 48.075 52.035 ;
        RECT 48.695 46.995 48.865 52.035 ;
        RECT 48.135 46.610 48.635 46.780 ;
        RECT 49.265 46.270 49.435 52.760 ;
        RECT 50.065 52.250 50.565 52.420 ;
        RECT 49.835 46.995 50.005 52.035 ;
        RECT 50.625 46.995 50.795 52.035 ;
        RECT 50.065 46.610 50.565 46.780 ;
        RECT 51.195 46.270 52.585 52.760 ;
        RECT 52.835 66.030 63.835 66.900 ;
        RECT 52.835 54.890 54.505 66.030 ;
        RECT 55.135 65.515 60.135 65.685 ;
        RECT 54.905 55.260 55.075 65.300 ;
        RECT 60.195 55.260 60.365 65.300 ;
        RECT 60.765 54.890 60.935 66.030 ;
        RECT 61.565 65.515 62.565 65.685 ;
        RECT 61.335 55.260 61.505 65.300 ;
        RECT 62.625 55.260 62.795 65.300 ;
        RECT 63.195 54.890 63.835 66.030 ;
        RECT 52.835 52.820 63.835 54.890 ;
        RECT 52.835 49.330 54.675 52.820 ;
        RECT 56.435 52.740 63.835 52.820 ;
        RECT 55.305 52.310 55.805 52.480 ;
        RECT 55.075 50.055 55.245 52.095 ;
        RECT 55.865 50.055 56.035 52.095 ;
        RECT 55.305 49.670 55.805 49.840 ;
        RECT 56.435 49.330 58.755 52.740 ;
        RECT 59.385 52.230 59.885 52.400 ;
        RECT 52.835 48.610 58.755 49.330 ;
        RECT 46.445 45.780 52.585 46.270 ;
        RECT 52.805 48.000 56.715 48.220 ;
        RECT 41.555 45.350 45.465 45.620 ;
        RECT 52.805 45.600 54.525 48.000 ;
        RECT 55.155 47.490 55.655 47.660 ;
        RECT 54.925 46.280 55.095 47.320 ;
        RECT 55.715 46.280 55.885 47.320 ;
        RECT 55.155 45.940 55.655 46.110 ;
        RECT 56.285 45.600 56.715 48.000 ;
        RECT 57.695 46.250 58.755 48.610 ;
        RECT 59.155 46.975 59.325 52.015 ;
        RECT 59.945 46.975 60.115 52.015 ;
        RECT 59.385 46.590 59.885 46.760 ;
        RECT 60.515 46.250 60.685 52.740 ;
        RECT 61.315 52.230 61.815 52.400 ;
        RECT 61.085 46.975 61.255 52.015 ;
        RECT 61.875 46.975 62.045 52.015 ;
        RECT 61.315 46.590 61.815 46.760 ;
        RECT 62.445 46.250 63.835 52.740 ;
        RECT 64.055 66.020 75.055 66.890 ;
        RECT 64.055 54.880 65.725 66.020 ;
        RECT 66.355 65.505 71.355 65.675 ;
        RECT 66.125 55.250 66.295 65.290 ;
        RECT 71.415 55.250 71.585 65.290 ;
        RECT 71.985 54.880 72.155 66.020 ;
        RECT 72.785 65.505 73.785 65.675 ;
        RECT 72.555 55.250 72.725 65.290 ;
        RECT 73.845 55.250 74.015 65.290 ;
        RECT 74.415 54.880 75.055 66.020 ;
        RECT 64.055 52.810 75.055 54.880 ;
        RECT 64.055 49.320 65.895 52.810 ;
        RECT 67.655 52.730 75.055 52.810 ;
        RECT 66.525 52.300 67.025 52.470 ;
        RECT 66.295 50.045 66.465 52.085 ;
        RECT 67.085 50.045 67.255 52.085 ;
        RECT 66.525 49.660 67.025 49.830 ;
        RECT 67.655 49.320 69.975 52.730 ;
        RECT 70.605 52.220 71.105 52.390 ;
        RECT 64.055 48.600 69.975 49.320 ;
        RECT 57.695 45.760 63.835 46.250 ;
        RECT 64.025 47.990 67.935 48.210 ;
        RECT 52.805 45.330 56.715 45.600 ;
        RECT 64.025 45.590 65.745 47.990 ;
        RECT 66.375 47.480 66.875 47.650 ;
        RECT 66.145 46.270 66.315 47.310 ;
        RECT 66.935 46.270 67.105 47.310 ;
        RECT 66.375 45.930 66.875 46.100 ;
        RECT 67.505 45.590 67.935 47.990 ;
        RECT 68.915 46.240 69.975 48.600 ;
        RECT 70.375 46.965 70.545 52.005 ;
        RECT 71.165 46.965 71.335 52.005 ;
        RECT 70.605 46.580 71.105 46.750 ;
        RECT 71.735 46.240 71.905 52.730 ;
        RECT 72.535 52.220 73.035 52.390 ;
        RECT 72.305 46.965 72.475 52.005 ;
        RECT 73.095 46.965 73.265 52.005 ;
        RECT 72.535 46.580 73.035 46.750 ;
        RECT 73.665 46.240 75.055 52.730 ;
        RECT 75.295 66.010 86.295 66.880 ;
        RECT 75.295 54.870 76.965 66.010 ;
        RECT 77.595 65.495 82.595 65.665 ;
        RECT 77.365 55.240 77.535 65.280 ;
        RECT 82.655 55.240 82.825 65.280 ;
        RECT 83.225 54.870 83.395 66.010 ;
        RECT 84.025 65.495 85.025 65.665 ;
        RECT 83.795 55.240 83.965 65.280 ;
        RECT 85.085 55.240 85.255 65.280 ;
        RECT 85.655 54.870 86.295 66.010 ;
        RECT 75.295 52.800 86.295 54.870 ;
        RECT 75.295 49.310 77.135 52.800 ;
        RECT 78.895 52.720 86.295 52.800 ;
        RECT 77.765 52.290 78.265 52.460 ;
        RECT 77.535 50.035 77.705 52.075 ;
        RECT 78.325 50.035 78.495 52.075 ;
        RECT 77.765 49.650 78.265 49.820 ;
        RECT 78.895 49.310 81.215 52.720 ;
        RECT 81.845 52.210 82.345 52.380 ;
        RECT 75.295 48.590 81.215 49.310 ;
        RECT 68.915 45.750 75.055 46.240 ;
        RECT 75.265 47.980 79.175 48.200 ;
        RECT 64.025 45.320 67.935 45.590 ;
        RECT 75.265 45.580 76.985 47.980 ;
        RECT 77.615 47.470 78.115 47.640 ;
        RECT 77.385 46.260 77.555 47.300 ;
        RECT 78.175 46.260 78.345 47.300 ;
        RECT 77.615 45.920 78.115 46.090 ;
        RECT 78.745 45.580 79.175 47.980 ;
        RECT 80.155 46.230 81.215 48.590 ;
        RECT 81.615 46.955 81.785 51.995 ;
        RECT 82.405 46.955 82.575 51.995 ;
        RECT 81.845 46.570 82.345 46.740 ;
        RECT 82.975 46.230 83.145 52.720 ;
        RECT 83.775 52.210 84.275 52.380 ;
        RECT 83.545 46.955 83.715 51.995 ;
        RECT 84.335 46.955 84.505 51.995 ;
        RECT 83.775 46.570 84.275 46.740 ;
        RECT 84.905 46.230 86.295 52.720 ;
        RECT 86.545 66.020 97.545 66.890 ;
        RECT 131.125 66.880 140.025 66.890 ;
        RECT 86.545 54.880 88.215 66.020 ;
        RECT 88.845 65.505 93.845 65.675 ;
        RECT 88.615 55.250 88.785 65.290 ;
        RECT 93.905 55.250 94.075 65.290 ;
        RECT 94.475 54.880 94.645 66.020 ;
        RECT 95.275 65.505 96.275 65.675 ;
        RECT 95.045 55.250 95.215 65.290 ;
        RECT 96.335 55.250 96.505 65.290 ;
        RECT 96.905 54.880 97.545 66.020 ;
        RECT 86.545 52.810 97.545 54.880 ;
        RECT 86.545 49.320 88.385 52.810 ;
        RECT 90.145 52.730 97.545 52.810 ;
        RECT 89.015 52.300 89.515 52.470 ;
        RECT 88.785 50.045 88.955 52.085 ;
        RECT 89.575 50.045 89.745 52.085 ;
        RECT 89.015 49.660 89.515 49.830 ;
        RECT 90.145 49.320 92.465 52.730 ;
        RECT 93.095 52.220 93.595 52.390 ;
        RECT 86.545 48.600 92.465 49.320 ;
        RECT 80.155 45.740 86.295 46.230 ;
        RECT 86.515 47.990 90.425 48.210 ;
        RECT 75.265 45.310 79.175 45.580 ;
        RECT 86.515 45.590 88.235 47.990 ;
        RECT 88.865 47.480 89.365 47.650 ;
        RECT 88.635 46.270 88.805 47.310 ;
        RECT 89.425 46.270 89.595 47.310 ;
        RECT 88.865 45.930 89.365 46.100 ;
        RECT 89.995 45.590 90.425 47.990 ;
        RECT 91.405 46.240 92.465 48.600 ;
        RECT 92.865 46.965 93.035 52.005 ;
        RECT 93.655 46.965 93.825 52.005 ;
        RECT 93.095 46.580 93.595 46.750 ;
        RECT 94.225 46.240 94.395 52.730 ;
        RECT 95.025 52.220 95.525 52.390 ;
        RECT 94.795 46.965 94.965 52.005 ;
        RECT 95.585 46.965 95.755 52.005 ;
        RECT 95.025 46.580 95.525 46.750 ;
        RECT 96.155 46.240 97.545 52.730 ;
        RECT 97.825 66.010 108.825 66.880 ;
        RECT 97.825 54.870 99.495 66.010 ;
        RECT 100.125 65.495 105.125 65.665 ;
        RECT 99.895 55.240 100.065 65.280 ;
        RECT 105.185 55.240 105.355 65.280 ;
        RECT 105.755 54.870 105.925 66.010 ;
        RECT 106.555 65.495 107.555 65.665 ;
        RECT 106.325 55.240 106.495 65.280 ;
        RECT 107.615 55.240 107.785 65.280 ;
        RECT 108.185 54.870 108.825 66.010 ;
        RECT 97.825 52.800 108.825 54.870 ;
        RECT 97.825 49.310 99.665 52.800 ;
        RECT 101.425 52.720 108.825 52.800 ;
        RECT 100.295 52.290 100.795 52.460 ;
        RECT 100.065 50.035 100.235 52.075 ;
        RECT 100.855 50.035 101.025 52.075 ;
        RECT 100.295 49.650 100.795 49.820 ;
        RECT 101.425 49.310 103.745 52.720 ;
        RECT 104.375 52.210 104.875 52.380 ;
        RECT 97.825 48.590 103.745 49.310 ;
        RECT 91.405 45.750 97.545 46.240 ;
        RECT 97.795 47.980 101.705 48.200 ;
        RECT 86.515 45.320 90.425 45.590 ;
        RECT 97.795 45.580 99.515 47.980 ;
        RECT 100.145 47.470 100.645 47.640 ;
        RECT 99.915 46.260 100.085 47.300 ;
        RECT 100.705 46.260 100.875 47.300 ;
        RECT 100.145 45.920 100.645 46.090 ;
        RECT 101.275 45.580 101.705 47.980 ;
        RECT 102.685 46.230 103.745 48.590 ;
        RECT 104.145 46.955 104.315 51.995 ;
        RECT 104.935 46.955 105.105 51.995 ;
        RECT 104.375 46.570 104.875 46.740 ;
        RECT 105.505 46.230 105.675 52.720 ;
        RECT 106.305 52.210 106.805 52.380 ;
        RECT 106.075 46.955 106.245 51.995 ;
        RECT 106.865 46.955 107.035 51.995 ;
        RECT 106.305 46.570 106.805 46.740 ;
        RECT 107.435 46.230 108.825 52.720 ;
        RECT 109.095 66.010 120.095 66.880 ;
        RECT 109.095 54.870 110.765 66.010 ;
        RECT 111.395 65.495 116.395 65.665 ;
        RECT 111.165 55.240 111.335 65.280 ;
        RECT 116.455 55.240 116.625 65.280 ;
        RECT 117.025 54.870 117.195 66.010 ;
        RECT 117.825 65.495 118.825 65.665 ;
        RECT 117.595 55.240 117.765 65.280 ;
        RECT 118.885 55.240 119.055 65.280 ;
        RECT 119.455 54.870 120.095 66.010 ;
        RECT 109.095 52.800 120.095 54.870 ;
        RECT 109.095 49.310 110.935 52.800 ;
        RECT 112.695 52.720 120.095 52.800 ;
        RECT 111.565 52.290 112.065 52.460 ;
        RECT 111.335 50.035 111.505 52.075 ;
        RECT 112.125 50.035 112.295 52.075 ;
        RECT 111.565 49.650 112.065 49.820 ;
        RECT 112.695 49.310 115.015 52.720 ;
        RECT 115.645 52.210 116.145 52.380 ;
        RECT 109.095 48.590 115.015 49.310 ;
        RECT 102.685 45.740 108.825 46.230 ;
        RECT 109.065 47.980 112.975 48.200 ;
        RECT 97.795 45.310 101.705 45.580 ;
        RECT 109.065 45.580 110.785 47.980 ;
        RECT 111.415 47.470 111.915 47.640 ;
        RECT 111.185 46.260 111.355 47.300 ;
        RECT 111.975 46.260 112.145 47.300 ;
        RECT 111.415 45.920 111.915 46.090 ;
        RECT 112.545 45.580 112.975 47.980 ;
        RECT 113.955 46.230 115.015 48.590 ;
        RECT 115.415 46.955 115.585 51.995 ;
        RECT 116.205 46.955 116.375 51.995 ;
        RECT 115.645 46.570 116.145 46.740 ;
        RECT 116.775 46.230 116.945 52.720 ;
        RECT 117.575 52.210 118.075 52.380 ;
        RECT 117.345 46.955 117.515 51.995 ;
        RECT 118.135 46.955 118.305 51.995 ;
        RECT 117.575 46.570 118.075 46.740 ;
        RECT 118.705 46.230 120.095 52.720 ;
        RECT 120.345 66.010 140.025 66.880 ;
        RECT 120.345 54.870 122.015 66.010 ;
        RECT 122.645 65.495 127.645 65.665 ;
        RECT 122.415 55.240 122.585 65.280 ;
        RECT 127.705 55.240 127.875 65.280 ;
        RECT 128.275 54.870 128.445 66.010 ;
        RECT 130.705 65.980 140.025 66.010 ;
        RECT 129.075 65.495 130.075 65.665 ;
        RECT 128.845 55.240 129.015 65.280 ;
        RECT 130.135 55.240 130.305 65.280 ;
        RECT 130.705 54.870 132.765 65.980 ;
        RECT 133.395 65.465 138.395 65.635 ;
        RECT 133.165 55.210 133.335 65.250 ;
        RECT 138.455 55.210 138.625 65.250 ;
        RECT 120.345 54.840 132.765 54.870 ;
        RECT 139.025 54.840 140.025 65.980 ;
        RECT 120.345 54.720 140.025 54.840 ;
        RECT 120.345 53.550 140.035 54.720 ;
        RECT 120.345 52.800 131.345 53.550 ;
        RECT 120.345 49.310 122.185 52.800 ;
        RECT 123.945 52.720 131.345 52.800 ;
        RECT 122.815 52.290 123.315 52.460 ;
        RECT 122.585 50.035 122.755 52.075 ;
        RECT 123.375 50.035 123.545 52.075 ;
        RECT 122.815 49.650 123.315 49.820 ;
        RECT 123.945 49.310 126.265 52.720 ;
        RECT 126.895 52.210 127.395 52.380 ;
        RECT 120.345 48.590 126.265 49.310 ;
        RECT 113.955 45.740 120.095 46.230 ;
        RECT 120.315 47.980 124.225 48.200 ;
        RECT 109.065 45.310 112.975 45.580 ;
        RECT 120.315 45.580 122.035 47.980 ;
        RECT 122.665 47.470 123.165 47.640 ;
        RECT 122.435 46.260 122.605 47.300 ;
        RECT 123.225 46.260 123.395 47.300 ;
        RECT 122.665 45.920 123.165 46.090 ;
        RECT 123.795 45.580 124.225 47.980 ;
        RECT 125.205 46.230 126.265 48.590 ;
        RECT 126.665 46.955 126.835 51.995 ;
        RECT 127.455 46.955 127.625 51.995 ;
        RECT 126.895 46.570 127.395 46.740 ;
        RECT 128.025 46.230 128.195 52.720 ;
        RECT 128.825 52.210 129.325 52.380 ;
        RECT 128.595 46.955 128.765 51.995 ;
        RECT 129.385 46.955 129.555 51.995 ;
        RECT 128.825 46.570 129.325 46.740 ;
        RECT 129.955 46.230 131.345 52.720 ;
        RECT 125.205 45.740 131.345 46.230 ;
        RECT 120.315 45.310 124.225 45.580 ;
        RECT 25.695 39.770 29.605 40.040 ;
        RECT 18.575 39.120 24.715 39.610 ;
        RECT 18.575 32.630 19.965 39.120 ;
        RECT 20.595 38.610 21.095 38.780 ;
        RECT 20.365 33.355 20.535 38.395 ;
        RECT 21.155 33.355 21.325 38.395 ;
        RECT 20.595 32.970 21.095 33.140 ;
        RECT 21.725 32.630 21.895 39.120 ;
        RECT 22.525 38.610 23.025 38.780 ;
        RECT 22.295 33.355 22.465 38.395 ;
        RECT 23.085 33.355 23.255 38.395 ;
        RECT 23.655 36.760 24.715 39.120 ;
        RECT 25.695 37.370 26.125 39.770 ;
        RECT 26.755 39.260 27.255 39.430 ;
        RECT 26.525 38.050 26.695 39.090 ;
        RECT 27.315 38.050 27.485 39.090 ;
        RECT 26.755 37.710 27.255 37.880 ;
        RECT 27.885 37.370 29.605 39.770 ;
        RECT 36.975 39.770 40.885 40.040 ;
        RECT 25.695 37.150 29.605 37.370 ;
        RECT 29.855 39.120 35.995 39.610 ;
        RECT 23.655 36.040 29.575 36.760 ;
        RECT 22.525 32.970 23.025 33.140 ;
        RECT 23.655 32.630 25.975 36.040 ;
        RECT 26.605 35.530 27.105 35.700 ;
        RECT 26.375 33.275 26.545 35.315 ;
        RECT 27.165 33.275 27.335 35.315 ;
        RECT 26.605 32.890 27.105 33.060 ;
        RECT 18.575 32.550 25.975 32.630 ;
        RECT 27.735 32.550 29.575 36.040 ;
        RECT 18.575 30.480 29.575 32.550 ;
        RECT 18.575 19.340 19.215 30.480 ;
        RECT 19.615 20.070 19.785 30.110 ;
        RECT 20.905 20.070 21.075 30.110 ;
        RECT 19.845 19.685 20.845 19.855 ;
        RECT 21.475 19.340 21.645 30.480 ;
        RECT 22.045 20.070 22.215 30.110 ;
        RECT 27.335 20.070 27.505 30.110 ;
        RECT 22.275 19.685 27.275 19.855 ;
        RECT 27.905 19.340 29.575 30.480 ;
        RECT 18.575 18.470 29.575 19.340 ;
        RECT 29.855 32.630 31.245 39.120 ;
        RECT 31.875 38.610 32.375 38.780 ;
        RECT 31.645 33.355 31.815 38.395 ;
        RECT 32.435 33.355 32.605 38.395 ;
        RECT 31.875 32.970 32.375 33.140 ;
        RECT 33.005 32.630 33.175 39.120 ;
        RECT 33.805 38.610 34.305 38.780 ;
        RECT 33.575 33.355 33.745 38.395 ;
        RECT 34.365 33.355 34.535 38.395 ;
        RECT 34.935 36.760 35.995 39.120 ;
        RECT 36.975 37.370 37.405 39.770 ;
        RECT 38.035 39.260 38.535 39.430 ;
        RECT 37.805 38.050 37.975 39.090 ;
        RECT 38.595 38.050 38.765 39.090 ;
        RECT 38.035 37.710 38.535 37.880 ;
        RECT 39.165 37.370 40.885 39.770 ;
        RECT 48.265 39.750 52.175 40.020 ;
        RECT 36.975 37.150 40.885 37.370 ;
        RECT 41.145 39.100 47.285 39.590 ;
        RECT 34.935 36.040 40.855 36.760 ;
        RECT 33.805 32.970 34.305 33.140 ;
        RECT 34.935 32.630 37.255 36.040 ;
        RECT 37.885 35.530 38.385 35.700 ;
        RECT 37.655 33.275 37.825 35.315 ;
        RECT 38.445 33.275 38.615 35.315 ;
        RECT 37.885 32.890 38.385 33.060 ;
        RECT 29.855 32.550 37.255 32.630 ;
        RECT 39.015 32.550 40.855 36.040 ;
        RECT 29.855 30.480 40.855 32.550 ;
        RECT 29.855 19.340 30.495 30.480 ;
        RECT 30.895 20.070 31.065 30.110 ;
        RECT 32.185 20.070 32.355 30.110 ;
        RECT 31.125 19.685 32.125 19.855 ;
        RECT 32.755 19.340 32.925 30.480 ;
        RECT 33.325 20.070 33.495 30.110 ;
        RECT 38.615 20.070 38.785 30.110 ;
        RECT 33.555 19.685 38.555 19.855 ;
        RECT 39.185 19.340 40.855 30.480 ;
        RECT 29.855 18.470 40.855 19.340 ;
        RECT 41.145 32.610 42.535 39.100 ;
        RECT 43.165 38.590 43.665 38.760 ;
        RECT 42.935 33.335 43.105 38.375 ;
        RECT 43.725 33.335 43.895 38.375 ;
        RECT 43.165 32.950 43.665 33.120 ;
        RECT 44.295 32.610 44.465 39.100 ;
        RECT 45.095 38.590 45.595 38.760 ;
        RECT 44.865 33.335 45.035 38.375 ;
        RECT 45.655 33.335 45.825 38.375 ;
        RECT 46.225 36.740 47.285 39.100 ;
        RECT 48.265 37.350 48.695 39.750 ;
        RECT 49.325 39.240 49.825 39.410 ;
        RECT 49.095 38.030 49.265 39.070 ;
        RECT 49.885 38.030 50.055 39.070 ;
        RECT 49.325 37.690 49.825 37.860 ;
        RECT 50.455 37.350 52.175 39.750 ;
        RECT 59.485 39.750 63.395 40.020 ;
        RECT 48.265 37.130 52.175 37.350 ;
        RECT 52.365 39.100 58.505 39.590 ;
        RECT 46.225 36.020 52.145 36.740 ;
        RECT 45.095 32.950 45.595 33.120 ;
        RECT 46.225 32.610 48.545 36.020 ;
        RECT 49.175 35.510 49.675 35.680 ;
        RECT 48.945 33.255 49.115 35.295 ;
        RECT 49.735 33.255 49.905 35.295 ;
        RECT 49.175 32.870 49.675 33.040 ;
        RECT 41.145 32.530 48.545 32.610 ;
        RECT 50.305 32.530 52.145 36.020 ;
        RECT 41.145 30.460 52.145 32.530 ;
        RECT 41.145 19.320 41.785 30.460 ;
        RECT 42.185 20.050 42.355 30.090 ;
        RECT 43.475 20.050 43.645 30.090 ;
        RECT 42.415 19.665 43.415 19.835 ;
        RECT 44.045 19.320 44.215 30.460 ;
        RECT 44.615 20.050 44.785 30.090 ;
        RECT 49.905 20.050 50.075 30.090 ;
        RECT 44.845 19.665 49.845 19.835 ;
        RECT 50.475 19.320 52.145 30.460 ;
        RECT 41.145 18.450 52.145 19.320 ;
        RECT 52.365 32.610 53.755 39.100 ;
        RECT 54.385 38.590 54.885 38.760 ;
        RECT 54.155 33.335 54.325 38.375 ;
        RECT 54.945 33.335 55.115 38.375 ;
        RECT 54.385 32.950 54.885 33.120 ;
        RECT 55.515 32.610 55.685 39.100 ;
        RECT 56.315 38.590 56.815 38.760 ;
        RECT 56.085 33.335 56.255 38.375 ;
        RECT 56.875 33.335 57.045 38.375 ;
        RECT 57.445 36.740 58.505 39.100 ;
        RECT 59.485 37.350 59.915 39.750 ;
        RECT 60.545 39.240 61.045 39.410 ;
        RECT 60.315 38.030 60.485 39.070 ;
        RECT 61.105 38.030 61.275 39.070 ;
        RECT 60.545 37.690 61.045 37.860 ;
        RECT 61.675 37.350 63.395 39.750 ;
        RECT 70.685 39.750 74.595 40.020 ;
        RECT 59.485 37.130 63.395 37.350 ;
        RECT 63.565 39.100 69.705 39.590 ;
        RECT 57.445 36.020 63.365 36.740 ;
        RECT 56.315 32.950 56.815 33.120 ;
        RECT 57.445 32.610 59.765 36.020 ;
        RECT 60.395 35.510 60.895 35.680 ;
        RECT 60.165 33.255 60.335 35.295 ;
        RECT 60.955 33.255 61.125 35.295 ;
        RECT 60.395 32.870 60.895 33.040 ;
        RECT 52.365 32.530 59.765 32.610 ;
        RECT 61.525 32.530 63.365 36.020 ;
        RECT 52.365 30.460 63.365 32.530 ;
        RECT 52.365 19.320 53.005 30.460 ;
        RECT 53.405 20.050 53.575 30.090 ;
        RECT 54.695 20.050 54.865 30.090 ;
        RECT 53.635 19.665 54.635 19.835 ;
        RECT 55.265 19.320 55.435 30.460 ;
        RECT 55.835 20.050 56.005 30.090 ;
        RECT 61.125 20.050 61.295 30.090 ;
        RECT 56.065 19.665 61.065 19.835 ;
        RECT 61.695 19.320 63.365 30.460 ;
        RECT 52.365 18.450 63.365 19.320 ;
        RECT 63.565 32.610 64.955 39.100 ;
        RECT 65.585 38.590 66.085 38.760 ;
        RECT 65.355 33.335 65.525 38.375 ;
        RECT 66.145 33.335 66.315 38.375 ;
        RECT 65.585 32.950 66.085 33.120 ;
        RECT 66.715 32.610 66.885 39.100 ;
        RECT 67.515 38.590 68.015 38.760 ;
        RECT 67.285 33.335 67.455 38.375 ;
        RECT 68.075 33.335 68.245 38.375 ;
        RECT 68.645 36.740 69.705 39.100 ;
        RECT 70.685 37.350 71.115 39.750 ;
        RECT 71.745 39.240 72.245 39.410 ;
        RECT 71.515 38.030 71.685 39.070 ;
        RECT 72.305 38.030 72.475 39.070 ;
        RECT 71.745 37.690 72.245 37.860 ;
        RECT 72.875 37.350 74.595 39.750 ;
        RECT 81.975 39.740 85.885 40.010 ;
        RECT 70.685 37.130 74.595 37.350 ;
        RECT 74.855 39.090 80.995 39.580 ;
        RECT 68.645 36.020 74.565 36.740 ;
        RECT 67.515 32.950 68.015 33.120 ;
        RECT 68.645 32.610 70.965 36.020 ;
        RECT 71.595 35.510 72.095 35.680 ;
        RECT 71.365 33.255 71.535 35.295 ;
        RECT 72.155 33.255 72.325 35.295 ;
        RECT 71.595 32.870 72.095 33.040 ;
        RECT 63.565 32.530 70.965 32.610 ;
        RECT 72.725 32.530 74.565 36.020 ;
        RECT 63.565 30.460 74.565 32.530 ;
        RECT 63.565 19.320 64.205 30.460 ;
        RECT 64.605 20.050 64.775 30.090 ;
        RECT 65.895 20.050 66.065 30.090 ;
        RECT 64.835 19.665 65.835 19.835 ;
        RECT 66.465 19.320 66.635 30.460 ;
        RECT 67.035 20.050 67.205 30.090 ;
        RECT 72.325 20.050 72.495 30.090 ;
        RECT 67.265 19.665 72.265 19.835 ;
        RECT 72.895 19.320 74.565 30.460 ;
        RECT 63.565 18.450 74.565 19.320 ;
        RECT 74.855 32.600 76.245 39.090 ;
        RECT 76.875 38.580 77.375 38.750 ;
        RECT 76.645 33.325 76.815 38.365 ;
        RECT 77.435 33.325 77.605 38.365 ;
        RECT 76.875 32.940 77.375 33.110 ;
        RECT 78.005 32.600 78.175 39.090 ;
        RECT 78.805 38.580 79.305 38.750 ;
        RECT 78.575 33.325 78.745 38.365 ;
        RECT 79.365 33.325 79.535 38.365 ;
        RECT 79.935 36.730 80.995 39.090 ;
        RECT 81.975 37.340 82.405 39.740 ;
        RECT 83.035 39.230 83.535 39.400 ;
        RECT 82.805 38.020 82.975 39.060 ;
        RECT 83.595 38.020 83.765 39.060 ;
        RECT 83.035 37.680 83.535 37.850 ;
        RECT 84.165 37.340 85.885 39.740 ;
        RECT 93.215 39.760 97.125 40.030 ;
        RECT 81.975 37.120 85.885 37.340 ;
        RECT 86.095 39.110 92.235 39.600 ;
        RECT 79.935 36.010 85.855 36.730 ;
        RECT 78.805 32.940 79.305 33.110 ;
        RECT 79.935 32.600 82.255 36.010 ;
        RECT 82.885 35.500 83.385 35.670 ;
        RECT 82.655 33.245 82.825 35.285 ;
        RECT 83.445 33.245 83.615 35.285 ;
        RECT 82.885 32.860 83.385 33.030 ;
        RECT 74.855 32.520 82.255 32.600 ;
        RECT 84.015 32.520 85.855 36.010 ;
        RECT 74.855 30.450 85.855 32.520 ;
        RECT 74.855 19.310 75.495 30.450 ;
        RECT 75.895 20.040 76.065 30.080 ;
        RECT 77.185 20.040 77.355 30.080 ;
        RECT 76.125 19.655 77.125 19.825 ;
        RECT 77.755 19.310 77.925 30.450 ;
        RECT 78.325 20.040 78.495 30.080 ;
        RECT 83.615 20.040 83.785 30.080 ;
        RECT 78.555 19.655 83.555 19.825 ;
        RECT 84.185 19.310 85.855 30.450 ;
        RECT 74.855 18.440 85.855 19.310 ;
        RECT 86.095 32.620 87.485 39.110 ;
        RECT 88.115 38.600 88.615 38.770 ;
        RECT 87.885 33.345 88.055 38.385 ;
        RECT 88.675 33.345 88.845 38.385 ;
        RECT 88.115 32.960 88.615 33.130 ;
        RECT 89.245 32.620 89.415 39.110 ;
        RECT 90.045 38.600 90.545 38.770 ;
        RECT 89.815 33.345 89.985 38.385 ;
        RECT 90.605 33.345 90.775 38.385 ;
        RECT 91.175 36.750 92.235 39.110 ;
        RECT 93.215 37.360 93.645 39.760 ;
        RECT 94.275 39.250 94.775 39.420 ;
        RECT 94.045 38.040 94.215 39.080 ;
        RECT 94.835 38.040 95.005 39.080 ;
        RECT 94.275 37.700 94.775 37.870 ;
        RECT 95.405 37.360 97.125 39.760 ;
        RECT 104.425 39.780 108.335 40.050 ;
        RECT 93.215 37.140 97.125 37.360 ;
        RECT 97.305 39.130 103.445 39.620 ;
        RECT 91.175 36.030 97.095 36.750 ;
        RECT 90.045 32.960 90.545 33.130 ;
        RECT 91.175 32.620 93.495 36.030 ;
        RECT 94.125 35.520 94.625 35.690 ;
        RECT 93.895 33.265 94.065 35.305 ;
        RECT 94.685 33.265 94.855 35.305 ;
        RECT 94.125 32.880 94.625 33.050 ;
        RECT 86.095 32.540 93.495 32.620 ;
        RECT 95.255 32.540 97.095 36.030 ;
        RECT 86.095 30.470 97.095 32.540 ;
        RECT 86.095 19.330 86.735 30.470 ;
        RECT 87.135 20.060 87.305 30.100 ;
        RECT 88.425 20.060 88.595 30.100 ;
        RECT 87.365 19.675 88.365 19.845 ;
        RECT 88.995 19.330 89.165 30.470 ;
        RECT 89.565 20.060 89.735 30.100 ;
        RECT 94.855 20.060 95.025 30.100 ;
        RECT 89.795 19.675 94.795 19.845 ;
        RECT 95.425 19.330 97.095 30.470 ;
        RECT 86.095 18.460 97.095 19.330 ;
        RECT 97.305 32.640 98.695 39.130 ;
        RECT 99.325 38.620 99.825 38.790 ;
        RECT 99.095 33.365 99.265 38.405 ;
        RECT 99.885 33.365 100.055 38.405 ;
        RECT 99.325 32.980 99.825 33.150 ;
        RECT 100.455 32.640 100.625 39.130 ;
        RECT 101.255 38.620 101.755 38.790 ;
        RECT 101.025 33.365 101.195 38.405 ;
        RECT 101.815 33.365 101.985 38.405 ;
        RECT 102.385 36.770 103.445 39.130 ;
        RECT 104.425 37.380 104.855 39.780 ;
        RECT 105.485 39.270 105.985 39.440 ;
        RECT 105.255 38.060 105.425 39.100 ;
        RECT 106.045 38.060 106.215 39.100 ;
        RECT 105.485 37.720 105.985 37.890 ;
        RECT 106.615 37.380 108.335 39.780 ;
        RECT 115.625 39.820 119.535 40.090 ;
        RECT 104.425 37.160 108.335 37.380 ;
        RECT 108.505 39.170 114.645 39.660 ;
        RECT 102.385 36.050 108.305 36.770 ;
        RECT 101.255 32.980 101.755 33.150 ;
        RECT 102.385 32.640 104.705 36.050 ;
        RECT 105.335 35.540 105.835 35.710 ;
        RECT 105.105 33.285 105.275 35.325 ;
        RECT 105.895 33.285 106.065 35.325 ;
        RECT 105.335 32.900 105.835 33.070 ;
        RECT 97.305 32.560 104.705 32.640 ;
        RECT 106.465 32.560 108.305 36.050 ;
        RECT 97.305 30.490 108.305 32.560 ;
        RECT 97.305 19.350 97.945 30.490 ;
        RECT 98.345 20.080 98.515 30.120 ;
        RECT 99.635 20.080 99.805 30.120 ;
        RECT 98.575 19.695 99.575 19.865 ;
        RECT 100.205 19.350 100.375 30.490 ;
        RECT 100.775 20.080 100.945 30.120 ;
        RECT 106.065 20.080 106.235 30.120 ;
        RECT 101.005 19.695 106.005 19.865 ;
        RECT 106.635 19.350 108.305 30.490 ;
        RECT 97.305 18.480 108.305 19.350 ;
        RECT 108.505 32.680 109.895 39.170 ;
        RECT 110.525 38.660 111.025 38.830 ;
        RECT 110.295 33.405 110.465 38.445 ;
        RECT 111.085 33.405 111.255 38.445 ;
        RECT 110.525 33.020 111.025 33.190 ;
        RECT 111.655 32.680 111.825 39.170 ;
        RECT 112.455 38.660 112.955 38.830 ;
        RECT 112.225 33.405 112.395 38.445 ;
        RECT 113.015 33.405 113.185 38.445 ;
        RECT 113.585 36.810 114.645 39.170 ;
        RECT 115.625 37.420 116.055 39.820 ;
        RECT 116.685 39.310 117.185 39.480 ;
        RECT 116.455 38.100 116.625 39.140 ;
        RECT 117.245 38.100 117.415 39.140 ;
        RECT 116.685 37.760 117.185 37.930 ;
        RECT 117.815 37.420 119.535 39.820 ;
        RECT 126.835 39.840 130.745 40.110 ;
        RECT 115.625 37.200 119.535 37.420 ;
        RECT 119.715 39.190 125.855 39.680 ;
        RECT 113.585 36.090 119.505 36.810 ;
        RECT 112.455 33.020 112.955 33.190 ;
        RECT 113.585 32.680 115.905 36.090 ;
        RECT 116.535 35.580 117.035 35.750 ;
        RECT 116.305 33.325 116.475 35.365 ;
        RECT 117.095 33.325 117.265 35.365 ;
        RECT 116.535 32.940 117.035 33.110 ;
        RECT 108.505 32.600 115.905 32.680 ;
        RECT 117.665 32.600 119.505 36.090 ;
        RECT 108.505 30.530 119.505 32.600 ;
        RECT 108.505 19.390 109.145 30.530 ;
        RECT 109.545 20.120 109.715 30.160 ;
        RECT 110.835 20.120 111.005 30.160 ;
        RECT 109.775 19.735 110.775 19.905 ;
        RECT 111.405 19.390 111.575 30.530 ;
        RECT 111.975 20.120 112.145 30.160 ;
        RECT 117.265 20.120 117.435 30.160 ;
        RECT 112.205 19.735 117.205 19.905 ;
        RECT 117.835 19.390 119.505 30.530 ;
        RECT 108.505 18.520 119.505 19.390 ;
        RECT 119.715 32.700 121.105 39.190 ;
        RECT 121.735 38.680 122.235 38.850 ;
        RECT 121.505 33.425 121.675 38.465 ;
        RECT 122.295 33.425 122.465 38.465 ;
        RECT 121.735 33.040 122.235 33.210 ;
        RECT 122.865 32.700 123.035 39.190 ;
        RECT 123.665 38.680 124.165 38.850 ;
        RECT 123.435 33.425 123.605 38.465 ;
        RECT 124.225 33.425 124.395 38.465 ;
        RECT 124.795 36.830 125.855 39.190 ;
        RECT 126.835 37.440 127.265 39.840 ;
        RECT 127.895 39.330 128.395 39.500 ;
        RECT 127.665 38.120 127.835 39.160 ;
        RECT 128.455 38.120 128.625 39.160 ;
        RECT 127.895 37.780 128.395 37.950 ;
        RECT 129.025 37.440 130.745 39.840 ;
        RECT 126.835 37.220 130.745 37.440 ;
        RECT 124.795 36.110 130.715 36.830 ;
        RECT 123.665 33.040 124.165 33.210 ;
        RECT 124.795 32.700 127.115 36.110 ;
        RECT 127.745 35.600 128.245 35.770 ;
        RECT 127.515 33.345 127.685 35.385 ;
        RECT 128.305 33.345 128.475 35.385 ;
        RECT 127.745 32.960 128.245 33.130 ;
        RECT 119.715 32.620 127.115 32.700 ;
        RECT 128.875 32.620 130.715 36.110 ;
        RECT 119.715 31.140 130.715 32.620 ;
        RECT 119.715 30.550 139.465 31.140 ;
        RECT 119.715 19.410 120.355 30.550 ;
        RECT 120.755 20.140 120.925 30.180 ;
        RECT 122.045 20.140 122.215 30.180 ;
        RECT 120.985 19.755 121.985 19.925 ;
        RECT 122.615 19.410 122.785 30.550 ;
        RECT 129.045 30.520 139.465 30.550 ;
        RECT 123.185 20.140 123.355 30.180 ;
        RECT 128.475 20.140 128.645 30.180 ;
        RECT 123.415 19.755 128.415 19.925 ;
        RECT 129.045 19.410 132.075 30.520 ;
        RECT 132.475 20.110 132.645 30.150 ;
        RECT 137.765 20.110 137.935 30.150 ;
        RECT 132.705 19.725 137.705 19.895 ;
        RECT 119.715 19.380 132.075 19.410 ;
        RECT 138.335 19.380 139.465 30.520 ;
        RECT 119.715 18.540 139.465 19.380 ;
        RECT 131.925 18.520 139.465 18.540 ;
      LAYER met1 ;
        RECT 135.340 223.880 136.790 225.180 ;
        RECT 10.650 214.195 118.610 214.675 ;
        RECT 11.430 211.475 118.610 211.955 ;
        RECT 57.615 210.935 57.905 210.980 ;
        RECT 60.735 210.935 61.025 210.980 ;
        RECT 62.625 210.935 62.915 210.980 ;
        RECT 57.615 210.795 62.915 210.935 ;
        RECT 57.615 210.750 57.905 210.795 ;
        RECT 60.735 210.750 61.025 210.795 ;
        RECT 62.625 210.750 62.915 210.795 ;
        RECT 51.520 209.915 51.840 209.975 ;
        RECT 56.535 209.960 56.825 210.275 ;
        RECT 57.615 210.255 57.905 210.300 ;
        RECT 61.195 210.255 61.485 210.300 ;
        RECT 63.030 210.255 63.320 210.300 ;
        RECT 57.615 210.115 63.320 210.255 ;
        RECT 57.615 210.070 57.905 210.115 ;
        RECT 61.195 210.070 61.485 210.115 ;
        RECT 63.030 210.070 63.320 210.115 ;
        RECT 63.480 210.055 63.800 210.315 ;
        RECT 69.000 210.055 69.320 210.315 ;
        RECT 56.235 209.915 56.825 209.960 ;
        RECT 59.475 209.915 60.125 209.960 ;
        RECT 51.520 209.775 60.125 209.915 ;
        RECT 51.520 209.715 51.840 209.775 ;
        RECT 56.235 209.730 56.525 209.775 ;
        RECT 59.475 209.730 60.125 209.775 ;
        RECT 62.115 209.915 62.405 209.960 ;
        RECT 62.560 209.915 62.880 209.975 ;
        RECT 62.115 209.775 62.880 209.915 ;
        RECT 62.115 209.730 62.405 209.775 ;
        RECT 62.560 209.715 62.880 209.775 ;
        RECT 54.740 209.375 55.060 209.635 ;
        RECT 68.540 209.375 68.860 209.635 ;
        RECT 10.650 208.755 118.610 209.235 ;
        RECT 51.520 208.355 51.840 208.615 ;
        RECT 52.915 208.215 53.205 208.260 ;
        RECT 55.775 208.215 56.065 208.260 ;
        RECT 59.015 208.215 59.665 208.260 ;
        RECT 52.915 208.075 59.665 208.215 ;
        RECT 52.915 208.030 53.205 208.075 ;
        RECT 55.775 208.030 56.365 208.075 ;
        RECT 59.015 208.030 59.665 208.075 ;
        RECT 66.355 208.215 66.645 208.260 ;
        RECT 68.540 208.215 68.860 208.275 ;
        RECT 69.595 208.215 70.245 208.260 ;
        RECT 66.355 208.075 70.245 208.215 ;
        RECT 66.355 208.030 66.945 208.075 ;
        RECT 51.995 207.875 52.285 207.920 ;
        RECT 52.455 207.875 52.745 207.920 ;
        RECT 51.995 207.735 52.745 207.875 ;
        RECT 51.995 207.690 52.285 207.735 ;
        RECT 52.455 207.690 52.745 207.735 ;
        RECT 56.075 207.715 56.365 208.030 ;
        RECT 57.155 207.875 57.445 207.920 ;
        RECT 60.735 207.875 61.025 207.920 ;
        RECT 62.570 207.875 62.860 207.920 ;
        RECT 57.155 207.735 62.860 207.875 ;
        RECT 57.155 207.690 57.445 207.735 ;
        RECT 60.735 207.690 61.025 207.735 ;
        RECT 62.570 207.690 62.860 207.735 ;
        RECT 66.655 207.715 66.945 208.030 ;
        RECT 68.540 208.015 68.860 208.075 ;
        RECT 69.595 208.030 70.245 208.075 ;
        RECT 92.920 208.215 93.240 208.275 ;
        RECT 93.955 208.215 94.245 208.260 ;
        RECT 97.195 208.215 97.845 208.260 ;
        RECT 92.920 208.075 97.845 208.215 ;
        RECT 92.920 208.015 93.240 208.075 ;
        RECT 93.955 208.030 94.545 208.075 ;
        RECT 97.195 208.030 97.845 208.075 ;
        RECT 67.735 207.875 68.025 207.920 ;
        RECT 71.315 207.875 71.605 207.920 ;
        RECT 73.150 207.875 73.440 207.920 ;
        RECT 67.735 207.735 73.440 207.875 ;
        RECT 67.735 207.690 68.025 207.735 ;
        RECT 71.315 207.690 71.605 207.735 ;
        RECT 73.150 207.690 73.440 207.735 ;
        RECT 94.255 207.715 94.545 208.030 ;
        RECT 95.335 207.875 95.625 207.920 ;
        RECT 98.915 207.875 99.205 207.920 ;
        RECT 100.750 207.875 101.040 207.920 ;
        RECT 95.335 207.735 101.040 207.875 ;
        RECT 95.335 207.690 95.625 207.735 ;
        RECT 98.915 207.690 99.205 207.735 ;
        RECT 100.750 207.690 101.040 207.735 ;
        RECT 52.530 207.535 52.670 207.690 ;
        RECT 58.880 207.535 59.200 207.595 ;
        RECT 52.530 207.395 59.200 207.535 ;
        RECT 58.880 207.335 59.200 207.395 ;
        RECT 61.640 207.335 61.960 207.595 ;
        RECT 63.035 207.535 63.325 207.580 ;
        RECT 63.480 207.535 63.800 207.595 ;
        RECT 63.035 207.395 63.800 207.535 ;
        RECT 63.035 207.350 63.325 207.395 ;
        RECT 63.480 207.335 63.800 207.395 ;
        RECT 72.220 207.335 72.540 207.595 ;
        RECT 73.615 207.535 73.905 207.580 ;
        RECT 84.640 207.535 84.960 207.595 ;
        RECT 73.615 207.395 84.960 207.535 ;
        RECT 73.615 207.350 73.905 207.395 ;
        RECT 84.640 207.335 84.960 207.395 ;
        RECT 99.820 207.335 100.140 207.595 ;
        RECT 101.215 207.535 101.505 207.580 ;
        RECT 101.660 207.535 101.980 207.595 ;
        RECT 101.215 207.395 101.980 207.535 ;
        RECT 101.215 207.350 101.505 207.395 ;
        RECT 101.660 207.335 101.980 207.395 ;
        RECT 57.155 207.195 57.445 207.240 ;
        RECT 60.275 207.195 60.565 207.240 ;
        RECT 62.165 207.195 62.455 207.240 ;
        RECT 57.155 207.055 62.455 207.195 ;
        RECT 57.155 207.010 57.445 207.055 ;
        RECT 60.275 207.010 60.565 207.055 ;
        RECT 62.165 207.010 62.455 207.055 ;
        RECT 67.735 207.195 68.025 207.240 ;
        RECT 70.855 207.195 71.145 207.240 ;
        RECT 72.745 207.195 73.035 207.240 ;
        RECT 67.735 207.055 73.035 207.195 ;
        RECT 67.735 207.010 68.025 207.055 ;
        RECT 70.855 207.010 71.145 207.055 ;
        RECT 72.745 207.010 73.035 207.055 ;
        RECT 95.335 207.195 95.625 207.240 ;
        RECT 98.455 207.195 98.745 207.240 ;
        RECT 100.345 207.195 100.635 207.240 ;
        RECT 95.335 207.055 100.635 207.195 ;
        RECT 95.335 207.010 95.625 207.055 ;
        RECT 98.455 207.010 98.745 207.055 ;
        RECT 100.345 207.010 100.635 207.055 ;
        RECT 54.295 206.855 54.585 206.900 ;
        RECT 56.580 206.855 56.900 206.915 ;
        RECT 54.295 206.715 56.900 206.855 ;
        RECT 54.295 206.670 54.585 206.715 ;
        RECT 56.580 206.655 56.900 206.715 ;
        RECT 60.720 206.855 61.040 206.915 ;
        RECT 64.875 206.855 65.165 206.900 ;
        RECT 60.720 206.715 65.165 206.855 ;
        RECT 60.720 206.655 61.040 206.715 ;
        RECT 64.875 206.670 65.165 206.715 ;
        RECT 90.620 206.855 90.940 206.915 ;
        RECT 92.475 206.855 92.765 206.900 ;
        RECT 90.620 206.715 92.765 206.855 ;
        RECT 90.620 206.655 90.940 206.715 ;
        RECT 92.475 206.670 92.765 206.715 ;
        RECT 11.430 206.035 118.610 206.515 ;
        RECT 62.100 205.880 62.420 205.895 ;
        RECT 62.100 205.835 62.450 205.880 ;
        RECT 61.950 205.695 62.450 205.835 ;
        RECT 62.100 205.650 62.450 205.695 ;
        RECT 69.935 205.835 70.225 205.880 ;
        RECT 72.220 205.835 72.540 205.895 ;
        RECT 69.935 205.695 72.540 205.835 ;
        RECT 69.935 205.650 70.225 205.695 ;
        RECT 62.100 205.635 62.420 205.650 ;
        RECT 72.220 205.635 72.540 205.695 ;
        RECT 53.375 205.495 53.665 205.540 ;
        RECT 62.560 205.495 62.880 205.555 ;
        RECT 63.495 205.495 63.785 205.540 ;
        RECT 65.320 205.495 65.640 205.555 ;
        RECT 53.375 205.355 59.340 205.495 ;
        RECT 53.375 205.310 53.665 205.355 ;
        RECT 59.200 205.215 59.340 205.355 ;
        RECT 62.560 205.355 63.785 205.495 ;
        RECT 62.560 205.295 62.880 205.355 ;
        RECT 63.495 205.310 63.785 205.355 ;
        RECT 64.030 205.355 65.640 205.495 ;
        RECT 56.580 205.155 56.900 205.215 ;
        RECT 57.390 205.155 57.680 205.200 ;
        RECT 56.580 205.015 57.680 205.155 ;
        RECT 59.200 205.155 59.660 205.215 ;
        RECT 64.030 205.155 64.170 205.355 ;
        RECT 65.320 205.295 65.640 205.355 ;
        RECT 95.795 205.495 96.085 205.540 ;
        RECT 98.915 205.495 99.205 205.540 ;
        RECT 100.805 205.495 101.095 205.540 ;
        RECT 95.795 205.355 101.095 205.495 ;
        RECT 95.795 205.310 96.085 205.355 ;
        RECT 98.915 205.310 99.205 205.355 ;
        RECT 100.805 205.310 101.095 205.355 ;
        RECT 59.200 205.015 64.170 205.155 ;
        RECT 64.875 205.155 65.165 205.200 ;
        RECT 67.635 205.155 67.925 205.200 ;
        RECT 64.875 205.015 67.925 205.155 ;
        RECT 56.580 204.955 56.900 205.015 ;
        RECT 57.390 204.970 57.680 205.015 ;
        RECT 59.340 204.955 59.660 205.015 ;
        RECT 64.875 204.970 65.165 205.015 ;
        RECT 67.635 204.970 67.925 205.015 ;
        RECT 54.295 204.815 54.585 204.860 ;
        RECT 54.740 204.815 55.060 204.875 ;
        RECT 54.295 204.675 55.060 204.815 ;
        RECT 54.295 204.630 54.585 204.675 ;
        RECT 54.370 204.475 54.510 204.630 ;
        RECT 54.740 204.615 55.060 204.675 ;
        RECT 56.135 204.815 56.425 204.860 ;
        RECT 57.975 204.815 58.265 204.860 ;
        RECT 56.135 204.675 59.340 204.815 ;
        RECT 56.135 204.630 56.425 204.675 ;
        RECT 57.975 204.630 58.265 204.675 ;
        RECT 58.435 204.475 58.725 204.520 ;
        RECT 54.370 204.335 58.725 204.475 ;
        RECT 59.200 204.475 59.340 204.675 ;
        RECT 59.800 204.615 60.120 204.875 ;
        RECT 60.720 204.475 61.040 204.535 ;
        RECT 59.200 204.335 61.040 204.475 ;
        RECT 58.435 204.290 58.725 204.335 ;
        RECT 60.720 204.275 61.040 204.335 ;
        RECT 63.035 204.475 63.325 204.520 ;
        RECT 64.950 204.475 65.090 204.970 ;
        RECT 65.320 204.615 65.640 204.875 ;
        RECT 66.240 204.815 66.560 204.875 ;
        RECT 67.175 204.815 67.465 204.860 ;
        RECT 66.240 204.675 67.465 204.815 ;
        RECT 66.240 204.615 66.560 204.675 ;
        RECT 67.175 204.630 67.465 204.675 ;
        RECT 68.080 204.815 68.400 204.875 ;
        RECT 69.475 204.815 69.765 204.860 ;
        RECT 68.080 204.675 69.765 204.815 ;
        RECT 68.080 204.615 68.400 204.675 ;
        RECT 69.475 204.630 69.765 204.675 ;
        RECT 83.720 204.815 84.040 204.875 ;
        RECT 84.195 204.815 84.485 204.860 ;
        RECT 83.720 204.675 84.485 204.815 ;
        RECT 83.720 204.615 84.040 204.675 ;
        RECT 84.195 204.630 84.485 204.675 ;
        RECT 91.095 204.815 91.385 204.860 ;
        RECT 93.380 204.815 93.700 204.875 ;
        RECT 91.095 204.675 93.700 204.815 ;
        RECT 91.095 204.630 91.385 204.675 ;
        RECT 93.380 204.615 93.700 204.675 ;
        RECT 94.715 204.520 95.005 204.835 ;
        RECT 95.795 204.815 96.085 204.860 ;
        RECT 99.375 204.815 99.665 204.860 ;
        RECT 101.210 204.815 101.500 204.860 ;
        RECT 95.795 204.675 101.500 204.815 ;
        RECT 95.795 204.630 96.085 204.675 ;
        RECT 99.375 204.630 99.665 204.675 ;
        RECT 101.210 204.630 101.500 204.675 ;
        RECT 101.660 204.815 101.980 204.875 ;
        RECT 103.960 204.815 104.280 204.875 ;
        RECT 101.660 204.675 104.280 204.815 ;
        RECT 101.660 204.615 101.980 204.675 ;
        RECT 103.960 204.615 104.280 204.675 ;
        RECT 63.035 204.335 65.090 204.475 ;
        RECT 91.555 204.475 91.845 204.520 ;
        RECT 94.415 204.475 95.005 204.520 ;
        RECT 97.655 204.475 98.305 204.520 ;
        RECT 91.555 204.335 98.305 204.475 ;
        RECT 63.035 204.290 63.325 204.335 ;
        RECT 91.555 204.290 91.845 204.335 ;
        RECT 94.415 204.290 94.705 204.335 ;
        RECT 97.655 204.290 98.305 204.335 ;
        RECT 98.900 204.475 99.220 204.535 ;
        RECT 100.295 204.475 100.585 204.520 ;
        RECT 98.900 204.335 100.585 204.475 ;
        RECT 98.900 204.275 99.220 204.335 ;
        RECT 100.295 204.290 100.585 204.335 ;
        RECT 55.200 203.935 55.520 204.195 ;
        RECT 56.595 204.135 56.885 204.180 ;
        RECT 57.960 204.135 58.280 204.195 ;
        RECT 56.595 203.995 58.280 204.135 ;
        RECT 56.595 203.950 56.885 203.995 ;
        RECT 57.960 203.935 58.280 203.995 ;
        RECT 61.180 203.935 61.500 204.195 ;
        RECT 62.035 204.135 62.325 204.180 ;
        RECT 62.560 204.135 62.880 204.195 ;
        RECT 62.035 203.995 62.880 204.135 ;
        RECT 62.035 203.950 62.325 203.995 ;
        RECT 62.560 203.935 62.880 203.995 ;
        RECT 85.115 204.135 85.405 204.180 ;
        RECT 86.020 204.135 86.340 204.195 ;
        RECT 85.115 203.995 86.340 204.135 ;
        RECT 85.115 203.950 85.405 203.995 ;
        RECT 86.020 203.935 86.340 203.995 ;
        RECT 92.935 204.135 93.225 204.180 ;
        RECT 93.840 204.135 94.160 204.195 ;
        RECT 92.935 203.995 94.160 204.135 ;
        RECT 92.935 203.950 93.225 203.995 ;
        RECT 93.840 203.935 94.160 203.995 ;
        RECT 10.650 203.315 118.610 203.795 ;
        RECT 55.200 203.115 55.520 203.175 ;
        RECT 55.200 202.975 60.490 203.115 ;
        RECT 55.200 202.915 55.520 202.975 ;
        RECT 56.135 202.775 56.425 202.820 ;
        RECT 56.580 202.775 56.900 202.835 ;
        RECT 56.135 202.635 56.900 202.775 ;
        RECT 56.135 202.590 56.425 202.635 ;
        RECT 56.580 202.575 56.900 202.635 ;
        RECT 57.975 202.775 58.265 202.820 ;
        RECT 59.800 202.775 60.120 202.835 ;
        RECT 57.975 202.635 60.120 202.775 ;
        RECT 60.350 202.775 60.490 202.975 ;
        RECT 60.720 202.915 61.040 203.175 ;
        RECT 62.100 203.115 62.420 203.175 ;
        RECT 62.575 203.115 62.865 203.160 ;
        RECT 62.100 202.975 62.865 203.115 ;
        RECT 62.100 202.915 62.420 202.975 ;
        RECT 62.575 202.930 62.865 202.975 ;
        RECT 63.020 203.115 63.340 203.175 ;
        RECT 65.335 203.115 65.625 203.160 ;
        RECT 63.020 202.975 65.625 203.115 ;
        RECT 63.020 202.915 63.340 202.975 ;
        RECT 65.335 202.930 65.625 202.975 ;
        RECT 80.055 203.115 80.345 203.160 ;
        RECT 80.055 202.975 88.090 203.115 ;
        RECT 80.055 202.930 80.345 202.975 ;
        RECT 61.640 202.775 61.960 202.835 ;
        RECT 67.175 202.775 67.465 202.820 ;
        RECT 68.080 202.775 68.400 202.835 ;
        RECT 60.350 202.635 68.400 202.775 ;
        RECT 57.975 202.590 58.265 202.635 ;
        RECT 59.800 202.575 60.120 202.635 ;
        RECT 61.640 202.575 61.960 202.635 ;
        RECT 67.175 202.590 67.465 202.635 ;
        RECT 68.080 202.575 68.400 202.635 ;
        RECT 78.675 202.775 78.965 202.820 ;
        RECT 81.535 202.775 81.825 202.820 ;
        RECT 84.775 202.775 85.425 202.820 ;
        RECT 78.675 202.635 85.425 202.775 ;
        RECT 78.675 202.590 78.965 202.635 ;
        RECT 81.535 202.590 82.125 202.635 ;
        RECT 84.775 202.590 85.425 202.635 ;
        RECT 86.020 202.775 86.340 202.835 ;
        RECT 87.415 202.775 87.705 202.820 ;
        RECT 86.020 202.635 87.705 202.775 ;
        RECT 87.950 202.775 88.090 202.975 ;
        RECT 92.920 202.915 93.240 203.175 ;
        RECT 98.900 202.915 99.220 203.175 ;
        RECT 99.820 203.115 100.140 203.175 ;
        RECT 100.295 203.115 100.585 203.160 ;
        RECT 99.820 202.975 100.585 203.115 ;
        RECT 99.820 202.915 100.140 202.975 ;
        RECT 100.295 202.930 100.585 202.975 ;
        RECT 95.695 202.775 95.985 202.820 ;
        RECT 87.950 202.635 95.985 202.775 ;
        RECT 56.670 202.435 56.810 202.575 ;
        RECT 60.275 202.435 60.565 202.480 ;
        RECT 56.670 202.295 60.565 202.435 ;
        RECT 60.275 202.250 60.565 202.295 ;
        RECT 61.180 202.435 61.500 202.495 ;
        RECT 63.495 202.435 63.785 202.480 ;
        RECT 61.180 202.295 63.785 202.435 ;
        RECT 61.180 202.235 61.500 202.295 ;
        RECT 63.495 202.250 63.785 202.295 ;
        RECT 66.240 202.235 66.560 202.495 ;
        RECT 69.000 202.435 69.320 202.495 ;
        RECT 78.215 202.435 78.505 202.480 ;
        RECT 69.000 202.295 78.505 202.435 ;
        RECT 69.000 202.235 69.320 202.295 ;
        RECT 78.215 202.250 78.505 202.295 ;
        RECT 81.835 202.275 82.125 202.590 ;
        RECT 86.020 202.575 86.340 202.635 ;
        RECT 87.415 202.590 87.705 202.635 ;
        RECT 93.010 202.495 93.150 202.635 ;
        RECT 95.695 202.590 95.985 202.635 ;
        RECT 82.915 202.435 83.205 202.480 ;
        RECT 86.495 202.435 86.785 202.480 ;
        RECT 88.330 202.435 88.620 202.480 ;
        RECT 92.475 202.435 92.765 202.480 ;
        RECT 82.915 202.295 88.620 202.435 ;
        RECT 82.915 202.250 83.205 202.295 ;
        RECT 86.495 202.250 86.785 202.295 ;
        RECT 88.330 202.250 88.620 202.295 ;
        RECT 89.330 202.295 92.765 202.435 ;
        RECT 66.330 202.095 66.470 202.235 ;
        RECT 60.810 201.955 66.470 202.095 ;
        RECT 57.975 201.755 58.265 201.800 ;
        RECT 59.340 201.755 59.660 201.815 ;
        RECT 57.975 201.615 59.660 201.755 ;
        RECT 57.975 201.570 58.265 201.615 ;
        RECT 59.340 201.555 59.660 201.615 ;
        RECT 60.810 201.475 60.950 201.955 ;
        RECT 56.595 201.415 56.885 201.460 ;
        RECT 60.720 201.415 61.040 201.475 ;
        RECT 56.595 201.275 61.040 201.415 ;
        RECT 56.595 201.230 56.885 201.275 ;
        RECT 60.720 201.215 61.040 201.275 ;
        RECT 61.655 201.415 61.945 201.460 ;
        RECT 62.100 201.415 62.420 201.475 ;
        RECT 61.655 201.275 62.420 201.415 ;
        RECT 78.290 201.415 78.430 202.250 ;
        RECT 85.560 202.095 85.880 202.155 ;
        RECT 88.795 202.095 89.085 202.140 ;
        RECT 85.560 201.955 89.085 202.095 ;
        RECT 85.560 201.895 85.880 201.955 ;
        RECT 88.795 201.910 89.085 201.955 ;
        RECT 82.915 201.755 83.205 201.800 ;
        RECT 86.035 201.755 86.325 201.800 ;
        RECT 87.925 201.755 88.215 201.800 ;
        RECT 82.915 201.615 88.215 201.755 ;
        RECT 82.915 201.570 83.205 201.615 ;
        RECT 86.035 201.570 86.325 201.615 ;
        RECT 87.925 201.570 88.215 201.615 ;
        RECT 89.330 201.415 89.470 202.295 ;
        RECT 92.475 202.250 92.765 202.295 ;
        RECT 92.550 202.095 92.690 202.250 ;
        RECT 92.920 202.235 93.240 202.495 ;
        RECT 93.840 202.435 94.160 202.495 ;
        RECT 97.995 202.435 98.285 202.480 ;
        RECT 93.840 202.295 95.450 202.435 ;
        RECT 93.840 202.235 94.160 202.295 ;
        RECT 93.380 202.095 93.700 202.155 ;
        RECT 92.550 201.955 93.700 202.095 ;
        RECT 93.380 201.895 93.700 201.955 ;
        RECT 94.760 201.895 95.080 202.155 ;
        RECT 95.310 202.140 95.450 202.295 ;
        RECT 97.610 202.295 98.285 202.435 ;
        RECT 95.235 202.095 95.525 202.140 ;
        RECT 96.600 202.095 96.920 202.155 ;
        RECT 95.235 201.955 96.920 202.095 ;
        RECT 95.235 201.910 95.525 201.955 ;
        RECT 96.600 201.895 96.920 201.955 ;
        RECT 97.610 201.800 97.750 202.295 ;
        RECT 97.995 202.250 98.285 202.295 ;
        RECT 99.360 202.235 99.680 202.495 ;
        RECT 97.535 201.570 97.825 201.800 ;
        RECT 78.290 201.275 89.470 201.415 ;
        RECT 61.655 201.230 61.945 201.275 ;
        RECT 62.100 201.215 62.420 201.275 ;
        RECT 11.430 200.595 118.610 201.075 ;
        RECT 69.000 200.395 69.320 200.455 ;
        RECT 59.200 200.255 69.320 200.395 ;
        RECT 59.200 200.115 59.340 200.255 ;
        RECT 69.000 200.195 69.320 200.255 ;
        RECT 98.455 200.395 98.745 200.440 ;
        RECT 99.360 200.395 99.680 200.455 ;
        RECT 98.455 200.255 99.680 200.395 ;
        RECT 98.455 200.210 98.745 200.255 ;
        RECT 99.360 200.195 99.680 200.255 ;
        RECT 53.325 200.055 53.615 200.100 ;
        RECT 55.215 200.055 55.505 200.100 ;
        RECT 58.335 200.055 58.625 200.100 ;
        RECT 53.325 199.915 58.625 200.055 ;
        RECT 53.325 199.870 53.615 199.915 ;
        RECT 55.215 199.870 55.505 199.915 ;
        RECT 58.335 199.870 58.625 199.915 ;
        RECT 58.880 199.915 59.340 200.115 ;
        RECT 63.480 200.055 63.800 200.115 ;
        RECT 62.190 199.915 63.800 200.055 ;
        RECT 58.880 199.855 59.200 199.915 ;
        RECT 62.190 199.715 62.330 199.915 ;
        RECT 63.480 199.855 63.800 199.915 ;
        RECT 79.550 200.055 79.840 200.100 ;
        RECT 82.330 200.055 82.620 200.100 ;
        RECT 84.190 200.055 84.480 200.100 ;
        RECT 79.550 199.915 84.480 200.055 ;
        RECT 79.550 199.870 79.840 199.915 ;
        RECT 82.330 199.870 82.620 199.915 ;
        RECT 84.190 199.870 84.480 199.915 ;
        RECT 43.330 199.575 47.610 199.715 ;
        RECT 43.330 199.420 43.470 199.575 ;
        RECT 43.255 199.190 43.545 199.420 ;
        RECT 46.000 199.175 46.320 199.435 ;
        RECT 47.470 199.420 47.610 199.575 ;
        RECT 52.530 199.575 62.330 199.715 ;
        RECT 52.530 199.435 52.670 199.575 ;
        RECT 95.220 199.515 95.540 199.775 ;
        RECT 47.395 199.375 47.685 199.420 ;
        RECT 47.840 199.375 48.160 199.435 ;
        RECT 47.395 199.235 48.160 199.375 ;
        RECT 47.395 199.190 47.685 199.235 ;
        RECT 47.840 199.175 48.160 199.235 ;
        RECT 52.440 199.175 52.760 199.435 ;
        RECT 52.920 199.375 53.210 199.420 ;
        RECT 54.755 199.375 55.045 199.420 ;
        RECT 58.335 199.375 58.625 199.420 ;
        RECT 52.920 199.235 58.625 199.375 ;
        RECT 52.920 199.190 53.210 199.235 ;
        RECT 54.755 199.190 55.045 199.235 ;
        RECT 58.335 199.190 58.625 199.235 ;
        RECT 53.835 198.850 54.125 199.080 ;
        RECT 56.115 199.035 56.765 199.080 ;
        RECT 57.500 199.035 57.820 199.095 ;
        RECT 59.415 199.080 59.705 199.395 ;
        RECT 60.260 199.375 60.580 199.435 ;
        RECT 62.575 199.375 62.865 199.420 ;
        RECT 63.480 199.375 63.800 199.435 ;
        RECT 60.260 199.235 63.800 199.375 ;
        RECT 60.260 199.175 60.580 199.235 ;
        RECT 62.575 199.190 62.865 199.235 ;
        RECT 63.480 199.175 63.800 199.235 ;
        RECT 79.550 199.375 79.840 199.420 ;
        RECT 82.815 199.375 83.105 199.420 ;
        RECT 84.180 199.375 84.500 199.435 ;
        RECT 79.550 199.235 82.085 199.375 ;
        RECT 79.550 199.190 79.840 199.235 ;
        RECT 59.415 199.035 60.005 199.080 ;
        RECT 56.115 198.895 60.005 199.035 ;
        RECT 56.115 198.850 56.765 198.895 ;
        RECT 40.020 198.695 40.340 198.755 ;
        RECT 42.795 198.695 43.085 198.740 ;
        RECT 40.020 198.555 43.085 198.695 ;
        RECT 40.020 198.495 40.340 198.555 ;
        RECT 42.795 198.510 43.085 198.555 ;
        RECT 44.160 198.695 44.480 198.755 ;
        RECT 45.095 198.695 45.385 198.740 ;
        RECT 44.160 198.555 45.385 198.695 ;
        RECT 44.160 198.495 44.480 198.555 ;
        RECT 45.095 198.510 45.385 198.555 ;
        RECT 46.935 198.695 47.225 198.740 ;
        RECT 47.380 198.695 47.700 198.755 ;
        RECT 46.935 198.555 47.700 198.695 ;
        RECT 53.910 198.695 54.050 198.850 ;
        RECT 57.500 198.835 57.820 198.895 ;
        RECT 59.715 198.850 60.005 198.895 ;
        RECT 77.690 199.035 77.980 199.080 ;
        RECT 79.120 199.035 79.440 199.095 ;
        RECT 81.870 199.080 82.085 199.235 ;
        RECT 82.815 199.235 84.500 199.375 ;
        RECT 82.815 199.190 83.105 199.235 ;
        RECT 84.180 199.175 84.500 199.235 ;
        RECT 84.655 199.375 84.945 199.420 ;
        RECT 85.560 199.375 85.880 199.435 ;
        RECT 84.655 199.235 85.880 199.375 ;
        RECT 84.655 199.190 84.945 199.235 ;
        RECT 85.560 199.175 85.880 199.235 ;
        RECT 100.740 199.175 101.060 199.435 ;
        RECT 80.950 199.035 81.240 199.080 ;
        RECT 77.690 198.895 81.240 199.035 ;
        RECT 77.690 198.850 77.980 198.895 ;
        RECT 79.120 198.835 79.440 198.895 ;
        RECT 80.950 198.850 81.240 198.895 ;
        RECT 81.870 199.035 82.160 199.080 ;
        RECT 83.730 199.035 84.020 199.080 ;
        RECT 81.870 198.895 84.020 199.035 ;
        RECT 81.870 198.850 82.160 198.895 ;
        RECT 83.730 198.850 84.020 198.895 ;
        RECT 90.620 199.035 90.940 199.095 ;
        RECT 96.155 199.035 96.445 199.080 ;
        RECT 99.360 199.035 99.680 199.095 ;
        RECT 90.620 198.895 99.680 199.035 ;
        RECT 90.620 198.835 90.940 198.895 ;
        RECT 96.155 198.850 96.445 198.895 ;
        RECT 99.360 198.835 99.680 198.895 ;
        RECT 58.420 198.695 58.740 198.755 ;
        RECT 75.900 198.740 76.220 198.755 ;
        RECT 53.910 198.555 58.740 198.695 ;
        RECT 46.935 198.510 47.225 198.555 ;
        RECT 47.380 198.495 47.700 198.555 ;
        RECT 58.420 198.495 58.740 198.555 ;
        RECT 75.685 198.510 76.220 198.740 ;
        RECT 75.900 198.495 76.220 198.510 ;
        RECT 96.600 198.495 96.920 198.755 ;
        RECT 101.675 198.695 101.965 198.740 ;
        RECT 102.580 198.695 102.900 198.755 ;
        RECT 101.675 198.555 102.900 198.695 ;
        RECT 101.675 198.510 101.965 198.555 ;
        RECT 102.580 198.495 102.900 198.555 ;
        RECT 10.650 197.875 118.610 198.355 ;
        RECT 57.500 197.475 57.820 197.735 ;
        RECT 58.420 197.475 58.740 197.735 ;
        RECT 59.340 197.475 59.660 197.735 ;
        RECT 62.575 197.490 62.865 197.720 ;
        RECT 63.020 197.675 63.340 197.735 ;
        RECT 79.135 197.675 79.425 197.720 ;
        RECT 63.020 197.535 68.310 197.675 ;
        RECT 40.020 197.380 40.340 197.395 ;
        RECT 34.060 197.335 34.350 197.380 ;
        RECT 35.920 197.335 36.210 197.380 ;
        RECT 34.060 197.195 36.210 197.335 ;
        RECT 34.060 197.150 34.350 197.195 ;
        RECT 35.920 197.150 36.210 197.195 ;
        RECT 36.840 197.335 37.130 197.380 ;
        RECT 40.020 197.335 40.390 197.380 ;
        RECT 36.840 197.195 40.390 197.335 ;
        RECT 36.840 197.150 37.130 197.195 ;
        RECT 40.020 197.150 40.390 197.195 ;
        RECT 45.030 197.335 45.320 197.380 ;
        RECT 47.380 197.335 47.700 197.395 ;
        RECT 48.290 197.335 48.580 197.380 ;
        RECT 45.030 197.195 48.580 197.335 ;
        RECT 45.030 197.150 45.320 197.195 ;
        RECT 35.995 196.995 36.210 197.150 ;
        RECT 40.020 197.135 40.340 197.150 ;
        RECT 47.380 197.135 47.700 197.195 ;
        RECT 48.290 197.150 48.580 197.195 ;
        RECT 49.210 197.335 49.500 197.380 ;
        RECT 51.070 197.335 51.360 197.380 ;
        RECT 49.210 197.195 51.360 197.335 ;
        RECT 59.430 197.335 59.570 197.475 ;
        RECT 62.650 197.335 62.790 197.490 ;
        RECT 63.020 197.475 63.340 197.535 ;
        RECT 68.170 197.380 68.310 197.535 ;
        RECT 79.135 197.535 82.570 197.675 ;
        RECT 79.135 197.490 79.425 197.535 ;
        RECT 67.015 197.335 67.305 197.380 ;
        RECT 59.430 197.195 61.870 197.335 ;
        RECT 62.650 197.195 67.305 197.335 ;
        RECT 49.210 197.150 49.500 197.195 ;
        RECT 51.070 197.150 51.360 197.195 ;
        RECT 38.240 196.995 38.530 197.040 ;
        RECT 35.995 196.855 38.530 196.995 ;
        RECT 38.240 196.810 38.530 196.855 ;
        RECT 46.890 196.995 47.180 197.040 ;
        RECT 49.210 196.995 49.425 197.150 ;
        RECT 61.730 197.055 61.870 197.195 ;
        RECT 67.015 197.150 67.305 197.195 ;
        RECT 68.095 197.150 68.385 197.380 ;
        RECT 81.895 197.335 82.185 197.380 ;
        RECT 76.910 197.195 82.185 197.335 ;
        RECT 46.890 196.855 49.425 196.995 ;
        RECT 46.890 196.810 47.180 196.855 ;
        RECT 50.140 196.795 50.460 197.055 ;
        RECT 56.580 196.995 56.900 197.055 ;
        RECT 57.055 196.995 57.345 197.040 ;
        RECT 58.880 196.995 59.200 197.055 ;
        RECT 56.580 196.855 59.200 196.995 ;
        RECT 56.580 196.795 56.900 196.855 ;
        RECT 57.055 196.810 57.345 196.855 ;
        RECT 58.880 196.795 59.200 196.855 ;
        RECT 59.355 196.810 59.645 197.040 ;
        RECT 33.120 196.455 33.440 196.715 ;
        RECT 34.975 196.655 35.265 196.700 ;
        RECT 44.160 196.655 44.480 196.715 ;
        RECT 34.975 196.515 44.480 196.655 ;
        RECT 34.975 196.470 35.265 196.515 ;
        RECT 44.160 196.455 44.480 196.515 ;
        RECT 44.620 196.655 44.940 196.715 ;
        RECT 51.995 196.655 52.285 196.700 ;
        RECT 52.440 196.655 52.760 196.715 ;
        RECT 44.620 196.515 52.760 196.655 ;
        RECT 59.430 196.655 59.570 196.810 ;
        RECT 60.260 196.795 60.580 197.055 ;
        RECT 60.720 196.795 61.040 197.055 ;
        RECT 61.180 196.795 61.500 197.055 ;
        RECT 61.640 196.795 61.960 197.055 ;
        RECT 63.940 196.795 64.260 197.055 ;
        RECT 64.400 196.995 64.720 197.055 ;
        RECT 65.780 196.995 66.100 197.055 ;
        RECT 64.400 196.855 66.100 196.995 ;
        RECT 64.400 196.795 64.720 196.855 ;
        RECT 65.780 196.795 66.100 196.855 ;
        RECT 74.060 196.795 74.380 197.055 ;
        RECT 75.900 196.995 76.220 197.055 ;
        RECT 76.910 197.040 77.050 197.195 ;
        RECT 81.895 197.150 82.185 197.195 ;
        RECT 76.835 196.995 77.125 197.040 ;
        RECT 75.900 196.855 77.125 196.995 ;
        RECT 75.900 196.795 76.220 196.855 ;
        RECT 76.835 196.810 77.125 196.855 ;
        RECT 77.280 196.795 77.600 197.055 ;
        RECT 82.430 196.995 82.570 197.535 ;
        RECT 83.720 197.475 84.040 197.735 ;
        RECT 84.180 197.475 84.500 197.735 ;
        RECT 94.315 197.335 94.605 197.380 ;
        RECT 96.715 197.335 97.005 197.380 ;
        RECT 99.955 197.335 100.605 197.380 ;
        RECT 94.315 197.195 100.605 197.335 ;
        RECT 94.315 197.150 94.605 197.195 ;
        RECT 96.715 197.150 97.305 197.195 ;
        RECT 99.955 197.150 100.605 197.195 ;
        RECT 85.115 196.995 85.405 197.040 ;
        RECT 82.430 196.855 85.405 196.995 ;
        RECT 85.115 196.810 85.405 196.855 ;
        RECT 93.380 196.995 93.700 197.055 ;
        RECT 93.855 196.995 94.145 197.040 ;
        RECT 93.380 196.855 94.145 196.995 ;
        RECT 93.380 196.795 93.700 196.855 ;
        RECT 93.855 196.810 94.145 196.855 ;
        RECT 97.015 196.835 97.305 197.150 ;
        RECT 102.580 197.135 102.900 197.395 ;
        RECT 98.095 196.995 98.385 197.040 ;
        RECT 101.675 196.995 101.965 197.040 ;
        RECT 103.510 196.995 103.800 197.040 ;
        RECT 98.095 196.855 103.800 196.995 ;
        RECT 98.095 196.810 98.385 196.855 ;
        RECT 101.675 196.810 101.965 196.855 ;
        RECT 103.510 196.810 103.800 196.855 ;
        RECT 103.960 196.795 104.280 197.055 ;
        RECT 59.430 196.515 66.470 196.655 ;
        RECT 44.620 196.455 44.940 196.515 ;
        RECT 51.995 196.470 52.285 196.515 ;
        RECT 52.440 196.455 52.760 196.515 ;
        RECT 66.330 196.360 66.470 196.515 ;
        RECT 74.520 196.455 74.840 196.715 ;
        RECT 76.375 196.470 76.665 196.700 ;
        RECT 80.515 196.470 80.805 196.700 ;
        RECT 81.435 196.655 81.725 196.700 ;
        RECT 92.920 196.655 93.240 196.715 ;
        RECT 81.435 196.515 93.240 196.655 ;
        RECT 81.435 196.470 81.725 196.515 ;
        RECT 33.600 196.315 33.890 196.360 ;
        RECT 35.460 196.315 35.750 196.360 ;
        RECT 38.240 196.315 38.530 196.360 ;
        RECT 33.600 196.175 38.530 196.315 ;
        RECT 33.600 196.130 33.890 196.175 ;
        RECT 35.460 196.130 35.750 196.175 ;
        RECT 38.240 196.130 38.530 196.175 ;
        RECT 42.105 196.315 42.395 196.360 ;
        RECT 46.890 196.315 47.180 196.360 ;
        RECT 49.670 196.315 49.960 196.360 ;
        RECT 51.530 196.315 51.820 196.360 ;
        RECT 42.105 196.175 44.390 196.315 ;
        RECT 42.105 196.130 42.395 196.175 ;
        RECT 44.250 196.035 44.390 196.175 ;
        RECT 46.890 196.175 51.820 196.315 ;
        RECT 46.890 196.130 47.180 196.175 ;
        RECT 49.670 196.130 49.960 196.175 ;
        RECT 51.530 196.130 51.820 196.175 ;
        RECT 66.255 196.130 66.545 196.360 ;
        RECT 67.620 196.315 67.940 196.375 ;
        RECT 66.790 196.175 67.940 196.315 ;
        RECT 43.025 195.975 43.315 196.020 ;
        RECT 43.700 195.975 44.020 196.035 ;
        RECT 43.025 195.835 44.020 195.975 ;
        RECT 43.025 195.790 43.315 195.835 ;
        RECT 43.700 195.775 44.020 195.835 ;
        RECT 44.160 195.775 44.480 196.035 ;
        RECT 61.640 195.975 61.960 196.035 ;
        RECT 63.955 195.975 64.245 196.020 ;
        RECT 66.790 195.975 66.930 196.175 ;
        RECT 67.620 196.115 67.940 196.175 ;
        RECT 73.600 196.315 73.920 196.375 ;
        RECT 76.450 196.315 76.590 196.470 ;
        RECT 80.590 196.315 80.730 196.470 ;
        RECT 92.920 196.455 93.240 196.515 ;
        RECT 91.080 196.315 91.400 196.375 ;
        RECT 73.600 196.175 91.400 196.315 ;
        RECT 73.600 196.115 73.920 196.175 ;
        RECT 91.080 196.115 91.400 196.175 ;
        RECT 98.095 196.315 98.385 196.360 ;
        RECT 101.215 196.315 101.505 196.360 ;
        RECT 103.105 196.315 103.395 196.360 ;
        RECT 98.095 196.175 103.395 196.315 ;
        RECT 98.095 196.130 98.385 196.175 ;
        RECT 101.215 196.130 101.505 196.175 ;
        RECT 103.105 196.130 103.395 196.175 ;
        RECT 61.640 195.835 66.930 195.975 ;
        RECT 67.175 195.975 67.465 196.020 ;
        RECT 68.540 195.975 68.860 196.035 ;
        RECT 67.175 195.835 68.860 195.975 ;
        RECT 61.640 195.775 61.960 195.835 ;
        RECT 63.955 195.790 64.245 195.835 ;
        RECT 67.175 195.790 67.465 195.835 ;
        RECT 68.540 195.775 68.860 195.835 ;
        RECT 94.760 195.975 95.080 196.035 ;
        RECT 95.235 195.975 95.525 196.020 ;
        RECT 94.760 195.835 95.525 195.975 ;
        RECT 94.760 195.775 95.080 195.835 ;
        RECT 95.235 195.790 95.525 195.835 ;
        RECT 11.430 195.155 118.610 195.635 ;
        RECT 46.000 194.755 46.320 195.015 ;
        RECT 49.695 194.955 49.985 195.000 ;
        RECT 50.140 194.955 50.460 195.015 ;
        RECT 49.695 194.815 50.460 194.955 ;
        RECT 49.695 194.770 49.985 194.815 ;
        RECT 50.140 194.755 50.460 194.815 ;
        RECT 63.495 194.955 63.785 195.000 ;
        RECT 63.940 194.955 64.260 195.015 ;
        RECT 63.495 194.815 64.260 194.955 ;
        RECT 63.495 194.770 63.785 194.815 ;
        RECT 63.940 194.755 64.260 194.815 ;
        RECT 64.415 194.770 64.705 195.000 ;
        RECT 79.580 194.955 79.900 195.015 ;
        RECT 81.435 194.955 81.725 195.000 ;
        RECT 79.580 194.815 81.725 194.955 ;
        RECT 30.935 194.615 31.225 194.660 ;
        RECT 34.055 194.615 34.345 194.660 ;
        RECT 35.945 194.615 36.235 194.660 ;
        RECT 64.490 194.615 64.630 194.770 ;
        RECT 79.580 194.755 79.900 194.815 ;
        RECT 81.435 194.770 81.725 194.815 ;
        RECT 100.740 194.955 101.060 195.015 ;
        RECT 102.595 194.955 102.885 195.000 ;
        RECT 100.740 194.815 102.885 194.955 ;
        RECT 100.740 194.755 101.060 194.815 ;
        RECT 102.595 194.770 102.885 194.815 ;
        RECT 66.700 194.615 67.020 194.675 ;
        RECT 75.410 194.615 75.700 194.660 ;
        RECT 78.190 194.615 78.480 194.660 ;
        RECT 80.050 194.615 80.340 194.660 ;
        RECT 30.935 194.475 36.235 194.615 ;
        RECT 30.935 194.430 31.225 194.475 ;
        RECT 34.055 194.430 34.345 194.475 ;
        RECT 35.945 194.430 36.235 194.475 ;
        RECT 60.350 194.475 64.630 194.615 ;
        RECT 65.410 194.475 69.230 194.615 ;
        RECT 36.815 194.275 37.105 194.320 ;
        RECT 40.940 194.275 41.260 194.335 ;
        RECT 36.815 194.135 41.260 194.275 ;
        RECT 36.815 194.090 37.105 194.135 ;
        RECT 40.940 194.075 41.260 194.135 ;
        RECT 43.255 194.275 43.545 194.320 ;
        RECT 48.300 194.275 48.620 194.335 ;
        RECT 43.255 194.135 48.620 194.275 ;
        RECT 43.255 194.090 43.545 194.135 ;
        RECT 48.300 194.075 48.620 194.135 ;
        RECT 60.350 193.995 60.490 194.475 ;
        RECT 65.410 194.275 65.550 194.475 ;
        RECT 66.700 194.415 67.020 194.475 ;
        RECT 64.490 194.135 65.550 194.275 ;
        RECT 65.780 194.275 66.100 194.335 ;
        RECT 69.090 194.320 69.230 194.475 ;
        RECT 75.410 194.475 80.340 194.615 ;
        RECT 75.410 194.430 75.700 194.475 ;
        RECT 78.190 194.430 78.480 194.475 ;
        RECT 80.050 194.430 80.340 194.475 ;
        RECT 86.940 194.615 87.260 194.675 ;
        RECT 88.335 194.615 88.625 194.660 ;
        RECT 86.940 194.475 88.625 194.615 ;
        RECT 86.940 194.415 87.260 194.475 ;
        RECT 88.335 194.430 88.625 194.475 ;
        RECT 65.780 194.135 67.390 194.275 ;
        RECT 29.900 193.955 30.220 193.995 ;
        RECT 29.855 193.735 30.220 193.955 ;
        RECT 30.935 193.935 31.225 193.980 ;
        RECT 34.515 193.935 34.805 193.980 ;
        RECT 36.350 193.935 36.640 193.980 ;
        RECT 30.935 193.795 36.640 193.935 ;
        RECT 30.935 193.750 31.225 193.795 ;
        RECT 34.515 193.750 34.805 193.795 ;
        RECT 36.350 193.750 36.640 193.795 ;
        RECT 38.655 193.935 38.945 193.980 ;
        RECT 40.020 193.935 40.340 193.995 ;
        RECT 38.655 193.795 40.340 193.935 ;
        RECT 38.655 193.750 38.945 193.795 ;
        RECT 40.020 193.735 40.340 193.795 ;
        RECT 43.715 193.935 44.005 193.980 ;
        RECT 44.160 193.935 44.480 193.995 ;
        RECT 43.715 193.795 44.480 193.935 ;
        RECT 43.715 193.750 44.005 193.795 ;
        RECT 44.160 193.735 44.480 193.795 ;
        RECT 48.760 193.735 49.080 193.995 ;
        RECT 60.260 193.735 60.580 193.995 ;
        RECT 60.720 193.935 61.040 193.995 ;
        RECT 64.490 193.980 64.630 194.135 ;
        RECT 65.780 194.075 66.100 194.135 ;
        RECT 64.415 193.935 64.705 193.980 ;
        RECT 66.240 193.935 66.560 193.995 ;
        RECT 67.250 193.980 67.390 194.135 ;
        RECT 69.015 194.090 69.305 194.320 ;
        RECT 80.500 194.275 80.820 194.335 ;
        RECT 85.560 194.275 85.880 194.335 ;
        RECT 80.500 194.135 85.880 194.275 ;
        RECT 80.500 194.075 80.820 194.135 ;
        RECT 85.560 194.075 85.880 194.135 ;
        RECT 91.080 194.275 91.400 194.335 ;
        RECT 95.220 194.275 95.540 194.335 ;
        RECT 99.375 194.275 99.665 194.320 ;
        RECT 91.080 194.135 99.665 194.275 ;
        RECT 91.080 194.075 91.400 194.135 ;
        RECT 95.220 194.075 95.540 194.135 ;
        RECT 99.375 194.090 99.665 194.135 ;
        RECT 60.720 193.795 64.705 193.935 ;
        RECT 60.720 193.735 61.040 193.795 ;
        RECT 64.415 193.750 64.705 193.795 ;
        RECT 64.950 193.795 66.930 193.935 ;
        RECT 29.855 193.640 30.145 193.735 ;
        RECT 29.555 193.595 30.145 193.640 ;
        RECT 32.795 193.595 33.445 193.640 ;
        RECT 29.555 193.455 33.445 193.595 ;
        RECT 29.555 193.410 29.845 193.455 ;
        RECT 32.795 193.410 33.445 193.455 ;
        RECT 35.420 193.395 35.740 193.655 ;
        RECT 61.180 193.595 61.500 193.655 ;
        RECT 64.950 193.595 65.090 193.795 ;
        RECT 66.240 193.735 66.560 193.795 ;
        RECT 61.180 193.455 65.090 193.595 ;
        RECT 66.790 193.595 66.930 193.795 ;
        RECT 67.175 193.750 67.465 193.980 ;
        RECT 67.620 193.735 67.940 193.995 ;
        RECT 75.410 193.935 75.700 193.980 ;
        RECT 75.410 193.795 77.945 193.935 ;
        RECT 75.410 193.750 75.700 193.795 ;
        RECT 73.550 193.595 73.840 193.640 ;
        RECT 74.520 193.595 74.840 193.655 ;
        RECT 77.730 193.640 77.945 193.795 ;
        RECT 78.660 193.735 78.980 193.995 ;
        RECT 81.895 193.935 82.185 193.980 ;
        RECT 82.800 193.935 83.120 193.995 ;
        RECT 81.895 193.795 83.120 193.935 ;
        RECT 81.895 193.750 82.185 193.795 ;
        RECT 82.800 193.735 83.120 193.795 ;
        RECT 76.810 193.595 77.100 193.640 ;
        RECT 66.790 193.455 68.310 193.595 ;
        RECT 61.180 193.395 61.500 193.455 ;
        RECT 28.060 193.255 28.380 193.315 ;
        RECT 31.280 193.255 31.600 193.315 ;
        RECT 28.060 193.115 31.600 193.255 ;
        RECT 28.060 193.055 28.380 193.115 ;
        RECT 31.280 193.055 31.600 193.115 ;
        RECT 39.560 193.055 39.880 193.315 ;
        RECT 43.700 193.255 44.020 193.315 ;
        RECT 44.175 193.255 44.465 193.300 ;
        RECT 43.700 193.115 44.465 193.255 ;
        RECT 43.700 193.055 44.020 193.115 ;
        RECT 44.175 193.070 44.465 193.115 ;
        RECT 63.035 193.255 63.325 193.300 ;
        RECT 67.620 193.255 67.940 193.315 ;
        RECT 68.170 193.300 68.310 193.455 ;
        RECT 73.550 193.455 77.100 193.595 ;
        RECT 73.550 193.410 73.840 193.455 ;
        RECT 74.520 193.395 74.840 193.455 ;
        RECT 76.810 193.410 77.100 193.455 ;
        RECT 77.730 193.595 78.020 193.640 ;
        RECT 79.590 193.595 79.880 193.640 ;
        RECT 77.730 193.455 79.880 193.595 ;
        RECT 77.730 193.410 78.020 193.455 ;
        RECT 79.590 193.410 79.880 193.455 ;
        RECT 85.100 193.595 85.420 193.655 ;
        RECT 90.635 193.595 90.925 193.640 ;
        RECT 85.100 193.455 90.925 193.595 ;
        RECT 85.100 193.395 85.420 193.455 ;
        RECT 90.635 193.410 90.925 193.455 ;
        RECT 93.380 193.595 93.700 193.655 ;
        RECT 96.155 193.595 96.445 193.640 ;
        RECT 100.295 193.595 100.585 193.640 ;
        RECT 93.380 193.455 96.445 193.595 ;
        RECT 93.380 193.395 93.700 193.455 ;
        RECT 96.155 193.410 96.445 193.455 ;
        RECT 96.690 193.455 100.585 193.595 ;
        RECT 63.035 193.115 67.940 193.255 ;
        RECT 63.035 193.070 63.325 193.115 ;
        RECT 67.620 193.055 67.940 193.115 ;
        RECT 68.095 193.070 68.385 193.300 ;
        RECT 68.540 193.055 68.860 193.315 ;
        RECT 71.300 193.300 71.620 193.315 ;
        RECT 71.300 193.070 71.835 193.300 ;
        RECT 88.320 193.255 88.640 193.315 ;
        RECT 90.175 193.255 90.465 193.300 ;
        RECT 88.320 193.115 90.465 193.255 ;
        RECT 71.300 193.055 71.620 193.070 ;
        RECT 88.320 193.055 88.640 193.115 ;
        RECT 90.175 193.070 90.465 193.115 ;
        RECT 94.760 193.255 95.080 193.315 ;
        RECT 96.690 193.300 96.830 193.455 ;
        RECT 100.295 193.410 100.585 193.455 ;
        RECT 96.615 193.255 96.905 193.300 ;
        RECT 94.760 193.115 96.905 193.255 ;
        RECT 94.760 193.055 95.080 193.115 ;
        RECT 96.615 193.070 96.905 193.115 ;
        RECT 97.980 193.255 98.300 193.315 ;
        RECT 98.455 193.255 98.745 193.300 ;
        RECT 97.980 193.115 98.745 193.255 ;
        RECT 97.980 193.055 98.300 193.115 ;
        RECT 98.455 193.070 98.745 193.115 ;
        RECT 99.360 193.255 99.680 193.315 ;
        RECT 100.755 193.255 101.045 193.300 ;
        RECT 99.360 193.115 101.045 193.255 ;
        RECT 99.360 193.055 99.680 193.115 ;
        RECT 100.755 193.070 101.045 193.115 ;
        RECT 10.650 192.435 118.610 192.915 ;
        RECT 19.320 192.235 19.640 192.295 ;
        RECT 19.320 192.095 29.670 192.235 ;
        RECT 19.320 192.035 19.640 192.095 ;
        RECT 23.475 191.895 23.765 191.940 ;
        RECT 25.775 191.895 26.065 191.940 ;
        RECT 23.475 191.755 26.065 191.895 ;
        RECT 23.475 191.710 23.765 191.755 ;
        RECT 25.775 191.710 26.065 191.755 ;
        RECT 20.715 191.555 21.005 191.600 ;
        RECT 28.060 191.555 28.380 191.615 ;
        RECT 29.530 191.600 29.670 192.095 ;
        RECT 29.900 192.035 30.220 192.295 ;
        RECT 43.700 192.235 44.020 192.295 ;
        RECT 46.935 192.235 47.225 192.280 ;
        RECT 43.700 192.095 47.225 192.235 ;
        RECT 43.700 192.035 44.020 192.095 ;
        RECT 46.935 192.050 47.225 192.095 ;
        RECT 48.760 192.235 49.080 192.295 ;
        RECT 49.235 192.235 49.525 192.280 ;
        RECT 67.175 192.235 67.465 192.280 ;
        RECT 48.760 192.095 49.525 192.235 ;
        RECT 48.760 192.035 49.080 192.095 ;
        RECT 49.235 192.050 49.525 192.095 ;
        RECT 65.410 192.095 67.465 192.235 ;
        RECT 31.295 191.895 31.585 191.940 ;
        RECT 33.695 191.895 33.985 191.940 ;
        RECT 36.935 191.895 37.585 191.940 ;
        RECT 31.295 191.755 37.585 191.895 ;
        RECT 31.295 191.710 31.585 191.755 ;
        RECT 33.695 191.710 34.285 191.755 ;
        RECT 36.935 191.710 37.585 191.755 ;
        RECT 20.715 191.415 28.380 191.555 ;
        RECT 20.715 191.370 21.005 191.415 ;
        RECT 28.060 191.355 28.380 191.415 ;
        RECT 29.455 191.555 29.745 191.600 ;
        RECT 30.835 191.555 31.125 191.600 ;
        RECT 29.455 191.415 31.125 191.555 ;
        RECT 29.455 191.370 29.745 191.415 ;
        RECT 30.835 191.370 31.125 191.415 ;
        RECT 33.995 191.395 34.285 191.710 ;
        RECT 39.560 191.695 39.880 191.955 ;
        RECT 46.000 191.895 46.320 191.955 ;
        RECT 47.840 191.895 48.160 191.955 ;
        RECT 65.410 191.940 65.550 192.095 ;
        RECT 67.175 192.050 67.465 192.095 ;
        RECT 71.300 192.235 71.620 192.295 ;
        RECT 74.995 192.235 75.285 192.280 ;
        RECT 77.280 192.235 77.600 192.295 ;
        RECT 71.300 192.095 77.600 192.235 ;
        RECT 71.300 192.035 71.620 192.095 ;
        RECT 74.995 192.050 75.285 192.095 ;
        RECT 77.280 192.035 77.600 192.095 ;
        RECT 78.660 192.035 78.980 192.295 ;
        RECT 57.055 191.895 57.345 191.940 ;
        RECT 59.455 191.895 59.745 191.940 ;
        RECT 62.695 191.895 63.345 191.940 ;
        RECT 46.000 191.755 51.290 191.895 ;
        RECT 46.000 191.695 46.320 191.755 ;
        RECT 47.840 191.695 48.160 191.755 ;
        RECT 35.075 191.555 35.365 191.600 ;
        RECT 38.655 191.555 38.945 191.600 ;
        RECT 40.490 191.555 40.780 191.600 ;
        RECT 35.075 191.415 40.780 191.555 ;
        RECT 35.075 191.370 35.365 191.415 ;
        RECT 38.655 191.370 38.945 191.415 ;
        RECT 40.490 191.370 40.780 191.415 ;
        RECT 47.380 191.355 47.700 191.615 ;
        RECT 51.150 191.600 51.290 191.755 ;
        RECT 57.055 191.755 63.345 191.895 ;
        RECT 57.055 191.710 57.345 191.755 ;
        RECT 59.455 191.710 60.045 191.755 ;
        RECT 62.695 191.710 63.345 191.755 ;
        RECT 65.335 191.710 65.625 191.940 ;
        RECT 80.500 191.895 80.820 191.955 ;
        RECT 66.790 191.755 80.820 191.895 ;
        RECT 51.075 191.370 51.365 191.600 ;
        RECT 51.995 191.370 52.285 191.600 ;
        RECT 24.855 191.030 25.145 191.260 ;
        RECT 25.315 191.215 25.605 191.260 ;
        RECT 25.760 191.215 26.080 191.275 ;
        RECT 30.360 191.215 30.680 191.275 ;
        RECT 25.315 191.075 30.680 191.215 ;
        RECT 25.315 191.030 25.605 191.075 ;
        RECT 24.930 190.875 25.070 191.030 ;
        RECT 25.760 191.015 26.080 191.075 ;
        RECT 30.360 191.015 30.680 191.075 ;
        RECT 40.940 191.215 41.260 191.275 ;
        RECT 44.620 191.215 44.940 191.275 ;
        RECT 40.940 191.075 44.940 191.215 ;
        RECT 40.940 191.015 41.260 191.075 ;
        RECT 44.620 191.015 44.940 191.075 ;
        RECT 46.475 191.215 46.765 191.260 ;
        RECT 48.300 191.215 48.620 191.275 ;
        RECT 46.475 191.075 48.620 191.215 ;
        RECT 46.475 191.030 46.765 191.075 ;
        RECT 48.300 191.015 48.620 191.075 ;
        RECT 50.140 191.215 50.460 191.275 ;
        RECT 52.070 191.215 52.210 191.370 ;
        RECT 56.580 191.355 56.900 191.615 ;
        RECT 59.755 191.395 60.045 191.710 ;
        RECT 66.790 191.600 66.930 191.755 ;
        RECT 80.500 191.695 80.820 191.755 ;
        RECT 83.275 191.895 83.565 191.940 ;
        RECT 85.675 191.895 85.965 191.940 ;
        RECT 88.915 191.895 89.565 191.940 ;
        RECT 83.275 191.755 89.565 191.895 ;
        RECT 83.275 191.710 83.565 191.755 ;
        RECT 85.675 191.710 86.265 191.755 ;
        RECT 88.915 191.710 89.565 191.755 ;
        RECT 91.080 191.895 91.400 191.955 ;
        RECT 91.555 191.895 91.845 191.940 ;
        RECT 91.080 191.755 91.845 191.895 ;
        RECT 60.835 191.555 61.125 191.600 ;
        RECT 64.415 191.555 64.705 191.600 ;
        RECT 66.250 191.555 66.540 191.600 ;
        RECT 60.835 191.415 66.540 191.555 ;
        RECT 60.835 191.370 61.125 191.415 ;
        RECT 64.415 191.370 64.705 191.415 ;
        RECT 66.250 191.370 66.540 191.415 ;
        RECT 66.715 191.370 67.005 191.600 ;
        RECT 67.620 191.555 67.940 191.615 ;
        RECT 69.015 191.555 69.305 191.600 ;
        RECT 67.620 191.415 69.305 191.555 ;
        RECT 67.620 191.355 67.940 191.415 ;
        RECT 69.015 191.370 69.305 191.415 ;
        RECT 73.140 191.555 73.460 191.615 ;
        RECT 75.455 191.555 75.745 191.600 ;
        RECT 77.755 191.555 78.045 191.600 ;
        RECT 73.140 191.415 75.745 191.555 ;
        RECT 73.140 191.355 73.460 191.415 ;
        RECT 75.455 191.370 75.745 191.415 ;
        RECT 77.370 191.415 78.045 191.555 ;
        RECT 50.140 191.075 52.210 191.215 ;
        RECT 50.140 191.015 50.460 191.075 ;
        RECT 68.540 191.015 68.860 191.275 ;
        RECT 73.600 191.215 73.920 191.275 ;
        RECT 74.075 191.215 74.365 191.260 ;
        RECT 73.600 191.075 74.365 191.215 ;
        RECT 73.600 191.015 73.920 191.075 ;
        RECT 74.075 191.030 74.365 191.075 ;
        RECT 34.500 190.875 34.820 190.935 ;
        RECT 77.370 190.920 77.510 191.415 ;
        RECT 77.755 191.370 78.045 191.415 ;
        RECT 82.800 191.355 83.120 191.615 ;
        RECT 85.975 191.395 86.265 191.710 ;
        RECT 91.080 191.695 91.400 191.755 ;
        RECT 91.555 191.710 91.845 191.755 ;
        RECT 94.875 191.895 95.165 191.940 ;
        RECT 98.115 191.895 98.765 191.940 ;
        RECT 94.875 191.755 98.765 191.895 ;
        RECT 94.875 191.710 95.465 191.755 ;
        RECT 98.115 191.710 98.765 191.755 ;
        RECT 95.175 191.615 95.465 191.710 ;
        RECT 87.055 191.555 87.345 191.600 ;
        RECT 90.635 191.555 90.925 191.600 ;
        RECT 92.470 191.555 92.760 191.600 ;
        RECT 87.055 191.415 92.760 191.555 ;
        RECT 87.055 191.370 87.345 191.415 ;
        RECT 90.635 191.370 90.925 191.415 ;
        RECT 92.470 191.370 92.760 191.415 ;
        RECT 95.175 191.395 95.540 191.615 ;
        RECT 95.220 191.355 95.540 191.395 ;
        RECT 96.255 191.555 96.545 191.600 ;
        RECT 99.835 191.555 100.125 191.600 ;
        RECT 101.670 191.555 101.960 191.600 ;
        RECT 96.255 191.415 101.960 191.555 ;
        RECT 96.255 191.370 96.545 191.415 ;
        RECT 99.835 191.370 100.125 191.415 ;
        RECT 101.670 191.370 101.960 191.415 ;
        RECT 102.135 191.555 102.425 191.600 ;
        RECT 103.960 191.555 104.280 191.615 ;
        RECT 102.135 191.415 104.280 191.555 ;
        RECT 102.135 191.370 102.425 191.415 ;
        RECT 103.960 191.355 104.280 191.415 ;
        RECT 109.495 191.555 109.785 191.600 ;
        RECT 110.860 191.555 111.180 191.615 ;
        RECT 109.495 191.415 111.180 191.555 ;
        RECT 109.495 191.370 109.785 191.415 ;
        RECT 110.860 191.355 111.180 191.415 ;
        RECT 85.560 191.215 85.880 191.275 ;
        RECT 92.935 191.215 93.225 191.260 ;
        RECT 85.560 191.075 93.225 191.215 ;
        RECT 85.560 191.015 85.880 191.075 ;
        RECT 92.935 191.030 93.225 191.075 ;
        RECT 98.900 191.215 99.220 191.275 ;
        RECT 100.755 191.215 101.045 191.260 ;
        RECT 98.900 191.075 101.045 191.215 ;
        RECT 98.900 191.015 99.220 191.075 ;
        RECT 100.755 191.030 101.045 191.075 ;
        RECT 24.930 190.735 34.820 190.875 ;
        RECT 34.500 190.675 34.820 190.735 ;
        RECT 35.075 190.875 35.365 190.920 ;
        RECT 38.195 190.875 38.485 190.920 ;
        RECT 40.085 190.875 40.375 190.920 ;
        RECT 35.075 190.735 40.375 190.875 ;
        RECT 35.075 190.690 35.365 190.735 ;
        RECT 38.195 190.690 38.485 190.735 ;
        RECT 40.085 190.690 40.375 190.735 ;
        RECT 60.835 190.875 61.125 190.920 ;
        RECT 63.955 190.875 64.245 190.920 ;
        RECT 65.845 190.875 66.135 190.920 ;
        RECT 60.835 190.735 66.135 190.875 ;
        RECT 60.835 190.690 61.125 190.735 ;
        RECT 63.955 190.690 64.245 190.735 ;
        RECT 65.845 190.690 66.135 190.735 ;
        RECT 77.295 190.690 77.585 190.920 ;
        RECT 87.055 190.875 87.345 190.920 ;
        RECT 90.175 190.875 90.465 190.920 ;
        RECT 92.065 190.875 92.355 190.920 ;
        RECT 87.055 190.735 92.355 190.875 ;
        RECT 87.055 190.690 87.345 190.735 ;
        RECT 90.175 190.690 90.465 190.735 ;
        RECT 92.065 190.690 92.355 190.735 ;
        RECT 96.255 190.875 96.545 190.920 ;
        RECT 99.375 190.875 99.665 190.920 ;
        RECT 101.265 190.875 101.555 190.920 ;
        RECT 96.255 190.735 101.555 190.875 ;
        RECT 96.255 190.690 96.545 190.735 ;
        RECT 99.375 190.690 99.665 190.735 ;
        RECT 101.265 190.690 101.555 190.735 ;
        RECT 26.680 190.535 27.000 190.595 ;
        RECT 27.615 190.535 27.905 190.580 ;
        RECT 26.680 190.395 27.905 190.535 ;
        RECT 26.680 190.335 27.000 190.395 ;
        RECT 27.615 190.350 27.905 190.395 ;
        RECT 32.215 190.535 32.505 190.580 ;
        RECT 35.880 190.535 36.200 190.595 ;
        RECT 32.215 190.395 36.200 190.535 ;
        RECT 32.215 190.350 32.505 190.395 ;
        RECT 35.880 190.335 36.200 190.395 ;
        RECT 49.680 190.535 50.000 190.595 ;
        RECT 50.615 190.535 50.905 190.580 ;
        RECT 49.680 190.395 50.905 190.535 ;
        RECT 49.680 190.335 50.000 190.395 ;
        RECT 50.615 190.350 50.905 190.395 ;
        RECT 52.915 190.535 53.205 190.580 ;
        RECT 53.820 190.535 54.140 190.595 ;
        RECT 52.915 190.395 54.140 190.535 ;
        RECT 52.915 190.350 53.205 190.395 ;
        RECT 53.820 190.335 54.140 190.395 ;
        RECT 57.975 190.535 58.265 190.580 ;
        RECT 60.260 190.535 60.580 190.595 ;
        RECT 63.020 190.535 63.340 190.595 ;
        RECT 57.975 190.395 63.340 190.535 ;
        RECT 57.975 190.350 58.265 190.395 ;
        RECT 60.260 190.335 60.580 190.395 ;
        RECT 63.020 190.335 63.340 190.395 ;
        RECT 84.195 190.535 84.485 190.580 ;
        RECT 85.100 190.535 85.420 190.595 ;
        RECT 84.195 190.395 85.420 190.535 ;
        RECT 84.195 190.350 84.485 190.395 ;
        RECT 85.100 190.335 85.420 190.395 ;
        RECT 93.380 190.335 93.700 190.595 ;
        RECT 109.035 190.535 109.325 190.580 ;
        RECT 109.480 190.535 109.800 190.595 ;
        RECT 109.035 190.395 109.800 190.535 ;
        RECT 109.035 190.350 109.325 190.395 ;
        RECT 109.480 190.335 109.800 190.395 ;
        RECT 11.430 189.715 118.610 190.195 ;
        RECT 20.715 189.515 21.005 189.560 ;
        RECT 25.760 189.515 26.080 189.575 ;
        RECT 20.715 189.375 26.080 189.515 ;
        RECT 20.715 189.330 21.005 189.375 ;
        RECT 25.760 189.315 26.080 189.375 ;
        RECT 31.755 189.515 32.045 189.560 ;
        RECT 35.420 189.515 35.740 189.575 ;
        RECT 31.755 189.375 35.740 189.515 ;
        RECT 31.755 189.330 32.045 189.375 ;
        RECT 35.420 189.315 35.740 189.375 ;
        RECT 40.020 189.315 40.340 189.575 ;
        RECT 78.660 189.515 78.980 189.575 ;
        RECT 82.800 189.515 83.120 189.575 ;
        RECT 78.660 189.375 83.120 189.515 ;
        RECT 78.660 189.315 78.980 189.375 ;
        RECT 82.800 189.315 83.120 189.375 ;
        RECT 88.320 189.315 88.640 189.575 ;
        RECT 94.775 189.515 95.065 189.560 ;
        RECT 95.220 189.515 95.540 189.575 ;
        RECT 94.775 189.375 95.540 189.515 ;
        RECT 94.775 189.330 95.065 189.375 ;
        RECT 95.220 189.315 95.540 189.375 ;
        RECT 98.900 189.315 99.220 189.575 ;
        RECT 23.575 189.175 23.865 189.220 ;
        RECT 26.695 189.175 26.985 189.220 ;
        RECT 28.585 189.175 28.875 189.220 ;
        RECT 23.575 189.035 28.875 189.175 ;
        RECT 23.575 188.990 23.865 189.035 ;
        RECT 26.695 188.990 26.985 189.035 ;
        RECT 28.585 188.990 28.875 189.035 ;
        RECT 31.280 189.175 31.600 189.235 ;
        RECT 50.570 189.175 50.860 189.220 ;
        RECT 53.350 189.175 53.640 189.220 ;
        RECT 55.210 189.175 55.500 189.220 ;
        RECT 31.280 189.035 34.730 189.175 ;
        RECT 31.280 188.975 31.600 189.035 ;
        RECT 29.440 188.835 29.760 188.895 ;
        RECT 33.120 188.835 33.440 188.895 ;
        RECT 34.590 188.880 34.730 189.035 ;
        RECT 50.570 189.035 55.500 189.175 ;
        RECT 50.570 188.990 50.860 189.035 ;
        RECT 53.350 188.990 53.640 189.035 ;
        RECT 55.210 188.990 55.500 189.035 ;
        RECT 87.875 189.175 88.165 189.220 ;
        RECT 91.080 189.175 91.400 189.235 ;
        RECT 87.875 189.035 91.400 189.175 ;
        RECT 87.875 188.990 88.165 189.035 ;
        RECT 91.080 188.975 91.400 189.035 ;
        RECT 102.580 189.175 102.900 189.235 ;
        RECT 105.815 189.175 106.105 189.220 ;
        RECT 102.580 189.035 106.105 189.175 ;
        RECT 102.580 188.975 102.900 189.035 ;
        RECT 105.815 188.990 106.105 189.035 ;
        RECT 108.675 189.175 108.965 189.220 ;
        RECT 111.795 189.175 112.085 189.220 ;
        RECT 113.685 189.175 113.975 189.220 ;
        RECT 108.675 189.035 113.975 189.175 ;
        RECT 108.675 188.990 108.965 189.035 ;
        RECT 111.795 188.990 112.085 189.035 ;
        RECT 113.685 188.990 113.975 189.035 ;
        RECT 29.440 188.695 33.440 188.835 ;
        RECT 29.440 188.635 29.760 188.695 ;
        RECT 33.120 188.635 33.440 188.695 ;
        RECT 34.515 188.650 34.805 188.880 ;
        RECT 34.960 188.835 35.280 188.895 ;
        RECT 35.435 188.835 35.725 188.880 ;
        RECT 37.275 188.835 37.565 188.880 ;
        RECT 48.300 188.835 48.620 188.895 ;
        RECT 34.960 188.695 48.620 188.835 ;
        RECT 34.960 188.635 35.280 188.695 ;
        RECT 35.435 188.650 35.725 188.695 ;
        RECT 37.275 188.650 37.565 188.695 ;
        RECT 48.300 188.635 48.620 188.695 ;
        RECT 53.820 188.635 54.140 188.895 ;
        RECT 56.580 188.835 56.900 188.895 ;
        RECT 64.875 188.835 65.165 188.880 ;
        RECT 56.580 188.695 65.165 188.835 ;
        RECT 56.580 188.635 56.900 188.695 ;
        RECT 64.875 188.650 65.165 188.695 ;
        RECT 73.600 188.835 73.920 188.895 ;
        RECT 82.815 188.835 83.105 188.880 ;
        RECT 110.860 188.835 111.180 188.895 ;
        RECT 73.600 188.695 83.105 188.835 ;
        RECT 73.600 188.635 73.920 188.695 ;
        RECT 82.815 188.650 83.105 188.695 ;
        RECT 100.830 188.695 111.180 188.835 ;
        RECT 19.320 188.295 19.640 188.555 ;
        RECT 22.495 188.200 22.785 188.515 ;
        RECT 23.575 188.495 23.865 188.540 ;
        RECT 27.155 188.495 27.445 188.540 ;
        RECT 28.990 188.495 29.280 188.540 ;
        RECT 23.575 188.355 29.280 188.495 ;
        RECT 23.575 188.310 23.865 188.355 ;
        RECT 27.155 188.310 27.445 188.355 ;
        RECT 28.990 188.310 29.280 188.355 ;
        RECT 30.835 188.495 31.125 188.540 ;
        RECT 45.095 188.495 45.385 188.540 ;
        RECT 46.000 188.495 46.320 188.555 ;
        RECT 30.835 188.355 32.430 188.495 ;
        RECT 30.835 188.310 31.125 188.355 ;
        RECT 19.795 188.155 20.085 188.200 ;
        RECT 22.195 188.155 22.785 188.200 ;
        RECT 25.435 188.155 26.085 188.200 ;
        RECT 19.795 188.015 26.085 188.155 ;
        RECT 19.795 187.970 20.085 188.015 ;
        RECT 22.195 187.970 22.485 188.015 ;
        RECT 25.435 187.970 26.085 188.015 ;
        RECT 28.060 187.955 28.380 188.215 ;
        RECT 32.290 187.860 32.430 188.355 ;
        RECT 45.095 188.355 46.320 188.495 ;
        RECT 45.095 188.310 45.385 188.355 ;
        RECT 46.000 188.295 46.320 188.355 ;
        RECT 50.570 188.495 50.860 188.540 ;
        RECT 50.570 188.355 53.105 188.495 ;
        RECT 50.570 188.310 50.860 188.355 ;
        RECT 38.195 188.155 38.485 188.200 ;
        RECT 44.160 188.155 44.480 188.215 ;
        RECT 46.705 188.155 46.995 188.200 ;
        RECT 47.840 188.155 48.160 188.215 ;
        RECT 38.195 188.015 44.480 188.155 ;
        RECT 38.195 187.970 38.485 188.015 ;
        RECT 44.160 187.955 44.480 188.015 ;
        RECT 45.170 188.015 48.160 188.155 ;
        RECT 32.215 187.630 32.505 187.860 ;
        RECT 34.055 187.815 34.345 187.860 ;
        RECT 35.880 187.815 36.200 187.875 ;
        RECT 37.735 187.815 38.025 187.860 ;
        RECT 34.055 187.675 38.025 187.815 ;
        RECT 34.055 187.630 34.345 187.675 ;
        RECT 35.880 187.615 36.200 187.675 ;
        RECT 37.735 187.630 38.025 187.675 ;
        RECT 42.780 187.815 43.100 187.875 ;
        RECT 45.170 187.815 45.310 188.015 ;
        RECT 46.705 187.970 46.995 188.015 ;
        RECT 47.840 187.955 48.160 188.015 ;
        RECT 48.710 188.155 49.000 188.200 ;
        RECT 49.680 188.155 50.000 188.215 ;
        RECT 52.890 188.200 53.105 188.355 ;
        RECT 55.660 188.295 55.980 188.555 ;
        RECT 62.560 188.495 62.880 188.555 ;
        RECT 63.955 188.495 64.245 188.540 ;
        RECT 62.560 188.355 64.245 188.495 ;
        RECT 62.560 188.295 62.880 188.355 ;
        RECT 63.955 188.310 64.245 188.355 ;
        RECT 74.060 188.495 74.380 188.555 ;
        RECT 74.995 188.495 75.285 188.540 ;
        RECT 78.660 188.495 78.980 188.555 ;
        RECT 74.060 188.355 78.980 188.495 ;
        RECT 74.060 188.295 74.380 188.355 ;
        RECT 74.995 188.310 75.285 188.355 ;
        RECT 78.660 188.295 78.980 188.355 ;
        RECT 80.960 188.295 81.280 188.555 ;
        RECT 86.940 188.295 87.260 188.555 ;
        RECT 90.160 188.495 90.480 188.555 ;
        RECT 91.095 188.495 91.385 188.540 ;
        RECT 93.380 188.495 93.700 188.555 ;
        RECT 90.160 188.355 93.700 188.495 ;
        RECT 90.160 188.295 90.480 188.355 ;
        RECT 91.095 188.310 91.385 188.355 ;
        RECT 93.380 188.295 93.700 188.355 ;
        RECT 93.840 188.495 94.160 188.555 ;
        RECT 94.315 188.495 94.605 188.540 ;
        RECT 93.840 188.355 94.605 188.495 ;
        RECT 93.840 188.295 94.160 188.355 ;
        RECT 94.315 188.310 94.605 188.355 ;
        RECT 97.980 188.295 98.300 188.555 ;
        RECT 100.280 188.495 100.600 188.555 ;
        RECT 100.830 188.540 100.970 188.695 ;
        RECT 110.860 188.635 111.180 188.695 ;
        RECT 100.755 188.495 101.045 188.540 ;
        RECT 100.280 188.355 101.045 188.495 ;
        RECT 100.280 188.295 100.600 188.355 ;
        RECT 100.755 188.310 101.045 188.355 ;
        RECT 102.595 188.495 102.885 188.540 ;
        RECT 103.040 188.495 103.360 188.555 ;
        RECT 102.595 188.355 103.360 188.495 ;
        RECT 102.595 188.310 102.885 188.355 ;
        RECT 103.040 188.295 103.360 188.355 ;
        RECT 51.970 188.155 52.260 188.200 ;
        RECT 48.710 188.015 52.260 188.155 ;
        RECT 48.710 187.970 49.000 188.015 ;
        RECT 49.680 187.955 50.000 188.015 ;
        RECT 51.970 187.970 52.260 188.015 ;
        RECT 52.890 188.155 53.180 188.200 ;
        RECT 54.750 188.155 55.040 188.200 ;
        RECT 52.890 188.015 55.040 188.155 ;
        RECT 52.890 187.970 53.180 188.015 ;
        RECT 54.750 187.970 55.040 188.015 ;
        RECT 79.120 187.955 79.440 188.215 ;
        RECT 79.580 188.155 79.900 188.215 ;
        RECT 107.595 188.200 107.885 188.515 ;
        RECT 108.675 188.495 108.965 188.540 ;
        RECT 112.255 188.495 112.545 188.540 ;
        RECT 114.090 188.495 114.380 188.540 ;
        RECT 108.675 188.355 114.380 188.495 ;
        RECT 108.675 188.310 108.965 188.355 ;
        RECT 112.255 188.310 112.545 188.355 ;
        RECT 114.090 188.310 114.380 188.355 ;
        RECT 114.540 188.295 114.860 188.555 ;
        RECT 83.735 188.155 84.025 188.200 ;
        RECT 79.580 188.015 84.025 188.155 ;
        RECT 79.580 187.955 79.900 188.015 ;
        RECT 83.735 187.970 84.025 188.015 ;
        RECT 107.295 188.155 107.885 188.200 ;
        RECT 109.480 188.155 109.800 188.215 ;
        RECT 110.535 188.155 111.185 188.200 ;
        RECT 107.295 188.015 111.185 188.155 ;
        RECT 107.295 187.970 107.585 188.015 ;
        RECT 109.480 187.955 109.800 188.015 ;
        RECT 110.535 187.970 111.185 188.015 ;
        RECT 113.160 187.955 113.480 188.215 ;
        RECT 42.780 187.675 45.310 187.815 ;
        RECT 42.780 187.615 43.100 187.675 ;
        RECT 45.540 187.615 45.860 187.875 ;
        RECT 74.520 187.615 74.840 187.875 ;
        RECT 77.740 187.815 78.060 187.875 ;
        RECT 80.055 187.815 80.345 187.860 ;
        RECT 77.740 187.675 80.345 187.815 ;
        RECT 77.740 187.615 78.060 187.675 ;
        RECT 80.055 187.630 80.345 187.675 ;
        RECT 84.195 187.815 84.485 187.860 ;
        RECT 85.100 187.815 85.420 187.875 ;
        RECT 84.195 187.675 85.420 187.815 ;
        RECT 84.195 187.630 84.485 187.675 ;
        RECT 85.100 187.615 85.420 187.675 ;
        RECT 86.035 187.815 86.325 187.860 ;
        RECT 88.320 187.815 88.640 187.875 ;
        RECT 86.035 187.675 88.640 187.815 ;
        RECT 86.035 187.630 86.325 187.675 ;
        RECT 88.320 187.615 88.640 187.675 ;
        RECT 101.200 187.615 101.520 187.875 ;
        RECT 105.355 187.815 105.645 187.860 ;
        RECT 106.260 187.815 106.580 187.875 ;
        RECT 105.355 187.675 106.580 187.815 ;
        RECT 105.355 187.630 105.645 187.675 ;
        RECT 106.260 187.615 106.580 187.675 ;
        RECT 10.650 186.995 118.610 187.475 ;
        RECT 27.615 186.795 27.905 186.840 ;
        RECT 28.060 186.795 28.380 186.855 ;
        RECT 27.615 186.655 28.380 186.795 ;
        RECT 27.615 186.610 27.905 186.655 ;
        RECT 28.060 186.595 28.380 186.655 ;
        RECT 47.840 186.795 48.160 186.855 ;
        RECT 49.235 186.795 49.525 186.840 ;
        RECT 47.840 186.655 49.525 186.795 ;
        RECT 47.840 186.595 48.160 186.655 ;
        RECT 49.235 186.610 49.525 186.655 ;
        RECT 50.140 186.795 50.460 186.855 ;
        RECT 51.535 186.795 51.825 186.840 ;
        RECT 50.140 186.655 51.825 186.795 ;
        RECT 50.140 186.595 50.460 186.655 ;
        RECT 51.535 186.610 51.825 186.655 ;
        RECT 61.640 186.795 61.960 186.855 ;
        RECT 65.320 186.795 65.640 186.855 ;
        RECT 61.640 186.655 65.640 186.795 ;
        RECT 61.640 186.595 61.960 186.655 ;
        RECT 65.320 186.595 65.640 186.655 ;
        RECT 104.895 186.610 105.185 186.840 ;
        RECT 113.160 186.795 113.480 186.855 ;
        RECT 115.015 186.795 115.305 186.840 ;
        RECT 106.350 186.655 112.010 186.795 ;
        RECT 48.760 186.455 49.080 186.515 ;
        RECT 49.695 186.455 49.985 186.500 ;
        RECT 66.700 186.455 67.020 186.515 ;
        RECT 69.000 186.455 69.320 186.515 ;
        RECT 48.760 186.315 49.985 186.455 ;
        RECT 48.760 186.255 49.080 186.315 ;
        RECT 49.695 186.270 49.985 186.315 ;
        RECT 65.870 186.315 69.320 186.455 ;
        RECT 65.870 186.175 66.010 186.315 ;
        RECT 66.700 186.255 67.020 186.315 ;
        RECT 69.000 186.255 69.320 186.315 ;
        RECT 71.875 186.455 72.165 186.500 ;
        RECT 74.520 186.455 74.840 186.515 ;
        RECT 75.115 186.455 75.765 186.500 ;
        RECT 71.875 186.315 75.765 186.455 ;
        RECT 71.875 186.270 72.465 186.315 ;
        RECT 26.680 185.915 27.000 186.175 ;
        RECT 38.655 186.115 38.945 186.160 ;
        RECT 39.100 186.115 39.420 186.175 ;
        RECT 38.655 185.975 39.420 186.115 ;
        RECT 38.655 185.930 38.945 185.975 ;
        RECT 39.100 185.915 39.420 185.975 ;
        RECT 50.140 186.115 50.460 186.175 ;
        RECT 51.995 186.115 52.285 186.160 ;
        RECT 50.140 185.975 52.285 186.115 ;
        RECT 50.140 185.915 50.460 185.975 ;
        RECT 51.995 185.930 52.285 185.975 ;
        RECT 60.720 186.115 61.040 186.175 ;
        RECT 63.480 186.115 63.800 186.175 ;
        RECT 64.860 186.115 65.180 186.175 ;
        RECT 60.720 185.975 65.180 186.115 ;
        RECT 60.720 185.915 61.040 185.975 ;
        RECT 63.480 185.915 63.800 185.975 ;
        RECT 64.860 185.915 65.180 185.975 ;
        RECT 65.320 185.915 65.640 186.175 ;
        RECT 65.780 185.915 66.100 186.175 ;
        RECT 66.240 185.915 66.560 186.175 ;
        RECT 67.635 185.930 67.925 186.160 ;
        RECT 72.175 185.955 72.465 186.270 ;
        RECT 74.520 186.255 74.840 186.315 ;
        RECT 75.115 186.270 75.765 186.315 ;
        RECT 77.740 186.255 78.060 186.515 ;
        RECT 79.120 186.455 79.440 186.515 ;
        RECT 81.535 186.455 81.825 186.500 ;
        RECT 84.775 186.455 85.425 186.500 ;
        RECT 79.120 186.315 85.425 186.455 ;
        RECT 79.120 186.255 79.440 186.315 ;
        RECT 81.535 186.270 82.125 186.315 ;
        RECT 84.775 186.270 85.425 186.315 ;
        RECT 73.255 186.115 73.545 186.160 ;
        RECT 76.835 186.115 77.125 186.160 ;
        RECT 78.670 186.115 78.960 186.160 ;
        RECT 73.255 185.975 78.960 186.115 ;
        RECT 73.255 185.930 73.545 185.975 ;
        RECT 76.835 185.930 77.125 185.975 ;
        RECT 78.670 185.930 78.960 185.975 ;
        RECT 81.835 185.955 82.125 186.270 ;
        RECT 87.400 186.255 87.720 186.515 ;
        RECT 103.040 186.255 103.360 186.515 ;
        RECT 104.970 186.455 105.110 186.610 ;
        RECT 106.350 186.455 106.490 186.655 ;
        RECT 104.970 186.315 106.490 186.455 ;
        RECT 107.295 186.455 107.585 186.500 ;
        RECT 110.535 186.455 111.185 186.500 ;
        RECT 107.295 186.315 111.185 186.455 ;
        RECT 111.870 186.455 112.010 186.655 ;
        RECT 113.160 186.655 115.305 186.795 ;
        RECT 113.160 186.595 113.480 186.655 ;
        RECT 115.015 186.610 115.305 186.655 ;
        RECT 111.870 186.315 116.150 186.455 ;
        RECT 107.295 186.270 107.885 186.315 ;
        RECT 110.535 186.270 111.185 186.315 ;
        RECT 82.915 186.115 83.205 186.160 ;
        RECT 86.495 186.115 86.785 186.160 ;
        RECT 88.330 186.115 88.620 186.160 ;
        RECT 82.915 185.975 88.620 186.115 ;
        RECT 82.915 185.930 83.205 185.975 ;
        RECT 86.495 185.930 86.785 185.975 ;
        RECT 88.330 185.930 88.620 185.975 ;
        RECT 48.300 185.575 48.620 185.835 ;
        RECT 62.560 185.775 62.880 185.835 ;
        RECT 67.710 185.775 67.850 185.930 ;
        RECT 100.280 185.915 100.600 186.175 ;
        RECT 101.200 186.115 101.520 186.175 ;
        RECT 107.595 186.115 107.885 186.270 ;
        RECT 116.010 186.160 116.150 186.315 ;
        RECT 101.200 185.975 107.885 186.115 ;
        RECT 101.200 185.915 101.520 185.975 ;
        RECT 107.595 185.955 107.885 185.975 ;
        RECT 108.675 186.115 108.965 186.160 ;
        RECT 112.255 186.115 112.545 186.160 ;
        RECT 114.090 186.115 114.380 186.160 ;
        RECT 108.675 185.975 114.380 186.115 ;
        RECT 108.675 185.930 108.965 185.975 ;
        RECT 112.255 185.930 112.545 185.975 ;
        RECT 114.090 185.930 114.380 185.975 ;
        RECT 115.935 185.930 116.225 186.160 ;
        RECT 62.560 185.635 67.850 185.775 ;
        RECT 69.015 185.775 69.305 185.820 ;
        RECT 74.060 185.775 74.380 185.835 ;
        RECT 69.015 185.635 74.380 185.775 ;
        RECT 62.560 185.575 62.880 185.635 ;
        RECT 69.015 185.590 69.305 185.635 ;
        RECT 74.060 185.575 74.380 185.635 ;
        RECT 79.135 185.775 79.425 185.820 ;
        RECT 85.560 185.775 85.880 185.835 ;
        RECT 88.795 185.775 89.085 185.820 ;
        RECT 79.135 185.635 89.085 185.775 ;
        RECT 79.135 185.590 79.425 185.635 ;
        RECT 85.560 185.575 85.880 185.635 ;
        RECT 88.795 185.590 89.085 185.635 ;
        RECT 102.120 185.575 102.440 185.835 ;
        RECT 102.580 185.575 102.900 185.835 ;
        RECT 113.160 185.575 113.480 185.835 ;
        RECT 114.540 185.775 114.860 185.835 ;
        RECT 116.380 185.775 116.700 185.835 ;
        RECT 114.540 185.635 116.700 185.775 ;
        RECT 114.540 185.575 114.860 185.635 ;
        RECT 116.380 185.575 116.700 185.635 ;
        RECT 73.255 185.435 73.545 185.480 ;
        RECT 76.375 185.435 76.665 185.480 ;
        RECT 78.265 185.435 78.555 185.480 ;
        RECT 73.255 185.295 78.555 185.435 ;
        RECT 73.255 185.250 73.545 185.295 ;
        RECT 76.375 185.250 76.665 185.295 ;
        RECT 78.265 185.250 78.555 185.295 ;
        RECT 82.915 185.435 83.205 185.480 ;
        RECT 86.035 185.435 86.325 185.480 ;
        RECT 87.925 185.435 88.215 185.480 ;
        RECT 82.915 185.295 88.215 185.435 ;
        RECT 82.915 185.250 83.205 185.295 ;
        RECT 86.035 185.250 86.325 185.295 ;
        RECT 87.925 185.250 88.215 185.295 ;
        RECT 108.675 185.435 108.965 185.480 ;
        RECT 111.795 185.435 112.085 185.480 ;
        RECT 113.685 185.435 113.975 185.480 ;
        RECT 108.675 185.295 113.975 185.435 ;
        RECT 108.675 185.250 108.965 185.295 ;
        RECT 111.795 185.250 112.085 185.295 ;
        RECT 113.685 185.250 113.975 185.295 ;
        RECT 44.620 185.095 44.940 185.155 ;
        RECT 45.095 185.095 45.385 185.140 ;
        RECT 44.620 184.955 45.385 185.095 ;
        RECT 44.620 184.895 44.940 184.955 ;
        RECT 45.095 184.910 45.385 184.955 ;
        RECT 52.915 185.095 53.205 185.140 ;
        RECT 53.360 185.095 53.680 185.155 ;
        RECT 52.915 184.955 53.680 185.095 ;
        RECT 52.915 184.910 53.205 184.955 ;
        RECT 53.360 184.895 53.680 184.955 ;
        RECT 59.800 185.095 60.120 185.155 ;
        RECT 63.955 185.095 64.245 185.140 ;
        RECT 59.800 184.955 64.245 185.095 ;
        RECT 59.800 184.895 60.120 184.955 ;
        RECT 63.955 184.910 64.245 184.955 ;
        RECT 65.320 185.095 65.640 185.155 ;
        RECT 69.460 185.095 69.780 185.155 ;
        RECT 65.320 184.955 69.780 185.095 ;
        RECT 65.320 184.895 65.640 184.955 ;
        RECT 69.460 184.895 69.780 184.955 ;
        RECT 70.395 185.095 70.685 185.140 ;
        RECT 72.680 185.095 73.000 185.155 ;
        RECT 70.395 184.955 73.000 185.095 ;
        RECT 70.395 184.910 70.685 184.955 ;
        RECT 72.680 184.895 73.000 184.955 ;
        RECT 74.060 185.095 74.380 185.155 ;
        RECT 79.580 185.095 79.900 185.155 ;
        RECT 80.055 185.095 80.345 185.140 ;
        RECT 74.060 184.955 80.345 185.095 ;
        RECT 74.060 184.895 74.380 184.955 ;
        RECT 79.580 184.895 79.900 184.955 ;
        RECT 80.055 184.910 80.345 184.955 ;
        RECT 98.440 185.095 98.760 185.155 ;
        RECT 99.835 185.095 100.125 185.140 ;
        RECT 98.440 184.955 100.125 185.095 ;
        RECT 98.440 184.895 98.760 184.955 ;
        RECT 99.835 184.910 100.125 184.955 ;
        RECT 103.040 185.095 103.360 185.155 ;
        RECT 105.815 185.095 106.105 185.140 ;
        RECT 106.720 185.095 107.040 185.155 ;
        RECT 103.040 184.955 107.040 185.095 ;
        RECT 103.040 184.895 103.360 184.955 ;
        RECT 105.815 184.910 106.105 184.955 ;
        RECT 106.720 184.895 107.040 184.955 ;
        RECT 11.430 184.275 118.610 184.755 ;
        RECT 48.300 184.075 48.620 184.135 ;
        RECT 61.180 184.075 61.500 184.135 ;
        RECT 39.190 183.935 48.620 184.075 ;
        RECT 27.255 183.735 27.545 183.780 ;
        RECT 30.375 183.735 30.665 183.780 ;
        RECT 32.265 183.735 32.555 183.780 ;
        RECT 27.255 183.595 32.555 183.735 ;
        RECT 27.255 183.550 27.545 183.595 ;
        RECT 30.375 183.550 30.665 183.595 ;
        RECT 32.265 183.550 32.555 183.595 ;
        RECT 33.120 183.195 33.440 183.455 ;
        RECT 34.040 183.395 34.360 183.455 ;
        RECT 37.735 183.395 38.025 183.440 ;
        RECT 39.190 183.395 39.330 183.935 ;
        RECT 48.300 183.875 48.620 183.935 ;
        RECT 59.430 183.935 61.500 184.075 ;
        RECT 40.495 183.550 40.785 183.780 ;
        RECT 46.000 183.735 46.320 183.795 ;
        RECT 49.220 183.735 49.540 183.795 ;
        RECT 43.790 183.595 49.540 183.735 ;
        RECT 34.040 183.255 39.330 183.395 ;
        RECT 34.040 183.195 34.360 183.255 ;
        RECT 37.735 183.210 38.025 183.255 ;
        RECT 20.700 183.055 21.020 183.115 ;
        RECT 26.175 183.055 26.465 183.075 ;
        RECT 20.700 182.915 26.465 183.055 ;
        RECT 20.700 182.855 21.020 182.915 ;
        RECT 26.175 182.760 26.465 182.915 ;
        RECT 27.255 183.055 27.545 183.100 ;
        RECT 30.835 183.055 31.125 183.100 ;
        RECT 32.670 183.055 32.960 183.100 ;
        RECT 27.255 182.915 32.960 183.055 ;
        RECT 40.570 183.055 40.710 183.550 ;
        RECT 42.335 183.055 42.625 183.100 ;
        RECT 40.570 182.915 42.625 183.055 ;
        RECT 27.255 182.870 27.545 182.915 ;
        RECT 30.835 182.870 31.125 182.915 ;
        RECT 32.670 182.870 32.960 182.915 ;
        RECT 42.335 182.870 42.625 182.915 ;
        RECT 43.240 182.855 43.560 183.115 ;
        RECT 43.790 183.100 43.930 183.595 ;
        RECT 46.000 183.535 46.320 183.595 ;
        RECT 49.220 183.535 49.540 183.595 ;
        RECT 50.110 183.735 50.400 183.780 ;
        RECT 52.890 183.735 53.180 183.780 ;
        RECT 54.750 183.735 55.040 183.780 ;
        RECT 50.110 183.595 55.040 183.735 ;
        RECT 50.110 183.550 50.400 183.595 ;
        RECT 52.890 183.550 53.180 183.595 ;
        RECT 54.750 183.550 55.040 183.595 ;
        RECT 44.710 183.255 53.130 183.395 ;
        RECT 44.710 183.115 44.850 183.255 ;
        RECT 43.715 182.870 44.005 183.100 ;
        RECT 44.620 182.855 44.940 183.115 ;
        RECT 50.110 183.055 50.400 183.100 ;
        RECT 52.990 183.055 53.130 183.255 ;
        RECT 53.360 183.195 53.680 183.455 ;
        RECT 59.430 183.440 59.570 183.935 ;
        RECT 61.180 183.875 61.500 183.935 ;
        RECT 64.860 184.075 65.180 184.135 ;
        RECT 75.455 184.075 75.745 184.120 ;
        RECT 80.960 184.075 81.280 184.135 ;
        RECT 64.860 183.935 68.770 184.075 ;
        RECT 64.860 183.875 65.180 183.935 ;
        RECT 62.575 183.735 62.865 183.780 ;
        RECT 66.700 183.735 67.020 183.795 ;
        RECT 59.890 183.595 67.020 183.735 ;
        RECT 59.890 183.440 60.030 183.595 ;
        RECT 62.575 183.550 62.865 183.595 ;
        RECT 66.700 183.535 67.020 183.595 ;
        RECT 59.355 183.210 59.645 183.440 ;
        RECT 59.815 183.210 60.105 183.440 ;
        RECT 60.720 183.195 61.040 183.455 ;
        RECT 61.180 183.395 61.500 183.455 ;
        RECT 65.335 183.395 65.625 183.440 ;
        RECT 65.780 183.395 66.100 183.455 ;
        RECT 61.180 183.255 66.100 183.395 ;
        RECT 61.180 183.195 61.500 183.255 ;
        RECT 65.335 183.210 65.625 183.255 ;
        RECT 65.780 183.195 66.100 183.255 ;
        RECT 66.255 183.395 66.545 183.440 ;
        RECT 67.160 183.395 67.480 183.455 ;
        RECT 68.630 183.440 68.770 183.935 ;
        RECT 75.455 183.935 81.280 184.075 ;
        RECT 75.455 183.890 75.745 183.935 ;
        RECT 80.960 183.875 81.280 183.935 ;
        RECT 82.800 184.075 83.120 184.135 ;
        RECT 82.800 183.935 86.710 184.075 ;
        RECT 82.800 183.875 83.120 183.935 ;
        RECT 78.215 183.735 78.505 183.780 ;
        RECT 86.020 183.735 86.340 183.795 ;
        RECT 78.215 183.595 86.340 183.735 ;
        RECT 86.570 183.735 86.710 183.935 ;
        RECT 87.400 183.875 87.720 184.135 ;
        RECT 100.280 184.075 100.600 184.135 ;
        RECT 90.250 183.935 100.600 184.075 ;
        RECT 90.250 183.735 90.390 183.935 ;
        RECT 100.280 183.875 100.600 183.935 ;
        RECT 102.120 184.075 102.440 184.135 ;
        RECT 106.260 184.075 106.580 184.135 ;
        RECT 111.795 184.075 112.085 184.120 ;
        RECT 113.160 184.075 113.480 184.135 ;
        RECT 102.120 183.935 105.110 184.075 ;
        RECT 102.120 183.875 102.440 183.935 ;
        RECT 86.570 183.595 90.390 183.735 ;
        RECT 78.215 183.550 78.505 183.595 ;
        RECT 86.020 183.535 86.340 183.595 ;
        RECT 66.255 183.255 67.480 183.395 ;
        RECT 66.255 183.210 66.545 183.255 ;
        RECT 67.160 183.195 67.480 183.255 ;
        RECT 68.555 183.210 68.845 183.440 ;
        RECT 69.000 183.195 69.320 183.455 ;
        RECT 69.460 183.195 69.780 183.455 ;
        RECT 72.695 183.395 72.985 183.440 ;
        RECT 73.600 183.395 73.920 183.455 ;
        RECT 72.695 183.255 73.920 183.395 ;
        RECT 72.695 183.210 72.985 183.255 ;
        RECT 73.600 183.195 73.920 183.255 ;
        RECT 55.215 183.055 55.505 183.100 ;
        RECT 55.660 183.055 55.980 183.115 ;
        RECT 50.110 182.915 52.645 183.055 ;
        RECT 52.990 182.915 55.980 183.055 ;
        RECT 50.110 182.870 50.400 182.915 ;
        RECT 25.875 182.715 26.465 182.760 ;
        RECT 29.115 182.715 29.765 182.760 ;
        RECT 25.875 182.575 29.765 182.715 ;
        RECT 25.875 182.530 26.165 182.575 ;
        RECT 29.115 182.530 29.765 182.575 ;
        RECT 31.755 182.715 32.045 182.760 ;
        RECT 38.195 182.715 38.485 182.760 ;
        RECT 45.080 182.715 45.400 182.775 ;
        RECT 31.755 182.575 32.890 182.715 ;
        RECT 31.755 182.530 32.045 182.575 ;
        RECT 32.750 182.435 32.890 182.575 ;
        RECT 38.195 182.575 45.400 182.715 ;
        RECT 38.195 182.530 38.485 182.575 ;
        RECT 45.080 182.515 45.400 182.575 ;
        RECT 45.540 182.715 45.860 182.775 ;
        RECT 52.430 182.760 52.645 182.915 ;
        RECT 55.215 182.870 55.505 182.915 ;
        RECT 55.660 182.855 55.980 182.915 ;
        RECT 60.275 182.870 60.565 183.100 ;
        RECT 60.810 183.055 60.950 183.195 ;
        RECT 63.020 183.055 63.340 183.115 ;
        RECT 68.095 183.055 68.385 183.100 ;
        RECT 60.810 182.915 62.790 183.055 ;
        RECT 48.250 182.715 48.540 182.760 ;
        RECT 51.510 182.715 51.800 182.760 ;
        RECT 45.540 182.575 51.800 182.715 ;
        RECT 45.540 182.515 45.860 182.575 ;
        RECT 48.250 182.530 48.540 182.575 ;
        RECT 51.510 182.530 51.800 182.575 ;
        RECT 52.430 182.715 52.720 182.760 ;
        RECT 54.290 182.715 54.580 182.760 ;
        RECT 52.430 182.575 54.580 182.715 ;
        RECT 52.430 182.530 52.720 182.575 ;
        RECT 54.290 182.530 54.580 182.575 ;
        RECT 24.380 182.175 24.700 182.435 ;
        RECT 32.660 182.175 32.980 182.435 ;
        RECT 36.800 182.375 37.120 182.435 ;
        RECT 38.655 182.375 38.945 182.420 ;
        RECT 36.800 182.235 38.945 182.375 ;
        RECT 36.800 182.175 37.120 182.235 ;
        RECT 38.655 182.190 38.945 182.235 ;
        RECT 39.560 182.375 39.880 182.435 ;
        RECT 41.415 182.375 41.705 182.420 ;
        RECT 39.560 182.235 41.705 182.375 ;
        RECT 39.560 182.175 39.880 182.235 ;
        RECT 41.415 182.190 41.705 182.235 ;
        RECT 46.245 182.375 46.535 182.420 ;
        RECT 48.760 182.375 49.080 182.435 ;
        RECT 46.245 182.235 49.080 182.375 ;
        RECT 60.350 182.375 60.490 182.870 ;
        RECT 61.640 182.515 61.960 182.775 ;
        RECT 62.650 182.760 62.790 182.915 ;
        RECT 63.020 182.915 68.385 183.055 ;
        RECT 63.020 182.855 63.340 182.915 ;
        RECT 68.095 182.870 68.385 182.915 ;
        RECT 73.140 182.855 73.460 183.115 ;
        RECT 84.640 182.855 84.960 183.115 ;
        RECT 88.320 182.855 88.640 183.115 ;
        RECT 88.780 183.055 89.100 183.115 ;
        RECT 88.780 182.915 89.470 183.055 ;
        RECT 88.780 182.855 89.100 182.915 ;
        RECT 62.575 182.530 62.865 182.760 ;
        RECT 64.875 182.715 65.165 182.760 ;
        RECT 65.320 182.715 65.640 182.775 ;
        RECT 64.875 182.575 65.640 182.715 ;
        RECT 64.875 182.530 65.165 182.575 ;
        RECT 61.180 182.375 61.500 182.435 ;
        RECT 64.950 182.375 65.090 182.530 ;
        RECT 65.320 182.515 65.640 182.575 ;
        RECT 67.175 182.715 67.465 182.760 ;
        RECT 67.620 182.715 67.940 182.775 ;
        RECT 67.175 182.575 67.940 182.715 ;
        RECT 89.330 182.715 89.470 182.915 ;
        RECT 89.700 182.855 90.020 183.115 ;
        RECT 90.250 183.100 90.390 183.595 ;
        RECT 99.475 183.735 99.765 183.780 ;
        RECT 102.595 183.735 102.885 183.780 ;
        RECT 104.485 183.735 104.775 183.780 ;
        RECT 99.475 183.595 104.775 183.735 ;
        RECT 104.970 183.735 105.110 183.935 ;
        RECT 106.260 183.935 107.410 184.075 ;
        RECT 106.260 183.875 106.580 183.935 ;
        RECT 104.970 183.595 106.950 183.735 ;
        RECT 99.475 183.550 99.765 183.595 ;
        RECT 102.595 183.550 102.885 183.595 ;
        RECT 104.485 183.550 104.775 183.595 ;
        RECT 95.220 183.395 95.540 183.455 ;
        RECT 96.155 183.395 96.445 183.440 ;
        RECT 95.220 183.255 96.445 183.395 ;
        RECT 95.220 183.195 95.540 183.255 ;
        RECT 96.155 183.210 96.445 183.255 ;
        RECT 103.960 183.395 104.280 183.455 ;
        RECT 105.355 183.395 105.645 183.440 ;
        RECT 106.260 183.395 106.580 183.455 ;
        RECT 106.810 183.440 106.950 183.595 ;
        RECT 107.270 183.440 107.410 183.935 ;
        RECT 111.795 183.935 113.480 184.075 ;
        RECT 111.795 183.890 112.085 183.935 ;
        RECT 113.160 183.875 113.480 183.935 ;
        RECT 109.495 183.550 109.785 183.780 ;
        RECT 103.960 183.255 106.580 183.395 ;
        RECT 103.960 183.195 104.280 183.255 ;
        RECT 105.355 183.210 105.645 183.255 ;
        RECT 106.260 183.195 106.580 183.255 ;
        RECT 106.735 183.210 107.025 183.440 ;
        RECT 107.195 183.210 107.485 183.440 ;
        RECT 90.175 182.870 90.465 183.100 ;
        RECT 90.620 183.055 90.940 183.115 ;
        RECT 91.095 183.055 91.385 183.100 ;
        RECT 92.935 183.055 93.225 183.100 ;
        RECT 90.620 182.915 91.385 183.055 ;
        RECT 90.620 182.855 90.940 182.915 ;
        RECT 91.095 182.870 91.385 182.915 ;
        RECT 91.630 182.915 93.225 183.055 ;
        RECT 91.630 182.715 91.770 182.915 ;
        RECT 92.935 182.870 93.225 182.915 ;
        RECT 93.380 183.055 93.700 183.115 ;
        RECT 93.855 183.055 94.145 183.100 ;
        RECT 93.380 182.915 94.145 183.055 ;
        RECT 93.380 182.855 93.700 182.915 ;
        RECT 93.855 182.870 94.145 182.915 ;
        RECT 94.300 182.855 94.620 183.115 ;
        RECT 94.775 183.055 95.065 183.100 ;
        RECT 97.520 183.055 97.840 183.115 ;
        RECT 98.440 183.075 98.760 183.115 ;
        RECT 94.775 182.915 97.840 183.055 ;
        RECT 94.775 182.870 95.065 182.915 ;
        RECT 97.520 182.855 97.840 182.915 ;
        RECT 98.395 182.855 98.760 183.075 ;
        RECT 99.475 183.055 99.765 183.100 ;
        RECT 103.055 183.055 103.345 183.100 ;
        RECT 104.890 183.055 105.180 183.100 ;
        RECT 99.475 182.915 105.180 183.055 ;
        RECT 106.810 183.055 106.950 183.210 ;
        RECT 107.640 183.195 107.960 183.455 ;
        RECT 107.730 183.055 107.870 183.195 ;
        RECT 106.810 182.915 107.870 183.055 ;
        RECT 109.570 183.055 109.710 183.550 ;
        RECT 110.875 183.055 111.165 183.100 ;
        RECT 109.570 182.915 111.165 183.055 ;
        RECT 99.475 182.870 99.765 182.915 ;
        RECT 103.055 182.870 103.345 182.915 ;
        RECT 104.890 182.870 105.180 182.915 ;
        RECT 110.875 182.870 111.165 182.915 ;
        RECT 98.395 182.760 98.685 182.855 ;
        RECT 89.330 182.575 91.770 182.715 ;
        RECT 98.095 182.715 98.685 182.760 ;
        RECT 101.335 182.715 101.985 182.760 ;
        RECT 98.095 182.575 101.985 182.715 ;
        RECT 67.175 182.530 67.465 182.575 ;
        RECT 67.620 182.515 67.940 182.575 ;
        RECT 98.095 182.530 98.385 182.575 ;
        RECT 101.335 182.530 101.985 182.575 ;
        RECT 103.975 182.715 104.265 182.760 ;
        RECT 105.800 182.715 106.120 182.775 ;
        RECT 103.975 182.575 106.120 182.715 ;
        RECT 103.975 182.530 104.265 182.575 ;
        RECT 105.800 182.515 106.120 182.575 ;
        RECT 60.350 182.235 65.090 182.375 ;
        RECT 73.615 182.375 73.905 182.420 ;
        RECT 74.060 182.375 74.380 182.435 ;
        RECT 73.615 182.235 74.380 182.375 ;
        RECT 46.245 182.190 46.535 182.235 ;
        RECT 48.760 182.175 49.080 182.235 ;
        RECT 61.180 182.175 61.500 182.235 ;
        RECT 73.615 182.190 73.905 182.235 ;
        RECT 74.060 182.175 74.380 182.235 ;
        RECT 92.015 182.375 92.305 182.420 ;
        RECT 93.380 182.375 93.700 182.435 ;
        RECT 92.015 182.235 93.700 182.375 ;
        RECT 92.015 182.190 92.305 182.235 ;
        RECT 93.380 182.175 93.700 182.235 ;
        RECT 96.615 182.375 96.905 182.420 ;
        RECT 98.900 182.375 99.220 182.435 ;
        RECT 107.655 182.375 107.945 182.420 ;
        RECT 96.615 182.235 107.945 182.375 ;
        RECT 96.615 182.190 96.905 182.235 ;
        RECT 98.900 182.175 99.220 182.235 ;
        RECT 107.655 182.190 107.945 182.235 ;
        RECT 10.650 181.555 118.610 182.035 ;
        RECT 26.695 181.355 26.985 181.400 ;
        RECT 24.930 181.215 26.985 181.355 ;
        RECT 24.930 181.060 25.070 181.215 ;
        RECT 26.695 181.170 26.985 181.215 ;
        RECT 32.215 181.170 32.505 181.400 ;
        RECT 16.575 181.015 16.865 181.060 ;
        RECT 18.975 181.015 19.265 181.060 ;
        RECT 22.215 181.015 22.865 181.060 ;
        RECT 16.575 180.875 22.865 181.015 ;
        RECT 16.575 180.830 16.865 180.875 ;
        RECT 18.975 180.830 19.565 180.875 ;
        RECT 22.215 180.830 22.865 180.875 ;
        RECT 24.855 180.830 25.145 181.060 ;
        RECT 29.440 181.015 29.760 181.075 ;
        RECT 26.310 180.875 29.760 181.015 ;
        RECT 16.115 180.675 16.405 180.720 ;
        RECT 16.115 180.535 19.090 180.675 ;
        RECT 16.115 180.490 16.405 180.535 ;
        RECT 18.950 180.395 19.090 180.535 ;
        RECT 19.275 180.515 19.565 180.830 ;
        RECT 26.310 180.720 26.450 180.875 ;
        RECT 29.440 180.815 29.760 180.875 ;
        RECT 20.355 180.675 20.645 180.720 ;
        RECT 23.935 180.675 24.225 180.720 ;
        RECT 25.770 180.675 26.060 180.720 ;
        RECT 20.355 180.535 26.060 180.675 ;
        RECT 20.355 180.490 20.645 180.535 ;
        RECT 23.935 180.490 24.225 180.535 ;
        RECT 25.770 180.490 26.060 180.535 ;
        RECT 26.235 180.490 26.525 180.720 ;
        RECT 27.600 180.475 27.920 180.735 ;
        RECT 29.915 180.675 30.205 180.720 ;
        RECT 28.150 180.535 30.205 180.675 ;
        RECT 18.860 180.135 19.180 180.395 ;
        RECT 24.380 180.335 24.700 180.395 ;
        RECT 27.140 180.335 27.460 180.395 ;
        RECT 28.150 180.335 28.290 180.535 ;
        RECT 29.915 180.490 30.205 180.535 ;
        RECT 30.360 180.475 30.680 180.735 ;
        RECT 32.290 180.675 32.430 181.170 ;
        RECT 32.660 181.155 32.980 181.415 ;
        RECT 45.080 181.355 45.400 181.415 ;
        RECT 46.245 181.355 46.535 181.400 ;
        RECT 47.380 181.355 47.700 181.415 ;
        RECT 50.140 181.355 50.460 181.415 ;
        RECT 51.075 181.355 51.365 181.400 ;
        RECT 45.080 181.215 49.450 181.355 ;
        RECT 45.080 181.155 45.400 181.215 ;
        RECT 46.245 181.170 46.535 181.215 ;
        RECT 47.380 181.155 47.700 181.215 ;
        RECT 38.200 181.015 38.490 181.060 ;
        RECT 40.060 181.015 40.350 181.060 ;
        RECT 38.200 180.875 40.350 181.015 ;
        RECT 38.200 180.830 38.490 180.875 ;
        RECT 40.060 180.830 40.350 180.875 ;
        RECT 40.980 181.015 41.270 181.060 ;
        RECT 43.240 181.015 43.560 181.075 ;
        RECT 49.310 181.060 49.450 181.215 ;
        RECT 50.140 181.215 51.365 181.355 ;
        RECT 50.140 181.155 50.460 181.215 ;
        RECT 51.075 181.170 51.365 181.215 ;
        RECT 57.515 181.355 57.805 181.400 ;
        RECT 94.300 181.355 94.620 181.415 ;
        RECT 57.515 181.215 94.620 181.355 ;
        RECT 57.515 181.170 57.805 181.215 ;
        RECT 44.240 181.015 44.530 181.060 ;
        RECT 40.980 180.875 44.530 181.015 ;
        RECT 40.980 180.830 41.270 180.875 ;
        RECT 33.595 180.675 33.885 180.720 ;
        RECT 32.290 180.535 33.885 180.675 ;
        RECT 33.595 180.490 33.885 180.535 ;
        RECT 39.115 180.675 39.405 180.720 ;
        RECT 39.560 180.675 39.880 180.735 ;
        RECT 39.115 180.535 39.880 180.675 ;
        RECT 40.135 180.675 40.350 180.830 ;
        RECT 43.240 180.815 43.560 180.875 ;
        RECT 44.240 180.830 44.530 180.875 ;
        RECT 49.235 180.830 49.525 181.060 ;
        RECT 49.680 181.015 50.000 181.075 ;
        RECT 57.590 181.015 57.730 181.170 ;
        RECT 94.300 181.155 94.620 181.215 ;
        RECT 97.535 181.355 97.825 181.400 ;
        RECT 103.960 181.355 104.280 181.415 ;
        RECT 97.535 181.215 104.280 181.355 ;
        RECT 97.535 181.170 97.825 181.215 ;
        RECT 103.960 181.155 104.280 181.215 ;
        RECT 49.680 180.875 57.730 181.015 ;
        RECT 60.720 181.015 61.040 181.075 ;
        RECT 66.240 181.015 66.560 181.075 ;
        RECT 60.720 180.875 64.630 181.015 ;
        RECT 49.680 180.815 50.000 180.875 ;
        RECT 60.720 180.815 61.040 180.875 ;
        RECT 42.380 180.675 42.670 180.720 ;
        RECT 40.135 180.535 42.670 180.675 ;
        RECT 39.115 180.490 39.405 180.535 ;
        RECT 39.560 180.475 39.880 180.535 ;
        RECT 42.380 180.490 42.670 180.535 ;
        RECT 57.960 180.675 58.280 180.735 ;
        RECT 58.435 180.675 58.725 180.720 ;
        RECT 57.960 180.535 58.725 180.675 ;
        RECT 57.960 180.475 58.280 180.535 ;
        RECT 58.435 180.490 58.725 180.535 ;
        RECT 62.575 180.675 62.865 180.720 ;
        RECT 63.020 180.675 63.340 180.735 ;
        RECT 64.490 180.720 64.630 180.875 ;
        RECT 64.950 180.875 66.560 181.015 ;
        RECT 64.950 180.720 65.090 180.875 ;
        RECT 66.240 180.815 66.560 180.875 ;
        RECT 70.855 181.015 71.145 181.060 ;
        RECT 73.600 181.015 73.920 181.075 ;
        RECT 70.855 180.875 73.920 181.015 ;
        RECT 70.855 180.830 71.145 180.875 ;
        RECT 73.600 180.815 73.920 180.875 ;
        RECT 87.515 181.015 87.805 181.060 ;
        RECT 89.700 181.015 90.020 181.075 ;
        RECT 90.755 181.015 91.405 181.060 ;
        RECT 87.515 180.875 91.405 181.015 ;
        RECT 87.515 180.830 88.105 180.875 ;
        RECT 62.575 180.535 63.340 180.675 ;
        RECT 62.575 180.490 62.865 180.535 ;
        RECT 63.020 180.475 63.340 180.535 ;
        RECT 64.415 180.490 64.705 180.720 ;
        RECT 64.875 180.490 65.165 180.720 ;
        RECT 65.335 180.675 65.625 180.720 ;
        RECT 66.700 180.675 67.020 180.735 ;
        RECT 65.335 180.535 67.020 180.675 ;
        RECT 65.335 180.490 65.625 180.535 ;
        RECT 66.700 180.475 67.020 180.535 ;
        RECT 68.080 180.675 68.400 180.735 ;
        RECT 69.015 180.675 69.305 180.720 ;
        RECT 68.080 180.535 69.305 180.675 ;
        RECT 68.080 180.475 68.400 180.535 ;
        RECT 69.015 180.490 69.305 180.535 ;
        RECT 84.195 180.675 84.485 180.720 ;
        RECT 86.020 180.675 86.340 180.735 ;
        RECT 84.195 180.535 86.340 180.675 ;
        RECT 84.195 180.490 84.485 180.535 ;
        RECT 86.020 180.475 86.340 180.535 ;
        RECT 87.815 180.515 88.105 180.830 ;
        RECT 89.700 180.815 90.020 180.875 ;
        RECT 90.755 180.830 91.405 180.875 ;
        RECT 93.380 180.815 93.700 181.075 ;
        RECT 103.500 181.015 103.820 181.075 ;
        RECT 103.500 180.875 106.030 181.015 ;
        RECT 103.500 180.815 103.820 180.875 ;
        RECT 88.895 180.675 89.185 180.720 ;
        RECT 92.475 180.675 92.765 180.720 ;
        RECT 94.310 180.675 94.600 180.720 ;
        RECT 88.895 180.535 94.600 180.675 ;
        RECT 88.895 180.490 89.185 180.535 ;
        RECT 92.475 180.490 92.765 180.535 ;
        RECT 94.310 180.490 94.600 180.535 ;
        RECT 103.960 180.475 104.280 180.735 ;
        RECT 105.890 180.720 106.030 180.875 ;
        RECT 105.815 180.490 106.105 180.720 ;
        RECT 106.720 180.475 107.040 180.735 ;
        RECT 107.180 180.475 107.500 180.735 ;
        RECT 107.655 180.675 107.945 180.720 ;
        RECT 108.100 180.675 108.420 180.735 ;
        RECT 107.655 180.535 108.420 180.675 ;
        RECT 107.655 180.490 107.945 180.535 ;
        RECT 108.100 180.475 108.420 180.535 ;
        RECT 110.415 180.490 110.705 180.720 ;
        RECT 24.380 180.195 28.290 180.335 ;
        RECT 28.520 180.335 28.840 180.395 ;
        RECT 29.455 180.335 29.745 180.380 ;
        RECT 34.040 180.335 34.360 180.395 ;
        RECT 28.520 180.195 34.360 180.335 ;
        RECT 24.380 180.135 24.700 180.195 ;
        RECT 27.140 180.135 27.460 180.195 ;
        RECT 28.520 180.135 28.840 180.195 ;
        RECT 29.455 180.150 29.745 180.195 ;
        RECT 34.040 180.135 34.360 180.195 ;
        RECT 37.275 180.335 37.565 180.380 ;
        RECT 44.620 180.335 44.940 180.395 ;
        RECT 37.275 180.195 44.940 180.335 ;
        RECT 37.275 180.150 37.565 180.195 ;
        RECT 44.620 180.135 44.940 180.195 ;
        RECT 48.300 180.135 48.620 180.395 ;
        RECT 48.760 180.135 49.080 180.395 ;
        RECT 65.795 180.150 66.085 180.380 ;
        RECT 86.110 180.335 86.250 180.475 ;
        RECT 94.775 180.335 95.065 180.380 ;
        RECT 86.110 180.195 95.065 180.335 ;
        RECT 94.775 180.150 95.065 180.195 ;
        RECT 101.200 180.335 101.520 180.395 ;
        RECT 110.490 180.335 110.630 180.490 ;
        RECT 110.860 180.475 111.180 180.735 ;
        RECT 112.700 180.475 113.020 180.735 ;
        RECT 101.200 180.195 110.630 180.335 ;
        RECT 20.355 179.995 20.645 180.040 ;
        RECT 23.475 179.995 23.765 180.040 ;
        RECT 25.365 179.995 25.655 180.040 ;
        RECT 20.355 179.855 25.655 179.995 ;
        RECT 20.355 179.810 20.645 179.855 ;
        RECT 23.475 179.810 23.765 179.855 ;
        RECT 25.365 179.810 25.655 179.855 ;
        RECT 37.740 179.995 38.030 180.040 ;
        RECT 39.600 179.995 39.890 180.040 ;
        RECT 42.380 179.995 42.670 180.040 ;
        RECT 37.740 179.855 42.670 179.995 ;
        RECT 37.740 179.810 38.030 179.855 ;
        RECT 39.600 179.810 39.890 179.855 ;
        RECT 42.380 179.810 42.670 179.855 ;
        RECT 57.500 179.995 57.820 180.055 ;
        RECT 60.720 179.995 61.040 180.055 ;
        RECT 57.500 179.855 61.040 179.995 ;
        RECT 57.500 179.795 57.820 179.855 ;
        RECT 60.720 179.795 61.040 179.855 ;
        RECT 61.180 179.995 61.500 180.055 ;
        RECT 65.870 179.995 66.010 180.150 ;
        RECT 101.200 180.135 101.520 180.195 ;
        RECT 61.180 179.855 66.010 179.995 ;
        RECT 88.895 179.995 89.185 180.040 ;
        RECT 92.015 179.995 92.305 180.040 ;
        RECT 93.905 179.995 94.195 180.040 ;
        RECT 88.895 179.855 94.195 179.995 ;
        RECT 61.180 179.795 61.500 179.855 ;
        RECT 88.895 179.810 89.185 179.855 ;
        RECT 92.015 179.810 92.305 179.855 ;
        RECT 93.905 179.810 94.195 179.855 ;
        RECT 105.800 179.995 106.120 180.055 ;
        RECT 109.495 179.995 109.785 180.040 ;
        RECT 105.800 179.855 109.785 179.995 ;
        RECT 105.800 179.795 106.120 179.855 ;
        RECT 109.495 179.810 109.785 179.855 ;
        RECT 17.495 179.655 17.785 179.700 ;
        RECT 22.080 179.655 22.400 179.715 ;
        RECT 17.495 179.515 22.400 179.655 ;
        RECT 17.495 179.470 17.785 179.515 ;
        RECT 22.080 179.455 22.400 179.515 ;
        RECT 62.560 179.655 62.880 179.715 ;
        RECT 63.035 179.655 63.325 179.700 ;
        RECT 62.560 179.515 63.325 179.655 ;
        RECT 62.560 179.455 62.880 179.515 ;
        RECT 63.035 179.470 63.325 179.515 ;
        RECT 66.700 179.455 67.020 179.715 ;
        RECT 86.035 179.655 86.325 179.700 ;
        RECT 87.860 179.655 88.180 179.715 ;
        RECT 86.035 179.515 88.180 179.655 ;
        RECT 86.035 179.470 86.325 179.515 ;
        RECT 87.860 179.455 88.180 179.515 ;
        RECT 100.280 179.655 100.600 179.715 ;
        RECT 107.180 179.655 107.500 179.715 ;
        RECT 100.280 179.515 107.500 179.655 ;
        RECT 100.280 179.455 100.600 179.515 ;
        RECT 107.180 179.455 107.500 179.515 ;
        RECT 108.560 179.655 108.880 179.715 ;
        RECT 109.035 179.655 109.325 179.700 ;
        RECT 108.560 179.515 109.325 179.655 ;
        RECT 108.560 179.455 108.880 179.515 ;
        RECT 109.035 179.470 109.325 179.515 ;
        RECT 111.320 179.455 111.640 179.715 ;
        RECT 113.635 179.655 113.925 179.700 ;
        RECT 115.000 179.655 115.320 179.715 ;
        RECT 113.635 179.515 115.320 179.655 ;
        RECT 113.635 179.470 113.925 179.515 ;
        RECT 115.000 179.455 115.320 179.515 ;
        RECT 11.430 178.835 118.610 179.315 ;
        RECT 20.700 178.435 21.020 178.695 ;
        RECT 27.600 178.635 27.920 178.695 ;
        RECT 28.995 178.635 29.285 178.680 ;
        RECT 27.600 178.495 29.285 178.635 ;
        RECT 27.600 178.435 27.920 178.495 ;
        RECT 28.995 178.450 29.285 178.495 ;
        RECT 48.300 178.635 48.620 178.695 ;
        RECT 51.535 178.635 51.825 178.680 ;
        RECT 48.300 178.495 51.825 178.635 ;
        RECT 48.300 178.435 48.620 178.495 ;
        RECT 51.535 178.450 51.825 178.495 ;
        RECT 57.500 178.435 57.820 178.695 ;
        RECT 60.720 178.635 61.040 178.695 ;
        RECT 89.700 178.635 90.020 178.695 ;
        RECT 60.720 178.495 90.020 178.635 ;
        RECT 60.720 178.435 61.040 178.495 ;
        RECT 89.700 178.435 90.020 178.495 ;
        RECT 90.175 178.635 90.465 178.680 ;
        RECT 90.620 178.635 90.940 178.695 ;
        RECT 90.175 178.495 90.940 178.635 ;
        RECT 90.175 178.450 90.465 178.495 ;
        RECT 90.620 178.435 90.940 178.495 ;
        RECT 101.200 178.435 101.520 178.695 ;
        RECT 101.660 178.635 101.980 178.695 ;
        RECT 108.100 178.635 108.420 178.695 ;
        RECT 101.660 178.495 108.420 178.635 ;
        RECT 101.660 178.435 101.980 178.495 ;
        RECT 108.100 178.435 108.420 178.495 ;
        RECT 24.855 178.295 25.145 178.340 ;
        RECT 36.800 178.295 37.120 178.355 ;
        RECT 47.840 178.295 48.160 178.355 ;
        RECT 49.680 178.295 50.000 178.355 ;
        RECT 24.855 178.155 37.120 178.295 ;
        RECT 24.855 178.110 25.145 178.155 ;
        RECT 36.800 178.095 37.120 178.155 ;
        RECT 47.010 178.155 50.000 178.295 ;
        RECT 26.235 177.955 26.525 178.000 ;
        RECT 28.520 177.955 28.840 178.015 ;
        RECT 26.235 177.815 28.840 177.955 ;
        RECT 26.235 177.770 26.525 177.815 ;
        RECT 28.520 177.755 28.840 177.815 ;
        RECT 30.360 177.955 30.680 178.015 ;
        RECT 30.360 177.815 37.030 177.955 ;
        RECT 30.360 177.755 30.680 177.815 ;
        RECT 19.320 177.615 19.640 177.675 ;
        RECT 20.255 177.615 20.545 177.660 ;
        RECT 19.320 177.475 20.545 177.615 ;
        RECT 19.320 177.415 19.640 177.475 ;
        RECT 20.255 177.430 20.545 177.475 ;
        RECT 22.080 177.415 22.400 177.675 ;
        RECT 27.140 177.415 27.460 177.675 ;
        RECT 35.420 177.615 35.740 177.675 ;
        RECT 35.895 177.615 36.185 177.660 ;
        RECT 35.420 177.475 36.185 177.615 ;
        RECT 35.420 177.415 35.740 177.475 ;
        RECT 35.895 177.430 36.185 177.475 ;
        RECT 36.340 177.415 36.660 177.675 ;
        RECT 36.890 177.660 37.030 177.815 ;
        RECT 36.815 177.430 37.105 177.660 ;
        RECT 37.735 177.615 38.025 177.660 ;
        RECT 39.560 177.615 39.880 177.675 ;
        RECT 47.010 177.660 47.150 178.155 ;
        RECT 47.840 178.095 48.160 178.155 ;
        RECT 49.680 178.095 50.000 178.155 ;
        RECT 57.590 177.955 57.730 178.435 ;
        RECT 59.340 178.295 59.660 178.355 ;
        RECT 59.815 178.295 60.105 178.340 ;
        RECT 71.760 178.295 72.080 178.355 ;
        RECT 59.340 178.155 72.080 178.295 ;
        RECT 59.340 178.095 59.660 178.155 ;
        RECT 59.815 178.110 60.105 178.155 ;
        RECT 71.760 178.095 72.080 178.155 ;
        RECT 80.010 178.295 80.300 178.340 ;
        RECT 82.790 178.295 83.080 178.340 ;
        RECT 84.650 178.295 84.940 178.340 ;
        RECT 99.820 178.295 100.140 178.355 ;
        RECT 110.515 178.295 110.805 178.340 ;
        RECT 113.635 178.295 113.925 178.340 ;
        RECT 115.525 178.295 115.815 178.340 ;
        RECT 80.010 178.155 84.940 178.295 ;
        RECT 80.010 178.110 80.300 178.155 ;
        RECT 82.790 178.110 83.080 178.155 ;
        RECT 84.650 178.110 84.940 178.155 ;
        RECT 87.490 178.155 100.140 178.295 ;
        RECT 47.930 177.815 57.730 177.955 ;
        RECT 57.960 177.955 58.280 178.015 ;
        RECT 62.115 177.955 62.405 178.000 ;
        RECT 57.960 177.815 62.405 177.955 ;
        RECT 37.735 177.475 39.880 177.615 ;
        RECT 37.735 177.430 38.025 177.475 ;
        RECT 39.560 177.415 39.880 177.475 ;
        RECT 46.475 177.430 46.765 177.660 ;
        RECT 46.935 177.430 47.225 177.660 ;
        RECT 22.170 176.935 22.310 177.415 ;
        RECT 30.360 177.275 30.680 177.335 ;
        RECT 34.040 177.275 34.360 177.335 ;
        RECT 36.430 177.275 36.570 177.415 ;
        RECT 30.360 177.135 36.570 177.275 ;
        RECT 46.550 177.275 46.690 177.430 ;
        RECT 47.380 177.415 47.700 177.675 ;
        RECT 47.930 177.275 48.070 177.815 ;
        RECT 57.960 177.755 58.280 177.815 ;
        RECT 62.115 177.770 62.405 177.815 ;
        RECT 63.035 177.955 63.325 178.000 ;
        RECT 65.780 177.955 66.100 178.015 ;
        RECT 63.035 177.815 66.100 177.955 ;
        RECT 63.035 177.770 63.325 177.815 ;
        RECT 65.780 177.755 66.100 177.815 ;
        RECT 66.700 177.755 67.020 178.015 ;
        RECT 73.155 177.955 73.445 178.000 ;
        RECT 80.500 177.955 80.820 178.015 ;
        RECT 87.490 178.000 87.630 178.155 ;
        RECT 87.415 177.955 87.705 178.000 ;
        RECT 73.155 177.815 87.705 177.955 ;
        RECT 73.155 177.770 73.445 177.815 ;
        RECT 80.500 177.755 80.820 177.815 ;
        RECT 87.415 177.770 87.705 177.815 ;
        RECT 87.860 177.955 88.180 178.015 ;
        RECT 92.920 177.955 93.240 178.015 ;
        RECT 98.530 178.000 98.670 178.155 ;
        RECT 99.820 178.095 100.140 178.155 ;
        RECT 101.750 178.155 104.190 178.295 ;
        RECT 87.860 177.815 93.240 177.955 ;
        RECT 87.860 177.755 88.180 177.815 ;
        RECT 92.920 177.755 93.240 177.815 ;
        RECT 98.455 177.770 98.745 178.000 ;
        RECT 98.900 177.955 99.220 178.015 ;
        RECT 101.750 177.955 101.890 178.155 ;
        RECT 98.900 177.815 101.890 177.955 ;
        RECT 98.900 177.755 99.220 177.815 ;
        RECT 48.315 177.615 48.605 177.660 ;
        RECT 49.680 177.615 50.000 177.675 ;
        RECT 48.315 177.475 50.000 177.615 ;
        RECT 48.315 177.430 48.605 177.475 ;
        RECT 49.680 177.415 50.000 177.475 ;
        RECT 56.595 177.615 56.885 177.660 ;
        RECT 58.050 177.615 58.190 177.755 ;
        RECT 56.595 177.475 58.190 177.615 ;
        RECT 58.435 177.615 58.725 177.660 ;
        RECT 58.880 177.615 59.200 177.675 ;
        RECT 58.435 177.475 59.200 177.615 ;
        RECT 56.595 177.430 56.885 177.475 ;
        RECT 58.435 177.430 58.725 177.475 ;
        RECT 58.880 177.415 59.200 177.475 ;
        RECT 61.640 177.415 61.960 177.675 ;
        RECT 62.560 177.615 62.880 177.675 ;
        RECT 63.495 177.615 63.785 177.660 ;
        RECT 62.560 177.475 63.785 177.615 ;
        RECT 62.560 177.415 62.880 177.475 ;
        RECT 63.495 177.430 63.785 177.475 ;
        RECT 64.875 177.615 65.165 177.660 ;
        RECT 66.790 177.615 66.930 177.755 ;
        RECT 68.095 177.615 68.385 177.660 ;
        RECT 64.875 177.475 68.385 177.615 ;
        RECT 64.875 177.430 65.165 177.475 ;
        RECT 68.095 177.430 68.385 177.475 ;
        RECT 80.010 177.615 80.300 177.660 ;
        RECT 80.010 177.475 82.545 177.615 ;
        RECT 80.010 177.430 80.300 177.475 ;
        RECT 46.550 177.135 48.070 177.275 ;
        RECT 52.915 177.275 53.205 177.320 ;
        RECT 63.955 177.275 64.245 177.320 ;
        RECT 71.775 177.275 72.065 177.320 ;
        RECT 52.915 177.135 72.065 177.275 ;
        RECT 30.360 177.075 30.680 177.135 ;
        RECT 34.040 177.075 34.360 177.135 ;
        RECT 47.470 176.995 47.610 177.135 ;
        RECT 52.915 177.090 53.205 177.135 ;
        RECT 63.955 177.090 64.245 177.135 ;
        RECT 71.775 177.090 72.065 177.135 ;
        RECT 78.150 177.275 78.440 177.320 ;
        RECT 79.580 177.275 79.900 177.335 ;
        RECT 82.330 177.320 82.545 177.475 ;
        RECT 83.260 177.415 83.580 177.675 ;
        RECT 85.115 177.615 85.405 177.660 ;
        RECT 86.020 177.615 86.340 177.675 ;
        RECT 85.115 177.475 86.340 177.615 ;
        RECT 85.115 177.430 85.405 177.475 ;
        RECT 86.020 177.415 86.340 177.475 ;
        RECT 96.155 177.615 96.445 177.660 ;
        RECT 99.375 177.615 99.665 177.660 ;
        RECT 96.155 177.475 99.665 177.615 ;
        RECT 96.155 177.430 96.445 177.475 ;
        RECT 99.375 177.430 99.665 177.475 ;
        RECT 101.660 177.615 101.980 177.675 ;
        RECT 104.050 177.660 104.190 178.155 ;
        RECT 110.515 178.155 115.815 178.295 ;
        RECT 110.515 178.110 110.805 178.155 ;
        RECT 113.635 178.110 113.925 178.155 ;
        RECT 115.525 178.110 115.815 178.155 ;
        RECT 115.000 177.755 115.320 178.015 ;
        RECT 103.055 177.615 103.345 177.660 ;
        RECT 101.660 177.475 103.345 177.615 ;
        RECT 101.660 177.415 101.980 177.475 ;
        RECT 103.055 177.430 103.345 177.475 ;
        RECT 103.515 177.430 103.805 177.660 ;
        RECT 103.975 177.430 104.265 177.660 ;
        RECT 104.895 177.430 105.185 177.660 ;
        RECT 81.410 177.275 81.700 177.320 ;
        RECT 78.150 177.135 81.700 177.275 ;
        RECT 78.150 177.090 78.440 177.135 ;
        RECT 79.580 177.075 79.900 177.135 ;
        RECT 81.410 177.090 81.700 177.135 ;
        RECT 82.330 177.275 82.620 177.320 ;
        RECT 84.190 177.275 84.480 177.320 ;
        RECT 82.330 177.135 84.480 177.275 ;
        RECT 82.330 177.090 82.620 177.135 ;
        RECT 84.190 177.090 84.480 177.135 ;
        RECT 100.280 177.275 100.600 177.335 ;
        RECT 103.590 177.275 103.730 177.430 ;
        RECT 100.280 177.135 103.730 177.275 ;
        RECT 100.280 177.075 100.600 177.135 ;
        RECT 26.695 176.935 26.985 176.980 ;
        RECT 31.740 176.935 32.060 176.995 ;
        RECT 22.170 176.795 32.060 176.935 ;
        RECT 26.695 176.750 26.985 176.795 ;
        RECT 31.740 176.735 32.060 176.795 ;
        RECT 34.515 176.935 34.805 176.980 ;
        RECT 34.960 176.935 35.280 176.995 ;
        RECT 34.515 176.795 35.280 176.935 ;
        RECT 34.515 176.750 34.805 176.795 ;
        RECT 34.960 176.735 35.280 176.795 ;
        RECT 45.080 176.735 45.400 176.995 ;
        RECT 47.380 176.735 47.700 176.995 ;
        RECT 55.660 176.735 55.980 176.995 ;
        RECT 63.480 176.935 63.800 176.995 ;
        RECT 65.795 176.935 66.085 176.980 ;
        RECT 63.480 176.795 66.085 176.935 ;
        RECT 63.480 176.735 63.800 176.795 ;
        RECT 65.795 176.750 66.085 176.795 ;
        RECT 66.240 176.935 66.560 176.995 ;
        RECT 76.360 176.980 76.680 176.995 ;
        RECT 67.175 176.935 67.465 176.980 ;
        RECT 76.145 176.935 76.680 176.980 ;
        RECT 88.335 176.935 88.625 176.980 ;
        RECT 66.240 176.795 67.465 176.935 ;
        RECT 75.925 176.795 88.625 176.935 ;
        RECT 66.240 176.735 66.560 176.795 ;
        RECT 67.175 176.750 67.465 176.795 ;
        RECT 76.145 176.750 76.680 176.795 ;
        RECT 88.335 176.750 88.625 176.795 ;
        RECT 101.200 176.935 101.520 176.995 ;
        RECT 101.675 176.935 101.965 176.980 ;
        RECT 101.200 176.795 101.965 176.935 ;
        RECT 76.360 176.735 76.680 176.750 ;
        RECT 101.200 176.735 101.520 176.795 ;
        RECT 101.675 176.750 101.965 176.795 ;
        RECT 103.500 176.935 103.820 176.995 ;
        RECT 104.970 176.935 105.110 177.430 ;
        RECT 106.260 177.415 106.580 177.675 ;
        RECT 109.435 177.320 109.725 177.635 ;
        RECT 110.515 177.615 110.805 177.660 ;
        RECT 114.095 177.615 114.385 177.660 ;
        RECT 115.930 177.615 116.220 177.660 ;
        RECT 110.515 177.475 116.220 177.615 ;
        RECT 110.515 177.430 110.805 177.475 ;
        RECT 114.095 177.430 114.385 177.475 ;
        RECT 115.930 177.430 116.220 177.475 ;
        RECT 116.380 177.415 116.700 177.675 ;
        RECT 109.135 177.275 109.725 177.320 ;
        RECT 111.320 177.275 111.640 177.335 ;
        RECT 112.375 177.275 113.025 177.320 ;
        RECT 109.135 177.135 113.025 177.275 ;
        RECT 109.135 177.090 109.425 177.135 ;
        RECT 111.320 177.075 111.640 177.135 ;
        RECT 112.375 177.090 113.025 177.135 ;
        RECT 103.500 176.795 105.110 176.935 ;
        RECT 107.655 176.935 107.945 176.980 ;
        RECT 108.100 176.935 108.420 176.995 ;
        RECT 107.655 176.795 108.420 176.935 ;
        RECT 103.500 176.735 103.820 176.795 ;
        RECT 107.655 176.750 107.945 176.795 ;
        RECT 108.100 176.735 108.420 176.795 ;
        RECT 10.650 176.115 118.610 176.595 ;
        RECT 35.420 175.915 35.740 175.975 ;
        RECT 31.370 175.775 35.740 175.915 ;
        RECT 19.320 175.575 19.640 175.635 ;
        RECT 23.460 175.575 23.780 175.635 ;
        RECT 27.140 175.575 27.460 175.635 ;
        RECT 19.320 175.435 26.910 175.575 ;
        RECT 19.320 175.375 19.640 175.435 ;
        RECT 23.460 175.375 23.780 175.435 ;
        RECT 20.240 175.035 20.560 175.295 ;
        RECT 26.770 175.280 26.910 175.435 ;
        RECT 27.140 175.435 30.130 175.575 ;
        RECT 27.140 175.375 27.460 175.435 ;
        RECT 29.990 175.280 30.130 175.435 ;
        RECT 26.695 175.050 26.985 175.280 ;
        RECT 28.995 175.050 29.285 175.280 ;
        RECT 29.915 175.050 30.205 175.280 ;
        RECT 29.070 174.555 29.210 175.050 ;
        RECT 30.360 175.035 30.680 175.295 ;
        RECT 30.835 175.235 31.125 175.280 ;
        RECT 31.370 175.235 31.510 175.775 ;
        RECT 35.420 175.715 35.740 175.775 ;
        RECT 36.340 175.915 36.660 175.975 ;
        RECT 37.720 175.915 38.040 175.975 ;
        RECT 36.340 175.775 38.040 175.915 ;
        RECT 36.340 175.715 36.660 175.775 ;
        RECT 37.720 175.715 38.040 175.775 ;
        RECT 46.000 175.715 46.320 175.975 ;
        RECT 76.360 175.915 76.680 175.975 ;
        RECT 76.835 175.915 77.125 175.960 ;
        RECT 76.360 175.775 77.125 175.915 ;
        RECT 76.360 175.715 76.680 175.775 ;
        RECT 76.835 175.730 77.125 175.775 ;
        RECT 83.260 175.915 83.580 175.975 ;
        RECT 84.195 175.915 84.485 175.960 ;
        RECT 83.260 175.775 84.485 175.915 ;
        RECT 83.260 175.715 83.580 175.775 ;
        RECT 84.195 175.730 84.485 175.775 ;
        RECT 110.415 175.915 110.705 175.960 ;
        RECT 112.700 175.915 113.020 175.975 ;
        RECT 110.415 175.775 113.020 175.915 ;
        RECT 110.415 175.730 110.705 175.775 ;
        RECT 112.700 175.715 113.020 175.775 ;
        RECT 31.740 175.575 32.060 175.635 ;
        RECT 41.860 175.575 42.180 175.635 ;
        RECT 59.340 175.575 59.660 175.635 ;
        RECT 31.740 175.435 38.870 175.575 ;
        RECT 31.740 175.375 32.060 175.435 ;
        RECT 30.835 175.095 31.510 175.235 ;
        RECT 30.835 175.050 31.125 175.095 ;
        RECT 32.660 175.035 32.980 175.295 ;
        RECT 33.595 175.050 33.885 175.280 ;
        RECT 31.280 174.895 31.600 174.955 ;
        RECT 33.670 174.895 33.810 175.050 ;
        RECT 34.040 175.035 34.360 175.295 ;
        RECT 34.515 175.235 34.805 175.280 ;
        RECT 35.420 175.235 35.740 175.295 ;
        RECT 37.735 175.235 38.025 175.280 ;
        RECT 34.515 175.095 38.025 175.235 ;
        RECT 34.515 175.050 34.805 175.095 ;
        RECT 35.420 175.035 35.740 175.095 ;
        RECT 31.280 174.755 33.810 174.895 ;
        RECT 31.280 174.695 31.600 174.755 ;
        RECT 36.340 174.695 36.660 174.955 ;
        RECT 36.890 174.895 37.030 175.095 ;
        RECT 37.735 175.050 38.025 175.095 ;
        RECT 38.180 175.035 38.500 175.295 ;
        RECT 38.730 175.280 38.870 175.435 ;
        RECT 39.190 175.435 59.660 175.575 ;
        RECT 38.655 175.050 38.945 175.280 ;
        RECT 39.190 174.895 39.330 175.435 ;
        RECT 41.860 175.375 42.180 175.435 ;
        RECT 59.340 175.375 59.660 175.435 ;
        RECT 62.560 175.575 62.880 175.635 ;
        RECT 79.580 175.575 79.900 175.635 ;
        RECT 80.975 175.575 81.265 175.620 ;
        RECT 62.560 175.435 68.770 175.575 ;
        RECT 62.560 175.375 62.880 175.435 ;
        RECT 39.560 175.035 39.880 175.295 ;
        RECT 42.335 175.050 42.625 175.280 ;
        RECT 42.780 175.235 43.100 175.295 ;
        RECT 43.255 175.235 43.545 175.280 ;
        RECT 42.780 175.095 43.545 175.235 ;
        RECT 36.890 174.755 39.330 174.895 ;
        RECT 32.660 174.555 32.980 174.615 ;
        RECT 39.560 174.555 39.880 174.615 ;
        RECT 29.070 174.415 39.880 174.555 ;
        RECT 32.660 174.355 32.980 174.415 ;
        RECT 39.560 174.355 39.880 174.415 ;
        RECT 21.160 174.015 21.480 174.275 ;
        RECT 27.140 174.015 27.460 174.275 ;
        RECT 31.740 174.215 32.060 174.275 ;
        RECT 32.215 174.215 32.505 174.260 ;
        RECT 31.740 174.075 32.505 174.215 ;
        RECT 31.740 174.015 32.060 174.075 ;
        RECT 32.215 174.030 32.505 174.075 ;
        RECT 35.895 174.215 36.185 174.260 ;
        RECT 36.340 174.215 36.660 174.275 ;
        RECT 35.895 174.075 36.660 174.215 ;
        RECT 42.410 174.215 42.550 175.050 ;
        RECT 42.780 175.035 43.100 175.095 ;
        RECT 43.255 175.050 43.545 175.095 ;
        RECT 43.715 175.050 44.005 175.280 ;
        RECT 44.175 175.235 44.465 175.280 ;
        RECT 47.380 175.235 47.700 175.295 ;
        RECT 44.175 175.095 47.700 175.235 ;
        RECT 44.175 175.050 44.465 175.095 ;
        RECT 43.790 174.555 43.930 175.050 ;
        RECT 47.380 175.035 47.700 175.095 ;
        RECT 47.840 175.035 48.160 175.295 ;
        RECT 48.315 175.235 48.605 175.280 ;
        RECT 48.760 175.235 49.080 175.295 ;
        RECT 48.315 175.095 49.080 175.235 ;
        RECT 48.315 175.050 48.605 175.095 ;
        RECT 48.760 175.035 49.080 175.095 ;
        RECT 49.235 175.235 49.525 175.280 ;
        RECT 52.900 175.235 53.220 175.295 ;
        RECT 49.235 175.095 53.220 175.235 ;
        RECT 49.235 175.050 49.525 175.095 ;
        RECT 45.555 174.895 45.845 174.940 ;
        RECT 46.920 174.895 47.240 174.955 ;
        RECT 45.555 174.755 47.240 174.895 ;
        RECT 45.555 174.710 45.845 174.755 ;
        RECT 46.920 174.695 47.240 174.755 ;
        RECT 46.000 174.555 46.320 174.615 ;
        RECT 47.930 174.555 48.070 175.035 ;
        RECT 43.790 174.415 48.070 174.555 ;
        RECT 46.000 174.355 46.320 174.415 ;
        RECT 49.310 174.215 49.450 175.050 ;
        RECT 52.900 175.035 53.220 175.095 ;
        RECT 58.435 175.235 58.725 175.280 ;
        RECT 59.800 175.235 60.120 175.295 ;
        RECT 58.435 175.095 60.120 175.235 ;
        RECT 58.435 175.050 58.725 175.095 ;
        RECT 59.800 175.035 60.120 175.095 ;
        RECT 61.640 175.235 61.960 175.295 ;
        RECT 64.030 175.280 64.170 175.435 ;
        RECT 62.115 175.235 62.405 175.280 ;
        RECT 61.640 175.095 62.405 175.235 ;
        RECT 61.640 175.035 61.960 175.095 ;
        RECT 62.115 175.050 62.405 175.095 ;
        RECT 63.955 175.050 64.245 175.280 ;
        RECT 64.415 175.050 64.705 175.280 ;
        RECT 64.490 174.895 64.630 175.050 ;
        RECT 65.780 175.035 66.100 175.295 ;
        RECT 66.700 175.235 67.020 175.295 ;
        RECT 67.175 175.235 67.465 175.280 ;
        RECT 66.700 175.095 67.465 175.235 ;
        RECT 66.700 175.035 67.020 175.095 ;
        RECT 67.175 175.050 67.465 175.095 ;
        RECT 68.630 174.940 68.770 175.435 ;
        RECT 79.580 175.435 81.265 175.575 ;
        RECT 79.580 175.375 79.900 175.435 ;
        RECT 80.975 175.390 81.265 175.435 ;
        RECT 91.490 175.575 91.780 175.620 ;
        RECT 92.920 175.575 93.240 175.635 ;
        RECT 94.750 175.575 95.040 175.620 ;
        RECT 91.490 175.435 95.040 175.575 ;
        RECT 91.490 175.390 91.780 175.435 ;
        RECT 92.920 175.375 93.240 175.435 ;
        RECT 94.750 175.390 95.040 175.435 ;
        RECT 95.670 175.575 95.960 175.620 ;
        RECT 97.530 175.575 97.820 175.620 ;
        RECT 106.260 175.575 106.580 175.635 ;
        RECT 116.380 175.575 116.700 175.635 ;
        RECT 95.670 175.435 97.820 175.575 ;
        RECT 95.670 175.390 95.960 175.435 ;
        RECT 97.530 175.390 97.820 175.435 ;
        RECT 98.070 175.435 116.700 175.575 ;
        RECT 70.395 175.235 70.685 175.280 ;
        RECT 70.285 175.095 70.685 175.235 ;
        RECT 70.395 175.050 70.685 175.095 ;
        RECT 76.820 175.235 77.140 175.295 ;
        RECT 77.295 175.235 77.585 175.280 ;
        RECT 80.500 175.235 80.820 175.295 ;
        RECT 76.820 175.095 77.585 175.235 ;
        RECT 59.430 174.755 64.630 174.895 ;
        RECT 68.555 174.895 68.845 174.940 ;
        RECT 70.470 174.895 70.610 175.050 ;
        RECT 76.820 175.035 77.140 175.095 ;
        RECT 77.295 175.050 77.585 175.095 ;
        RECT 78.750 175.095 80.820 175.235 ;
        RECT 70.840 174.895 71.160 174.955 ;
        RECT 68.555 174.755 71.160 174.895 ;
        RECT 59.430 174.600 59.570 174.755 ;
        RECT 68.555 174.710 68.845 174.755 ;
        RECT 70.840 174.695 71.160 174.755 ;
        RECT 75.440 174.895 75.760 174.955 ;
        RECT 76.375 174.895 76.665 174.940 ;
        RECT 78.750 174.895 78.890 175.095 ;
        RECT 80.500 175.035 80.820 175.095 ;
        RECT 81.420 175.035 81.740 175.295 ;
        RECT 81.880 175.035 82.200 175.295 ;
        RECT 83.275 175.050 83.565 175.280 ;
        RECT 93.350 175.235 93.640 175.280 ;
        RECT 95.670 175.235 95.885 175.390 ;
        RECT 93.350 175.095 95.885 175.235 ;
        RECT 98.070 175.225 98.210 175.435 ;
        RECT 106.260 175.375 106.580 175.435 ;
        RECT 116.380 175.375 116.700 175.435 ;
        RECT 98.455 175.225 98.745 175.280 ;
        RECT 93.350 175.050 93.640 175.095 ;
        RECT 98.070 175.085 98.745 175.225 ;
        RECT 98.455 175.050 98.745 175.085 ;
        RECT 98.900 175.235 99.220 175.295 ;
        RECT 101.660 175.235 101.980 175.295 ;
        RECT 98.900 175.095 101.980 175.235 ;
        RECT 83.350 174.895 83.490 175.050 ;
        RECT 98.900 175.035 99.220 175.095 ;
        RECT 101.660 175.035 101.980 175.095 ;
        RECT 102.135 175.050 102.425 175.280 ;
        RECT 75.440 174.755 78.890 174.895 ;
        RECT 79.210 174.755 83.490 174.895 ;
        RECT 96.615 174.895 96.905 174.940 ;
        RECT 97.060 174.895 97.380 174.955 ;
        RECT 100.280 174.895 100.600 174.955 ;
        RECT 102.210 174.895 102.350 175.050 ;
        RECT 102.580 175.035 102.900 175.295 ;
        RECT 103.500 175.035 103.820 175.295 ;
        RECT 108.575 175.235 108.865 175.280 ;
        RECT 104.050 175.095 108.865 175.235 ;
        RECT 96.615 174.755 97.380 174.895 ;
        RECT 75.440 174.695 75.760 174.755 ;
        RECT 76.375 174.710 76.665 174.755 ;
        RECT 59.355 174.370 59.645 174.600 ;
        RECT 60.720 174.355 61.040 174.615 ;
        RECT 79.210 174.600 79.350 174.755 ;
        RECT 96.615 174.710 96.905 174.755 ;
        RECT 97.060 174.695 97.380 174.755 ;
        RECT 98.990 174.755 102.350 174.895 ;
        RECT 102.670 174.895 102.810 175.035 ;
        RECT 104.050 174.895 104.190 175.095 ;
        RECT 108.575 175.050 108.865 175.095 ;
        RECT 102.670 174.755 104.190 174.895 ;
        RECT 63.110 174.415 78.890 174.555 ;
        RECT 42.410 174.075 49.450 174.215 ;
        RECT 58.880 174.215 59.200 174.275 ;
        RECT 61.195 174.215 61.485 174.260 ;
        RECT 58.880 174.075 61.485 174.215 ;
        RECT 35.895 174.030 36.185 174.075 ;
        RECT 36.340 174.015 36.660 174.075 ;
        RECT 58.880 174.015 59.200 174.075 ;
        RECT 61.195 174.030 61.485 174.075 ;
        RECT 62.560 174.215 62.880 174.275 ;
        RECT 63.110 174.260 63.250 174.415 ;
        RECT 63.035 174.215 63.325 174.260 ;
        RECT 62.560 174.075 63.325 174.215 ;
        RECT 62.560 174.015 62.880 174.075 ;
        RECT 63.035 174.030 63.325 174.075 ;
        RECT 68.080 174.015 68.400 174.275 ;
        RECT 69.460 174.015 69.780 174.275 ;
        RECT 78.750 174.215 78.890 174.415 ;
        RECT 79.135 174.370 79.425 174.600 ;
        RECT 88.780 174.555 89.100 174.615 ;
        RECT 92.000 174.555 92.320 174.615 ;
        RECT 82.430 174.415 92.320 174.555 ;
        RECT 82.430 174.215 82.570 174.415 ;
        RECT 88.780 174.355 89.100 174.415 ;
        RECT 92.000 174.355 92.320 174.415 ;
        RECT 93.350 174.555 93.640 174.600 ;
        RECT 96.130 174.555 96.420 174.600 ;
        RECT 97.990 174.555 98.280 174.600 ;
        RECT 93.350 174.415 98.280 174.555 ;
        RECT 93.350 174.370 93.640 174.415 ;
        RECT 96.130 174.370 96.420 174.415 ;
        RECT 97.990 174.370 98.280 174.415 ;
        RECT 98.990 174.275 99.130 174.755 ;
        RECT 100.280 174.695 100.600 174.755 ;
        RECT 107.180 174.695 107.500 174.955 ;
        RECT 108.100 174.695 108.420 174.955 ;
        RECT 99.820 174.555 100.140 174.615 ;
        RECT 107.270 174.555 107.410 174.695 ;
        RECT 99.820 174.415 107.410 174.555 ;
        RECT 135.635 174.550 136.775 223.880 ;
        RECT 138.130 223.810 139.580 225.110 ;
        RECT 143.180 223.840 144.630 225.140 ;
        RECT 99.820 174.355 100.140 174.415 ;
        RECT 78.750 174.075 82.570 174.215 ;
        RECT 82.815 174.215 83.105 174.260 ;
        RECT 84.180 174.215 84.500 174.275 ;
        RECT 82.815 174.075 84.500 174.215 ;
        RECT 82.815 174.030 83.105 174.075 ;
        RECT 84.180 174.015 84.500 174.075 ;
        RECT 89.240 174.260 89.560 174.275 ;
        RECT 89.240 174.030 89.775 174.260 ;
        RECT 90.620 174.215 90.940 174.275 ;
        RECT 94.300 174.215 94.620 174.275 ;
        RECT 98.900 174.215 99.220 174.275 ;
        RECT 90.620 174.075 99.220 174.215 ;
        RECT 89.240 174.015 89.560 174.030 ;
        RECT 90.620 174.015 90.940 174.075 ;
        RECT 94.300 174.015 94.620 174.075 ;
        RECT 98.900 174.015 99.220 174.075 ;
        RECT 100.295 174.215 100.585 174.260 ;
        RECT 100.740 174.215 101.060 174.275 ;
        RECT 100.295 174.075 101.060 174.215 ;
        RECT 100.295 174.030 100.585 174.075 ;
        RECT 100.740 174.015 101.060 174.075 ;
        RECT 11.430 173.395 118.610 173.875 ;
        RECT 135.580 173.430 136.830 174.550 ;
        RECT 135.635 173.420 136.775 173.430 ;
        RECT 29.440 173.195 29.760 173.255 ;
        RECT 55.660 173.195 55.980 173.255 ;
        RECT 27.690 173.055 34.270 173.195 ;
        RECT 18.515 172.855 18.805 172.900 ;
        RECT 21.635 172.855 21.925 172.900 ;
        RECT 23.525 172.855 23.815 172.900 ;
        RECT 18.515 172.715 23.815 172.855 ;
        RECT 18.515 172.670 18.805 172.715 ;
        RECT 21.635 172.670 21.925 172.715 ;
        RECT 23.525 172.670 23.815 172.715 ;
        RECT 19.320 172.515 19.640 172.575 ;
        RECT 14.810 172.375 19.640 172.515 ;
        RECT 14.810 172.235 14.950 172.375 ;
        RECT 19.320 172.315 19.640 172.375 ;
        RECT 21.160 172.515 21.480 172.575 ;
        RECT 23.015 172.515 23.305 172.560 ;
        RECT 21.160 172.375 23.305 172.515 ;
        RECT 21.160 172.315 21.480 172.375 ;
        RECT 23.015 172.330 23.305 172.375 ;
        RECT 24.395 172.515 24.685 172.560 ;
        RECT 25.760 172.515 26.080 172.575 ;
        RECT 27.690 172.515 27.830 173.055 ;
        RECT 29.440 172.995 29.760 173.055 ;
        RECT 28.175 172.855 28.465 172.900 ;
        RECT 31.295 172.855 31.585 172.900 ;
        RECT 33.185 172.855 33.475 172.900 ;
        RECT 28.175 172.715 33.475 172.855 ;
        RECT 28.175 172.670 28.465 172.715 ;
        RECT 31.295 172.670 31.585 172.715 ;
        RECT 33.185 172.670 33.475 172.715 ;
        RECT 34.130 172.560 34.270 173.055 ;
        RECT 48.390 173.055 55.980 173.195 ;
        RECT 42.780 172.855 43.100 172.915 ;
        RECT 48.390 172.855 48.530 173.055 ;
        RECT 55.660 172.995 55.980 173.055 ;
        RECT 57.960 173.195 58.280 173.255 ;
        RECT 62.560 173.195 62.880 173.255 ;
        RECT 69.460 173.195 69.780 173.255 ;
        RECT 81.420 173.195 81.740 173.255 ;
        RECT 91.080 173.195 91.400 173.255 ;
        RECT 57.960 173.055 62.880 173.195 ;
        RECT 57.960 172.995 58.280 173.055 ;
        RECT 62.560 172.995 62.880 173.055 ;
        RECT 68.630 173.055 77.050 173.195 ;
        RECT 42.780 172.715 48.530 172.855 ;
        RECT 49.680 172.855 50.000 172.915 ;
        RECT 68.630 172.855 68.770 173.055 ;
        RECT 69.460 172.995 69.780 173.055 ;
        RECT 76.360 172.855 76.680 172.915 ;
        RECT 49.680 172.715 68.770 172.855 ;
        RECT 42.780 172.655 43.100 172.715 ;
        RECT 49.680 172.655 50.000 172.715 ;
        RECT 24.395 172.375 27.830 172.515 ;
        RECT 24.395 172.330 24.685 172.375 ;
        RECT 25.760 172.315 26.080 172.375 ;
        RECT 34.055 172.330 34.345 172.560 ;
        RECT 35.880 172.515 36.200 172.575 ;
        RECT 35.880 172.375 37.950 172.515 ;
        RECT 35.880 172.315 36.200 172.375 ;
        RECT 14.720 171.975 15.040 172.235 ;
        RECT 17.435 171.880 17.725 172.195 ;
        RECT 18.515 172.175 18.805 172.220 ;
        RECT 22.095 172.175 22.385 172.220 ;
        RECT 23.930 172.175 24.220 172.220 ;
        RECT 27.140 172.195 27.460 172.235 ;
        RECT 18.515 172.035 24.220 172.175 ;
        RECT 18.515 171.990 18.805 172.035 ;
        RECT 22.095 171.990 22.385 172.035 ;
        RECT 23.930 171.990 24.220 172.035 ;
        RECT 27.095 171.975 27.460 172.195 ;
        RECT 28.175 172.175 28.465 172.220 ;
        RECT 31.755 172.175 32.045 172.220 ;
        RECT 33.590 172.175 33.880 172.220 ;
        RECT 28.175 172.035 33.880 172.175 ;
        RECT 28.175 171.990 28.465 172.035 ;
        RECT 31.755 171.990 32.045 172.035 ;
        RECT 33.590 171.990 33.880 172.035 ;
        RECT 35.420 172.175 35.740 172.235 ;
        RECT 36.815 172.175 37.105 172.220 ;
        RECT 35.420 172.035 37.105 172.175 ;
        RECT 35.420 171.975 35.740 172.035 ;
        RECT 36.815 171.990 37.105 172.035 ;
        RECT 37.260 171.975 37.580 172.235 ;
        RECT 37.810 172.220 37.950 172.375 ;
        RECT 45.630 172.375 47.150 172.515 ;
        RECT 37.735 171.990 38.025 172.220 ;
        RECT 38.655 172.175 38.945 172.220 ;
        RECT 39.560 172.175 39.880 172.235 ;
        RECT 38.655 172.035 39.880 172.175 ;
        RECT 38.655 171.990 38.945 172.035 ;
        RECT 39.560 171.975 39.880 172.035 ;
        RECT 44.160 171.975 44.480 172.235 ;
        RECT 45.630 172.220 45.770 172.375 ;
        RECT 45.555 171.990 45.845 172.220 ;
        RECT 46.000 171.975 46.320 172.235 ;
        RECT 46.475 171.990 46.765 172.220 ;
        RECT 27.095 171.880 27.385 171.975 ;
        RECT 14.275 171.835 14.565 171.880 ;
        RECT 17.135 171.835 17.725 171.880 ;
        RECT 20.375 171.835 21.025 171.880 ;
        RECT 14.275 171.695 21.025 171.835 ;
        RECT 14.275 171.650 14.565 171.695 ;
        RECT 17.135 171.650 17.425 171.695 ;
        RECT 20.375 171.650 21.025 171.695 ;
        RECT 26.795 171.835 27.385 171.880 ;
        RECT 30.035 171.835 30.685 171.880 ;
        RECT 26.795 171.695 30.685 171.835 ;
        RECT 26.795 171.650 27.085 171.695 ;
        RECT 30.035 171.650 30.685 171.695 ;
        RECT 32.675 171.835 32.965 171.880 ;
        RECT 34.040 171.835 34.360 171.895 ;
        RECT 32.675 171.695 34.360 171.835 ;
        RECT 37.350 171.835 37.490 171.975 ;
        RECT 42.780 171.835 43.100 171.895 ;
        RECT 37.350 171.695 43.100 171.835 ;
        RECT 44.250 171.835 44.390 171.975 ;
        RECT 46.550 171.835 46.690 171.990 ;
        RECT 44.250 171.695 46.690 171.835 ;
        RECT 32.675 171.650 32.965 171.695 ;
        RECT 34.040 171.635 34.360 171.695 ;
        RECT 42.780 171.635 43.100 171.695 ;
        RECT 15.655 171.495 15.945 171.540 ;
        RECT 17.940 171.495 18.260 171.555 ;
        RECT 15.655 171.355 18.260 171.495 ;
        RECT 15.655 171.310 15.945 171.355 ;
        RECT 17.940 171.295 18.260 171.355 ;
        RECT 25.315 171.495 25.605 171.540 ;
        RECT 26.220 171.495 26.540 171.555 ;
        RECT 25.315 171.355 26.540 171.495 ;
        RECT 25.315 171.310 25.605 171.355 ;
        RECT 26.220 171.295 26.540 171.355 ;
        RECT 33.120 171.495 33.440 171.555 ;
        RECT 35.435 171.495 35.725 171.540 ;
        RECT 33.120 171.355 35.725 171.495 ;
        RECT 33.120 171.295 33.440 171.355 ;
        RECT 35.435 171.310 35.725 171.355 ;
        RECT 41.400 171.495 41.720 171.555 ;
        RECT 44.175 171.495 44.465 171.540 ;
        RECT 41.400 171.355 44.465 171.495 ;
        RECT 47.010 171.495 47.150 172.375 ;
        RECT 68.630 172.235 68.770 172.715 ;
        RECT 69.550 172.715 76.680 172.855 ;
        RECT 47.395 171.990 47.685 172.220 ;
        RECT 49.220 172.175 49.540 172.235 ;
        RECT 49.695 172.175 49.985 172.220 ;
        RECT 49.220 172.035 49.985 172.175 ;
        RECT 47.470 171.835 47.610 171.990 ;
        RECT 49.220 171.975 49.540 172.035 ;
        RECT 49.695 171.990 49.985 172.035 ;
        RECT 68.540 171.975 68.860 172.235 ;
        RECT 69.550 172.220 69.690 172.715 ;
        RECT 76.360 172.655 76.680 172.715 ;
        RECT 70.010 172.375 74.290 172.515 ;
        RECT 70.010 172.220 70.150 172.375 ;
        RECT 69.475 171.990 69.765 172.220 ;
        RECT 69.935 171.990 70.225 172.220 ;
        RECT 70.395 172.175 70.685 172.220 ;
        RECT 72.220 172.175 72.540 172.235 ;
        RECT 74.150 172.220 74.290 172.375 ;
        RECT 73.615 172.175 73.905 172.220 ;
        RECT 70.395 172.035 73.905 172.175 ;
        RECT 70.395 171.990 70.685 172.035 ;
        RECT 52.900 171.835 53.220 171.895 ;
        RECT 57.960 171.835 58.280 171.895 ;
        RECT 70.010 171.835 70.150 171.990 ;
        RECT 72.220 171.975 72.540 172.035 ;
        RECT 73.615 171.990 73.905 172.035 ;
        RECT 74.075 171.990 74.365 172.220 ;
        RECT 74.535 171.990 74.825 172.220 ;
        RECT 74.980 172.175 75.300 172.235 ;
        RECT 75.455 172.175 75.745 172.220 ;
        RECT 76.910 172.175 77.050 173.055 ;
        RECT 81.420 173.055 91.400 173.195 ;
        RECT 81.420 172.995 81.740 173.055 ;
        RECT 80.055 172.515 80.345 172.560 ;
        RECT 80.500 172.515 80.820 172.575 ;
        RECT 80.055 172.375 80.820 172.515 ;
        RECT 80.055 172.330 80.345 172.375 ;
        RECT 80.500 172.315 80.820 172.375 ;
        RECT 74.980 172.035 77.050 172.175 ;
        RECT 77.280 172.175 77.600 172.235 ;
        RECT 78.675 172.175 78.965 172.220 ;
        RECT 82.430 172.175 82.570 173.055 ;
        RECT 91.080 172.995 91.400 173.055 ;
        RECT 92.000 173.195 92.320 173.255 ;
        RECT 101.660 173.195 101.980 173.255 ;
        RECT 103.500 173.195 103.820 173.255 ;
        RECT 92.000 173.055 103.820 173.195 ;
        RECT 92.000 172.995 92.320 173.055 ;
        RECT 101.660 172.995 101.980 173.055 ;
        RECT 103.500 172.995 103.820 173.055 ;
        RECT 82.815 172.670 83.105 172.900 ;
        RECT 89.240 172.855 89.560 172.915 ;
        RECT 92.460 172.855 92.780 172.915 ;
        RECT 108.990 172.855 109.280 172.900 ;
        RECT 111.770 172.855 112.060 172.900 ;
        RECT 113.630 172.855 113.920 172.900 ;
        RECT 89.240 172.715 92.780 172.855 ;
        RECT 82.890 172.515 83.030 172.670 ;
        RECT 89.240 172.655 89.560 172.715 ;
        RECT 92.460 172.655 92.780 172.715 ;
        RECT 93.470 172.715 102.350 172.855 ;
        RECT 82.890 172.375 84.410 172.515 ;
        RECT 83.275 172.175 83.565 172.220 ;
        RECT 77.280 172.035 83.565 172.175 ;
        RECT 84.270 172.185 84.410 172.375 ;
        RECT 84.655 172.185 84.945 172.220 ;
        RECT 84.270 172.045 84.945 172.185 ;
        RECT 47.470 171.695 58.280 171.835 ;
        RECT 52.900 171.635 53.220 171.695 ;
        RECT 57.960 171.635 58.280 171.695 ;
        RECT 59.200 171.695 70.150 171.835 ;
        RECT 71.775 171.835 72.065 171.880 ;
        RECT 74.610 171.835 74.750 171.990 ;
        RECT 74.980 171.975 75.300 172.035 ;
        RECT 75.455 171.990 75.745 172.035 ;
        RECT 77.280 171.975 77.600 172.035 ;
        RECT 78.675 171.990 78.965 172.035 ;
        RECT 83.275 171.990 83.565 172.035 ;
        RECT 84.655 171.990 84.945 172.045 ;
        RECT 80.975 171.835 81.265 171.880 ;
        RECT 89.330 171.835 89.470 172.655 ;
        RECT 93.470 172.515 93.610 172.715 ;
        RECT 91.170 172.375 93.610 172.515 ;
        RECT 89.700 172.175 90.020 172.235 ;
        RECT 90.175 172.175 90.465 172.220 ;
        RECT 89.700 172.035 90.465 172.175 ;
        RECT 89.700 171.975 90.020 172.035 ;
        RECT 90.175 171.990 90.465 172.035 ;
        RECT 71.775 171.695 73.830 171.835 ;
        RECT 74.610 171.695 89.470 171.835 ;
        RECT 47.380 171.495 47.700 171.555 ;
        RECT 47.010 171.355 47.700 171.495 ;
        RECT 41.400 171.295 41.720 171.355 ;
        RECT 44.175 171.310 44.465 171.355 ;
        RECT 47.380 171.295 47.700 171.355 ;
        RECT 49.680 171.495 50.000 171.555 ;
        RECT 50.155 171.495 50.445 171.540 ;
        RECT 49.680 171.355 50.445 171.495 ;
        RECT 49.680 171.295 50.000 171.355 ;
        RECT 50.155 171.310 50.445 171.355 ;
        RECT 55.660 171.495 55.980 171.555 ;
        RECT 59.200 171.495 59.340 171.695 ;
        RECT 69.550 171.555 69.690 171.695 ;
        RECT 71.775 171.650 72.065 171.695 ;
        RECT 73.690 171.555 73.830 171.695 ;
        RECT 80.975 171.650 81.265 171.695 ;
        RECT 55.660 171.355 59.340 171.495 ;
        RECT 61.180 171.495 61.500 171.555 ;
        RECT 68.080 171.495 68.400 171.555 ;
        RECT 61.180 171.355 68.400 171.495 ;
        RECT 55.660 171.295 55.980 171.355 ;
        RECT 61.180 171.295 61.500 171.355 ;
        RECT 68.080 171.295 68.400 171.355 ;
        RECT 69.460 171.295 69.780 171.555 ;
        RECT 72.220 171.295 72.540 171.555 ;
        RECT 73.600 171.295 73.920 171.555 ;
        RECT 78.215 171.495 78.505 171.540 ;
        RECT 79.580 171.495 79.900 171.555 ;
        RECT 78.215 171.355 79.900 171.495 ;
        RECT 78.215 171.310 78.505 171.355 ;
        RECT 79.580 171.295 79.900 171.355 ;
        RECT 80.500 171.295 80.820 171.555 ;
        RECT 83.720 171.295 84.040 171.555 ;
        RECT 85.575 171.495 85.865 171.540 ;
        RECT 87.400 171.495 87.720 171.555 ;
        RECT 85.575 171.355 87.720 171.495 ;
        RECT 85.575 171.310 85.865 171.355 ;
        RECT 87.400 171.295 87.720 171.355 ;
        RECT 88.795 171.495 89.085 171.540 ;
        RECT 89.700 171.495 90.020 171.555 ;
        RECT 88.795 171.355 90.020 171.495 ;
        RECT 90.250 171.495 90.390 171.990 ;
        RECT 90.620 171.975 90.940 172.235 ;
        RECT 91.170 172.220 91.310 172.375 ;
        RECT 91.095 171.990 91.385 172.220 ;
        RECT 92.000 171.975 92.320 172.235 ;
        RECT 93.470 172.175 93.610 172.375 ;
        RECT 93.855 172.515 94.145 172.560 ;
        RECT 99.820 172.515 100.140 172.575 ;
        RECT 102.210 172.560 102.350 172.715 ;
        RECT 108.990 172.715 113.920 172.855 ;
        RECT 108.990 172.670 109.280 172.715 ;
        RECT 111.770 172.670 112.060 172.715 ;
        RECT 113.630 172.670 113.920 172.715 ;
        RECT 101.215 172.515 101.505 172.560 ;
        RECT 93.855 172.375 101.505 172.515 ;
        RECT 93.855 172.330 94.145 172.375 ;
        RECT 99.820 172.315 100.140 172.375 ;
        RECT 101.215 172.330 101.505 172.375 ;
        RECT 102.135 172.515 102.425 172.560 ;
        RECT 105.125 172.515 105.415 172.560 ;
        RECT 102.135 172.375 105.415 172.515 ;
        RECT 102.135 172.330 102.425 172.375 ;
        RECT 105.125 172.330 105.415 172.375 ;
        RECT 114.095 172.515 114.385 172.560 ;
        RECT 116.380 172.515 116.700 172.575 ;
        RECT 114.095 172.375 116.700 172.515 ;
        RECT 114.095 172.330 114.385 172.375 ;
        RECT 116.380 172.315 116.700 172.375 ;
        RECT 94.775 172.175 95.065 172.220 ;
        RECT 98.440 172.175 98.760 172.235 ;
        RECT 93.470 172.035 95.065 172.175 ;
        RECT 94.775 171.990 95.065 172.035 ;
        RECT 95.770 172.035 98.760 172.175 ;
        RECT 92.460 171.835 92.780 171.895 ;
        RECT 94.315 171.835 94.605 171.880 ;
        RECT 92.460 171.695 94.605 171.835 ;
        RECT 92.460 171.635 92.780 171.695 ;
        RECT 94.315 171.650 94.605 171.695 ;
        RECT 95.770 171.495 95.910 172.035 ;
        RECT 98.440 171.975 98.760 172.035 ;
        RECT 98.900 171.975 99.220 172.235 ;
        RECT 99.375 171.990 99.665 172.220 ;
        RECT 100.295 172.175 100.585 172.220 ;
        RECT 101.660 172.175 101.980 172.235 ;
        RECT 100.295 172.035 101.980 172.175 ;
        RECT 100.295 171.990 100.585 172.035 ;
        RECT 99.450 171.835 99.590 171.990 ;
        RECT 101.660 171.975 101.980 172.035 ;
        RECT 102.595 172.175 102.885 172.220 ;
        RECT 108.100 172.175 108.420 172.235 ;
        RECT 102.595 172.035 108.420 172.175 ;
        RECT 102.595 171.990 102.885 172.035 ;
        RECT 102.670 171.835 102.810 171.990 ;
        RECT 108.100 171.975 108.420 172.035 ;
        RECT 108.990 172.175 109.280 172.220 ;
        RECT 108.990 172.035 111.525 172.175 ;
        RECT 108.990 171.990 109.280 172.035 ;
        RECT 107.180 171.880 107.500 171.895 ;
        RECT 111.310 171.880 111.525 172.035 ;
        RECT 112.240 171.975 112.560 172.235 ;
        RECT 115.460 171.975 115.780 172.235 ;
        RECT 133.700 172.190 134.930 172.680 ;
        RECT 133.700 171.930 136.690 172.190 ;
        RECT 138.330 171.930 139.470 223.810 ;
        RECT 99.450 171.695 102.810 171.835 ;
        RECT 107.130 171.835 107.500 171.880 ;
        RECT 110.390 171.835 110.680 171.880 ;
        RECT 107.130 171.695 110.680 171.835 ;
        RECT 107.130 171.650 107.500 171.695 ;
        RECT 110.390 171.650 110.680 171.695 ;
        RECT 111.310 171.835 111.600 171.880 ;
        RECT 113.170 171.835 113.460 171.880 ;
        RECT 111.310 171.695 113.460 171.835 ;
        RECT 111.310 171.650 111.600 171.695 ;
        RECT 113.170 171.650 113.460 171.695 ;
        RECT 113.620 171.835 113.940 171.895 ;
        RECT 114.555 171.835 114.845 171.880 ;
        RECT 113.620 171.695 114.845 171.835 ;
        RECT 107.180 171.635 107.500 171.650 ;
        RECT 113.620 171.635 113.940 171.695 ;
        RECT 114.555 171.650 114.845 171.695 ;
        RECT 90.250 171.355 95.910 171.495 ;
        RECT 88.795 171.310 89.085 171.355 ;
        RECT 89.700 171.295 90.020 171.355 ;
        RECT 96.600 171.295 96.920 171.555 ;
        RECT 97.075 171.495 97.365 171.540 ;
        RECT 97.520 171.495 97.840 171.555 ;
        RECT 97.075 171.355 97.840 171.495 ;
        RECT 97.075 171.310 97.365 171.355 ;
        RECT 97.520 171.295 97.840 171.355 ;
        RECT 104.435 171.495 104.725 171.540 ;
        RECT 109.020 171.495 109.340 171.555 ;
        RECT 104.435 171.355 109.340 171.495 ;
        RECT 104.435 171.310 104.725 171.355 ;
        RECT 109.020 171.295 109.340 171.355 ;
        RECT 10.650 170.675 118.610 171.155 ;
        RECT 133.700 170.790 139.470 171.930 ;
        RECT 133.700 170.600 136.690 170.790 ;
        RECT 18.415 170.475 18.705 170.520 ;
        RECT 20.240 170.475 20.560 170.535 ;
        RECT 18.415 170.335 20.560 170.475 ;
        RECT 18.415 170.290 18.705 170.335 ;
        RECT 20.240 170.275 20.560 170.335 ;
        RECT 21.175 170.475 21.465 170.520 ;
        RECT 25.760 170.475 26.080 170.535 ;
        RECT 61.180 170.475 61.500 170.535 ;
        RECT 21.175 170.335 26.080 170.475 ;
        RECT 21.175 170.290 21.465 170.335 ;
        RECT 25.760 170.275 26.080 170.335 ;
        RECT 34.590 170.335 53.130 170.475 ;
        RECT 15.640 170.135 15.960 170.195 ;
        RECT 16.575 170.135 16.865 170.180 ;
        RECT 15.640 169.995 16.865 170.135 ;
        RECT 15.640 169.935 15.960 169.995 ;
        RECT 16.575 169.950 16.865 169.995 ;
        RECT 27.600 169.935 27.920 170.195 ;
        RECT 34.590 170.180 34.730 170.335 ;
        RECT 34.515 169.950 34.805 170.180 ;
        RECT 48.295 170.135 48.945 170.180 ;
        RECT 49.680 170.135 50.000 170.195 ;
        RECT 51.895 170.135 52.185 170.180 ;
        RECT 48.295 169.995 52.185 170.135 ;
        RECT 52.990 170.135 53.130 170.335 ;
        RECT 53.910 170.335 61.500 170.475 ;
        RECT 53.910 170.135 54.050 170.335 ;
        RECT 61.180 170.275 61.500 170.335 ;
        RECT 69.460 170.475 69.780 170.535 ;
        RECT 76.820 170.475 77.140 170.535 ;
        RECT 92.920 170.475 93.240 170.535 ;
        RECT 93.395 170.475 93.685 170.520 ;
        RECT 69.460 170.335 73.830 170.475 ;
        RECT 69.460 170.275 69.780 170.335 ;
        RECT 64.415 170.135 64.705 170.180 ;
        RECT 52.990 169.995 54.050 170.135 ;
        RECT 58.510 169.995 64.705 170.135 ;
        RECT 48.295 169.950 48.945 169.995 ;
        RECT 49.680 169.935 50.000 169.995 ;
        RECT 51.595 169.950 52.185 169.995 ;
        RECT 14.275 169.795 14.565 169.840 ;
        RECT 14.720 169.795 15.040 169.855 ;
        RECT 21.160 169.795 21.480 169.855 ;
        RECT 14.275 169.655 15.040 169.795 ;
        RECT 14.275 169.610 14.565 169.655 ;
        RECT 14.720 169.595 15.040 169.655 ;
        RECT 15.730 169.655 21.480 169.795 ;
        RECT 15.730 169.500 15.870 169.655 ;
        RECT 21.160 169.595 21.480 169.655 ;
        RECT 29.440 169.595 29.760 169.855 ;
        RECT 30.375 169.795 30.665 169.840 ;
        RECT 36.355 169.795 36.645 169.840 ;
        RECT 30.375 169.655 36.645 169.795 ;
        RECT 30.375 169.610 30.665 169.655 ;
        RECT 36.355 169.610 36.645 169.655 ;
        RECT 37.735 169.610 38.025 169.840 ;
        RECT 41.860 169.795 42.180 169.855 ;
        RECT 42.335 169.795 42.625 169.840 ;
        RECT 41.860 169.655 42.625 169.795 ;
        RECT 15.655 169.270 15.945 169.500 ;
        RECT 16.115 169.455 16.405 169.500 ;
        RECT 17.940 169.455 18.260 169.515 ;
        RECT 21.620 169.455 21.940 169.515 ;
        RECT 16.115 169.315 21.940 169.455 ;
        RECT 16.115 169.270 16.405 169.315 ;
        RECT 17.940 169.255 18.260 169.315 ;
        RECT 21.620 169.255 21.940 169.315 ;
        RECT 23.460 169.455 23.780 169.515 ;
        RECT 30.450 169.455 30.590 169.610 ;
        RECT 23.460 169.315 30.590 169.455 ;
        RECT 37.810 169.455 37.950 169.610 ;
        RECT 41.860 169.595 42.180 169.655 ;
        RECT 42.335 169.610 42.625 169.655 ;
        RECT 42.780 169.595 43.100 169.855 ;
        RECT 43.255 169.795 43.545 169.840 ;
        RECT 43.700 169.795 44.020 169.855 ;
        RECT 43.255 169.655 44.020 169.795 ;
        RECT 43.255 169.610 43.545 169.655 ;
        RECT 43.700 169.595 44.020 169.655 ;
        RECT 44.160 169.595 44.480 169.855 ;
        RECT 45.100 169.795 45.390 169.840 ;
        RECT 46.935 169.795 47.225 169.840 ;
        RECT 50.515 169.795 50.805 169.840 ;
        RECT 45.100 169.655 50.805 169.795 ;
        RECT 45.100 169.610 45.390 169.655 ;
        RECT 46.935 169.610 47.225 169.655 ;
        RECT 50.515 169.610 50.805 169.655 ;
        RECT 51.595 169.635 51.885 169.950 ;
        RECT 37.810 169.315 38.410 169.455 ;
        RECT 23.460 169.255 23.780 169.315 ;
        RECT 13.815 169.115 14.105 169.160 ;
        RECT 16.560 169.115 16.880 169.175 ;
        RECT 13.815 168.975 16.880 169.115 ;
        RECT 13.815 168.930 14.105 168.975 ;
        RECT 16.560 168.915 16.880 168.975 ;
        RECT 30.835 169.115 31.125 169.160 ;
        RECT 32.200 169.115 32.520 169.175 ;
        RECT 30.835 168.975 32.520 169.115 ;
        RECT 30.835 168.930 31.125 168.975 ;
        RECT 32.200 168.915 32.520 168.975 ;
        RECT 32.660 168.775 32.980 168.835 ;
        RECT 33.135 168.775 33.425 168.820 ;
        RECT 32.660 168.635 33.425 168.775 ;
        RECT 38.270 168.775 38.410 169.315 ;
        RECT 44.620 169.255 44.940 169.515 ;
        RECT 46.000 169.255 46.320 169.515 ;
        RECT 49.680 169.455 50.000 169.515 ;
        RECT 53.375 169.455 53.665 169.500 ;
        RECT 49.680 169.315 53.665 169.455 ;
        RECT 49.680 169.255 50.000 169.315 ;
        RECT 53.375 169.270 53.665 169.315 ;
        RECT 40.940 168.915 41.260 169.175 ;
        RECT 39.560 168.775 39.880 168.835 ;
        RECT 38.270 168.635 39.880 168.775 ;
        RECT 44.710 168.775 44.850 169.255 ;
        RECT 45.505 169.115 45.795 169.160 ;
        RECT 47.395 169.115 47.685 169.160 ;
        RECT 50.515 169.115 50.805 169.160 ;
        RECT 45.505 168.975 50.805 169.115 ;
        RECT 45.505 168.930 45.795 168.975 ;
        RECT 47.395 168.930 47.685 168.975 ;
        RECT 50.515 168.930 50.805 168.975 ;
        RECT 51.060 169.115 51.380 169.175 ;
        RECT 58.510 169.115 58.650 169.995 ;
        RECT 64.415 169.950 64.705 169.995 ;
        RECT 59.355 169.610 59.645 169.840 ;
        RECT 60.720 169.795 61.040 169.855 ;
        RECT 63.940 169.795 64.260 169.855 ;
        RECT 60.720 169.655 64.260 169.795 ;
        RECT 59.430 169.455 59.570 169.610 ;
        RECT 60.720 169.595 61.040 169.655 ;
        RECT 63.940 169.595 64.260 169.655 ;
        RECT 64.490 169.455 64.630 169.950 ;
        RECT 65.780 169.795 66.100 169.855 ;
        RECT 67.635 169.795 67.925 169.840 ;
        RECT 65.780 169.655 67.925 169.795 ;
        RECT 65.780 169.595 66.100 169.655 ;
        RECT 67.635 169.610 67.925 169.655 ;
        RECT 68.095 169.795 68.385 169.840 ;
        RECT 68.540 169.795 68.860 169.855 ;
        RECT 68.095 169.655 68.860 169.795 ;
        RECT 68.095 169.610 68.385 169.655 ;
        RECT 68.540 169.595 68.860 169.655 ;
        RECT 69.000 169.595 69.320 169.855 ;
        RECT 69.460 169.595 69.780 169.855 ;
        RECT 69.935 169.795 70.225 169.840 ;
        RECT 71.760 169.795 72.080 169.855 ;
        RECT 73.690 169.840 73.830 170.335 ;
        RECT 74.150 170.335 77.140 170.475 ;
        RECT 74.150 169.840 74.290 170.335 ;
        RECT 76.820 170.275 77.140 170.335 ;
        RECT 77.370 170.335 90.390 170.475 ;
        RECT 77.370 170.135 77.510 170.335 ;
        RECT 74.610 169.995 77.510 170.135 ;
        RECT 82.290 170.135 82.580 170.180 ;
        RECT 83.720 170.135 84.040 170.195 ;
        RECT 85.550 170.135 85.840 170.180 ;
        RECT 82.290 169.995 85.840 170.135 ;
        RECT 73.055 169.795 73.345 169.840 ;
        RECT 69.935 169.745 72.910 169.795 ;
        RECT 73.055 169.745 73.370 169.795 ;
        RECT 69.935 169.655 73.370 169.745 ;
        RECT 69.935 169.610 70.225 169.655 ;
        RECT 71.760 169.595 72.080 169.655 ;
        RECT 72.770 169.605 73.370 169.655 ;
        RECT 73.615 169.610 73.905 169.840 ;
        RECT 74.075 169.610 74.365 169.840 ;
        RECT 74.610 169.455 74.750 169.995 ;
        RECT 82.290 169.950 82.580 169.995 ;
        RECT 83.720 169.935 84.040 169.995 ;
        RECT 85.550 169.950 85.840 169.995 ;
        RECT 86.470 170.135 86.760 170.180 ;
        RECT 88.330 170.135 88.620 170.180 ;
        RECT 86.470 169.995 88.620 170.135 ;
        RECT 86.470 169.950 86.760 169.995 ;
        RECT 88.330 169.950 88.620 169.995 ;
        RECT 74.980 169.595 75.300 169.855 ;
        RECT 80.500 169.840 80.820 169.855 ;
        RECT 77.295 169.795 77.585 169.840 ;
        RECT 80.285 169.795 80.820 169.840 ;
        RECT 76.910 169.655 80.820 169.795 ;
        RECT 59.430 169.315 63.250 169.455 ;
        RECT 64.490 169.315 74.750 169.455 ;
        RECT 75.440 169.455 75.760 169.515 ;
        RECT 75.915 169.455 76.205 169.500 ;
        RECT 75.440 169.315 76.205 169.455 ;
        RECT 63.110 169.175 63.250 169.315 ;
        RECT 75.440 169.255 75.760 169.315 ;
        RECT 75.915 169.270 76.205 169.315 ;
        RECT 51.060 168.975 58.650 169.115 ;
        RECT 51.060 168.915 51.380 168.975 ;
        RECT 58.880 168.915 59.200 169.175 ;
        RECT 63.020 169.115 63.340 169.175 ;
        RECT 65.780 169.115 66.100 169.175 ;
        RECT 63.020 168.975 66.100 169.115 ;
        RECT 63.020 168.915 63.340 168.975 ;
        RECT 65.780 168.915 66.100 168.975 ;
        RECT 67.160 168.915 67.480 169.175 ;
        RECT 71.315 168.930 71.605 169.160 ;
        RECT 53.820 168.775 54.140 168.835 ;
        RECT 44.710 168.635 54.140 168.775 ;
        RECT 32.660 168.575 32.980 168.635 ;
        RECT 33.135 168.590 33.425 168.635 ;
        RECT 39.560 168.575 39.880 168.635 ;
        RECT 53.820 168.575 54.140 168.635 ;
        RECT 55.200 168.775 55.520 168.835 ;
        RECT 61.655 168.775 61.945 168.820 ;
        RECT 64.400 168.775 64.720 168.835 ;
        RECT 55.200 168.635 64.720 168.775 ;
        RECT 71.390 168.775 71.530 168.930 ;
        RECT 71.760 168.915 72.080 169.175 ;
        RECT 72.680 169.115 73.000 169.175 ;
        RECT 76.910 169.115 77.050 169.655 ;
        RECT 77.295 169.610 77.585 169.655 ;
        RECT 80.285 169.610 80.820 169.655 ;
        RECT 84.150 169.795 84.440 169.840 ;
        RECT 86.470 169.795 86.685 169.950 ;
        RECT 84.150 169.655 86.685 169.795 ;
        RECT 84.150 169.610 84.440 169.655 ;
        RECT 80.500 169.595 80.820 169.610 ;
        RECT 87.400 169.595 87.720 169.855 ;
        RECT 86.020 169.455 86.340 169.515 ;
        RECT 89.255 169.455 89.545 169.500 ;
        RECT 86.020 169.315 89.545 169.455 ;
        RECT 90.250 169.455 90.390 170.335 ;
        RECT 92.920 170.335 93.685 170.475 ;
        RECT 92.920 170.275 93.240 170.335 ;
        RECT 93.395 170.290 93.685 170.335 ;
        RECT 97.060 170.275 97.380 170.535 ;
        RECT 106.735 170.475 107.025 170.520 ;
        RECT 107.180 170.475 107.500 170.535 ;
        RECT 106.735 170.335 107.500 170.475 ;
        RECT 106.735 170.290 107.025 170.335 ;
        RECT 107.180 170.275 107.500 170.335 ;
        RECT 111.335 170.475 111.625 170.520 ;
        RECT 112.240 170.475 112.560 170.535 ;
        RECT 111.335 170.335 112.560 170.475 ;
        RECT 111.335 170.290 111.625 170.335 ;
        RECT 112.240 170.275 112.560 170.335 ;
        RECT 90.620 170.135 90.940 170.195 ;
        RECT 109.020 170.135 109.340 170.195 ;
        RECT 90.620 169.995 106.490 170.135 ;
        RECT 90.620 169.935 90.940 169.995 ;
        RECT 93.930 169.840 94.070 169.995 ;
        RECT 106.350 169.855 106.490 169.995 ;
        RECT 109.020 169.995 110.630 170.135 ;
        RECT 133.700 170.120 134.930 170.600 ;
        RECT 109.020 169.935 109.340 169.995 ;
        RECT 93.855 169.610 94.145 169.840 ;
        RECT 96.155 169.795 96.445 169.840 ;
        RECT 96.600 169.795 96.920 169.855 ;
        RECT 96.155 169.655 96.920 169.795 ;
        RECT 96.155 169.610 96.445 169.655 ;
        RECT 96.600 169.595 96.920 169.655 ;
        RECT 106.260 169.795 106.580 169.855 ;
        RECT 110.490 169.840 110.630 169.995 ;
        RECT 108.575 169.795 108.865 169.840 ;
        RECT 106.260 169.655 108.865 169.795 ;
        RECT 106.260 169.595 106.580 169.655 ;
        RECT 108.575 169.610 108.865 169.655 ;
        RECT 109.955 169.610 110.245 169.840 ;
        RECT 110.415 169.610 110.705 169.840 ;
        RECT 110.030 169.455 110.170 169.610 ;
        RECT 113.620 169.455 113.940 169.515 ;
        RECT 90.250 169.315 113.940 169.455 ;
        RECT 86.020 169.255 86.340 169.315 ;
        RECT 89.255 169.270 89.545 169.315 ;
        RECT 113.620 169.255 113.940 169.315 ;
        RECT 72.680 168.975 77.050 169.115 ;
        RECT 79.135 169.115 79.425 169.160 ;
        RECT 81.880 169.115 82.200 169.175 ;
        RECT 79.135 168.975 82.200 169.115 ;
        RECT 72.680 168.915 73.000 168.975 ;
        RECT 79.135 168.930 79.425 168.975 ;
        RECT 81.880 168.915 82.200 168.975 ;
        RECT 84.150 169.115 84.440 169.160 ;
        RECT 86.930 169.115 87.220 169.160 ;
        RECT 88.790 169.115 89.080 169.160 ;
        RECT 84.150 168.975 89.080 169.115 ;
        RECT 84.150 168.930 84.440 168.975 ;
        RECT 86.930 168.930 87.220 168.975 ;
        RECT 88.790 168.930 89.080 168.975 ;
        RECT 75.440 168.775 75.760 168.835 ;
        RECT 71.390 168.635 75.760 168.775 ;
        RECT 55.200 168.575 55.520 168.635 ;
        RECT 61.655 168.590 61.945 168.635 ;
        RECT 64.400 168.575 64.720 168.635 ;
        RECT 75.440 168.575 75.760 168.635 ;
        RECT 97.060 168.775 97.380 168.835 ;
        RECT 99.360 168.775 99.680 168.835 ;
        RECT 97.060 168.635 99.680 168.775 ;
        RECT 97.060 168.575 97.380 168.635 ;
        RECT 99.360 168.575 99.680 168.635 ;
        RECT 11.430 167.955 118.610 168.435 ;
        RECT 21.160 167.755 21.480 167.815 ;
        RECT 21.160 167.615 26.450 167.755 ;
        RECT 21.160 167.555 21.480 167.615 ;
        RECT 14.735 167.230 15.025 167.460 ;
        RECT 18.515 167.415 18.805 167.460 ;
        RECT 21.635 167.415 21.925 167.460 ;
        RECT 23.525 167.415 23.815 167.460 ;
        RECT 18.515 167.275 23.815 167.415 ;
        RECT 18.515 167.230 18.805 167.275 ;
        RECT 21.635 167.230 21.925 167.275 ;
        RECT 23.525 167.230 23.815 167.275 ;
        RECT 14.810 167.075 14.950 167.230 ;
        RECT 23.015 167.075 23.305 167.120 ;
        RECT 14.810 166.935 23.305 167.075 ;
        RECT 23.015 166.890 23.305 166.935 ;
        RECT 24.395 167.075 24.685 167.120 ;
        RECT 25.760 167.075 26.080 167.135 ;
        RECT 26.310 167.120 26.450 167.615 ;
        RECT 34.040 167.555 34.360 167.815 ;
        RECT 39.100 167.755 39.420 167.815 ;
        RECT 76.820 167.800 77.140 167.815 ;
        RECT 39.100 167.615 65.090 167.755 ;
        RECT 39.100 167.555 39.420 167.615 ;
        RECT 29.455 167.415 29.745 167.460 ;
        RECT 40.020 167.415 40.340 167.475 ;
        RECT 43.240 167.415 43.560 167.475 ;
        RECT 44.160 167.415 44.480 167.475 ;
        RECT 64.950 167.460 65.090 167.615 ;
        RECT 76.820 167.570 77.355 167.800 ;
        RECT 76.820 167.555 77.140 167.570 ;
        RECT 29.455 167.275 35.190 167.415 ;
        RECT 29.455 167.230 29.745 167.275 ;
        RECT 24.395 166.935 26.080 167.075 ;
        RECT 24.395 166.890 24.685 166.935 ;
        RECT 25.760 166.875 26.080 166.935 ;
        RECT 26.235 167.075 26.525 167.120 ;
        RECT 30.375 167.075 30.665 167.120 ;
        RECT 32.660 167.075 32.980 167.135 ;
        RECT 33.580 167.075 33.900 167.135 ;
        RECT 26.235 166.935 33.900 167.075 ;
        RECT 26.235 166.890 26.525 166.935 ;
        RECT 30.375 166.890 30.665 166.935 ;
        RECT 32.660 166.875 32.980 166.935 ;
        RECT 33.580 166.875 33.900 166.935 ;
        RECT 35.050 166.780 35.190 167.275 ;
        RECT 40.020 167.275 44.480 167.415 ;
        RECT 40.020 167.215 40.340 167.275 ;
        RECT 43.240 167.215 43.560 167.275 ;
        RECT 44.160 167.215 44.480 167.275 ;
        RECT 57.470 167.415 57.760 167.460 ;
        RECT 60.250 167.415 60.540 167.460 ;
        RECT 62.110 167.415 62.400 167.460 ;
        RECT 57.470 167.275 62.400 167.415 ;
        RECT 57.470 167.230 57.760 167.275 ;
        RECT 60.250 167.230 60.540 167.275 ;
        RECT 62.110 167.230 62.400 167.275 ;
        RECT 64.875 167.415 65.165 167.460 ;
        RECT 74.520 167.415 74.840 167.475 ;
        RECT 64.875 167.275 74.840 167.415 ;
        RECT 64.875 167.230 65.165 167.275 ;
        RECT 74.520 167.215 74.840 167.275 ;
        RECT 80.930 167.415 81.220 167.460 ;
        RECT 83.710 167.415 84.000 167.460 ;
        RECT 85.570 167.415 85.860 167.460 ;
        RECT 80.930 167.275 85.860 167.415 ;
        RECT 80.930 167.230 81.220 167.275 ;
        RECT 83.710 167.230 84.000 167.275 ;
        RECT 85.570 167.230 85.860 167.275 ;
        RECT 48.300 167.075 48.620 167.135 ;
        RECT 51.995 167.075 52.285 167.120 ;
        RECT 48.300 166.935 52.285 167.075 ;
        RECT 48.300 166.875 48.620 166.935 ;
        RECT 51.995 166.890 52.285 166.935 ;
        RECT 54.280 167.075 54.600 167.135 ;
        RECT 60.735 167.075 61.025 167.120 ;
        RECT 54.280 166.935 61.025 167.075 ;
        RECT 54.280 166.875 54.600 166.935 ;
        RECT 60.735 166.890 61.025 166.935 ;
        RECT 63.480 167.075 63.800 167.135 ;
        RECT 63.480 166.935 67.390 167.075 ;
        RECT 63.480 166.875 63.800 166.935 ;
        RECT 13.815 166.735 14.105 166.780 ;
        RECT 13.815 166.595 16.330 166.735 ;
        RECT 13.815 166.550 14.105 166.595 ;
        RECT 15.640 165.855 15.960 166.115 ;
        RECT 16.190 166.055 16.330 166.595 ;
        RECT 16.560 166.395 16.880 166.455 ;
        RECT 17.435 166.440 17.725 166.755 ;
        RECT 18.515 166.735 18.805 166.780 ;
        RECT 22.095 166.735 22.385 166.780 ;
        RECT 23.930 166.735 24.220 166.780 ;
        RECT 27.615 166.735 27.905 166.780 ;
        RECT 18.515 166.595 24.220 166.735 ;
        RECT 18.515 166.550 18.805 166.595 ;
        RECT 22.095 166.550 22.385 166.595 ;
        RECT 23.930 166.550 24.220 166.595 ;
        RECT 24.470 166.595 34.730 166.735 ;
        RECT 17.135 166.395 17.725 166.440 ;
        RECT 20.375 166.395 21.025 166.440 ;
        RECT 16.560 166.255 21.025 166.395 ;
        RECT 16.560 166.195 16.880 166.255 ;
        RECT 17.135 166.210 17.425 166.255 ;
        RECT 20.375 166.210 21.025 166.255 ;
        RECT 21.620 166.395 21.940 166.455 ;
        RECT 24.470 166.395 24.610 166.595 ;
        RECT 27.615 166.550 27.905 166.595 ;
        RECT 21.620 166.255 24.610 166.395 ;
        RECT 26.220 166.395 26.540 166.455 ;
        RECT 27.155 166.395 27.445 166.440 ;
        RECT 31.755 166.395 32.045 166.440 ;
        RECT 34.040 166.395 34.360 166.455 ;
        RECT 26.220 166.255 34.360 166.395 ;
        RECT 34.590 166.395 34.730 166.595 ;
        RECT 34.975 166.550 35.265 166.780 ;
        RECT 39.560 166.735 39.880 166.795 ;
        RECT 47.395 166.735 47.685 166.780 ;
        RECT 50.140 166.735 50.460 166.795 ;
        RECT 39.560 166.595 50.460 166.735 ;
        RECT 39.560 166.535 39.880 166.595 ;
        RECT 47.395 166.550 47.685 166.595 ;
        RECT 50.140 166.535 50.460 166.595 ;
        RECT 51.075 166.735 51.365 166.780 ;
        RECT 52.900 166.735 53.220 166.795 ;
        RECT 53.605 166.735 53.895 166.780 ;
        RECT 51.075 166.595 53.895 166.735 ;
        RECT 51.075 166.550 51.365 166.595 ;
        RECT 52.900 166.535 53.220 166.595 ;
        RECT 53.605 166.550 53.895 166.595 ;
        RECT 57.470 166.735 57.760 166.780 ;
        RECT 57.470 166.595 60.005 166.735 ;
        RECT 57.470 166.550 57.760 166.595 ;
        RECT 40.480 166.395 40.800 166.455 ;
        RECT 34.590 166.255 40.800 166.395 ;
        RECT 21.620 166.195 21.940 166.255 ;
        RECT 26.220 166.195 26.540 166.255 ;
        RECT 27.155 166.210 27.445 166.255 ;
        RECT 31.755 166.210 32.045 166.255 ;
        RECT 34.040 166.195 34.360 166.255 ;
        RECT 40.480 166.195 40.800 166.255 ;
        RECT 46.015 166.395 46.305 166.440 ;
        RECT 48.760 166.395 49.080 166.455 ;
        RECT 58.880 166.440 59.200 166.455 ;
        RECT 46.015 166.255 49.080 166.395 ;
        RECT 46.015 166.210 46.305 166.255 ;
        RECT 48.760 166.195 49.080 166.255 ;
        RECT 55.610 166.395 55.900 166.440 ;
        RECT 58.870 166.395 59.200 166.440 ;
        RECT 55.610 166.255 59.200 166.395 ;
        RECT 55.610 166.210 55.900 166.255 ;
        RECT 58.870 166.210 59.200 166.255 ;
        RECT 59.790 166.440 60.005 166.595 ;
        RECT 62.575 166.550 62.865 166.780 ;
        RECT 59.790 166.395 60.080 166.440 ;
        RECT 61.650 166.395 61.940 166.440 ;
        RECT 59.790 166.255 61.940 166.395 ;
        RECT 59.790 166.210 60.080 166.255 ;
        RECT 61.650 166.210 61.940 166.255 ;
        RECT 58.880 166.195 59.200 166.210 ;
        RECT 18.400 166.055 18.720 166.115 ;
        RECT 16.190 165.915 18.720 166.055 ;
        RECT 18.400 165.855 18.720 165.915 ;
        RECT 31.280 165.855 31.600 166.115 ;
        RECT 33.595 166.055 33.885 166.100 ;
        RECT 34.500 166.055 34.820 166.115 ;
        RECT 33.595 165.915 34.820 166.055 ;
        RECT 33.595 165.870 33.885 165.915 ;
        RECT 34.500 165.855 34.820 165.915 ;
        RECT 49.220 165.855 49.540 166.115 ;
        RECT 49.680 166.055 50.000 166.115 ;
        RECT 51.535 166.055 51.825 166.100 ;
        RECT 49.680 165.915 51.825 166.055 ;
        RECT 49.680 165.855 50.000 165.915 ;
        RECT 51.535 165.870 51.825 165.915 ;
        RECT 53.820 166.055 54.140 166.115 ;
        RECT 62.650 166.055 62.790 166.550 ;
        RECT 63.940 166.535 64.260 166.795 ;
        RECT 67.250 166.780 67.390 166.935 ;
        RECT 84.180 166.875 84.500 167.135 ;
        RECT 67.175 166.735 67.465 166.780 ;
        RECT 69.015 166.735 69.305 166.780 ;
        RECT 67.175 166.595 69.305 166.735 ;
        RECT 67.175 166.550 67.465 166.595 ;
        RECT 69.015 166.550 69.305 166.595 ;
        RECT 80.930 166.735 81.220 166.780 ;
        RECT 80.930 166.595 83.465 166.735 ;
        RECT 80.930 166.550 81.220 166.595 ;
        RECT 64.400 166.395 64.720 166.455 ;
        RECT 79.070 166.395 79.360 166.440 ;
        RECT 79.580 166.395 79.900 166.455 ;
        RECT 83.250 166.440 83.465 166.595 ;
        RECT 86.020 166.535 86.340 166.795 ;
        RECT 92.920 166.735 93.240 166.795 ;
        RECT 93.855 166.735 94.145 166.780 ;
        RECT 92.920 166.595 94.145 166.735 ;
        RECT 92.920 166.535 93.240 166.595 ;
        RECT 93.855 166.550 94.145 166.595 ;
        RECT 94.760 166.535 95.080 166.795 ;
        RECT 95.235 166.550 95.525 166.780 ;
        RECT 95.695 166.550 95.985 166.780 ;
        RECT 82.330 166.395 82.620 166.440 ;
        RECT 64.400 166.255 78.890 166.395 ;
        RECT 64.400 166.195 64.720 166.255 ;
        RECT 53.820 165.915 62.790 166.055 ;
        RECT 53.820 165.855 54.140 165.915 ;
        RECT 68.080 165.855 68.400 166.115 ;
        RECT 69.920 165.855 70.240 166.115 ;
        RECT 78.750 166.055 78.890 166.255 ;
        RECT 79.070 166.255 82.620 166.395 ;
        RECT 79.070 166.210 79.360 166.255 ;
        RECT 79.580 166.195 79.900 166.255 ;
        RECT 82.330 166.210 82.620 166.255 ;
        RECT 83.250 166.395 83.540 166.440 ;
        RECT 85.110 166.395 85.400 166.440 ;
        RECT 95.310 166.395 95.450 166.550 ;
        RECT 83.250 166.255 85.400 166.395 ;
        RECT 83.250 166.210 83.540 166.255 ;
        RECT 85.110 166.210 85.400 166.255 ;
        RECT 93.930 166.255 95.450 166.395 ;
        RECT 93.930 166.115 94.070 166.255 ;
        RECT 90.620 166.055 90.940 166.115 ;
        RECT 78.750 165.915 90.940 166.055 ;
        RECT 90.620 165.855 90.940 165.915 ;
        RECT 93.840 165.855 94.160 166.115 ;
        RECT 94.300 166.055 94.620 166.115 ;
        RECT 95.770 166.055 95.910 166.550 ;
        RECT 94.300 165.915 95.910 166.055 ;
        RECT 97.075 166.055 97.365 166.100 ;
        RECT 97.980 166.055 98.300 166.115 ;
        RECT 97.075 165.915 98.300 166.055 ;
        RECT 94.300 165.855 94.620 165.915 ;
        RECT 97.075 165.870 97.365 165.915 ;
        RECT 97.980 165.855 98.300 165.915 ;
        RECT 10.650 165.235 118.610 165.715 ;
        RECT 135.580 165.470 136.830 166.590 ;
        RECT 15.640 165.035 15.960 165.095 ;
        RECT 15.640 164.895 16.330 165.035 ;
        RECT 15.640 164.835 15.960 164.895 ;
        RECT 16.190 164.695 16.330 164.895 ;
        RECT 18.400 164.835 18.720 165.095 ;
        RECT 20.715 165.035 21.005 165.080 ;
        RECT 43.700 165.035 44.020 165.095 ;
        RECT 20.715 164.895 44.020 165.035 ;
        RECT 20.715 164.850 21.005 164.895 ;
        RECT 20.790 164.695 20.930 164.850 ;
        RECT 43.700 164.835 44.020 164.895 ;
        RECT 46.000 165.035 46.320 165.095 ;
        RECT 47.395 165.035 47.685 165.080 ;
        RECT 46.000 164.895 47.685 165.035 ;
        RECT 46.000 164.835 46.320 164.895 ;
        RECT 47.395 164.850 47.685 164.895 ;
        RECT 60.260 164.835 60.580 165.095 ;
        RECT 62.115 165.035 62.405 165.080 ;
        RECT 90.160 165.035 90.480 165.095 ;
        RECT 62.115 164.895 72.910 165.035 ;
        RECT 62.115 164.850 62.405 164.895 ;
        RECT 32.200 164.740 32.520 164.755 ;
        RECT 16.190 164.555 20.930 164.695 ;
        RECT 29.460 164.695 29.750 164.740 ;
        RECT 31.320 164.695 31.610 164.740 ;
        RECT 29.460 164.555 31.610 164.695 ;
        RECT 29.460 164.510 29.750 164.555 ;
        RECT 31.320 164.510 31.610 164.555 ;
        RECT 14.720 164.355 15.040 164.415 ;
        RECT 15.655 164.355 15.945 164.400 ;
        RECT 14.720 164.215 15.945 164.355 ;
        RECT 14.720 164.155 15.040 164.215 ;
        RECT 15.655 164.170 15.945 164.215 ;
        RECT 17.020 164.155 17.340 164.415 ;
        RECT 20.255 164.355 20.545 164.400 ;
        RECT 20.700 164.355 21.020 164.415 ;
        RECT 20.255 164.215 21.020 164.355 ;
        RECT 20.255 164.170 20.545 164.215 ;
        RECT 20.700 164.155 21.020 164.215 ;
        RECT 25.760 164.355 26.080 164.415 ;
        RECT 28.535 164.355 28.825 164.400 ;
        RECT 25.760 164.215 28.825 164.355 ;
        RECT 31.395 164.355 31.610 164.510 ;
        RECT 32.200 164.695 32.530 164.740 ;
        RECT 35.500 164.695 35.790 164.740 ;
        RECT 46.460 164.695 46.780 164.755 ;
        RECT 55.200 164.695 55.520 164.755 ;
        RECT 59.815 164.695 60.105 164.740 ;
        RECT 62.805 164.695 63.095 164.740 ;
        RECT 32.200 164.555 35.790 164.695 ;
        RECT 32.200 164.510 32.530 164.555 ;
        RECT 35.500 164.510 35.790 164.555 ;
        RECT 45.630 164.555 55.520 164.695 ;
        RECT 32.200 164.495 32.520 164.510 ;
        RECT 33.640 164.355 33.930 164.400 ;
        RECT 31.395 164.215 33.930 164.355 ;
        RECT 25.760 164.155 26.080 164.215 ;
        RECT 28.535 164.170 28.825 164.215 ;
        RECT 33.640 164.170 33.930 164.215 ;
        RECT 40.020 164.155 40.340 164.415 ;
        RECT 40.480 164.355 40.800 164.415 ;
        RECT 40.955 164.355 41.245 164.400 ;
        RECT 40.480 164.215 41.245 164.355 ;
        RECT 40.480 164.155 40.800 164.215 ;
        RECT 40.955 164.170 41.245 164.215 ;
        RECT 41.415 164.170 41.705 164.400 ;
        RECT 21.160 163.815 21.480 164.075 ;
        RECT 30.360 163.815 30.680 164.075 ;
        RECT 37.505 164.015 37.795 164.060 ;
        RECT 38.180 164.015 38.500 164.075 ;
        RECT 37.505 163.875 38.500 164.015 ;
        RECT 41.490 164.015 41.630 164.170 ;
        RECT 41.860 164.155 42.180 164.415 ;
        RECT 43.700 164.155 44.020 164.415 ;
        RECT 44.620 164.155 44.940 164.415 ;
        RECT 45.630 164.400 45.770 164.555 ;
        RECT 46.460 164.495 46.780 164.555 ;
        RECT 55.200 164.495 55.520 164.555 ;
        RECT 57.130 164.555 63.095 164.695 ;
        RECT 45.095 164.170 45.385 164.400 ;
        RECT 45.555 164.170 45.845 164.400 ;
        RECT 48.315 164.355 48.605 164.400 ;
        RECT 49.220 164.355 49.540 164.415 ;
        RECT 48.315 164.215 49.540 164.355 ;
        RECT 48.315 164.170 48.605 164.215 ;
        RECT 45.170 164.015 45.310 164.170 ;
        RECT 49.220 164.155 49.540 164.215 ;
        RECT 54.740 164.355 55.060 164.415 ;
        RECT 56.135 164.355 56.425 164.400 ;
        RECT 54.740 164.215 56.425 164.355 ;
        RECT 54.740 164.155 55.060 164.215 ;
        RECT 56.135 164.170 56.425 164.215 ;
        RECT 56.580 164.155 56.900 164.415 ;
        RECT 57.130 164.400 57.270 164.555 ;
        RECT 59.815 164.510 60.105 164.555 ;
        RECT 62.805 164.510 63.095 164.555 ;
        RECT 64.810 164.695 65.100 164.740 ;
        RECT 67.160 164.695 67.480 164.755 ;
        RECT 68.070 164.695 68.360 164.740 ;
        RECT 64.810 164.555 68.360 164.695 ;
        RECT 64.810 164.510 65.100 164.555 ;
        RECT 67.160 164.495 67.480 164.555 ;
        RECT 68.070 164.510 68.360 164.555 ;
        RECT 68.990 164.695 69.280 164.740 ;
        RECT 70.850 164.695 71.140 164.740 ;
        RECT 68.990 164.555 71.140 164.695 ;
        RECT 68.990 164.510 69.280 164.555 ;
        RECT 70.850 164.510 71.140 164.555 ;
        RECT 57.055 164.170 57.345 164.400 ;
        RECT 57.960 164.155 58.280 164.415 ;
        RECT 66.670 164.355 66.960 164.400 ;
        RECT 68.990 164.355 69.205 164.510 ;
        RECT 66.670 164.215 69.205 164.355 ;
        RECT 66.670 164.170 66.960 164.215 ;
        RECT 69.935 164.170 70.225 164.400 ;
        RECT 71.775 164.355 72.065 164.400 ;
        RECT 72.770 164.355 72.910 164.895 ;
        RECT 89.790 164.895 90.480 165.035 ;
        RECT 73.155 164.355 73.445 164.400 ;
        RECT 71.775 164.215 72.450 164.355 ;
        RECT 72.770 164.215 73.445 164.355 ;
        RECT 71.775 164.170 72.065 164.215 ;
        RECT 41.490 163.875 45.310 164.015 ;
        RECT 51.995 164.015 52.285 164.060 ;
        RECT 52.900 164.015 53.220 164.075 ;
        RECT 51.995 163.875 53.220 164.015 ;
        RECT 37.505 163.830 37.795 163.875 ;
        RECT 38.180 163.815 38.500 163.875 ;
        RECT 44.250 163.735 44.390 163.875 ;
        RECT 51.995 163.830 52.285 163.875 ;
        RECT 52.900 163.815 53.220 163.875 ;
        RECT 59.355 164.015 59.645 164.060 ;
        RECT 60.260 164.015 60.580 164.075 ;
        RECT 59.355 163.875 60.580 164.015 ;
        RECT 70.010 164.015 70.150 164.170 ;
        RECT 72.310 164.015 72.450 164.215 ;
        RECT 73.155 164.170 73.445 164.215 ;
        RECT 88.780 164.155 89.100 164.415 ;
        RECT 89.790 164.400 89.930 164.895 ;
        RECT 90.160 164.835 90.480 164.895 ;
        RECT 90.620 165.035 90.940 165.095 ;
        RECT 94.300 165.035 94.620 165.095 ;
        RECT 102.135 165.035 102.425 165.080 ;
        RECT 113.160 165.035 113.480 165.095 ;
        RECT 90.620 164.895 98.210 165.035 ;
        RECT 90.620 164.835 90.940 164.895 ;
        RECT 94.300 164.835 94.620 164.895 ;
        RECT 94.760 164.695 95.080 164.755 ;
        RECT 94.760 164.555 97.750 164.695 ;
        RECT 94.760 164.495 95.080 164.555 ;
        RECT 89.715 164.170 90.005 164.400 ;
        RECT 90.160 164.155 90.480 164.415 ;
        RECT 90.620 164.155 90.940 164.415 ;
        RECT 92.475 164.170 92.765 164.400 ;
        RECT 86.020 164.015 86.340 164.075 ;
        RECT 70.010 163.875 71.990 164.015 ;
        RECT 72.310 163.875 86.340 164.015 ;
        RECT 88.870 164.015 89.010 164.155 ;
        RECT 92.550 164.015 92.690 164.170 ;
        RECT 93.380 164.155 93.700 164.415 ;
        RECT 93.840 164.155 94.160 164.415 ;
        RECT 94.300 164.155 94.620 164.415 ;
        RECT 96.155 164.170 96.445 164.400 ;
        RECT 92.920 164.015 93.240 164.075 ;
        RECT 96.230 164.015 96.370 164.170 ;
        RECT 97.060 164.155 97.380 164.415 ;
        RECT 97.610 164.400 97.750 164.555 ;
        RECT 98.070 164.400 98.210 164.895 ;
        RECT 102.135 164.895 113.480 165.035 ;
        RECT 102.135 164.850 102.425 164.895 ;
        RECT 113.160 164.835 113.480 164.895 ;
        RECT 108.675 164.695 108.965 164.740 ;
        RECT 111.915 164.695 112.565 164.740 ;
        RECT 106.350 164.555 112.565 164.695 ;
        RECT 97.535 164.170 97.825 164.400 ;
        RECT 97.995 164.170 98.285 164.400 ;
        RECT 99.820 164.155 100.140 164.415 ;
        RECT 101.200 164.155 101.520 164.415 ;
        RECT 105.800 164.155 106.120 164.415 ;
        RECT 106.350 164.400 106.490 164.555 ;
        RECT 108.675 164.510 109.265 164.555 ;
        RECT 111.915 164.510 112.565 164.555 ;
        RECT 106.275 164.170 106.565 164.400 ;
        RECT 108.975 164.195 109.265 164.510 ;
        RECT 110.055 164.355 110.345 164.400 ;
        RECT 113.635 164.355 113.925 164.400 ;
        RECT 115.470 164.355 115.760 164.400 ;
        RECT 110.055 164.215 115.760 164.355 ;
        RECT 110.055 164.170 110.345 164.215 ;
        RECT 113.635 164.170 113.925 164.215 ;
        RECT 115.470 164.170 115.760 164.215 ;
        RECT 88.870 163.875 96.370 164.015 ;
        RECT 96.600 164.015 96.920 164.075 ;
        RECT 100.755 164.015 101.045 164.060 ;
        RECT 96.600 163.875 101.045 164.015 ;
        RECT 59.355 163.830 59.645 163.875 ;
        RECT 60.260 163.815 60.580 163.875 ;
        RECT 29.000 163.675 29.290 163.720 ;
        RECT 30.860 163.675 31.150 163.720 ;
        RECT 33.640 163.675 33.930 163.720 ;
        RECT 29.000 163.535 33.930 163.675 ;
        RECT 29.000 163.490 29.290 163.535 ;
        RECT 30.860 163.490 31.150 163.535 ;
        RECT 33.640 163.490 33.930 163.535 ;
        RECT 44.160 163.675 44.480 163.735 ;
        RECT 66.670 163.675 66.960 163.720 ;
        RECT 69.450 163.675 69.740 163.720 ;
        RECT 71.310 163.675 71.600 163.720 ;
        RECT 44.160 163.535 55.430 163.675 ;
        RECT 44.160 163.475 44.480 163.535 ;
        RECT 16.100 163.135 16.420 163.395 ;
        RECT 17.955 163.335 18.245 163.380 ;
        RECT 23.000 163.335 23.320 163.395 ;
        RECT 17.955 163.195 23.320 163.335 ;
        RECT 17.955 163.150 18.245 163.195 ;
        RECT 23.000 163.135 23.320 163.195 ;
        RECT 34.040 163.335 34.360 163.395 ;
        RECT 37.720 163.335 38.040 163.395 ;
        RECT 34.040 163.195 38.040 163.335 ;
        RECT 34.040 163.135 34.360 163.195 ;
        RECT 37.720 163.135 38.040 163.195 ;
        RECT 43.240 163.135 43.560 163.395 ;
        RECT 46.460 163.335 46.780 163.395 ;
        RECT 46.935 163.335 47.225 163.380 ;
        RECT 46.460 163.195 47.225 163.335 ;
        RECT 46.460 163.135 46.780 163.195 ;
        RECT 46.935 163.150 47.225 163.195 ;
        RECT 47.380 163.335 47.700 163.395 ;
        RECT 48.775 163.335 49.065 163.380 ;
        RECT 47.380 163.195 49.065 163.335 ;
        RECT 47.380 163.135 47.700 163.195 ;
        RECT 48.775 163.150 49.065 163.195 ;
        RECT 49.220 163.335 49.540 163.395 ;
        RECT 54.755 163.335 55.045 163.380 ;
        RECT 49.220 163.195 55.045 163.335 ;
        RECT 55.290 163.335 55.430 163.535 ;
        RECT 66.670 163.535 71.600 163.675 ;
        RECT 71.850 163.675 71.990 163.875 ;
        RECT 86.020 163.815 86.340 163.875 ;
        RECT 92.920 163.815 93.240 163.875 ;
        RECT 96.600 163.815 96.920 163.875 ;
        RECT 100.755 163.830 101.045 163.875 ;
        RECT 114.540 163.815 114.860 164.075 ;
        RECT 115.935 164.015 116.225 164.060 ;
        RECT 116.380 164.015 116.700 164.075 ;
        RECT 115.935 163.875 116.700 164.015 ;
        RECT 115.935 163.830 116.225 163.875 ;
        RECT 116.380 163.815 116.700 163.875 ;
        RECT 72.235 163.675 72.525 163.720 ;
        RECT 93.840 163.675 94.160 163.735 ;
        RECT 94.760 163.675 95.080 163.735 ;
        RECT 71.850 163.535 72.525 163.675 ;
        RECT 66.670 163.490 66.960 163.535 ;
        RECT 69.450 163.490 69.740 163.535 ;
        RECT 71.310 163.490 71.600 163.535 ;
        RECT 72.235 163.490 72.525 163.535 ;
        RECT 90.250 163.535 95.080 163.675 ;
        RECT 90.250 163.395 90.390 163.535 ;
        RECT 93.840 163.475 94.160 163.535 ;
        RECT 94.760 163.475 95.080 163.535 ;
        RECT 110.055 163.675 110.345 163.720 ;
        RECT 113.175 163.675 113.465 163.720 ;
        RECT 115.065 163.675 115.355 163.720 ;
        RECT 110.055 163.535 115.355 163.675 ;
        RECT 110.055 163.490 110.345 163.535 ;
        RECT 113.175 163.490 113.465 163.535 ;
        RECT 115.065 163.490 115.355 163.535 ;
        RECT 69.920 163.335 70.240 163.395 ;
        RECT 90.160 163.335 90.480 163.395 ;
        RECT 55.290 163.195 90.480 163.335 ;
        RECT 49.220 163.135 49.540 163.195 ;
        RECT 54.755 163.150 55.045 163.195 ;
        RECT 69.920 163.135 70.240 163.195 ;
        RECT 90.160 163.135 90.480 163.195 ;
        RECT 92.015 163.335 92.305 163.380 ;
        RECT 93.380 163.335 93.700 163.395 ;
        RECT 92.015 163.195 93.700 163.335 ;
        RECT 92.015 163.150 92.305 163.195 ;
        RECT 93.380 163.135 93.700 163.195 ;
        RECT 95.680 163.135 96.000 163.395 ;
        RECT 99.360 163.135 99.680 163.395 ;
        RECT 100.280 163.135 100.600 163.395 ;
        RECT 107.180 163.135 107.500 163.395 ;
        RECT 11.430 162.515 118.610 162.995 ;
        RECT 31.280 162.315 31.600 162.375 ;
        RECT 32.200 162.315 32.520 162.375 ;
        RECT 38.180 162.315 38.500 162.375 ;
        RECT 50.155 162.315 50.445 162.360 ;
        RECT 54.280 162.315 54.600 162.375 ;
        RECT 31.280 162.175 43.010 162.315 ;
        RECT 31.280 162.115 31.600 162.175 ;
        RECT 32.200 162.115 32.520 162.175 ;
        RECT 38.180 162.115 38.500 162.175 ;
        RECT 18.515 161.975 18.805 162.020 ;
        RECT 21.635 161.975 21.925 162.020 ;
        RECT 23.525 161.975 23.815 162.020 ;
        RECT 18.515 161.835 23.815 161.975 ;
        RECT 18.515 161.790 18.805 161.835 ;
        RECT 21.635 161.790 21.925 161.835 ;
        RECT 23.525 161.790 23.815 161.835 ;
        RECT 30.360 161.975 30.680 162.035 ;
        RECT 33.595 161.975 33.885 162.020 ;
        RECT 42.320 161.975 42.640 162.035 ;
        RECT 30.360 161.835 33.885 161.975 ;
        RECT 30.360 161.775 30.680 161.835 ;
        RECT 33.595 161.790 33.885 161.835 ;
        RECT 37.350 161.835 42.640 161.975 ;
        RECT 15.655 161.635 15.945 161.680 ;
        RECT 20.700 161.635 21.020 161.695 ;
        RECT 15.655 161.495 21.020 161.635 ;
        RECT 15.655 161.450 15.945 161.495 ;
        RECT 20.700 161.435 21.020 161.495 ;
        RECT 23.000 161.435 23.320 161.695 ;
        RECT 24.395 161.635 24.685 161.680 ;
        RECT 25.760 161.635 26.080 161.695 ;
        RECT 24.395 161.495 26.080 161.635 ;
        RECT 24.395 161.450 24.685 161.495 ;
        RECT 25.760 161.435 26.080 161.495 ;
        RECT 16.100 160.955 16.420 161.015 ;
        RECT 17.435 161.000 17.725 161.315 ;
        RECT 18.515 161.295 18.805 161.340 ;
        RECT 22.095 161.295 22.385 161.340 ;
        RECT 23.930 161.295 24.220 161.340 ;
        RECT 18.515 161.155 24.220 161.295 ;
        RECT 18.515 161.110 18.805 161.155 ;
        RECT 22.095 161.110 22.385 161.155 ;
        RECT 23.930 161.110 24.220 161.155 ;
        RECT 34.500 161.095 34.820 161.355 ;
        RECT 37.350 161.340 37.490 161.835 ;
        RECT 42.320 161.775 42.640 161.835 ;
        RECT 37.720 161.635 38.040 161.695 ;
        RECT 42.870 161.635 43.010 162.175 ;
        RECT 50.155 162.175 54.600 162.315 ;
        RECT 50.155 162.130 50.445 162.175 ;
        RECT 54.280 162.115 54.600 162.175 ;
        RECT 58.510 162.175 61.410 162.315 ;
        RECT 58.510 161.975 58.650 162.175 ;
        RECT 48.850 161.835 58.650 161.975 ;
        RECT 61.270 161.975 61.410 162.175 ;
        RECT 94.300 162.115 94.620 162.375 ;
        RECT 96.600 162.115 96.920 162.375 ;
        RECT 100.295 162.315 100.585 162.360 ;
        RECT 103.040 162.315 103.360 162.375 ;
        RECT 100.295 162.175 103.360 162.315 ;
        RECT 100.295 162.130 100.585 162.175 ;
        RECT 103.040 162.115 103.360 162.175 ;
        RECT 114.540 162.315 114.860 162.375 ;
        RECT 115.015 162.315 115.305 162.360 ;
        RECT 114.540 162.175 115.305 162.315 ;
        RECT 114.540 162.115 114.860 162.175 ;
        RECT 115.015 162.130 115.305 162.175 ;
        RECT 66.240 161.975 66.560 162.035 ;
        RECT 61.270 161.835 66.560 161.975 ;
        RECT 37.720 161.495 38.410 161.635 ;
        RECT 42.870 161.495 44.850 161.635 ;
        RECT 37.720 161.435 38.040 161.495 ;
        RECT 38.270 161.340 38.410 161.495 ;
        RECT 37.275 161.110 37.565 161.340 ;
        RECT 38.195 161.110 38.485 161.340 ;
        RECT 38.640 161.095 38.960 161.355 ;
        RECT 39.100 161.095 39.420 161.355 ;
        RECT 40.020 161.095 40.340 161.355 ;
        RECT 41.860 161.295 42.180 161.355 ;
        RECT 43.715 161.295 44.005 161.340 ;
        RECT 41.860 161.155 44.005 161.295 ;
        RECT 41.860 161.095 42.180 161.155 ;
        RECT 43.715 161.110 44.005 161.155 ;
        RECT 44.160 161.095 44.480 161.355 ;
        RECT 44.710 161.340 44.850 161.495 ;
        RECT 44.635 161.110 44.925 161.340 ;
        RECT 45.555 161.110 45.845 161.340 ;
        RECT 17.135 160.955 17.725 161.000 ;
        RECT 20.375 160.955 21.025 161.000 ;
        RECT 16.100 160.815 21.025 160.955 ;
        RECT 16.100 160.755 16.420 160.815 ;
        RECT 17.135 160.770 17.425 160.815 ;
        RECT 20.375 160.770 21.025 160.815 ;
        RECT 35.880 160.955 36.200 161.015 ;
        RECT 39.190 160.955 39.330 161.095 ;
        RECT 35.880 160.815 39.330 160.955 ;
        RECT 40.110 160.955 40.250 161.095 ;
        RECT 45.630 160.955 45.770 161.110 ;
        RECT 47.380 161.095 47.700 161.355 ;
        RECT 48.300 161.095 48.620 161.355 ;
        RECT 48.850 161.340 48.990 161.835 ;
        RECT 66.240 161.775 66.560 161.835 ;
        RECT 68.555 161.790 68.845 162.020 ;
        RECT 94.390 161.975 94.530 162.115 ;
        RECT 99.820 161.975 100.140 162.035 ;
        RECT 101.675 161.975 101.965 162.020 ;
        RECT 108.560 161.975 108.880 162.035 ;
        RECT 94.390 161.835 95.450 161.975 ;
        RECT 50.140 161.635 50.460 161.695 ;
        RECT 50.140 161.495 54.050 161.635 ;
        RECT 50.140 161.435 50.460 161.495 ;
        RECT 48.775 161.110 49.065 161.340 ;
        RECT 49.220 161.095 49.540 161.355 ;
        RECT 51.980 161.095 52.300 161.355 ;
        RECT 52.440 161.095 52.760 161.355 ;
        RECT 52.900 161.095 53.220 161.355 ;
        RECT 53.910 161.340 54.050 161.495 ;
        RECT 54.280 161.435 54.600 161.695 ;
        RECT 54.830 161.495 58.190 161.635 ;
        RECT 53.835 161.110 54.125 161.340 ;
        RECT 54.830 161.295 54.970 161.495 ;
        RECT 54.370 161.155 54.970 161.295 ;
        RECT 54.370 160.955 54.510 161.155 ;
        RECT 55.675 161.110 55.965 161.340 ;
        RECT 40.110 160.815 54.510 160.955 ;
        RECT 54.740 160.955 55.060 161.015 ;
        RECT 55.750 160.955 55.890 161.110 ;
        RECT 56.120 161.095 56.440 161.355 ;
        RECT 56.595 161.295 56.885 161.340 ;
        RECT 56.595 161.155 57.270 161.295 ;
        RECT 56.595 161.110 56.885 161.155 ;
        RECT 54.740 160.815 55.890 160.955 ;
        RECT 57.130 160.955 57.270 161.155 ;
        RECT 57.500 161.095 57.820 161.355 ;
        RECT 58.050 161.295 58.190 161.495 ;
        RECT 60.260 161.435 60.580 161.695 ;
        RECT 68.630 161.635 68.770 161.790 ;
        RECT 85.100 161.635 85.420 161.695 ;
        RECT 93.840 161.635 94.160 161.695 ;
        RECT 68.630 161.495 73.140 161.635 ;
        RECT 68.630 161.295 68.770 161.495 ;
        RECT 58.050 161.155 68.770 161.295 ;
        RECT 69.460 161.295 69.780 161.355 ;
        RECT 70.840 161.295 71.160 161.355 ;
        RECT 69.460 161.155 71.160 161.295 ;
        RECT 69.460 161.095 69.780 161.155 ;
        RECT 70.840 161.095 71.160 161.155 ;
        RECT 59.800 160.955 60.120 161.015 ;
        RECT 61.195 160.955 61.485 161.000 ;
        RECT 57.130 160.815 61.485 160.955 ;
        RECT 73.000 160.955 73.140 161.495 ;
        RECT 85.100 161.495 89.930 161.635 ;
        RECT 85.100 161.435 85.420 161.495 ;
        RECT 84.640 161.095 84.960 161.355 ;
        RECT 88.780 161.095 89.100 161.355 ;
        RECT 89.790 161.340 89.930 161.495 ;
        RECT 93.840 161.495 94.990 161.635 ;
        RECT 93.840 161.435 94.160 161.495 ;
        RECT 89.715 161.110 90.005 161.340 ;
        RECT 90.160 161.095 90.480 161.355 ;
        RECT 90.620 161.095 90.940 161.355 ;
        RECT 93.395 161.110 93.685 161.340 ;
        RECT 88.870 160.955 89.010 161.095 ;
        RECT 93.470 160.955 93.610 161.110 ;
        RECT 94.300 161.095 94.620 161.355 ;
        RECT 94.850 161.340 94.990 161.495 ;
        RECT 95.310 161.340 95.450 161.835 ;
        RECT 99.820 161.835 101.965 161.975 ;
        RECT 99.820 161.775 100.140 161.835 ;
        RECT 101.675 161.790 101.965 161.835 ;
        RECT 104.050 161.835 108.880 161.975 ;
        RECT 99.360 161.435 99.680 161.695 ;
        RECT 104.050 161.635 104.190 161.835 ;
        RECT 108.560 161.775 108.880 161.835 ;
        RECT 109.495 161.790 109.785 162.020 ;
        RECT 100.370 161.495 104.190 161.635 ;
        RECT 106.735 161.635 107.025 161.680 ;
        RECT 107.640 161.635 107.960 161.695 ;
        RECT 106.735 161.495 107.960 161.635 ;
        RECT 109.570 161.635 109.710 161.790 ;
        RECT 109.570 161.495 114.310 161.635 ;
        RECT 100.370 161.340 100.510 161.495 ;
        RECT 106.735 161.450 107.025 161.495 ;
        RECT 107.640 161.435 107.960 161.495 ;
        RECT 94.775 161.110 95.065 161.340 ;
        RECT 95.235 161.110 95.525 161.340 ;
        RECT 100.295 161.110 100.585 161.340 ;
        RECT 102.580 161.295 102.900 161.355 ;
        RECT 103.055 161.295 103.345 161.340 ;
        RECT 102.580 161.155 103.345 161.295 ;
        RECT 102.580 161.095 102.900 161.155 ;
        RECT 103.055 161.110 103.345 161.155 ;
        RECT 103.515 161.110 103.805 161.340 ;
        RECT 103.975 161.110 104.265 161.340 ;
        RECT 104.420 161.295 104.740 161.355 ;
        RECT 104.895 161.295 105.185 161.340 ;
        RECT 104.420 161.155 105.185 161.295 ;
        RECT 73.000 160.815 93.610 160.955 ;
        RECT 35.880 160.755 36.200 160.815 ;
        RECT 54.740 160.755 55.060 160.815 ;
        RECT 59.800 160.755 60.120 160.815 ;
        RECT 61.195 160.770 61.485 160.815 ;
        RECT 98.900 160.755 99.220 161.015 ;
        RECT 102.120 160.955 102.440 161.015 ;
        RECT 103.590 160.955 103.730 161.110 ;
        RECT 102.120 160.815 103.730 160.955 ;
        RECT 104.050 160.955 104.190 161.110 ;
        RECT 104.420 161.095 104.740 161.155 ;
        RECT 104.895 161.110 105.185 161.155 ;
        RECT 106.260 161.295 106.580 161.355 ;
        RECT 110.415 161.295 110.705 161.340 ;
        RECT 106.260 161.155 110.705 161.295 ;
        RECT 106.260 161.095 106.580 161.155 ;
        RECT 110.415 161.110 110.705 161.155 ;
        RECT 112.700 161.095 113.020 161.355 ;
        RECT 114.170 161.340 114.310 161.495 ;
        RECT 114.095 161.110 114.385 161.340 ;
        RECT 104.050 160.815 107.410 160.955 ;
        RECT 102.120 160.755 102.440 160.815 ;
        RECT 107.270 160.675 107.410 160.815 ;
        RECT 40.020 160.615 40.340 160.675 ;
        RECT 40.495 160.615 40.785 160.660 ;
        RECT 40.020 160.475 40.785 160.615 ;
        RECT 40.020 160.415 40.340 160.475 ;
        RECT 40.495 160.430 40.785 160.475 ;
        RECT 42.320 160.415 42.640 160.675 ;
        RECT 42.780 160.615 43.100 160.675 ;
        RECT 50.615 160.615 50.905 160.660 ;
        RECT 42.780 160.475 50.905 160.615 ;
        RECT 42.780 160.415 43.100 160.475 ;
        RECT 50.615 160.430 50.905 160.475 ;
        RECT 55.660 160.615 55.980 160.675 ;
        RECT 61.655 160.615 61.945 160.660 ;
        RECT 55.660 160.475 61.945 160.615 ;
        RECT 55.660 160.415 55.980 160.475 ;
        RECT 61.655 160.430 61.945 160.475 ;
        RECT 63.495 160.615 63.785 160.660 ;
        RECT 70.840 160.615 71.160 160.675 ;
        RECT 63.495 160.475 71.160 160.615 ;
        RECT 63.495 160.430 63.785 160.475 ;
        RECT 70.840 160.415 71.160 160.475 ;
        RECT 85.575 160.615 85.865 160.660 ;
        RECT 87.400 160.615 87.720 160.675 ;
        RECT 85.575 160.475 87.720 160.615 ;
        RECT 85.575 160.430 85.865 160.475 ;
        RECT 87.400 160.415 87.720 160.475 ;
        RECT 92.015 160.615 92.305 160.660 ;
        RECT 92.920 160.615 93.240 160.675 ;
        RECT 92.015 160.475 93.240 160.615 ;
        RECT 92.015 160.430 92.305 160.475 ;
        RECT 92.920 160.415 93.240 160.475 ;
        RECT 101.215 160.615 101.505 160.660 ;
        RECT 103.500 160.615 103.820 160.675 ;
        RECT 101.215 160.475 103.820 160.615 ;
        RECT 101.215 160.430 101.505 160.475 ;
        RECT 103.500 160.415 103.820 160.475 ;
        RECT 107.180 160.415 107.500 160.675 ;
        RECT 107.655 160.615 107.945 160.660 ;
        RECT 108.100 160.615 108.420 160.675 ;
        RECT 107.655 160.475 108.420 160.615 ;
        RECT 107.655 160.430 107.945 160.475 ;
        RECT 108.100 160.415 108.420 160.475 ;
        RECT 110.860 160.415 111.180 160.675 ;
        RECT 113.635 160.615 113.925 160.660 ;
        RECT 114.540 160.615 114.860 160.675 ;
        RECT 113.635 160.475 114.860 160.615 ;
        RECT 113.635 160.430 113.925 160.475 ;
        RECT 114.540 160.415 114.860 160.475 ;
        RECT 10.650 159.795 118.610 160.275 ;
        RECT 17.020 159.595 17.340 159.655 ;
        RECT 18.415 159.595 18.705 159.640 ;
        RECT 17.020 159.455 18.705 159.595 ;
        RECT 17.020 159.395 17.340 159.455 ;
        RECT 18.415 159.410 18.705 159.455 ;
        RECT 32.200 159.395 32.520 159.655 ;
        RECT 34.055 159.595 34.345 159.640 ;
        RECT 37.735 159.595 38.025 159.640 ;
        RECT 34.055 159.455 35.650 159.595 ;
        RECT 34.055 159.410 34.345 159.455 ;
        RECT 27.600 159.255 27.920 159.315 ;
        RECT 27.600 159.115 32.890 159.255 ;
        RECT 27.600 159.055 27.920 159.115 ;
        RECT 20.240 158.715 20.560 158.975 ;
        RECT 26.680 158.915 27.000 158.975 ;
        RECT 30.360 158.915 30.680 158.975 ;
        RECT 31.755 158.915 32.045 158.960 ;
        RECT 26.680 158.775 32.045 158.915 ;
        RECT 32.750 158.915 32.890 159.115 ;
        RECT 35.510 158.960 35.650 159.455 ;
        RECT 35.970 159.455 38.025 159.595 ;
        RECT 32.750 158.775 34.270 158.915 ;
        RECT 26.680 158.715 27.000 158.775 ;
        RECT 30.360 158.715 30.680 158.775 ;
        RECT 31.755 158.730 32.045 158.775 ;
        RECT 20.700 158.375 21.020 158.635 ;
        RECT 21.160 158.375 21.480 158.635 ;
        RECT 31.295 158.575 31.585 158.620 ;
        RECT 32.660 158.575 32.980 158.635 ;
        RECT 33.580 158.575 33.900 158.635 ;
        RECT 31.295 158.435 33.900 158.575 ;
        RECT 34.130 158.575 34.270 158.775 ;
        RECT 35.435 158.730 35.725 158.960 ;
        RECT 35.970 158.575 36.110 159.455 ;
        RECT 37.735 159.410 38.025 159.455 ;
        RECT 43.240 159.595 43.560 159.655 ;
        RECT 50.140 159.595 50.460 159.655 ;
        RECT 57.500 159.595 57.820 159.655 ;
        RECT 68.540 159.595 68.860 159.655 ;
        RECT 43.240 159.455 48.530 159.595 ;
        RECT 43.240 159.395 43.560 159.455 ;
        RECT 40.020 159.055 40.340 159.315 ;
        RECT 42.780 159.055 43.100 159.315 ;
        RECT 38.655 158.915 38.945 158.960 ;
        RECT 38.655 158.775 40.710 158.915 ;
        RECT 38.655 158.730 38.945 158.775 ;
        RECT 34.130 158.435 36.110 158.575 ;
        RECT 39.575 158.575 39.865 158.620 ;
        RECT 40.020 158.575 40.340 158.635 ;
        RECT 39.575 158.435 40.340 158.575 ;
        RECT 40.570 158.575 40.710 158.775 ;
        RECT 41.400 158.715 41.720 158.975 ;
        RECT 41.875 158.915 42.165 158.960 ;
        RECT 42.320 158.915 42.640 158.975 ;
        RECT 41.875 158.775 42.640 158.915 ;
        RECT 41.875 158.730 42.165 158.775 ;
        RECT 42.320 158.715 42.640 158.775 ;
        RECT 43.255 158.915 43.545 158.960 ;
        RECT 43.700 158.915 44.020 158.975 ;
        RECT 43.255 158.775 44.020 158.915 ;
        RECT 43.255 158.730 43.545 158.775 ;
        RECT 43.700 158.715 44.020 158.775 ;
        RECT 44.160 158.715 44.480 158.975 ;
        RECT 44.620 158.715 44.940 158.975 ;
        RECT 45.095 158.915 45.385 158.960 ;
        RECT 46.000 158.915 46.320 158.975 ;
        RECT 45.095 158.775 46.320 158.915 ;
        RECT 45.095 158.730 45.385 158.775 ;
        RECT 46.000 158.715 46.320 158.775 ;
        RECT 46.920 158.915 47.240 158.975 ;
        RECT 48.390 158.960 48.530 159.455 ;
        RECT 50.140 159.455 68.860 159.595 ;
        RECT 50.140 159.395 50.460 159.455 ;
        RECT 57.500 159.395 57.820 159.455 ;
        RECT 68.540 159.395 68.860 159.455 ;
        RECT 86.020 159.595 86.340 159.655 ;
        RECT 98.900 159.595 99.220 159.655 ;
        RECT 101.675 159.595 101.965 159.640 ;
        RECT 86.020 159.455 89.010 159.595 ;
        RECT 86.020 159.395 86.340 159.455 ;
        RECT 49.235 159.255 49.525 159.300 ;
        RECT 54.280 159.255 54.600 159.315 ;
        RECT 49.235 159.115 54.600 159.255 ;
        RECT 49.235 159.070 49.525 159.115 ;
        RECT 54.280 159.055 54.600 159.115 ;
        RECT 78.675 159.255 78.965 159.300 ;
        RECT 81.535 159.255 81.825 159.300 ;
        RECT 84.775 159.255 85.425 159.300 ;
        RECT 78.675 159.115 85.425 159.255 ;
        RECT 78.675 159.070 78.965 159.115 ;
        RECT 81.535 159.070 82.125 159.115 ;
        RECT 84.775 159.070 85.425 159.115 ;
        RECT 73.615 158.975 73.905 158.990 ;
        RECT 47.855 158.915 48.145 158.960 ;
        RECT 46.920 158.775 48.145 158.915 ;
        RECT 46.920 158.715 47.240 158.775 ;
        RECT 47.855 158.730 48.145 158.775 ;
        RECT 48.315 158.730 48.605 158.960 ;
        RECT 64.875 158.915 65.165 158.960 ;
        RECT 65.780 158.915 66.100 158.975 ;
        RECT 64.875 158.775 66.100 158.915 ;
        RECT 64.875 158.730 65.165 158.775 ;
        RECT 65.780 158.715 66.100 158.775 ;
        RECT 66.700 158.715 67.020 158.975 ;
        RECT 69.460 158.715 69.780 158.975 ;
        RECT 70.840 158.715 71.160 158.975 ;
        RECT 72.680 158.715 73.000 158.975 ;
        RECT 73.600 158.715 73.920 158.975 ;
        RECT 74.075 158.730 74.365 158.960 ;
        RECT 74.520 158.915 74.840 158.975 ;
        RECT 76.820 158.915 77.140 158.975 ;
        RECT 74.520 158.775 77.140 158.915 ;
        RECT 42.780 158.575 43.100 158.635 ;
        RECT 46.475 158.575 46.765 158.620 ;
        RECT 40.570 158.435 42.550 158.575 ;
        RECT 31.295 158.390 31.585 158.435 ;
        RECT 32.660 158.375 32.980 158.435 ;
        RECT 33.580 158.375 33.900 158.435 ;
        RECT 39.575 158.390 39.865 158.435 ;
        RECT 40.020 158.375 40.340 158.435 ;
        RECT 28.980 158.235 29.300 158.295 ;
        RECT 40.495 158.235 40.785 158.280 ;
        RECT 28.980 158.095 40.785 158.235 ;
        RECT 42.410 158.235 42.550 158.435 ;
        RECT 42.780 158.435 46.765 158.575 ;
        RECT 42.780 158.375 43.100 158.435 ;
        RECT 46.475 158.390 46.765 158.435 ;
        RECT 68.080 158.575 68.400 158.635 ;
        RECT 74.150 158.575 74.290 158.730 ;
        RECT 74.520 158.715 74.840 158.775 ;
        RECT 76.820 158.715 77.140 158.775 ;
        RECT 77.280 158.915 77.600 158.975 ;
        RECT 79.135 158.915 79.425 158.960 ;
        RECT 77.280 158.775 79.425 158.915 ;
        RECT 77.280 158.715 77.600 158.775 ;
        RECT 79.135 158.730 79.425 158.775 ;
        RECT 81.835 158.755 82.125 159.070 ;
        RECT 87.400 159.055 87.720 159.315 ;
        RECT 88.870 158.960 89.010 159.455 ;
        RECT 98.900 159.455 101.965 159.595 ;
        RECT 98.900 159.395 99.220 159.455 ;
        RECT 101.675 159.410 101.965 159.455 ;
        RECT 96.615 159.255 96.905 159.300 ;
        RECT 97.075 159.255 97.365 159.300 ;
        RECT 108.100 159.255 108.420 159.315 ;
        RECT 96.615 159.115 97.365 159.255 ;
        RECT 96.615 159.070 96.905 159.115 ;
        RECT 97.075 159.070 97.365 159.115 ;
        RECT 97.610 159.115 108.420 159.255 ;
        RECT 82.915 158.915 83.205 158.960 ;
        RECT 86.495 158.915 86.785 158.960 ;
        RECT 88.330 158.915 88.620 158.960 ;
        RECT 82.915 158.775 88.620 158.915 ;
        RECT 82.915 158.730 83.205 158.775 ;
        RECT 86.495 158.730 86.785 158.775 ;
        RECT 88.330 158.730 88.620 158.775 ;
        RECT 88.795 158.730 89.085 158.960 ;
        RECT 95.220 158.715 95.540 158.975 ;
        RECT 95.680 158.715 96.000 158.975 ;
        RECT 68.080 158.435 74.290 158.575 ;
        RECT 68.080 158.375 68.400 158.435 ;
        RECT 49.220 158.235 49.540 158.295 ;
        RECT 42.410 158.095 44.390 158.235 ;
        RECT 28.980 158.035 29.300 158.095 ;
        RECT 40.495 158.050 40.785 158.095 ;
        RECT 33.580 157.895 33.900 157.955 ;
        RECT 34.515 157.895 34.805 157.940 ;
        RECT 33.580 157.755 34.805 157.895 ;
        RECT 33.580 157.695 33.900 157.755 ;
        RECT 34.515 157.710 34.805 157.755 ;
        RECT 39.100 157.695 39.420 157.955 ;
        RECT 42.795 157.895 43.085 157.940 ;
        RECT 43.240 157.895 43.560 157.955 ;
        RECT 42.795 157.755 43.560 157.895 ;
        RECT 44.250 157.895 44.390 158.095 ;
        RECT 46.550 158.095 49.540 158.235 ;
        RECT 46.550 157.895 46.690 158.095 ;
        RECT 49.220 158.035 49.540 158.095 ;
        RECT 52.440 158.235 52.760 158.295 ;
        RECT 56.120 158.235 56.440 158.295 ;
        RECT 65.795 158.235 66.085 158.280 ;
        RECT 74.150 158.235 74.290 158.435 ;
        RECT 80.055 158.575 80.345 158.620 ;
        RECT 97.610 158.575 97.750 159.115 ;
        RECT 98.455 158.730 98.745 158.960 ;
        RECT 80.055 158.435 97.750 158.575 ;
        RECT 80.055 158.390 80.345 158.435 ;
        RECT 81.970 158.295 82.110 158.435 ;
        RECT 74.980 158.235 75.300 158.295 ;
        RECT 52.440 158.095 73.830 158.235 ;
        RECT 74.150 158.095 75.300 158.235 ;
        RECT 52.440 158.035 52.760 158.095 ;
        RECT 56.120 158.035 56.440 158.095 ;
        RECT 65.795 158.050 66.085 158.095 ;
        RECT 44.250 157.755 46.690 157.895 ;
        RECT 42.795 157.710 43.085 157.755 ;
        RECT 43.240 157.695 43.560 157.755 ;
        RECT 46.920 157.695 47.240 157.955 ;
        RECT 47.840 157.695 48.160 157.955 ;
        RECT 58.435 157.895 58.725 157.940 ;
        RECT 59.340 157.895 59.660 157.955 ;
        RECT 58.435 157.755 59.660 157.895 ;
        RECT 58.435 157.710 58.725 157.755 ;
        RECT 59.340 157.695 59.660 157.755 ;
        RECT 64.400 157.895 64.720 157.955 ;
        RECT 69.935 157.895 70.225 157.940 ;
        RECT 64.400 157.755 70.225 157.895 ;
        RECT 73.690 157.895 73.830 158.095 ;
        RECT 74.980 158.035 75.300 158.095 ;
        RECT 75.530 158.095 81.650 158.235 ;
        RECT 75.530 157.895 75.670 158.095 ;
        RECT 73.690 157.755 75.670 157.895 ;
        RECT 75.915 157.895 76.205 157.940 ;
        RECT 76.360 157.895 76.680 157.955 ;
        RECT 75.915 157.755 76.680 157.895 ;
        RECT 81.510 157.895 81.650 158.095 ;
        RECT 81.880 158.035 82.200 158.295 ;
        RECT 82.915 158.235 83.205 158.280 ;
        RECT 86.035 158.235 86.325 158.280 ;
        RECT 87.925 158.235 88.215 158.280 ;
        RECT 98.530 158.235 98.670 158.730 ;
        RECT 98.900 158.715 99.220 158.975 ;
        RECT 99.450 158.960 99.590 159.115 ;
        RECT 108.100 159.055 108.420 159.115 ;
        RECT 109.430 159.255 109.720 159.300 ;
        RECT 110.860 159.255 111.180 159.315 ;
        RECT 112.690 159.255 112.980 159.300 ;
        RECT 109.430 159.115 112.980 159.255 ;
        RECT 109.430 159.070 109.720 159.115 ;
        RECT 110.860 159.055 111.180 159.115 ;
        RECT 112.690 159.070 112.980 159.115 ;
        RECT 113.610 159.255 113.900 159.300 ;
        RECT 115.470 159.255 115.760 159.300 ;
        RECT 113.610 159.115 115.760 159.255 ;
        RECT 113.610 159.070 113.900 159.115 ;
        RECT 115.470 159.070 115.760 159.115 ;
        RECT 99.375 158.730 99.665 158.960 ;
        RECT 99.820 158.915 100.140 158.975 ;
        RECT 100.295 158.915 100.585 158.960 ;
        RECT 99.820 158.775 100.585 158.915 ;
        RECT 99.820 158.715 100.140 158.775 ;
        RECT 100.295 158.730 100.585 158.775 ;
        RECT 102.580 158.915 102.900 158.975 ;
        RECT 103.055 158.915 103.345 158.960 ;
        RECT 102.580 158.775 103.345 158.915 ;
        RECT 102.580 158.715 102.900 158.775 ;
        RECT 103.055 158.730 103.345 158.775 ;
        RECT 103.515 158.730 103.805 158.960 ;
        RECT 103.975 158.730 104.265 158.960 ;
        RECT 104.420 158.915 104.740 158.975 ;
        RECT 104.895 158.915 105.185 158.960 ;
        RECT 104.420 158.775 105.185 158.915 ;
        RECT 98.990 158.575 99.130 158.715 ;
        RECT 102.120 158.575 102.440 158.635 ;
        RECT 103.590 158.575 103.730 158.730 ;
        RECT 98.990 158.435 103.730 158.575 ;
        RECT 104.050 158.575 104.190 158.730 ;
        RECT 104.420 158.715 104.740 158.775 ;
        RECT 104.895 158.730 105.185 158.775 ;
        RECT 111.290 158.915 111.580 158.960 ;
        RECT 113.610 158.915 113.825 159.070 ;
        RECT 111.290 158.775 113.825 158.915 ;
        RECT 111.290 158.730 111.580 158.775 ;
        RECT 114.540 158.715 114.860 158.975 ;
        RECT 116.380 158.715 116.700 158.975 ;
        RECT 104.050 158.435 107.640 158.575 ;
        RECT 102.120 158.375 102.440 158.435 ;
        RECT 102.580 158.235 102.900 158.295 ;
        RECT 82.915 158.095 88.215 158.235 ;
        RECT 82.915 158.050 83.205 158.095 ;
        RECT 86.035 158.050 86.325 158.095 ;
        RECT 87.925 158.050 88.215 158.095 ;
        RECT 93.930 158.095 98.210 158.235 ;
        RECT 98.530 158.095 102.900 158.235 ;
        RECT 93.930 157.955 94.070 158.095 ;
        RECT 93.840 157.895 94.160 157.955 ;
        RECT 81.510 157.755 94.160 157.895 ;
        RECT 64.400 157.695 64.720 157.755 ;
        RECT 69.935 157.710 70.225 157.755 ;
        RECT 75.915 157.710 76.205 157.755 ;
        RECT 76.360 157.695 76.680 157.755 ;
        RECT 93.840 157.695 94.160 157.755 ;
        RECT 94.300 157.695 94.620 157.955 ;
        RECT 96.615 157.895 96.905 157.940 ;
        RECT 97.060 157.895 97.380 157.955 ;
        RECT 96.615 157.755 97.380 157.895 ;
        RECT 98.070 157.895 98.210 158.095 ;
        RECT 102.580 158.035 102.900 158.095 ;
        RECT 98.900 157.895 99.220 157.955 ;
        RECT 107.500 157.940 107.640 158.435 ;
        RECT 111.290 158.235 111.580 158.280 ;
        RECT 114.070 158.235 114.360 158.280 ;
        RECT 115.930 158.235 116.220 158.280 ;
        RECT 111.290 158.095 116.220 158.235 ;
        RECT 111.290 158.050 111.580 158.095 ;
        RECT 114.070 158.050 114.360 158.095 ;
        RECT 115.930 158.050 116.220 158.095 ;
        RECT 98.070 157.755 99.220 157.895 ;
        RECT 96.615 157.710 96.905 157.755 ;
        RECT 97.060 157.695 97.380 157.755 ;
        RECT 98.900 157.695 99.220 157.755 ;
        RECT 107.425 157.895 107.715 157.940 ;
        RECT 109.020 157.895 109.340 157.955 ;
        RECT 107.425 157.755 109.340 157.895 ;
        RECT 107.425 157.710 107.715 157.755 ;
        RECT 109.020 157.695 109.340 157.755 ;
        RECT 11.430 157.075 118.610 157.555 ;
        RECT 20.700 156.875 21.020 156.935 ;
        RECT 20.700 156.735 24.150 156.875 ;
        RECT 20.700 156.675 21.020 156.735 ;
        RECT 23.460 156.335 23.780 156.595 ;
        RECT 24.010 156.535 24.150 156.735 ;
        RECT 26.680 156.675 27.000 156.935 ;
        RECT 44.160 156.875 44.480 156.935 ;
        RECT 27.230 156.735 44.480 156.875 ;
        RECT 27.230 156.535 27.370 156.735 ;
        RECT 44.160 156.675 44.480 156.735 ;
        RECT 46.920 156.675 47.240 156.935 ;
        RECT 57.285 156.875 57.575 156.920 ;
        RECT 59.800 156.875 60.120 156.935 ;
        RECT 57.285 156.735 60.120 156.875 ;
        RECT 57.285 156.690 57.575 156.735 ;
        RECT 59.800 156.675 60.120 156.735 ;
        RECT 66.700 156.875 67.020 156.935 ;
        RECT 67.635 156.875 67.925 156.920 ;
        RECT 66.700 156.735 67.925 156.875 ;
        RECT 66.700 156.675 67.020 156.735 ;
        RECT 67.635 156.690 67.925 156.735 ;
        RECT 68.540 156.875 68.860 156.935 ;
        RECT 74.060 156.875 74.380 156.935 ;
        RECT 80.960 156.875 81.280 156.935 ;
        RECT 68.540 156.735 74.380 156.875 ;
        RECT 68.540 156.675 68.860 156.735 ;
        RECT 74.060 156.675 74.380 156.735 ;
        RECT 79.900 156.735 81.280 156.875 ;
        RECT 24.010 156.395 27.370 156.535 ;
        RECT 29.555 156.535 29.845 156.580 ;
        RECT 32.675 156.535 32.965 156.580 ;
        RECT 34.565 156.535 34.855 156.580 ;
        RECT 29.555 156.395 34.855 156.535 ;
        RECT 29.555 156.350 29.845 156.395 ;
        RECT 32.675 156.350 32.965 156.395 ;
        RECT 34.565 156.350 34.855 156.395 ;
        RECT 61.150 156.535 61.440 156.580 ;
        RECT 63.930 156.535 64.220 156.580 ;
        RECT 65.790 156.535 66.080 156.580 ;
        RECT 61.150 156.395 66.080 156.535 ;
        RECT 61.150 156.350 61.440 156.395 ;
        RECT 63.930 156.350 64.220 156.395 ;
        RECT 65.790 156.350 66.080 156.395 ;
        RECT 66.240 156.535 66.560 156.595 ;
        RECT 68.080 156.535 68.400 156.595 ;
        RECT 71.775 156.535 72.065 156.580 ;
        RECT 79.900 156.535 80.040 156.735 ;
        RECT 80.960 156.675 81.280 156.735 ;
        RECT 84.195 156.875 84.485 156.920 ;
        RECT 84.640 156.875 84.960 156.935 ;
        RECT 84.195 156.735 84.960 156.875 ;
        RECT 84.195 156.690 84.485 156.735 ;
        RECT 84.640 156.675 84.960 156.735 ;
        RECT 98.440 156.675 98.760 156.935 ;
        RECT 110.875 156.875 111.165 156.920 ;
        RECT 112.700 156.875 113.020 156.935 ;
        RECT 110.875 156.735 113.020 156.875 ;
        RECT 110.875 156.690 111.165 156.735 ;
        RECT 112.700 156.675 113.020 156.735 ;
        RECT 66.240 156.395 68.770 156.535 ;
        RECT 66.240 156.335 66.560 156.395 ;
        RECT 68.080 156.335 68.400 156.395 ;
        RECT 23.550 156.195 23.690 156.335 ;
        RECT 33.580 156.195 33.900 156.255 ;
        RECT 34.055 156.195 34.345 156.240 ;
        RECT 18.490 156.055 25.530 156.195 ;
        RECT 18.490 155.900 18.630 156.055 ;
        RECT 18.415 155.670 18.705 155.900 ;
        RECT 21.620 155.855 21.940 155.915 ;
        RECT 25.390 155.900 25.530 156.055 ;
        RECT 33.580 156.055 34.345 156.195 ;
        RECT 33.580 155.995 33.900 156.055 ;
        RECT 34.055 156.010 34.345 156.055 ;
        RECT 46.460 155.995 46.780 156.255 ;
        RECT 48.300 156.195 48.620 156.255 ;
        RECT 50.155 156.195 50.445 156.240 ;
        RECT 56.120 156.195 56.440 156.255 ;
        RECT 48.300 156.055 50.445 156.195 ;
        RECT 48.300 155.995 48.620 156.055 ;
        RECT 50.155 156.010 50.445 156.055 ;
        RECT 55.290 156.055 56.440 156.195 ;
        RECT 23.475 155.855 23.765 155.900 ;
        RECT 21.620 155.715 23.765 155.855 ;
        RECT 21.620 155.655 21.940 155.715 ;
        RECT 23.475 155.670 23.765 155.715 ;
        RECT 25.315 155.670 25.605 155.900 ;
        RECT 28.475 155.560 28.765 155.875 ;
        RECT 29.555 155.855 29.845 155.900 ;
        RECT 33.135 155.855 33.425 155.900 ;
        RECT 34.970 155.855 35.260 155.900 ;
        RECT 29.555 155.715 35.260 155.855 ;
        RECT 29.555 155.670 29.845 155.715 ;
        RECT 33.135 155.670 33.425 155.715 ;
        RECT 34.970 155.670 35.260 155.715 ;
        RECT 35.420 155.655 35.740 155.915 ;
        RECT 45.540 155.655 45.860 155.915 ;
        RECT 48.775 155.855 49.065 155.900 ;
        RECT 49.220 155.855 49.540 155.915 ;
        RECT 48.775 155.715 49.540 155.855 ;
        RECT 48.775 155.670 49.065 155.715 ;
        RECT 49.220 155.655 49.540 155.715 ;
        RECT 49.680 155.855 50.000 155.915 ;
        RECT 51.075 155.855 51.365 155.900 ;
        RECT 49.680 155.715 51.365 155.855 ;
        RECT 49.680 155.655 50.000 155.715 ;
        RECT 51.075 155.670 51.365 155.715 ;
        RECT 54.740 155.655 55.060 155.915 ;
        RECT 55.290 155.900 55.430 156.055 ;
        RECT 56.120 155.995 56.440 156.055 ;
        RECT 64.400 155.995 64.720 156.255 ;
        RECT 68.630 156.240 68.770 156.395 ;
        RECT 71.775 156.395 80.040 156.535 ;
        RECT 94.300 156.535 94.620 156.595 ;
        RECT 111.780 156.535 112.100 156.595 ;
        RECT 94.300 156.395 112.100 156.535 ;
        RECT 71.775 156.350 72.065 156.395 ;
        RECT 94.300 156.335 94.620 156.395 ;
        RECT 111.780 156.335 112.100 156.395 ;
        RECT 65.870 156.055 67.390 156.195 ;
        RECT 55.215 155.670 55.505 155.900 ;
        RECT 55.660 155.655 55.980 155.915 ;
        RECT 56.595 155.855 56.885 155.900 ;
        RECT 57.500 155.855 57.820 155.915 ;
        RECT 56.595 155.715 57.820 155.855 ;
        RECT 56.595 155.670 56.885 155.715 ;
        RECT 57.500 155.655 57.820 155.715 ;
        RECT 61.150 155.855 61.440 155.900 ;
        RECT 61.150 155.715 63.685 155.855 ;
        RECT 61.150 155.670 61.440 155.715 ;
        RECT 62.560 155.560 62.880 155.575 ;
        RECT 25.775 155.515 26.065 155.560 ;
        RECT 28.175 155.515 28.765 155.560 ;
        RECT 31.415 155.515 32.065 155.560 ;
        RECT 25.775 155.375 32.065 155.515 ;
        RECT 25.775 155.330 26.065 155.375 ;
        RECT 28.175 155.330 28.465 155.375 ;
        RECT 31.415 155.330 32.065 155.375 ;
        RECT 46.935 155.515 47.225 155.560 ;
        RECT 53.375 155.515 53.665 155.560 ;
        RECT 46.935 155.375 53.665 155.515 ;
        RECT 46.935 155.330 47.225 155.375 ;
        RECT 53.375 155.330 53.665 155.375 ;
        RECT 59.290 155.515 59.580 155.560 ;
        RECT 62.550 155.515 62.880 155.560 ;
        RECT 59.290 155.375 62.880 155.515 ;
        RECT 59.290 155.330 59.580 155.375 ;
        RECT 62.550 155.330 62.880 155.375 ;
        RECT 63.470 155.560 63.685 155.715 ;
        RECT 63.470 155.515 63.760 155.560 ;
        RECT 65.330 155.515 65.620 155.560 ;
        RECT 63.470 155.375 65.620 155.515 ;
        RECT 63.470 155.330 63.760 155.375 ;
        RECT 65.330 155.330 65.620 155.375 ;
        RECT 62.560 155.315 62.880 155.330 ;
        RECT 17.940 154.975 18.260 155.235 ;
        RECT 20.700 155.175 21.020 155.235 ;
        RECT 22.555 155.175 22.845 155.220 ;
        RECT 20.700 155.035 22.845 155.175 ;
        RECT 20.700 154.975 21.020 155.035 ;
        RECT 22.555 154.990 22.845 155.035 ;
        RECT 44.620 154.975 44.940 155.235 ;
        RECT 48.315 155.175 48.605 155.220 ;
        RECT 48.760 155.175 49.080 155.235 ;
        RECT 48.315 155.035 49.080 155.175 ;
        RECT 48.315 154.990 48.605 155.035 ;
        RECT 48.760 154.975 49.080 155.035 ;
        RECT 50.140 155.175 50.460 155.235 ;
        RECT 50.615 155.175 50.905 155.220 ;
        RECT 50.140 155.035 50.905 155.175 ;
        RECT 50.140 154.975 50.460 155.035 ;
        RECT 50.615 154.990 50.905 155.035 ;
        RECT 52.915 155.175 53.205 155.220 ;
        RECT 55.200 155.175 55.520 155.235 ;
        RECT 52.915 155.035 55.520 155.175 ;
        RECT 52.915 154.990 53.205 155.035 ;
        RECT 55.200 154.975 55.520 155.035 ;
        RECT 62.100 155.175 62.420 155.235 ;
        RECT 65.870 155.175 66.010 156.055 ;
        RECT 67.250 155.900 67.390 156.055 ;
        RECT 68.555 156.010 68.845 156.240 ;
        RECT 69.015 156.195 69.305 156.240 ;
        RECT 69.460 156.195 69.780 156.255 ;
        RECT 75.900 156.195 76.220 156.255 ;
        RECT 69.015 156.055 69.780 156.195 ;
        RECT 69.015 156.010 69.305 156.055 ;
        RECT 69.460 155.995 69.780 156.055 ;
        RECT 73.690 156.055 76.220 156.195 ;
        RECT 66.255 155.670 66.545 155.900 ;
        RECT 67.175 155.670 67.465 155.900 ;
        RECT 66.330 155.515 66.470 155.670 ;
        RECT 70.380 155.655 70.700 155.915 ;
        RECT 70.840 155.855 71.160 155.915 ;
        RECT 72.680 155.855 73.000 155.915 ;
        RECT 73.690 155.900 73.830 156.055 ;
        RECT 75.900 155.995 76.220 156.055 ;
        RECT 80.960 155.995 81.280 156.255 ;
        RECT 81.880 155.995 82.200 156.255 ;
        RECT 93.380 156.195 93.700 156.255 ;
        RECT 97.995 156.195 98.285 156.240 ;
        RECT 93.380 156.055 98.285 156.195 ;
        RECT 93.380 155.995 93.700 156.055 ;
        RECT 97.995 156.010 98.285 156.055 ;
        RECT 99.820 156.195 100.140 156.255 ;
        RECT 103.960 156.195 104.280 156.255 ;
        RECT 99.820 156.055 104.650 156.195 ;
        RECT 99.820 155.995 100.140 156.055 ;
        RECT 103.960 155.995 104.280 156.055 ;
        RECT 70.840 155.715 73.000 155.855 ;
        RECT 70.840 155.655 71.160 155.715 ;
        RECT 72.680 155.655 73.000 155.715 ;
        RECT 73.615 155.670 73.905 155.900 ;
        RECT 74.060 155.855 74.380 155.915 ;
        RECT 74.765 155.855 75.055 155.900 ;
        RECT 76.820 155.855 77.140 155.915 ;
        RECT 74.060 155.715 74.575 155.855 ;
        RECT 74.765 155.715 77.140 155.855 ;
        RECT 74.060 155.655 74.380 155.715 ;
        RECT 74.765 155.670 75.055 155.715 ;
        RECT 76.820 155.655 77.140 155.715 ;
        RECT 97.520 155.655 97.840 155.915 ;
        RECT 102.580 155.655 102.900 155.915 ;
        RECT 104.510 155.900 104.650 156.055 ;
        RECT 107.640 155.995 107.960 156.255 ;
        RECT 103.055 155.670 103.345 155.900 ;
        RECT 103.515 155.670 103.805 155.900 ;
        RECT 104.435 155.670 104.725 155.900 ;
        RECT 107.180 155.855 107.500 155.915 ;
        RECT 109.035 155.855 109.325 155.900 ;
        RECT 107.180 155.715 109.325 155.855 ;
        RECT 66.330 155.375 73.830 155.515 ;
        RECT 62.100 155.035 66.010 155.175 ;
        RECT 69.000 155.175 69.320 155.235 ;
        RECT 70.380 155.175 70.700 155.235 ;
        RECT 69.000 155.035 70.700 155.175 ;
        RECT 73.690 155.175 73.830 155.375 ;
        RECT 98.900 155.315 99.220 155.575 ;
        RECT 102.120 155.515 102.440 155.575 ;
        RECT 103.130 155.515 103.270 155.670 ;
        RECT 102.120 155.375 103.270 155.515 ;
        RECT 103.590 155.515 103.730 155.670 ;
        RECT 107.180 155.655 107.500 155.715 ;
        RECT 109.035 155.670 109.325 155.715 ;
        RECT 108.100 155.515 108.420 155.575 ;
        RECT 103.590 155.375 108.420 155.515 ;
        RECT 102.120 155.315 102.440 155.375 ;
        RECT 108.100 155.315 108.420 155.375 ;
        RECT 74.980 155.175 75.300 155.235 ;
        RECT 73.690 155.035 75.300 155.175 ;
        RECT 62.100 154.975 62.420 155.035 ;
        RECT 69.000 154.975 69.320 155.035 ;
        RECT 70.380 154.975 70.700 155.035 ;
        RECT 74.980 154.975 75.300 155.035 ;
        RECT 75.900 154.975 76.220 155.235 ;
        RECT 81.880 155.175 82.200 155.235 ;
        RECT 82.355 155.175 82.645 155.220 ;
        RECT 81.880 155.035 82.645 155.175 ;
        RECT 81.880 154.975 82.200 155.035 ;
        RECT 82.355 154.990 82.645 155.035 ;
        RECT 95.680 155.175 96.000 155.235 ;
        RECT 96.615 155.175 96.905 155.220 ;
        RECT 95.680 155.035 96.905 155.175 ;
        RECT 95.680 154.975 96.000 155.035 ;
        RECT 96.615 154.990 96.905 155.035 ;
        RECT 99.360 155.175 99.680 155.235 ;
        RECT 101.215 155.175 101.505 155.220 ;
        RECT 99.360 155.035 101.505 155.175 ;
        RECT 99.360 154.975 99.680 155.035 ;
        RECT 101.215 154.990 101.505 155.035 ;
        RECT 108.575 155.175 108.865 155.220 ;
        RECT 109.020 155.175 109.340 155.235 ;
        RECT 108.575 155.035 109.340 155.175 ;
        RECT 108.575 154.990 108.865 155.035 ;
        RECT 109.020 154.975 109.340 155.035 ;
        RECT 10.650 154.355 118.610 154.835 ;
        RECT 36.800 153.955 37.120 154.215 ;
        RECT 38.180 154.155 38.500 154.215 ;
        RECT 53.360 154.155 53.680 154.215 ;
        RECT 65.780 154.155 66.100 154.215 ;
        RECT 67.175 154.155 67.465 154.200 ;
        RECT 38.180 154.015 39.330 154.155 ;
        RECT 38.180 153.955 38.500 154.015 ;
        RECT 17.940 153.860 18.260 153.875 ;
        RECT 14.835 153.815 15.125 153.860 ;
        RECT 17.940 153.815 18.725 153.860 ;
        RECT 14.835 153.675 18.725 153.815 ;
        RECT 14.835 153.630 15.425 153.675 ;
        RECT 15.135 153.315 15.425 153.630 ;
        RECT 17.940 153.630 18.725 153.675 ;
        RECT 17.940 153.615 18.260 153.630 ;
        RECT 20.700 153.615 21.020 153.875 ;
        RECT 26.220 153.815 26.540 153.875 ;
        RECT 32.200 153.815 32.520 153.875 ;
        RECT 35.420 153.815 35.740 153.875 ;
        RECT 22.170 153.675 35.740 153.815 ;
        RECT 36.890 153.815 37.030 153.955 ;
        RECT 39.190 153.815 39.330 154.015 ;
        RECT 53.360 154.015 65.090 154.155 ;
        RECT 53.360 153.955 53.680 154.015 ;
        RECT 46.410 153.815 46.700 153.860 ;
        RECT 48.760 153.815 49.080 153.875 ;
        RECT 49.670 153.815 49.960 153.860 ;
        RECT 36.890 153.675 37.950 153.815 ;
        RECT 22.170 153.520 22.310 153.675 ;
        RECT 26.220 153.615 26.540 153.675 ;
        RECT 32.200 153.615 32.520 153.675 ;
        RECT 35.420 153.615 35.740 153.675 ;
        RECT 37.810 153.535 37.950 153.675 ;
        RECT 39.190 153.675 43.930 153.815 ;
        RECT 16.215 153.475 16.505 153.520 ;
        RECT 19.795 153.475 20.085 153.520 ;
        RECT 21.630 153.475 21.920 153.520 ;
        RECT 16.215 153.335 21.920 153.475 ;
        RECT 16.215 153.290 16.505 153.335 ;
        RECT 19.795 153.290 20.085 153.335 ;
        RECT 21.630 153.290 21.920 153.335 ;
        RECT 22.095 153.290 22.385 153.520 ;
        RECT 30.360 153.275 30.680 153.535 ;
        RECT 35.880 153.475 36.200 153.535 ;
        RECT 36.800 153.475 37.120 153.535 ;
        RECT 37.275 153.475 37.565 153.520 ;
        RECT 35.880 153.335 37.565 153.475 ;
        RECT 35.880 153.275 36.200 153.335 ;
        RECT 36.800 153.275 37.120 153.335 ;
        RECT 37.275 153.290 37.565 153.335 ;
        RECT 37.720 153.275 38.040 153.535 ;
        RECT 39.190 153.520 39.330 153.675 ;
        RECT 43.790 153.535 43.930 153.675 ;
        RECT 46.410 153.675 49.960 153.815 ;
        RECT 46.410 153.630 46.700 153.675 ;
        RECT 48.760 153.615 49.080 153.675 ;
        RECT 49.670 153.630 49.960 153.675 ;
        RECT 50.590 153.815 50.880 153.860 ;
        RECT 52.450 153.815 52.740 153.860 ;
        RECT 50.590 153.675 52.740 153.815 ;
        RECT 50.590 153.630 50.880 153.675 ;
        RECT 52.450 153.630 52.740 153.675 ;
        RECT 38.195 153.290 38.485 153.520 ;
        RECT 39.115 153.290 39.405 153.520 ;
        RECT 39.575 153.475 39.865 153.520 ;
        RECT 40.020 153.475 40.340 153.535 ;
        RECT 39.575 153.335 40.340 153.475 ;
        RECT 39.575 153.290 39.865 153.335 ;
        RECT 13.355 153.135 13.645 153.180 ;
        RECT 20.240 153.135 20.560 153.195 ;
        RECT 13.355 152.995 20.560 153.135 ;
        RECT 13.355 152.950 13.645 152.995 ;
        RECT 20.240 152.935 20.560 152.995 ;
        RECT 23.015 153.135 23.305 153.180 ;
        RECT 30.820 153.135 31.140 153.195 ;
        RECT 23.015 152.995 31.140 153.135 ;
        RECT 23.015 152.950 23.305 152.995 ;
        RECT 30.820 152.935 31.140 152.995 ;
        RECT 31.295 153.135 31.585 153.180 ;
        RECT 33.120 153.135 33.440 153.195 ;
        RECT 31.295 152.995 33.440 153.135 ;
        RECT 31.295 152.950 31.585 152.995 ;
        RECT 33.120 152.935 33.440 152.995 ;
        RECT 16.215 152.795 16.505 152.840 ;
        RECT 19.335 152.795 19.625 152.840 ;
        RECT 21.225 152.795 21.515 152.840 ;
        RECT 16.215 152.655 21.515 152.795 ;
        RECT 16.215 152.610 16.505 152.655 ;
        RECT 19.335 152.610 19.625 152.655 ;
        RECT 21.225 152.610 21.515 152.655 ;
        RECT 22.540 152.795 22.860 152.855 ;
        RECT 38.270 152.795 38.410 153.290 ;
        RECT 40.020 153.275 40.340 153.335 ;
        RECT 43.700 153.475 44.020 153.535 ;
        RECT 48.270 153.475 48.560 153.520 ;
        RECT 50.590 153.475 50.805 153.630 ;
        RECT 52.900 153.475 53.220 153.535 ;
        RECT 43.700 153.335 45.310 153.475 ;
        RECT 43.700 153.275 44.020 153.335 ;
        RECT 40.940 152.935 41.260 153.195 ;
        RECT 42.320 153.135 42.640 153.195 ;
        RECT 44.620 153.135 44.940 153.195 ;
        RECT 42.320 152.995 44.940 153.135 ;
        RECT 45.170 153.135 45.310 153.335 ;
        RECT 48.270 153.335 50.805 153.475 ;
        RECT 51.150 153.335 53.220 153.475 ;
        RECT 48.270 153.290 48.560 153.335 ;
        RECT 51.150 153.135 51.290 153.335 ;
        RECT 52.900 153.275 53.220 153.335 ;
        RECT 53.375 153.475 53.665 153.520 ;
        RECT 53.820 153.475 54.140 153.535 ;
        RECT 53.375 153.335 54.140 153.475 ;
        RECT 53.375 153.290 53.665 153.335 ;
        RECT 53.820 153.275 54.140 153.335 ;
        RECT 55.200 153.275 55.520 153.535 ;
        RECT 59.295 153.490 59.585 153.520 ;
        RECT 59.295 153.475 60.030 153.490 ;
        RECT 61.195 153.475 61.485 153.520 ;
        RECT 62.100 153.475 62.420 153.535 ;
        RECT 59.295 153.350 62.420 153.475 ;
        RECT 59.295 153.290 59.585 153.350 ;
        RECT 59.890 153.335 62.420 153.350 ;
        RECT 61.195 153.290 61.485 153.335 ;
        RECT 62.100 153.275 62.420 153.335 ;
        RECT 45.170 152.995 51.290 153.135 ;
        RECT 51.535 153.135 51.825 153.180 ;
        RECT 60.260 153.135 60.580 153.195 ;
        RECT 63.955 153.135 64.245 153.180 ;
        RECT 51.535 152.995 54.510 153.135 ;
        RECT 42.320 152.935 42.640 152.995 ;
        RECT 44.620 152.935 44.940 152.995 ;
        RECT 51.535 152.950 51.825 152.995 ;
        RECT 54.370 152.840 54.510 152.995 ;
        RECT 60.260 152.995 64.245 153.135 ;
        RECT 60.260 152.935 60.580 152.995 ;
        RECT 63.955 152.950 64.245 152.995 ;
        RECT 22.540 152.655 38.410 152.795 ;
        RECT 48.270 152.795 48.560 152.840 ;
        RECT 51.050 152.795 51.340 152.840 ;
        RECT 52.910 152.795 53.200 152.840 ;
        RECT 48.270 152.655 53.200 152.795 ;
        RECT 22.540 152.595 22.860 152.655 ;
        RECT 48.270 152.610 48.560 152.655 ;
        RECT 51.050 152.610 51.340 152.655 ;
        RECT 52.910 152.610 53.200 152.655 ;
        RECT 54.295 152.610 54.585 152.840 ;
        RECT 64.950 152.795 65.090 154.015 ;
        RECT 65.780 154.015 67.465 154.155 ;
        RECT 65.780 153.955 66.100 154.015 ;
        RECT 67.175 153.970 67.465 154.015 ;
        RECT 70.855 154.155 71.145 154.200 ;
        RECT 73.140 154.155 73.460 154.215 ;
        RECT 70.855 154.015 72.450 154.155 ;
        RECT 70.855 153.970 71.145 154.015 ;
        RECT 65.335 153.815 65.625 153.860 ;
        RECT 69.000 153.815 69.320 153.875 ;
        RECT 65.335 153.675 69.320 153.815 ;
        RECT 65.335 153.630 65.625 153.675 ;
        RECT 69.000 153.615 69.320 153.675 ;
        RECT 66.255 153.475 66.545 153.520 ;
        RECT 67.160 153.475 67.480 153.535 ;
        RECT 66.255 153.335 67.480 153.475 ;
        RECT 66.255 153.290 66.545 153.335 ;
        RECT 67.160 153.275 67.480 153.335 ;
        RECT 68.095 153.475 68.385 153.520 ;
        RECT 69.460 153.475 69.780 153.535 ;
        RECT 69.935 153.475 70.225 153.520 ;
        RECT 68.095 153.335 70.225 153.475 ;
        RECT 68.095 153.290 68.385 153.335 ;
        RECT 69.460 153.275 69.780 153.335 ;
        RECT 69.935 153.290 70.225 153.335 ;
        RECT 71.775 153.290 72.065 153.520 ;
        RECT 70.840 153.135 71.160 153.195 ;
        RECT 71.850 153.135 71.990 153.290 ;
        RECT 69.090 152.995 71.990 153.135 ;
        RECT 72.310 153.135 72.450 154.015 ;
        RECT 72.770 154.015 73.460 154.155 ;
        RECT 72.770 153.520 72.910 154.015 ;
        RECT 73.140 153.955 73.460 154.015 ;
        RECT 74.060 154.155 74.380 154.215 ;
        RECT 75.900 154.155 76.220 154.215 ;
        RECT 74.060 154.015 76.220 154.155 ;
        RECT 74.060 153.955 74.380 154.015 ;
        RECT 75.900 153.955 76.220 154.015 ;
        RECT 80.285 154.155 80.575 154.200 ;
        RECT 81.420 154.155 81.740 154.215 ;
        RECT 80.285 154.015 81.740 154.155 ;
        RECT 80.285 153.970 80.575 154.015 ;
        RECT 81.420 153.955 81.740 154.015 ;
        RECT 81.970 154.015 89.470 154.155 ;
        RECT 74.520 153.815 74.840 153.875 ;
        RECT 73.230 153.675 74.840 153.815 ;
        RECT 73.230 153.535 73.370 153.675 ;
        RECT 74.520 153.615 74.840 153.675 ;
        RECT 74.980 153.815 75.300 153.875 ;
        RECT 81.970 153.815 82.110 154.015 ;
        RECT 85.560 153.860 85.880 153.875 ;
        RECT 74.980 153.675 82.110 153.815 ;
        RECT 82.290 153.815 82.580 153.860 ;
        RECT 85.550 153.815 85.880 153.860 ;
        RECT 82.290 153.675 85.880 153.815 ;
        RECT 74.980 153.615 75.300 153.675 ;
        RECT 82.290 153.630 82.580 153.675 ;
        RECT 85.550 153.630 85.880 153.675 ;
        RECT 85.560 153.615 85.880 153.630 ;
        RECT 86.470 153.815 86.760 153.860 ;
        RECT 88.330 153.815 88.620 153.860 ;
        RECT 86.470 153.675 88.620 153.815 ;
        RECT 86.470 153.630 86.760 153.675 ;
        RECT 88.330 153.630 88.620 153.675 ;
        RECT 72.695 153.290 72.985 153.520 ;
        RECT 73.140 153.275 73.460 153.535 ;
        RECT 73.600 153.475 73.920 153.535 ;
        RECT 76.820 153.475 77.140 153.535 ;
        RECT 73.600 153.335 77.140 153.475 ;
        RECT 73.600 153.275 73.920 153.335 ;
        RECT 76.820 153.275 77.140 153.335 ;
        RECT 84.150 153.475 84.440 153.520 ;
        RECT 86.470 153.475 86.685 153.630 ;
        RECT 89.330 153.535 89.470 154.015 ;
        RECT 98.900 153.955 99.220 154.215 ;
        RECT 102.120 154.155 102.440 154.215 ;
        RECT 100.830 154.015 102.440 154.155 ;
        RECT 92.475 153.815 92.765 153.860 ;
        RECT 92.935 153.815 93.225 153.860 ;
        RECT 92.475 153.675 93.225 153.815 ;
        RECT 92.475 153.630 92.765 153.675 ;
        RECT 92.935 153.630 93.225 153.675 ;
        RECT 93.840 153.815 94.160 153.875 ;
        RECT 100.830 153.815 100.970 154.015 ;
        RECT 102.120 153.955 102.440 154.015 ;
        RECT 108.100 154.155 108.420 154.215 ;
        RECT 108.575 154.155 108.865 154.200 ;
        RECT 108.100 154.015 108.865 154.155 ;
        RECT 108.100 153.955 108.420 154.015 ;
        RECT 108.575 153.970 108.865 154.015 ;
        RECT 109.020 153.955 109.340 154.215 ;
        RECT 93.840 153.675 100.970 153.815 ;
        RECT 93.840 153.615 94.160 153.675 ;
        RECT 84.150 153.335 86.685 153.475 ;
        RECT 84.150 153.290 84.440 153.335 ;
        RECT 89.240 153.275 89.560 153.535 ;
        RECT 89.700 153.475 90.020 153.535 ;
        RECT 94.850 153.520 94.990 153.675 ;
        RECT 91.095 153.475 91.385 153.520 ;
        RECT 94.315 153.475 94.605 153.520 ;
        RECT 89.700 153.335 91.385 153.475 ;
        RECT 89.700 153.275 90.020 153.335 ;
        RECT 91.095 153.290 91.385 153.335 ;
        RECT 93.930 153.335 94.605 153.475 ;
        RECT 77.280 153.135 77.600 153.195 ;
        RECT 72.310 152.995 77.600 153.135 ;
        RECT 69.090 152.840 69.230 152.995 ;
        RECT 70.840 152.935 71.160 152.995 ;
        RECT 77.280 152.935 77.600 152.995 ;
        RECT 87.400 152.935 87.720 153.195 ;
        RECT 92.015 153.135 92.305 153.180 ;
        RECT 92.920 153.135 93.240 153.195 ;
        RECT 92.015 152.995 93.240 153.135 ;
        RECT 92.015 152.950 92.305 152.995 ;
        RECT 92.920 152.935 93.240 152.995 ;
        RECT 69.015 152.795 69.305 152.840 ;
        RECT 84.150 152.795 84.440 152.840 ;
        RECT 86.930 152.795 87.220 152.840 ;
        RECT 88.790 152.795 89.080 152.840 ;
        RECT 93.930 152.795 94.070 153.335 ;
        RECT 94.315 153.290 94.605 153.335 ;
        RECT 94.775 153.290 95.065 153.520 ;
        RECT 95.235 153.290 95.525 153.520 ;
        RECT 96.140 153.475 96.460 153.535 ;
        RECT 98.900 153.475 99.220 153.535 ;
        RECT 100.830 153.520 100.970 153.675 ;
        RECT 100.295 153.475 100.585 153.520 ;
        RECT 96.140 153.335 98.670 153.475 ;
        RECT 95.310 153.135 95.450 153.290 ;
        RECT 96.140 153.275 96.460 153.335 ;
        RECT 98.530 153.135 98.670 153.335 ;
        RECT 98.900 153.335 100.585 153.475 ;
        RECT 98.900 153.275 99.220 153.335 ;
        RECT 100.295 153.290 100.585 153.335 ;
        RECT 100.755 153.290 101.045 153.520 ;
        RECT 101.215 153.475 101.505 153.520 ;
        RECT 101.660 153.475 101.980 153.535 ;
        RECT 101.215 153.335 101.980 153.475 ;
        RECT 101.215 153.290 101.505 153.335 ;
        RECT 101.660 153.275 101.980 153.335 ;
        RECT 102.135 153.290 102.425 153.520 ;
        RECT 99.820 153.135 100.140 153.195 ;
        RECT 102.210 153.135 102.350 153.290 ;
        RECT 113.620 153.275 113.940 153.535 ;
        RECT 95.310 152.995 96.370 153.135 ;
        RECT 98.530 152.995 102.350 153.135 ;
        RECT 96.230 152.855 96.370 152.995 ;
        RECT 99.820 152.935 100.140 152.995 ;
        RECT 107.640 152.935 107.960 153.195 ;
        RECT 109.480 153.135 109.800 153.195 ;
        RECT 112.255 153.135 112.545 153.180 ;
        RECT 109.480 152.995 112.545 153.135 ;
        RECT 109.480 152.935 109.800 152.995 ;
        RECT 112.255 152.950 112.545 152.995 ;
        RECT 64.950 152.655 69.305 152.795 ;
        RECT 69.015 152.610 69.305 152.655 ;
        RECT 73.000 152.655 83.950 152.795 ;
        RECT 25.760 152.255 26.080 152.515 ;
        RECT 28.535 152.455 28.825 152.500 ;
        RECT 29.900 152.455 30.220 152.515 ;
        RECT 28.535 152.315 30.220 152.455 ;
        RECT 28.535 152.270 28.825 152.315 ;
        RECT 29.900 152.255 30.220 152.315 ;
        RECT 35.880 152.255 36.200 152.515 ;
        RECT 44.620 152.500 44.940 152.515 ;
        RECT 44.405 152.270 44.940 152.500 ;
        RECT 44.620 152.255 44.940 152.270 ;
        RECT 45.540 152.455 45.860 152.515 ;
        RECT 60.275 152.455 60.565 152.500 ;
        RECT 61.180 152.455 61.500 152.515 ;
        RECT 45.540 152.315 61.500 152.455 ;
        RECT 45.540 152.255 45.860 152.315 ;
        RECT 60.275 152.270 60.565 152.315 ;
        RECT 61.180 152.255 61.500 152.315 ;
        RECT 62.100 152.455 62.420 152.515 ;
        RECT 73.000 152.455 73.140 152.655 ;
        RECT 62.100 152.315 73.140 152.455 ;
        RECT 62.100 152.255 62.420 152.315 ;
        RECT 74.980 152.255 75.300 152.515 ;
        RECT 83.810 152.455 83.950 152.655 ;
        RECT 84.150 152.655 89.080 152.795 ;
        RECT 84.150 152.610 84.440 152.655 ;
        RECT 86.930 152.610 87.220 152.655 ;
        RECT 88.790 152.610 89.080 152.655 ;
        RECT 89.790 152.655 94.070 152.795 ;
        RECT 89.790 152.455 89.930 152.655 ;
        RECT 83.810 152.315 89.930 152.455 ;
        RECT 90.160 152.255 90.480 152.515 ;
        RECT 90.620 152.455 90.940 152.515 ;
        RECT 91.095 152.455 91.385 152.500 ;
        RECT 90.620 152.315 91.385 152.455 ;
        RECT 93.930 152.455 94.070 152.655 ;
        RECT 96.140 152.595 96.460 152.855 ;
        RECT 98.900 152.455 99.220 152.515 ;
        RECT 102.580 152.455 102.900 152.515 ;
        RECT 93.930 152.315 102.900 152.455 ;
        RECT 90.620 152.255 90.940 152.315 ;
        RECT 91.095 152.270 91.385 152.315 ;
        RECT 98.900 152.255 99.220 152.315 ;
        RECT 102.580 152.255 102.900 152.315 ;
        RECT 110.875 152.455 111.165 152.500 ;
        RECT 116.840 152.455 117.160 152.515 ;
        RECT 110.875 152.315 117.160 152.455 ;
        RECT 110.875 152.270 111.165 152.315 ;
        RECT 116.840 152.255 117.160 152.315 ;
        RECT 11.430 151.635 118.610 152.115 ;
        RECT 21.620 151.235 21.940 151.495 ;
        RECT 30.360 151.435 30.680 151.495 ;
        RECT 37.260 151.435 37.580 151.495 ;
        RECT 46.460 151.435 46.780 151.495 ;
        RECT 62.560 151.435 62.880 151.495 ;
        RECT 63.495 151.435 63.785 151.480 ;
        RECT 30.360 151.295 37.580 151.435 ;
        RECT 30.360 151.235 30.680 151.295 ;
        RECT 37.260 151.235 37.580 151.295 ;
        RECT 46.090 151.295 59.340 151.435 ;
        RECT 21.160 151.095 21.480 151.155 ;
        RECT 24.380 151.095 24.700 151.155 ;
        RECT 18.950 150.955 24.700 151.095 ;
        RECT 18.950 150.800 19.090 150.955 ;
        RECT 21.160 150.895 21.480 150.955 ;
        RECT 24.380 150.895 24.700 150.955 ;
        RECT 26.335 151.095 26.625 151.140 ;
        RECT 29.455 151.095 29.745 151.140 ;
        RECT 31.345 151.095 31.635 151.140 ;
        RECT 26.335 150.955 31.635 151.095 ;
        RECT 26.335 150.910 26.625 150.955 ;
        RECT 29.455 150.910 29.745 150.955 ;
        RECT 31.345 150.910 31.635 150.955 ;
        RECT 34.500 151.095 34.820 151.155 ;
        RECT 38.180 151.095 38.500 151.155 ;
        RECT 34.500 150.955 38.500 151.095 ;
        RECT 34.500 150.895 34.820 150.955 ;
        RECT 38.180 150.895 38.500 150.955 ;
        RECT 18.875 150.570 19.165 150.800 ;
        RECT 19.335 150.755 19.625 150.800 ;
        RECT 20.240 150.755 20.560 150.815 ;
        RECT 22.540 150.755 22.860 150.815 ;
        RECT 19.335 150.615 22.860 150.755 ;
        RECT 19.335 150.570 19.625 150.615 ;
        RECT 20.240 150.555 20.560 150.615 ;
        RECT 22.540 150.555 22.860 150.615 ;
        RECT 23.475 150.755 23.765 150.800 ;
        RECT 30.360 150.755 30.680 150.815 ;
        RECT 23.475 150.615 30.680 150.755 ;
        RECT 23.475 150.570 23.765 150.615 ;
        RECT 30.360 150.555 30.680 150.615 ;
        RECT 32.200 150.555 32.520 150.815 ;
        RECT 40.940 150.755 41.260 150.815 ;
        RECT 32.750 150.615 41.260 150.755 ;
        RECT 22.095 150.230 22.385 150.460 ;
        RECT 15.640 150.075 15.960 150.135 ;
        RECT 22.170 150.075 22.310 150.230 ;
        RECT 25.255 150.120 25.545 150.435 ;
        RECT 26.335 150.415 26.625 150.460 ;
        RECT 29.915 150.415 30.205 150.460 ;
        RECT 31.750 150.415 32.040 150.460 ;
        RECT 32.750 150.415 32.890 150.615 ;
        RECT 40.940 150.555 41.260 150.615 ;
        RECT 26.335 150.275 32.040 150.415 ;
        RECT 26.335 150.230 26.625 150.275 ;
        RECT 29.915 150.230 30.205 150.275 ;
        RECT 31.750 150.230 32.040 150.275 ;
        RECT 32.290 150.275 32.890 150.415 ;
        RECT 35.420 150.415 35.740 150.475 ;
        RECT 36.355 150.415 36.645 150.460 ;
        RECT 35.420 150.275 36.645 150.415 ;
        RECT 15.640 149.935 22.310 150.075 ;
        RECT 15.640 149.875 15.960 149.935 ;
        RECT 19.780 149.535 20.100 149.795 ;
        RECT 22.170 149.735 22.310 149.935 ;
        RECT 22.555 150.075 22.845 150.120 ;
        RECT 24.955 150.075 25.545 150.120 ;
        RECT 28.195 150.075 28.845 150.120 ;
        RECT 22.555 149.935 28.845 150.075 ;
        RECT 22.555 149.890 22.845 149.935 ;
        RECT 24.955 149.890 25.245 149.935 ;
        RECT 28.195 149.890 28.845 149.935 ;
        RECT 30.820 149.875 31.140 150.135 ;
        RECT 23.460 149.735 23.780 149.795 ;
        RECT 32.290 149.735 32.430 150.275 ;
        RECT 35.420 150.215 35.740 150.275 ;
        RECT 36.355 150.230 36.645 150.275 ;
        RECT 36.815 150.230 37.105 150.460 ;
        RECT 36.890 150.075 37.030 150.230 ;
        RECT 37.260 150.215 37.580 150.475 ;
        RECT 38.180 150.215 38.500 150.475 ;
        RECT 45.540 150.215 45.860 150.475 ;
        RECT 46.090 150.460 46.230 151.295 ;
        RECT 46.460 151.235 46.780 151.295 ;
        RECT 48.300 151.095 48.620 151.155 ;
        RECT 59.200 151.095 59.340 151.295 ;
        RECT 62.560 151.295 63.785 151.435 ;
        RECT 62.560 151.235 62.880 151.295 ;
        RECT 63.495 151.250 63.785 151.295 ;
        RECT 85.560 151.235 85.880 151.495 ;
        RECT 87.400 151.235 87.720 151.495 ;
        RECT 100.280 151.235 100.600 151.495 ;
        RECT 65.780 151.095 66.100 151.155 ;
        RECT 48.300 150.955 50.370 151.095 ;
        RECT 59.200 150.955 66.100 151.095 ;
        RECT 48.300 150.895 48.620 150.955 ;
        RECT 49.680 150.755 50.000 150.815 ;
        RECT 50.230 150.800 50.370 150.955 ;
        RECT 65.780 150.895 66.100 150.955 ;
        RECT 71.300 151.095 71.620 151.155 ;
        RECT 74.535 151.095 74.825 151.140 ;
        RECT 71.300 150.955 74.825 151.095 ;
        RECT 71.300 150.895 71.620 150.955 ;
        RECT 74.535 150.910 74.825 150.955 ;
        RECT 84.195 150.910 84.485 151.140 ;
        RECT 106.505 151.095 106.795 151.140 ;
        RECT 107.180 151.095 107.500 151.155 ;
        RECT 106.505 150.955 107.500 151.095 ;
        RECT 106.505 150.910 106.795 150.955 ;
        RECT 46.550 150.615 50.000 150.755 ;
        RECT 46.550 150.460 46.690 150.615 ;
        RECT 49.680 150.555 50.000 150.615 ;
        RECT 50.155 150.570 50.445 150.800 ;
        RECT 65.870 150.755 66.010 150.895 ;
        RECT 65.870 150.615 77.050 150.755 ;
        RECT 76.910 150.475 77.050 150.615 ;
        RECT 80.960 150.555 81.280 150.815 ;
        RECT 81.880 150.555 82.200 150.815 ;
        RECT 84.270 150.755 84.410 150.910 ;
        RECT 107.180 150.895 107.500 150.955 ;
        RECT 110.370 151.095 110.660 151.140 ;
        RECT 113.150 151.095 113.440 151.140 ;
        RECT 115.010 151.095 115.300 151.140 ;
        RECT 110.370 150.955 115.300 151.095 ;
        RECT 110.370 150.910 110.660 150.955 ;
        RECT 113.150 150.910 113.440 150.955 ;
        RECT 115.010 150.910 115.300 150.955 ;
        RECT 97.980 150.755 98.300 150.815 ;
        RECT 99.835 150.755 100.125 150.800 ;
        RECT 84.270 150.615 86.710 150.755 ;
        RECT 46.015 150.230 46.305 150.460 ;
        RECT 46.475 150.230 46.765 150.460 ;
        RECT 47.395 150.415 47.685 150.460 ;
        RECT 48.760 150.415 49.080 150.475 ;
        RECT 47.395 150.275 49.080 150.415 ;
        RECT 47.395 150.230 47.685 150.275 ;
        RECT 48.760 150.215 49.080 150.275 ;
        RECT 60.720 150.415 61.040 150.475 ;
        RECT 63.020 150.415 63.340 150.475 ;
        RECT 63.955 150.415 64.245 150.460 ;
        RECT 60.720 150.275 64.245 150.415 ;
        RECT 60.720 150.215 61.040 150.275 ;
        RECT 63.020 150.215 63.340 150.275 ;
        RECT 63.955 150.230 64.245 150.275 ;
        RECT 70.840 150.415 71.160 150.475 ;
        RECT 71.315 150.415 71.605 150.460 ;
        RECT 70.840 150.275 71.605 150.415 ;
        RECT 70.840 150.215 71.160 150.275 ;
        RECT 71.315 150.230 71.605 150.275 ;
        RECT 71.760 150.415 72.080 150.475 ;
        RECT 72.235 150.415 72.525 150.460 ;
        RECT 71.760 150.275 72.525 150.415 ;
        RECT 71.760 150.215 72.080 150.275 ;
        RECT 72.235 150.230 72.525 150.275 ;
        RECT 72.680 150.215 73.000 150.475 ;
        RECT 73.155 150.415 73.445 150.460 ;
        RECT 73.600 150.415 73.920 150.475 ;
        RECT 73.155 150.275 73.920 150.415 ;
        RECT 73.155 150.230 73.445 150.275 ;
        RECT 73.600 150.215 73.920 150.275 ;
        RECT 76.375 150.230 76.665 150.460 ;
        RECT 37.720 150.075 38.040 150.135 ;
        RECT 39.560 150.075 39.880 150.135 ;
        RECT 36.890 149.935 39.880 150.075 ;
        RECT 37.720 149.875 38.040 149.935 ;
        RECT 39.560 149.875 39.880 149.935 ;
        RECT 44.620 150.075 44.940 150.135 ;
        RECT 50.140 150.075 50.460 150.135 ;
        RECT 51.535 150.075 51.825 150.120 ;
        RECT 44.620 149.935 51.825 150.075 ;
        RECT 44.620 149.875 44.940 149.935 ;
        RECT 50.140 149.875 50.460 149.935 ;
        RECT 51.535 149.890 51.825 149.935 ;
        RECT 61.180 150.075 61.500 150.135 ;
        RECT 75.900 150.075 76.220 150.135 ;
        RECT 76.450 150.075 76.590 150.230 ;
        RECT 76.820 150.215 77.140 150.475 ;
        RECT 77.295 150.230 77.585 150.460 ;
        RECT 77.740 150.415 78.060 150.475 ;
        RECT 78.215 150.415 78.505 150.460 ;
        RECT 77.740 150.275 78.505 150.415 ;
        RECT 61.180 149.935 76.590 150.075 ;
        RECT 77.370 150.075 77.510 150.230 ;
        RECT 77.740 150.215 78.060 150.275 ;
        RECT 78.215 150.230 78.505 150.275 ;
        RECT 81.970 150.075 82.110 150.555 ;
        RECT 86.020 150.215 86.340 150.475 ;
        RECT 86.570 150.460 86.710 150.615 ;
        RECT 97.980 150.615 100.125 150.755 ;
        RECT 97.980 150.555 98.300 150.615 ;
        RECT 99.835 150.570 100.125 150.615 ;
        RECT 86.495 150.230 86.785 150.460 ;
        RECT 99.360 150.215 99.680 150.475 ;
        RECT 100.740 150.215 101.060 150.475 ;
        RECT 104.895 150.415 105.185 150.460 ;
        RECT 106.260 150.415 106.580 150.475 ;
        RECT 104.895 150.275 106.580 150.415 ;
        RECT 104.895 150.230 105.185 150.275 ;
        RECT 106.260 150.215 106.580 150.275 ;
        RECT 110.370 150.415 110.660 150.460 ;
        RECT 110.370 150.275 112.905 150.415 ;
        RECT 110.370 150.230 110.660 150.275 ;
        RECT 77.370 149.935 82.110 150.075 ;
        RECT 106.720 150.075 107.040 150.135 ;
        RECT 112.690 150.120 112.905 150.275 ;
        RECT 113.620 150.215 113.940 150.475 ;
        RECT 115.460 150.215 115.780 150.475 ;
        RECT 116.840 150.215 117.160 150.475 ;
        RECT 108.510 150.075 108.800 150.120 ;
        RECT 111.770 150.075 112.060 150.120 ;
        RECT 106.720 149.935 112.060 150.075 ;
        RECT 61.180 149.875 61.500 149.935 ;
        RECT 75.900 149.875 76.220 149.935 ;
        RECT 106.720 149.875 107.040 149.935 ;
        RECT 108.510 149.890 108.800 149.935 ;
        RECT 111.770 149.890 112.060 149.935 ;
        RECT 112.690 150.075 112.980 150.120 ;
        RECT 114.550 150.075 114.840 150.120 ;
        RECT 112.690 149.935 114.840 150.075 ;
        RECT 112.690 149.890 112.980 149.935 ;
        RECT 114.550 149.890 114.840 149.935 ;
        RECT 22.170 149.595 32.430 149.735 ;
        RECT 34.040 149.735 34.360 149.795 ;
        RECT 34.975 149.735 35.265 149.780 ;
        RECT 34.040 149.595 35.265 149.735 ;
        RECT 23.460 149.535 23.780 149.595 ;
        RECT 34.040 149.535 34.360 149.595 ;
        RECT 34.975 149.550 35.265 149.595 ;
        RECT 35.420 149.735 35.740 149.795 ;
        RECT 44.175 149.735 44.465 149.780 ;
        RECT 35.420 149.595 44.465 149.735 ;
        RECT 35.420 149.535 35.740 149.595 ;
        RECT 44.175 149.550 44.465 149.595 ;
        RECT 47.380 149.735 47.700 149.795 ;
        RECT 51.075 149.735 51.365 149.780 ;
        RECT 47.380 149.595 51.365 149.735 ;
        RECT 47.380 149.535 47.700 149.595 ;
        RECT 51.075 149.550 51.365 149.595 ;
        RECT 53.375 149.735 53.665 149.780 ;
        RECT 55.200 149.735 55.520 149.795 ;
        RECT 53.375 149.595 55.520 149.735 ;
        RECT 53.375 149.550 53.665 149.595 ;
        RECT 55.200 149.535 55.520 149.595 ;
        RECT 74.520 149.735 74.840 149.795 ;
        RECT 74.995 149.735 75.285 149.780 ;
        RECT 74.520 149.595 75.285 149.735 ;
        RECT 74.520 149.535 74.840 149.595 ;
        RECT 74.995 149.550 75.285 149.595 ;
        RECT 82.340 149.535 82.660 149.795 ;
        RECT 101.200 149.735 101.520 149.795 ;
        RECT 101.675 149.735 101.965 149.780 ;
        RECT 101.200 149.595 101.965 149.735 ;
        RECT 101.200 149.535 101.520 149.595 ;
        RECT 101.675 149.550 101.965 149.595 ;
        RECT 105.340 149.535 105.660 149.795 ;
        RECT 115.000 149.735 115.320 149.795 ;
        RECT 115.935 149.735 116.225 149.780 ;
        RECT 115.000 149.595 116.225 149.735 ;
        RECT 115.000 149.535 115.320 149.595 ;
        RECT 115.935 149.550 116.225 149.595 ;
        RECT 10.650 148.915 118.610 149.395 ;
        RECT 25.300 148.515 25.620 148.775 ;
        RECT 30.820 148.515 31.140 148.775 ;
        RECT 34.500 148.715 34.820 148.775 ;
        RECT 38.180 148.715 38.500 148.775 ;
        RECT 45.540 148.715 45.860 148.775 ;
        RECT 31.830 148.575 38.500 148.715 ;
        RECT 14.260 148.375 14.580 148.435 ;
        RECT 15.295 148.375 15.585 148.420 ;
        RECT 18.535 148.375 19.185 148.420 ;
        RECT 14.260 148.235 19.185 148.375 ;
        RECT 14.260 148.175 14.580 148.235 ;
        RECT 15.295 148.190 15.885 148.235 ;
        RECT 18.535 148.190 19.185 148.235 ;
        RECT 25.775 148.375 26.065 148.420 ;
        RECT 25.775 148.235 27.830 148.375 ;
        RECT 25.775 148.190 26.065 148.235 ;
        RECT 15.595 147.875 15.885 148.190 ;
        RECT 16.675 148.035 16.965 148.080 ;
        RECT 20.255 148.035 20.545 148.080 ;
        RECT 22.090 148.035 22.380 148.080 ;
        RECT 16.675 147.895 22.380 148.035 ;
        RECT 16.675 147.850 16.965 147.895 ;
        RECT 20.255 147.850 20.545 147.895 ;
        RECT 22.090 147.850 22.380 147.895 ;
        RECT 22.555 148.035 22.845 148.080 ;
        RECT 27.140 148.035 27.460 148.095 ;
        RECT 22.555 147.895 27.460 148.035 ;
        RECT 22.555 147.850 22.845 147.895 ;
        RECT 27.140 147.835 27.460 147.895 ;
        RECT 17.940 147.695 18.260 147.755 ;
        RECT 21.175 147.695 21.465 147.740 ;
        RECT 17.940 147.555 21.465 147.695 ;
        RECT 17.940 147.495 18.260 147.555 ;
        RECT 21.175 147.510 21.465 147.555 ;
        RECT 24.380 147.695 24.700 147.755 ;
        RECT 26.235 147.695 26.525 147.740 ;
        RECT 24.380 147.555 26.525 147.695 ;
        RECT 24.380 147.495 24.700 147.555 ;
        RECT 26.235 147.510 26.525 147.555 ;
        RECT 16.675 147.355 16.965 147.400 ;
        RECT 19.795 147.355 20.085 147.400 ;
        RECT 21.685 147.355 21.975 147.400 ;
        RECT 16.675 147.215 21.975 147.355 ;
        RECT 16.675 147.170 16.965 147.215 ;
        RECT 19.795 147.170 20.085 147.215 ;
        RECT 21.685 147.170 21.975 147.215 ;
        RECT 22.540 147.355 22.860 147.415 ;
        RECT 27.690 147.355 27.830 148.235 ;
        RECT 29.900 147.835 30.220 148.095 ;
        RECT 31.295 148.035 31.585 148.080 ;
        RECT 31.830 148.035 31.970 148.575 ;
        RECT 34.500 148.515 34.820 148.575 ;
        RECT 38.180 148.515 38.500 148.575 ;
        RECT 41.950 148.575 45.860 148.715 ;
        RECT 33.210 148.235 37.030 148.375 ;
        RECT 31.295 147.895 31.970 148.035 ;
        RECT 31.295 147.850 31.585 147.895 ;
        RECT 32.200 147.835 32.520 148.095 ;
        RECT 32.660 147.835 32.980 148.095 ;
        RECT 33.210 148.080 33.350 148.235 ;
        RECT 36.890 148.095 37.030 148.235 ;
        RECT 33.135 147.850 33.425 148.080 ;
        RECT 34.500 148.035 34.820 148.095 ;
        RECT 34.975 148.035 35.265 148.080 ;
        RECT 34.500 147.895 35.265 148.035 ;
        RECT 34.500 147.835 34.820 147.895 ;
        RECT 34.975 147.850 35.265 147.895 ;
        RECT 35.895 147.850 36.185 148.080 ;
        RECT 36.355 147.850 36.645 148.080 ;
        RECT 30.360 147.695 30.680 147.755 ;
        RECT 35.970 147.695 36.110 147.850 ;
        RECT 30.360 147.555 36.110 147.695 ;
        RECT 36.430 147.695 36.570 147.850 ;
        RECT 36.800 147.835 37.120 148.095 ;
        RECT 41.950 148.080 42.090 148.575 ;
        RECT 45.540 148.515 45.860 148.575 ;
        RECT 80.960 148.715 81.280 148.775 ;
        RECT 96.140 148.715 96.460 148.775 ;
        RECT 99.835 148.715 100.125 148.760 ;
        RECT 80.960 148.575 93.610 148.715 ;
        RECT 80.960 148.515 81.280 148.575 ;
        RECT 44.620 148.375 44.940 148.435 ;
        RECT 49.680 148.420 50.000 148.435 ;
        RECT 42.870 148.235 44.940 148.375 ;
        RECT 42.870 148.080 43.010 148.235 ;
        RECT 44.620 148.175 44.940 148.235 ;
        RECT 46.410 148.375 46.700 148.420 ;
        RECT 49.670 148.375 50.000 148.420 ;
        RECT 46.410 148.235 50.000 148.375 ;
        RECT 46.410 148.190 46.700 148.235 ;
        RECT 49.670 148.190 50.000 148.235 ;
        RECT 49.680 148.175 50.000 148.190 ;
        RECT 50.590 148.375 50.880 148.420 ;
        RECT 52.450 148.375 52.740 148.420 ;
        RECT 50.590 148.235 52.740 148.375 ;
        RECT 50.590 148.190 50.880 148.235 ;
        RECT 52.450 148.190 52.740 148.235 ;
        RECT 41.875 147.850 42.165 148.080 ;
        RECT 42.335 147.850 42.625 148.080 ;
        RECT 42.795 147.850 43.085 148.080 ;
        RECT 43.715 147.850 44.005 148.080 ;
        RECT 48.270 148.035 48.560 148.080 ;
        RECT 50.590 148.035 50.805 148.190 ;
        RECT 74.520 148.175 74.840 148.435 ;
        RECT 86.480 148.420 86.800 148.435 ;
        RECT 83.210 148.375 83.500 148.420 ;
        RECT 86.470 148.375 86.800 148.420 ;
        RECT 83.210 148.235 86.800 148.375 ;
        RECT 83.210 148.190 83.500 148.235 ;
        RECT 86.470 148.190 86.800 148.235 ;
        RECT 86.480 148.175 86.800 148.190 ;
        RECT 87.390 148.375 87.680 148.420 ;
        RECT 89.250 148.375 89.540 148.420 ;
        RECT 87.390 148.235 89.540 148.375 ;
        RECT 87.390 148.190 87.680 148.235 ;
        RECT 89.250 148.190 89.540 148.235 ;
        RECT 48.270 147.895 50.805 148.035 ;
        RECT 51.535 148.035 51.825 148.080 ;
        RECT 51.535 147.895 54.510 148.035 ;
        RECT 48.270 147.850 48.560 147.895 ;
        RECT 51.535 147.850 51.825 147.895 ;
        RECT 39.560 147.695 39.880 147.755 ;
        RECT 36.430 147.555 39.880 147.695 ;
        RECT 30.360 147.495 30.680 147.555 ;
        RECT 31.280 147.355 31.600 147.415 ;
        RECT 22.540 147.215 31.600 147.355 ;
        RECT 22.540 147.155 22.860 147.215 ;
        RECT 31.280 147.155 31.600 147.215 ;
        RECT 32.660 147.355 32.980 147.415 ;
        RECT 36.430 147.355 36.570 147.555 ;
        RECT 39.560 147.495 39.880 147.555 ;
        RECT 32.660 147.215 36.570 147.355 ;
        RECT 42.410 147.355 42.550 147.850 ;
        RECT 43.790 147.695 43.930 147.850 ;
        RECT 48.760 147.695 49.080 147.755 ;
        RECT 43.790 147.555 49.080 147.695 ;
        RECT 48.760 147.495 49.080 147.555 ;
        RECT 53.360 147.495 53.680 147.755 ;
        RECT 46.460 147.355 46.780 147.415 ;
        RECT 54.370 147.400 54.510 147.895 ;
        RECT 55.200 147.835 55.520 148.095 ;
        RECT 57.515 148.035 57.805 148.080 ;
        RECT 55.750 147.895 57.805 148.035 ;
        RECT 42.410 147.215 46.780 147.355 ;
        RECT 32.660 147.155 32.980 147.215 ;
        RECT 46.460 147.155 46.780 147.215 ;
        RECT 48.270 147.355 48.560 147.400 ;
        RECT 51.050 147.355 51.340 147.400 ;
        RECT 52.910 147.355 53.200 147.400 ;
        RECT 48.270 147.215 53.200 147.355 ;
        RECT 48.270 147.170 48.560 147.215 ;
        RECT 51.050 147.170 51.340 147.215 ;
        RECT 52.910 147.170 53.200 147.215 ;
        RECT 54.295 147.170 54.585 147.400 ;
        RECT 13.800 146.815 14.120 147.075 ;
        RECT 23.460 146.815 23.780 147.075 ;
        RECT 33.120 147.015 33.440 147.075 ;
        RECT 34.515 147.015 34.805 147.060 ;
        RECT 33.120 146.875 34.805 147.015 ;
        RECT 33.120 146.815 33.440 146.875 ;
        RECT 34.515 146.830 34.805 146.875 ;
        RECT 36.800 147.015 37.120 147.075 ;
        RECT 38.195 147.015 38.485 147.060 ;
        RECT 36.800 146.875 38.485 147.015 ;
        RECT 36.800 146.815 37.120 146.875 ;
        RECT 38.195 146.830 38.485 146.875 ;
        RECT 40.480 146.815 40.800 147.075 ;
        RECT 44.405 147.015 44.695 147.060 ;
        RECT 47.380 147.015 47.700 147.075 ;
        RECT 44.405 146.875 47.700 147.015 ;
        RECT 44.405 146.830 44.695 146.875 ;
        RECT 47.380 146.815 47.700 146.875 ;
        RECT 49.220 147.015 49.540 147.075 ;
        RECT 55.750 147.015 55.890 147.895 ;
        RECT 57.515 147.850 57.805 147.895 ;
        RECT 66.255 148.035 66.545 148.080 ;
        RECT 67.620 148.035 67.940 148.095 ;
        RECT 66.255 147.895 67.940 148.035 ;
        RECT 66.255 147.850 66.545 147.895 ;
        RECT 67.620 147.835 67.940 147.895 ;
        RECT 73.140 147.835 73.460 148.095 ;
        RECT 85.070 148.035 85.360 148.080 ;
        RECT 87.390 148.035 87.605 148.190 ;
        RECT 85.070 147.895 87.605 148.035 ;
        RECT 85.070 147.850 85.360 147.895 ;
        RECT 74.060 147.495 74.380 147.755 ;
        RECT 88.320 147.495 88.640 147.755 ;
        RECT 89.240 147.695 89.560 147.755 ;
        RECT 90.175 147.695 90.465 147.740 ;
        RECT 89.240 147.555 90.465 147.695 ;
        RECT 93.470 147.695 93.610 148.575 ;
        RECT 96.140 148.575 100.125 148.715 ;
        RECT 96.140 148.515 96.460 148.575 ;
        RECT 99.835 148.530 100.125 148.575 ;
        RECT 106.720 148.515 107.040 148.775 ;
        RECT 108.100 148.760 108.420 148.775 ;
        RECT 107.885 148.530 108.420 148.760 ;
        RECT 108.100 148.515 108.420 148.530 ;
        RECT 100.295 148.375 100.585 148.420 ;
        RECT 101.660 148.375 101.980 148.435 ;
        RECT 105.340 148.375 105.660 148.435 ;
        RECT 109.890 148.375 110.180 148.420 ;
        RECT 113.150 148.375 113.440 148.420 ;
        RECT 100.295 148.235 104.190 148.375 ;
        RECT 100.295 148.190 100.585 148.235 ;
        RECT 101.660 148.175 101.980 148.235 ;
        RECT 94.850 147.895 99.130 148.035 ;
        RECT 94.850 147.740 94.990 147.895 ;
        RECT 98.990 147.755 99.130 147.895 ;
        RECT 94.775 147.695 95.065 147.740 ;
        RECT 93.470 147.555 95.065 147.695 ;
        RECT 89.240 147.495 89.560 147.555 ;
        RECT 90.175 147.510 90.465 147.555 ;
        RECT 94.775 147.510 95.065 147.555 ;
        RECT 95.695 147.510 95.985 147.740 ;
        RECT 70.840 147.355 71.160 147.415 ;
        RECT 81.205 147.355 81.495 147.400 ;
        RECT 82.340 147.355 82.660 147.415 ;
        RECT 70.840 147.215 73.370 147.355 ;
        RECT 70.840 147.155 71.160 147.215 ;
        RECT 49.220 146.875 55.890 147.015 ;
        RECT 49.220 146.815 49.540 146.875 ;
        RECT 57.960 146.815 58.280 147.075 ;
        RECT 63.480 147.015 63.800 147.075 ;
        RECT 65.335 147.015 65.625 147.060 ;
        RECT 63.480 146.875 65.625 147.015 ;
        RECT 63.480 146.815 63.800 146.875 ;
        RECT 65.335 146.830 65.625 146.875 ;
        RECT 71.760 147.015 72.080 147.075 ;
        RECT 73.230 147.060 73.370 147.215 ;
        RECT 81.205 147.215 82.660 147.355 ;
        RECT 81.205 147.170 81.495 147.215 ;
        RECT 82.340 147.155 82.660 147.215 ;
        RECT 85.070 147.355 85.360 147.400 ;
        RECT 87.850 147.355 88.140 147.400 ;
        RECT 89.710 147.355 90.000 147.400 ;
        RECT 85.070 147.215 90.000 147.355 ;
        RECT 85.070 147.170 85.360 147.215 ;
        RECT 87.850 147.170 88.140 147.215 ;
        RECT 89.710 147.170 90.000 147.215 ;
        RECT 92.920 147.355 93.240 147.415 ;
        RECT 95.770 147.355 95.910 147.510 ;
        RECT 98.900 147.495 99.220 147.755 ;
        RECT 104.050 147.695 104.190 148.235 ;
        RECT 105.340 148.235 113.440 148.375 ;
        RECT 105.340 148.175 105.660 148.235 ;
        RECT 109.890 148.190 110.180 148.235 ;
        RECT 113.150 148.190 113.440 148.235 ;
        RECT 114.070 148.375 114.360 148.420 ;
        RECT 115.930 148.375 116.220 148.420 ;
        RECT 114.070 148.235 116.220 148.375 ;
        RECT 114.070 148.190 114.360 148.235 ;
        RECT 115.930 148.190 116.220 148.235 ;
        RECT 106.260 147.835 106.580 148.095 ;
        RECT 111.750 148.035 112.040 148.080 ;
        RECT 114.070 148.035 114.285 148.190 ;
        RECT 111.750 147.895 114.285 148.035 ;
        RECT 111.750 147.850 112.040 147.895 ;
        RECT 115.000 147.835 115.320 148.095 ;
        RECT 107.180 147.695 107.500 147.755 ;
        RECT 104.050 147.555 107.500 147.695 ;
        RECT 107.180 147.495 107.500 147.555 ;
        RECT 115.460 147.695 115.780 147.755 ;
        RECT 116.855 147.695 117.145 147.740 ;
        RECT 115.460 147.555 117.145 147.695 ;
        RECT 115.460 147.495 115.780 147.555 ;
        RECT 116.855 147.510 117.145 147.555 ;
        RECT 92.920 147.215 95.910 147.355 ;
        RECT 111.750 147.355 112.040 147.400 ;
        RECT 114.530 147.355 114.820 147.400 ;
        RECT 116.390 147.355 116.680 147.400 ;
        RECT 111.750 147.215 116.680 147.355 ;
        RECT 92.920 147.155 93.240 147.215 ;
        RECT 111.750 147.170 112.040 147.215 ;
        RECT 114.530 147.170 114.820 147.215 ;
        RECT 116.390 147.170 116.680 147.215 ;
        RECT 72.235 147.015 72.525 147.060 ;
        RECT 71.760 146.875 72.525 147.015 ;
        RECT 71.760 146.815 72.080 146.875 ;
        RECT 72.235 146.830 72.525 146.875 ;
        RECT 73.155 146.830 73.445 147.060 ;
        RECT 97.980 146.815 98.300 147.075 ;
        RECT 102.120 146.815 102.440 147.075 ;
        RECT 11.430 146.195 118.610 146.675 ;
        RECT 14.260 145.795 14.580 146.055 ;
        RECT 17.940 145.795 18.260 146.055 ;
        RECT 18.415 145.995 18.705 146.040 ;
        RECT 22.540 145.995 22.860 146.055 ;
        RECT 18.415 145.855 22.860 145.995 ;
        RECT 18.415 145.810 18.705 145.855 ;
        RECT 22.540 145.795 22.860 145.855 ;
        RECT 31.280 145.995 31.600 146.055 ;
        RECT 33.135 145.995 33.425 146.040 ;
        RECT 31.280 145.855 33.425 145.995 ;
        RECT 31.280 145.795 31.600 145.855 ;
        RECT 33.135 145.810 33.425 145.855 ;
        RECT 49.680 145.995 50.000 146.055 ;
        RECT 51.075 145.995 51.365 146.040 ;
        RECT 49.680 145.855 51.365 145.995 ;
        RECT 49.680 145.795 50.000 145.855 ;
        RECT 51.075 145.810 51.365 145.855 ;
        RECT 55.905 145.995 56.195 146.040 ;
        RECT 57.500 145.995 57.820 146.055 ;
        RECT 55.905 145.855 57.820 145.995 ;
        RECT 55.905 145.810 56.195 145.855 ;
        RECT 57.500 145.795 57.820 145.855 ;
        RECT 72.680 145.995 73.000 146.055 ;
        RECT 73.155 145.995 73.445 146.040 ;
        RECT 72.680 145.855 73.445 145.995 ;
        RECT 72.680 145.795 73.000 145.855 ;
        RECT 73.155 145.810 73.445 145.855 ;
        RECT 86.035 145.995 86.325 146.040 ;
        RECT 86.480 145.995 86.800 146.055 ;
        RECT 86.035 145.855 86.800 145.995 ;
        RECT 86.035 145.810 86.325 145.855 ;
        RECT 86.480 145.795 86.800 145.855 ;
        RECT 87.875 145.995 88.165 146.040 ;
        RECT 88.320 145.995 88.640 146.055 ;
        RECT 87.875 145.855 88.640 145.995 ;
        RECT 87.875 145.810 88.165 145.855 ;
        RECT 88.320 145.795 88.640 145.855 ;
        RECT 95.465 145.995 95.755 146.040 ;
        RECT 96.140 145.995 96.460 146.055 ;
        RECT 95.465 145.855 96.460 145.995 ;
        RECT 95.465 145.810 95.755 145.855 ;
        RECT 96.140 145.795 96.460 145.855 ;
        RECT 112.255 145.995 112.545 146.040 ;
        RECT 113.620 145.995 113.940 146.055 ;
        RECT 112.255 145.855 113.940 145.995 ;
        RECT 112.255 145.810 112.545 145.855 ;
        RECT 113.620 145.795 113.940 145.855 ;
        RECT 21.275 145.655 21.565 145.700 ;
        RECT 24.395 145.655 24.685 145.700 ;
        RECT 26.285 145.655 26.575 145.700 ;
        RECT 33.580 145.655 33.900 145.715 ;
        RECT 37.720 145.655 38.040 145.715 ;
        RECT 21.275 145.515 26.575 145.655 ;
        RECT 21.275 145.470 21.565 145.515 ;
        RECT 24.395 145.470 24.685 145.515 ;
        RECT 26.285 145.470 26.575 145.515 ;
        RECT 33.210 145.515 33.900 145.655 ;
        RECT 27.140 145.115 27.460 145.375 ;
        RECT 14.735 144.975 15.025 145.020 ;
        RECT 15.640 144.975 15.960 145.035 ;
        RECT 14.735 144.835 15.960 144.975 ;
        RECT 14.735 144.790 15.025 144.835 ;
        RECT 15.640 144.775 15.960 144.835 ;
        RECT 17.020 144.775 17.340 145.035 ;
        RECT 33.210 145.020 33.350 145.515 ;
        RECT 33.580 145.455 33.900 145.515 ;
        RECT 36.430 145.515 38.040 145.655 ;
        RECT 20.195 144.680 20.485 144.995 ;
        RECT 21.275 144.975 21.565 145.020 ;
        RECT 24.855 144.975 25.145 145.020 ;
        RECT 26.690 144.975 26.980 145.020 ;
        RECT 21.275 144.835 26.980 144.975 ;
        RECT 21.275 144.790 21.565 144.835 ;
        RECT 24.855 144.790 25.145 144.835 ;
        RECT 26.690 144.790 26.980 144.835 ;
        RECT 33.135 144.790 33.425 145.020 ;
        RECT 33.595 144.975 33.885 145.020 ;
        RECT 34.040 144.975 34.360 145.035 ;
        RECT 33.595 144.835 34.360 144.975 ;
        RECT 33.595 144.790 33.885 144.835 ;
        RECT 34.040 144.775 34.360 144.835 ;
        RECT 34.515 144.975 34.805 145.020 ;
        RECT 35.420 144.975 35.740 145.035 ;
        RECT 36.430 145.020 36.570 145.515 ;
        RECT 37.720 145.455 38.040 145.515 ;
        RECT 59.770 145.655 60.060 145.700 ;
        RECT 62.550 145.655 62.840 145.700 ;
        RECT 64.410 145.655 64.700 145.700 ;
        RECT 59.770 145.515 64.700 145.655 ;
        RECT 59.770 145.470 60.060 145.515 ;
        RECT 62.550 145.470 62.840 145.515 ;
        RECT 64.410 145.470 64.700 145.515 ;
        RECT 75.900 145.455 76.220 145.715 ;
        RECT 85.115 145.470 85.405 145.700 ;
        RECT 99.330 145.655 99.620 145.700 ;
        RECT 102.110 145.655 102.400 145.700 ;
        RECT 103.970 145.655 104.260 145.700 ;
        RECT 99.330 145.515 104.260 145.655 ;
        RECT 99.330 145.470 99.620 145.515 ;
        RECT 102.110 145.470 102.400 145.515 ;
        RECT 103.970 145.470 104.260 145.515 ;
        RECT 109.955 145.470 110.245 145.700 ;
        RECT 39.560 145.315 39.880 145.375 ;
        RECT 36.890 145.175 39.880 145.315 ;
        RECT 36.890 145.020 37.030 145.175 ;
        RECT 39.560 145.115 39.880 145.175 ;
        RECT 53.360 145.315 53.680 145.375 ;
        RECT 53.360 145.175 62.790 145.315 ;
        RECT 53.360 145.115 53.680 145.175 ;
        RECT 34.515 144.835 35.740 144.975 ;
        RECT 34.515 144.790 34.805 144.835 ;
        RECT 35.420 144.775 35.740 144.835 ;
        RECT 36.355 144.790 36.645 145.020 ;
        RECT 36.815 144.790 37.105 145.020 ;
        RECT 37.260 144.775 37.580 145.035 ;
        RECT 38.180 144.775 38.500 145.035 ;
        RECT 45.540 144.975 45.860 145.035 ;
        RECT 46.015 144.975 46.305 145.020 ;
        RECT 45.540 144.835 46.305 144.975 ;
        RECT 45.540 144.775 45.860 144.835 ;
        RECT 46.015 144.790 46.305 144.835 ;
        RECT 46.460 144.775 46.780 145.035 ;
        RECT 46.935 144.975 47.225 145.020 ;
        RECT 47.380 144.975 47.700 145.035 ;
        RECT 46.935 144.835 47.700 144.975 ;
        RECT 46.935 144.790 47.225 144.835 ;
        RECT 47.380 144.775 47.700 144.835 ;
        RECT 47.855 144.975 48.145 145.020 ;
        RECT 48.760 144.975 49.080 145.035 ;
        RECT 47.855 144.835 49.080 144.975 ;
        RECT 47.855 144.790 48.145 144.835 ;
        RECT 48.760 144.775 49.080 144.835 ;
        RECT 49.220 144.975 49.540 145.035 ;
        RECT 51.535 144.975 51.825 145.020 ;
        RECT 54.295 144.975 54.585 145.020 ;
        RECT 49.220 144.835 54.585 144.975 ;
        RECT 49.220 144.775 49.540 144.835 ;
        RECT 51.535 144.790 51.825 144.835 ;
        RECT 54.295 144.790 54.585 144.835 ;
        RECT 59.770 144.975 60.060 145.020 ;
        RECT 62.650 144.975 62.790 145.175 ;
        RECT 63.020 145.115 63.340 145.375 ;
        RECT 71.300 145.315 71.620 145.375 ;
        RECT 72.695 145.315 72.985 145.360 ;
        RECT 75.990 145.315 76.130 145.455 ;
        RECT 71.300 145.175 72.985 145.315 ;
        RECT 71.300 145.115 71.620 145.175 ;
        RECT 72.695 145.130 72.985 145.175 ;
        RECT 75.530 145.175 76.130 145.315 ;
        RECT 80.960 145.315 81.280 145.375 ;
        RECT 81.895 145.315 82.185 145.360 ;
        RECT 80.960 145.175 82.185 145.315 ;
        RECT 85.190 145.315 85.330 145.470 ;
        RECT 98.900 145.315 99.220 145.375 ;
        RECT 106.735 145.315 107.025 145.360 ;
        RECT 107.640 145.315 107.960 145.375 ;
        RECT 85.190 145.175 87.170 145.315 ;
        RECT 64.875 144.975 65.165 145.020 ;
        RECT 65.780 144.975 66.100 145.035 ;
        RECT 59.770 144.835 62.305 144.975 ;
        RECT 62.650 144.835 66.100 144.975 ;
        RECT 59.770 144.790 60.060 144.835 ;
        RECT 16.115 144.635 16.405 144.680 ;
        RECT 19.895 144.635 20.485 144.680 ;
        RECT 23.135 144.635 23.785 144.680 ;
        RECT 16.115 144.495 23.785 144.635 ;
        RECT 16.115 144.450 16.405 144.495 ;
        RECT 19.895 144.450 20.185 144.495 ;
        RECT 23.135 144.450 23.785 144.495 ;
        RECT 25.760 144.435 26.080 144.695 ;
        RECT 56.120 144.635 56.440 144.695 ;
        RECT 57.960 144.680 58.280 144.695 ;
        RECT 62.090 144.680 62.305 144.835 ;
        RECT 64.875 144.790 65.165 144.835 ;
        RECT 65.780 144.775 66.100 144.835 ;
        RECT 72.220 144.775 72.540 145.035 ;
        RECT 75.530 145.020 75.670 145.175 ;
        RECT 80.960 145.115 81.280 145.175 ;
        RECT 81.895 145.130 82.185 145.175 ;
        RECT 75.455 144.790 75.745 145.020 ;
        RECT 75.915 144.790 76.205 145.020 ;
        RECT 76.375 144.790 76.665 145.020 ;
        RECT 77.295 144.975 77.585 145.020 ;
        RECT 77.740 144.975 78.060 145.035 ;
        RECT 77.295 144.835 78.060 144.975 ;
        RECT 77.295 144.790 77.585 144.835 ;
        RECT 37.350 144.495 56.440 144.635 ;
        RECT 32.215 144.295 32.505 144.340 ;
        RECT 32.660 144.295 32.980 144.355 ;
        RECT 32.215 144.155 32.980 144.295 ;
        RECT 32.215 144.110 32.505 144.155 ;
        RECT 32.660 144.095 32.980 144.155 ;
        RECT 33.580 144.295 33.900 144.355 ;
        RECT 34.975 144.295 35.265 144.340 ;
        RECT 33.580 144.155 35.265 144.295 ;
        RECT 33.580 144.095 33.900 144.155 ;
        RECT 34.975 144.110 35.265 144.155 ;
        RECT 35.420 144.295 35.740 144.355 ;
        RECT 37.350 144.295 37.490 144.495 ;
        RECT 56.120 144.435 56.440 144.495 ;
        RECT 57.910 144.635 58.280 144.680 ;
        RECT 61.170 144.635 61.460 144.680 ;
        RECT 57.910 144.495 61.460 144.635 ;
        RECT 57.910 144.450 58.280 144.495 ;
        RECT 61.170 144.450 61.460 144.495 ;
        RECT 62.090 144.635 62.380 144.680 ;
        RECT 63.950 144.635 64.240 144.680 ;
        RECT 62.090 144.495 64.240 144.635 ;
        RECT 62.090 144.450 62.380 144.495 ;
        RECT 63.950 144.450 64.240 144.495 ;
        RECT 73.615 144.635 73.905 144.680 ;
        RECT 74.075 144.635 74.365 144.680 ;
        RECT 73.615 144.495 74.365 144.635 ;
        RECT 73.615 144.450 73.905 144.495 ;
        RECT 74.075 144.450 74.365 144.495 ;
        RECT 57.960 144.435 58.280 144.450 ;
        RECT 35.420 144.155 37.490 144.295 ;
        RECT 44.160 144.295 44.480 144.355 ;
        RECT 44.635 144.295 44.925 144.340 ;
        RECT 44.160 144.155 44.925 144.295 ;
        RECT 35.420 144.095 35.740 144.155 ;
        RECT 44.160 144.095 44.480 144.155 ;
        RECT 44.635 144.110 44.925 144.155 ;
        RECT 54.740 144.095 55.060 144.355 ;
        RECT 69.920 144.295 70.240 144.355 ;
        RECT 71.315 144.295 71.605 144.340 ;
        RECT 69.920 144.155 71.605 144.295 ;
        RECT 69.920 144.095 70.240 144.155 ;
        RECT 71.315 144.110 71.605 144.155 ;
        RECT 73.140 144.295 73.460 144.355 ;
        RECT 75.990 144.295 76.130 144.790 ;
        RECT 76.450 144.635 76.590 144.790 ;
        RECT 77.740 144.775 78.060 144.835 ;
        RECT 86.020 144.975 86.340 145.035 ;
        RECT 87.030 145.020 87.170 145.175 ;
        RECT 98.900 145.175 107.960 145.315 ;
        RECT 98.900 145.115 99.220 145.175 ;
        RECT 106.735 145.130 107.025 145.175 ;
        RECT 107.640 145.115 107.960 145.175 ;
        RECT 86.495 144.975 86.785 145.020 ;
        RECT 86.020 144.835 86.785 144.975 ;
        RECT 86.020 144.775 86.340 144.835 ;
        RECT 86.495 144.790 86.785 144.835 ;
        RECT 86.955 144.790 87.245 145.020 ;
        RECT 82.340 144.635 82.660 144.695 ;
        RECT 82.815 144.635 83.105 144.680 ;
        RECT 76.450 144.495 83.105 144.635 ;
        RECT 86.570 144.635 86.710 144.790 ;
        RECT 93.840 144.775 94.160 145.035 ;
        RECT 99.330 144.975 99.620 145.020 ;
        RECT 99.330 144.835 101.865 144.975 ;
        RECT 99.330 144.790 99.620 144.835 ;
        RECT 93.930 144.635 94.070 144.775 ;
        RECT 101.650 144.680 101.865 144.835 ;
        RECT 102.580 144.775 102.900 145.035 ;
        RECT 104.420 144.975 104.740 145.035 ;
        RECT 104.420 144.835 107.640 144.975 ;
        RECT 104.420 144.775 104.740 144.835 ;
        RECT 86.570 144.495 94.070 144.635 ;
        RECT 94.315 144.635 94.605 144.680 ;
        RECT 97.470 144.635 97.760 144.680 ;
        RECT 100.730 144.635 101.020 144.680 ;
        RECT 94.315 144.495 101.020 144.635 ;
        RECT 82.340 144.435 82.660 144.495 ;
        RECT 82.815 144.450 83.105 144.495 ;
        RECT 94.315 144.450 94.605 144.495 ;
        RECT 97.470 144.450 97.760 144.495 ;
        RECT 100.730 144.450 101.020 144.495 ;
        RECT 101.650 144.635 101.940 144.680 ;
        RECT 103.510 144.635 103.800 144.680 ;
        RECT 101.650 144.495 103.800 144.635 ;
        RECT 107.500 144.635 107.640 144.835 ;
        RECT 108.100 144.775 108.420 145.035 ;
        RECT 110.030 144.975 110.170 145.470 ;
        RECT 111.335 144.975 111.625 145.020 ;
        RECT 110.030 144.835 111.625 144.975 ;
        RECT 111.335 144.790 111.625 144.835 ;
        RECT 115.460 144.635 115.780 144.695 ;
        RECT 107.500 144.495 115.780 144.635 ;
        RECT 101.650 144.450 101.940 144.495 ;
        RECT 103.510 144.450 103.800 144.495 ;
        RECT 115.460 144.435 115.780 144.495 ;
        RECT 76.820 144.295 77.140 144.355 ;
        RECT 73.140 144.155 77.140 144.295 ;
        RECT 73.140 144.095 73.460 144.155 ;
        RECT 76.820 144.095 77.140 144.155 ;
        RECT 83.260 144.095 83.580 144.355 ;
        RECT 107.180 144.295 107.500 144.355 ;
        RECT 107.655 144.295 107.945 144.340 ;
        RECT 107.180 144.155 107.945 144.295 ;
        RECT 107.180 144.095 107.500 144.155 ;
        RECT 107.655 144.110 107.945 144.155 ;
        RECT 10.650 143.475 118.610 143.955 ;
        RECT 17.020 143.275 17.340 143.335 ;
        RECT 18.875 143.275 19.165 143.320 ;
        RECT 17.020 143.135 19.165 143.275 ;
        RECT 17.020 143.075 17.340 143.135 ;
        RECT 18.875 143.090 19.165 143.135 ;
        RECT 20.715 143.275 21.005 143.320 ;
        RECT 22.540 143.275 22.860 143.335 ;
        RECT 20.715 143.135 22.860 143.275 ;
        RECT 20.715 143.090 21.005 143.135 ;
        RECT 22.540 143.075 22.860 143.135 ;
        RECT 25.315 143.275 25.605 143.320 ;
        RECT 25.760 143.275 26.080 143.335 ;
        RECT 25.315 143.135 26.080 143.275 ;
        RECT 25.315 143.090 25.605 143.135 ;
        RECT 25.760 143.075 26.080 143.135 ;
        RECT 31.280 143.275 31.600 143.335 ;
        RECT 34.500 143.275 34.820 143.335 ;
        RECT 31.280 143.135 34.820 143.275 ;
        RECT 31.280 143.075 31.600 143.135 ;
        RECT 34.500 143.075 34.820 143.135 ;
        RECT 35.420 143.075 35.740 143.335 ;
        RECT 44.160 143.275 44.480 143.335 ;
        RECT 37.350 143.135 44.480 143.275 ;
        RECT 16.575 142.935 16.865 142.980 ;
        RECT 19.780 142.935 20.100 142.995 ;
        RECT 16.575 142.795 20.100 142.935 ;
        RECT 16.575 142.750 16.865 142.795 ;
        RECT 19.780 142.735 20.100 142.795 ;
        RECT 21.175 142.935 21.465 142.980 ;
        RECT 32.200 142.935 32.520 142.995 ;
        RECT 21.175 142.795 32.520 142.935 ;
        RECT 21.175 142.750 21.465 142.795 ;
        RECT 13.800 142.595 14.120 142.655 ;
        RECT 21.250 142.595 21.390 142.750 ;
        RECT 32.200 142.735 32.520 142.795 ;
        RECT 32.675 142.935 32.965 142.980 ;
        RECT 37.350 142.935 37.490 143.135 ;
        RECT 44.160 143.075 44.480 143.135 ;
        RECT 47.380 143.275 47.700 143.335 ;
        RECT 51.535 143.275 51.825 143.320 ;
        RECT 77.740 143.275 78.060 143.335 ;
        RECT 47.380 143.135 51.825 143.275 ;
        RECT 47.380 143.075 47.700 143.135 ;
        RECT 51.535 143.090 51.825 143.135 ;
        RECT 52.070 143.135 78.060 143.275 ;
        RECT 32.675 142.795 37.490 142.935 ;
        RECT 37.735 142.935 38.025 142.980 ;
        RECT 40.480 142.935 40.800 142.995 ;
        RECT 37.735 142.795 40.800 142.935 ;
        RECT 32.675 142.750 32.965 142.795 ;
        RECT 37.735 142.750 38.025 142.795 ;
        RECT 40.480 142.735 40.800 142.795 ;
        RECT 46.460 142.935 46.780 142.995 ;
        RECT 48.760 142.935 49.080 142.995 ;
        RECT 52.070 142.935 52.210 143.135 ;
        RECT 46.460 142.795 48.070 142.935 ;
        RECT 46.460 142.735 46.780 142.795 ;
        RECT 13.800 142.455 21.390 142.595 ;
        RECT 23.460 142.595 23.780 142.655 ;
        RECT 24.395 142.595 24.685 142.640 ;
        RECT 23.460 142.455 24.685 142.595 ;
        RECT 13.800 142.395 14.120 142.455 ;
        RECT 23.460 142.395 23.780 142.455 ;
        RECT 24.395 142.410 24.685 142.455 ;
        RECT 33.580 142.395 33.900 142.655 ;
        RECT 34.055 142.595 34.345 142.640 ;
        RECT 34.960 142.595 35.280 142.655 ;
        RECT 34.055 142.455 35.280 142.595 ;
        RECT 34.055 142.410 34.345 142.455 ;
        RECT 34.960 142.395 35.280 142.455 ;
        RECT 36.340 142.395 36.660 142.655 ;
        RECT 36.800 142.395 37.120 142.655 ;
        RECT 45.540 142.595 45.860 142.655 ;
        RECT 47.380 142.595 47.700 142.655 ;
        RECT 47.930 142.640 48.070 142.795 ;
        RECT 48.760 142.795 52.210 142.935 ;
        RECT 54.740 142.935 55.060 142.995 ;
        RECT 57.910 142.935 58.200 142.980 ;
        RECT 61.170 142.935 61.460 142.980 ;
        RECT 54.740 142.795 61.460 142.935 ;
        RECT 48.760 142.735 49.080 142.795 ;
        RECT 49.310 142.640 49.450 142.795 ;
        RECT 54.740 142.735 55.060 142.795 ;
        RECT 57.910 142.750 58.200 142.795 ;
        RECT 61.170 142.750 61.460 142.795 ;
        RECT 62.090 142.935 62.380 142.980 ;
        RECT 63.950 142.935 64.240 142.980 ;
        RECT 62.090 142.795 64.240 142.935 ;
        RECT 62.090 142.750 62.380 142.795 ;
        RECT 63.950 142.750 64.240 142.795 ;
        RECT 45.540 142.455 47.700 142.595 ;
        RECT 45.540 142.395 45.860 142.455 ;
        RECT 47.380 142.395 47.700 142.455 ;
        RECT 47.855 142.410 48.145 142.640 ;
        RECT 48.315 142.410 48.605 142.640 ;
        RECT 49.235 142.410 49.525 142.640 ;
        RECT 59.770 142.595 60.060 142.640 ;
        RECT 62.090 142.595 62.305 142.750 ;
        RECT 70.930 142.640 71.070 143.135 ;
        RECT 77.740 143.075 78.060 143.135 ;
        RECT 86.495 143.090 86.785 143.320 ;
        RECT 92.245 143.275 92.535 143.320 ;
        RECT 92.920 143.275 93.240 143.335 ;
        RECT 87.490 143.135 93.240 143.275 ;
        RECT 83.260 142.935 83.580 142.995 ;
        RECT 84.195 142.935 84.485 142.980 ;
        RECT 71.850 142.795 84.485 142.935 ;
        RECT 71.850 142.640 71.990 142.795 ;
        RECT 83.260 142.735 83.580 142.795 ;
        RECT 84.195 142.750 84.485 142.795 ;
        RECT 59.770 142.455 62.305 142.595 ;
        RECT 59.770 142.410 60.060 142.455 ;
        RECT 70.855 142.410 71.145 142.640 ;
        RECT 71.775 142.410 72.065 142.640 ;
        RECT 72.235 142.410 72.525 142.640 ;
        RECT 72.695 142.595 72.985 142.640 ;
        RECT 75.900 142.595 76.220 142.655 ;
        RECT 72.695 142.455 76.220 142.595 ;
        RECT 72.695 142.410 72.985 142.455 ;
        RECT 21.160 142.255 21.480 142.315 ;
        RECT 21.635 142.255 21.925 142.300 ;
        RECT 21.160 142.115 21.925 142.255 ;
        RECT 21.160 142.055 21.480 142.115 ;
        RECT 21.635 142.070 21.925 142.115 ;
        RECT 34.975 141.915 35.265 141.960 ;
        RECT 48.390 141.915 48.530 142.410 ;
        RECT 48.760 142.255 49.080 142.315 ;
        RECT 50.140 142.255 50.460 142.315 ;
        RECT 48.760 142.115 50.460 142.255 ;
        RECT 48.760 142.055 49.080 142.115 ;
        RECT 50.140 142.055 50.460 142.115 ;
        RECT 51.075 142.070 51.365 142.300 ;
        RECT 61.180 142.255 61.500 142.315 ;
        RECT 63.035 142.255 63.325 142.300 ;
        RECT 61.180 142.115 63.325 142.255 ;
        RECT 51.150 141.915 51.290 142.070 ;
        RECT 61.180 142.055 61.500 142.115 ;
        RECT 63.035 142.070 63.325 142.115 ;
        RECT 64.875 142.255 65.165 142.300 ;
        RECT 65.780 142.255 66.100 142.315 ;
        RECT 64.875 142.115 66.100 142.255 ;
        RECT 72.310 142.255 72.450 142.410 ;
        RECT 75.900 142.395 76.220 142.455 ;
        RECT 76.375 142.410 76.665 142.640 ;
        RECT 76.835 142.410 77.125 142.640 ;
        RECT 73.140 142.255 73.460 142.315 ;
        RECT 72.310 142.115 73.460 142.255 ;
        RECT 64.875 142.070 65.165 142.115 ;
        RECT 65.780 142.055 66.100 142.115 ;
        RECT 73.140 142.055 73.460 142.115 ;
        RECT 74.535 142.070 74.825 142.300 ;
        RECT 55.905 141.915 56.195 141.960 ;
        RECT 57.960 141.915 58.280 141.975 ;
        RECT 34.975 141.775 46.690 141.915 ;
        RECT 48.390 141.775 58.280 141.915 ;
        RECT 34.975 141.730 35.265 141.775 ;
        RECT 32.660 141.375 32.980 141.635 ;
        RECT 34.040 141.575 34.360 141.635 ;
        RECT 36.355 141.575 36.645 141.620 ;
        RECT 34.040 141.435 36.645 141.575 ;
        RECT 34.040 141.375 34.360 141.435 ;
        RECT 36.355 141.390 36.645 141.435 ;
        RECT 43.700 141.575 44.020 141.635 ;
        RECT 46.015 141.575 46.305 141.620 ;
        RECT 43.700 141.435 46.305 141.575 ;
        RECT 46.550 141.575 46.690 141.775 ;
        RECT 55.905 141.730 56.195 141.775 ;
        RECT 57.960 141.715 58.280 141.775 ;
        RECT 59.770 141.915 60.060 141.960 ;
        RECT 62.550 141.915 62.840 141.960 ;
        RECT 64.410 141.915 64.700 141.960 ;
        RECT 59.770 141.775 64.700 141.915 ;
        RECT 59.770 141.730 60.060 141.775 ;
        RECT 62.550 141.730 62.840 141.775 ;
        RECT 64.410 141.730 64.700 141.775 ;
        RECT 71.760 141.915 72.080 141.975 ;
        RECT 74.610 141.915 74.750 142.070 ;
        RECT 71.760 141.775 74.750 141.915 ;
        RECT 76.450 141.915 76.590 142.410 ;
        RECT 76.910 142.255 77.050 142.410 ;
        RECT 77.740 142.395 78.060 142.655 ;
        RECT 84.655 142.595 84.945 142.640 ;
        RECT 78.290 142.455 84.945 142.595 ;
        RECT 86.570 142.595 86.710 143.090 ;
        RECT 86.955 142.595 87.245 142.640 ;
        RECT 86.570 142.455 87.245 142.595 ;
        RECT 78.290 142.255 78.430 142.455 ;
        RECT 84.655 142.410 84.945 142.455 ;
        RECT 86.955 142.410 87.245 142.455 ;
        RECT 76.910 142.115 78.430 142.255 ;
        RECT 80.960 142.255 81.280 142.315 ;
        RECT 83.275 142.255 83.565 142.300 ;
        RECT 80.960 142.115 83.565 142.255 ;
        RECT 84.730 142.255 84.870 142.410 ;
        RECT 87.490 142.255 87.630 143.135 ;
        RECT 92.245 143.090 92.535 143.135 ;
        RECT 92.920 143.075 93.240 143.135 ;
        RECT 102.580 143.075 102.900 143.335 ;
        RECT 94.250 142.935 94.540 142.980 ;
        RECT 96.600 142.935 96.920 142.995 ;
        RECT 97.510 142.935 97.800 142.980 ;
        RECT 94.250 142.795 97.800 142.935 ;
        RECT 94.250 142.750 94.540 142.795 ;
        RECT 96.600 142.735 96.920 142.795 ;
        RECT 97.510 142.750 97.800 142.795 ;
        RECT 98.430 142.935 98.720 142.980 ;
        RECT 100.290 142.935 100.580 142.980 ;
        RECT 104.420 142.935 104.740 142.995 ;
        RECT 98.430 142.795 100.580 142.935 ;
        RECT 98.430 142.750 98.720 142.795 ;
        RECT 100.290 142.750 100.580 142.795 ;
        RECT 101.290 142.795 104.740 142.935 ;
        RECT 96.110 142.595 96.400 142.640 ;
        RECT 98.430 142.595 98.645 142.750 ;
        RECT 101.290 142.640 101.430 142.795 ;
        RECT 104.420 142.735 104.740 142.795 ;
        RECT 96.110 142.455 98.645 142.595 ;
        RECT 96.110 142.410 96.400 142.455 ;
        RECT 101.215 142.410 101.505 142.640 ;
        RECT 101.675 142.595 101.965 142.640 ;
        RECT 102.120 142.595 102.440 142.655 ;
        RECT 101.675 142.455 102.440 142.595 ;
        RECT 101.675 142.410 101.965 142.455 ;
        RECT 102.120 142.395 102.440 142.455 ;
        RECT 84.730 142.115 87.630 142.255 ;
        RECT 80.960 142.055 81.280 142.115 ;
        RECT 83.275 142.070 83.565 142.115 ;
        RECT 99.360 142.055 99.680 142.315 ;
        RECT 76.820 141.915 77.140 141.975 ;
        RECT 76.450 141.775 77.140 141.915 ;
        RECT 71.760 141.715 72.080 141.775 ;
        RECT 76.820 141.715 77.140 141.775 ;
        RECT 96.110 141.915 96.400 141.960 ;
        RECT 98.890 141.915 99.180 141.960 ;
        RECT 100.750 141.915 101.040 141.960 ;
        RECT 96.110 141.775 101.040 141.915 ;
        RECT 96.110 141.730 96.400 141.775 ;
        RECT 98.890 141.730 99.180 141.775 ;
        RECT 100.750 141.730 101.040 141.775 ;
        RECT 52.900 141.575 53.220 141.635 ;
        RECT 46.550 141.435 53.220 141.575 ;
        RECT 43.700 141.375 44.020 141.435 ;
        RECT 46.015 141.390 46.305 141.435 ;
        RECT 52.900 141.375 53.220 141.435 ;
        RECT 53.375 141.575 53.665 141.620 ;
        RECT 58.420 141.575 58.740 141.635 ;
        RECT 53.375 141.435 58.740 141.575 ;
        RECT 53.375 141.390 53.665 141.435 ;
        RECT 58.420 141.375 58.740 141.435 ;
        RECT 74.075 141.575 74.365 141.620 ;
        RECT 74.520 141.575 74.840 141.635 ;
        RECT 74.075 141.435 74.840 141.575 ;
        RECT 74.075 141.390 74.365 141.435 ;
        RECT 74.520 141.375 74.840 141.435 ;
        RECT 87.875 141.575 88.165 141.620 ;
        RECT 88.320 141.575 88.640 141.635 ;
        RECT 87.875 141.435 88.640 141.575 ;
        RECT 87.875 141.390 88.165 141.435 ;
        RECT 88.320 141.375 88.640 141.435 ;
        RECT 11.430 140.755 118.610 141.235 ;
        RECT 135.635 141.220 136.775 165.470 ;
        RECT 34.960 140.355 35.280 140.615 ;
        RECT 35.420 140.355 35.740 140.615 ;
        RECT 36.800 140.355 37.120 140.615 ;
        RECT 45.080 140.355 45.400 140.615 ;
        RECT 51.520 140.555 51.840 140.615 ;
        RECT 60.260 140.555 60.580 140.615 ;
        RECT 47.930 140.415 51.840 140.555 ;
        RECT 33.120 140.215 33.440 140.275 ;
        RECT 33.120 140.075 37.030 140.215 ;
        RECT 33.120 140.015 33.440 140.075 ;
        RECT 31.740 139.875 32.060 139.935 ;
        RECT 34.515 139.875 34.805 139.920 ;
        RECT 35.880 139.875 36.200 139.935 ;
        RECT 36.890 139.920 37.030 140.075 ;
        RECT 31.740 139.735 34.270 139.875 ;
        RECT 31.740 139.675 32.060 139.735 ;
        RECT 33.580 139.335 33.900 139.595 ;
        RECT 34.130 139.535 34.270 139.735 ;
        RECT 34.515 139.735 36.200 139.875 ;
        RECT 34.515 139.690 34.805 139.735 ;
        RECT 35.880 139.675 36.200 139.735 ;
        RECT 36.815 139.690 37.105 139.920 ;
        RECT 42.780 139.875 43.100 139.935 ;
        RECT 45.095 139.875 45.385 139.920 ;
        RECT 42.780 139.735 45.385 139.875 ;
        RECT 42.780 139.675 43.100 139.735 ;
        RECT 45.095 139.690 45.385 139.735 ;
        RECT 46.460 139.875 46.780 139.935 ;
        RECT 47.930 139.875 48.070 140.415 ;
        RECT 51.520 140.355 51.840 140.415 ;
        RECT 59.200 140.415 60.580 140.555 ;
        RECT 50.140 140.215 50.460 140.275 ;
        RECT 59.200 140.215 59.340 140.415 ;
        RECT 60.260 140.355 60.580 140.415 ;
        RECT 61.180 140.355 61.500 140.615 ;
        RECT 62.575 140.555 62.865 140.600 ;
        RECT 63.020 140.555 63.340 140.615 ;
        RECT 62.575 140.415 63.340 140.555 ;
        RECT 62.575 140.370 62.865 140.415 ;
        RECT 63.020 140.355 63.340 140.415 ;
        RECT 70.840 140.355 71.160 140.615 ;
        RECT 73.140 140.355 73.460 140.615 ;
        RECT 81.205 140.555 81.495 140.600 ;
        RECT 83.260 140.555 83.580 140.615 ;
        RECT 81.205 140.415 83.580 140.555 ;
        RECT 81.205 140.370 81.495 140.415 ;
        RECT 83.260 140.355 83.580 140.415 ;
        RECT 96.155 140.555 96.445 140.600 ;
        RECT 96.600 140.555 96.920 140.615 ;
        RECT 96.155 140.415 96.920 140.555 ;
        RECT 96.155 140.370 96.445 140.415 ;
        RECT 96.600 140.355 96.920 140.415 ;
        RECT 98.915 140.555 99.205 140.600 ;
        RECT 99.360 140.555 99.680 140.615 ;
        RECT 98.915 140.415 99.680 140.555 ;
        RECT 98.915 140.370 99.205 140.415 ;
        RECT 99.360 140.355 99.680 140.415 ;
        RECT 50.140 140.075 59.340 140.215 ;
        RECT 50.140 140.015 50.460 140.075 ;
        RECT 56.670 139.920 56.810 140.075 ;
        RECT 59.815 140.030 60.105 140.260 ;
        RECT 75.440 140.215 75.760 140.275 ;
        RECT 73.230 140.075 75.760 140.215 ;
        RECT 46.460 139.735 48.070 139.875 ;
        RECT 46.460 139.675 46.780 139.735 ;
        RECT 36.355 139.535 36.645 139.580 ;
        RECT 34.130 139.395 36.645 139.535 ;
        RECT 36.355 139.350 36.645 139.395 ;
        RECT 37.735 139.535 38.025 139.580 ;
        RECT 43.700 139.535 44.020 139.595 ;
        RECT 37.735 139.395 44.020 139.535 ;
        RECT 37.735 139.350 38.025 139.395 ;
        RECT 43.700 139.335 44.020 139.395 ;
        RECT 44.175 139.535 44.465 139.580 ;
        RECT 44.620 139.535 44.940 139.595 ;
        RECT 44.175 139.395 44.940 139.535 ;
        RECT 44.175 139.350 44.465 139.395 ;
        RECT 44.620 139.335 44.940 139.395 ;
        RECT 47.380 139.335 47.700 139.595 ;
        RECT 47.930 139.580 48.070 139.735 ;
        RECT 48.390 139.735 55.430 139.875 ;
        RECT 48.390 139.580 48.530 139.735 ;
        RECT 47.855 139.350 48.145 139.580 ;
        RECT 48.315 139.350 48.605 139.580 ;
        RECT 49.220 139.535 49.540 139.595 ;
        RECT 49.220 139.395 50.830 139.535 ;
        RECT 49.220 139.335 49.540 139.395 ;
        RECT 34.975 139.195 35.265 139.240 ;
        RECT 45.555 139.195 45.845 139.240 ;
        RECT 49.695 139.195 49.985 139.240 ;
        RECT 34.975 139.055 44.390 139.195 ;
        RECT 34.975 139.010 35.265 139.055 ;
        RECT 32.675 138.855 32.965 138.900 ;
        RECT 41.860 138.855 42.180 138.915 ;
        RECT 32.675 138.715 42.180 138.855 ;
        RECT 32.675 138.670 32.965 138.715 ;
        RECT 41.860 138.655 42.180 138.715 ;
        RECT 43.255 138.855 43.545 138.900 ;
        RECT 43.700 138.855 44.020 138.915 ;
        RECT 43.255 138.715 44.020 138.855 ;
        RECT 44.250 138.855 44.390 139.055 ;
        RECT 45.555 139.055 49.985 139.195 ;
        RECT 45.555 139.010 45.845 139.055 ;
        RECT 49.695 139.010 49.985 139.055 ;
        RECT 46.015 138.855 46.305 138.900 ;
        RECT 44.250 138.715 46.305 138.855 ;
        RECT 50.690 138.855 50.830 139.395 ;
        RECT 51.060 139.335 51.380 139.595 ;
        RECT 51.520 139.335 51.840 139.595 ;
        RECT 51.995 139.350 52.285 139.580 ;
        RECT 52.440 139.535 52.760 139.595 ;
        RECT 52.915 139.535 53.205 139.580 ;
        RECT 52.440 139.395 53.205 139.535 ;
        RECT 55.290 139.535 55.430 139.735 ;
        RECT 56.595 139.690 56.885 139.920 ;
        RECT 59.890 139.875 60.030 140.030 ;
        RECT 59.890 139.735 61.870 139.875 ;
        RECT 57.500 139.535 57.820 139.595 ;
        RECT 55.290 139.395 57.820 139.535 ;
        RECT 52.070 139.195 52.210 139.350 ;
        RECT 52.440 139.335 52.760 139.395 ;
        RECT 52.915 139.350 53.205 139.395 ;
        RECT 57.500 139.335 57.820 139.395 ;
        RECT 57.960 139.335 58.280 139.595 ;
        RECT 58.420 139.535 58.740 139.595 ;
        RECT 61.730 139.580 61.870 139.735 ;
        RECT 60.275 139.535 60.565 139.580 ;
        RECT 58.420 139.395 60.565 139.535 ;
        RECT 58.420 139.335 58.740 139.395 ;
        RECT 60.275 139.350 60.565 139.395 ;
        RECT 61.655 139.350 61.945 139.580 ;
        RECT 70.380 139.335 70.700 139.595 ;
        RECT 70.855 139.350 71.145 139.580 ;
        RECT 59.800 139.195 60.120 139.255 ;
        RECT 52.070 139.055 60.120 139.195 ;
        RECT 70.930 139.195 71.070 139.350 ;
        RECT 71.760 139.335 72.080 139.595 ;
        RECT 73.230 139.580 73.370 140.075 ;
        RECT 75.440 140.015 75.760 140.075 ;
        RECT 85.070 140.215 85.360 140.260 ;
        RECT 87.850 140.215 88.140 140.260 ;
        RECT 89.710 140.215 90.000 140.260 ;
        RECT 135.580 140.230 136.830 141.220 ;
        RECT 85.070 140.075 90.000 140.215 ;
        RECT 135.635 140.155 136.775 140.230 ;
        RECT 85.070 140.030 85.360 140.075 ;
        RECT 87.850 140.030 88.140 140.075 ;
        RECT 89.710 140.030 90.000 140.075 ;
        RECT 74.075 139.875 74.365 139.920 ;
        RECT 74.980 139.875 75.300 139.935 ;
        RECT 74.075 139.735 75.300 139.875 ;
        RECT 74.075 139.690 74.365 139.735 ;
        RECT 74.980 139.675 75.300 139.735 ;
        RECT 88.320 139.675 88.640 139.935 ;
        RECT 89.240 139.875 89.560 139.935 ;
        RECT 90.175 139.875 90.465 139.920 ;
        RECT 89.240 139.735 90.465 139.875 ;
        RECT 89.240 139.675 89.560 139.735 ;
        RECT 90.175 139.690 90.465 139.735 ;
        RECT 93.840 139.875 94.160 139.935 ;
        RECT 93.840 139.735 109.710 139.875 ;
        RECT 93.840 139.675 94.160 139.735 ;
        RECT 73.155 139.350 73.445 139.580 ;
        RECT 74.520 139.335 74.840 139.595 ;
        RECT 96.690 139.580 96.830 139.735 ;
        RECT 109.570 139.595 109.710 139.735 ;
        RECT 85.070 139.535 85.360 139.580 ;
        RECT 85.070 139.395 87.605 139.535 ;
        RECT 85.070 139.350 85.360 139.395 ;
        RECT 76.360 139.195 76.680 139.255 ;
        RECT 86.480 139.240 86.800 139.255 ;
        RECT 70.930 139.055 76.680 139.195 ;
        RECT 59.800 138.995 60.120 139.055 ;
        RECT 76.360 138.995 76.680 139.055 ;
        RECT 83.210 139.195 83.500 139.240 ;
        RECT 86.470 139.195 86.800 139.240 ;
        RECT 83.210 139.055 86.800 139.195 ;
        RECT 83.210 139.010 83.500 139.055 ;
        RECT 86.470 139.010 86.800 139.055 ;
        RECT 87.390 139.240 87.605 139.395 ;
        RECT 96.615 139.350 96.905 139.580 ;
        RECT 97.980 139.335 98.300 139.595 ;
        RECT 109.480 139.335 109.800 139.595 ;
        RECT 110.860 139.335 111.180 139.595 ;
        RECT 87.390 139.195 87.680 139.240 ;
        RECT 89.250 139.195 89.540 139.240 ;
        RECT 87.390 139.055 89.540 139.195 ;
        RECT 87.390 139.010 87.680 139.055 ;
        RECT 89.250 139.010 89.540 139.055 ;
        RECT 132.510 139.190 135.210 140.010 ;
        RECT 143.370 139.390 144.510 223.840 ;
        RECT 137.240 139.380 144.510 139.390 ;
        RECT 136.210 139.190 144.510 139.380 ;
        RECT 86.480 138.995 86.800 139.010 ;
        RECT 51.980 138.855 52.300 138.915 ;
        RECT 50.690 138.715 52.300 138.855 ;
        RECT 43.255 138.670 43.545 138.715 ;
        RECT 43.700 138.655 44.020 138.715 ;
        RECT 46.015 138.670 46.305 138.715 ;
        RECT 51.980 138.655 52.300 138.715 ;
        RECT 69.475 138.855 69.765 138.900 ;
        RECT 70.380 138.855 70.700 138.915 ;
        RECT 69.475 138.715 70.700 138.855 ;
        RECT 69.475 138.670 69.765 138.715 ;
        RECT 70.380 138.655 70.700 138.715 ;
        RECT 72.235 138.855 72.525 138.900 ;
        RECT 75.900 138.855 76.220 138.915 ;
        RECT 72.235 138.715 76.220 138.855 ;
        RECT 72.235 138.670 72.525 138.715 ;
        RECT 75.900 138.655 76.220 138.715 ;
        RECT 109.940 138.655 110.260 138.915 ;
        RECT 111.795 138.855 112.085 138.900 ;
        RECT 113.620 138.855 113.940 138.915 ;
        RECT 111.795 138.715 113.940 138.855 ;
        RECT 111.795 138.670 112.085 138.715 ;
        RECT 113.620 138.655 113.940 138.715 ;
        RECT 132.510 138.530 144.510 139.190 ;
        RECT 10.650 138.035 118.610 138.515 ;
        RECT 132.510 138.190 135.210 138.530 ;
        RECT 136.210 138.250 144.510 138.530 ;
        RECT 136.210 138.240 138.350 138.250 ;
        RECT 31.755 137.835 32.045 137.880 ;
        RECT 32.660 137.835 32.980 137.895 ;
        RECT 31.755 137.695 32.980 137.835 ;
        RECT 31.755 137.650 32.045 137.695 ;
        RECT 32.660 137.635 32.980 137.695 ;
        RECT 34.040 137.635 34.360 137.895 ;
        RECT 34.500 137.635 34.820 137.895 ;
        RECT 36.800 137.835 37.120 137.895 ;
        RECT 38.655 137.835 38.945 137.880 ;
        RECT 36.800 137.695 38.945 137.835 ;
        RECT 36.800 137.635 37.120 137.695 ;
        RECT 38.655 137.650 38.945 137.695 ;
        RECT 57.500 137.835 57.820 137.895 ;
        RECT 59.355 137.835 59.645 137.880 ;
        RECT 57.500 137.695 59.645 137.835 ;
        RECT 57.500 137.635 57.820 137.695 ;
        RECT 59.355 137.650 59.645 137.695 ;
        RECT 61.195 137.650 61.485 137.880 ;
        RECT 71.300 137.835 71.620 137.895 ;
        RECT 72.235 137.835 72.525 137.880 ;
        RECT 71.300 137.695 72.525 137.835 ;
        RECT 14.260 137.495 14.580 137.555 ;
        RECT 15.590 137.495 15.880 137.540 ;
        RECT 18.850 137.495 19.140 137.540 ;
        RECT 14.260 137.355 19.140 137.495 ;
        RECT 14.260 137.295 14.580 137.355 ;
        RECT 15.590 137.310 15.880 137.355 ;
        RECT 18.850 137.310 19.140 137.355 ;
        RECT 19.770 137.495 20.060 137.540 ;
        RECT 21.630 137.495 21.920 137.540 ;
        RECT 19.770 137.355 21.920 137.495 ;
        RECT 19.770 137.310 20.060 137.355 ;
        RECT 21.630 137.310 21.920 137.355 ;
        RECT 35.510 137.355 37.950 137.495 ;
        RECT 17.450 137.155 17.740 137.200 ;
        RECT 19.770 137.155 19.985 137.310 ;
        RECT 17.450 137.015 19.985 137.155 ;
        RECT 22.555 137.155 22.845 137.200 ;
        RECT 26.680 137.155 27.000 137.215 ;
        RECT 22.555 137.015 27.000 137.155 ;
        RECT 17.450 136.970 17.740 137.015 ;
        RECT 22.555 136.970 22.845 137.015 ;
        RECT 26.680 136.955 27.000 137.015 ;
        RECT 27.155 137.155 27.445 137.200 ;
        RECT 28.060 137.155 28.380 137.215 ;
        RECT 35.510 137.200 35.650 137.355 ;
        RECT 37.810 137.215 37.950 137.355 ;
        RECT 27.155 137.015 28.380 137.155 ;
        RECT 27.155 136.970 27.445 137.015 ;
        RECT 28.060 136.955 28.380 137.015 ;
        RECT 30.835 137.155 31.125 137.200 ;
        RECT 33.135 137.155 33.425 137.200 ;
        RECT 35.435 137.155 35.725 137.200 ;
        RECT 30.835 137.015 35.725 137.155 ;
        RECT 30.835 136.970 31.125 137.015 ;
        RECT 33.135 136.970 33.425 137.015 ;
        RECT 35.435 136.970 35.725 137.015 ;
        RECT 35.880 136.955 36.200 137.215 ;
        RECT 37.720 136.955 38.040 137.215 ;
        RECT 58.895 137.155 59.185 137.200 ;
        RECT 59.800 137.155 60.120 137.215 ;
        RECT 58.895 137.015 60.120 137.155 ;
        RECT 61.270 137.155 61.410 137.650 ;
        RECT 71.300 137.635 71.620 137.695 ;
        RECT 72.235 137.650 72.525 137.695 ;
        RECT 72.680 137.635 73.000 137.895 ;
        RECT 86.035 137.835 86.325 137.880 ;
        RECT 86.480 137.835 86.800 137.895 ;
        RECT 86.035 137.695 86.800 137.835 ;
        RECT 86.035 137.650 86.325 137.695 ;
        RECT 86.480 137.635 86.800 137.695 ;
        RECT 97.060 137.635 97.380 137.895 ;
        RECT 99.820 137.835 100.140 137.895 ;
        RECT 102.135 137.835 102.425 137.880 ;
        RECT 99.820 137.695 102.425 137.835 ;
        RECT 99.820 137.635 100.140 137.695 ;
        RECT 102.135 137.650 102.425 137.695 ;
        RECT 63.480 137.495 63.800 137.555 ;
        RECT 66.255 137.495 66.545 137.540 ;
        RECT 80.040 137.495 80.360 137.555 ;
        RECT 92.015 137.495 92.305 137.540 ;
        RECT 63.480 137.355 66.545 137.495 ;
        RECT 63.480 137.295 63.800 137.355 ;
        RECT 64.490 137.200 64.630 137.355 ;
        RECT 66.255 137.310 66.545 137.355 ;
        RECT 70.930 137.355 92.305 137.495 ;
        RECT 70.930 137.200 71.070 137.355 ;
        RECT 80.040 137.295 80.360 137.355 ;
        RECT 92.015 137.310 92.305 137.355 ;
        RECT 92.475 137.495 92.765 137.540 ;
        RECT 108.510 137.495 108.800 137.540 ;
        RECT 109.940 137.495 110.260 137.555 ;
        RECT 111.770 137.495 112.060 137.540 ;
        RECT 92.475 137.355 98.670 137.495 ;
        RECT 92.475 137.310 92.765 137.355 ;
        RECT 62.575 137.155 62.865 137.200 ;
        RECT 64.415 137.155 64.705 137.200 ;
        RECT 61.270 137.015 62.865 137.155 ;
        RECT 64.305 137.015 64.705 137.155 ;
        RECT 58.895 136.970 59.185 137.015 ;
        RECT 59.800 136.955 60.120 137.015 ;
        RECT 62.575 136.970 62.865 137.015 ;
        RECT 64.415 136.970 64.705 137.015 ;
        RECT 70.855 136.970 71.145 137.200 ;
        RECT 71.315 137.155 71.605 137.200 ;
        RECT 73.615 137.155 73.905 137.200 ;
        RECT 71.315 137.015 73.905 137.155 ;
        RECT 71.315 136.970 71.605 137.015 ;
        RECT 73.615 136.970 73.905 137.015 ;
        RECT 81.880 137.155 82.200 137.215 ;
        RECT 84.195 137.155 84.485 137.200 ;
        RECT 81.880 137.015 84.485 137.155 ;
        RECT 17.940 136.815 18.260 136.875 ;
        RECT 20.715 136.815 21.005 136.860 ;
        RECT 17.940 136.675 21.005 136.815 ;
        RECT 17.940 136.615 18.260 136.675 ;
        RECT 20.715 136.630 21.005 136.675 ;
        RECT 21.160 136.815 21.480 136.875 ;
        RECT 29.915 136.815 30.205 136.860 ;
        RECT 21.160 136.675 30.205 136.815 ;
        RECT 21.160 136.615 21.480 136.675 ;
        RECT 29.915 136.630 30.205 136.675 ;
        RECT 30.360 136.815 30.680 136.875 ;
        RECT 32.215 136.815 32.505 136.860 ;
        RECT 30.360 136.675 32.505 136.815 ;
        RECT 30.360 136.615 30.680 136.675 ;
        RECT 32.215 136.630 32.505 136.675 ;
        RECT 36.815 136.630 37.105 136.860 ;
        RECT 58.435 136.815 58.725 136.860 ;
        RECT 60.260 136.815 60.580 136.875 ;
        RECT 71.390 136.815 71.530 136.970 ;
        RECT 81.880 136.955 82.200 137.015 ;
        RECT 84.195 136.970 84.485 137.015 ;
        RECT 86.495 137.155 86.785 137.200 ;
        RECT 93.840 137.155 94.160 137.215 ;
        RECT 98.530 137.200 98.670 137.355 ;
        RECT 108.510 137.355 112.060 137.495 ;
        RECT 108.510 137.310 108.800 137.355 ;
        RECT 109.940 137.295 110.260 137.355 ;
        RECT 111.770 137.310 112.060 137.355 ;
        RECT 112.690 137.495 112.980 137.540 ;
        RECT 114.550 137.495 114.840 137.540 ;
        RECT 112.690 137.355 114.840 137.495 ;
        RECT 112.690 137.310 112.980 137.355 ;
        RECT 114.550 137.310 114.840 137.355 ;
        RECT 96.615 137.155 96.905 137.200 ;
        RECT 86.495 137.015 94.160 137.155 ;
        RECT 86.495 136.970 86.785 137.015 ;
        RECT 93.840 136.955 94.160 137.015 ;
        RECT 94.390 137.015 96.905 137.155 ;
        RECT 58.435 136.675 60.580 136.815 ;
        RECT 58.435 136.630 58.725 136.675 ;
        RECT 17.450 136.475 17.740 136.520 ;
        RECT 20.230 136.475 20.520 136.520 ;
        RECT 22.090 136.475 22.380 136.520 ;
        RECT 17.450 136.335 22.380 136.475 ;
        RECT 17.450 136.290 17.740 136.335 ;
        RECT 20.230 136.290 20.520 136.335 ;
        RECT 22.090 136.290 22.380 136.335 ;
        RECT 26.680 136.475 27.000 136.535 ;
        RECT 36.890 136.475 37.030 136.630 ;
        RECT 60.260 136.615 60.580 136.675 ;
        RECT 67.250 136.675 71.530 136.815 ;
        RECT 74.535 136.815 74.825 136.860 ;
        RECT 75.440 136.815 75.760 136.875 ;
        RECT 74.535 136.675 75.760 136.815 ;
        RECT 26.680 136.335 37.030 136.475 ;
        RECT 26.680 136.275 27.000 136.335 ;
        RECT 67.250 136.195 67.390 136.675 ;
        RECT 74.535 136.630 74.825 136.675 ;
        RECT 75.440 136.615 75.760 136.675 ;
        RECT 91.555 136.815 91.845 136.860 ;
        RECT 93.380 136.815 93.700 136.875 ;
        RECT 91.555 136.675 93.700 136.815 ;
        RECT 91.555 136.630 91.845 136.675 ;
        RECT 93.380 136.615 93.700 136.675 ;
        RECT 94.390 136.520 94.530 137.015 ;
        RECT 96.615 136.970 96.905 137.015 ;
        RECT 97.995 136.970 98.285 137.200 ;
        RECT 98.455 137.155 98.745 137.200 ;
        RECT 99.360 137.155 99.680 137.215 ;
        RECT 98.455 137.015 99.680 137.155 ;
        RECT 98.455 136.970 98.745 137.015 ;
        RECT 98.070 136.815 98.210 136.970 ;
        RECT 99.360 136.955 99.680 137.015 ;
        RECT 102.580 137.155 102.900 137.215 ;
        RECT 103.055 137.155 103.345 137.200 ;
        RECT 102.580 137.015 103.345 137.155 ;
        RECT 102.580 136.955 102.900 137.015 ;
        RECT 103.055 136.970 103.345 137.015 ;
        RECT 110.370 137.155 110.660 137.200 ;
        RECT 112.690 137.155 112.905 137.310 ;
        RECT 110.370 137.015 112.905 137.155 ;
        RECT 110.370 136.970 110.660 137.015 ;
        RECT 113.620 136.955 113.940 137.215 ;
        RECT 102.670 136.815 102.810 136.955 ;
        RECT 106.260 136.860 106.580 136.875 ;
        RECT 98.070 136.675 102.810 136.815 ;
        RECT 103.975 136.815 104.265 136.860 ;
        RECT 106.260 136.815 106.795 136.860 ;
        RECT 103.975 136.675 106.795 136.815 ;
        RECT 103.975 136.630 104.265 136.675 ;
        RECT 106.260 136.630 106.795 136.675 ;
        RECT 106.260 136.615 106.580 136.630 ;
        RECT 115.460 136.615 115.780 136.875 ;
        RECT 94.315 136.290 94.605 136.520 ;
        RECT 110.370 136.475 110.660 136.520 ;
        RECT 113.150 136.475 113.440 136.520 ;
        RECT 115.010 136.475 115.300 136.520 ;
        RECT 110.370 136.335 115.300 136.475 ;
        RECT 110.370 136.290 110.660 136.335 ;
        RECT 113.150 136.290 113.440 136.335 ;
        RECT 115.010 136.290 115.300 136.335 ;
        RECT 13.585 136.135 13.875 136.180 ;
        RECT 21.160 136.135 21.480 136.195 ;
        RECT 13.585 135.995 21.480 136.135 ;
        RECT 13.585 135.950 13.875 135.995 ;
        RECT 21.160 135.935 21.480 135.995 ;
        RECT 25.760 136.135 26.080 136.195 ;
        RECT 26.235 136.135 26.525 136.180 ;
        RECT 25.760 135.995 26.525 136.135 ;
        RECT 25.760 135.935 26.080 135.995 ;
        RECT 26.235 135.950 26.525 135.995 ;
        RECT 63.495 136.135 63.785 136.180 ;
        RECT 64.400 136.135 64.720 136.195 ;
        RECT 63.495 135.995 64.720 136.135 ;
        RECT 63.495 135.950 63.785 135.995 ;
        RECT 64.400 135.935 64.720 135.995 ;
        RECT 65.335 136.135 65.625 136.180 ;
        RECT 65.780 136.135 66.100 136.195 ;
        RECT 65.335 135.995 66.100 136.135 ;
        RECT 65.335 135.950 65.625 135.995 ;
        RECT 65.780 135.935 66.100 135.995 ;
        RECT 66.715 136.135 67.005 136.180 ;
        RECT 67.160 136.135 67.480 136.195 ;
        RECT 66.715 135.995 67.480 136.135 ;
        RECT 66.715 135.950 67.005 135.995 ;
        RECT 67.160 135.935 67.480 135.995 ;
        RECT 83.735 136.135 84.025 136.180 ;
        RECT 84.180 136.135 84.500 136.195 ;
        RECT 83.735 135.995 84.500 136.135 ;
        RECT 83.735 135.950 84.025 135.995 ;
        RECT 84.180 135.935 84.500 135.995 ;
        RECT 94.760 136.135 95.080 136.195 ;
        RECT 95.695 136.135 95.985 136.180 ;
        RECT 94.760 135.995 95.985 136.135 ;
        RECT 94.760 135.935 95.080 135.995 ;
        RECT 95.695 135.950 95.985 135.995 ;
        RECT 11.430 135.315 118.610 135.795 ;
        RECT 14.260 134.915 14.580 135.175 ;
        RECT 17.940 134.915 18.260 135.175 ;
        RECT 28.060 134.915 28.380 135.175 ;
        RECT 40.940 135.115 41.260 135.175 ;
        RECT 57.285 135.115 57.575 135.160 ;
        RECT 59.800 135.115 60.120 135.175 ;
        RECT 69.460 135.115 69.780 135.175 ;
        RECT 40.940 134.975 47.150 135.115 ;
        RECT 40.940 134.915 41.260 134.975 ;
        RECT 22.510 134.775 22.800 134.820 ;
        RECT 25.290 134.775 25.580 134.820 ;
        RECT 27.150 134.775 27.440 134.820 ;
        RECT 22.510 134.635 27.440 134.775 ;
        RECT 22.510 134.590 22.800 134.635 ;
        RECT 25.290 134.590 25.580 134.635 ;
        RECT 27.150 134.590 27.440 134.635 ;
        RECT 36.340 134.775 36.660 134.835 ;
        RECT 37.720 134.775 38.040 134.835 ;
        RECT 47.010 134.775 47.150 134.975 ;
        RECT 57.285 134.975 60.120 135.115 ;
        RECT 57.285 134.930 57.575 134.975 ;
        RECT 59.800 134.915 60.120 134.975 ;
        RECT 60.810 134.975 69.780 135.115 ;
        RECT 60.810 134.775 60.950 134.975 ;
        RECT 69.460 134.915 69.780 134.975 ;
        RECT 70.840 134.915 71.160 135.175 ;
        RECT 73.140 134.915 73.460 135.175 ;
        RECT 108.115 135.115 108.405 135.160 ;
        RECT 110.860 135.115 111.180 135.175 ;
        RECT 108.115 134.975 111.180 135.115 ;
        RECT 108.115 134.930 108.405 134.975 ;
        RECT 110.860 134.915 111.180 134.975 ;
        RECT 36.340 134.635 46.690 134.775 ;
        RECT 47.010 134.635 60.950 134.775 ;
        RECT 61.150 134.775 61.440 134.820 ;
        RECT 63.930 134.775 64.220 134.820 ;
        RECT 65.790 134.775 66.080 134.820 ;
        RECT 61.150 134.635 66.080 134.775 ;
        RECT 36.340 134.575 36.660 134.635 ;
        RECT 37.720 134.575 38.040 134.635 ;
        RECT 25.760 134.235 26.080 134.495 ;
        RECT 31.280 134.435 31.600 134.495 ;
        RECT 33.135 134.435 33.425 134.480 ;
        RECT 31.280 134.295 33.425 134.435 ;
        RECT 31.280 134.235 31.600 134.295 ;
        RECT 33.135 134.250 33.425 134.295 ;
        RECT 38.270 134.295 40.250 134.435 ;
        RECT 14.720 134.095 15.040 134.155 ;
        RECT 15.655 134.095 15.945 134.140 ;
        RECT 14.720 133.955 15.945 134.095 ;
        RECT 14.720 133.895 15.040 133.955 ;
        RECT 15.655 133.910 15.945 133.955 ;
        RECT 17.035 134.095 17.325 134.140 ;
        RECT 18.400 134.095 18.720 134.155 ;
        RECT 17.035 133.955 18.720 134.095 ;
        RECT 17.035 133.910 17.325 133.955 ;
        RECT 18.400 133.895 18.720 133.955 ;
        RECT 22.510 134.095 22.800 134.140 ;
        RECT 27.140 134.095 27.460 134.155 ;
        RECT 27.615 134.095 27.905 134.140 ;
        RECT 22.510 133.955 25.045 134.095 ;
        RECT 22.510 133.910 22.800 133.955 ;
        RECT 24.830 133.800 25.045 133.955 ;
        RECT 27.140 133.955 27.905 134.095 ;
        RECT 27.140 133.895 27.460 133.955 ;
        RECT 27.615 133.910 27.905 133.955 ;
        RECT 29.915 134.095 30.205 134.140 ;
        RECT 30.360 134.095 30.680 134.155 ;
        RECT 38.270 134.095 38.410 134.295 ;
        RECT 29.915 133.955 30.680 134.095 ;
        RECT 29.915 133.910 30.205 133.955 ;
        RECT 30.360 133.895 30.680 133.955 ;
        RECT 36.890 133.955 38.410 134.095 ;
        RECT 38.655 134.095 38.945 134.140 ;
        RECT 39.100 134.095 39.420 134.155 ;
        RECT 38.655 133.955 39.420 134.095 ;
        RECT 36.890 133.815 37.030 133.955 ;
        RECT 38.655 133.910 38.945 133.955 ;
        RECT 39.100 133.895 39.420 133.955 ;
        RECT 39.575 133.910 39.865 134.140 ;
        RECT 16.115 133.755 16.405 133.800 ;
        RECT 20.650 133.755 20.940 133.800 ;
        RECT 23.910 133.755 24.200 133.800 ;
        RECT 16.115 133.615 24.200 133.755 ;
        RECT 16.115 133.570 16.405 133.615 ;
        RECT 20.650 133.570 20.940 133.615 ;
        RECT 23.910 133.570 24.200 133.615 ;
        RECT 24.830 133.755 25.120 133.800 ;
        RECT 26.690 133.755 26.980 133.800 ;
        RECT 24.830 133.615 26.980 133.755 ;
        RECT 24.830 133.570 25.120 133.615 ;
        RECT 26.690 133.570 26.980 133.615 ;
        RECT 34.055 133.755 34.345 133.800 ;
        RECT 36.800 133.755 37.120 133.815 ;
        RECT 34.055 133.615 37.120 133.755 ;
        RECT 34.055 133.570 34.345 133.615 ;
        RECT 36.800 133.555 37.120 133.615 ;
        RECT 18.860 133.460 19.180 133.475 ;
        RECT 18.645 133.230 19.180 133.460 ;
        RECT 30.375 133.415 30.665 133.460 ;
        RECT 31.740 133.415 32.060 133.475 ;
        RECT 34.515 133.415 34.805 133.460 ;
        RECT 35.880 133.415 36.200 133.475 ;
        RECT 30.375 133.275 36.200 133.415 ;
        RECT 30.375 133.230 30.665 133.275 ;
        RECT 18.860 133.215 19.180 133.230 ;
        RECT 31.740 133.215 32.060 133.275 ;
        RECT 34.515 133.230 34.805 133.275 ;
        RECT 35.880 133.215 36.200 133.275 ;
        RECT 36.355 133.415 36.645 133.460 ;
        RECT 39.100 133.415 39.420 133.475 ;
        RECT 36.355 133.275 39.420 133.415 ;
        RECT 39.650 133.415 39.790 133.910 ;
        RECT 40.110 133.755 40.250 134.295 ;
        RECT 40.480 134.235 40.800 134.495 ;
        RECT 41.875 133.910 42.165 134.140 ;
        RECT 42.335 133.910 42.625 134.140 ;
        RECT 41.950 133.755 42.090 133.910 ;
        RECT 40.110 133.615 42.090 133.755 ;
        RECT 42.410 133.755 42.550 133.910 ;
        RECT 43.240 133.895 43.560 134.155 ;
        RECT 44.160 133.895 44.480 134.155 ;
        RECT 44.620 133.895 44.940 134.155 ;
        RECT 45.080 134.095 45.400 134.155 ;
        RECT 46.015 134.095 46.305 134.140 ;
        RECT 45.080 133.955 46.305 134.095 ;
        RECT 46.550 134.095 46.690 134.635 ;
        RECT 61.150 134.590 61.440 134.635 ;
        RECT 63.930 134.590 64.220 134.635 ;
        RECT 65.790 134.590 66.080 134.635 ;
        RECT 83.690 134.775 83.980 134.820 ;
        RECT 86.470 134.775 86.760 134.820 ;
        RECT 88.330 134.775 88.620 134.820 ;
        RECT 83.690 134.635 88.620 134.775 ;
        RECT 83.690 134.590 83.980 134.635 ;
        RECT 86.470 134.590 86.760 134.635 ;
        RECT 88.330 134.590 88.620 134.635 ;
        RECT 93.400 134.775 93.690 134.820 ;
        RECT 95.260 134.775 95.550 134.820 ;
        RECT 98.040 134.775 98.330 134.820 ;
        RECT 93.400 134.635 98.330 134.775 ;
        RECT 93.400 134.590 93.690 134.635 ;
        RECT 95.260 134.590 95.550 134.635 ;
        RECT 98.040 134.590 98.330 134.635 ;
        RECT 47.380 134.435 47.700 134.495 ;
        RECT 47.855 134.435 48.145 134.480 ;
        RECT 47.380 134.295 48.145 134.435 ;
        RECT 47.380 134.235 47.700 134.295 ;
        RECT 47.855 134.250 48.145 134.295 ;
        RECT 60.720 134.235 61.040 134.495 ;
        RECT 64.400 134.235 64.720 134.495 ;
        RECT 72.695 134.435 72.985 134.480 ;
        RECT 72.695 134.295 74.750 134.435 ;
        RECT 72.695 134.250 72.985 134.295 ;
        RECT 46.935 134.095 47.225 134.140 ;
        RECT 56.595 134.095 56.885 134.140 ;
        RECT 60.810 134.095 60.950 134.235 ;
        RECT 74.610 134.155 74.750 134.295 ;
        RECT 76.360 134.235 76.680 134.495 ;
        RECT 88.795 134.435 89.085 134.480 ;
        RECT 89.240 134.435 89.560 134.495 ;
        RECT 92.935 134.435 93.225 134.480 ;
        RECT 88.795 134.295 93.225 134.435 ;
        RECT 88.795 134.250 89.085 134.295 ;
        RECT 89.240 134.235 89.560 134.295 ;
        RECT 92.935 134.250 93.225 134.295 ;
        RECT 93.840 134.235 94.160 134.495 ;
        RECT 94.760 134.235 95.080 134.495 ;
        RECT 105.355 134.435 105.645 134.480 ;
        RECT 107.640 134.435 107.960 134.495 ;
        RECT 135.660 134.480 136.800 134.510 ;
        RECT 109.035 134.435 109.325 134.480 ;
        RECT 95.310 134.295 109.325 134.435 ;
        RECT 46.550 133.955 48.530 134.095 ;
        RECT 45.080 133.895 45.400 133.955 ;
        RECT 46.015 133.910 46.305 133.955 ;
        RECT 46.935 133.910 47.225 133.955 ;
        RECT 44.710 133.755 44.850 133.895 ;
        RECT 42.410 133.615 44.850 133.755 ;
        RECT 45.555 133.755 45.845 133.800 ;
        RECT 47.840 133.755 48.160 133.815 ;
        RECT 45.555 133.615 48.160 133.755 ;
        RECT 42.410 133.415 42.550 133.615 ;
        RECT 45.555 133.570 45.845 133.615 ;
        RECT 47.840 133.555 48.160 133.615 ;
        RECT 39.650 133.275 42.550 133.415 ;
        RECT 48.390 133.415 48.530 133.955 ;
        RECT 56.595 133.955 60.950 134.095 ;
        RECT 61.150 134.095 61.440 134.140 ;
        RECT 61.150 133.955 63.685 134.095 ;
        RECT 56.595 133.910 56.885 133.955 ;
        RECT 61.150 133.910 61.440 133.955 ;
        RECT 63.470 133.800 63.685 133.955 ;
        RECT 66.240 133.895 66.560 134.155 ;
        RECT 67.160 134.095 67.480 134.155 ;
        RECT 71.775 134.095 72.065 134.140 ;
        RECT 74.075 134.095 74.365 134.140 ;
        RECT 67.160 133.955 74.365 134.095 ;
        RECT 67.160 133.895 67.480 133.955 ;
        RECT 71.775 133.910 72.065 133.955 ;
        RECT 74.075 133.910 74.365 133.955 ;
        RECT 74.520 133.895 74.840 134.155 ;
        RECT 74.980 133.895 75.300 134.155 ;
        RECT 80.040 134.140 80.360 134.155 ;
        RECT 77.295 134.095 77.585 134.140 ;
        RECT 79.825 134.095 80.360 134.140 ;
        RECT 77.295 133.955 80.360 134.095 ;
        RECT 77.295 133.910 77.585 133.955 ;
        RECT 79.825 133.910 80.360 133.955 ;
        RECT 83.690 134.095 83.980 134.140 ;
        RECT 83.690 133.955 86.225 134.095 ;
        RECT 83.690 133.910 83.980 133.955 ;
        RECT 80.040 133.895 80.360 133.910 ;
        RECT 56.135 133.755 56.425 133.800 ;
        RECT 59.290 133.755 59.580 133.800 ;
        RECT 62.550 133.755 62.840 133.800 ;
        RECT 56.135 133.615 62.840 133.755 ;
        RECT 56.135 133.570 56.425 133.615 ;
        RECT 59.290 133.570 59.580 133.615 ;
        RECT 62.550 133.570 62.840 133.615 ;
        RECT 63.470 133.755 63.760 133.800 ;
        RECT 65.330 133.755 65.620 133.800 ;
        RECT 63.470 133.615 65.620 133.755 ;
        RECT 63.470 133.570 63.760 133.615 ;
        RECT 65.330 133.570 65.620 133.615 ;
        RECT 65.780 133.755 66.100 133.815 ;
        RECT 66.700 133.755 67.020 133.815 ;
        RECT 67.635 133.755 67.925 133.800 ;
        RECT 65.780 133.615 67.925 133.755 ;
        RECT 65.780 133.555 66.100 133.615 ;
        RECT 66.700 133.555 67.020 133.615 ;
        RECT 67.635 133.570 67.925 133.615 ;
        RECT 81.830 133.755 82.120 133.800 ;
        RECT 84.180 133.755 84.500 133.815 ;
        RECT 86.010 133.800 86.225 133.955 ;
        RECT 86.940 133.895 87.260 134.155 ;
        RECT 91.095 134.095 91.385 134.140 ;
        RECT 93.930 134.095 94.070 134.235 ;
        RECT 91.095 133.955 94.070 134.095 ;
        RECT 94.300 134.095 94.620 134.155 ;
        RECT 95.310 134.095 95.450 134.295 ;
        RECT 105.355 134.250 105.645 134.295 ;
        RECT 107.640 134.235 107.960 134.295 ;
        RECT 109.035 134.250 109.325 134.295 ;
        RECT 98.040 134.095 98.330 134.140 ;
        RECT 94.300 133.955 95.450 134.095 ;
        RECT 95.795 133.955 98.330 134.095 ;
        RECT 91.095 133.910 91.385 133.955 ;
        RECT 94.300 133.895 94.620 133.955 ;
        RECT 95.795 133.800 96.010 133.955 ;
        RECT 98.040 133.910 98.330 133.955 ;
        RECT 99.360 134.095 99.680 134.155 ;
        RECT 101.905 134.095 102.195 134.140 ;
        RECT 105.815 134.095 106.105 134.140 ;
        RECT 99.360 133.955 106.105 134.095 ;
        RECT 99.360 133.895 99.680 133.955 ;
        RECT 101.905 133.910 102.195 133.955 ;
        RECT 105.815 133.910 106.105 133.955 ;
        RECT 106.260 134.095 106.580 134.155 ;
        RECT 109.955 134.095 110.245 134.140 ;
        RECT 106.260 133.955 110.245 134.095 ;
        RECT 106.260 133.895 106.580 133.955 ;
        RECT 109.955 133.910 110.245 133.955 ;
        RECT 85.090 133.755 85.380 133.800 ;
        RECT 81.830 133.615 85.380 133.755 ;
        RECT 81.830 133.570 82.120 133.615 ;
        RECT 84.180 133.555 84.500 133.615 ;
        RECT 85.090 133.570 85.380 133.615 ;
        RECT 86.010 133.755 86.300 133.800 ;
        RECT 87.870 133.755 88.160 133.800 ;
        RECT 86.010 133.615 88.160 133.755 ;
        RECT 86.010 133.570 86.300 133.615 ;
        RECT 87.870 133.570 88.160 133.615 ;
        RECT 93.860 133.755 94.150 133.800 ;
        RECT 95.720 133.755 96.010 133.800 ;
        RECT 96.640 133.755 96.930 133.800 ;
        RECT 99.900 133.755 100.190 133.800 ;
        RECT 93.860 133.615 96.010 133.755 ;
        RECT 93.860 133.570 94.150 133.615 ;
        RECT 95.720 133.570 96.010 133.615 ;
        RECT 96.230 133.615 100.190 133.755 ;
        RECT 67.160 133.415 67.480 133.475 ;
        RECT 48.390 133.275 67.480 133.415 ;
        RECT 36.355 133.230 36.645 133.275 ;
        RECT 39.100 133.215 39.420 133.275 ;
        RECT 67.160 133.215 67.480 133.275 ;
        RECT 68.095 133.415 68.385 133.460 ;
        RECT 68.540 133.415 68.860 133.475 ;
        RECT 68.095 133.275 68.860 133.415 ;
        RECT 68.095 133.230 68.385 133.275 ;
        RECT 68.540 133.215 68.860 133.275 ;
        RECT 75.440 133.415 75.760 133.475 ;
        RECT 76.835 133.415 77.125 133.460 ;
        RECT 75.440 133.275 77.125 133.415 ;
        RECT 75.440 133.215 75.760 133.275 ;
        RECT 76.835 133.230 77.125 133.275 ;
        RECT 79.135 133.415 79.425 133.460 ;
        RECT 82.340 133.415 82.660 133.475 ;
        RECT 79.135 133.275 82.660 133.415 ;
        RECT 79.135 133.230 79.425 133.275 ;
        RECT 82.340 133.215 82.660 133.275 ;
        RECT 91.555 133.415 91.845 133.460 ;
        RECT 96.230 133.415 96.370 133.615 ;
        RECT 96.640 133.570 96.930 133.615 ;
        RECT 99.900 133.570 100.190 133.615 ;
        RECT 91.555 133.275 96.370 133.415 ;
        RECT 91.555 133.230 91.845 133.275 ;
        RECT 110.400 133.215 110.720 133.475 ;
        RECT 112.255 133.415 112.545 133.460 ;
        RECT 112.700 133.415 113.020 133.475 ;
        RECT 112.255 133.275 113.020 133.415 ;
        RECT 135.590 133.400 136.850 134.480 ;
        RECT 112.255 133.230 112.545 133.275 ;
        RECT 112.700 133.215 113.020 133.275 ;
        RECT 10.650 132.595 118.610 133.075 ;
        RECT 18.400 132.195 18.720 132.455 ;
        RECT 20.255 132.395 20.545 132.440 ;
        RECT 21.160 132.395 21.480 132.455 ;
        RECT 20.255 132.255 21.480 132.395 ;
        RECT 20.255 132.210 20.545 132.255 ;
        RECT 15.655 132.055 15.945 132.100 ;
        RECT 20.330 132.055 20.470 132.210 ;
        RECT 21.160 132.195 21.480 132.255 ;
        RECT 28.765 132.395 29.055 132.440 ;
        RECT 31.740 132.395 32.060 132.455 ;
        RECT 28.765 132.255 32.060 132.395 ;
        RECT 28.765 132.210 29.055 132.255 ;
        RECT 31.740 132.195 32.060 132.255 ;
        RECT 38.195 132.210 38.485 132.440 ;
        RECT 46.920 132.395 47.240 132.455 ;
        RECT 48.315 132.395 48.605 132.440 ;
        RECT 59.800 132.395 60.120 132.455 ;
        RECT 61.195 132.395 61.485 132.440 ;
        RECT 68.540 132.395 68.860 132.455 ;
        RECT 85.115 132.395 85.405 132.440 ;
        RECT 86.940 132.395 87.260 132.455 ;
        RECT 46.920 132.255 48.605 132.395 ;
        RECT 15.655 131.915 20.470 132.055 ;
        RECT 27.155 132.055 27.445 132.100 ;
        RECT 30.770 132.055 31.060 132.100 ;
        RECT 34.030 132.055 34.320 132.100 ;
        RECT 27.155 131.915 34.320 132.055 ;
        RECT 15.655 131.870 15.945 131.915 ;
        RECT 27.155 131.870 27.445 131.915 ;
        RECT 30.770 131.870 31.060 131.915 ;
        RECT 34.030 131.870 34.320 131.915 ;
        RECT 34.950 132.055 35.240 132.100 ;
        RECT 36.810 132.055 37.100 132.100 ;
        RECT 34.950 131.915 37.100 132.055 ;
        RECT 34.950 131.870 35.240 131.915 ;
        RECT 36.810 131.870 37.100 131.915 ;
        RECT 16.100 131.515 16.420 131.775 ;
        RECT 26.220 131.715 26.540 131.775 ;
        RECT 26.695 131.715 26.985 131.760 ;
        RECT 18.490 131.575 21.850 131.715 ;
        RECT 15.195 131.375 15.485 131.420 ;
        RECT 18.490 131.375 18.630 131.575 ;
        RECT 15.195 131.235 18.630 131.375 ;
        RECT 18.860 131.375 19.180 131.435 ;
        RECT 21.710 131.420 21.850 131.575 ;
        RECT 26.220 131.575 26.985 131.715 ;
        RECT 26.220 131.515 26.540 131.575 ;
        RECT 26.695 131.530 26.985 131.575 ;
        RECT 32.630 131.715 32.920 131.760 ;
        RECT 34.950 131.715 35.165 131.870 ;
        RECT 32.630 131.575 35.165 131.715 ;
        RECT 35.895 131.715 36.185 131.760 ;
        RECT 38.270 131.715 38.410 132.210 ;
        RECT 46.920 132.195 47.240 132.255 ;
        RECT 48.315 132.210 48.605 132.255 ;
        RECT 49.310 132.255 59.340 132.395 ;
        RECT 44.620 132.055 44.940 132.115 ;
        RECT 49.310 132.055 49.450 132.255 ;
        RECT 44.620 131.915 49.450 132.055 ;
        RECT 59.200 132.055 59.340 132.255 ;
        RECT 59.800 132.255 61.485 132.395 ;
        RECT 59.800 132.195 60.120 132.255 ;
        RECT 61.195 132.210 61.485 132.255 ;
        RECT 67.710 132.255 84.870 132.395 ;
        RECT 67.710 132.055 67.850 132.255 ;
        RECT 68.540 132.195 68.860 132.255 ;
        RECT 69.015 132.055 69.305 132.100 ;
        RECT 59.200 131.915 67.850 132.055 ;
        RECT 68.630 131.915 69.305 132.055 ;
        RECT 44.620 131.855 44.940 131.915 ;
        RECT 35.895 131.575 38.410 131.715 ;
        RECT 32.630 131.530 32.920 131.575 ;
        RECT 35.895 131.530 36.185 131.575 ;
        RECT 39.100 131.515 39.420 131.775 ;
        RECT 49.310 131.760 49.450 131.915 ;
        RECT 49.235 131.530 49.525 131.760 ;
        RECT 58.435 131.715 58.725 131.760 ;
        RECT 64.415 131.715 64.705 131.760 ;
        RECT 58.435 131.575 62.790 131.715 ;
        RECT 58.435 131.530 58.725 131.575 ;
        RECT 20.715 131.375 21.005 131.420 ;
        RECT 18.860 131.235 21.005 131.375 ;
        RECT 15.195 131.190 15.485 131.235 ;
        RECT 18.860 131.175 19.180 131.235 ;
        RECT 20.715 131.190 21.005 131.235 ;
        RECT 21.635 131.375 21.925 131.420 ;
        RECT 25.760 131.375 26.080 131.435 ;
        RECT 21.635 131.235 26.080 131.375 ;
        RECT 21.635 131.190 21.925 131.235 ;
        RECT 20.790 131.035 20.930 131.190 ;
        RECT 25.760 131.175 26.080 131.235 ;
        RECT 27.140 131.375 27.460 131.435 ;
        RECT 37.735 131.375 38.025 131.420 ;
        RECT 27.140 131.235 38.025 131.375 ;
        RECT 27.140 131.175 27.460 131.235 ;
        RECT 37.735 131.190 38.025 131.235 ;
        RECT 50.140 131.175 50.460 131.435 ;
        RECT 60.260 131.175 60.580 131.435 ;
        RECT 60.735 131.190 61.025 131.420 ;
        RECT 30.360 131.035 30.680 131.095 ;
        RECT 20.790 130.895 30.680 131.035 ;
        RECT 30.360 130.835 30.680 130.895 ;
        RECT 32.630 131.035 32.920 131.080 ;
        RECT 35.410 131.035 35.700 131.080 ;
        RECT 37.270 131.035 37.560 131.080 ;
        RECT 32.630 130.895 37.560 131.035 ;
        RECT 32.630 130.850 32.920 130.895 ;
        RECT 35.410 130.850 35.700 130.895 ;
        RECT 37.270 130.850 37.560 130.895 ;
        RECT 55.660 131.035 55.980 131.095 ;
        RECT 60.810 131.035 60.950 131.190 ;
        RECT 55.660 130.895 60.950 131.035 ;
        RECT 55.660 130.835 55.980 130.895 ;
        RECT 17.940 130.495 18.260 130.755 ;
        RECT 57.040 130.495 57.360 130.755 ;
        RECT 62.650 130.695 62.790 131.575 ;
        RECT 63.110 131.575 64.705 131.715 ;
        RECT 63.110 131.080 63.250 131.575 ;
        RECT 64.415 131.530 64.705 131.575 ;
        RECT 66.700 131.515 67.020 131.775 ;
        RECT 65.795 131.375 66.085 131.420 ;
        RECT 68.080 131.375 68.400 131.435 ;
        RECT 65.795 131.235 68.400 131.375 ;
        RECT 65.795 131.190 66.085 131.235 ;
        RECT 68.080 131.175 68.400 131.235 ;
        RECT 63.035 130.850 63.325 131.080 ;
        RECT 67.635 131.035 67.925 131.080 ;
        RECT 68.630 131.035 68.770 131.915 ;
        RECT 69.015 131.870 69.305 131.915 ;
        RECT 75.440 131.515 75.760 131.775 ;
        RECT 80.975 131.715 81.265 131.760 ;
        RECT 77.370 131.575 81.265 131.715 ;
        RECT 70.395 131.375 70.685 131.420 ;
        RECT 74.535 131.375 74.825 131.420 ;
        RECT 70.395 131.235 74.825 131.375 ;
        RECT 70.395 131.190 70.685 131.235 ;
        RECT 74.535 131.190 74.825 131.235 ;
        RECT 74.980 131.375 75.300 131.435 ;
        RECT 76.820 131.375 77.140 131.435 ;
        RECT 74.980 131.235 77.140 131.375 ;
        RECT 64.950 130.895 68.770 131.035 ;
        RECT 74.610 131.035 74.750 131.190 ;
        RECT 74.980 131.175 75.300 131.235 ;
        RECT 76.820 131.175 77.140 131.235 ;
        RECT 76.360 131.035 76.680 131.095 ;
        RECT 77.370 131.080 77.510 131.575 ;
        RECT 80.975 131.530 81.265 131.575 ;
        RECT 82.340 131.715 82.660 131.775 ;
        RECT 84.195 131.715 84.485 131.760 ;
        RECT 82.340 131.575 84.485 131.715 ;
        RECT 84.730 131.715 84.870 132.255 ;
        RECT 85.115 132.255 87.260 132.395 ;
        RECT 85.115 132.210 85.405 132.255 ;
        RECT 86.940 132.195 87.260 132.255 ;
        RECT 90.620 132.395 90.940 132.455 ;
        RECT 91.095 132.395 91.385 132.440 ;
        RECT 90.620 132.255 91.385 132.395 ;
        RECT 90.620 132.195 90.940 132.255 ;
        RECT 91.095 132.210 91.385 132.255 ;
        RECT 97.995 132.395 98.285 132.440 ;
        RECT 98.440 132.395 98.760 132.455 ;
        RECT 97.995 132.255 98.760 132.395 ;
        RECT 97.995 132.210 98.285 132.255 ;
        RECT 98.440 132.195 98.760 132.255 ;
        RECT 100.280 132.195 100.600 132.455 ;
        RECT 102.595 132.395 102.885 132.440 ;
        RECT 103.040 132.395 103.360 132.455 ;
        RECT 102.595 132.255 103.360 132.395 ;
        RECT 102.595 132.210 102.885 132.255 ;
        RECT 103.040 132.195 103.360 132.255 ;
        RECT 112.240 132.100 112.560 132.115 ;
        RECT 108.970 132.055 109.260 132.100 ;
        RECT 112.230 132.055 112.560 132.100 ;
        RECT 92.090 131.915 99.130 132.055 ;
        RECT 92.090 131.760 92.230 131.915 ;
        RECT 98.990 131.760 99.130 131.915 ;
        RECT 108.970 131.915 112.560 132.055 ;
        RECT 108.970 131.870 109.260 131.915 ;
        RECT 112.230 131.870 112.560 131.915 ;
        RECT 112.240 131.855 112.560 131.870 ;
        RECT 113.150 132.055 113.440 132.100 ;
        RECT 115.010 132.055 115.300 132.100 ;
        RECT 113.150 131.915 115.300 132.055 ;
        RECT 113.150 131.870 113.440 131.915 ;
        RECT 115.010 131.870 115.300 131.915 ;
        RECT 92.015 131.715 92.305 131.760 ;
        RECT 95.235 131.715 95.525 131.760 ;
        RECT 84.730 131.575 92.305 131.715 ;
        RECT 82.340 131.515 82.660 131.575 ;
        RECT 84.195 131.530 84.485 131.575 ;
        RECT 92.015 131.530 92.305 131.575 ;
        RECT 93.010 131.575 95.525 131.715 ;
        RECT 88.320 131.375 88.640 131.435 ;
        RECT 93.010 131.420 93.150 131.575 ;
        RECT 95.235 131.530 95.525 131.575 ;
        RECT 98.915 131.715 99.205 131.760 ;
        RECT 101.215 131.715 101.505 131.760 ;
        RECT 102.580 131.715 102.900 131.775 ;
        RECT 103.515 131.715 103.805 131.760 ;
        RECT 98.915 131.575 103.805 131.715 ;
        RECT 98.915 131.530 99.205 131.575 ;
        RECT 101.215 131.530 101.505 131.575 ;
        RECT 102.580 131.515 102.900 131.575 ;
        RECT 103.515 131.530 103.805 131.575 ;
        RECT 110.830 131.715 111.120 131.760 ;
        RECT 113.150 131.715 113.365 131.870 ;
        RECT 110.830 131.575 113.365 131.715 ;
        RECT 115.460 131.715 115.780 131.775 ;
        RECT 115.935 131.715 116.225 131.760 ;
        RECT 115.460 131.575 116.225 131.715 ;
        RECT 110.830 131.530 111.120 131.575 ;
        RECT 115.460 131.515 115.780 131.575 ;
        RECT 115.935 131.530 116.225 131.575 ;
        RECT 92.935 131.375 93.225 131.420 ;
        RECT 88.320 131.235 93.225 131.375 ;
        RECT 88.320 131.175 88.640 131.235 ;
        RECT 92.935 131.190 93.225 131.235 ;
        RECT 94.300 131.175 94.620 131.435 ;
        RECT 94.775 131.375 95.065 131.420 ;
        RECT 99.835 131.375 100.125 131.420 ;
        RECT 94.775 131.235 100.125 131.375 ;
        RECT 94.775 131.190 95.065 131.235 ;
        RECT 99.835 131.190 100.125 131.235 ;
        RECT 102.135 131.375 102.425 131.420 ;
        RECT 103.040 131.375 103.360 131.435 ;
        RECT 102.135 131.235 103.360 131.375 ;
        RECT 102.135 131.190 102.425 131.235 ;
        RECT 74.610 130.895 76.680 131.035 ;
        RECT 64.950 130.695 65.090 130.895 ;
        RECT 67.635 130.850 67.925 130.895 ;
        RECT 76.360 130.835 76.680 130.895 ;
        RECT 77.295 130.850 77.585 131.080 ;
        RECT 98.900 131.035 99.220 131.095 ;
        RECT 99.910 131.035 100.050 131.190 ;
        RECT 103.040 131.175 103.360 131.235 ;
        RECT 104.435 131.375 104.725 131.420 ;
        RECT 106.965 131.375 107.255 131.420 ;
        RECT 110.400 131.375 110.720 131.435 ;
        RECT 104.435 131.235 110.720 131.375 ;
        RECT 104.435 131.190 104.725 131.235 ;
        RECT 106.965 131.190 107.255 131.235 ;
        RECT 110.400 131.175 110.720 131.235 ;
        RECT 114.080 131.175 114.400 131.435 ;
        RECT 98.900 130.895 100.050 131.035 ;
        RECT 110.830 131.035 111.120 131.080 ;
        RECT 113.610 131.035 113.900 131.080 ;
        RECT 115.470 131.035 115.760 131.080 ;
        RECT 110.830 130.895 115.760 131.035 ;
        RECT 98.900 130.835 99.220 130.895 ;
        RECT 110.830 130.850 111.120 130.895 ;
        RECT 113.610 130.850 113.900 130.895 ;
        RECT 115.470 130.850 115.760 130.895 ;
        RECT 62.650 130.555 65.090 130.695 ;
        RECT 65.320 130.495 65.640 130.755 ;
        RECT 80.040 130.495 80.360 130.755 ;
        RECT 96.140 130.695 96.460 130.755 ;
        RECT 97.075 130.695 97.365 130.740 ;
        RECT 96.140 130.555 97.365 130.695 ;
        RECT 96.140 130.495 96.460 130.555 ;
        RECT 97.075 130.510 97.365 130.555 ;
        RECT 11.430 129.875 118.610 130.355 ;
        RECT 34.960 129.675 35.280 129.735 ;
        RECT 35.895 129.675 36.185 129.720 ;
        RECT 34.960 129.535 36.185 129.675 ;
        RECT 34.960 129.475 35.280 129.535 ;
        RECT 35.895 129.490 36.185 129.535 ;
        RECT 55.660 129.675 55.980 129.735 ;
        RECT 57.285 129.675 57.575 129.720 ;
        RECT 55.660 129.535 57.575 129.675 ;
        RECT 55.660 129.475 55.980 129.535 ;
        RECT 57.285 129.490 57.575 129.535 ;
        RECT 70.625 129.675 70.915 129.720 ;
        RECT 75.440 129.675 75.760 129.735 ;
        RECT 70.625 129.535 75.760 129.675 ;
        RECT 70.625 129.490 70.915 129.535 ;
        RECT 75.440 129.475 75.760 129.535 ;
        RECT 82.355 129.675 82.645 129.720 ;
        RECT 89.240 129.675 89.560 129.735 ;
        RECT 82.355 129.535 89.560 129.675 ;
        RECT 82.355 129.490 82.645 129.535 ;
        RECT 45.970 129.335 46.260 129.380 ;
        RECT 48.750 129.335 49.040 129.380 ;
        RECT 50.610 129.335 50.900 129.380 ;
        RECT 45.970 129.195 50.900 129.335 ;
        RECT 45.970 129.150 46.260 129.195 ;
        RECT 48.750 129.150 49.040 129.195 ;
        RECT 50.610 129.150 50.900 129.195 ;
        RECT 51.520 129.335 51.840 129.395 ;
        RECT 53.375 129.335 53.665 129.380 ;
        RECT 51.520 129.195 53.665 129.335 ;
        RECT 51.520 129.135 51.840 129.195 ;
        RECT 53.375 129.150 53.665 129.195 ;
        RECT 61.150 129.335 61.440 129.380 ;
        RECT 63.930 129.335 64.220 129.380 ;
        RECT 65.790 129.335 66.080 129.380 ;
        RECT 61.150 129.195 66.080 129.335 ;
        RECT 61.150 129.150 61.440 129.195 ;
        RECT 63.930 129.150 64.220 129.195 ;
        RECT 65.790 129.150 66.080 129.195 ;
        RECT 74.490 129.335 74.780 129.380 ;
        RECT 77.270 129.335 77.560 129.380 ;
        RECT 79.130 129.335 79.420 129.380 ;
        RECT 82.430 129.335 82.570 129.490 ;
        RECT 89.240 129.475 89.560 129.535 ;
        RECT 111.795 129.675 112.085 129.720 ;
        RECT 112.240 129.675 112.560 129.735 ;
        RECT 111.795 129.535 112.560 129.675 ;
        RECT 111.795 129.490 112.085 129.535 ;
        RECT 112.240 129.475 112.560 129.535 ;
        RECT 113.635 129.675 113.925 129.720 ;
        RECT 114.080 129.675 114.400 129.735 ;
        RECT 113.635 129.535 114.400 129.675 ;
        RECT 113.635 129.490 113.925 129.535 ;
        RECT 114.080 129.475 114.400 129.535 ;
        RECT 107.640 129.335 107.960 129.395 ;
        RECT 74.490 129.195 79.420 129.335 ;
        RECT 74.490 129.150 74.780 129.195 ;
        RECT 77.270 129.150 77.560 129.195 ;
        RECT 79.130 129.150 79.420 129.195 ;
        RECT 79.670 129.195 82.570 129.335 ;
        RECT 106.810 129.195 107.960 129.335 ;
        RECT 16.100 128.995 16.420 129.055 ;
        RECT 21.175 128.995 21.465 129.040 ;
        RECT 25.760 128.995 26.080 129.055 ;
        RECT 31.280 128.995 31.600 129.055 ;
        RECT 37.735 128.995 38.025 129.040 ;
        RECT 45.540 128.995 45.860 129.055 ;
        RECT 16.100 128.855 20.470 128.995 ;
        RECT 16.100 128.795 16.420 128.855 ;
        RECT 14.720 128.455 15.040 128.715 ;
        RECT 16.575 128.655 16.865 128.700 ;
        RECT 17.940 128.655 18.260 128.715 ;
        RECT 20.330 128.700 20.470 128.855 ;
        RECT 21.175 128.855 45.860 128.995 ;
        RECT 21.175 128.810 21.465 128.855 ;
        RECT 25.760 128.795 26.080 128.855 ;
        RECT 31.280 128.795 31.600 128.855 ;
        RECT 37.735 128.810 38.025 128.855 ;
        RECT 45.540 128.795 45.860 128.855 ;
        RECT 51.075 128.995 51.365 129.040 ;
        RECT 53.820 128.995 54.140 129.055 ;
        RECT 64.415 128.995 64.705 129.040 ;
        RECT 65.320 128.995 65.640 129.055 ;
        RECT 79.670 129.040 79.810 129.195 ;
        RECT 51.075 128.855 64.170 128.995 ;
        RECT 51.075 128.810 51.365 128.855 ;
        RECT 53.820 128.795 54.140 128.855 ;
        RECT 16.575 128.515 18.260 128.655 ;
        RECT 16.575 128.470 16.865 128.515 ;
        RECT 17.940 128.455 18.260 128.515 ;
        RECT 20.255 128.655 20.545 128.700 ;
        RECT 26.680 128.655 27.000 128.715 ;
        RECT 20.255 128.515 27.000 128.655 ;
        RECT 20.255 128.470 20.545 128.515 ;
        RECT 26.680 128.455 27.000 128.515 ;
        RECT 29.900 128.655 30.220 128.715 ;
        RECT 34.055 128.655 34.345 128.700 ;
        RECT 29.900 128.515 34.345 128.655 ;
        RECT 29.900 128.455 30.220 128.515 ;
        RECT 34.055 128.470 34.345 128.515 ;
        RECT 34.975 128.655 35.265 128.700 ;
        RECT 36.340 128.655 36.660 128.715 ;
        RECT 34.975 128.515 36.660 128.655 ;
        RECT 34.975 128.470 35.265 128.515 ;
        RECT 36.340 128.455 36.660 128.515 ;
        RECT 40.480 128.455 40.800 128.715 ;
        RECT 45.970 128.655 46.260 128.700 ;
        RECT 45.970 128.515 48.505 128.655 ;
        RECT 45.970 128.470 46.260 128.515 ;
        RECT 38.195 128.315 38.485 128.360 ;
        RECT 39.100 128.315 39.420 128.375 ;
        RECT 40.570 128.315 40.710 128.455 ;
        RECT 42.105 128.315 42.395 128.360 ;
        RECT 38.195 128.175 42.395 128.315 ;
        RECT 38.195 128.130 38.485 128.175 ;
        RECT 39.100 128.115 39.420 128.175 ;
        RECT 42.105 128.130 42.395 128.175 ;
        RECT 43.240 128.315 43.560 128.375 ;
        RECT 48.290 128.360 48.505 128.515 ;
        RECT 49.220 128.455 49.540 128.715 ;
        RECT 52.455 128.655 52.745 128.700 ;
        RECT 53.360 128.655 53.680 128.715 ;
        RECT 52.455 128.515 53.680 128.655 ;
        RECT 52.455 128.470 52.745 128.515 ;
        RECT 53.360 128.455 53.680 128.515 ;
        RECT 54.280 128.455 54.600 128.715 ;
        RECT 56.210 128.700 56.350 128.855 ;
        RECT 56.135 128.470 56.425 128.700 ;
        RECT 61.150 128.655 61.440 128.700 ;
        RECT 64.030 128.655 64.170 128.855 ;
        RECT 64.415 128.855 65.640 128.995 ;
        RECT 64.415 128.810 64.705 128.855 ;
        RECT 65.320 128.795 65.640 128.855 ;
        RECT 79.595 128.810 79.885 129.040 ;
        RECT 81.880 128.995 82.200 129.055 ;
        RECT 106.810 129.040 106.950 129.195 ;
        RECT 107.640 129.135 107.960 129.195 ;
        RECT 109.495 129.335 109.785 129.380 ;
        RECT 110.860 129.335 111.180 129.395 ;
        RECT 109.495 129.195 111.180 129.335 ;
        RECT 109.495 129.150 109.785 129.195 ;
        RECT 110.860 129.135 111.180 129.195 ;
        RECT 81.880 128.855 89.470 128.995 ;
        RECT 81.880 128.795 82.200 128.855 ;
        RECT 66.240 128.655 66.560 128.715 ;
        RECT 61.150 128.515 63.685 128.655 ;
        RECT 64.030 128.515 66.560 128.655 ;
        RECT 61.150 128.470 61.440 128.515 ;
        RECT 62.560 128.360 62.880 128.375 ;
        RECT 44.110 128.315 44.400 128.360 ;
        RECT 47.370 128.315 47.660 128.360 ;
        RECT 43.240 128.175 47.660 128.315 ;
        RECT 43.240 128.115 43.560 128.175 ;
        RECT 44.110 128.130 44.400 128.175 ;
        RECT 47.370 128.130 47.660 128.175 ;
        RECT 48.290 128.315 48.580 128.360 ;
        RECT 50.150 128.315 50.440 128.360 ;
        RECT 48.290 128.175 50.440 128.315 ;
        RECT 48.290 128.130 48.580 128.175 ;
        RECT 50.150 128.130 50.440 128.175 ;
        RECT 59.290 128.315 59.580 128.360 ;
        RECT 62.550 128.315 62.880 128.360 ;
        RECT 59.290 128.175 62.880 128.315 ;
        RECT 59.290 128.130 59.580 128.175 ;
        RECT 62.550 128.130 62.880 128.175 ;
        RECT 63.470 128.360 63.685 128.515 ;
        RECT 66.240 128.455 66.560 128.515 ;
        RECT 74.490 128.655 74.780 128.700 ;
        RECT 77.755 128.655 78.045 128.700 ;
        RECT 80.040 128.655 80.360 128.715 ;
        RECT 74.490 128.515 77.025 128.655 ;
        RECT 74.490 128.470 74.780 128.515 ;
        RECT 63.470 128.315 63.760 128.360 ;
        RECT 65.330 128.315 65.620 128.360 ;
        RECT 63.470 128.175 65.620 128.315 ;
        RECT 63.470 128.130 63.760 128.175 ;
        RECT 65.330 128.130 65.620 128.175 ;
        RECT 72.630 128.315 72.920 128.360 ;
        RECT 74.060 128.315 74.380 128.375 ;
        RECT 76.810 128.360 77.025 128.515 ;
        RECT 77.755 128.515 80.360 128.655 ;
        RECT 77.755 128.470 78.045 128.515 ;
        RECT 80.040 128.455 80.360 128.515 ;
        RECT 88.780 128.455 89.100 128.715 ;
        RECT 89.330 128.700 89.470 128.855 ;
        RECT 106.735 128.810 107.025 129.040 ;
        RECT 107.195 128.995 107.485 129.040 ;
        RECT 110.400 128.995 110.720 129.055 ;
        RECT 107.195 128.855 110.720 128.995 ;
        RECT 107.195 128.810 107.485 128.855 ;
        RECT 110.400 128.795 110.720 128.855 ;
        RECT 89.255 128.470 89.545 128.700 ;
        RECT 95.220 128.455 95.540 128.715 ;
        RECT 103.040 128.655 103.360 128.715 ;
        RECT 107.655 128.655 107.945 128.700 ;
        RECT 103.040 128.515 107.945 128.655 ;
        RECT 103.040 128.455 103.360 128.515 ;
        RECT 107.655 128.470 107.945 128.515 ;
        RECT 109.020 128.655 109.340 128.715 ;
        RECT 112.255 128.655 112.545 128.700 ;
        RECT 109.020 128.515 112.545 128.655 ;
        RECT 109.020 128.455 109.340 128.515 ;
        RECT 112.255 128.470 112.545 128.515 ;
        RECT 112.700 128.455 113.020 128.715 ;
        RECT 75.890 128.315 76.180 128.360 ;
        RECT 72.630 128.175 76.180 128.315 ;
        RECT 72.630 128.130 72.920 128.175 ;
        RECT 62.560 128.115 62.880 128.130 ;
        RECT 74.060 128.115 74.380 128.175 ;
        RECT 75.890 128.130 76.180 128.175 ;
        RECT 76.810 128.315 77.100 128.360 ;
        RECT 78.670 128.315 78.960 128.360 ;
        RECT 76.810 128.175 78.960 128.315 ;
        RECT 88.870 128.315 89.010 128.455 ;
        RECT 96.615 128.315 96.905 128.360 ;
        RECT 88.870 128.175 96.905 128.315 ;
        RECT 76.810 128.130 77.100 128.175 ;
        RECT 78.670 128.130 78.960 128.175 ;
        RECT 96.615 128.130 96.905 128.175 ;
        RECT 105.355 128.315 105.645 128.360 ;
        RECT 106.720 128.315 107.040 128.375 ;
        RECT 105.355 128.175 107.640 128.315 ;
        RECT 105.355 128.130 105.645 128.175 ;
        RECT 106.720 128.115 107.040 128.175 ;
        RECT 14.275 127.975 14.565 128.020 ;
        RECT 16.100 127.975 16.420 128.035 ;
        RECT 14.275 127.835 16.420 127.975 ;
        RECT 14.275 127.790 14.565 127.835 ;
        RECT 16.100 127.775 16.420 127.835 ;
        RECT 17.480 127.775 17.800 128.035 ;
        RECT 17.940 127.775 18.260 128.035 ;
        RECT 19.320 127.975 19.640 128.035 ;
        RECT 19.795 127.975 20.085 128.020 ;
        RECT 19.320 127.835 20.085 127.975 ;
        RECT 19.320 127.775 19.640 127.835 ;
        RECT 19.795 127.790 20.085 127.835 ;
        RECT 36.800 127.975 37.120 128.035 ;
        RECT 38.655 127.975 38.945 128.020 ;
        RECT 36.800 127.835 38.945 127.975 ;
        RECT 36.800 127.775 37.120 127.835 ;
        RECT 38.655 127.790 38.945 127.835 ;
        RECT 40.495 127.975 40.785 128.020 ;
        RECT 40.940 127.975 41.260 128.035 ;
        RECT 40.495 127.835 41.260 127.975 ;
        RECT 40.495 127.790 40.785 127.835 ;
        RECT 40.940 127.775 41.260 127.835 ;
        RECT 49.680 127.975 50.000 128.035 ;
        RECT 51.995 127.975 52.285 128.020 ;
        RECT 49.680 127.835 52.285 127.975 ;
        RECT 49.680 127.775 50.000 127.835 ;
        RECT 51.995 127.790 52.285 127.835 ;
        RECT 89.700 127.775 90.020 128.035 ;
        RECT 96.155 127.975 96.445 128.020 ;
        RECT 100.280 127.975 100.600 128.035 ;
        RECT 96.155 127.835 100.600 127.975 ;
        RECT 107.500 127.975 107.640 128.175 ;
        RECT 110.875 127.975 111.165 128.020 ;
        RECT 115.460 127.975 115.780 128.035 ;
        RECT 107.500 127.835 115.780 127.975 ;
        RECT 96.155 127.790 96.445 127.835 ;
        RECT 100.280 127.775 100.600 127.835 ;
        RECT 110.875 127.790 111.165 127.835 ;
        RECT 115.460 127.775 115.780 127.835 ;
        RECT 10.650 127.155 118.610 127.635 ;
        RECT 19.780 126.955 20.100 127.015 ;
        RECT 29.900 126.955 30.220 127.015 ;
        RECT 19.780 126.815 30.220 126.955 ;
        RECT 19.780 126.755 20.100 126.815 ;
        RECT 29.900 126.755 30.220 126.815 ;
        RECT 34.285 126.955 34.575 127.000 ;
        RECT 36.800 126.955 37.120 127.015 ;
        RECT 34.285 126.815 37.120 126.955 ;
        RECT 34.285 126.770 34.575 126.815 ;
        RECT 36.800 126.755 37.120 126.815 ;
        RECT 50.140 126.955 50.460 127.015 ;
        RECT 56.135 126.955 56.425 127.000 ;
        RECT 50.140 126.815 56.425 126.955 ;
        RECT 50.140 126.755 50.460 126.815 ;
        RECT 56.135 126.770 56.425 126.815 ;
        RECT 62.560 126.955 62.880 127.015 ;
        RECT 63.495 126.955 63.785 127.000 ;
        RECT 62.560 126.815 63.785 126.955 ;
        RECT 62.560 126.755 62.880 126.815 ;
        RECT 63.495 126.770 63.785 126.815 ;
        RECT 74.060 126.755 74.380 127.015 ;
        RECT 74.520 126.955 74.840 127.015 ;
        RECT 76.835 126.955 77.125 127.000 ;
        RECT 79.580 126.955 79.900 127.015 ;
        RECT 85.115 126.955 85.405 127.000 ;
        RECT 94.300 126.955 94.620 127.015 ;
        RECT 74.520 126.815 85.405 126.955 ;
        RECT 74.520 126.755 74.840 126.815 ;
        RECT 76.835 126.770 77.125 126.815 ;
        RECT 79.580 126.755 79.900 126.815 ;
        RECT 85.115 126.770 85.405 126.815 ;
        RECT 88.870 126.815 94.620 126.955 ;
        RECT 16.100 126.660 16.420 126.675 ;
        RECT 16.050 126.615 16.420 126.660 ;
        RECT 19.310 126.615 19.600 126.660 ;
        RECT 16.050 126.475 19.600 126.615 ;
        RECT 16.050 126.430 16.420 126.475 ;
        RECT 19.310 126.430 19.600 126.475 ;
        RECT 20.230 126.615 20.520 126.660 ;
        RECT 22.090 126.615 22.380 126.660 ;
        RECT 27.140 126.615 27.460 126.675 ;
        RECT 20.230 126.475 22.380 126.615 ;
        RECT 20.230 126.430 20.520 126.475 ;
        RECT 22.090 126.430 22.380 126.475 ;
        RECT 23.090 126.475 27.460 126.615 ;
        RECT 16.100 126.415 16.420 126.430 ;
        RECT 17.910 126.275 18.200 126.320 ;
        RECT 20.230 126.275 20.445 126.430 ;
        RECT 23.090 126.320 23.230 126.475 ;
        RECT 27.140 126.415 27.460 126.475 ;
        RECT 36.290 126.615 36.580 126.660 ;
        RECT 37.720 126.615 38.040 126.675 ;
        RECT 49.680 126.660 50.000 126.675 ;
        RECT 39.550 126.615 39.840 126.660 ;
        RECT 36.290 126.475 39.840 126.615 ;
        RECT 36.290 126.430 36.580 126.475 ;
        RECT 37.720 126.415 38.040 126.475 ;
        RECT 39.550 126.430 39.840 126.475 ;
        RECT 40.470 126.615 40.760 126.660 ;
        RECT 42.330 126.615 42.620 126.660 ;
        RECT 40.470 126.475 42.620 126.615 ;
        RECT 40.470 126.430 40.760 126.475 ;
        RECT 42.330 126.430 42.620 126.475 ;
        RECT 46.410 126.615 46.700 126.660 ;
        RECT 49.670 126.615 50.000 126.660 ;
        RECT 46.410 126.475 50.000 126.615 ;
        RECT 46.410 126.430 46.700 126.475 ;
        RECT 49.670 126.430 50.000 126.475 ;
        RECT 17.910 126.135 20.445 126.275 ;
        RECT 17.910 126.090 18.200 126.135 ;
        RECT 23.015 126.090 23.305 126.320 ;
        RECT 23.935 126.275 24.225 126.320 ;
        RECT 26.220 126.275 26.540 126.335 ;
        RECT 23.935 126.135 26.540 126.275 ;
        RECT 23.935 126.090 24.225 126.135 ;
        RECT 14.045 125.935 14.335 125.980 ;
        RECT 15.640 125.935 15.960 125.995 ;
        RECT 14.045 125.795 15.960 125.935 ;
        RECT 14.045 125.750 14.335 125.795 ;
        RECT 15.640 125.735 15.960 125.795 ;
        RECT 17.480 125.935 17.800 125.995 ;
        RECT 21.175 125.935 21.465 125.980 ;
        RECT 17.480 125.795 21.465 125.935 ;
        RECT 17.480 125.735 17.800 125.795 ;
        RECT 21.175 125.750 21.465 125.795 ;
        RECT 17.910 125.595 18.200 125.640 ;
        RECT 20.690 125.595 20.980 125.640 ;
        RECT 22.550 125.595 22.840 125.640 ;
        RECT 17.910 125.455 22.840 125.595 ;
        RECT 17.910 125.410 18.200 125.455 ;
        RECT 20.690 125.410 20.980 125.455 ;
        RECT 22.550 125.410 22.840 125.455 ;
        RECT 14.720 125.255 15.040 125.315 ;
        RECT 24.010 125.255 24.150 126.090 ;
        RECT 26.220 126.075 26.540 126.135 ;
        RECT 30.360 126.075 30.680 126.335 ;
        RECT 38.150 126.275 38.440 126.320 ;
        RECT 40.470 126.275 40.685 126.430 ;
        RECT 49.680 126.415 50.000 126.430 ;
        RECT 50.590 126.615 50.880 126.660 ;
        RECT 52.450 126.615 52.740 126.660 ;
        RECT 84.655 126.615 84.945 126.660 ;
        RECT 87.645 126.615 87.935 126.660 ;
        RECT 88.320 126.615 88.640 126.675 ;
        RECT 50.590 126.475 52.740 126.615 ;
        RECT 50.590 126.430 50.880 126.475 ;
        RECT 52.450 126.430 52.740 126.475 ;
        RECT 73.690 126.475 77.970 126.615 ;
        RECT 38.150 126.135 40.685 126.275 ;
        RECT 38.150 126.090 38.440 126.135 ;
        RECT 41.400 126.075 41.720 126.335 ;
        RECT 44.160 126.320 44.480 126.335 ;
        RECT 44.160 126.090 44.695 126.320 ;
        RECT 48.270 126.275 48.560 126.320 ;
        RECT 50.590 126.275 50.805 126.430 ;
        RECT 48.270 126.135 50.805 126.275 ;
        RECT 48.270 126.090 48.560 126.135 ;
        RECT 44.160 126.075 44.480 126.090 ;
        RECT 51.520 126.075 51.840 126.335 ;
        RECT 56.595 126.275 56.885 126.320 ;
        RECT 52.070 126.135 56.885 126.275 ;
        RECT 29.455 125.750 29.745 125.980 ;
        RECT 40.480 125.935 40.800 125.995 ;
        RECT 43.255 125.935 43.545 125.980 ;
        RECT 40.480 125.795 43.545 125.935 ;
        RECT 29.530 125.595 29.670 125.750 ;
        RECT 40.480 125.735 40.800 125.795 ;
        RECT 43.255 125.750 43.545 125.795 ;
        RECT 47.380 125.935 47.700 125.995 ;
        RECT 52.070 125.935 52.210 126.135 ;
        RECT 56.595 126.090 56.885 126.135 ;
        RECT 60.720 126.275 61.040 126.335 ;
        RECT 63.955 126.275 64.245 126.320 ;
        RECT 60.720 126.135 64.245 126.275 ;
        RECT 60.720 126.075 61.040 126.135 ;
        RECT 63.955 126.090 64.245 126.135 ;
        RECT 69.460 126.275 69.780 126.335 ;
        RECT 73.690 126.320 73.830 126.475 ;
        RECT 72.235 126.275 72.525 126.320 ;
        RECT 73.615 126.275 73.905 126.320 ;
        RECT 69.460 126.135 73.905 126.275 ;
        RECT 69.460 126.075 69.780 126.135 ;
        RECT 72.235 126.090 72.525 126.135 ;
        RECT 73.615 126.090 73.905 126.135 ;
        RECT 76.820 126.275 77.140 126.335 ;
        RECT 77.295 126.275 77.585 126.320 ;
        RECT 76.820 126.135 77.585 126.275 ;
        RECT 77.830 126.275 77.970 126.475 ;
        RECT 84.655 126.475 88.640 126.615 ;
        RECT 84.655 126.430 84.945 126.475 ;
        RECT 87.645 126.430 87.935 126.475 ;
        RECT 88.320 126.415 88.640 126.475 ;
        RECT 81.880 126.275 82.200 126.335 ;
        RECT 88.870 126.275 89.010 126.815 ;
        RECT 94.300 126.755 94.620 126.815 ;
        RECT 95.220 126.955 95.540 127.015 ;
        RECT 100.755 126.955 101.045 127.000 ;
        RECT 95.220 126.815 101.045 126.955 ;
        RECT 95.220 126.755 95.540 126.815 ;
        RECT 100.755 126.770 101.045 126.815 ;
        RECT 103.040 126.955 103.360 127.015 ;
        RECT 106.045 126.955 106.335 127.000 ;
        RECT 103.040 126.815 106.335 126.955 ;
        RECT 103.040 126.755 103.360 126.815 ;
        RECT 106.045 126.770 106.335 126.815 ;
        RECT 89.700 126.660 90.020 126.675 ;
        RECT 89.650 126.615 90.020 126.660 ;
        RECT 92.910 126.615 93.200 126.660 ;
        RECT 89.650 126.475 93.200 126.615 ;
        RECT 89.650 126.430 90.020 126.475 ;
        RECT 92.910 126.430 93.200 126.475 ;
        RECT 93.830 126.615 94.120 126.660 ;
        RECT 95.690 126.615 95.980 126.660 ;
        RECT 93.830 126.475 95.980 126.615 ;
        RECT 93.830 126.430 94.120 126.475 ;
        RECT 95.690 126.430 95.980 126.475 ;
        RECT 98.900 126.615 99.220 126.675 ;
        RECT 102.595 126.615 102.885 126.660 ;
        RECT 98.900 126.475 102.885 126.615 ;
        RECT 89.700 126.415 90.020 126.430 ;
        RECT 77.830 126.135 82.200 126.275 ;
        RECT 76.820 126.075 77.140 126.135 ;
        RECT 77.295 126.090 77.585 126.135 ;
        RECT 81.880 126.075 82.200 126.135 ;
        RECT 84.270 126.135 89.010 126.275 ;
        RECT 91.510 126.275 91.800 126.320 ;
        RECT 93.830 126.275 94.045 126.430 ;
        RECT 98.900 126.415 99.220 126.475 ;
        RECT 102.595 126.430 102.885 126.475 ;
        RECT 108.050 126.615 108.340 126.660 ;
        RECT 109.480 126.615 109.800 126.675 ;
        RECT 111.310 126.615 111.600 126.660 ;
        RECT 108.050 126.475 111.600 126.615 ;
        RECT 108.050 126.430 108.340 126.475 ;
        RECT 109.480 126.415 109.800 126.475 ;
        RECT 111.310 126.430 111.600 126.475 ;
        RECT 112.230 126.615 112.520 126.660 ;
        RECT 114.090 126.615 114.380 126.660 ;
        RECT 112.230 126.475 114.380 126.615 ;
        RECT 112.230 126.430 112.520 126.475 ;
        RECT 114.090 126.430 114.380 126.475 ;
        RECT 91.510 126.135 94.045 126.275 ;
        RECT 47.380 125.795 52.210 125.935 ;
        RECT 53.375 125.935 53.665 125.980 ;
        RECT 53.820 125.935 54.140 125.995 ;
        RECT 53.375 125.795 54.140 125.935 ;
        RECT 47.380 125.735 47.700 125.795 ;
        RECT 53.375 125.750 53.665 125.795 ;
        RECT 53.820 125.735 54.140 125.795 ;
        RECT 57.040 125.735 57.360 125.995 ;
        RECT 76.360 125.935 76.680 125.995 ;
        RECT 84.270 125.980 84.410 126.135 ;
        RECT 91.510 126.090 91.800 126.135 ;
        RECT 94.760 126.075 95.080 126.335 ;
        RECT 99.375 126.090 99.665 126.320 ;
        RECT 109.910 126.275 110.200 126.320 ;
        RECT 112.230 126.275 112.445 126.430 ;
        RECT 109.910 126.135 112.445 126.275 ;
        RECT 115.015 126.275 115.305 126.320 ;
        RECT 115.460 126.275 115.780 126.335 ;
        RECT 115.015 126.135 115.780 126.275 ;
        RECT 109.910 126.090 110.200 126.135 ;
        RECT 115.015 126.090 115.305 126.135 ;
        RECT 84.195 125.935 84.485 125.980 ;
        RECT 76.360 125.795 84.485 125.935 ;
        RECT 76.360 125.735 76.680 125.795 ;
        RECT 84.195 125.750 84.485 125.795 ;
        RECT 89.240 125.935 89.560 125.995 ;
        RECT 96.615 125.935 96.905 125.980 ;
        RECT 89.240 125.795 96.905 125.935 ;
        RECT 89.240 125.735 89.560 125.795 ;
        RECT 96.615 125.750 96.905 125.795 ;
        RECT 31.280 125.595 31.600 125.655 ;
        RECT 29.530 125.455 31.600 125.595 ;
        RECT 31.280 125.395 31.600 125.455 ;
        RECT 38.150 125.595 38.440 125.640 ;
        RECT 40.930 125.595 41.220 125.640 ;
        RECT 42.790 125.595 43.080 125.640 ;
        RECT 38.150 125.455 43.080 125.595 ;
        RECT 38.150 125.410 38.440 125.455 ;
        RECT 40.930 125.410 41.220 125.455 ;
        RECT 42.790 125.410 43.080 125.455 ;
        RECT 48.270 125.595 48.560 125.640 ;
        RECT 51.050 125.595 51.340 125.640 ;
        RECT 52.910 125.595 53.200 125.640 ;
        RECT 57.130 125.595 57.270 125.735 ;
        RECT 48.270 125.455 53.200 125.595 ;
        RECT 48.270 125.410 48.560 125.455 ;
        RECT 51.050 125.410 51.340 125.455 ;
        RECT 52.910 125.410 53.200 125.455 ;
        RECT 53.450 125.455 57.270 125.595 ;
        RECT 91.510 125.595 91.800 125.640 ;
        RECT 94.290 125.595 94.580 125.640 ;
        RECT 96.150 125.595 96.440 125.640 ;
        RECT 91.510 125.455 96.440 125.595 ;
        RECT 99.450 125.595 99.590 126.090 ;
        RECT 115.460 126.075 115.780 126.135 ;
        RECT 103.975 125.935 104.265 125.980 ;
        RECT 107.640 125.935 107.960 125.995 ;
        RECT 103.975 125.795 107.960 125.935 ;
        RECT 103.975 125.750 104.265 125.795 ;
        RECT 107.640 125.735 107.960 125.795 ;
        RECT 113.160 125.735 113.480 125.995 ;
        RECT 109.020 125.595 109.340 125.655 ;
        RECT 99.450 125.455 109.340 125.595 ;
        RECT 14.720 125.115 24.150 125.255 ;
        RECT 24.395 125.255 24.685 125.300 ;
        RECT 25.760 125.255 26.080 125.315 ;
        RECT 24.395 125.115 26.080 125.255 ;
        RECT 14.720 125.055 15.040 125.115 ;
        RECT 24.395 125.070 24.685 125.115 ;
        RECT 25.760 125.055 26.080 125.115 ;
        RECT 32.200 125.055 32.520 125.315 ;
        RECT 45.540 125.255 45.860 125.315 ;
        RECT 49.680 125.255 50.000 125.315 ;
        RECT 53.450 125.255 53.590 125.455 ;
        RECT 91.510 125.410 91.800 125.455 ;
        RECT 94.290 125.410 94.580 125.455 ;
        RECT 96.150 125.410 96.440 125.455 ;
        RECT 109.020 125.395 109.340 125.455 ;
        RECT 109.910 125.595 110.200 125.640 ;
        RECT 112.690 125.595 112.980 125.640 ;
        RECT 114.550 125.595 114.840 125.640 ;
        RECT 109.910 125.455 114.840 125.595 ;
        RECT 109.910 125.410 110.200 125.455 ;
        RECT 112.690 125.410 112.980 125.455 ;
        RECT 114.550 125.410 114.840 125.455 ;
        RECT 45.540 125.115 53.590 125.255 ;
        RECT 54.295 125.255 54.585 125.300 ;
        RECT 55.660 125.255 55.980 125.315 ;
        RECT 54.295 125.115 55.980 125.255 ;
        RECT 45.540 125.055 45.860 125.115 ;
        RECT 49.680 125.055 50.000 125.115 ;
        RECT 54.295 125.070 54.585 125.115 ;
        RECT 55.660 125.055 55.980 125.115 ;
        RECT 72.680 125.055 73.000 125.315 ;
        RECT 77.280 125.255 77.600 125.315 ;
        RECT 79.135 125.255 79.425 125.300 ;
        RECT 77.280 125.115 79.425 125.255 ;
        RECT 77.280 125.055 77.600 125.115 ;
        RECT 79.135 125.070 79.425 125.115 ;
        RECT 82.340 125.055 82.660 125.315 ;
        RECT 86.940 125.055 87.260 125.315 ;
        RECT 99.820 125.055 100.140 125.315 ;
        RECT 11.430 124.435 118.610 124.915 ;
        RECT 15.885 124.235 16.175 124.280 ;
        RECT 19.320 124.235 19.640 124.295 ;
        RECT 15.885 124.095 19.640 124.235 ;
        RECT 15.885 124.050 16.175 124.095 ;
        RECT 19.320 124.035 19.640 124.095 ;
        RECT 25.545 124.235 25.835 124.280 ;
        RECT 30.360 124.235 30.680 124.295 ;
        RECT 25.545 124.095 37.490 124.235 ;
        RECT 25.545 124.050 25.835 124.095 ;
        RECT 30.360 124.035 30.680 124.095 ;
        RECT 19.750 123.895 20.040 123.940 ;
        RECT 22.530 123.895 22.820 123.940 ;
        RECT 24.390 123.895 24.680 123.940 ;
        RECT 19.750 123.755 24.680 123.895 ;
        RECT 19.750 123.710 20.040 123.755 ;
        RECT 22.530 123.710 22.820 123.755 ;
        RECT 24.390 123.710 24.680 123.755 ;
        RECT 29.410 123.895 29.700 123.940 ;
        RECT 32.190 123.895 32.480 123.940 ;
        RECT 34.050 123.895 34.340 123.940 ;
        RECT 29.410 123.755 34.340 123.895 ;
        RECT 37.350 123.895 37.490 124.095 ;
        RECT 37.720 124.035 38.040 124.295 ;
        RECT 41.400 124.235 41.720 124.295 ;
        RECT 42.335 124.235 42.625 124.280 ;
        RECT 41.400 124.095 42.625 124.235 ;
        RECT 41.400 124.035 41.720 124.095 ;
        RECT 42.335 124.050 42.625 124.095 ;
        RECT 43.240 124.035 43.560 124.295 ;
        RECT 50.140 124.235 50.460 124.295 ;
        RECT 53.605 124.235 53.895 124.280 ;
        RECT 50.140 124.095 53.895 124.235 ;
        RECT 50.140 124.035 50.460 124.095 ;
        RECT 53.605 124.050 53.895 124.095 ;
        RECT 68.080 124.235 68.400 124.295 ;
        RECT 70.855 124.235 71.145 124.280 ;
        RECT 68.080 124.095 71.145 124.235 ;
        RECT 68.080 124.035 68.400 124.095 ;
        RECT 70.855 124.050 71.145 124.095 ;
        RECT 72.465 124.235 72.755 124.280 ;
        RECT 76.820 124.235 77.140 124.295 ;
        RECT 72.465 124.095 77.140 124.235 ;
        RECT 72.465 124.050 72.755 124.095 ;
        RECT 76.820 124.035 77.140 124.095 ;
        RECT 79.580 124.235 79.900 124.295 ;
        RECT 82.125 124.235 82.415 124.280 ;
        RECT 79.580 124.095 82.415 124.235 ;
        RECT 79.580 124.035 79.900 124.095 ;
        RECT 82.125 124.050 82.415 124.095 ;
        RECT 94.760 124.235 95.080 124.295 ;
        RECT 95.235 124.235 95.525 124.280 ;
        RECT 94.760 124.095 95.525 124.235 ;
        RECT 94.760 124.035 95.080 124.095 ;
        RECT 95.235 124.050 95.525 124.095 ;
        RECT 96.845 124.235 97.135 124.280 ;
        RECT 98.900 124.235 99.220 124.295 ;
        RECT 96.845 124.095 99.220 124.235 ;
        RECT 96.845 124.050 97.135 124.095 ;
        RECT 98.900 124.035 99.220 124.095 ;
        RECT 109.480 124.035 109.800 124.295 ;
        RECT 111.795 124.235 112.085 124.280 ;
        RECT 113.160 124.235 113.480 124.295 ;
        RECT 111.795 124.095 113.480 124.235 ;
        RECT 111.795 124.050 112.085 124.095 ;
        RECT 113.160 124.035 113.480 124.095 ;
        RECT 47.380 123.895 47.700 123.955 ;
        RECT 37.350 123.755 47.700 123.895 ;
        RECT 29.410 123.710 29.700 123.755 ;
        RECT 32.190 123.710 32.480 123.755 ;
        RECT 34.050 123.710 34.340 123.755 ;
        RECT 47.380 123.695 47.700 123.755 ;
        RECT 57.470 123.895 57.760 123.940 ;
        RECT 60.250 123.895 60.540 123.940 ;
        RECT 62.110 123.895 62.400 123.940 ;
        RECT 57.470 123.755 62.400 123.895 ;
        RECT 57.470 123.710 57.760 123.755 ;
        RECT 60.250 123.710 60.540 123.755 ;
        RECT 62.110 123.710 62.400 123.755 ;
        RECT 76.330 123.895 76.620 123.940 ;
        RECT 79.110 123.895 79.400 123.940 ;
        RECT 80.970 123.895 81.260 123.940 ;
        RECT 76.330 123.755 81.260 123.895 ;
        RECT 76.330 123.710 76.620 123.755 ;
        RECT 79.110 123.710 79.400 123.755 ;
        RECT 80.970 123.710 81.260 123.755 ;
        RECT 85.990 123.895 86.280 123.940 ;
        RECT 88.770 123.895 89.060 123.940 ;
        RECT 90.630 123.895 90.920 123.940 ;
        RECT 85.990 123.755 90.920 123.895 ;
        RECT 85.990 123.710 86.280 123.755 ;
        RECT 88.770 123.710 89.060 123.755 ;
        RECT 90.630 123.710 90.920 123.755 ;
        RECT 100.710 123.895 101.000 123.940 ;
        RECT 103.490 123.895 103.780 123.940 ;
        RECT 105.350 123.895 105.640 123.940 ;
        RECT 100.710 123.755 105.640 123.895 ;
        RECT 100.710 123.710 101.000 123.755 ;
        RECT 103.490 123.710 103.780 123.755 ;
        RECT 105.350 123.710 105.640 123.755 ;
        RECT 18.400 123.555 18.720 123.615 ;
        RECT 23.015 123.555 23.305 123.600 ;
        RECT 18.400 123.415 23.305 123.555 ;
        RECT 18.400 123.355 18.720 123.415 ;
        RECT 23.015 123.370 23.305 123.415 ;
        RECT 24.840 123.555 25.160 123.615 ;
        RECT 27.140 123.555 27.460 123.615 ;
        RECT 24.840 123.415 32.430 123.555 ;
        RECT 24.840 123.355 25.160 123.415 ;
        RECT 27.140 123.355 27.460 123.415 ;
        RECT 14.720 123.015 15.040 123.275 ;
        RECT 19.750 123.215 20.040 123.260 ;
        RECT 29.410 123.215 29.700 123.260 ;
        RECT 32.290 123.215 32.430 123.415 ;
        RECT 32.660 123.355 32.980 123.615 ;
        RECT 53.360 123.555 53.680 123.615 ;
        RECT 37.810 123.415 53.680 123.555 ;
        RECT 34.515 123.215 34.805 123.260 ;
        RECT 19.750 123.075 22.285 123.215 ;
        RECT 19.750 123.030 20.040 123.075 ;
        RECT 22.070 122.920 22.285 123.075 ;
        RECT 29.410 123.075 31.945 123.215 ;
        RECT 32.290 123.075 34.805 123.215 ;
        RECT 29.410 123.030 29.700 123.075 ;
        RECT 14.275 122.875 14.565 122.920 ;
        RECT 17.890 122.875 18.180 122.920 ;
        RECT 21.150 122.875 21.440 122.920 ;
        RECT 14.275 122.735 21.440 122.875 ;
        RECT 14.275 122.690 14.565 122.735 ;
        RECT 17.890 122.690 18.180 122.735 ;
        RECT 21.150 122.690 21.440 122.735 ;
        RECT 22.070 122.875 22.360 122.920 ;
        RECT 23.930 122.875 24.220 122.920 ;
        RECT 22.070 122.735 24.220 122.875 ;
        RECT 22.070 122.690 22.360 122.735 ;
        RECT 23.930 122.690 24.220 122.735 ;
        RECT 25.760 122.875 26.080 122.935 ;
        RECT 31.730 122.920 31.945 123.075 ;
        RECT 34.515 123.030 34.805 123.075 ;
        RECT 37.275 123.215 37.565 123.260 ;
        RECT 37.810 123.215 37.950 123.415 ;
        RECT 37.275 123.075 37.950 123.215 ;
        RECT 40.940 123.215 41.260 123.275 ;
        RECT 42.870 123.260 43.010 123.415 ;
        RECT 53.360 123.355 53.680 123.415 ;
        RECT 53.820 123.555 54.140 123.615 ;
        RECT 53.820 123.415 60.490 123.555 ;
        RECT 53.820 123.355 54.140 123.415 ;
        RECT 41.415 123.215 41.705 123.260 ;
        RECT 40.940 123.075 41.705 123.215 ;
        RECT 37.275 123.030 37.565 123.075 ;
        RECT 27.550 122.875 27.840 122.920 ;
        RECT 30.810 122.875 31.100 122.920 ;
        RECT 25.760 122.735 31.100 122.875 ;
        RECT 25.760 122.675 26.080 122.735 ;
        RECT 27.550 122.690 27.840 122.735 ;
        RECT 30.810 122.690 31.100 122.735 ;
        RECT 31.730 122.875 32.020 122.920 ;
        RECT 33.590 122.875 33.880 122.920 ;
        RECT 31.730 122.735 33.880 122.875 ;
        RECT 31.730 122.690 32.020 122.735 ;
        RECT 33.590 122.690 33.880 122.735 ;
        RECT 26.220 122.535 26.540 122.595 ;
        RECT 37.350 122.535 37.490 123.030 ;
        RECT 40.940 123.015 41.260 123.075 ;
        RECT 41.415 123.030 41.705 123.075 ;
        RECT 42.795 123.030 43.085 123.260 ;
        RECT 52.900 123.015 53.220 123.275 ;
        RECT 57.470 123.215 57.760 123.260 ;
        RECT 60.350 123.215 60.490 123.415 ;
        RECT 60.720 123.355 61.040 123.615 ;
        RECT 81.435 123.555 81.725 123.600 ;
        RECT 85.560 123.555 85.880 123.615 ;
        RECT 89.700 123.555 90.020 123.615 ;
        RECT 91.095 123.555 91.385 123.600 ;
        RECT 81.435 123.415 91.385 123.555 ;
        RECT 81.435 123.370 81.725 123.415 ;
        RECT 85.560 123.355 85.880 123.415 ;
        RECT 89.700 123.355 90.020 123.415 ;
        RECT 91.095 123.370 91.385 123.415 ;
        RECT 100.280 123.555 100.600 123.615 ;
        RECT 103.975 123.555 104.265 123.600 ;
        RECT 100.280 123.415 104.265 123.555 ;
        RECT 100.280 123.355 100.600 123.415 ;
        RECT 103.975 123.370 104.265 123.415 ;
        RECT 62.575 123.215 62.865 123.260 ;
        RECT 57.470 123.075 60.005 123.215 ;
        RECT 60.350 123.075 62.865 123.215 ;
        RECT 57.470 123.030 57.760 123.075 ;
        RECT 54.740 122.875 55.060 122.935 ;
        RECT 59.790 122.920 60.005 123.075 ;
        RECT 62.575 123.030 62.865 123.075 ;
        RECT 71.315 123.030 71.605 123.260 ;
        RECT 76.330 123.215 76.620 123.260 ;
        RECT 76.330 123.075 78.865 123.215 ;
        RECT 76.330 123.030 76.620 123.075 ;
        RECT 55.610 122.875 55.900 122.920 ;
        RECT 58.870 122.875 59.160 122.920 ;
        RECT 54.740 122.735 59.160 122.875 ;
        RECT 54.740 122.675 55.060 122.735 ;
        RECT 55.610 122.690 55.900 122.735 ;
        RECT 58.870 122.690 59.160 122.735 ;
        RECT 59.790 122.875 60.080 122.920 ;
        RECT 61.650 122.875 61.940 122.920 ;
        RECT 59.790 122.735 61.940 122.875 ;
        RECT 59.790 122.690 60.080 122.735 ;
        RECT 61.650 122.690 61.940 122.735 ;
        RECT 26.220 122.395 37.490 122.535 ;
        RECT 26.220 122.335 26.540 122.395 ;
        RECT 45.540 122.335 45.860 122.595 ;
        RECT 71.390 122.535 71.530 123.030 ;
        RECT 72.680 122.875 73.000 122.935 ;
        RECT 78.650 122.920 78.865 123.075 ;
        RECT 79.580 123.015 79.900 123.275 ;
        RECT 85.990 123.215 86.280 123.260 ;
        RECT 85.990 123.075 88.525 123.215 ;
        RECT 85.990 123.030 86.280 123.075 ;
        RECT 74.470 122.875 74.760 122.920 ;
        RECT 77.730 122.875 78.020 122.920 ;
        RECT 72.680 122.735 78.020 122.875 ;
        RECT 72.680 122.675 73.000 122.735 ;
        RECT 74.470 122.690 74.760 122.735 ;
        RECT 77.730 122.690 78.020 122.735 ;
        RECT 78.650 122.875 78.940 122.920 ;
        RECT 80.510 122.875 80.800 122.920 ;
        RECT 78.650 122.735 80.800 122.875 ;
        RECT 78.650 122.690 78.940 122.735 ;
        RECT 80.510 122.690 80.800 122.735 ;
        RECT 82.340 122.875 82.660 122.935 ;
        RECT 88.310 122.920 88.525 123.075 ;
        RECT 89.240 123.015 89.560 123.275 ;
        RECT 96.140 123.015 96.460 123.275 ;
        RECT 100.710 123.215 101.000 123.260 ;
        RECT 105.815 123.215 106.105 123.260 ;
        RECT 106.720 123.215 107.040 123.275 ;
        RECT 100.710 123.075 103.245 123.215 ;
        RECT 100.710 123.030 101.000 123.075 ;
        RECT 84.130 122.875 84.420 122.920 ;
        RECT 87.390 122.875 87.680 122.920 ;
        RECT 82.340 122.735 87.680 122.875 ;
        RECT 82.340 122.675 82.660 122.735 ;
        RECT 84.130 122.690 84.420 122.735 ;
        RECT 87.390 122.690 87.680 122.735 ;
        RECT 88.310 122.875 88.600 122.920 ;
        RECT 90.170 122.875 90.460 122.920 ;
        RECT 88.310 122.735 90.460 122.875 ;
        RECT 88.310 122.690 88.600 122.735 ;
        RECT 90.170 122.690 90.460 122.735 ;
        RECT 98.850 122.875 99.140 122.920 ;
        RECT 99.820 122.875 100.140 122.935 ;
        RECT 103.030 122.920 103.245 123.075 ;
        RECT 105.815 123.075 107.040 123.215 ;
        RECT 105.815 123.030 106.105 123.075 ;
        RECT 106.720 123.015 107.040 123.075 ;
        RECT 109.020 123.015 109.340 123.275 ;
        RECT 110.860 123.015 111.180 123.275 ;
        RECT 102.110 122.875 102.400 122.920 ;
        RECT 98.850 122.735 102.400 122.875 ;
        RECT 98.850 122.690 99.140 122.735 ;
        RECT 99.820 122.675 100.140 122.735 ;
        RECT 102.110 122.690 102.400 122.735 ;
        RECT 103.030 122.875 103.320 122.920 ;
        RECT 104.890 122.875 105.180 122.920 ;
        RECT 103.030 122.735 105.180 122.875 ;
        RECT 103.030 122.690 103.320 122.735 ;
        RECT 104.890 122.690 105.180 122.735 ;
        RECT 115.920 122.535 116.240 122.595 ;
        RECT 71.390 122.395 116.240 122.535 ;
        RECT 115.920 122.335 116.240 122.395 ;
        RECT 10.650 121.715 118.610 122.195 ;
        RECT 18.400 121.315 18.720 121.575 ;
        RECT 21.175 121.515 21.465 121.560 ;
        RECT 24.840 121.515 25.160 121.575 ;
        RECT 21.175 121.375 25.160 121.515 ;
        RECT 21.175 121.330 21.465 121.375 ;
        RECT 24.840 121.315 25.160 121.375 ;
        RECT 32.660 121.315 32.980 121.575 ;
        RECT 44.160 121.515 44.480 121.575 ;
        RECT 46.015 121.515 46.305 121.560 ;
        RECT 44.160 121.375 46.305 121.515 ;
        RECT 44.160 121.315 44.480 121.375 ;
        RECT 46.015 121.330 46.305 121.375 ;
        RECT 50.140 121.515 50.460 121.575 ;
        RECT 50.615 121.515 50.905 121.560 ;
        RECT 50.140 121.375 50.905 121.515 ;
        RECT 27.600 120.975 27.920 121.235 ;
        RECT 46.090 121.175 46.230 121.330 ;
        RECT 50.140 121.315 50.460 121.375 ;
        RECT 50.615 121.330 50.905 121.375 ;
        RECT 52.915 121.515 53.205 121.560 ;
        RECT 54.280 121.515 54.600 121.575 ;
        RECT 52.915 121.375 54.600 121.515 ;
        RECT 52.915 121.330 53.205 121.375 ;
        RECT 54.280 121.315 54.600 121.375 ;
        RECT 54.740 121.315 55.060 121.575 ;
        RECT 56.595 121.515 56.885 121.560 ;
        RECT 60.720 121.515 61.040 121.575 ;
        RECT 56.595 121.375 61.040 121.515 ;
        RECT 56.595 121.330 56.885 121.375 ;
        RECT 60.720 121.315 61.040 121.375 ;
        RECT 79.135 121.515 79.425 121.560 ;
        RECT 79.580 121.515 79.900 121.575 ;
        RECT 79.135 121.375 79.900 121.515 ;
        RECT 79.135 121.330 79.425 121.375 ;
        RECT 79.580 121.315 79.900 121.375 ;
        RECT 89.240 121.315 89.560 121.575 ;
        RECT 115.920 121.315 116.240 121.575 ;
        RECT 51.075 121.175 51.365 121.220 ;
        RECT 46.090 121.035 51.365 121.175 ;
        RECT 51.075 120.990 51.365 121.035 ;
        RECT 53.360 121.175 53.680 121.235 ;
        RECT 57.975 121.175 58.265 121.220 ;
        RECT 53.360 121.035 58.265 121.175 ;
        RECT 53.360 120.975 53.680 121.035 ;
        RECT 17.495 120.835 17.785 120.880 ;
        RECT 17.940 120.835 18.260 120.895 ;
        RECT 17.495 120.695 18.260 120.835 ;
        RECT 17.495 120.650 17.785 120.695 ;
        RECT 17.940 120.635 18.260 120.695 ;
        RECT 31.755 120.835 32.045 120.880 ;
        RECT 32.200 120.835 32.520 120.895 ;
        RECT 31.755 120.695 32.520 120.835 ;
        RECT 31.755 120.650 32.045 120.695 ;
        RECT 32.200 120.635 32.520 120.695 ;
        RECT 39.100 120.835 39.420 120.895 ;
        RECT 54.370 120.880 54.510 121.035 ;
        RECT 57.975 120.990 58.265 121.035 ;
        RECT 46.475 120.835 46.765 120.880 ;
        RECT 39.100 120.695 46.765 120.835 ;
        RECT 39.100 120.635 39.420 120.695 ;
        RECT 46.475 120.650 46.765 120.695 ;
        RECT 54.295 120.650 54.585 120.880 ;
        RECT 55.660 120.635 55.980 120.895 ;
        RECT 59.355 120.835 59.645 120.880 ;
        RECT 60.260 120.835 60.580 120.895 ;
        RECT 59.355 120.695 60.580 120.835 ;
        RECT 59.355 120.650 59.645 120.695 ;
        RECT 60.260 120.635 60.580 120.695 ;
        RECT 72.680 120.635 73.000 120.895 ;
        RECT 73.155 120.835 73.445 120.880 ;
        RECT 74.060 120.835 74.380 120.895 ;
        RECT 73.155 120.695 74.380 120.835 ;
        RECT 73.155 120.650 73.445 120.695 ;
        RECT 74.060 120.635 74.380 120.695 ;
        RECT 77.280 120.835 77.600 120.895 ;
        RECT 78.215 120.835 78.505 120.880 ;
        RECT 77.280 120.695 78.505 120.835 ;
        RECT 77.280 120.635 77.600 120.695 ;
        RECT 78.215 120.650 78.505 120.695 ;
        RECT 86.940 120.835 87.260 120.895 ;
        RECT 88.335 120.835 88.625 120.880 ;
        RECT 86.940 120.695 88.625 120.835 ;
        RECT 86.940 120.635 87.260 120.695 ;
        RECT 88.335 120.650 88.625 120.695 ;
        RECT 110.875 120.650 111.165 120.880 ;
        RECT 45.555 120.495 45.845 120.540 ;
        RECT 49.680 120.495 50.000 120.555 ;
        RECT 45.555 120.355 50.000 120.495 ;
        RECT 45.555 120.310 45.845 120.355 ;
        RECT 49.680 120.295 50.000 120.355 ;
        RECT 107.180 120.495 107.500 120.555 ;
        RECT 110.950 120.495 111.090 120.650 ;
        RECT 111.320 120.635 111.640 120.895 ;
        RECT 111.780 120.835 112.100 120.895 ;
        RECT 113.175 120.835 113.465 120.880 ;
        RECT 111.780 120.695 113.465 120.835 ;
        RECT 111.780 120.635 112.100 120.695 ;
        RECT 113.175 120.650 113.465 120.695 ;
        RECT 116.840 120.635 117.160 120.895 ;
        RECT 107.180 120.355 111.090 120.495 ;
        RECT 107.180 120.295 107.500 120.355 ;
        RECT 48.300 119.615 48.620 119.875 ;
        RECT 108.100 119.815 108.420 119.875 ;
        RECT 114.095 119.815 114.385 119.860 ;
        RECT 108.100 119.675 114.385 119.815 ;
        RECT 108.100 119.615 108.420 119.675 ;
        RECT 114.095 119.630 114.385 119.675 ;
        RECT 11.430 118.995 118.610 119.475 ;
        RECT 35.420 118.795 35.740 118.855 ;
        RECT 35.420 118.655 47.150 118.795 ;
        RECT 35.420 118.595 35.740 118.655 ;
        RECT 34.615 118.455 34.905 118.500 ;
        RECT 37.735 118.455 38.025 118.500 ;
        RECT 39.625 118.455 39.915 118.500 ;
        RECT 34.615 118.315 39.915 118.455 ;
        RECT 34.615 118.270 34.905 118.315 ;
        RECT 37.735 118.270 38.025 118.315 ;
        RECT 39.625 118.270 39.915 118.315 ;
        RECT 30.375 118.115 30.665 118.160 ;
        RECT 34.040 118.115 34.360 118.175 ;
        RECT 30.375 117.975 34.360 118.115 ;
        RECT 30.375 117.930 30.665 117.975 ;
        RECT 34.040 117.915 34.360 117.975 ;
        RECT 39.100 118.115 39.420 118.175 ;
        RECT 40.480 118.115 40.800 118.175 ;
        RECT 39.100 117.975 40.800 118.115 ;
        RECT 39.100 117.915 39.420 117.975 ;
        RECT 40.480 117.915 40.800 117.975 ;
        RECT 24.855 117.775 25.145 117.820 ;
        RECT 28.980 117.775 29.300 117.835 ;
        RECT 24.855 117.635 29.300 117.775 ;
        RECT 24.855 117.590 25.145 117.635 ;
        RECT 28.980 117.575 29.300 117.635 ;
        RECT 30.360 117.435 30.680 117.495 ;
        RECT 33.535 117.480 33.825 117.795 ;
        RECT 34.615 117.775 34.905 117.820 ;
        RECT 38.195 117.775 38.485 117.820 ;
        RECT 40.030 117.775 40.320 117.820 ;
        RECT 34.615 117.635 40.320 117.775 ;
        RECT 34.615 117.590 34.905 117.635 ;
        RECT 38.195 117.590 38.485 117.635 ;
        RECT 40.030 117.590 40.320 117.635 ;
        RECT 41.860 117.775 42.180 117.835 ;
        RECT 42.335 117.775 42.625 117.820 ;
        RECT 41.860 117.635 42.625 117.775 ;
        RECT 41.860 117.575 42.180 117.635 ;
        RECT 42.335 117.590 42.625 117.635 ;
        RECT 43.700 117.575 44.020 117.835 ;
        RECT 47.010 117.820 47.150 118.655 ;
        RECT 49.220 118.595 49.540 118.855 ;
        RECT 107.180 118.795 107.500 118.855 ;
        RECT 108.560 118.795 108.880 118.855 ;
        RECT 107.180 118.655 108.880 118.795 ;
        RECT 107.180 118.595 107.500 118.655 ;
        RECT 108.560 118.595 108.880 118.655 ;
        RECT 69.920 118.455 70.240 118.515 ;
        RECT 107.270 118.455 107.410 118.595 ;
        RECT 69.920 118.315 74.290 118.455 ;
        RECT 69.920 118.255 70.240 118.315 ;
        RECT 71.315 118.115 71.605 118.160 ;
        RECT 73.600 118.115 73.920 118.175 ;
        RECT 69.550 117.975 73.920 118.115 ;
        RECT 46.935 117.590 47.225 117.820 ;
        RECT 48.300 117.575 48.620 117.835 ;
        RECT 57.515 117.775 57.805 117.820 ;
        RECT 59.340 117.775 59.660 117.835 ;
        RECT 59.815 117.775 60.105 117.820 ;
        RECT 57.515 117.635 60.105 117.775 ;
        RECT 57.515 117.590 57.805 117.635 ;
        RECT 59.340 117.575 59.660 117.635 ;
        RECT 59.815 117.590 60.105 117.635 ;
        RECT 60.260 117.775 60.580 117.835 ;
        RECT 61.195 117.775 61.485 117.820 ;
        RECT 60.260 117.635 61.485 117.775 ;
        RECT 60.260 117.575 60.580 117.635 ;
        RECT 61.195 117.590 61.485 117.635 ;
        RECT 61.640 117.775 61.960 117.835 ;
        RECT 69.550 117.820 69.690 117.975 ;
        RECT 71.315 117.930 71.605 117.975 ;
        RECT 73.600 117.915 73.920 117.975 ;
        RECT 63.495 117.775 63.785 117.820 ;
        RECT 61.640 117.635 63.785 117.775 ;
        RECT 33.235 117.435 33.825 117.480 ;
        RECT 36.475 117.435 37.125 117.480 ;
        RECT 30.360 117.295 37.125 117.435 ;
        RECT 30.360 117.235 30.680 117.295 ;
        RECT 33.235 117.250 33.525 117.295 ;
        RECT 36.475 117.250 37.125 117.295 ;
        RECT 39.115 117.435 39.405 117.480 ;
        RECT 61.270 117.435 61.410 117.590 ;
        RECT 61.640 117.575 61.960 117.635 ;
        RECT 63.495 117.590 63.785 117.635 ;
        RECT 69.475 117.590 69.765 117.820 ;
        RECT 69.935 117.590 70.225 117.820 ;
        RECT 72.220 117.775 72.540 117.835 ;
        RECT 74.150 117.820 74.290 118.315 ;
        RECT 103.130 118.315 107.410 118.455 ;
        RECT 107.605 118.455 107.895 118.500 ;
        RECT 109.495 118.455 109.785 118.500 ;
        RECT 112.615 118.455 112.905 118.500 ;
        RECT 107.605 118.315 112.905 118.455 ;
        RECT 93.380 118.115 93.700 118.175 ;
        RECT 103.130 118.115 103.270 118.315 ;
        RECT 107.605 118.270 107.895 118.315 ;
        RECT 109.495 118.270 109.785 118.315 ;
        RECT 112.615 118.270 112.905 118.315 ;
        RECT 93.380 117.975 103.270 118.115 ;
        RECT 93.380 117.915 93.700 117.975 ;
        RECT 72.695 117.775 72.985 117.820 ;
        RECT 72.220 117.635 72.985 117.775 ;
        RECT 70.010 117.435 70.150 117.590 ;
        RECT 72.220 117.575 72.540 117.635 ;
        RECT 72.695 117.590 72.985 117.635 ;
        RECT 74.075 117.590 74.365 117.820 ;
        RECT 75.900 117.775 76.220 117.835 ;
        RECT 77.755 117.775 78.045 117.820 ;
        RECT 75.900 117.635 78.045 117.775 ;
        RECT 75.900 117.575 76.220 117.635 ;
        RECT 77.755 117.590 78.045 117.635 ;
        RECT 85.115 117.590 85.405 117.820 ;
        RECT 95.680 117.775 96.000 117.835 ;
        RECT 100.830 117.820 100.970 117.975 ;
        RECT 97.995 117.775 98.285 117.820 ;
        RECT 95.680 117.635 98.285 117.775 ;
        RECT 39.115 117.295 43.010 117.435 ;
        RECT 61.270 117.295 70.150 117.435 ;
        RECT 70.380 117.435 70.700 117.495 ;
        RECT 85.190 117.435 85.330 117.590 ;
        RECT 95.680 117.575 96.000 117.635 ;
        RECT 97.995 117.590 98.285 117.635 ;
        RECT 100.755 117.590 101.045 117.820 ;
        RECT 101.200 117.575 101.520 117.835 ;
        RECT 103.130 117.775 103.270 117.975 ;
        RECT 103.500 118.115 103.820 118.175 ;
        RECT 103.500 117.975 105.570 118.115 ;
        RECT 103.500 117.915 103.820 117.975 ;
        RECT 105.430 117.820 105.570 117.975 ;
        RECT 108.100 117.915 108.420 118.175 ;
        RECT 103.975 117.775 104.265 117.820 ;
        RECT 103.130 117.635 104.265 117.775 ;
        RECT 103.975 117.590 104.265 117.635 ;
        RECT 105.355 117.590 105.645 117.820 ;
        RECT 106.720 117.575 107.040 117.835 ;
        RECT 107.200 117.775 107.490 117.820 ;
        RECT 109.035 117.775 109.325 117.820 ;
        RECT 112.615 117.775 112.905 117.820 ;
        RECT 107.200 117.635 112.905 117.775 ;
        RECT 107.200 117.590 107.490 117.635 ;
        RECT 109.035 117.590 109.325 117.635 ;
        RECT 112.615 117.590 112.905 117.635 ;
        RECT 70.380 117.295 85.330 117.435 ;
        RECT 110.395 117.435 111.045 117.480 ;
        RECT 111.320 117.435 111.640 117.495 ;
        RECT 113.695 117.480 113.985 117.795 ;
        RECT 113.695 117.435 114.285 117.480 ;
        RECT 110.395 117.295 114.285 117.435 ;
        RECT 39.115 117.250 39.405 117.295 ;
        RECT 23.460 117.095 23.780 117.155 ;
        RECT 23.935 117.095 24.225 117.140 ;
        RECT 23.460 116.955 24.225 117.095 ;
        RECT 23.460 116.895 23.780 116.955 ;
        RECT 23.935 116.910 24.225 116.955 ;
        RECT 41.400 116.895 41.720 117.155 ;
        RECT 42.870 117.140 43.010 117.295 ;
        RECT 70.380 117.235 70.700 117.295 ;
        RECT 110.395 117.250 111.045 117.295 ;
        RECT 111.320 117.235 111.640 117.295 ;
        RECT 113.995 117.250 114.285 117.295 ;
        RECT 116.855 117.435 117.145 117.480 ;
        RECT 117.300 117.435 117.620 117.495 ;
        RECT 116.855 117.295 117.620 117.435 ;
        RECT 116.855 117.250 117.145 117.295 ;
        RECT 117.300 117.235 117.620 117.295 ;
        RECT 42.795 116.910 43.085 117.140 ;
        RECT 47.855 117.095 48.145 117.140 ;
        RECT 51.980 117.095 52.300 117.155 ;
        RECT 47.855 116.955 52.300 117.095 ;
        RECT 47.855 116.910 48.145 116.955 ;
        RECT 51.980 116.895 52.300 116.955 ;
        RECT 57.960 116.895 58.280 117.155 ;
        RECT 64.415 117.095 64.705 117.140 ;
        RECT 66.240 117.095 66.560 117.155 ;
        RECT 64.415 116.955 66.560 117.095 ;
        RECT 64.415 116.910 64.705 116.955 ;
        RECT 66.240 116.895 66.560 116.955 ;
        RECT 69.000 116.895 69.320 117.155 ;
        RECT 73.600 116.895 73.920 117.155 ;
        RECT 74.995 117.095 75.285 117.140 ;
        RECT 76.360 117.095 76.680 117.155 ;
        RECT 74.995 116.955 76.680 117.095 ;
        RECT 74.995 116.910 75.285 116.955 ;
        RECT 76.360 116.895 76.680 116.955 ;
        RECT 78.675 117.095 78.965 117.140 ;
        RECT 79.580 117.095 79.900 117.155 ;
        RECT 78.675 116.955 79.900 117.095 ;
        RECT 78.675 116.910 78.965 116.955 ;
        RECT 79.580 116.895 79.900 116.955 ;
        RECT 86.035 117.095 86.325 117.140 ;
        RECT 88.780 117.095 89.100 117.155 ;
        RECT 86.035 116.955 89.100 117.095 ;
        RECT 86.035 116.910 86.325 116.955 ;
        RECT 88.780 116.895 89.100 116.955 ;
        RECT 98.900 116.895 99.220 117.155 ;
        RECT 100.280 116.895 100.600 117.155 ;
        RECT 102.120 116.895 102.440 117.155 ;
        RECT 103.960 117.095 104.280 117.155 ;
        RECT 104.435 117.095 104.725 117.140 ;
        RECT 103.960 116.955 104.725 117.095 ;
        RECT 103.960 116.895 104.280 116.955 ;
        RECT 104.435 116.910 104.725 116.955 ;
        RECT 106.275 117.095 106.565 117.140 ;
        RECT 112.240 117.095 112.560 117.155 ;
        RECT 106.275 116.955 112.560 117.095 ;
        RECT 106.275 116.910 106.565 116.955 ;
        RECT 112.240 116.895 112.560 116.955 ;
        RECT 10.650 116.275 118.610 116.755 ;
        RECT 26.695 116.075 26.985 116.120 ;
        RECT 24.930 115.935 26.985 116.075 ;
        RECT 17.480 115.735 17.800 115.795 ;
        RECT 24.930 115.780 25.070 115.935 ;
        RECT 26.695 115.890 26.985 115.935 ;
        RECT 30.360 115.875 30.680 116.135 ;
        RECT 73.600 116.075 73.920 116.135 ;
        RECT 84.180 116.075 84.500 116.135 ;
        RECT 73.600 115.935 77.050 116.075 ;
        RECT 73.600 115.875 73.920 115.935 ;
        RECT 18.975 115.735 19.265 115.780 ;
        RECT 22.215 115.735 22.865 115.780 ;
        RECT 17.480 115.595 22.865 115.735 ;
        RECT 17.480 115.535 17.800 115.595 ;
        RECT 18.975 115.550 19.565 115.595 ;
        RECT 22.215 115.550 22.865 115.595 ;
        RECT 24.855 115.550 25.145 115.780 ;
        RECT 35.535 115.735 35.825 115.780 ;
        RECT 38.180 115.735 38.500 115.795 ;
        RECT 38.775 115.735 39.425 115.780 ;
        RECT 35.535 115.595 39.425 115.735 ;
        RECT 35.535 115.550 36.125 115.595 ;
        RECT 19.275 115.235 19.565 115.550 ;
        RECT 20.355 115.395 20.645 115.440 ;
        RECT 23.935 115.395 24.225 115.440 ;
        RECT 25.770 115.395 26.060 115.440 ;
        RECT 20.355 115.255 26.060 115.395 ;
        RECT 20.355 115.210 20.645 115.255 ;
        RECT 23.935 115.210 24.225 115.255 ;
        RECT 25.770 115.210 26.060 115.255 ;
        RECT 26.235 115.395 26.525 115.440 ;
        RECT 27.140 115.395 27.460 115.455 ;
        RECT 26.235 115.255 27.460 115.395 ;
        RECT 26.235 115.210 26.525 115.255 ;
        RECT 27.140 115.195 27.460 115.255 ;
        RECT 27.615 115.395 27.905 115.440 ;
        RECT 28.060 115.395 28.380 115.455 ;
        RECT 27.615 115.255 28.380 115.395 ;
        RECT 27.615 115.210 27.905 115.255 ;
        RECT 28.060 115.195 28.380 115.255 ;
        RECT 28.535 115.395 28.825 115.440 ;
        RECT 29.900 115.395 30.220 115.455 ;
        RECT 28.535 115.255 30.220 115.395 ;
        RECT 28.535 115.210 28.825 115.255 ;
        RECT 29.900 115.195 30.220 115.255 ;
        RECT 32.200 115.195 32.520 115.455 ;
        RECT 35.835 115.235 36.125 115.550 ;
        RECT 38.180 115.535 38.500 115.595 ;
        RECT 38.775 115.550 39.425 115.595 ;
        RECT 41.400 115.535 41.720 115.795 ;
        RECT 46.115 115.735 46.405 115.780 ;
        RECT 48.300 115.735 48.620 115.795 ;
        RECT 49.355 115.735 50.005 115.780 ;
        RECT 46.115 115.595 50.005 115.735 ;
        RECT 46.115 115.550 46.705 115.595 ;
        RECT 36.915 115.395 37.205 115.440 ;
        RECT 40.495 115.395 40.785 115.440 ;
        RECT 42.330 115.395 42.620 115.440 ;
        RECT 36.915 115.255 42.620 115.395 ;
        RECT 36.915 115.210 37.205 115.255 ;
        RECT 40.495 115.210 40.785 115.255 ;
        RECT 42.330 115.210 42.620 115.255 ;
        RECT 42.795 115.395 43.085 115.440 ;
        RECT 45.540 115.395 45.860 115.455 ;
        RECT 42.795 115.255 45.860 115.395 ;
        RECT 42.795 115.210 43.085 115.255 ;
        RECT 45.540 115.195 45.860 115.255 ;
        RECT 46.415 115.235 46.705 115.550 ;
        RECT 48.300 115.535 48.620 115.595 ;
        RECT 49.355 115.550 50.005 115.595 ;
        RECT 51.980 115.535 52.300 115.795 ;
        RECT 57.960 115.735 58.280 115.795 ;
        RECT 60.375 115.735 60.665 115.780 ;
        RECT 63.615 115.735 64.265 115.780 ;
        RECT 57.960 115.595 64.265 115.735 ;
        RECT 57.960 115.535 58.280 115.595 ;
        RECT 60.375 115.550 60.965 115.595 ;
        RECT 63.615 115.550 64.265 115.595 ;
        RECT 47.495 115.395 47.785 115.440 ;
        RECT 51.075 115.395 51.365 115.440 ;
        RECT 52.910 115.395 53.200 115.440 ;
        RECT 47.495 115.255 53.200 115.395 ;
        RECT 47.495 115.210 47.785 115.255 ;
        RECT 51.075 115.210 51.365 115.255 ;
        RECT 52.910 115.210 53.200 115.255 ;
        RECT 55.200 115.195 55.520 115.455 ;
        RECT 56.120 115.195 56.440 115.455 ;
        RECT 60.675 115.235 60.965 115.550 ;
        RECT 66.240 115.535 66.560 115.795 ;
        RECT 67.620 115.735 67.940 115.795 ;
        RECT 68.095 115.735 68.385 115.780 ;
        RECT 67.620 115.595 68.385 115.735 ;
        RECT 67.620 115.535 67.940 115.595 ;
        RECT 68.095 115.550 68.385 115.595 ;
        RECT 69.000 115.735 69.320 115.795 ;
        RECT 76.910 115.780 77.050 115.935 ;
        RECT 80.130 115.935 84.500 116.075 ;
        RECT 80.130 115.780 80.270 115.935 ;
        RECT 84.180 115.875 84.500 115.935 ;
        RECT 86.480 115.780 86.800 115.795 ;
        RECT 70.955 115.735 71.245 115.780 ;
        RECT 74.195 115.735 74.845 115.780 ;
        RECT 69.000 115.595 74.845 115.735 ;
        RECT 69.000 115.535 69.320 115.595 ;
        RECT 70.955 115.550 71.545 115.595 ;
        RECT 74.195 115.550 74.845 115.595 ;
        RECT 76.835 115.550 77.125 115.780 ;
        RECT 80.055 115.550 80.345 115.780 ;
        RECT 82.915 115.735 83.205 115.780 ;
        RECT 86.155 115.735 86.805 115.780 ;
        RECT 82.915 115.595 86.805 115.735 ;
        RECT 82.915 115.550 83.505 115.595 ;
        RECT 86.155 115.550 86.805 115.595 ;
        RECT 61.755 115.395 62.045 115.440 ;
        RECT 65.335 115.395 65.625 115.440 ;
        RECT 67.170 115.395 67.460 115.440 ;
        RECT 61.755 115.255 67.460 115.395 ;
        RECT 61.755 115.210 62.045 115.255 ;
        RECT 65.335 115.210 65.625 115.255 ;
        RECT 67.170 115.210 67.460 115.255 ;
        RECT 71.255 115.235 71.545 115.550 ;
        RECT 72.335 115.395 72.625 115.440 ;
        RECT 75.915 115.395 76.205 115.440 ;
        RECT 77.750 115.395 78.040 115.440 ;
        RECT 72.335 115.255 78.040 115.395 ;
        RECT 72.335 115.210 72.625 115.255 ;
        RECT 75.915 115.210 76.205 115.255 ;
        RECT 77.750 115.210 78.040 115.255 ;
        RECT 83.215 115.235 83.505 115.550 ;
        RECT 86.480 115.535 86.800 115.550 ;
        RECT 88.780 115.535 89.100 115.795 ;
        RECT 90.160 115.735 90.480 115.795 ;
        RECT 97.635 115.735 97.925 115.780 ;
        RECT 100.280 115.735 100.600 115.795 ;
        RECT 100.875 115.735 101.525 115.780 ;
        RECT 90.160 115.595 93.150 115.735 ;
        RECT 90.160 115.535 90.480 115.595 ;
        RECT 93.010 115.440 93.150 115.595 ;
        RECT 97.635 115.595 101.525 115.735 ;
        RECT 97.635 115.550 98.225 115.595 ;
        RECT 84.295 115.395 84.585 115.440 ;
        RECT 87.875 115.395 88.165 115.440 ;
        RECT 89.710 115.395 90.000 115.440 ;
        RECT 84.295 115.255 90.000 115.395 ;
        RECT 84.295 115.210 84.585 115.255 ;
        RECT 87.875 115.210 88.165 115.255 ;
        RECT 89.710 115.210 90.000 115.255 ;
        RECT 92.935 115.210 93.225 115.440 ;
        RECT 93.380 115.195 93.700 115.455 ;
        RECT 97.935 115.235 98.225 115.550 ;
        RECT 100.280 115.535 100.600 115.595 ;
        RECT 100.875 115.550 101.525 115.595 ;
        RECT 102.120 115.735 102.440 115.795 ;
        RECT 103.515 115.735 103.805 115.780 ;
        RECT 102.120 115.595 103.805 115.735 ;
        RECT 102.120 115.535 102.440 115.595 ;
        RECT 103.515 115.550 103.805 115.595 ;
        RECT 106.735 115.735 107.025 115.780 ;
        RECT 109.595 115.735 109.885 115.780 ;
        RECT 110.400 115.735 110.720 115.795 ;
        RECT 112.835 115.735 113.485 115.780 ;
        RECT 106.735 115.595 107.640 115.735 ;
        RECT 106.735 115.550 107.025 115.595 ;
        RECT 99.015 115.395 99.305 115.440 ;
        RECT 102.595 115.395 102.885 115.440 ;
        RECT 104.430 115.395 104.720 115.440 ;
        RECT 99.015 115.255 104.720 115.395 ;
        RECT 99.015 115.210 99.305 115.255 ;
        RECT 102.595 115.210 102.885 115.255 ;
        RECT 104.430 115.210 104.720 115.255 ;
        RECT 16.115 115.055 16.405 115.100 ;
        RECT 17.940 115.055 18.260 115.115 ;
        RECT 16.115 114.915 18.260 115.055 ;
        RECT 16.115 114.870 16.405 114.915 ;
        RECT 17.940 114.855 18.260 114.915 ;
        RECT 32.675 115.055 32.965 115.100 ;
        RECT 39.560 115.055 39.880 115.115 ;
        RECT 32.675 114.915 39.880 115.055 ;
        RECT 32.675 114.870 32.965 114.915 ;
        RECT 39.560 114.855 39.880 114.915 ;
        RECT 43.255 114.870 43.545 115.100 ;
        RECT 45.630 115.055 45.770 115.195 ;
        RECT 53.375 115.055 53.665 115.100 ;
        RECT 53.820 115.055 54.140 115.115 ;
        RECT 45.630 114.915 54.140 115.055 ;
        RECT 53.375 114.870 53.665 114.915 ;
        RECT 20.355 114.715 20.645 114.760 ;
        RECT 23.475 114.715 23.765 114.760 ;
        RECT 25.365 114.715 25.655 114.760 ;
        RECT 20.355 114.575 25.655 114.715 ;
        RECT 20.355 114.530 20.645 114.575 ;
        RECT 23.475 114.530 23.765 114.575 ;
        RECT 25.365 114.530 25.655 114.575 ;
        RECT 36.915 114.715 37.205 114.760 ;
        RECT 40.035 114.715 40.325 114.760 ;
        RECT 41.925 114.715 42.215 114.760 ;
        RECT 36.915 114.575 42.215 114.715 ;
        RECT 43.330 114.715 43.470 114.870 ;
        RECT 53.820 114.855 54.140 114.915 ;
        RECT 57.515 115.055 57.805 115.100 ;
        RECT 61.180 115.055 61.500 115.115 ;
        RECT 57.515 114.915 61.500 115.055 ;
        RECT 57.515 114.870 57.805 114.915 ;
        RECT 61.180 114.855 61.500 114.915 ;
        RECT 64.400 115.055 64.720 115.115 ;
        RECT 67.635 115.055 67.925 115.100 ;
        RECT 64.400 114.915 67.925 115.055 ;
        RECT 64.400 114.855 64.720 114.915 ;
        RECT 67.635 114.870 67.925 114.915 ;
        RECT 78.215 115.055 78.505 115.100 ;
        RECT 80.040 115.055 80.360 115.115 ;
        RECT 85.560 115.055 85.880 115.115 ;
        RECT 90.175 115.055 90.465 115.100 ;
        RECT 78.215 114.915 90.465 115.055 ;
        RECT 78.215 114.870 78.505 114.915 ;
        RECT 80.040 114.855 80.360 114.915 ;
        RECT 85.560 114.855 85.880 114.915 ;
        RECT 90.175 114.870 90.465 114.915 ;
        RECT 94.775 115.055 95.065 115.100 ;
        RECT 100.740 115.055 101.060 115.115 ;
        RECT 94.775 114.915 101.060 115.055 ;
        RECT 94.775 114.870 95.065 114.915 ;
        RECT 100.740 114.855 101.060 114.915 ;
        RECT 103.040 115.055 103.360 115.115 ;
        RECT 104.895 115.055 105.185 115.100 ;
        RECT 106.720 115.055 107.040 115.115 ;
        RECT 103.040 114.915 107.040 115.055 ;
        RECT 107.500 115.055 107.640 115.595 ;
        RECT 109.595 115.595 113.485 115.735 ;
        RECT 109.595 115.550 110.185 115.595 ;
        RECT 109.895 115.235 110.185 115.550 ;
        RECT 110.400 115.535 110.720 115.595 ;
        RECT 112.835 115.550 113.485 115.595 ;
        RECT 115.000 115.735 115.320 115.795 ;
        RECT 115.475 115.735 115.765 115.780 ;
        RECT 115.000 115.595 115.765 115.735 ;
        RECT 115.000 115.535 115.320 115.595 ;
        RECT 115.475 115.550 115.765 115.595 ;
        RECT 110.975 115.395 111.265 115.440 ;
        RECT 114.555 115.395 114.845 115.440 ;
        RECT 116.390 115.395 116.680 115.440 ;
        RECT 110.975 115.255 116.680 115.395 ;
        RECT 110.975 115.210 111.265 115.255 ;
        RECT 114.555 115.210 114.845 115.255 ;
        RECT 116.390 115.210 116.680 115.255 ;
        RECT 111.780 115.055 112.100 115.115 ;
        RECT 107.500 114.915 112.100 115.055 ;
        RECT 103.040 114.855 103.360 114.915 ;
        RECT 104.895 114.870 105.185 114.915 ;
        RECT 106.720 114.855 107.040 114.915 ;
        RECT 111.780 114.855 112.100 114.915 ;
        RECT 115.460 115.055 115.780 115.115 ;
        RECT 116.855 115.055 117.145 115.100 ;
        RECT 115.460 114.915 117.145 115.055 ;
        RECT 115.460 114.855 115.780 114.915 ;
        RECT 116.855 114.870 117.145 114.915 ;
        RECT 45.540 114.715 45.860 114.775 ;
        RECT 43.330 114.575 45.860 114.715 ;
        RECT 36.915 114.530 37.205 114.575 ;
        RECT 40.035 114.530 40.325 114.575 ;
        RECT 41.925 114.530 42.215 114.575 ;
        RECT 45.540 114.515 45.860 114.575 ;
        RECT 47.495 114.715 47.785 114.760 ;
        RECT 50.615 114.715 50.905 114.760 ;
        RECT 52.505 114.715 52.795 114.760 ;
        RECT 47.495 114.575 52.795 114.715 ;
        RECT 47.495 114.530 47.785 114.575 ;
        RECT 50.615 114.530 50.905 114.575 ;
        RECT 52.505 114.530 52.795 114.575 ;
        RECT 61.755 114.715 62.045 114.760 ;
        RECT 64.875 114.715 65.165 114.760 ;
        RECT 66.765 114.715 67.055 114.760 ;
        RECT 61.755 114.575 67.055 114.715 ;
        RECT 61.755 114.530 62.045 114.575 ;
        RECT 64.875 114.530 65.165 114.575 ;
        RECT 66.765 114.530 67.055 114.575 ;
        RECT 72.335 114.715 72.625 114.760 ;
        RECT 75.455 114.715 75.745 114.760 ;
        RECT 77.345 114.715 77.635 114.760 ;
        RECT 72.335 114.575 77.635 114.715 ;
        RECT 72.335 114.530 72.625 114.575 ;
        RECT 75.455 114.530 75.745 114.575 ;
        RECT 77.345 114.530 77.635 114.575 ;
        RECT 84.295 114.715 84.585 114.760 ;
        RECT 87.415 114.715 87.705 114.760 ;
        RECT 89.305 114.715 89.595 114.760 ;
        RECT 84.295 114.575 89.595 114.715 ;
        RECT 84.295 114.530 84.585 114.575 ;
        RECT 87.415 114.530 87.705 114.575 ;
        RECT 89.305 114.530 89.595 114.575 ;
        RECT 99.015 114.715 99.305 114.760 ;
        RECT 102.135 114.715 102.425 114.760 ;
        RECT 104.025 114.715 104.315 114.760 ;
        RECT 99.015 114.575 104.315 114.715 ;
        RECT 99.015 114.530 99.305 114.575 ;
        RECT 102.135 114.530 102.425 114.575 ;
        RECT 104.025 114.530 104.315 114.575 ;
        RECT 110.975 114.715 111.265 114.760 ;
        RECT 114.095 114.715 114.385 114.760 ;
        RECT 115.985 114.715 116.275 114.760 ;
        RECT 110.975 114.575 116.275 114.715 ;
        RECT 110.975 114.530 111.265 114.575 ;
        RECT 114.095 114.530 114.385 114.575 ;
        RECT 115.985 114.530 116.275 114.575 ;
        RECT 28.995 114.375 29.285 114.420 ;
        RECT 29.440 114.375 29.760 114.435 ;
        RECT 28.995 114.235 29.760 114.375 ;
        RECT 28.995 114.190 29.285 114.235 ;
        RECT 29.440 114.175 29.760 114.235 ;
        RECT 31.280 114.175 31.600 114.435 ;
        RECT 52.900 114.375 53.220 114.435 ;
        RECT 54.295 114.375 54.585 114.420 ;
        RECT 52.900 114.235 54.585 114.375 ;
        RECT 52.900 114.175 53.220 114.235 ;
        RECT 54.295 114.190 54.585 114.235 ;
        RECT 57.040 114.175 57.360 114.435 ;
        RECT 90.620 114.375 90.940 114.435 ;
        RECT 92.015 114.375 92.305 114.420 ;
        RECT 90.620 114.235 92.305 114.375 ;
        RECT 90.620 114.175 90.940 114.235 ;
        RECT 92.015 114.190 92.305 114.235 ;
        RECT 93.840 114.175 94.160 114.435 ;
        RECT 11.430 113.555 118.610 114.035 ;
        RECT 16.115 113.355 16.405 113.400 ;
        RECT 17.480 113.355 17.800 113.415 ;
        RECT 16.115 113.215 17.800 113.355 ;
        RECT 16.115 113.170 16.405 113.215 ;
        RECT 17.480 113.155 17.800 113.215 ;
        RECT 38.180 113.355 38.500 113.415 ;
        RECT 38.655 113.355 38.945 113.400 ;
        RECT 38.180 113.215 38.945 113.355 ;
        RECT 38.180 113.155 38.500 113.215 ;
        RECT 38.655 113.170 38.945 113.215 ;
        RECT 53.820 113.355 54.140 113.415 ;
        RECT 64.400 113.355 64.720 113.415 ;
        RECT 53.820 113.215 64.720 113.355 ;
        RECT 53.820 113.155 54.140 113.215 ;
        RECT 64.400 113.155 64.720 113.215 ;
        RECT 79.580 113.355 79.900 113.415 ;
        RECT 86.480 113.355 86.800 113.415 ;
        RECT 89.255 113.355 89.545 113.400 ;
        RECT 79.580 113.215 80.270 113.355 ;
        RECT 79.580 113.155 79.900 113.215 ;
        RECT 21.275 113.015 21.565 113.060 ;
        RECT 24.395 113.015 24.685 113.060 ;
        RECT 26.285 113.015 26.575 113.060 ;
        RECT 31.280 113.015 31.600 113.075 ;
        RECT 21.275 112.875 26.575 113.015 ;
        RECT 21.275 112.830 21.565 112.875 ;
        RECT 24.395 112.830 24.685 112.875 ;
        RECT 26.285 112.830 26.575 112.875 ;
        RECT 26.770 112.875 31.600 113.015 ;
        RECT 17.035 112.675 17.325 112.720 ;
        RECT 23.000 112.675 23.320 112.735 ;
        RECT 17.035 112.535 23.320 112.675 ;
        RECT 17.035 112.490 17.325 112.535 ;
        RECT 23.000 112.475 23.320 112.535 ;
        RECT 25.775 112.675 26.065 112.720 ;
        RECT 26.770 112.675 26.910 112.875 ;
        RECT 31.280 112.815 31.600 112.875 ;
        RECT 31.855 113.015 32.145 113.060 ;
        RECT 34.975 113.015 35.265 113.060 ;
        RECT 36.865 113.015 37.155 113.060 ;
        RECT 39.100 113.015 39.420 113.075 ;
        RECT 31.855 112.875 37.155 113.015 ;
        RECT 31.855 112.830 32.145 112.875 ;
        RECT 34.975 112.830 35.265 112.875 ;
        RECT 36.865 112.830 37.155 112.875 ;
        RECT 37.810 112.875 39.420 113.015 ;
        RECT 25.775 112.535 26.910 112.675 ;
        RECT 27.140 112.675 27.460 112.735 ;
        RECT 37.810 112.720 37.950 112.875 ;
        RECT 39.100 112.815 39.420 112.875 ;
        RECT 47.955 113.015 48.245 113.060 ;
        RECT 51.075 113.015 51.365 113.060 ;
        RECT 52.965 113.015 53.255 113.060 ;
        RECT 47.955 112.875 53.255 113.015 ;
        RECT 47.955 112.830 48.245 112.875 ;
        RECT 51.075 112.830 51.365 112.875 ;
        RECT 52.965 112.830 53.255 112.875 ;
        RECT 58.535 113.015 58.825 113.060 ;
        RECT 61.655 113.015 61.945 113.060 ;
        RECT 63.545 113.015 63.835 113.060 ;
        RECT 58.535 112.875 63.835 113.015 ;
        RECT 58.535 112.830 58.825 112.875 ;
        RECT 61.655 112.830 61.945 112.875 ;
        RECT 63.545 112.830 63.835 112.875 ;
        RECT 71.875 113.015 72.165 113.060 ;
        RECT 74.995 113.015 75.285 113.060 ;
        RECT 76.885 113.015 77.175 113.060 ;
        RECT 71.875 112.875 77.175 113.015 ;
        RECT 71.875 112.830 72.165 112.875 ;
        RECT 74.995 112.830 75.285 112.875 ;
        RECT 76.885 112.830 77.175 112.875 ;
        RECT 37.735 112.675 38.025 112.720 ;
        RECT 27.140 112.535 38.025 112.675 ;
        RECT 25.775 112.490 26.065 112.535 ;
        RECT 27.140 112.475 27.460 112.535 ;
        RECT 37.735 112.490 38.025 112.535 ;
        RECT 43.715 112.675 44.005 112.720 ;
        RECT 50.140 112.675 50.460 112.735 ;
        RECT 43.715 112.535 50.460 112.675 ;
        RECT 43.715 112.490 44.005 112.535 ;
        RECT 50.140 112.475 50.460 112.535 ;
        RECT 53.820 112.475 54.140 112.735 ;
        RECT 57.040 112.675 57.360 112.735 ;
        RECT 63.035 112.675 63.325 112.720 ;
        RECT 57.040 112.535 63.325 112.675 ;
        RECT 57.040 112.475 57.360 112.535 ;
        RECT 63.035 112.490 63.325 112.535 ;
        RECT 64.400 112.475 64.720 112.735 ;
        RECT 67.635 112.675 67.925 112.720 ;
        RECT 73.140 112.675 73.460 112.735 ;
        RECT 67.635 112.535 73.460 112.675 ;
        RECT 67.635 112.490 67.925 112.535 ;
        RECT 73.140 112.475 73.460 112.535 ;
        RECT 76.360 112.475 76.680 112.735 ;
        RECT 78.215 112.675 78.505 112.720 ;
        RECT 79.580 112.675 79.900 112.735 ;
        RECT 78.215 112.535 79.900 112.675 ;
        RECT 80.130 112.675 80.270 113.215 ;
        RECT 86.480 113.215 89.545 113.355 ;
        RECT 86.480 113.155 86.800 113.215 ;
        RECT 89.255 113.170 89.545 113.215 ;
        RECT 115.000 113.155 115.320 113.415 ;
        RECT 82.455 113.015 82.745 113.060 ;
        RECT 85.575 113.015 85.865 113.060 ;
        RECT 87.465 113.015 87.755 113.060 ;
        RECT 82.455 112.875 87.755 113.015 ;
        RECT 82.455 112.830 82.745 112.875 ;
        RECT 85.575 112.830 85.865 112.875 ;
        RECT 87.465 112.830 87.755 112.875 ;
        RECT 97.175 113.015 97.465 113.060 ;
        RECT 100.295 113.015 100.585 113.060 ;
        RECT 102.185 113.015 102.475 113.060 ;
        RECT 97.175 112.875 102.475 113.015 ;
        RECT 97.175 112.830 97.465 112.875 ;
        RECT 100.295 112.830 100.585 112.875 ;
        RECT 102.185 112.830 102.475 112.875 ;
        RECT 107.755 113.015 108.045 113.060 ;
        RECT 110.875 113.015 111.165 113.060 ;
        RECT 112.765 113.015 113.055 113.060 ;
        RECT 107.755 112.875 113.055 113.015 ;
        RECT 107.755 112.830 108.045 112.875 ;
        RECT 110.875 112.830 111.165 112.875 ;
        RECT 112.765 112.830 113.055 112.875 ;
        RECT 86.955 112.675 87.245 112.720 ;
        RECT 80.130 112.535 87.245 112.675 ;
        RECT 78.215 112.490 78.505 112.535 ;
        RECT 79.580 112.475 79.900 112.535 ;
        RECT 86.955 112.490 87.245 112.535 ;
        RECT 98.900 112.675 99.220 112.735 ;
        RECT 101.675 112.675 101.965 112.720 ;
        RECT 98.900 112.535 101.965 112.675 ;
        RECT 98.900 112.475 99.220 112.535 ;
        RECT 101.675 112.490 101.965 112.535 ;
        RECT 103.040 112.475 103.360 112.735 ;
        RECT 103.515 112.675 103.805 112.720 ;
        RECT 106.260 112.675 106.580 112.735 ;
        RECT 103.515 112.535 106.580 112.675 ;
        RECT 103.515 112.490 103.805 112.535 ;
        RECT 106.260 112.475 106.580 112.535 ;
        RECT 112.240 112.475 112.560 112.735 ;
        RECT 113.635 112.675 113.925 112.720 ;
        RECT 115.460 112.675 115.780 112.735 ;
        RECT 113.635 112.535 115.780 112.675 ;
        RECT 113.635 112.490 113.925 112.535 ;
        RECT 115.460 112.475 115.780 112.535 ;
        RECT 14.735 112.335 15.025 112.380 ;
        RECT 15.655 112.335 15.945 112.380 ;
        RECT 14.735 112.195 15.945 112.335 ;
        RECT 14.735 112.150 15.025 112.195 ;
        RECT 15.655 112.150 15.945 112.195 ;
        RECT 14.260 111.455 14.580 111.715 ;
        RECT 15.730 111.655 15.870 112.150 ;
        RECT 20.195 112.040 20.485 112.355 ;
        RECT 21.275 112.335 21.565 112.380 ;
        RECT 24.855 112.335 25.145 112.380 ;
        RECT 26.690 112.335 26.980 112.380 ;
        RECT 21.275 112.195 26.980 112.335 ;
        RECT 21.275 112.150 21.565 112.195 ;
        RECT 24.855 112.150 25.145 112.195 ;
        RECT 26.690 112.150 26.980 112.195 ;
        RECT 19.895 111.995 20.485 112.040 ;
        RECT 23.135 111.995 23.785 112.040 ;
        RECT 25.300 111.995 25.620 112.055 ;
        RECT 19.895 111.855 25.620 111.995 ;
        RECT 19.895 111.810 20.185 111.855 ;
        RECT 23.135 111.810 23.785 111.855 ;
        RECT 25.300 111.795 25.620 111.855 ;
        RECT 27.615 111.995 27.905 112.040 ;
        RECT 28.980 111.995 29.300 112.055 ;
        RECT 27.615 111.855 29.300 111.995 ;
        RECT 27.615 111.810 27.905 111.855 ;
        RECT 28.980 111.795 29.300 111.855 ;
        RECT 29.440 111.995 29.760 112.055 ;
        RECT 30.775 112.040 31.065 112.355 ;
        RECT 31.855 112.335 32.145 112.380 ;
        RECT 35.435 112.335 35.725 112.380 ;
        RECT 37.270 112.335 37.560 112.380 ;
        RECT 31.855 112.195 37.560 112.335 ;
        RECT 31.855 112.150 32.145 112.195 ;
        RECT 35.435 112.150 35.725 112.195 ;
        RECT 37.270 112.150 37.560 112.195 ;
        RECT 39.100 112.135 39.420 112.395 ;
        RECT 40.495 112.335 40.785 112.380 ;
        RECT 42.320 112.335 42.640 112.395 ;
        RECT 40.495 112.195 42.640 112.335 ;
        RECT 40.495 112.150 40.785 112.195 ;
        RECT 42.320 112.135 42.640 112.195 ;
        RECT 46.875 112.040 47.165 112.355 ;
        RECT 47.955 112.335 48.245 112.380 ;
        RECT 51.535 112.335 51.825 112.380 ;
        RECT 53.370 112.335 53.660 112.380 ;
        RECT 47.955 112.195 53.660 112.335 ;
        RECT 47.955 112.150 48.245 112.195 ;
        RECT 51.535 112.150 51.825 112.195 ;
        RECT 53.370 112.150 53.660 112.195 ;
        RECT 30.475 111.995 31.065 112.040 ;
        RECT 33.715 111.995 34.365 112.040 ;
        RECT 29.440 111.855 34.365 111.995 ;
        RECT 29.440 111.795 29.760 111.855 ;
        RECT 30.475 111.810 30.765 111.855 ;
        RECT 33.715 111.810 34.365 111.855 ;
        RECT 36.355 111.810 36.645 112.040 ;
        RECT 46.575 111.995 47.165 112.040 ;
        RECT 49.815 111.995 50.465 112.040 ;
        RECT 51.980 111.995 52.300 112.055 ;
        RECT 46.575 111.855 52.300 111.995 ;
        RECT 46.575 111.810 46.865 111.855 ;
        RECT 49.815 111.810 50.465 111.855 ;
        RECT 29.900 111.655 30.220 111.715 ;
        RECT 15.730 111.515 30.220 111.655 ;
        RECT 36.430 111.655 36.570 111.810 ;
        RECT 51.980 111.795 52.300 111.855 ;
        RECT 52.455 111.995 52.745 112.040 ;
        RECT 52.900 111.995 53.220 112.055 ;
        RECT 52.455 111.855 53.220 111.995 ;
        RECT 52.455 111.810 52.745 111.855 ;
        RECT 52.900 111.795 53.220 111.855 ;
        RECT 54.295 111.995 54.585 112.040 ;
        RECT 56.580 111.995 56.900 112.055 ;
        RECT 57.455 112.040 57.745 112.355 ;
        RECT 58.535 112.335 58.825 112.380 ;
        RECT 62.115 112.335 62.405 112.380 ;
        RECT 63.950 112.335 64.240 112.380 ;
        RECT 58.535 112.195 64.240 112.335 ;
        RECT 58.535 112.150 58.825 112.195 ;
        RECT 62.115 112.150 62.405 112.195 ;
        RECT 63.950 112.150 64.240 112.195 ;
        RECT 54.295 111.855 56.900 111.995 ;
        RECT 54.295 111.810 54.585 111.855 ;
        RECT 56.580 111.795 56.900 111.855 ;
        RECT 57.155 111.995 57.745 112.040 ;
        RECT 57.960 111.995 58.280 112.055 ;
        RECT 70.795 112.040 71.085 112.355 ;
        RECT 71.875 112.335 72.165 112.380 ;
        RECT 75.455 112.335 75.745 112.380 ;
        RECT 77.290 112.335 77.580 112.380 ;
        RECT 71.875 112.195 77.580 112.335 ;
        RECT 71.875 112.150 72.165 112.195 ;
        RECT 75.455 112.150 75.745 112.195 ;
        RECT 77.290 112.150 77.580 112.195 ;
        RECT 77.755 112.335 78.045 112.380 ;
        RECT 80.040 112.335 80.360 112.395 ;
        RECT 77.755 112.195 80.360 112.335 ;
        RECT 77.755 112.150 78.045 112.195 ;
        RECT 80.040 112.135 80.360 112.195 ;
        RECT 60.395 111.995 61.045 112.040 ;
        RECT 57.155 111.855 61.045 111.995 ;
        RECT 57.155 111.810 57.445 111.855 ;
        RECT 57.960 111.795 58.280 111.855 ;
        RECT 60.395 111.810 61.045 111.855 ;
        RECT 70.495 111.995 71.085 112.040 ;
        RECT 72.680 111.995 73.000 112.055 ;
        RECT 73.735 111.995 74.385 112.040 ;
        RECT 70.495 111.855 74.385 111.995 ;
        RECT 70.495 111.810 70.785 111.855 ;
        RECT 72.680 111.795 73.000 111.855 ;
        RECT 73.735 111.810 74.385 111.855 ;
        RECT 78.660 111.995 78.980 112.055 ;
        RECT 81.375 112.040 81.665 112.355 ;
        RECT 82.455 112.335 82.745 112.380 ;
        RECT 86.035 112.335 86.325 112.380 ;
        RECT 87.870 112.335 88.160 112.380 ;
        RECT 82.455 112.195 88.160 112.335 ;
        RECT 82.455 112.150 82.745 112.195 ;
        RECT 86.035 112.150 86.325 112.195 ;
        RECT 87.870 112.150 88.160 112.195 ;
        RECT 88.335 112.150 88.625 112.380 ;
        RECT 89.700 112.335 90.020 112.395 ;
        RECT 91.095 112.335 91.385 112.380 ;
        RECT 93.380 112.335 93.700 112.395 ;
        RECT 89.700 112.195 93.700 112.335 ;
        RECT 81.075 111.995 81.665 112.040 ;
        RECT 84.315 111.995 84.965 112.040 ;
        RECT 78.660 111.855 84.965 111.995 ;
        RECT 78.660 111.795 78.980 111.855 ;
        RECT 81.075 111.810 81.365 111.855 ;
        RECT 84.315 111.810 84.965 111.855 ;
        RECT 85.560 111.995 85.880 112.055 ;
        RECT 88.410 111.995 88.550 112.150 ;
        RECT 89.700 112.135 90.020 112.195 ;
        RECT 91.095 112.150 91.385 112.195 ;
        RECT 93.380 112.135 93.700 112.195 ;
        RECT 93.840 112.335 94.160 112.395 ;
        RECT 96.095 112.335 96.385 112.355 ;
        RECT 93.840 112.195 96.385 112.335 ;
        RECT 93.840 112.135 94.160 112.195 ;
        RECT 85.560 111.855 88.550 111.995 ;
        RECT 92.935 111.995 93.225 112.040 ;
        RECT 95.220 111.995 95.540 112.055 ;
        RECT 96.095 112.040 96.385 112.195 ;
        RECT 97.175 112.335 97.465 112.380 ;
        RECT 100.755 112.335 101.045 112.380 ;
        RECT 102.590 112.335 102.880 112.380 ;
        RECT 97.175 112.195 102.880 112.335 ;
        RECT 97.175 112.150 97.465 112.195 ;
        RECT 100.755 112.150 101.045 112.195 ;
        RECT 102.590 112.150 102.880 112.195 ;
        RECT 92.935 111.855 95.540 111.995 ;
        RECT 85.560 111.795 85.880 111.855 ;
        RECT 92.935 111.810 93.225 111.855 ;
        RECT 95.220 111.795 95.540 111.855 ;
        RECT 95.795 111.995 96.385 112.040 ;
        RECT 99.035 111.995 99.685 112.040 ;
        RECT 95.795 111.855 99.685 111.995 ;
        RECT 95.795 111.810 96.085 111.855 ;
        RECT 99.035 111.810 99.685 111.855 ;
        RECT 103.960 111.995 104.280 112.055 ;
        RECT 106.675 112.040 106.965 112.355 ;
        RECT 107.755 112.335 108.045 112.380 ;
        RECT 111.335 112.335 111.625 112.380 ;
        RECT 113.170 112.335 113.460 112.380 ;
        RECT 107.755 112.195 113.460 112.335 ;
        RECT 107.755 112.150 108.045 112.195 ;
        RECT 111.335 112.150 111.625 112.195 ;
        RECT 113.170 112.150 113.460 112.195 ;
        RECT 114.080 112.135 114.400 112.395 ;
        RECT 106.375 111.995 106.965 112.040 ;
        RECT 109.615 111.995 110.265 112.040 ;
        RECT 103.960 111.855 110.265 111.995 ;
        RECT 103.960 111.795 104.280 111.855 ;
        RECT 106.375 111.810 106.665 111.855 ;
        RECT 109.615 111.810 110.265 111.855 ;
        RECT 39.575 111.655 39.865 111.700 ;
        RECT 36.430 111.515 39.865 111.655 ;
        RECT 29.900 111.455 30.220 111.515 ;
        RECT 39.575 111.470 39.865 111.515 ;
        RECT 88.320 111.655 88.640 111.715 ;
        RECT 90.635 111.655 90.925 111.700 ;
        RECT 88.320 111.515 90.925 111.655 ;
        RECT 88.320 111.455 88.640 111.515 ;
        RECT 90.635 111.470 90.925 111.515 ;
        RECT 10.650 110.835 118.610 111.315 ;
        RECT 23.460 110.635 23.780 110.695 ;
        RECT 25.300 110.635 25.620 110.695 ;
        RECT 26.695 110.635 26.985 110.680 ;
        RECT 23.460 110.495 24.610 110.635 ;
        RECT 23.460 110.435 23.780 110.495 ;
        RECT 14.260 110.295 14.580 110.355 ;
        RECT 24.470 110.340 24.610 110.495 ;
        RECT 25.300 110.495 26.985 110.635 ;
        RECT 25.300 110.435 25.620 110.495 ;
        RECT 26.695 110.450 26.985 110.495 ;
        RECT 47.855 110.635 48.145 110.680 ;
        RECT 48.300 110.635 48.620 110.695 ;
        RECT 47.855 110.495 48.620 110.635 ;
        RECT 47.855 110.450 48.145 110.495 ;
        RECT 48.300 110.435 48.620 110.495 ;
        RECT 51.980 110.435 52.300 110.695 ;
        RECT 57.960 110.635 58.280 110.695 ;
        RECT 58.895 110.635 59.185 110.680 ;
        RECT 57.960 110.495 59.185 110.635 ;
        RECT 57.960 110.435 58.280 110.495 ;
        RECT 58.895 110.450 59.185 110.495 ;
        RECT 78.660 110.435 78.980 110.695 ;
        RECT 89.700 110.635 90.020 110.695 ;
        RECT 84.270 110.495 90.020 110.635 ;
        RECT 18.515 110.295 18.805 110.340 ;
        RECT 21.755 110.295 22.405 110.340 ;
        RECT 14.260 110.155 22.405 110.295 ;
        RECT 14.260 110.095 14.580 110.155 ;
        RECT 18.515 110.110 19.105 110.155 ;
        RECT 21.755 110.110 22.405 110.155 ;
        RECT 24.395 110.110 24.685 110.340 ;
        RECT 18.815 109.795 19.105 110.110 ;
        RECT 19.895 109.955 20.185 110.000 ;
        RECT 23.475 109.955 23.765 110.000 ;
        RECT 25.310 109.955 25.600 110.000 ;
        RECT 19.895 109.815 25.600 109.955 ;
        RECT 19.895 109.770 20.185 109.815 ;
        RECT 23.475 109.770 23.765 109.815 ;
        RECT 25.310 109.770 25.600 109.815 ;
        RECT 25.775 109.955 26.065 110.000 ;
        RECT 26.680 109.955 27.000 110.015 ;
        RECT 25.775 109.815 27.000 109.955 ;
        RECT 25.775 109.770 26.065 109.815 ;
        RECT 26.680 109.755 27.000 109.815 ;
        RECT 27.155 109.955 27.445 110.000 ;
        RECT 29.900 109.955 30.220 110.015 ;
        RECT 39.100 109.955 39.420 110.015 ;
        RECT 48.315 109.955 48.605 110.000 ;
        RECT 52.455 109.955 52.745 110.000 ;
        RECT 59.340 109.955 59.660 110.015 ;
        RECT 27.155 109.815 59.660 109.955 ;
        RECT 27.155 109.770 27.445 109.815 ;
        RECT 29.900 109.755 30.220 109.815 ;
        RECT 39.100 109.755 39.420 109.815 ;
        RECT 48.315 109.770 48.605 109.815 ;
        RECT 52.455 109.770 52.745 109.815 ;
        RECT 59.340 109.755 59.660 109.815 ;
        RECT 74.060 109.955 74.380 110.015 ;
        RECT 78.215 109.955 78.505 110.000 ;
        RECT 84.270 109.955 84.410 110.495 ;
        RECT 89.700 110.435 90.020 110.495 ;
        RECT 110.400 110.635 110.720 110.695 ;
        RECT 110.875 110.635 111.165 110.680 ;
        RECT 110.400 110.495 111.165 110.635 ;
        RECT 110.400 110.435 110.720 110.495 ;
        RECT 110.875 110.450 111.165 110.495 ;
        RECT 88.320 110.340 88.640 110.355 ;
        RECT 84.755 110.295 85.045 110.340 ;
        RECT 87.995 110.295 88.645 110.340 ;
        RECT 84.755 110.155 88.645 110.295 ;
        RECT 84.755 110.110 85.345 110.155 ;
        RECT 87.995 110.110 88.645 110.155 ;
        RECT 74.060 109.815 84.410 109.955 ;
        RECT 74.060 109.755 74.380 109.815 ;
        RECT 78.215 109.770 78.505 109.815 ;
        RECT 85.055 109.795 85.345 110.110 ;
        RECT 88.320 110.095 88.640 110.110 ;
        RECT 90.620 110.095 90.940 110.355 ;
        RECT 86.135 109.955 86.425 110.000 ;
        RECT 89.715 109.955 90.005 110.000 ;
        RECT 91.550 109.955 91.840 110.000 ;
        RECT 86.135 109.815 91.840 109.955 ;
        RECT 86.135 109.770 86.425 109.815 ;
        RECT 89.715 109.770 90.005 109.815 ;
        RECT 91.550 109.770 91.840 109.815 ;
        RECT 108.560 109.955 108.880 110.015 ;
        RECT 110.415 109.955 110.705 110.000 ;
        RECT 108.560 109.815 110.705 109.955 ;
        RECT 108.560 109.755 108.880 109.815 ;
        RECT 110.415 109.770 110.705 109.815 ;
        RECT 12.420 109.615 12.740 109.675 ;
        RECT 15.655 109.615 15.945 109.660 ;
        RECT 12.420 109.475 15.945 109.615 ;
        RECT 12.420 109.415 12.740 109.475 ;
        RECT 15.655 109.430 15.945 109.475 ;
        RECT 81.895 109.615 82.185 109.660 ;
        RECT 85.560 109.615 85.880 109.675 ;
        RECT 92.015 109.615 92.305 109.660 ;
        RECT 81.895 109.475 85.330 109.615 ;
        RECT 81.895 109.430 82.185 109.475 ;
        RECT 19.895 109.275 20.185 109.320 ;
        RECT 23.015 109.275 23.305 109.320 ;
        RECT 24.905 109.275 25.195 109.320 ;
        RECT 19.895 109.135 25.195 109.275 ;
        RECT 19.895 109.090 20.185 109.135 ;
        RECT 23.015 109.090 23.305 109.135 ;
        RECT 24.905 109.090 25.195 109.135 ;
        RECT 85.190 108.935 85.330 109.475 ;
        RECT 85.560 109.475 92.305 109.615 ;
        RECT 85.560 109.415 85.880 109.475 ;
        RECT 92.015 109.430 92.305 109.475 ;
        RECT 86.135 109.275 86.425 109.320 ;
        RECT 89.255 109.275 89.545 109.320 ;
        RECT 91.145 109.275 91.435 109.320 ;
        RECT 86.135 109.135 91.435 109.275 ;
        RECT 86.135 109.090 86.425 109.135 ;
        RECT 89.255 109.090 89.545 109.135 ;
        RECT 91.145 109.090 91.435 109.135 ;
        RECT 89.700 108.935 90.020 108.995 ;
        RECT 85.190 108.795 90.020 108.935 ;
        RECT 89.700 108.735 90.020 108.795 ;
        RECT 11.430 108.115 118.610 108.595 ;
        RECT 135.660 106.690 136.800 133.400 ;
        RECT 133.100 106.600 136.850 106.690 ;
        RECT 129.700 105.630 136.850 106.600 ;
        RECT 133.100 105.500 136.850 105.630 ;
        RECT 133.330 76.630 136.060 77.830 ;
        RECT 137.920 77.810 143.450 77.960 ;
        RECT 21.115 74.380 23.065 74.390 ;
        RECT 19.415 73.240 23.065 74.380 ;
        RECT 19.415 73.230 21.125 73.240 ;
        RECT 28.135 73.230 30.305 74.410 ;
        RECT 32.315 74.390 34.265 74.400 ;
        RECT 30.615 73.250 34.265 74.390 ;
        RECT 30.615 73.240 32.325 73.250 ;
        RECT 39.425 73.200 41.595 74.380 ;
        RECT 43.535 74.360 45.485 74.370 ;
        RECT 41.835 73.220 45.485 74.360 ;
        RECT 54.785 74.340 56.735 74.350 ;
        RECT 41.835 73.210 43.545 73.220 ;
        RECT 3.910 73.080 6.100 73.190 ;
        RECT 50.005 73.140 52.175 74.320 ;
        RECT 53.085 73.200 56.735 74.340 ;
        RECT 53.085 73.190 54.795 73.200 ;
        RECT 61.425 73.170 63.595 74.350 ;
        RECT 66.005 74.330 67.955 74.340 ;
        RECT 64.305 73.190 67.955 74.330 ;
        RECT 64.305 73.180 66.015 73.190 ;
        RECT 72.535 73.180 74.705 74.360 ;
        RECT 77.245 74.320 79.195 74.330 ;
        RECT 75.545 73.180 79.195 74.320 ;
        RECT 75.545 73.170 77.255 73.180 ;
        RECT 83.805 73.170 85.975 74.350 ;
        RECT 88.495 74.330 90.445 74.340 ;
        RECT 86.795 73.190 90.445 74.330 ;
        RECT 99.775 74.320 101.725 74.330 ;
        RECT 86.795 73.180 88.505 73.190 ;
        RECT 94.995 73.110 97.165 74.290 ;
        RECT 98.075 73.180 101.725 74.320 ;
        RECT 98.075 73.170 99.785 73.180 ;
        RECT 106.405 73.160 108.575 74.340 ;
        RECT 111.045 74.320 112.995 74.330 ;
        RECT 109.345 73.180 112.995 74.320 ;
        RECT 109.345 73.170 111.055 73.180 ;
        RECT 117.605 73.160 119.775 74.340 ;
        RECT 122.295 74.320 124.245 74.330 ;
        RECT 120.595 73.180 124.245 74.320 ;
        RECT 129.455 73.240 131.625 74.420 ;
        RECT 120.595 73.170 122.305 73.180 ;
        RECT 3.910 72.820 12.240 73.080 ;
        RECT 29.635 72.840 43.235 72.850 ;
        RECT 18.435 72.820 43.235 72.840 ;
        RECT 3.910 72.800 54.455 72.820 ;
        RECT 3.910 72.790 65.705 72.800 ;
        RECT 133.960 72.790 135.640 76.630 ;
        RECT 137.190 76.610 143.450 77.810 ;
        RECT 137.920 75.460 143.450 76.610 ;
        RECT 3.910 72.780 76.925 72.790 ;
        RECT 85.815 72.780 99.415 72.790 ;
        RECT 132.085 72.780 140.600 72.790 ;
        RECT 3.910 71.700 140.600 72.780 ;
        RECT 3.910 71.690 32.035 71.700 ;
        RECT 3.910 71.670 19.135 71.690 ;
        RECT 40.855 71.670 140.600 71.700 ;
        RECT 3.910 71.500 12.240 71.670 ;
        RECT 52.105 71.650 140.600 71.670 ;
        RECT 63.325 71.640 140.600 71.650 ;
        RECT 74.565 71.630 88.165 71.640 ;
        RECT 97.095 71.630 133.215 71.640 ;
        RECT 3.910 71.370 6.100 71.500 ;
        RECT 10.800 71.180 11.950 71.500 ;
        RECT 10.800 69.480 11.915 71.180 ;
        RECT 29.635 71.170 43.285 71.180 ;
        RECT 15.510 71.155 17.040 71.160 ;
        RECT 18.435 71.155 43.285 71.170 ;
        RECT 12.285 71.150 43.285 71.155 ;
        RECT 12.285 71.130 54.505 71.150 ;
        RECT 141.810 71.140 143.230 75.460 ;
        RECT 12.285 71.120 65.755 71.130 ;
        RECT 12.285 71.110 76.975 71.120 ;
        RECT 85.815 71.110 99.465 71.120 ;
        RECT 140.220 71.110 143.240 71.140 ;
        RECT 12.285 70.030 143.240 71.110 ;
        RECT 12.285 70.020 32.085 70.030 ;
        RECT 12.285 70.005 19.375 70.020 ;
        RECT 10.800 13.800 11.950 69.480 ;
        RECT 12.320 15.450 13.470 70.005 ;
        RECT 15.510 68.660 17.040 70.005 ;
        RECT 40.855 70.000 143.240 70.030 ;
        RECT 52.105 69.980 143.240 70.000 ;
        RECT 63.325 69.970 143.240 69.980 ;
        RECT 74.565 69.960 88.215 69.970 ;
        RECT 97.095 69.960 143.240 69.970 ;
        RECT 140.220 69.910 143.240 69.960 ;
        RECT 29.645 69.670 43.315 69.680 ;
        RECT 18.445 69.650 43.315 69.670 ;
        RECT 18.445 69.630 54.535 69.650 ;
        RECT 18.445 69.620 65.785 69.630 ;
        RECT 139.590 69.620 150.610 69.640 ;
        RECT 18.445 69.610 77.005 69.620 ;
        RECT 85.825 69.610 99.495 69.620 ;
        RECT 132.155 69.610 150.610 69.620 ;
        RECT 18.445 69.570 150.610 69.610 ;
        RECT 18.445 68.530 150.740 69.570 ;
        RECT 18.445 68.520 32.115 68.530 ;
        RECT 40.865 68.500 150.740 68.530 ;
        RECT 52.115 68.490 143.320 68.500 ;
        RECT 52.115 68.480 140.670 68.490 ;
        RECT 63.335 68.470 140.670 68.480 ;
        RECT 74.575 68.460 88.245 68.470 ;
        RECT 97.105 68.460 133.295 68.470 ;
        RECT 141.080 68.450 142.300 68.490 ;
        RECT 149.360 68.470 150.740 68.500 ;
        RECT 29.655 68.100 43.325 68.110 ;
        RECT 13.950 68.080 43.325 68.100 ;
        RECT 13.950 68.060 54.545 68.080 ;
        RECT 13.950 68.050 65.795 68.060 ;
        RECT 13.950 68.040 77.015 68.050 ;
        RECT 85.835 68.040 99.505 68.050 ;
        RECT 139.530 68.040 143.320 68.060 ;
        RECT 13.950 66.960 152.870 68.040 ;
        RECT 13.950 66.950 32.125 66.960 ;
        RECT 13.950 18.530 15.100 66.950 ;
        RECT 40.875 66.930 152.870 66.960 ;
        RECT 52.125 66.910 152.870 66.930 ;
        RECT 63.345 66.900 152.870 66.910 ;
        RECT 74.585 66.890 88.255 66.900 ;
        RECT 97.115 66.890 143.320 66.900 ;
        RECT 141.030 66.770 142.490 66.890 ;
        RECT 21.405 65.510 26.555 65.790 ;
        RECT 27.815 65.490 28.965 65.800 ;
        RECT 32.605 65.520 37.755 65.800 ;
        RECT 39.015 65.500 40.165 65.810 ;
        RECT 43.825 65.490 48.975 65.770 ;
        RECT 50.235 65.470 51.385 65.780 ;
        RECT 149.460 65.760 150.600 65.780 ;
        RECT 55.075 65.470 60.225 65.750 ;
        RECT 61.485 65.450 62.635 65.760 ;
        RECT 66.295 65.460 71.445 65.740 ;
        RECT 72.705 65.440 73.855 65.750 ;
        RECT 77.535 65.450 82.685 65.730 ;
        RECT 83.945 65.430 85.095 65.740 ;
        RECT 88.785 65.460 93.935 65.740 ;
        RECT 95.195 65.440 96.345 65.750 ;
        RECT 100.065 65.450 105.215 65.730 ;
        RECT 106.475 65.430 107.625 65.740 ;
        RECT 111.335 65.450 116.485 65.730 ;
        RECT 117.745 65.430 118.895 65.740 ;
        RECT 122.585 65.450 127.735 65.730 ;
        RECT 128.995 65.430 130.145 65.740 ;
        RECT 133.315 65.430 138.455 65.690 ;
        RECT 21.205 65.140 21.435 65.320 ;
        RECT 26.495 65.190 26.725 65.320 ;
        RECT 21.125 55.220 21.485 65.140 ;
        RECT 26.435 55.240 26.805 65.190 ;
        RECT 27.635 65.150 27.865 65.320 ;
        RECT 27.565 55.200 27.935 65.150 ;
        RECT 28.925 65.140 29.155 65.320 ;
        RECT 32.405 65.150 32.635 65.330 ;
        RECT 37.695 65.200 37.925 65.330 ;
        RECT 28.835 55.250 29.255 65.140 ;
        RECT 32.325 55.230 32.685 65.150 ;
        RECT 37.635 55.250 38.005 65.200 ;
        RECT 38.835 65.160 39.065 65.330 ;
        RECT 38.765 55.210 39.135 65.160 ;
        RECT 40.125 65.150 40.355 65.330 ;
        RECT 40.035 55.260 40.455 65.150 ;
        RECT 43.625 65.120 43.855 65.300 ;
        RECT 48.915 65.170 49.145 65.300 ;
        RECT 43.545 55.200 43.905 65.120 ;
        RECT 48.855 55.220 49.225 65.170 ;
        RECT 50.055 65.130 50.285 65.300 ;
        RECT 49.985 55.180 50.355 65.130 ;
        RECT 51.345 65.120 51.575 65.300 ;
        RECT 51.255 55.230 51.675 65.120 ;
        RECT 54.875 65.100 55.105 65.280 ;
        RECT 60.165 65.150 60.395 65.280 ;
        RECT 54.795 55.180 55.155 65.100 ;
        RECT 60.105 55.200 60.475 65.150 ;
        RECT 61.305 65.110 61.535 65.280 ;
        RECT 61.235 55.160 61.605 65.110 ;
        RECT 62.595 65.100 62.825 65.280 ;
        RECT 62.505 55.210 62.925 65.100 ;
        RECT 66.095 65.090 66.325 65.270 ;
        RECT 71.385 65.140 71.615 65.270 ;
        RECT 66.015 55.170 66.375 65.090 ;
        RECT 71.325 55.190 71.695 65.140 ;
        RECT 72.525 65.100 72.755 65.270 ;
        RECT 72.455 55.150 72.825 65.100 ;
        RECT 73.815 65.090 74.045 65.270 ;
        RECT 73.725 55.200 74.145 65.090 ;
        RECT 77.335 65.080 77.565 65.260 ;
        RECT 82.625 65.130 82.855 65.260 ;
        RECT 77.255 55.160 77.615 65.080 ;
        RECT 82.565 55.180 82.935 65.130 ;
        RECT 83.765 65.090 83.995 65.260 ;
        RECT 83.695 55.140 84.065 65.090 ;
        RECT 85.055 65.080 85.285 65.260 ;
        RECT 88.585 65.090 88.815 65.270 ;
        RECT 93.875 65.140 94.105 65.270 ;
        RECT 84.965 55.190 85.385 65.080 ;
        RECT 88.505 55.170 88.865 65.090 ;
        RECT 93.815 55.190 94.185 65.140 ;
        RECT 95.015 65.100 95.245 65.270 ;
        RECT 94.945 55.150 95.315 65.100 ;
        RECT 96.305 65.090 96.535 65.270 ;
        RECT 96.215 55.200 96.635 65.090 ;
        RECT 99.865 65.080 100.095 65.260 ;
        RECT 105.155 65.130 105.385 65.260 ;
        RECT 99.785 55.160 100.145 65.080 ;
        RECT 105.095 55.180 105.465 65.130 ;
        RECT 106.295 65.090 106.525 65.260 ;
        RECT 106.225 55.140 106.595 65.090 ;
        RECT 107.585 65.080 107.815 65.260 ;
        RECT 111.135 65.080 111.365 65.260 ;
        RECT 116.425 65.130 116.655 65.260 ;
        RECT 107.495 55.190 107.915 65.080 ;
        RECT 111.055 55.160 111.415 65.080 ;
        RECT 116.365 55.180 116.735 65.130 ;
        RECT 117.565 65.090 117.795 65.260 ;
        RECT 117.495 55.140 117.865 65.090 ;
        RECT 118.855 65.080 119.085 65.260 ;
        RECT 122.385 65.080 122.615 65.260 ;
        RECT 127.675 65.130 127.905 65.260 ;
        RECT 118.765 55.190 119.185 65.080 ;
        RECT 122.305 55.160 122.665 65.080 ;
        RECT 127.615 55.180 127.985 65.130 ;
        RECT 128.815 65.090 129.045 65.260 ;
        RECT 128.745 55.140 129.115 65.090 ;
        RECT 130.105 65.080 130.335 65.260 ;
        RECT 133.135 65.130 133.365 65.230 ;
        RECT 130.015 55.190 130.435 65.080 ;
        RECT 133.005 55.240 133.405 65.130 ;
        RECT 138.425 65.100 138.655 65.230 ;
        RECT 133.135 55.230 133.365 55.240 ;
        RECT 138.345 55.130 138.725 65.100 ;
        RECT 149.340 64.660 150.720 65.760 ;
        RECT 20.815 54.230 25.555 54.530 ;
        RECT 32.015 54.240 36.755 54.540 ;
        RECT 43.235 54.210 47.975 54.510 ;
        RECT 54.485 54.190 59.225 54.490 ;
        RECT 65.705 54.180 70.445 54.480 ;
        RECT 76.945 54.170 81.685 54.470 ;
        RECT 88.195 54.180 92.935 54.480 ;
        RECT 99.475 54.170 104.215 54.470 ;
        RECT 110.745 54.170 115.485 54.470 ;
        RECT 121.995 54.170 126.735 54.470 ;
        RECT 21.655 52.320 22.115 52.550 ;
        RECT 25.625 52.280 26.255 52.560 ;
        RECT 25.735 52.240 26.195 52.280 ;
        RECT 27.665 52.240 28.125 52.470 ;
        RECT 32.855 52.330 33.315 52.560 ;
        RECT 36.825 52.290 37.455 52.570 ;
        RECT 36.935 52.250 37.395 52.290 ;
        RECT 38.865 52.250 39.325 52.480 ;
        RECT 44.075 52.300 44.535 52.530 ;
        RECT 48.045 52.260 48.675 52.540 ;
        RECT 48.155 52.220 48.615 52.260 ;
        RECT 50.085 52.220 50.545 52.450 ;
        RECT 55.325 52.280 55.785 52.510 ;
        RECT 59.295 52.240 59.925 52.520 ;
        RECT 59.405 52.200 59.865 52.240 ;
        RECT 61.335 52.200 61.795 52.430 ;
        RECT 66.545 52.270 67.005 52.500 ;
        RECT 70.515 52.230 71.145 52.510 ;
        RECT 70.625 52.190 71.085 52.230 ;
        RECT 72.555 52.190 73.015 52.420 ;
        RECT 77.785 52.260 78.245 52.490 ;
        RECT 81.755 52.220 82.385 52.500 ;
        RECT 81.865 52.180 82.325 52.220 ;
        RECT 83.795 52.180 84.255 52.410 ;
        RECT 89.035 52.270 89.495 52.500 ;
        RECT 93.005 52.230 93.635 52.510 ;
        RECT 93.115 52.190 93.575 52.230 ;
        RECT 95.045 52.190 95.505 52.420 ;
        RECT 100.315 52.260 100.775 52.490 ;
        RECT 104.285 52.220 104.915 52.500 ;
        RECT 104.395 52.180 104.855 52.220 ;
        RECT 106.325 52.180 106.785 52.410 ;
        RECT 111.585 52.260 112.045 52.490 ;
        RECT 115.555 52.220 116.185 52.500 ;
        RECT 115.665 52.180 116.125 52.220 ;
        RECT 117.595 52.180 118.055 52.410 ;
        RECT 122.835 52.260 123.295 52.490 ;
        RECT 126.805 52.220 127.435 52.500 ;
        RECT 126.915 52.180 127.375 52.220 ;
        RECT 128.845 52.180 129.305 52.410 ;
        RECT 21.375 52.010 21.605 52.115 ;
        RECT 21.245 50.290 21.615 52.010 ;
        RECT 22.165 51.890 22.395 52.115 ;
        RECT 25.455 51.980 25.685 52.035 ;
        RECT 21.375 50.115 21.605 50.290 ;
        RECT 22.155 50.210 22.525 51.890 ;
        RECT 22.165 50.115 22.395 50.210 ;
        RECT 21.525 49.670 22.245 49.930 ;
        RECT 19.295 46.650 20.065 47.720 ;
        RECT 21.385 47.490 22.105 47.750 ;
        RECT 21.225 47.200 21.455 47.340 ;
        RECT 21.085 46.430 21.475 47.200 ;
        RECT 22.015 47.190 22.245 47.340 ;
        RECT 22.005 46.450 22.375 47.190 ;
        RECT 25.305 47.010 25.735 51.980 ;
        RECT 26.245 51.970 26.475 52.035 ;
        RECT 27.385 51.970 27.615 52.035 ;
        RECT 26.185 46.970 26.585 51.970 ;
        RECT 27.265 46.970 27.665 51.970 ;
        RECT 28.175 51.940 28.405 52.035 ;
        RECT 32.575 52.020 32.805 52.125 ;
        RECT 28.115 46.970 28.545 51.940 ;
        RECT 32.445 50.300 32.815 52.020 ;
        RECT 33.365 51.900 33.595 52.125 ;
        RECT 36.655 51.990 36.885 52.045 ;
        RECT 32.575 50.125 32.805 50.300 ;
        RECT 33.355 50.220 33.725 51.900 ;
        RECT 33.365 50.125 33.595 50.220 ;
        RECT 32.725 49.680 33.445 49.940 ;
        RECT 25.735 46.600 26.195 46.830 ;
        RECT 27.665 46.710 28.125 46.830 ;
        RECT 27.515 46.600 28.125 46.710 ;
        RECT 30.495 46.660 31.265 47.730 ;
        RECT 32.585 47.500 33.305 47.760 ;
        RECT 32.425 47.210 32.655 47.350 ;
        RECT 21.225 46.340 21.455 46.430 ;
        RECT 22.015 46.340 22.245 46.450 ;
        RECT 27.515 46.430 28.095 46.600 ;
        RECT 32.285 46.440 32.675 47.210 ;
        RECT 33.215 47.200 33.445 47.350 ;
        RECT 33.205 46.460 33.575 47.200 ;
        RECT 36.505 47.020 36.935 51.990 ;
        RECT 37.445 51.980 37.675 52.045 ;
        RECT 38.585 51.980 38.815 52.045 ;
        RECT 37.385 46.980 37.785 51.980 ;
        RECT 38.465 46.980 38.865 51.980 ;
        RECT 39.375 51.950 39.605 52.045 ;
        RECT 43.795 51.990 44.025 52.095 ;
        RECT 39.315 46.980 39.745 51.950 ;
        RECT 43.665 50.270 44.035 51.990 ;
        RECT 44.585 51.870 44.815 52.095 ;
        RECT 47.875 51.960 48.105 52.015 ;
        RECT 43.795 50.095 44.025 50.270 ;
        RECT 44.575 50.190 44.945 51.870 ;
        RECT 44.585 50.095 44.815 50.190 ;
        RECT 43.945 49.650 44.665 49.910 ;
        RECT 36.935 46.610 37.395 46.840 ;
        RECT 38.865 46.720 39.325 46.840 ;
        RECT 38.715 46.610 39.325 46.720 ;
        RECT 41.715 46.630 42.485 47.700 ;
        RECT 43.805 47.470 44.525 47.730 ;
        RECT 43.645 47.180 43.875 47.320 ;
        RECT 32.425 46.350 32.655 46.440 ;
        RECT 33.215 46.350 33.445 46.460 ;
        RECT 38.715 46.440 39.295 46.610 ;
        RECT 43.505 46.410 43.895 47.180 ;
        RECT 44.435 47.170 44.665 47.320 ;
        RECT 44.425 46.430 44.795 47.170 ;
        RECT 47.725 46.990 48.155 51.960 ;
        RECT 48.665 51.950 48.895 52.015 ;
        RECT 49.805 51.950 50.035 52.015 ;
        RECT 48.605 46.950 49.005 51.950 ;
        RECT 49.685 46.950 50.085 51.950 ;
        RECT 50.595 51.920 50.825 52.015 ;
        RECT 55.045 51.970 55.275 52.075 ;
        RECT 50.535 46.950 50.965 51.920 ;
        RECT 54.915 50.250 55.285 51.970 ;
        RECT 55.835 51.850 56.065 52.075 ;
        RECT 59.125 51.940 59.355 51.995 ;
        RECT 55.045 50.075 55.275 50.250 ;
        RECT 55.825 50.170 56.195 51.850 ;
        RECT 55.835 50.075 56.065 50.170 ;
        RECT 55.195 49.630 55.915 49.890 ;
        RECT 48.155 46.580 48.615 46.810 ;
        RECT 50.085 46.690 50.545 46.810 ;
        RECT 49.935 46.580 50.545 46.690 ;
        RECT 52.965 46.610 53.735 47.680 ;
        RECT 55.055 47.450 55.775 47.710 ;
        RECT 54.895 47.160 55.125 47.300 ;
        RECT 43.645 46.320 43.875 46.410 ;
        RECT 44.435 46.320 44.665 46.430 ;
        RECT 49.935 46.410 50.515 46.580 ;
        RECT 54.755 46.390 55.145 47.160 ;
        RECT 55.685 47.150 55.915 47.300 ;
        RECT 55.675 46.410 56.045 47.150 ;
        RECT 58.975 46.970 59.405 51.940 ;
        RECT 59.915 51.930 60.145 51.995 ;
        RECT 61.055 51.930 61.285 51.995 ;
        RECT 59.855 46.930 60.255 51.930 ;
        RECT 60.935 46.930 61.335 51.930 ;
        RECT 61.845 51.900 62.075 51.995 ;
        RECT 66.265 51.960 66.495 52.065 ;
        RECT 61.785 46.930 62.215 51.900 ;
        RECT 66.135 50.240 66.505 51.960 ;
        RECT 67.055 51.840 67.285 52.065 ;
        RECT 70.345 51.930 70.575 51.985 ;
        RECT 66.265 50.065 66.495 50.240 ;
        RECT 67.045 50.160 67.415 51.840 ;
        RECT 67.055 50.065 67.285 50.160 ;
        RECT 66.415 49.620 67.135 49.880 ;
        RECT 59.405 46.560 59.865 46.790 ;
        RECT 61.335 46.670 61.795 46.790 ;
        RECT 61.185 46.560 61.795 46.670 ;
        RECT 64.185 46.600 64.955 47.670 ;
        RECT 66.275 47.440 66.995 47.700 ;
        RECT 66.115 47.150 66.345 47.290 ;
        RECT 54.895 46.300 55.125 46.390 ;
        RECT 55.685 46.300 55.915 46.410 ;
        RECT 61.185 46.390 61.765 46.560 ;
        RECT 65.975 46.380 66.365 47.150 ;
        RECT 66.905 47.140 67.135 47.290 ;
        RECT 66.895 46.400 67.265 47.140 ;
        RECT 70.195 46.960 70.625 51.930 ;
        RECT 71.135 51.920 71.365 51.985 ;
        RECT 72.275 51.920 72.505 51.985 ;
        RECT 71.075 46.920 71.475 51.920 ;
        RECT 72.155 46.920 72.555 51.920 ;
        RECT 73.065 51.890 73.295 51.985 ;
        RECT 77.505 51.950 77.735 52.055 ;
        RECT 73.005 46.920 73.435 51.890 ;
        RECT 77.375 50.230 77.745 51.950 ;
        RECT 78.295 51.830 78.525 52.055 ;
        RECT 81.585 51.920 81.815 51.975 ;
        RECT 77.505 50.055 77.735 50.230 ;
        RECT 78.285 50.150 78.655 51.830 ;
        RECT 78.295 50.055 78.525 50.150 ;
        RECT 77.655 49.610 78.375 49.870 ;
        RECT 70.625 46.550 71.085 46.780 ;
        RECT 72.555 46.660 73.015 46.780 ;
        RECT 72.405 46.550 73.015 46.660 ;
        RECT 75.425 46.590 76.195 47.660 ;
        RECT 77.515 47.430 78.235 47.690 ;
        RECT 77.355 47.140 77.585 47.280 ;
        RECT 66.115 46.290 66.345 46.380 ;
        RECT 66.905 46.290 67.135 46.400 ;
        RECT 72.405 46.380 72.985 46.550 ;
        RECT 77.215 46.370 77.605 47.140 ;
        RECT 78.145 47.130 78.375 47.280 ;
        RECT 78.135 46.390 78.505 47.130 ;
        RECT 81.435 46.950 81.865 51.920 ;
        RECT 82.375 51.910 82.605 51.975 ;
        RECT 83.515 51.910 83.745 51.975 ;
        RECT 82.315 46.910 82.715 51.910 ;
        RECT 83.395 46.910 83.795 51.910 ;
        RECT 84.305 51.880 84.535 51.975 ;
        RECT 88.755 51.960 88.985 52.065 ;
        RECT 84.245 46.910 84.675 51.880 ;
        RECT 88.625 50.240 88.995 51.960 ;
        RECT 89.545 51.840 89.775 52.065 ;
        RECT 92.835 51.930 93.065 51.985 ;
        RECT 88.755 50.065 88.985 50.240 ;
        RECT 89.535 50.160 89.905 51.840 ;
        RECT 89.545 50.065 89.775 50.160 ;
        RECT 88.905 49.620 89.625 49.880 ;
        RECT 81.865 46.540 82.325 46.770 ;
        RECT 83.795 46.650 84.255 46.770 ;
        RECT 83.645 46.540 84.255 46.650 ;
        RECT 86.675 46.600 87.445 47.670 ;
        RECT 88.765 47.440 89.485 47.700 ;
        RECT 88.605 47.150 88.835 47.290 ;
        RECT 77.355 46.280 77.585 46.370 ;
        RECT 78.145 46.280 78.375 46.390 ;
        RECT 83.645 46.370 84.225 46.540 ;
        RECT 88.465 46.380 88.855 47.150 ;
        RECT 89.395 47.140 89.625 47.290 ;
        RECT 89.385 46.400 89.755 47.140 ;
        RECT 92.685 46.960 93.115 51.930 ;
        RECT 93.625 51.920 93.855 51.985 ;
        RECT 94.765 51.920 94.995 51.985 ;
        RECT 93.565 46.920 93.965 51.920 ;
        RECT 94.645 46.920 95.045 51.920 ;
        RECT 95.555 51.890 95.785 51.985 ;
        RECT 100.035 51.950 100.265 52.055 ;
        RECT 95.495 46.920 95.925 51.890 ;
        RECT 99.905 50.230 100.275 51.950 ;
        RECT 100.825 51.830 101.055 52.055 ;
        RECT 104.115 51.920 104.345 51.975 ;
        RECT 100.035 50.055 100.265 50.230 ;
        RECT 100.815 50.150 101.185 51.830 ;
        RECT 100.825 50.055 101.055 50.150 ;
        RECT 100.185 49.610 100.905 49.870 ;
        RECT 93.115 46.550 93.575 46.780 ;
        RECT 95.045 46.660 95.505 46.780 ;
        RECT 94.895 46.550 95.505 46.660 ;
        RECT 97.955 46.590 98.725 47.660 ;
        RECT 100.045 47.430 100.765 47.690 ;
        RECT 99.885 47.140 100.115 47.280 ;
        RECT 88.605 46.290 88.835 46.380 ;
        RECT 89.395 46.290 89.625 46.400 ;
        RECT 94.895 46.380 95.475 46.550 ;
        RECT 99.745 46.370 100.135 47.140 ;
        RECT 100.675 47.130 100.905 47.280 ;
        RECT 100.665 46.390 101.035 47.130 ;
        RECT 103.965 46.950 104.395 51.920 ;
        RECT 104.905 51.910 105.135 51.975 ;
        RECT 106.045 51.910 106.275 51.975 ;
        RECT 104.845 46.910 105.245 51.910 ;
        RECT 105.925 46.910 106.325 51.910 ;
        RECT 106.835 51.880 107.065 51.975 ;
        RECT 111.305 51.950 111.535 52.055 ;
        RECT 106.775 46.910 107.205 51.880 ;
        RECT 111.175 50.230 111.545 51.950 ;
        RECT 112.095 51.830 112.325 52.055 ;
        RECT 115.385 51.920 115.615 51.975 ;
        RECT 111.305 50.055 111.535 50.230 ;
        RECT 112.085 50.150 112.455 51.830 ;
        RECT 112.095 50.055 112.325 50.150 ;
        RECT 111.455 49.610 112.175 49.870 ;
        RECT 104.395 46.540 104.855 46.770 ;
        RECT 106.325 46.650 106.785 46.770 ;
        RECT 106.175 46.540 106.785 46.650 ;
        RECT 109.225 46.590 109.995 47.660 ;
        RECT 111.315 47.430 112.035 47.690 ;
        RECT 111.155 47.140 111.385 47.280 ;
        RECT 99.885 46.280 100.115 46.370 ;
        RECT 100.675 46.280 100.905 46.390 ;
        RECT 106.175 46.370 106.755 46.540 ;
        RECT 111.015 46.370 111.405 47.140 ;
        RECT 111.945 47.130 112.175 47.280 ;
        RECT 111.935 46.390 112.305 47.130 ;
        RECT 115.235 46.950 115.665 51.920 ;
        RECT 116.175 51.910 116.405 51.975 ;
        RECT 117.315 51.910 117.545 51.975 ;
        RECT 116.115 46.910 116.515 51.910 ;
        RECT 117.195 46.910 117.595 51.910 ;
        RECT 118.105 51.880 118.335 51.975 ;
        RECT 122.555 51.950 122.785 52.055 ;
        RECT 118.045 46.910 118.475 51.880 ;
        RECT 122.425 50.230 122.795 51.950 ;
        RECT 123.345 51.830 123.575 52.055 ;
        RECT 126.635 51.920 126.865 51.975 ;
        RECT 122.555 50.055 122.785 50.230 ;
        RECT 123.335 50.150 123.705 51.830 ;
        RECT 123.345 50.055 123.575 50.150 ;
        RECT 122.705 49.610 123.425 49.870 ;
        RECT 115.665 46.540 116.125 46.770 ;
        RECT 117.595 46.650 118.055 46.770 ;
        RECT 117.445 46.540 118.055 46.650 ;
        RECT 120.475 46.590 121.245 47.660 ;
        RECT 122.565 47.430 123.285 47.690 ;
        RECT 122.405 47.140 122.635 47.280 ;
        RECT 111.155 46.280 111.385 46.370 ;
        RECT 111.945 46.280 112.175 46.390 ;
        RECT 117.445 46.370 118.025 46.540 ;
        RECT 122.265 46.370 122.655 47.140 ;
        RECT 123.195 47.130 123.425 47.280 ;
        RECT 123.185 46.390 123.555 47.130 ;
        RECT 126.485 46.950 126.915 51.920 ;
        RECT 127.425 51.910 127.655 51.975 ;
        RECT 128.565 51.910 128.795 51.975 ;
        RECT 127.365 46.910 127.765 51.910 ;
        RECT 128.445 46.910 128.845 51.910 ;
        RECT 129.355 51.880 129.585 51.975 ;
        RECT 129.295 46.910 129.725 51.880 ;
        RECT 126.915 46.540 127.375 46.770 ;
        RECT 128.845 46.650 129.305 46.770 ;
        RECT 128.695 46.540 129.305 46.650 ;
        RECT 122.405 46.280 122.635 46.370 ;
        RECT 123.195 46.280 123.425 46.390 ;
        RECT 128.695 46.370 129.275 46.540 ;
        RECT 21.505 45.950 21.965 46.180 ;
        RECT 32.705 45.960 33.165 46.190 ;
        RECT 43.925 45.930 44.385 46.160 ;
        RECT 55.175 45.910 55.635 46.140 ;
        RECT 66.395 45.900 66.855 46.130 ;
        RECT 77.635 45.890 78.095 46.120 ;
        RECT 88.885 45.900 89.345 46.130 ;
        RECT 100.165 45.890 100.625 46.120 ;
        RECT 111.435 45.890 111.895 46.120 ;
        RECT 122.685 45.890 123.145 46.120 ;
        RECT 29.055 45.020 41.225 45.030 ;
        RECT 17.855 45.005 41.225 45.020 ;
        RECT 15.900 45.000 41.225 45.005 ;
        RECT 15.900 44.980 52.445 45.000 ;
        RECT 15.900 44.970 63.695 44.980 ;
        RECT 15.900 44.960 74.915 44.970 ;
        RECT 85.235 44.960 97.405 44.970 ;
        RECT 15.900 43.880 131.205 44.960 ;
        RECT 15.900 43.870 30.025 43.880 ;
        RECT 15.900 43.855 18.690 43.870 ;
        RECT 15.900 41.620 17.050 43.855 ;
        RECT 40.275 43.850 131.205 43.880 ;
        RECT 51.525 43.830 131.205 43.850 ;
        RECT 62.745 43.820 131.205 43.830 ;
        RECT 73.985 43.810 86.155 43.820 ;
        RECT 96.515 43.810 131.205 43.820 ;
        RECT 29.015 43.330 41.185 43.340 ;
        RECT 17.815 43.310 41.185 43.330 ;
        RECT 142.830 43.320 144.150 43.340 ;
        RECT 17.815 43.290 52.405 43.310 ;
        RECT 140.750 43.300 144.150 43.320 ;
        RECT 17.815 43.280 63.655 43.290 ;
        RECT 119.895 43.280 144.150 43.300 ;
        RECT 17.815 43.270 74.875 43.280 ;
        RECT 85.195 43.270 97.365 43.280 ;
        RECT 108.685 43.270 144.150 43.280 ;
        RECT 17.815 42.180 144.150 43.270 ;
        RECT 18.755 42.150 144.150 42.180 ;
        RECT 18.755 42.120 131.165 42.150 ;
        RECT 18.755 42.090 109.655 42.120 ;
        RECT 18.755 42.080 98.445 42.090 ;
        RECT 41.325 42.070 98.445 42.080 ;
        RECT 142.830 42.070 144.150 42.150 ;
        RECT 41.325 42.060 87.205 42.070 ;
        RECT 75.035 42.050 87.205 42.060 ;
        RECT 15.900 41.540 19.685 41.620 ;
        RECT 142.070 41.610 146.210 41.640 ;
        RECT 119.855 41.590 146.210 41.610 ;
        RECT 108.645 41.550 146.210 41.590 ;
        RECT 15.900 41.520 42.165 41.540 ;
        RECT 97.445 41.530 146.210 41.550 ;
        RECT 15.900 41.510 75.875 41.520 ;
        RECT 86.235 41.510 146.210 41.530 ;
        RECT 15.900 40.500 146.210 41.510 ;
        RECT 15.900 40.480 142.320 40.500 ;
        RECT 15.900 40.470 140.920 40.480 ;
        RECT 18.715 40.460 140.920 40.470 ;
        RECT 142.070 40.460 142.250 40.480 ;
        RECT 18.715 40.440 120.815 40.460 ;
        RECT 18.715 40.400 109.615 40.440 ;
        RECT 18.715 40.390 98.405 40.400 ;
        RECT 41.285 40.380 98.405 40.390 ;
        RECT 41.285 40.370 87.165 40.380 ;
        RECT 74.995 40.360 87.165 40.370 ;
        RECT 26.775 39.230 27.235 39.460 ;
        RECT 38.055 39.230 38.515 39.460 ;
        RECT 49.345 39.210 49.805 39.440 ;
        RECT 60.565 39.210 61.025 39.440 ;
        RECT 71.765 39.210 72.225 39.440 ;
        RECT 83.055 39.200 83.515 39.430 ;
        RECT 94.295 39.220 94.755 39.450 ;
        RECT 105.505 39.240 105.965 39.470 ;
        RECT 116.705 39.280 117.165 39.510 ;
        RECT 127.915 39.300 128.375 39.530 ;
        RECT 20.645 38.810 21.225 38.980 ;
        RECT 26.495 38.960 26.725 39.070 ;
        RECT 27.285 38.980 27.515 39.070 ;
        RECT 20.615 38.700 21.225 38.810 ;
        RECT 20.615 38.580 21.075 38.700 ;
        RECT 22.545 38.580 23.005 38.810 ;
        RECT 20.195 33.470 20.625 38.440 ;
        RECT 20.335 33.375 20.565 33.470 ;
        RECT 21.075 33.440 21.475 38.440 ;
        RECT 22.155 33.440 22.555 38.440 ;
        RECT 21.125 33.375 21.355 33.440 ;
        RECT 22.265 33.375 22.495 33.440 ;
        RECT 23.005 33.430 23.435 38.400 ;
        RECT 26.365 38.220 26.735 38.960 ;
        RECT 26.495 38.070 26.725 38.220 ;
        RECT 27.265 38.210 27.655 38.980 ;
        RECT 31.925 38.810 32.505 38.980 ;
        RECT 37.775 38.960 38.005 39.070 ;
        RECT 38.565 38.980 38.795 39.070 ;
        RECT 27.285 38.070 27.515 38.210 ;
        RECT 26.635 37.660 27.355 37.920 ;
        RECT 28.675 37.690 29.445 38.760 ;
        RECT 31.895 38.700 32.505 38.810 ;
        RECT 31.895 38.580 32.355 38.700 ;
        RECT 33.825 38.580 34.285 38.810 ;
        RECT 26.495 35.480 27.215 35.740 ;
        RECT 26.345 35.200 26.575 35.295 ;
        RECT 26.215 33.520 26.585 35.200 ;
        RECT 27.135 35.120 27.365 35.295 ;
        RECT 23.055 33.375 23.285 33.430 ;
        RECT 26.345 33.295 26.575 33.520 ;
        RECT 27.125 33.400 27.495 35.120 ;
        RECT 31.475 33.470 31.905 38.440 ;
        RECT 27.135 33.295 27.365 33.400 ;
        RECT 31.615 33.375 31.845 33.470 ;
        RECT 32.355 33.440 32.755 38.440 ;
        RECT 33.435 33.440 33.835 38.440 ;
        RECT 32.405 33.375 32.635 33.440 ;
        RECT 33.545 33.375 33.775 33.440 ;
        RECT 34.285 33.430 34.715 38.400 ;
        RECT 37.645 38.220 38.015 38.960 ;
        RECT 37.775 38.070 38.005 38.220 ;
        RECT 38.545 38.210 38.935 38.980 ;
        RECT 43.215 38.790 43.795 38.960 ;
        RECT 49.065 38.940 49.295 39.050 ;
        RECT 49.855 38.960 50.085 39.050 ;
        RECT 38.565 38.070 38.795 38.210 ;
        RECT 37.915 37.660 38.635 37.920 ;
        RECT 39.955 37.690 40.725 38.760 ;
        RECT 43.185 38.680 43.795 38.790 ;
        RECT 43.185 38.560 43.645 38.680 ;
        RECT 45.115 38.560 45.575 38.790 ;
        RECT 37.775 35.480 38.495 35.740 ;
        RECT 37.625 35.200 37.855 35.295 ;
        RECT 37.495 33.520 37.865 35.200 ;
        RECT 38.415 35.120 38.645 35.295 ;
        RECT 34.335 33.375 34.565 33.430 ;
        RECT 37.625 33.295 37.855 33.520 ;
        RECT 38.405 33.400 38.775 35.120 ;
        RECT 42.765 33.450 43.195 38.420 ;
        RECT 38.415 33.295 38.645 33.400 ;
        RECT 42.905 33.355 43.135 33.450 ;
        RECT 43.645 33.420 44.045 38.420 ;
        RECT 44.725 33.420 45.125 38.420 ;
        RECT 43.695 33.355 43.925 33.420 ;
        RECT 44.835 33.355 45.065 33.420 ;
        RECT 45.575 33.410 46.005 38.380 ;
        RECT 48.935 38.200 49.305 38.940 ;
        RECT 49.065 38.050 49.295 38.200 ;
        RECT 49.835 38.190 50.225 38.960 ;
        RECT 54.435 38.790 55.015 38.960 ;
        RECT 60.285 38.940 60.515 39.050 ;
        RECT 61.075 38.960 61.305 39.050 ;
        RECT 49.855 38.050 50.085 38.190 ;
        RECT 49.205 37.640 49.925 37.900 ;
        RECT 51.245 37.670 52.015 38.740 ;
        RECT 54.405 38.680 55.015 38.790 ;
        RECT 54.405 38.560 54.865 38.680 ;
        RECT 56.335 38.560 56.795 38.790 ;
        RECT 49.065 35.460 49.785 35.720 ;
        RECT 48.915 35.180 49.145 35.275 ;
        RECT 48.785 33.500 49.155 35.180 ;
        RECT 49.705 35.100 49.935 35.275 ;
        RECT 45.625 33.355 45.855 33.410 ;
        RECT 48.915 33.275 49.145 33.500 ;
        RECT 49.695 33.380 50.065 35.100 ;
        RECT 53.985 33.450 54.415 38.420 ;
        RECT 49.705 33.275 49.935 33.380 ;
        RECT 54.125 33.355 54.355 33.450 ;
        RECT 54.865 33.420 55.265 38.420 ;
        RECT 55.945 33.420 56.345 38.420 ;
        RECT 54.915 33.355 55.145 33.420 ;
        RECT 56.055 33.355 56.285 33.420 ;
        RECT 56.795 33.410 57.225 38.380 ;
        RECT 60.155 38.200 60.525 38.940 ;
        RECT 60.285 38.050 60.515 38.200 ;
        RECT 61.055 38.190 61.445 38.960 ;
        RECT 65.635 38.790 66.215 38.960 ;
        RECT 71.485 38.940 71.715 39.050 ;
        RECT 72.275 38.960 72.505 39.050 ;
        RECT 61.075 38.050 61.305 38.190 ;
        RECT 60.425 37.640 61.145 37.900 ;
        RECT 62.465 37.670 63.235 38.740 ;
        RECT 65.605 38.680 66.215 38.790 ;
        RECT 65.605 38.560 66.065 38.680 ;
        RECT 67.535 38.560 67.995 38.790 ;
        RECT 60.285 35.460 61.005 35.720 ;
        RECT 60.135 35.180 60.365 35.275 ;
        RECT 60.005 33.500 60.375 35.180 ;
        RECT 60.925 35.100 61.155 35.275 ;
        RECT 56.845 33.355 57.075 33.410 ;
        RECT 60.135 33.275 60.365 33.500 ;
        RECT 60.915 33.380 61.285 35.100 ;
        RECT 65.185 33.450 65.615 38.420 ;
        RECT 60.925 33.275 61.155 33.380 ;
        RECT 65.325 33.355 65.555 33.450 ;
        RECT 66.065 33.420 66.465 38.420 ;
        RECT 67.145 33.420 67.545 38.420 ;
        RECT 66.115 33.355 66.345 33.420 ;
        RECT 67.255 33.355 67.485 33.420 ;
        RECT 67.995 33.410 68.425 38.380 ;
        RECT 71.355 38.200 71.725 38.940 ;
        RECT 71.485 38.050 71.715 38.200 ;
        RECT 72.255 38.190 72.645 38.960 ;
        RECT 76.925 38.780 77.505 38.950 ;
        RECT 82.775 38.930 83.005 39.040 ;
        RECT 83.565 38.950 83.795 39.040 ;
        RECT 72.275 38.050 72.505 38.190 ;
        RECT 71.625 37.640 72.345 37.900 ;
        RECT 73.665 37.670 74.435 38.740 ;
        RECT 76.895 38.670 77.505 38.780 ;
        RECT 76.895 38.550 77.355 38.670 ;
        RECT 78.825 38.550 79.285 38.780 ;
        RECT 71.485 35.460 72.205 35.720 ;
        RECT 71.335 35.180 71.565 35.275 ;
        RECT 71.205 33.500 71.575 35.180 ;
        RECT 72.125 35.100 72.355 35.275 ;
        RECT 68.045 33.355 68.275 33.410 ;
        RECT 71.335 33.275 71.565 33.500 ;
        RECT 72.115 33.380 72.485 35.100 ;
        RECT 76.475 33.440 76.905 38.410 ;
        RECT 72.125 33.275 72.355 33.380 ;
        RECT 76.615 33.345 76.845 33.440 ;
        RECT 77.355 33.410 77.755 38.410 ;
        RECT 78.435 33.410 78.835 38.410 ;
        RECT 77.405 33.345 77.635 33.410 ;
        RECT 78.545 33.345 78.775 33.410 ;
        RECT 79.285 33.400 79.715 38.370 ;
        RECT 82.645 38.190 83.015 38.930 ;
        RECT 82.775 38.040 83.005 38.190 ;
        RECT 83.545 38.180 83.935 38.950 ;
        RECT 88.165 38.800 88.745 38.970 ;
        RECT 94.015 38.950 94.245 39.060 ;
        RECT 94.805 38.970 95.035 39.060 ;
        RECT 83.565 38.040 83.795 38.180 ;
        RECT 82.915 37.630 83.635 37.890 ;
        RECT 84.955 37.660 85.725 38.730 ;
        RECT 88.135 38.690 88.745 38.800 ;
        RECT 88.135 38.570 88.595 38.690 ;
        RECT 90.065 38.570 90.525 38.800 ;
        RECT 82.775 35.450 83.495 35.710 ;
        RECT 82.625 35.170 82.855 35.265 ;
        RECT 82.495 33.490 82.865 35.170 ;
        RECT 83.415 35.090 83.645 35.265 ;
        RECT 79.335 33.345 79.565 33.400 ;
        RECT 82.625 33.265 82.855 33.490 ;
        RECT 83.405 33.370 83.775 35.090 ;
        RECT 87.715 33.460 88.145 38.430 ;
        RECT 83.415 33.265 83.645 33.370 ;
        RECT 87.855 33.365 88.085 33.460 ;
        RECT 88.595 33.430 88.995 38.430 ;
        RECT 89.675 33.430 90.075 38.430 ;
        RECT 88.645 33.365 88.875 33.430 ;
        RECT 89.785 33.365 90.015 33.430 ;
        RECT 90.525 33.420 90.955 38.390 ;
        RECT 93.885 38.210 94.255 38.950 ;
        RECT 94.015 38.060 94.245 38.210 ;
        RECT 94.785 38.200 95.175 38.970 ;
        RECT 99.375 38.820 99.955 38.990 ;
        RECT 105.225 38.970 105.455 39.080 ;
        RECT 106.015 38.990 106.245 39.080 ;
        RECT 94.805 38.060 95.035 38.200 ;
        RECT 94.155 37.650 94.875 37.910 ;
        RECT 96.195 37.680 96.965 38.750 ;
        RECT 99.345 38.710 99.955 38.820 ;
        RECT 99.345 38.590 99.805 38.710 ;
        RECT 101.275 38.590 101.735 38.820 ;
        RECT 94.015 35.470 94.735 35.730 ;
        RECT 93.865 35.190 94.095 35.285 ;
        RECT 93.735 33.510 94.105 35.190 ;
        RECT 94.655 35.110 94.885 35.285 ;
        RECT 90.575 33.365 90.805 33.420 ;
        RECT 93.865 33.285 94.095 33.510 ;
        RECT 94.645 33.390 95.015 35.110 ;
        RECT 98.925 33.480 99.355 38.450 ;
        RECT 94.655 33.285 94.885 33.390 ;
        RECT 99.065 33.385 99.295 33.480 ;
        RECT 99.805 33.450 100.205 38.450 ;
        RECT 100.885 33.450 101.285 38.450 ;
        RECT 99.855 33.385 100.085 33.450 ;
        RECT 100.995 33.385 101.225 33.450 ;
        RECT 101.735 33.440 102.165 38.410 ;
        RECT 105.095 38.230 105.465 38.970 ;
        RECT 105.225 38.080 105.455 38.230 ;
        RECT 105.995 38.220 106.385 38.990 ;
        RECT 110.575 38.860 111.155 39.030 ;
        RECT 116.425 39.010 116.655 39.120 ;
        RECT 117.215 39.030 117.445 39.120 ;
        RECT 106.015 38.080 106.245 38.220 ;
        RECT 105.365 37.670 106.085 37.930 ;
        RECT 107.405 37.700 108.175 38.770 ;
        RECT 110.545 38.750 111.155 38.860 ;
        RECT 110.545 38.630 111.005 38.750 ;
        RECT 112.475 38.630 112.935 38.860 ;
        RECT 105.225 35.490 105.945 35.750 ;
        RECT 105.075 35.210 105.305 35.305 ;
        RECT 104.945 33.530 105.315 35.210 ;
        RECT 105.865 35.130 106.095 35.305 ;
        RECT 101.785 33.385 102.015 33.440 ;
        RECT 105.075 33.305 105.305 33.530 ;
        RECT 105.855 33.410 106.225 35.130 ;
        RECT 110.125 33.520 110.555 38.490 ;
        RECT 110.265 33.425 110.495 33.520 ;
        RECT 111.005 33.490 111.405 38.490 ;
        RECT 112.085 33.490 112.485 38.490 ;
        RECT 111.055 33.425 111.285 33.490 ;
        RECT 112.195 33.425 112.425 33.490 ;
        RECT 112.935 33.480 113.365 38.450 ;
        RECT 116.295 38.270 116.665 39.010 ;
        RECT 116.425 38.120 116.655 38.270 ;
        RECT 117.195 38.260 117.585 39.030 ;
        RECT 121.785 38.880 122.365 39.050 ;
        RECT 127.635 39.030 127.865 39.140 ;
        RECT 128.425 39.050 128.655 39.140 ;
        RECT 117.215 38.120 117.445 38.260 ;
        RECT 116.565 37.710 117.285 37.970 ;
        RECT 118.605 37.740 119.375 38.810 ;
        RECT 121.755 38.770 122.365 38.880 ;
        RECT 121.755 38.650 122.215 38.770 ;
        RECT 123.685 38.650 124.145 38.880 ;
        RECT 116.425 35.530 117.145 35.790 ;
        RECT 116.275 35.250 116.505 35.345 ;
        RECT 116.145 33.570 116.515 35.250 ;
        RECT 117.065 35.170 117.295 35.345 ;
        RECT 112.985 33.425 113.215 33.480 ;
        RECT 105.865 33.305 106.095 33.410 ;
        RECT 116.275 33.345 116.505 33.570 ;
        RECT 117.055 33.450 117.425 35.170 ;
        RECT 121.335 33.540 121.765 38.510 ;
        RECT 117.065 33.345 117.295 33.450 ;
        RECT 121.475 33.445 121.705 33.540 ;
        RECT 122.215 33.510 122.615 38.510 ;
        RECT 123.295 33.510 123.695 38.510 ;
        RECT 122.265 33.445 122.495 33.510 ;
        RECT 123.405 33.445 123.635 33.510 ;
        RECT 124.145 33.500 124.575 38.470 ;
        RECT 127.505 38.290 127.875 39.030 ;
        RECT 127.635 38.140 127.865 38.290 ;
        RECT 128.405 38.280 128.795 39.050 ;
        RECT 128.425 38.140 128.655 38.280 ;
        RECT 127.775 37.730 128.495 37.990 ;
        RECT 129.815 37.760 130.585 38.830 ;
        RECT 142.850 37.630 144.170 38.900 ;
        RECT 127.635 35.550 128.355 35.810 ;
        RECT 127.485 35.270 127.715 35.365 ;
        RECT 127.355 33.590 127.725 35.270 ;
        RECT 128.275 35.190 128.505 35.365 ;
        RECT 124.195 33.445 124.425 33.500 ;
        RECT 127.485 33.365 127.715 33.590 ;
        RECT 128.265 33.470 128.635 35.190 ;
        RECT 128.275 33.365 128.505 33.470 ;
        RECT 20.615 32.940 21.075 33.170 ;
        RECT 22.545 33.130 23.005 33.170 ;
        RECT 22.485 32.850 23.115 33.130 ;
        RECT 26.625 32.860 27.085 33.090 ;
        RECT 31.895 32.940 32.355 33.170 ;
        RECT 33.825 33.130 34.285 33.170 ;
        RECT 33.765 32.850 34.395 33.130 ;
        RECT 37.905 32.860 38.365 33.090 ;
        RECT 43.185 32.920 43.645 33.150 ;
        RECT 45.115 33.110 45.575 33.150 ;
        RECT 45.055 32.830 45.685 33.110 ;
        RECT 49.195 32.840 49.655 33.070 ;
        RECT 54.405 32.920 54.865 33.150 ;
        RECT 56.335 33.110 56.795 33.150 ;
        RECT 56.275 32.830 56.905 33.110 ;
        RECT 60.415 32.840 60.875 33.070 ;
        RECT 65.605 32.920 66.065 33.150 ;
        RECT 67.535 33.110 67.995 33.150 ;
        RECT 67.475 32.830 68.105 33.110 ;
        RECT 71.615 32.840 72.075 33.070 ;
        RECT 76.895 32.910 77.355 33.140 ;
        RECT 78.825 33.100 79.285 33.140 ;
        RECT 78.765 32.820 79.395 33.100 ;
        RECT 82.905 32.830 83.365 33.060 ;
        RECT 88.135 32.930 88.595 33.160 ;
        RECT 90.065 33.120 90.525 33.160 ;
        RECT 90.005 32.840 90.635 33.120 ;
        RECT 94.145 32.850 94.605 33.080 ;
        RECT 99.345 32.950 99.805 33.180 ;
        RECT 101.275 33.140 101.735 33.180 ;
        RECT 101.215 32.860 101.845 33.140 ;
        RECT 105.355 32.870 105.815 33.100 ;
        RECT 110.545 32.990 111.005 33.220 ;
        RECT 112.475 33.180 112.935 33.220 ;
        RECT 112.415 32.900 113.045 33.180 ;
        RECT 116.555 32.910 117.015 33.140 ;
        RECT 121.755 33.010 122.215 33.240 ;
        RECT 123.685 33.200 124.145 33.240 ;
        RECT 123.625 32.920 124.255 33.200 ;
        RECT 127.765 32.930 128.225 33.160 ;
        RECT 23.185 30.880 27.925 31.180 ;
        RECT 34.465 30.880 39.205 31.180 ;
        RECT 45.755 30.860 50.495 31.160 ;
        RECT 56.975 30.860 61.715 31.160 ;
        RECT 68.175 30.860 72.915 31.160 ;
        RECT 79.465 30.850 84.205 31.150 ;
        RECT 90.705 30.870 95.445 31.170 ;
        RECT 101.915 30.890 106.655 31.190 ;
        RECT 113.115 30.930 117.855 31.230 ;
        RECT 124.325 30.950 129.065 31.250 ;
        RECT 19.485 20.270 19.905 30.160 ;
        RECT 19.585 20.090 19.815 20.270 ;
        RECT 20.805 20.260 21.175 30.210 ;
        RECT 20.875 20.090 21.105 20.260 ;
        RECT 21.935 20.220 22.305 30.170 ;
        RECT 27.255 20.270 27.615 30.190 ;
        RECT 30.765 20.270 31.185 30.160 ;
        RECT 22.015 20.090 22.245 20.220 ;
        RECT 27.305 20.090 27.535 20.270 ;
        RECT 30.865 20.090 31.095 20.270 ;
        RECT 32.085 20.260 32.455 30.210 ;
        RECT 32.155 20.090 32.385 20.260 ;
        RECT 33.215 20.220 33.585 30.170 ;
        RECT 38.535 20.270 38.895 30.190 ;
        RECT 33.295 20.090 33.525 20.220 ;
        RECT 38.585 20.090 38.815 20.270 ;
        RECT 42.055 20.250 42.475 30.140 ;
        RECT 42.155 20.070 42.385 20.250 ;
        RECT 43.375 20.240 43.745 30.190 ;
        RECT 43.445 20.070 43.675 20.240 ;
        RECT 44.505 20.200 44.875 30.150 ;
        RECT 49.825 20.250 50.185 30.170 ;
        RECT 53.275 20.250 53.695 30.140 ;
        RECT 44.585 20.070 44.815 20.200 ;
        RECT 49.875 20.070 50.105 20.250 ;
        RECT 53.375 20.070 53.605 20.250 ;
        RECT 54.595 20.240 54.965 30.190 ;
        RECT 54.665 20.070 54.895 20.240 ;
        RECT 55.725 20.200 56.095 30.150 ;
        RECT 61.045 20.250 61.405 30.170 ;
        RECT 64.475 20.250 64.895 30.140 ;
        RECT 55.805 20.070 56.035 20.200 ;
        RECT 61.095 20.070 61.325 20.250 ;
        RECT 64.575 20.070 64.805 20.250 ;
        RECT 65.795 20.240 66.165 30.190 ;
        RECT 65.865 20.070 66.095 20.240 ;
        RECT 66.925 20.200 67.295 30.150 ;
        RECT 72.245 20.250 72.605 30.170 ;
        RECT 67.005 20.070 67.235 20.200 ;
        RECT 72.295 20.070 72.525 20.250 ;
        RECT 75.765 20.240 76.185 30.130 ;
        RECT 75.865 20.060 76.095 20.240 ;
        RECT 77.085 20.230 77.455 30.180 ;
        RECT 77.155 20.060 77.385 20.230 ;
        RECT 78.215 20.190 78.585 30.140 ;
        RECT 83.535 20.240 83.895 30.160 ;
        RECT 87.005 20.260 87.425 30.150 ;
        RECT 78.295 20.060 78.525 20.190 ;
        RECT 83.585 20.060 83.815 20.240 ;
        RECT 87.105 20.080 87.335 20.260 ;
        RECT 88.325 20.250 88.695 30.200 ;
        RECT 88.395 20.080 88.625 20.250 ;
        RECT 89.455 20.210 89.825 30.160 ;
        RECT 94.775 20.260 95.135 30.180 ;
        RECT 98.215 20.280 98.635 30.170 ;
        RECT 89.535 20.080 89.765 20.210 ;
        RECT 94.825 20.080 95.055 20.260 ;
        RECT 98.315 20.100 98.545 20.280 ;
        RECT 99.535 20.270 99.905 30.220 ;
        RECT 99.605 20.100 99.835 20.270 ;
        RECT 100.665 20.230 101.035 30.180 ;
        RECT 105.985 20.280 106.345 30.200 ;
        RECT 109.415 20.320 109.835 30.210 ;
        RECT 100.745 20.100 100.975 20.230 ;
        RECT 106.035 20.100 106.265 20.280 ;
        RECT 109.515 20.140 109.745 20.320 ;
        RECT 110.735 20.310 111.105 30.260 ;
        RECT 110.805 20.140 111.035 20.310 ;
        RECT 111.865 20.270 112.235 30.220 ;
        RECT 117.185 20.320 117.545 30.240 ;
        RECT 120.625 20.340 121.045 30.230 ;
        RECT 111.945 20.140 112.175 20.270 ;
        RECT 117.235 20.140 117.465 20.320 ;
        RECT 120.725 20.160 120.955 20.340 ;
        RECT 121.945 20.330 122.315 30.280 ;
        RECT 122.015 20.160 122.245 20.330 ;
        RECT 123.075 20.290 123.445 30.240 ;
        RECT 128.395 20.340 128.755 30.260 ;
        RECT 123.155 20.160 123.385 20.290 ;
        RECT 128.445 20.160 128.675 20.340 ;
        RECT 132.345 20.170 132.755 30.180 ;
        RECT 137.735 30.120 137.965 30.130 ;
        RECT 132.445 20.130 132.675 20.170 ;
        RECT 137.665 20.080 138.055 30.120 ;
        RECT 19.775 19.610 20.925 19.920 ;
        RECT 22.185 19.620 27.335 19.900 ;
        RECT 31.055 19.610 32.205 19.920 ;
        RECT 33.465 19.620 38.615 19.900 ;
        RECT 42.345 19.590 43.495 19.900 ;
        RECT 44.755 19.600 49.905 19.880 ;
        RECT 53.565 19.590 54.715 19.900 ;
        RECT 55.975 19.600 61.125 19.880 ;
        RECT 64.765 19.590 65.915 19.900 ;
        RECT 67.175 19.600 72.325 19.880 ;
        RECT 76.055 19.580 77.205 19.890 ;
        RECT 78.465 19.590 83.615 19.870 ;
        RECT 87.295 19.600 88.445 19.910 ;
        RECT 89.705 19.610 94.855 19.890 ;
        RECT 98.505 19.620 99.655 19.930 ;
        RECT 100.915 19.630 106.065 19.910 ;
        RECT 109.705 19.660 110.855 19.970 ;
        RECT 112.115 19.670 117.265 19.950 ;
        RECT 120.915 19.680 122.065 19.990 ;
        RECT 123.325 19.690 128.475 19.970 ;
        RECT 132.635 19.640 138.025 19.930 ;
        RECT 142.940 19.110 144.080 37.630 ;
        RECT 13.940 18.460 17.635 18.530 ;
        RECT 117.755 18.510 131.425 18.530 ;
        RECT 106.545 18.470 131.425 18.510 ;
        RECT 13.940 18.440 41.565 18.460 ;
        RECT 95.345 18.450 131.425 18.470 ;
        RECT 13.940 18.430 75.275 18.440 ;
        RECT 84.135 18.430 131.425 18.450 ;
        RECT 13.940 17.380 131.425 18.430 ;
        RECT 142.890 17.990 144.140 19.110 ;
        RECT 145.070 18.880 146.210 40.500 ;
        RECT 145.030 17.960 146.250 18.880 ;
        RECT 13.950 17.370 15.100 17.380 ;
        RECT 16.615 17.360 120.215 17.380 ;
        RECT 16.615 17.320 109.015 17.360 ;
        RECT 16.615 17.310 97.805 17.320 ;
        RECT 39.185 17.300 97.805 17.310 ;
        RECT 39.185 17.290 86.565 17.300 ;
        RECT 72.895 17.280 86.565 17.290 ;
        RECT 117.765 16.950 140.620 16.960 ;
        RECT 142.040 16.950 148.010 16.980 ;
        RECT 117.765 16.940 148.010 16.950 ;
        RECT 106.555 16.900 148.010 16.940 ;
        RECT 16.625 16.870 41.575 16.890 ;
        RECT 95.355 16.880 148.010 16.900 ;
        RECT 16.625 16.860 75.285 16.870 ;
        RECT 84.145 16.860 148.010 16.880 ;
        RECT 16.625 15.840 148.010 16.860 ;
        RECT 16.625 15.820 142.660 15.840 ;
        RECT 16.625 15.810 140.620 15.820 ;
        RECT 142.040 15.810 142.660 15.820 ;
        RECT 16.625 15.790 120.225 15.810 ;
        RECT 16.625 15.750 109.025 15.790 ;
        RECT 16.625 15.740 97.815 15.750 ;
        RECT 39.195 15.730 97.815 15.740 ;
        RECT 39.195 15.720 86.575 15.730 ;
        RECT 72.905 15.710 86.575 15.720 ;
        RECT 131.215 15.460 132.585 15.470 ;
        RECT 12.290 15.390 17.625 15.450 ;
        RECT 117.795 15.440 132.785 15.460 ;
        RECT 106.585 15.400 132.785 15.440 ;
        RECT 12.290 15.370 41.585 15.390 ;
        RECT 95.385 15.380 132.785 15.400 ;
        RECT 12.290 15.360 75.295 15.370 ;
        RECT 84.175 15.360 132.785 15.380 ;
        RECT 12.290 14.320 132.785 15.360 ;
        RECT 142.905 15.040 144.045 15.050 ;
        RECT 12.290 14.310 131.445 14.320 ;
        RECT 12.290 14.300 120.235 14.310 ;
        RECT 12.320 14.280 13.470 14.300 ;
        RECT 16.655 14.290 120.235 14.300 ;
        RECT 16.655 14.250 109.035 14.290 ;
        RECT 16.655 14.240 97.825 14.250 ;
        RECT 39.225 14.230 97.825 14.240 ;
        RECT 39.225 14.220 86.585 14.230 ;
        RECT 72.935 14.210 86.585 14.220 ;
        RECT 142.850 13.920 144.100 15.040 ;
        RECT 145.020 14.870 146.160 14.980 ;
        RECT 144.980 13.950 146.200 14.870 ;
        RECT 16.965 13.800 17.435 13.810 ;
        RECT 10.800 13.780 17.435 13.800 ;
        RECT 10.800 13.720 17.555 13.780 ;
        RECT 117.845 13.770 131.445 13.790 ;
        RECT 106.635 13.730 131.445 13.770 ;
        RECT 10.800 13.700 41.585 13.720 ;
        RECT 95.435 13.710 131.445 13.730 ;
        RECT 10.800 13.690 75.295 13.700 ;
        RECT 84.225 13.690 131.445 13.710 ;
        RECT 10.800 12.650 131.445 13.690 ;
        RECT 16.705 12.640 131.445 12.650 ;
        RECT 16.705 12.620 120.235 12.640 ;
        RECT 16.705 12.580 109.035 12.620 ;
        RECT 16.705 12.570 97.825 12.580 ;
        RECT 39.275 12.560 97.825 12.570 ;
        RECT 39.275 12.550 86.585 12.560 ;
        RECT 72.985 12.540 86.585 12.550 ;
        RECT 128.755 12.240 130.465 12.250 ;
        RECT 117.545 12.220 119.255 12.230 ;
        RECT 106.345 12.180 108.055 12.190 ;
        RECT 27.615 12.170 29.325 12.180 ;
        RECT 38.895 12.170 40.605 12.180 ;
        RECT 25.675 11.030 29.325 12.170 ;
        RECT 36.955 11.030 40.605 12.170 ;
        RECT 95.135 12.160 96.845 12.170 ;
        RECT 50.185 12.150 51.895 12.160 ;
        RECT 61.405 12.150 63.115 12.160 ;
        RECT 72.605 12.150 74.315 12.160 ;
        RECT 25.675 11.020 27.625 11.030 ;
        RECT 36.955 11.020 38.905 11.030 ;
        RECT 48.245 11.010 51.895 12.150 ;
        RECT 59.465 11.010 63.115 12.150 ;
        RECT 70.665 11.010 74.315 12.150 ;
        RECT 83.895 12.140 85.605 12.150 ;
        RECT 48.245 11.000 50.195 11.010 ;
        RECT 59.465 11.000 61.415 11.010 ;
        RECT 70.665 11.000 72.615 11.010 ;
        RECT 81.955 11.000 85.605 12.140 ;
        RECT 93.195 11.020 96.845 12.160 ;
        RECT 104.405 11.040 108.055 12.180 ;
        RECT 115.605 11.080 119.255 12.220 ;
        RECT 126.815 11.100 130.465 12.240 ;
        RECT 126.815 11.090 128.765 11.100 ;
        RECT 115.605 11.070 117.555 11.080 ;
        RECT 104.405 11.030 106.355 11.040 ;
        RECT 93.195 11.010 95.145 11.020 ;
        RECT 81.955 10.990 83.905 11.000 ;
        RECT 142.905 8.580 144.045 13.920 ;
        RECT 74.420 7.440 144.045 8.580 ;
        RECT 74.420 1.410 75.560 7.440 ;
        RECT 145.020 6.630 146.160 13.950 ;
        RECT 93.650 5.490 146.160 6.630 ;
        RECT 93.650 1.480 94.790 5.490 ;
        RECT 146.870 4.560 148.010 15.840 ;
        RECT 113.130 3.420 148.010 4.560 ;
        RECT 113.130 1.610 114.270 3.420 ;
        RECT 149.460 2.770 150.600 64.660 ;
        RECT 131.940 1.880 150.600 2.770 ;
        RECT 131.800 1.630 150.600 1.880 ;
        RECT 74.290 0.160 75.680 1.410 ;
        RECT 93.500 0.230 94.890 1.480 ;
        RECT 112.900 0.360 114.290 1.610 ;
        RECT 131.800 1.380 133.490 1.630 ;
        RECT 151.730 1.420 152.870 66.900 ;
        RECT 131.800 0.430 133.540 1.380 ;
        RECT 113.130 0.330 114.270 0.360 ;
        RECT 151.600 0.300 152.970 1.420 ;
        RECT 93.650 0.150 94.790 0.230 ;
      LAYER met2 ;
        RECT 135.390 223.830 136.740 225.230 ;
        RECT 138.180 223.760 139.530 225.160 ;
        RECT 143.230 223.790 144.580 225.190 ;
        RECT 10.680 214.250 12.220 214.620 ;
        RECT 37.470 214.250 39.010 214.620 ;
        RECT 64.260 214.250 65.800 214.620 ;
        RECT 91.050 214.250 92.590 214.620 ;
        RECT 24.075 211.530 25.615 211.900 ;
        RECT 50.865 211.530 52.405 211.900 ;
        RECT 77.655 211.530 79.195 211.900 ;
        RECT 104.445 211.530 105.985 211.900 ;
        RECT 63.510 210.025 63.770 210.345 ;
        RECT 69.030 210.025 69.290 210.345 ;
        RECT 51.550 209.685 51.810 210.005 ;
        RECT 62.590 209.685 62.850 210.005 ;
        RECT 10.680 208.810 12.220 209.180 ;
        RECT 37.470 208.810 39.010 209.180 ;
        RECT 51.610 208.645 51.750 209.685 ;
        RECT 54.770 209.345 55.030 209.665 ;
        RECT 51.550 208.325 51.810 208.645 ;
        RECT 24.075 206.090 25.615 206.460 ;
        RECT 50.865 206.090 52.405 206.460 ;
        RECT 54.830 204.905 54.970 209.345 ;
        RECT 58.910 207.305 59.170 207.625 ;
        RECT 61.670 207.305 61.930 207.625 ;
        RECT 56.610 206.625 56.870 206.945 ;
        RECT 56.670 205.245 56.810 206.625 ;
        RECT 56.610 204.925 56.870 205.245 ;
        RECT 54.770 204.585 55.030 204.905 ;
        RECT 55.230 203.905 55.490 204.225 ;
        RECT 10.680 203.370 12.220 203.740 ;
        RECT 37.470 203.370 39.010 203.740 ;
        RECT 55.290 203.205 55.430 203.905 ;
        RECT 55.230 202.885 55.490 203.205 ;
        RECT 56.670 202.865 56.810 204.925 ;
        RECT 57.990 203.905 58.250 204.225 ;
        RECT 56.610 202.545 56.870 202.865 ;
        RECT 24.075 200.650 25.615 201.020 ;
        RECT 50.865 200.650 52.405 201.020 ;
        RECT 46.030 199.145 46.290 199.465 ;
        RECT 47.870 199.145 48.130 199.465 ;
        RECT 52.470 199.145 52.730 199.465 ;
        RECT 40.050 198.465 40.310 198.785 ;
        RECT 44.190 198.465 44.450 198.785 ;
        RECT 10.680 197.930 12.220 198.300 ;
        RECT 37.470 197.930 39.010 198.300 ;
        RECT 40.110 197.425 40.250 198.465 ;
        RECT 40.050 197.105 40.310 197.425 ;
        RECT 44.250 196.745 44.390 198.465 ;
        RECT 33.150 196.425 33.410 196.745 ;
        RECT 44.190 196.425 44.450 196.745 ;
        RECT 44.650 196.425 44.910 196.745 ;
        RECT 24.075 195.210 25.615 195.580 ;
        RECT 29.930 193.705 30.190 194.025 ;
        RECT 28.090 193.025 28.350 193.345 ;
        RECT 10.680 192.490 12.220 192.860 ;
        RECT 19.350 192.005 19.610 192.325 ;
        RECT 19.410 188.585 19.550 192.005 ;
        RECT 28.150 191.645 28.290 193.025 ;
        RECT 29.990 192.325 30.130 193.705 ;
        RECT 31.310 193.025 31.570 193.345 ;
        RECT 29.930 192.005 30.190 192.325 ;
        RECT 28.090 191.325 28.350 191.645 ;
        RECT 25.790 190.985 26.050 191.305 ;
        RECT 30.390 190.985 30.650 191.305 ;
        RECT 24.075 189.770 25.615 190.140 ;
        RECT 25.850 189.605 25.990 190.985 ;
        RECT 26.710 190.305 26.970 190.625 ;
        RECT 25.790 189.285 26.050 189.605 ;
        RECT 19.350 188.265 19.610 188.585 ;
        RECT 10.680 187.050 12.220 187.420 ;
        RECT 10.680 181.610 12.220 181.980 ;
        RECT 18.890 180.335 19.150 180.425 ;
        RECT 19.410 180.335 19.550 188.265 ;
        RECT 26.770 186.205 26.910 190.305 ;
        RECT 29.470 188.605 29.730 188.925 ;
        RECT 28.090 187.925 28.350 188.245 ;
        RECT 28.150 186.885 28.290 187.925 ;
        RECT 28.090 186.565 28.350 186.885 ;
        RECT 26.710 185.885 26.970 186.205 ;
        RECT 24.075 184.330 25.615 184.700 ;
        RECT 20.730 182.825 20.990 183.145 ;
        RECT 18.890 180.195 19.550 180.335 ;
        RECT 18.890 180.105 19.150 180.195 ;
        RECT 19.410 177.705 19.550 180.195 ;
        RECT 20.790 178.725 20.930 182.825 ;
        RECT 24.410 182.145 24.670 182.465 ;
        RECT 24.470 180.425 24.610 182.145 ;
        RECT 29.530 181.105 29.670 188.605 ;
        RECT 29.470 180.785 29.730 181.105 ;
        RECT 27.630 180.445 27.890 180.765 ;
        RECT 24.410 180.105 24.670 180.425 ;
        RECT 27.170 180.105 27.430 180.425 ;
        RECT 22.110 179.425 22.370 179.745 ;
        RECT 20.730 178.405 20.990 178.725 ;
        RECT 22.170 177.705 22.310 179.425 ;
        RECT 24.075 178.890 25.615 179.260 ;
        RECT 27.230 177.705 27.370 180.105 ;
        RECT 27.690 178.725 27.830 180.445 ;
        RECT 28.550 180.105 28.810 180.425 ;
        RECT 27.630 178.405 27.890 178.725 ;
        RECT 28.610 178.045 28.750 180.105 ;
        RECT 28.550 177.725 28.810 178.045 ;
        RECT 19.350 177.385 19.610 177.705 ;
        RECT 22.110 177.385 22.370 177.705 ;
        RECT 27.170 177.385 27.430 177.705 ;
        RECT 10.680 176.170 12.220 176.540 ;
        RECT 19.410 175.665 19.550 177.385 ;
        RECT 27.230 175.665 27.370 177.385 ;
        RECT 19.350 175.345 19.610 175.665 ;
        RECT 23.490 175.345 23.750 175.665 ;
        RECT 27.170 175.345 27.430 175.665 ;
        RECT 19.410 172.605 19.550 175.345 ;
        RECT 20.270 175.005 20.530 175.325 ;
        RECT 19.350 172.285 19.610 172.605 ;
        RECT 14.750 171.945 15.010 172.265 ;
        RECT 10.680 170.730 12.220 171.100 ;
        RECT 14.810 169.885 14.950 171.945 ;
        RECT 17.970 171.265 18.230 171.585 ;
        RECT 15.670 169.905 15.930 170.225 ;
        RECT 14.750 169.565 15.010 169.885 ;
        RECT 10.680 165.290 12.220 165.660 ;
        RECT 14.810 164.445 14.950 169.565 ;
        RECT 15.730 166.145 15.870 169.905 ;
        RECT 18.030 169.545 18.170 171.265 ;
        RECT 20.330 170.565 20.470 175.005 ;
        RECT 21.190 173.985 21.450 174.305 ;
        RECT 21.250 172.605 21.390 173.985 ;
        RECT 21.190 172.285 21.450 172.605 ;
        RECT 20.270 170.245 20.530 170.565 ;
        RECT 21.190 169.565 21.450 169.885 ;
        RECT 17.970 169.225 18.230 169.545 ;
        RECT 16.590 168.885 16.850 169.205 ;
        RECT 16.650 166.485 16.790 168.885 ;
        RECT 21.250 167.845 21.390 169.565 ;
        RECT 23.550 169.545 23.690 175.345 ;
        RECT 27.620 175.150 27.900 175.520 ;
        RECT 27.170 173.985 27.430 174.305 ;
        RECT 24.075 173.450 25.615 173.820 ;
        RECT 25.790 172.285 26.050 172.605 ;
        RECT 25.850 170.565 25.990 172.285 ;
        RECT 27.230 172.265 27.370 173.985 ;
        RECT 27.170 171.945 27.430 172.265 ;
        RECT 26.250 171.265 26.510 171.585 ;
        RECT 25.790 170.245 26.050 170.565 ;
        RECT 21.650 169.225 21.910 169.545 ;
        RECT 23.490 169.225 23.750 169.545 ;
        RECT 21.190 167.525 21.450 167.845 ;
        RECT 16.590 166.165 16.850 166.485 ;
        RECT 15.670 165.825 15.930 166.145 ;
        RECT 18.430 165.825 18.690 166.145 ;
        RECT 15.730 165.125 15.870 165.825 ;
        RECT 18.490 165.125 18.630 165.825 ;
        RECT 15.670 164.805 15.930 165.125 ;
        RECT 18.430 164.805 18.690 165.125 ;
        RECT 14.750 164.125 15.010 164.445 ;
        RECT 17.050 164.125 17.310 164.445 ;
        RECT 20.730 164.125 20.990 164.445 ;
        RECT 16.130 163.105 16.390 163.425 ;
        RECT 16.190 161.045 16.330 163.105 ;
        RECT 16.130 160.725 16.390 161.045 ;
        RECT 10.680 159.850 12.220 160.220 ;
        RECT 17.110 159.685 17.250 164.125 ;
        RECT 20.790 161.725 20.930 164.125 ;
        RECT 21.250 164.105 21.390 167.525 ;
        RECT 21.710 166.485 21.850 169.225 ;
        RECT 24.075 168.010 25.615 168.380 ;
        RECT 25.850 167.165 25.990 170.245 ;
        RECT 25.790 166.845 26.050 167.165 ;
        RECT 21.650 166.165 21.910 166.485 ;
        RECT 25.850 164.445 25.990 166.845 ;
        RECT 26.310 166.485 26.450 171.265 ;
        RECT 27.690 170.225 27.830 175.150 ;
        RECT 29.530 173.285 29.670 180.785 ;
        RECT 30.450 180.765 30.590 190.985 ;
        RECT 31.370 189.265 31.510 193.025 ;
        RECT 31.310 188.945 31.570 189.265 ;
        RECT 30.390 180.445 30.650 180.765 ;
        RECT 30.450 178.045 30.590 180.445 ;
        RECT 30.390 177.725 30.650 178.045 ;
        RECT 30.390 177.045 30.650 177.365 ;
        RECT 30.450 175.325 30.590 177.045 ;
        RECT 30.390 175.005 30.650 175.325 ;
        RECT 31.370 174.985 31.510 188.945 ;
        RECT 33.210 188.925 33.350 196.425 ;
        RECT 43.730 195.745 43.990 196.065 ;
        RECT 44.190 195.745 44.450 196.065 ;
        RECT 40.970 194.045 41.230 194.365 ;
        RECT 40.050 193.705 40.310 194.025 ;
        RECT 35.450 193.365 35.710 193.685 ;
        RECT 34.530 190.645 34.790 190.965 ;
        RECT 34.590 190.365 34.730 190.645 ;
        RECT 34.590 190.225 35.190 190.365 ;
        RECT 35.050 188.925 35.190 190.225 ;
        RECT 35.510 189.605 35.650 193.365 ;
        RECT 39.590 193.025 39.850 193.345 ;
        RECT 37.470 192.490 39.010 192.860 ;
        RECT 39.650 191.985 39.790 193.025 ;
        RECT 39.590 191.665 39.850 191.985 ;
        RECT 35.910 190.305 36.170 190.625 ;
        RECT 35.450 189.285 35.710 189.605 ;
        RECT 33.150 188.605 33.410 188.925 ;
        RECT 34.990 188.605 35.250 188.925 ;
        RECT 33.210 183.485 33.350 188.605 ;
        RECT 35.970 187.905 36.110 190.305 ;
        RECT 40.110 189.605 40.250 193.705 ;
        RECT 41.030 191.305 41.170 194.045 ;
        RECT 43.790 193.345 43.930 195.745 ;
        RECT 44.250 194.025 44.390 195.745 ;
        RECT 44.190 193.705 44.450 194.025 ;
        RECT 43.730 193.025 43.990 193.345 ;
        RECT 43.790 192.325 43.930 193.025 ;
        RECT 43.730 192.005 43.990 192.325 ;
        RECT 40.970 190.985 41.230 191.305 ;
        RECT 40.050 189.285 40.310 189.605 ;
        RECT 35.910 187.585 36.170 187.905 ;
        RECT 42.810 187.585 43.070 187.905 ;
        RECT 33.150 183.165 33.410 183.485 ;
        RECT 34.070 183.165 34.330 183.485 ;
        RECT 32.690 182.145 32.950 182.465 ;
        RECT 32.750 181.445 32.890 182.145 ;
        RECT 32.690 181.125 32.950 181.445 ;
        RECT 34.130 180.425 34.270 183.165 ;
        RECT 34.070 180.105 34.330 180.425 ;
        RECT 35.450 177.385 35.710 177.705 ;
        RECT 34.070 177.045 34.330 177.365 ;
        RECT 31.770 176.705 32.030 177.025 ;
        RECT 31.830 175.665 31.970 176.705 ;
        RECT 31.770 175.345 32.030 175.665 ;
        RECT 34.130 175.325 34.270 177.045 ;
        RECT 34.990 176.705 35.250 177.025 ;
        RECT 32.690 175.005 32.950 175.325 ;
        RECT 34.070 175.005 34.330 175.325 ;
        RECT 31.310 174.665 31.570 174.985 ;
        RECT 32.750 174.645 32.890 175.005 ;
        RECT 32.690 174.325 32.950 174.645 ;
        RECT 31.770 173.985 32.030 174.305 ;
        RECT 29.470 172.965 29.730 173.285 ;
        RECT 27.630 169.905 27.890 170.225 ;
        RECT 29.530 169.885 29.670 172.965 ;
        RECT 29.470 169.565 29.730 169.885 ;
        RECT 26.250 166.165 26.510 166.485 ;
        RECT 31.310 165.825 31.570 166.145 ;
        RECT 25.790 164.125 26.050 164.445 ;
        RECT 21.190 163.785 21.450 164.105 ;
        RECT 20.730 161.405 20.990 161.725 ;
        RECT 17.050 159.365 17.310 159.685 ;
        RECT 20.270 158.685 20.530 159.005 ;
        RECT 17.970 154.945 18.230 155.265 ;
        RECT 10.680 154.410 12.220 154.780 ;
        RECT 18.030 153.905 18.170 154.945 ;
        RECT 17.970 153.585 18.230 153.905 ;
        RECT 20.330 153.225 20.470 158.685 ;
        RECT 20.790 158.665 20.930 161.405 ;
        RECT 21.250 158.665 21.390 163.785 ;
        RECT 23.030 163.105 23.290 163.425 ;
        RECT 23.090 161.725 23.230 163.105 ;
        RECT 24.075 162.570 25.615 162.940 ;
        RECT 25.850 161.725 25.990 164.125 ;
        RECT 30.390 163.785 30.650 164.105 ;
        RECT 30.450 162.065 30.590 163.785 ;
        RECT 31.370 162.405 31.510 165.825 ;
        RECT 31.310 162.085 31.570 162.405 ;
        RECT 30.390 161.745 30.650 162.065 ;
        RECT 23.030 161.405 23.290 161.725 ;
        RECT 25.790 161.405 26.050 161.725 ;
        RECT 20.730 158.345 20.990 158.665 ;
        RECT 21.190 158.345 21.450 158.665 ;
        RECT 20.790 156.965 20.930 158.345 ;
        RECT 20.730 156.645 20.990 156.965 ;
        RECT 20.730 154.945 20.990 155.265 ;
        RECT 20.790 153.905 20.930 154.945 ;
        RECT 20.730 153.585 20.990 153.905 ;
        RECT 20.270 152.905 20.530 153.225 ;
        RECT 20.330 150.845 20.470 152.905 ;
        RECT 21.250 151.185 21.390 158.345 ;
        RECT 24.075 157.130 25.615 157.500 ;
        RECT 23.490 156.305 23.750 156.625 ;
        RECT 21.650 155.625 21.910 155.945 ;
        RECT 21.710 151.525 21.850 155.625 ;
        RECT 22.570 152.565 22.830 152.885 ;
        RECT 21.650 151.205 21.910 151.525 ;
        RECT 21.190 150.865 21.450 151.185 ;
        RECT 20.270 150.525 20.530 150.845 ;
        RECT 15.670 149.845 15.930 150.165 ;
        RECT 10.680 148.970 12.220 149.340 ;
        RECT 14.290 148.145 14.550 148.465 ;
        RECT 13.830 146.785 14.090 147.105 ;
        RECT 10.680 143.530 12.220 143.900 ;
        RECT 13.890 142.685 14.030 146.785 ;
        RECT 14.350 146.085 14.490 148.145 ;
        RECT 14.290 145.765 14.550 146.085 ;
        RECT 15.730 145.065 15.870 149.845 ;
        RECT 19.810 149.505 20.070 149.825 ;
        RECT 17.970 147.465 18.230 147.785 ;
        RECT 18.030 146.085 18.170 147.465 ;
        RECT 17.970 145.765 18.230 146.085 ;
        RECT 15.670 144.745 15.930 145.065 ;
        RECT 17.050 144.745 17.310 145.065 ;
        RECT 17.110 143.365 17.250 144.745 ;
        RECT 17.050 143.045 17.310 143.365 ;
        RECT 19.870 143.025 20.010 149.505 ;
        RECT 19.810 142.705 20.070 143.025 ;
        RECT 13.830 142.365 14.090 142.685 ;
        RECT 21.250 142.345 21.390 150.865 ;
        RECT 22.630 150.845 22.770 152.565 ;
        RECT 22.570 150.525 22.830 150.845 ;
        RECT 23.550 149.825 23.690 156.305 ;
        RECT 25.850 155.125 25.990 161.405 ;
        RECT 27.630 159.025 27.890 159.345 ;
        RECT 26.710 158.685 26.970 159.005 ;
        RECT 26.770 156.965 26.910 158.685 ;
        RECT 26.710 156.645 26.970 156.965 ;
        RECT 25.850 154.985 26.450 155.125 ;
        RECT 26.310 153.905 26.450 154.985 ;
        RECT 26.250 153.585 26.510 153.905 ;
        RECT 25.790 152.225 26.050 152.545 ;
        RECT 24.075 151.690 25.615 152.060 ;
        RECT 24.410 150.865 24.670 151.185 ;
        RECT 23.490 149.505 23.750 149.825 ;
        RECT 24.470 147.785 24.610 150.865 ;
        RECT 25.850 150.415 25.990 152.225 ;
        RECT 25.390 150.275 25.990 150.415 ;
        RECT 25.390 148.805 25.530 150.275 ;
        RECT 25.330 148.485 25.590 148.805 ;
        RECT 27.170 147.805 27.430 148.125 ;
        RECT 24.410 147.465 24.670 147.785 ;
        RECT 22.570 147.125 22.830 147.445 ;
        RECT 22.630 146.085 22.770 147.125 ;
        RECT 23.490 146.785 23.750 147.105 ;
        RECT 22.570 145.765 22.830 146.085 ;
        RECT 22.630 143.365 22.770 145.765 ;
        RECT 22.570 143.045 22.830 143.365 ;
        RECT 23.550 142.685 23.690 146.785 ;
        RECT 24.075 146.250 25.615 146.620 ;
        RECT 27.230 145.405 27.370 147.805 ;
        RECT 27.170 145.085 27.430 145.405 ;
        RECT 25.790 144.405 26.050 144.725 ;
        RECT 25.850 143.365 25.990 144.405 ;
        RECT 25.790 143.045 26.050 143.365 ;
        RECT 23.490 142.365 23.750 142.685 ;
        RECT 21.190 142.025 21.450 142.345 ;
        RECT 24.075 140.810 25.615 141.180 ;
        RECT 10.680 138.090 12.220 138.460 ;
        RECT 14.290 137.265 14.550 137.585 ;
        RECT 14.350 135.205 14.490 137.265 ;
        RECT 26.710 137.155 26.970 137.245 ;
        RECT 27.230 137.155 27.370 145.085 ;
        RECT 26.710 137.015 27.370 137.155 ;
        RECT 26.710 136.925 26.970 137.015 ;
        RECT 17.970 136.585 18.230 136.905 ;
        RECT 21.190 136.585 21.450 136.905 ;
        RECT 18.030 135.205 18.170 136.585 ;
        RECT 21.250 136.225 21.390 136.585 ;
        RECT 26.710 136.245 26.970 136.565 ;
        RECT 21.190 135.905 21.450 136.225 ;
        RECT 25.790 135.905 26.050 136.225 ;
        RECT 14.290 134.885 14.550 135.205 ;
        RECT 17.970 134.885 18.230 135.205 ;
        RECT 14.750 133.865 15.010 134.185 ;
        RECT 18.430 133.865 18.690 134.185 ;
        RECT 10.680 132.650 12.220 133.020 ;
        RECT 14.810 128.745 14.950 133.865 ;
        RECT 18.490 132.485 18.630 133.865 ;
        RECT 18.890 133.185 19.150 133.505 ;
        RECT 18.430 132.165 18.690 132.485 ;
        RECT 16.130 131.485 16.390 131.805 ;
        RECT 16.190 129.085 16.330 131.485 ;
        RECT 18.950 131.465 19.090 133.185 ;
        RECT 21.250 132.485 21.390 135.905 ;
        RECT 24.075 135.370 25.615 135.740 ;
        RECT 25.850 134.525 25.990 135.905 ;
        RECT 25.790 134.205 26.050 134.525 ;
        RECT 21.190 132.165 21.450 132.485 ;
        RECT 26.250 131.485 26.510 131.805 ;
        RECT 18.890 131.145 19.150 131.465 ;
        RECT 25.790 131.145 26.050 131.465 ;
        RECT 17.970 130.465 18.230 130.785 ;
        RECT 16.130 128.765 16.390 129.085 ;
        RECT 14.750 128.425 15.010 128.745 ;
        RECT 16.190 128.485 16.330 128.765 ;
        RECT 18.030 128.745 18.170 130.465 ;
        RECT 24.075 129.930 25.615 130.300 ;
        RECT 25.850 129.085 25.990 131.145 ;
        RECT 25.790 128.765 26.050 129.085 ;
        RECT 10.680 127.210 12.220 127.580 ;
        RECT 14.810 125.345 14.950 128.425 ;
        RECT 15.730 128.345 16.330 128.485 ;
        RECT 17.970 128.425 18.230 128.745 ;
        RECT 15.730 126.025 15.870 128.345 ;
        RECT 16.130 127.745 16.390 128.065 ;
        RECT 17.510 127.745 17.770 128.065 ;
        RECT 17.970 127.745 18.230 128.065 ;
        RECT 19.350 127.745 19.610 128.065 ;
        RECT 16.190 126.705 16.330 127.745 ;
        RECT 16.130 126.385 16.390 126.705 ;
        RECT 17.570 126.025 17.710 127.745 ;
        RECT 15.670 125.705 15.930 126.025 ;
        RECT 17.510 125.705 17.770 126.025 ;
        RECT 14.750 125.025 15.010 125.345 ;
        RECT 14.810 123.305 14.950 125.025 ;
        RECT 14.750 122.985 15.010 123.305 ;
        RECT 10.680 121.770 12.220 122.140 ;
        RECT 18.030 120.925 18.170 127.745 ;
        RECT 19.410 127.125 19.550 127.745 ;
        RECT 19.410 127.045 20.010 127.125 ;
        RECT 19.410 126.985 20.070 127.045 ;
        RECT 19.410 124.325 19.550 126.985 ;
        RECT 19.810 126.725 20.070 126.985 ;
        RECT 26.310 126.365 26.450 131.485 ;
        RECT 26.770 128.745 26.910 136.245 ;
        RECT 27.230 134.185 27.370 137.015 ;
        RECT 27.690 134.605 27.830 159.025 ;
        RECT 30.390 158.685 30.650 159.005 ;
        RECT 29.010 158.005 29.270 158.325 ;
        RECT 28.090 136.925 28.350 137.245 ;
        RECT 28.150 135.205 28.290 136.925 ;
        RECT 28.090 134.885 28.350 135.205 ;
        RECT 27.690 134.465 28.290 134.605 ;
        RECT 27.170 133.865 27.430 134.185 ;
        RECT 27.230 131.465 27.370 133.865 ;
        RECT 27.170 131.145 27.430 131.465 ;
        RECT 26.710 128.425 26.970 128.745 ;
        RECT 27.230 126.705 27.370 131.145 ;
        RECT 27.170 126.385 27.430 126.705 ;
        RECT 26.250 126.045 26.510 126.365 ;
        RECT 25.790 125.025 26.050 125.345 ;
        RECT 24.075 124.490 25.615 124.860 ;
        RECT 19.350 124.005 19.610 124.325 ;
        RECT 18.430 123.325 18.690 123.645 ;
        RECT 24.870 123.325 25.130 123.645 ;
        RECT 18.490 121.605 18.630 123.325 ;
        RECT 24.930 121.605 25.070 123.325 ;
        RECT 25.850 122.965 25.990 125.025 ;
        RECT 25.790 122.645 26.050 122.965 ;
        RECT 26.310 122.625 26.450 126.045 ;
        RECT 27.230 123.645 27.370 126.385 ;
        RECT 27.170 123.325 27.430 123.645 ;
        RECT 26.250 122.305 26.510 122.625 ;
        RECT 18.430 121.285 18.690 121.605 ;
        RECT 24.870 121.285 25.130 121.605 ;
        RECT 17.970 120.605 18.230 120.925 ;
        RECT 24.075 119.050 25.615 119.420 ;
        RECT 23.490 116.865 23.750 117.185 ;
        RECT 10.680 116.330 12.220 116.700 ;
        RECT 17.510 115.505 17.770 115.825 ;
        RECT 17.570 113.445 17.710 115.505 ;
        RECT 17.970 114.825 18.230 115.145 ;
        RECT 17.510 113.125 17.770 113.445 ;
        RECT 14.290 111.425 14.550 111.745 ;
        RECT 10.680 110.890 12.220 111.260 ;
        RECT 14.350 110.385 14.490 111.425 ;
        RECT 14.290 110.065 14.550 110.385 ;
        RECT 12.450 109.385 12.710 109.705 ;
        RECT 12.510 106.285 12.650 109.385 ;
        RECT 18.030 106.285 18.170 114.825 ;
        RECT 23.030 112.445 23.290 112.765 ;
        RECT 23.090 110.125 23.230 112.445 ;
        RECT 23.550 110.725 23.690 116.865 ;
        RECT 27.230 115.485 27.370 123.325 ;
        RECT 27.620 122.790 27.900 123.160 ;
        RECT 27.690 121.265 27.830 122.790 ;
        RECT 27.630 120.945 27.890 121.265 ;
        RECT 28.150 115.485 28.290 134.465 ;
        RECT 29.070 117.865 29.210 158.005 ;
        RECT 30.450 153.565 30.590 158.685 ;
        RECT 30.390 153.245 30.650 153.565 ;
        RECT 29.930 152.225 30.190 152.545 ;
        RECT 29.990 148.125 30.130 152.225 ;
        RECT 30.450 151.525 30.590 153.245 ;
        RECT 30.850 152.905 31.110 153.225 ;
        RECT 30.390 151.205 30.650 151.525 ;
        RECT 30.910 150.925 31.050 152.905 ;
        RECT 30.450 150.845 31.050 150.925 ;
        RECT 30.390 150.785 31.050 150.845 ;
        RECT 30.390 150.525 30.650 150.785 ;
        RECT 29.930 147.805 30.190 148.125 ;
        RECT 30.450 147.785 30.590 150.525 ;
        RECT 30.850 149.845 31.110 150.165 ;
        RECT 30.910 148.805 31.050 149.845 ;
        RECT 30.850 148.485 31.110 148.805 ;
        RECT 30.390 147.465 30.650 147.785 ;
        RECT 31.310 147.125 31.570 147.445 ;
        RECT 31.370 146.960 31.510 147.125 ;
        RECT 31.300 146.590 31.580 146.960 ;
        RECT 31.310 145.765 31.570 146.085 ;
        RECT 31.370 143.365 31.510 145.765 ;
        RECT 31.310 143.045 31.570 143.365 ;
        RECT 31.830 139.965 31.970 173.985 ;
        RECT 34.070 171.605 34.330 171.925 ;
        RECT 33.150 171.265 33.410 171.585 ;
        RECT 32.230 168.885 32.490 169.205 ;
        RECT 32.290 164.785 32.430 168.885 ;
        RECT 32.690 168.545 32.950 168.865 ;
        RECT 32.750 167.165 32.890 168.545 ;
        RECT 32.690 166.845 32.950 167.165 ;
        RECT 32.230 164.465 32.490 164.785 ;
        RECT 32.230 162.085 32.490 162.405 ;
        RECT 32.290 159.685 32.430 162.085 ;
        RECT 32.230 159.365 32.490 159.685 ;
        RECT 32.690 158.345 32.950 158.665 ;
        RECT 32.750 155.125 32.890 158.345 ;
        RECT 33.210 155.685 33.350 171.265 ;
        RECT 34.130 167.845 34.270 171.605 ;
        RECT 34.070 167.525 34.330 167.845 ;
        RECT 33.610 166.845 33.870 167.165 ;
        RECT 33.670 158.665 33.810 166.845 ;
        RECT 34.070 166.165 34.330 166.485 ;
        RECT 34.130 163.425 34.270 166.165 ;
        RECT 34.530 165.825 34.790 166.145 ;
        RECT 34.070 163.105 34.330 163.425 ;
        RECT 34.590 161.385 34.730 165.825 ;
        RECT 34.530 161.065 34.790 161.385 ;
        RECT 33.610 158.345 33.870 158.665 ;
        RECT 33.610 157.665 33.870 157.985 ;
        RECT 33.670 156.285 33.810 157.665 ;
        RECT 33.610 155.965 33.870 156.285 ;
        RECT 33.210 155.545 33.810 155.685 ;
        RECT 32.750 154.985 33.350 155.125 ;
        RECT 32.230 153.585 32.490 153.905 ;
        RECT 32.290 150.845 32.430 153.585 ;
        RECT 33.210 153.225 33.350 154.985 ;
        RECT 33.150 152.905 33.410 153.225 ;
        RECT 32.230 150.525 32.490 150.845 ;
        RECT 32.230 147.805 32.490 148.125 ;
        RECT 32.690 147.805 32.950 148.125 ;
        RECT 32.290 143.025 32.430 147.805 ;
        RECT 32.750 147.445 32.890 147.805 ;
        RECT 32.690 147.125 32.950 147.445 ;
        RECT 33.150 146.785 33.410 147.105 ;
        RECT 32.690 144.065 32.950 144.385 ;
        RECT 32.230 142.705 32.490 143.025 ;
        RECT 32.750 142.200 32.890 144.065 ;
        RECT 32.680 141.830 32.960 142.200 ;
        RECT 32.690 141.345 32.950 141.665 ;
        RECT 31.770 139.645 32.030 139.965 ;
        RECT 32.750 137.925 32.890 141.345 ;
        RECT 33.210 140.305 33.350 146.785 ;
        RECT 33.670 145.745 33.810 155.545 ;
        RECT 34.530 150.865 34.790 151.185 ;
        RECT 34.070 149.505 34.330 149.825 ;
        RECT 33.610 145.425 33.870 145.745 ;
        RECT 34.130 145.065 34.270 149.505 ;
        RECT 34.590 148.805 34.730 150.865 ;
        RECT 34.530 148.485 34.790 148.805 ;
        RECT 34.590 148.125 34.730 148.485 ;
        RECT 34.530 147.805 34.790 148.125 ;
        RECT 34.070 144.745 34.330 145.065 ;
        RECT 33.610 144.065 33.870 144.385 ;
        RECT 33.670 142.685 33.810 144.065 ;
        RECT 34.530 143.045 34.790 143.365 ;
        RECT 33.610 142.365 33.870 142.685 ;
        RECT 34.070 141.345 34.330 141.665 ;
        RECT 33.600 140.470 33.880 140.840 ;
        RECT 33.150 139.985 33.410 140.305 ;
        RECT 33.670 139.625 33.810 140.470 ;
        RECT 33.610 139.305 33.870 139.625 ;
        RECT 34.130 137.925 34.270 141.345 ;
        RECT 34.590 137.925 34.730 143.045 ;
        RECT 35.050 142.685 35.190 176.705 ;
        RECT 35.510 176.005 35.650 177.385 ;
        RECT 35.450 175.685 35.710 176.005 ;
        RECT 35.510 175.325 35.650 175.685 ;
        RECT 35.450 175.005 35.710 175.325 ;
        RECT 35.510 172.265 35.650 175.005 ;
        RECT 35.970 172.605 36.110 187.585 ;
        RECT 37.470 187.050 39.010 187.420 ;
        RECT 39.130 185.885 39.390 186.205 ;
        RECT 36.830 182.145 37.090 182.465 ;
        RECT 36.890 178.385 37.030 182.145 ;
        RECT 37.470 181.610 39.010 181.980 ;
        RECT 36.830 178.065 37.090 178.385 ;
        RECT 36.370 177.385 36.630 177.705 ;
        RECT 36.430 176.005 36.570 177.385 ;
        RECT 37.470 176.170 39.010 176.540 ;
        RECT 36.370 175.685 36.630 176.005 ;
        RECT 37.750 175.685 38.010 176.005 ;
        RECT 37.810 175.235 37.950 175.685 ;
        RECT 39.190 175.520 39.330 185.885 ;
        RECT 39.590 182.145 39.850 182.465 ;
        RECT 39.650 180.765 39.790 182.145 ;
        RECT 39.590 180.445 39.850 180.765 ;
        RECT 39.590 177.385 39.850 177.705 ;
        RECT 38.210 175.235 38.470 175.325 ;
        RECT 37.810 175.095 38.470 175.235 ;
        RECT 39.120 175.150 39.400 175.520 ;
        RECT 39.650 175.325 39.790 177.385 ;
        RECT 41.890 175.345 42.150 175.665 ;
        RECT 36.370 174.840 36.630 174.985 ;
        RECT 36.360 174.470 36.640 174.840 ;
        RECT 36.370 173.985 36.630 174.305 ;
        RECT 35.910 172.285 36.170 172.605 ;
        RECT 35.450 171.945 35.710 172.265 ;
        RECT 35.910 160.725 36.170 161.045 ;
        RECT 35.450 155.625 35.710 155.945 ;
        RECT 35.510 153.905 35.650 155.625 ;
        RECT 35.450 153.585 35.710 153.905 ;
        RECT 35.970 153.565 36.110 160.725 ;
        RECT 35.910 153.245 36.170 153.565 ;
        RECT 35.970 152.965 36.110 153.245 ;
        RECT 35.510 152.825 36.110 152.965 ;
        RECT 35.510 150.505 35.650 152.825 ;
        RECT 35.910 152.225 36.170 152.545 ;
        RECT 35.450 150.185 35.710 150.505 ;
        RECT 35.450 149.505 35.710 149.825 ;
        RECT 35.510 145.065 35.650 149.505 ;
        RECT 35.450 144.745 35.710 145.065 ;
        RECT 35.450 144.065 35.710 144.385 ;
        RECT 35.510 143.365 35.650 144.065 ;
        RECT 35.450 143.045 35.710 143.365 ;
        RECT 34.990 142.365 35.250 142.685 ;
        RECT 34.990 140.325 35.250 140.645 ;
        RECT 35.450 140.325 35.710 140.645 ;
        RECT 32.690 137.605 32.950 137.925 ;
        RECT 34.070 137.605 34.330 137.925 ;
        RECT 34.530 137.605 34.790 137.925 ;
        RECT 30.390 136.585 30.650 136.905 ;
        RECT 30.450 134.185 30.590 136.585 ;
        RECT 31.310 134.205 31.570 134.525 ;
        RECT 30.390 133.865 30.650 134.185 ;
        RECT 30.450 131.125 30.590 133.865 ;
        RECT 30.390 130.805 30.650 131.125 ;
        RECT 31.370 129.085 31.510 134.205 ;
        RECT 31.770 133.185 32.030 133.505 ;
        RECT 31.830 132.485 31.970 133.185 ;
        RECT 31.770 132.165 32.030 132.485 ;
        RECT 35.050 129.765 35.190 140.325 ;
        RECT 34.990 129.445 35.250 129.765 ;
        RECT 31.310 128.765 31.570 129.085 ;
        RECT 29.930 128.425 30.190 128.745 ;
        RECT 29.990 127.045 30.130 128.425 ;
        RECT 29.930 126.725 30.190 127.045 ;
        RECT 30.390 126.045 30.650 126.365 ;
        RECT 30.450 124.325 30.590 126.045 ;
        RECT 31.370 125.685 31.510 128.765 ;
        RECT 31.310 125.365 31.570 125.685 ;
        RECT 32.230 125.025 32.490 125.345 ;
        RECT 30.390 124.005 30.650 124.325 ;
        RECT 32.290 120.925 32.430 125.025 ;
        RECT 32.690 123.325 32.950 123.645 ;
        RECT 32.750 121.605 32.890 123.325 ;
        RECT 32.690 121.285 32.950 121.605 ;
        RECT 32.230 120.605 32.490 120.925 ;
        RECT 32.220 120.070 32.500 120.440 ;
        RECT 29.010 117.545 29.270 117.865 ;
        RECT 30.390 117.205 30.650 117.525 ;
        RECT 30.450 116.165 30.590 117.205 ;
        RECT 30.390 115.845 30.650 116.165 ;
        RECT 32.290 115.485 32.430 120.070 ;
        RECT 35.510 118.885 35.650 140.325 ;
        RECT 35.970 139.965 36.110 152.225 ;
        RECT 36.430 142.685 36.570 173.985 ;
        RECT 37.810 173.365 37.950 175.095 ;
        RECT 38.210 175.005 38.470 175.095 ;
        RECT 39.590 175.005 39.850 175.325 ;
        RECT 39.650 174.840 39.790 175.005 ;
        RECT 39.580 174.470 39.860 174.840 ;
        RECT 39.590 174.325 39.850 174.470 ;
        RECT 37.350 173.225 37.950 173.365 ;
        RECT 37.350 172.265 37.490 173.225 ;
        RECT 39.650 172.265 39.790 174.325 ;
        RECT 37.290 171.945 37.550 172.265 ;
        RECT 39.590 171.945 39.850 172.265 ;
        RECT 41.430 171.265 41.690 171.585 ;
        RECT 37.470 170.730 39.010 171.100 ;
        RECT 40.970 168.885 41.230 169.205 ;
        RECT 39.590 168.545 39.850 168.865 ;
        RECT 39.130 167.525 39.390 167.845 ;
        RECT 37.470 165.290 39.010 165.660 ;
        RECT 38.210 163.785 38.470 164.105 ;
        RECT 37.750 163.105 38.010 163.425 ;
        RECT 37.810 161.725 37.950 163.105 ;
        RECT 38.270 162.405 38.410 163.785 ;
        RECT 38.210 162.085 38.470 162.405 ;
        RECT 37.750 161.405 38.010 161.725 ;
        RECT 39.190 161.385 39.330 167.525 ;
        RECT 39.650 166.825 39.790 168.545 ;
        RECT 40.050 167.185 40.310 167.505 ;
        RECT 39.590 166.505 39.850 166.825 ;
        RECT 38.670 161.240 38.930 161.385 ;
        RECT 36.820 160.870 37.100 161.240 ;
        RECT 38.660 160.870 38.940 161.240 ;
        RECT 39.130 161.065 39.390 161.385 ;
        RECT 36.890 154.245 37.030 160.870 ;
        RECT 37.470 159.850 39.010 160.220 ;
        RECT 39.130 157.665 39.390 157.985 ;
        RECT 37.470 154.410 39.010 154.780 ;
        RECT 36.830 153.925 37.090 154.245 ;
        RECT 38.210 153.925 38.470 154.245 ;
        RECT 36.830 153.245 37.090 153.565 ;
        RECT 37.750 153.245 38.010 153.565 ;
        RECT 36.890 148.125 37.030 153.245 ;
        RECT 37.290 151.205 37.550 151.525 ;
        RECT 37.350 150.505 37.490 151.205 ;
        RECT 37.290 150.185 37.550 150.505 ;
        RECT 37.810 150.165 37.950 153.245 ;
        RECT 38.270 151.185 38.410 153.925 ;
        RECT 38.210 150.865 38.470 151.185 ;
        RECT 38.270 150.505 38.410 150.865 ;
        RECT 38.210 150.185 38.470 150.505 ;
        RECT 37.750 149.845 38.010 150.165 ;
        RECT 37.470 148.970 39.010 149.340 ;
        RECT 38.210 148.485 38.470 148.805 ;
        RECT 36.830 148.035 37.090 148.125 ;
        RECT 36.830 147.895 37.950 148.035 ;
        RECT 36.830 147.805 37.090 147.895 ;
        RECT 36.830 146.785 37.090 147.105 ;
        RECT 36.890 142.685 37.030 146.785 ;
        RECT 37.280 146.590 37.560 146.960 ;
        RECT 37.350 145.065 37.490 146.590 ;
        RECT 37.810 145.745 37.950 147.895 ;
        RECT 37.750 145.425 38.010 145.745 ;
        RECT 38.270 145.065 38.410 148.485 ;
        RECT 37.290 144.745 37.550 145.065 ;
        RECT 38.210 144.745 38.470 145.065 ;
        RECT 37.470 143.530 39.010 143.900 ;
        RECT 36.370 142.365 36.630 142.685 ;
        RECT 36.830 142.365 37.090 142.685 ;
        RECT 36.830 140.325 37.090 140.645 ;
        RECT 35.910 139.645 36.170 139.965 ;
        RECT 36.890 137.925 37.030 140.325 ;
        RECT 37.470 138.090 39.010 138.460 ;
        RECT 36.830 137.605 37.090 137.925 ;
        RECT 35.910 136.925 36.170 137.245 ;
        RECT 37.750 136.925 38.010 137.245 ;
        RECT 35.970 133.505 36.110 136.925 ;
        RECT 37.810 134.865 37.950 136.925 ;
        RECT 36.370 134.545 36.630 134.865 ;
        RECT 37.750 134.545 38.010 134.865 ;
        RECT 35.910 133.185 36.170 133.505 ;
        RECT 36.430 128.745 36.570 134.545 ;
        RECT 39.190 134.185 39.330 157.665 ;
        RECT 39.650 155.125 39.790 166.505 ;
        RECT 40.110 164.445 40.250 167.185 ;
        RECT 40.510 166.165 40.770 166.485 ;
        RECT 40.570 164.445 40.710 166.165 ;
        RECT 40.050 164.125 40.310 164.445 ;
        RECT 40.510 164.125 40.770 164.445 ;
        RECT 40.110 161.385 40.250 164.125 ;
        RECT 40.050 161.065 40.310 161.385 ;
        RECT 40.050 160.385 40.310 160.705 ;
        RECT 40.110 159.345 40.250 160.385 ;
        RECT 40.050 159.025 40.310 159.345 ;
        RECT 40.050 158.405 40.310 158.665 ;
        RECT 41.030 158.405 41.170 168.885 ;
        RECT 41.490 159.005 41.630 171.265 ;
        RECT 41.950 169.885 42.090 175.345 ;
        RECT 42.870 175.325 43.010 187.585 ;
        RECT 43.270 182.825 43.530 183.145 ;
        RECT 43.330 181.105 43.470 182.825 ;
        RECT 43.270 180.785 43.530 181.105 ;
        RECT 42.810 175.005 43.070 175.325 ;
        RECT 42.810 172.625 43.070 172.945 ;
        RECT 42.870 171.925 43.010 172.625 ;
        RECT 42.810 171.605 43.070 171.925 ;
        RECT 42.870 169.885 43.010 171.605 ;
        RECT 43.790 169.885 43.930 192.005 ;
        RECT 44.250 188.245 44.390 193.705 ;
        RECT 44.710 191.305 44.850 196.425 ;
        RECT 46.090 195.045 46.230 199.145 ;
        RECT 47.410 198.465 47.670 198.785 ;
        RECT 47.470 197.425 47.610 198.465 ;
        RECT 47.410 197.105 47.670 197.425 ;
        RECT 46.030 194.725 46.290 195.045 ;
        RECT 47.930 191.985 48.070 199.145 ;
        RECT 50.170 196.765 50.430 197.085 ;
        RECT 50.230 195.045 50.370 196.765 ;
        RECT 52.530 196.745 52.670 199.145 ;
        RECT 57.530 198.805 57.790 199.125 ;
        RECT 57.590 197.765 57.730 198.805 ;
        RECT 57.530 197.445 57.790 197.765 ;
        RECT 56.610 196.765 56.870 197.085 ;
        RECT 52.470 196.425 52.730 196.745 ;
        RECT 50.865 195.210 52.405 195.580 ;
        RECT 50.170 194.725 50.430 195.045 ;
        RECT 48.330 194.045 48.590 194.365 ;
        RECT 46.030 191.665 46.290 191.985 ;
        RECT 47.870 191.665 48.130 191.985 ;
        RECT 44.650 190.985 44.910 191.305 ;
        RECT 44.190 187.925 44.450 188.245 ;
        RECT 44.250 172.265 44.390 187.925 ;
        RECT 44.710 185.185 44.850 190.985 ;
        RECT 46.090 188.585 46.230 191.665 ;
        RECT 47.410 191.325 47.670 191.645 ;
        RECT 46.030 188.265 46.290 188.585 ;
        RECT 45.570 187.585 45.830 187.905 ;
        RECT 44.650 184.865 44.910 185.185 ;
        RECT 44.710 183.145 44.850 184.865 ;
        RECT 44.650 182.825 44.910 183.145 ;
        RECT 44.710 180.425 44.850 182.825 ;
        RECT 45.630 182.805 45.770 187.585 ;
        RECT 46.090 183.825 46.230 188.265 ;
        RECT 47.470 188.155 47.610 191.325 ;
        RECT 48.390 191.305 48.530 194.045 ;
        RECT 48.790 193.705 49.050 194.025 ;
        RECT 48.850 192.325 48.990 193.705 ;
        RECT 48.790 192.005 49.050 192.325 ;
        RECT 56.670 191.645 56.810 196.765 ;
        RECT 56.610 191.325 56.870 191.645 ;
        RECT 48.330 190.985 48.590 191.305 ;
        RECT 50.170 190.985 50.430 191.305 ;
        RECT 48.390 188.925 48.530 190.985 ;
        RECT 49.710 190.305 49.970 190.625 ;
        RECT 48.330 188.605 48.590 188.925 ;
        RECT 47.870 188.155 48.130 188.245 ;
        RECT 47.470 188.015 48.130 188.155 ;
        RECT 47.870 187.925 48.130 188.015 ;
        RECT 47.930 186.885 48.070 187.925 ;
        RECT 47.870 186.565 48.130 186.885 ;
        RECT 48.390 185.865 48.530 188.605 ;
        RECT 49.770 188.245 49.910 190.305 ;
        RECT 49.710 187.925 49.970 188.245 ;
        RECT 50.230 186.885 50.370 190.985 ;
        RECT 53.850 190.305 54.110 190.625 ;
        RECT 50.865 189.770 52.405 190.140 ;
        RECT 53.910 188.925 54.050 190.305 ;
        RECT 56.670 188.925 56.810 191.325 ;
        RECT 53.850 188.605 54.110 188.925 ;
        RECT 56.610 188.605 56.870 188.925 ;
        RECT 55.690 188.265 55.950 188.585 ;
        RECT 50.170 186.565 50.430 186.885 ;
        RECT 48.790 186.225 49.050 186.545 ;
        RECT 48.330 185.545 48.590 185.865 ;
        RECT 48.390 184.165 48.530 185.545 ;
        RECT 48.330 183.845 48.590 184.165 ;
        RECT 46.030 183.505 46.290 183.825 ;
        RECT 45.110 182.485 45.370 182.805 ;
        RECT 45.570 182.485 45.830 182.805 ;
        RECT 45.170 181.445 45.310 182.485 ;
        RECT 45.110 181.125 45.370 181.445 ;
        RECT 47.410 181.125 47.670 181.445 ;
        RECT 44.650 180.105 44.910 180.425 ;
        RECT 44.190 171.945 44.450 172.265 ;
        RECT 41.890 169.565 42.150 169.885 ;
        RECT 42.810 169.565 43.070 169.885 ;
        RECT 43.730 169.565 43.990 169.885 ;
        RECT 44.190 169.565 44.450 169.885 ;
        RECT 44.250 167.505 44.390 169.565 ;
        RECT 44.710 169.545 44.850 180.105 ;
        RECT 47.470 177.705 47.610 181.125 ;
        RECT 48.390 180.425 48.530 183.845 ;
        RECT 48.850 182.465 48.990 186.225 ;
        RECT 50.170 185.885 50.430 186.205 ;
        RECT 49.250 183.505 49.510 183.825 ;
        RECT 48.790 182.145 49.050 182.465 ;
        RECT 48.850 180.425 48.990 182.145 ;
        RECT 48.330 180.105 48.590 180.425 ;
        RECT 48.790 180.105 49.050 180.425 ;
        RECT 48.390 178.725 48.530 180.105 ;
        RECT 48.330 178.405 48.590 178.725 ;
        RECT 47.870 178.065 48.130 178.385 ;
        RECT 47.410 177.385 47.670 177.705 ;
        RECT 45.110 176.705 45.370 177.025 ;
        RECT 47.410 176.705 47.670 177.025 ;
        RECT 44.650 169.225 44.910 169.545 ;
        RECT 43.270 167.185 43.530 167.505 ;
        RECT 44.190 167.185 44.450 167.505 ;
        RECT 41.880 164.270 42.160 164.640 ;
        RECT 43.330 164.355 43.470 167.185 ;
        RECT 43.730 165.035 43.990 165.125 ;
        RECT 43.730 164.895 44.850 165.035 ;
        RECT 43.730 164.805 43.990 164.895 ;
        RECT 44.710 164.445 44.850 164.895 ;
        RECT 43.730 164.355 43.990 164.445 ;
        RECT 41.890 164.125 42.150 164.270 ;
        RECT 43.330 164.215 43.990 164.355 ;
        RECT 43.730 164.125 43.990 164.215 ;
        RECT 44.650 164.125 44.910 164.445 ;
        RECT 41.950 161.385 42.090 164.125 ;
        RECT 44.190 163.445 44.450 163.765 ;
        RECT 43.270 163.105 43.530 163.425 ;
        RECT 42.350 161.920 42.610 162.065 ;
        RECT 42.340 161.550 42.620 161.920 ;
        RECT 41.890 161.065 42.150 161.385 ;
        RECT 42.350 160.385 42.610 160.705 ;
        RECT 42.810 160.385 43.070 160.705 ;
        RECT 42.410 159.005 42.550 160.385 ;
        RECT 42.870 159.345 43.010 160.385 ;
        RECT 43.330 159.685 43.470 163.105 ;
        RECT 44.250 161.385 44.390 163.445 ;
        RECT 44.190 161.125 44.450 161.385 ;
        RECT 44.190 161.065 44.850 161.125 ;
        RECT 44.250 160.985 44.850 161.065 ;
        RECT 43.270 159.365 43.530 159.685 ;
        RECT 42.810 159.025 43.070 159.345 ;
        RECT 44.710 159.005 44.850 160.985 ;
        RECT 41.430 158.685 41.690 159.005 ;
        RECT 42.350 158.685 42.610 159.005 ;
        RECT 43.730 158.685 43.990 159.005 ;
        RECT 44.190 158.685 44.450 159.005 ;
        RECT 44.650 158.685 44.910 159.005 ;
        RECT 40.050 158.345 41.170 158.405 ;
        RECT 42.810 158.345 43.070 158.665 ;
        RECT 40.110 158.265 41.170 158.345 ;
        RECT 39.650 154.985 40.250 155.125 ;
        RECT 40.110 153.565 40.250 154.985 ;
        RECT 40.050 153.245 40.310 153.565 ;
        RECT 40.970 152.905 41.230 153.225 ;
        RECT 42.350 152.905 42.610 153.225 ;
        RECT 41.030 150.845 41.170 152.905 ;
        RECT 40.970 150.525 41.230 150.845 ;
        RECT 39.590 149.845 39.850 150.165 ;
        RECT 39.650 147.785 39.790 149.845 ;
        RECT 39.590 147.465 39.850 147.785 ;
        RECT 39.650 145.405 39.790 147.465 ;
        RECT 40.510 146.785 40.770 147.105 ;
        RECT 39.590 145.085 39.850 145.405 ;
        RECT 40.570 143.025 40.710 146.785 ;
        RECT 40.510 142.705 40.770 143.025 ;
        RECT 41.030 135.205 41.170 150.525 ;
        RECT 41.890 138.625 42.150 138.945 ;
        RECT 40.970 134.885 41.230 135.205 ;
        RECT 40.510 134.205 40.770 134.525 ;
        RECT 39.130 133.865 39.390 134.185 ;
        RECT 36.830 133.525 37.090 133.845 ;
        RECT 36.370 128.425 36.630 128.745 ;
        RECT 36.890 128.065 37.030 133.525 ;
        RECT 39.130 133.185 39.390 133.505 ;
        RECT 37.470 132.650 39.010 133.020 ;
        RECT 39.190 131.805 39.330 133.185 ;
        RECT 39.130 131.485 39.390 131.805 ;
        RECT 40.570 128.745 40.710 134.205 ;
        RECT 40.510 128.425 40.770 128.745 ;
        RECT 39.130 128.085 39.390 128.405 ;
        RECT 36.830 127.745 37.090 128.065 ;
        RECT 36.890 127.045 37.030 127.745 ;
        RECT 37.470 127.210 39.010 127.580 ;
        RECT 36.830 126.725 37.090 127.045 ;
        RECT 37.750 126.385 38.010 126.705 ;
        RECT 37.810 124.325 37.950 126.385 ;
        RECT 37.750 124.005 38.010 124.325 ;
        RECT 37.470 121.770 39.010 122.140 ;
        RECT 39.190 120.925 39.330 128.085 ;
        RECT 40.970 127.745 41.230 128.065 ;
        RECT 40.510 125.705 40.770 126.025 ;
        RECT 39.130 120.605 39.390 120.925 ;
        RECT 35.450 118.565 35.710 118.885 ;
        RECT 34.130 118.205 34.730 118.285 ;
        RECT 40.570 118.205 40.710 125.705 ;
        RECT 41.030 123.305 41.170 127.745 ;
        RECT 41.430 126.045 41.690 126.365 ;
        RECT 41.490 124.325 41.630 126.045 ;
        RECT 41.430 124.005 41.690 124.325 ;
        RECT 40.970 122.985 41.230 123.305 ;
        RECT 34.070 118.145 34.730 118.205 ;
        RECT 34.070 117.885 34.330 118.145 ;
        RECT 27.170 115.165 27.430 115.485 ;
        RECT 28.090 115.165 28.350 115.485 ;
        RECT 29.930 115.165 30.190 115.485 ;
        RECT 32.230 115.165 32.490 115.485 ;
        RECT 24.075 113.610 25.615 113.980 ;
        RECT 27.230 112.765 27.370 115.165 ;
        RECT 29.470 114.145 29.730 114.465 ;
        RECT 27.170 112.445 27.430 112.765 ;
        RECT 25.330 111.765 25.590 112.085 ;
        RECT 25.390 110.725 25.530 111.765 ;
        RECT 23.490 110.405 23.750 110.725 ;
        RECT 25.330 110.405 25.590 110.725 ;
        RECT 23.090 109.985 23.690 110.125 ;
        RECT 23.550 106.285 23.690 109.985 ;
        RECT 26.710 109.955 26.970 110.045 ;
        RECT 27.230 109.955 27.370 112.445 ;
        RECT 29.530 112.085 29.670 114.145 ;
        RECT 29.010 111.765 29.270 112.085 ;
        RECT 29.470 111.765 29.730 112.085 ;
        RECT 26.710 109.815 27.370 109.955 ;
        RECT 26.710 109.725 26.970 109.815 ;
        RECT 24.075 108.170 25.615 108.540 ;
        RECT 29.070 106.285 29.210 111.765 ;
        RECT 29.990 111.745 30.130 115.165 ;
        RECT 31.310 114.145 31.570 114.465 ;
        RECT 31.370 113.105 31.510 114.145 ;
        RECT 31.310 112.785 31.570 113.105 ;
        RECT 29.930 111.425 30.190 111.745 ;
        RECT 29.990 110.045 30.130 111.425 ;
        RECT 29.930 109.725 30.190 110.045 ;
        RECT 34.590 106.285 34.730 118.145 ;
        RECT 39.130 117.885 39.390 118.205 ;
        RECT 40.510 117.885 40.770 118.205 ;
        RECT 37.470 116.330 39.010 116.700 ;
        RECT 38.210 115.505 38.470 115.825 ;
        RECT 38.270 113.445 38.410 115.505 ;
        RECT 38.210 113.125 38.470 113.445 ;
        RECT 39.190 113.105 39.330 117.885 ;
        RECT 41.950 117.865 42.090 138.625 ;
        RECT 41.890 117.545 42.150 117.865 ;
        RECT 41.430 116.865 41.690 117.185 ;
        RECT 41.490 115.825 41.630 116.865 ;
        RECT 41.430 115.505 41.690 115.825 ;
        RECT 39.590 115.055 39.850 115.145 ;
        RECT 39.590 114.915 40.250 115.055 ;
        RECT 39.590 114.825 39.850 114.915 ;
        RECT 39.130 112.785 39.390 113.105 ;
        RECT 39.130 112.105 39.390 112.425 ;
        RECT 37.470 110.890 39.010 111.260 ;
        RECT 39.190 110.045 39.330 112.105 ;
        RECT 39.130 109.725 39.390 110.045 ;
        RECT 40.110 106.285 40.250 114.915 ;
        RECT 42.410 112.425 42.550 152.905 ;
        RECT 42.870 139.965 43.010 158.345 ;
        RECT 43.270 157.665 43.530 157.985 ;
        RECT 42.810 139.645 43.070 139.965 ;
        RECT 43.330 134.185 43.470 157.665 ;
        RECT 43.790 153.565 43.930 158.685 ;
        RECT 44.250 156.965 44.390 158.685 ;
        RECT 44.190 156.645 44.450 156.965 ;
        RECT 44.650 154.945 44.910 155.265 ;
        RECT 43.730 153.245 43.990 153.565 ;
        RECT 44.710 153.225 44.850 154.945 ;
        RECT 44.650 152.905 44.910 153.225 ;
        RECT 44.650 152.225 44.910 152.545 ;
        RECT 44.710 150.165 44.850 152.225 ;
        RECT 44.650 149.845 44.910 150.165 ;
        RECT 44.710 148.465 44.850 149.845 ;
        RECT 44.650 148.145 44.910 148.465 ;
        RECT 45.170 147.525 45.310 176.705 ;
        RECT 46.030 175.915 46.290 176.005 ;
        RECT 45.630 175.775 46.290 175.915 ;
        RECT 45.630 155.945 45.770 175.775 ;
        RECT 46.030 175.685 46.290 175.775 ;
        RECT 47.470 175.325 47.610 176.705 ;
        RECT 47.930 175.325 48.070 178.065 ;
        RECT 48.850 175.325 48.990 180.105 ;
        RECT 47.410 175.005 47.670 175.325 ;
        RECT 47.870 175.005 48.130 175.325 ;
        RECT 48.790 175.005 49.050 175.325 ;
        RECT 46.950 174.665 47.210 174.985 ;
        RECT 46.030 174.325 46.290 174.645 ;
        RECT 46.090 172.265 46.230 174.325 ;
        RECT 46.030 171.945 46.290 172.265 ;
        RECT 46.030 169.225 46.290 169.545 ;
        RECT 46.090 165.125 46.230 169.225 ;
        RECT 46.030 164.805 46.290 165.125 ;
        RECT 46.490 164.640 46.750 164.785 ;
        RECT 46.480 164.525 46.760 164.640 ;
        RECT 46.090 164.385 46.760 164.525 ;
        RECT 46.090 159.005 46.230 164.385 ;
        RECT 46.480 164.270 46.760 164.385 ;
        RECT 46.490 163.105 46.750 163.425 ;
        RECT 46.030 158.685 46.290 159.005 ;
        RECT 46.550 156.285 46.690 163.105 ;
        RECT 47.010 159.005 47.150 174.665 ;
        RECT 47.470 171.585 47.610 175.005 ;
        RECT 49.310 172.265 49.450 183.505 ;
        RECT 50.230 181.445 50.370 185.885 ;
        RECT 53.390 184.865 53.650 185.185 ;
        RECT 50.865 184.330 52.405 184.700 ;
        RECT 53.450 183.485 53.590 184.865 ;
        RECT 53.390 183.165 53.650 183.485 ;
        RECT 55.750 183.145 55.890 188.265 ;
        RECT 55.690 182.825 55.950 183.145 ;
        RECT 50.170 181.125 50.430 181.445 ;
        RECT 49.710 180.785 49.970 181.105 ;
        RECT 49.770 178.385 49.910 180.785 ;
        RECT 58.050 180.765 58.190 203.905 ;
        RECT 58.970 200.145 59.110 207.305 ;
        RECT 60.750 206.625 61.010 206.945 ;
        RECT 59.370 204.925 59.630 205.245 ;
        RECT 59.430 201.845 59.570 204.925 ;
        RECT 59.830 204.585 60.090 204.905 ;
        RECT 59.890 202.865 60.030 204.585 ;
        RECT 60.810 204.565 60.950 206.625 ;
        RECT 60.750 204.245 61.010 204.565 ;
        RECT 60.810 203.205 60.950 204.245 ;
        RECT 61.210 203.905 61.470 204.225 ;
        RECT 60.750 202.885 61.010 203.205 ;
        RECT 59.830 202.545 60.090 202.865 ;
        RECT 59.370 201.525 59.630 201.845 ;
        RECT 58.910 199.825 59.170 200.145 ;
        RECT 58.450 198.465 58.710 198.785 ;
        RECT 58.510 197.765 58.650 198.465 ;
        RECT 58.450 197.445 58.710 197.765 ;
        RECT 58.970 197.085 59.110 199.825 ;
        RECT 59.430 197.765 59.570 201.525 ;
        RECT 59.890 199.885 60.030 202.545 ;
        RECT 61.270 202.525 61.410 203.905 ;
        RECT 61.730 203.285 61.870 207.305 ;
        RECT 62.130 205.605 62.390 205.925 ;
        RECT 62.190 204.645 62.330 205.605 ;
        RECT 62.650 205.585 62.790 209.685 ;
        RECT 63.570 207.625 63.710 210.025 ;
        RECT 68.570 209.345 68.830 209.665 ;
        RECT 64.260 208.810 65.800 209.180 ;
        RECT 68.630 208.305 68.770 209.345 ;
        RECT 68.570 207.985 68.830 208.305 ;
        RECT 63.510 207.305 63.770 207.625 ;
        RECT 62.590 205.265 62.850 205.585 ;
        RECT 62.190 204.505 63.250 204.645 ;
        RECT 62.590 203.905 62.850 204.225 ;
        RECT 61.730 203.205 62.330 203.285 ;
        RECT 61.730 203.145 62.390 203.205 ;
        RECT 62.130 202.885 62.390 203.145 ;
        RECT 61.670 202.545 61.930 202.865 ;
        RECT 61.210 202.205 61.470 202.525 ;
        RECT 60.750 201.185 61.010 201.505 ;
        RECT 59.890 199.745 60.490 199.885 ;
        RECT 60.350 199.465 60.490 199.745 ;
        RECT 60.290 199.145 60.550 199.465 ;
        RECT 59.370 197.445 59.630 197.765 ;
        RECT 60.350 197.085 60.490 199.145 ;
        RECT 60.810 197.085 60.950 201.185 ;
        RECT 61.730 197.675 61.870 202.545 ;
        RECT 62.130 201.185 62.390 201.505 ;
        RECT 61.270 197.535 61.870 197.675 ;
        RECT 61.270 197.085 61.410 197.535 ;
        RECT 58.910 196.765 59.170 197.085 ;
        RECT 60.290 196.765 60.550 197.085 ;
        RECT 60.750 196.765 61.010 197.085 ;
        RECT 61.210 196.765 61.470 197.085 ;
        RECT 61.670 196.765 61.930 197.085 ;
        RECT 60.810 194.025 60.950 196.765 ;
        RECT 60.290 193.705 60.550 194.025 ;
        RECT 60.750 193.705 61.010 194.025 ;
        RECT 60.350 190.625 60.490 193.705 ;
        RECT 61.270 193.685 61.410 196.765 ;
        RECT 61.730 196.065 61.870 196.765 ;
        RECT 61.670 195.745 61.930 196.065 ;
        RECT 61.210 193.365 61.470 193.685 ;
        RECT 60.290 190.305 60.550 190.625 ;
        RECT 61.730 186.885 61.870 195.745 ;
        RECT 61.670 186.565 61.930 186.885 ;
        RECT 60.750 185.885 61.010 186.205 ;
        RECT 59.830 184.865 60.090 185.185 ;
        RECT 57.990 180.445 58.250 180.765 ;
        RECT 57.530 179.765 57.790 180.085 ;
        RECT 50.865 178.890 52.405 179.260 ;
        RECT 57.590 178.725 57.730 179.765 ;
        RECT 57.530 178.405 57.790 178.725 ;
        RECT 49.710 178.065 49.970 178.385 ;
        RECT 58.050 178.045 58.190 180.445 ;
        RECT 59.370 178.065 59.630 178.385 ;
        RECT 57.990 177.725 58.250 178.045 ;
        RECT 49.710 177.385 49.970 177.705 ;
        RECT 58.910 177.385 59.170 177.705 ;
        RECT 49.770 174.840 49.910 177.385 ;
        RECT 55.690 176.705 55.950 177.025 ;
        RECT 52.930 175.005 53.190 175.325 ;
        RECT 49.700 174.470 49.980 174.840 ;
        RECT 49.770 172.945 49.910 174.470 ;
        RECT 50.865 173.450 52.405 173.820 ;
        RECT 49.710 172.625 49.970 172.945 ;
        RECT 49.250 171.945 49.510 172.265 ;
        RECT 47.410 171.265 47.670 171.585 ;
        RECT 49.310 169.965 49.450 171.945 ;
        RECT 52.990 171.925 53.130 175.005 ;
        RECT 55.750 173.285 55.890 176.705 ;
        RECT 58.440 175.150 58.720 175.520 ;
        RECT 55.690 172.965 55.950 173.285 ;
        RECT 57.990 172.965 58.250 173.285 ;
        RECT 52.930 171.605 53.190 171.925 ;
        RECT 55.750 171.585 55.890 172.965 ;
        RECT 58.050 171.925 58.190 172.965 ;
        RECT 57.990 171.605 58.250 171.925 ;
        RECT 49.710 171.265 49.970 171.585 ;
        RECT 55.690 171.265 55.950 171.585 ;
        RECT 49.770 170.225 49.910 171.265 ;
        RECT 48.850 169.825 49.450 169.965 ;
        RECT 49.710 169.905 49.970 170.225 ;
        RECT 48.330 166.845 48.590 167.165 ;
        RECT 47.410 163.105 47.670 163.425 ;
        RECT 47.470 161.385 47.610 163.105 ;
        RECT 48.390 161.385 48.530 166.845 ;
        RECT 48.850 166.485 48.990 169.825 ;
        RECT 49.710 169.225 49.970 169.545 ;
        RECT 48.790 166.165 49.050 166.485 ;
        RECT 47.410 161.065 47.670 161.385 ;
        RECT 48.330 161.065 48.590 161.385 ;
        RECT 46.950 158.685 47.210 159.005 ;
        RECT 46.950 157.840 47.210 157.985 ;
        RECT 46.940 157.470 47.220 157.840 ;
        RECT 47.870 157.665 48.130 157.985 ;
        RECT 46.950 156.645 47.210 156.965 ;
        RECT 46.490 155.965 46.750 156.285 ;
        RECT 45.570 155.625 45.830 155.945 ;
        RECT 45.570 152.225 45.830 152.545 ;
        RECT 45.630 150.505 45.770 152.225 ;
        RECT 46.490 151.205 46.750 151.525 ;
        RECT 45.570 150.185 45.830 150.505 ;
        RECT 45.630 148.805 45.770 150.185 ;
        RECT 45.570 148.485 45.830 148.805 ;
        RECT 44.710 147.385 45.310 147.525 ;
        RECT 44.190 144.065 44.450 144.385 ;
        RECT 44.250 143.365 44.390 144.065 ;
        RECT 44.190 143.045 44.450 143.365 ;
        RECT 43.730 141.345 43.990 141.665 ;
        RECT 43.790 139.625 43.930 141.345 ;
        RECT 44.710 139.625 44.850 147.385 ;
        RECT 45.630 145.065 45.770 148.485 ;
        RECT 46.550 147.445 46.690 151.205 ;
        RECT 46.490 147.125 46.750 147.445 ;
        RECT 46.550 145.065 46.690 147.125 ;
        RECT 45.570 144.745 45.830 145.065 ;
        RECT 46.490 144.745 46.750 145.065 ;
        RECT 45.630 142.685 45.770 144.745 ;
        RECT 46.550 143.025 46.690 144.745 ;
        RECT 46.490 142.705 46.750 143.025 ;
        RECT 45.570 142.365 45.830 142.685 ;
        RECT 45.110 140.325 45.370 140.645 ;
        RECT 43.730 139.305 43.990 139.625 ;
        RECT 44.650 139.305 44.910 139.625 ;
        RECT 43.730 138.625 43.990 138.945 ;
        RECT 43.270 133.865 43.530 134.185 ;
        RECT 43.270 128.085 43.530 128.405 ;
        RECT 43.330 124.325 43.470 128.085 ;
        RECT 43.270 124.005 43.530 124.325 ;
        RECT 43.790 117.865 43.930 138.625 ;
        RECT 45.170 134.185 45.310 140.325 ;
        RECT 46.550 139.965 46.690 142.705 ;
        RECT 46.490 139.645 46.750 139.965 ;
        RECT 44.190 133.865 44.450 134.185 ;
        RECT 44.650 133.865 44.910 134.185 ;
        RECT 45.110 133.865 45.370 134.185 ;
        RECT 44.250 126.365 44.390 133.865 ;
        RECT 44.710 132.145 44.850 133.865 ;
        RECT 47.010 132.485 47.150 156.645 ;
        RECT 47.410 149.505 47.670 149.825 ;
        RECT 47.470 147.105 47.610 149.505 ;
        RECT 47.410 146.785 47.670 147.105 ;
        RECT 47.470 145.065 47.610 146.785 ;
        RECT 47.410 144.745 47.670 145.065 ;
        RECT 47.470 143.365 47.610 144.745 ;
        RECT 47.410 143.045 47.670 143.365 ;
        RECT 47.410 142.365 47.670 142.685 ;
        RECT 47.470 139.625 47.610 142.365 ;
        RECT 47.410 139.480 47.670 139.625 ;
        RECT 47.400 139.110 47.680 139.480 ;
        RECT 47.410 134.205 47.670 134.525 ;
        RECT 46.950 132.165 47.210 132.485 ;
        RECT 44.650 131.825 44.910 132.145 ;
        RECT 45.570 128.765 45.830 129.085 ;
        RECT 44.190 126.045 44.450 126.365 ;
        RECT 44.250 121.605 44.390 126.045 ;
        RECT 45.630 125.345 45.770 128.765 ;
        RECT 47.470 126.025 47.610 134.205 ;
        RECT 47.930 133.845 48.070 157.665 ;
        RECT 48.390 156.285 48.530 161.065 ;
        RECT 48.850 157.725 48.990 166.165 ;
        RECT 49.770 166.145 49.910 169.225 ;
        RECT 51.090 168.925 51.350 169.205 ;
        RECT 50.230 168.885 51.350 168.925 ;
        RECT 50.230 168.785 51.290 168.885 ;
        RECT 50.230 166.825 50.370 168.785 ;
        RECT 53.850 168.545 54.110 168.865 ;
        RECT 55.230 168.545 55.490 168.865 ;
        RECT 50.865 168.010 52.405 168.380 ;
        RECT 50.170 166.505 50.430 166.825 ;
        RECT 52.930 166.505 53.190 166.825 ;
        RECT 49.250 165.825 49.510 166.145 ;
        RECT 49.710 165.825 49.970 166.145 ;
        RECT 49.310 164.445 49.450 165.825 ;
        RECT 49.250 164.125 49.510 164.445 ;
        RECT 49.250 163.105 49.510 163.425 ;
        RECT 49.310 161.385 49.450 163.105 ;
        RECT 49.250 161.065 49.510 161.385 ;
        RECT 49.310 158.325 49.450 161.065 ;
        RECT 49.250 158.005 49.510 158.325 ;
        RECT 48.850 157.585 49.450 157.725 ;
        RECT 48.330 155.965 48.590 156.285 ;
        RECT 48.390 151.185 48.530 155.965 ;
        RECT 49.310 155.945 49.450 157.585 ;
        RECT 49.770 155.945 49.910 165.825 ;
        RECT 52.990 164.105 53.130 166.505 ;
        RECT 53.910 166.145 54.050 168.545 ;
        RECT 54.310 166.845 54.570 167.165 ;
        RECT 53.850 165.825 54.110 166.145 ;
        RECT 52.930 163.785 53.190 164.105 ;
        RECT 50.865 162.570 52.405 162.940 ;
        RECT 50.160 161.550 50.440 161.920 ;
        RECT 50.170 161.405 50.430 161.550 ;
        RECT 50.230 159.685 50.370 161.405 ;
        RECT 52.990 161.385 53.130 163.785 ;
        RECT 52.010 161.240 52.270 161.385 ;
        RECT 52.000 160.870 52.280 161.240 ;
        RECT 52.470 161.065 52.730 161.385 ;
        RECT 52.930 161.065 53.190 161.385 ;
        RECT 50.170 159.365 50.430 159.685 ;
        RECT 52.530 158.325 52.670 161.065 ;
        RECT 52.470 158.005 52.730 158.325 ;
        RECT 50.865 157.130 52.405 157.500 ;
        RECT 49.250 155.625 49.510 155.945 ;
        RECT 49.710 155.625 49.970 155.945 ;
        RECT 48.790 154.945 49.050 155.265 ;
        RECT 48.850 153.905 48.990 154.945 ;
        RECT 48.790 153.585 49.050 153.905 ;
        RECT 48.330 150.865 48.590 151.185 ;
        RECT 48.390 142.255 48.530 150.865 ;
        RECT 48.790 150.185 49.050 150.505 ;
        RECT 48.850 147.785 48.990 150.185 ;
        RECT 48.790 147.465 49.050 147.785 ;
        RECT 48.850 145.065 48.990 147.465 ;
        RECT 49.310 147.105 49.450 155.625 ;
        RECT 49.770 150.845 49.910 155.625 ;
        RECT 50.170 154.945 50.430 155.265 ;
        RECT 49.710 150.525 49.970 150.845 ;
        RECT 50.230 150.165 50.370 154.945 ;
        RECT 53.390 153.925 53.650 154.245 ;
        RECT 52.930 153.475 53.190 153.565 ;
        RECT 53.450 153.475 53.590 153.925 ;
        RECT 53.910 153.565 54.050 165.825 ;
        RECT 54.370 162.405 54.510 166.845 ;
        RECT 55.290 164.785 55.430 168.545 ;
        RECT 55.230 164.465 55.490 164.785 ;
        RECT 58.050 164.445 58.190 171.605 ;
        RECT 54.770 164.125 55.030 164.445 ;
        RECT 56.610 164.125 56.870 164.445 ;
        RECT 57.990 164.125 58.250 164.445 ;
        RECT 54.310 162.085 54.570 162.405 ;
        RECT 54.310 161.405 54.570 161.725 ;
        RECT 54.370 159.345 54.510 161.405 ;
        RECT 54.830 161.240 54.970 164.125 ;
        RECT 56.150 161.295 56.410 161.385 ;
        RECT 56.670 161.295 56.810 164.125 ;
        RECT 54.760 160.870 55.040 161.240 ;
        RECT 56.150 161.155 56.810 161.295 ;
        RECT 56.150 161.065 56.410 161.155 ;
        RECT 57.530 161.065 57.790 161.385 ;
        RECT 54.770 160.725 55.030 160.870 ;
        RECT 54.310 159.025 54.570 159.345 ;
        RECT 54.830 155.945 54.970 160.725 ;
        RECT 55.690 160.385 55.950 160.705 ;
        RECT 55.750 155.945 55.890 160.385 ;
        RECT 56.210 158.325 56.350 161.065 ;
        RECT 57.590 159.685 57.730 161.065 ;
        RECT 57.530 159.365 57.790 159.685 ;
        RECT 56.150 158.005 56.410 158.325 ;
        RECT 56.210 156.285 56.350 158.005 ;
        RECT 56.150 155.965 56.410 156.285 ;
        RECT 57.590 155.945 57.730 159.365 ;
        RECT 58.510 157.840 58.650 175.150 ;
        RECT 58.970 174.305 59.110 177.385 ;
        RECT 59.430 175.665 59.570 178.065 ;
        RECT 59.370 175.345 59.630 175.665 ;
        RECT 59.890 175.325 60.030 184.865 ;
        RECT 60.810 183.485 60.950 185.885 ;
        RECT 61.210 183.845 61.470 184.165 ;
        RECT 61.270 183.485 61.410 183.845 ;
        RECT 60.750 183.165 61.010 183.485 ;
        RECT 61.210 183.165 61.470 183.485 ;
        RECT 60.810 181.105 60.950 183.165 ;
        RECT 61.670 182.485 61.930 182.805 ;
        RECT 61.210 182.145 61.470 182.465 ;
        RECT 60.750 180.785 61.010 181.105 ;
        RECT 61.270 180.085 61.410 182.145 ;
        RECT 60.750 179.765 61.010 180.085 ;
        RECT 61.210 179.765 61.470 180.085 ;
        RECT 60.810 178.725 60.950 179.765 ;
        RECT 60.750 178.405 61.010 178.725 ;
        RECT 61.730 177.705 61.870 182.485 ;
        RECT 61.670 177.385 61.930 177.705 ;
        RECT 61.730 175.325 61.870 177.385 ;
        RECT 59.830 175.005 60.090 175.325 ;
        RECT 61.670 175.005 61.930 175.325 ;
        RECT 60.750 174.325 61.010 174.645 ;
        RECT 58.910 173.985 59.170 174.305 ;
        RECT 60.810 169.885 60.950 174.325 ;
        RECT 61.210 171.265 61.470 171.585 ;
        RECT 61.270 170.565 61.410 171.265 ;
        RECT 61.210 170.245 61.470 170.565 ;
        RECT 60.750 169.565 61.010 169.885 ;
        RECT 58.910 168.885 59.170 169.205 ;
        RECT 58.970 166.485 59.110 168.885 ;
        RECT 58.910 166.165 59.170 166.485 ;
        RECT 60.290 164.805 60.550 165.125 ;
        RECT 60.350 164.525 60.490 164.805 ;
        RECT 59.890 164.385 60.490 164.525 ;
        RECT 59.890 161.045 60.030 164.385 ;
        RECT 60.290 163.785 60.550 164.105 ;
        RECT 60.350 161.725 60.490 163.785 ;
        RECT 60.290 161.405 60.550 161.725 ;
        RECT 59.830 160.725 60.090 161.045 ;
        RECT 59.370 157.840 59.630 157.985 ;
        RECT 58.440 157.470 58.720 157.840 ;
        RECT 59.360 157.470 59.640 157.840 ;
        RECT 59.890 156.965 60.030 160.725 ;
        RECT 59.830 156.645 60.090 156.965 ;
        RECT 54.770 155.625 55.030 155.945 ;
        RECT 55.690 155.625 55.950 155.945 ;
        RECT 57.530 155.625 57.790 155.945 ;
        RECT 52.930 153.335 53.590 153.475 ;
        RECT 52.930 153.245 53.190 153.335 ;
        RECT 53.850 153.245 54.110 153.565 ;
        RECT 54.830 153.080 54.970 155.625 ;
        RECT 55.230 154.945 55.490 155.265 ;
        RECT 55.290 153.565 55.430 154.945 ;
        RECT 55.230 153.245 55.490 153.565 ;
        RECT 54.760 152.710 55.040 153.080 ;
        RECT 50.865 151.690 52.405 152.060 ;
        RECT 50.170 149.845 50.430 150.165 ;
        RECT 55.230 149.505 55.490 149.825 ;
        RECT 49.710 148.145 49.970 148.465 ;
        RECT 49.250 146.785 49.510 147.105 ;
        RECT 49.310 145.065 49.450 146.785 ;
        RECT 49.770 146.085 49.910 148.145 ;
        RECT 55.290 148.125 55.430 149.505 ;
        RECT 55.230 147.805 55.490 148.125 ;
        RECT 53.390 147.465 53.650 147.785 ;
        RECT 50.865 146.250 52.405 146.620 ;
        RECT 49.710 145.765 49.970 146.085 ;
        RECT 53.450 145.405 53.590 147.465 ;
        RECT 53.390 145.085 53.650 145.405 ;
        RECT 48.790 144.745 49.050 145.065 ;
        RECT 49.250 144.745 49.510 145.065 ;
        RECT 48.850 143.025 48.990 144.745 ;
        RECT 54.770 144.065 55.030 144.385 ;
        RECT 54.830 143.025 54.970 144.065 ;
        RECT 48.790 142.765 49.050 143.025 ;
        RECT 48.790 142.705 49.450 142.765 ;
        RECT 54.770 142.705 55.030 143.025 ;
        RECT 48.850 142.625 49.450 142.705 ;
        RECT 48.790 142.255 49.050 142.345 ;
        RECT 48.390 142.115 49.050 142.255 ;
        RECT 48.790 142.025 49.050 142.115 ;
        RECT 49.310 139.625 49.450 142.625 ;
        RECT 50.170 142.025 50.430 142.345 ;
        RECT 50.230 140.305 50.370 142.025 ;
        RECT 52.930 141.405 53.190 141.665 ;
        RECT 52.930 141.345 55.430 141.405 ;
        RECT 52.990 141.265 55.430 141.345 ;
        RECT 50.865 140.810 52.405 141.180 ;
        RECT 51.550 140.325 51.810 140.645 ;
        RECT 50.170 139.985 50.430 140.305 ;
        RECT 51.610 139.625 51.750 140.325 ;
        RECT 49.250 139.305 49.510 139.625 ;
        RECT 51.090 139.480 51.350 139.625 ;
        RECT 51.080 139.110 51.360 139.480 ;
        RECT 51.550 139.305 51.810 139.625 ;
        RECT 52.470 139.365 52.730 139.625 ;
        RECT 52.070 139.305 52.730 139.365 ;
        RECT 52.070 139.225 52.670 139.305 ;
        RECT 52.070 138.945 52.210 139.225 ;
        RECT 52.010 138.625 52.270 138.945 ;
        RECT 50.865 135.370 52.405 135.740 ;
        RECT 47.870 133.525 48.130 133.845 ;
        RECT 50.170 131.145 50.430 131.465 ;
        RECT 49.250 128.425 49.510 128.745 ;
        RECT 47.410 125.705 47.670 126.025 ;
        RECT 45.570 125.025 45.830 125.345 ;
        RECT 47.470 123.985 47.610 125.705 ;
        RECT 47.410 123.665 47.670 123.985 ;
        RECT 45.570 122.305 45.830 122.625 ;
        RECT 44.190 121.285 44.450 121.605 ;
        RECT 43.730 117.545 43.990 117.865 ;
        RECT 45.630 115.485 45.770 122.305 ;
        RECT 48.330 119.585 48.590 119.905 ;
        RECT 48.390 117.865 48.530 119.585 ;
        RECT 49.310 118.885 49.450 128.425 ;
        RECT 49.710 127.745 49.970 128.065 ;
        RECT 49.770 126.705 49.910 127.745 ;
        RECT 50.230 127.045 50.370 131.145 ;
        RECT 50.865 129.930 52.405 130.300 ;
        RECT 51.550 129.105 51.810 129.425 ;
        RECT 50.170 126.725 50.430 127.045 ;
        RECT 49.710 126.385 49.970 126.705 ;
        RECT 49.710 125.025 49.970 125.345 ;
        RECT 49.770 120.585 49.910 125.025 ;
        RECT 50.230 124.325 50.370 126.725 ;
        RECT 51.610 126.365 51.750 129.105 ;
        RECT 53.850 128.765 54.110 129.085 ;
        RECT 53.390 128.425 53.650 128.745 ;
        RECT 52.920 126.870 53.200 127.240 ;
        RECT 51.550 126.045 51.810 126.365 ;
        RECT 50.865 124.490 52.405 124.860 ;
        RECT 50.170 124.005 50.430 124.325 ;
        RECT 50.230 121.605 50.370 124.005 ;
        RECT 52.990 123.305 53.130 126.870 ;
        RECT 53.450 123.645 53.590 128.425 ;
        RECT 53.910 126.025 54.050 128.765 ;
        RECT 54.310 128.425 54.570 128.745 ;
        RECT 53.850 125.705 54.110 126.025 ;
        RECT 53.910 123.645 54.050 125.705 ;
        RECT 53.390 123.325 53.650 123.645 ;
        RECT 53.850 123.325 54.110 123.645 ;
        RECT 52.930 123.160 53.190 123.305 ;
        RECT 52.920 122.790 53.200 123.160 ;
        RECT 50.170 121.285 50.430 121.605 ;
        RECT 53.450 121.265 53.590 123.325 ;
        RECT 53.390 120.945 53.650 121.265 ;
        RECT 49.710 120.265 49.970 120.585 ;
        RECT 50.865 119.050 52.405 119.420 ;
        RECT 49.250 118.565 49.510 118.885 ;
        RECT 48.330 117.545 48.590 117.865 ;
        RECT 52.010 116.865 52.270 117.185 ;
        RECT 52.070 115.825 52.210 116.865 ;
        RECT 48.330 115.505 48.590 115.825 ;
        RECT 52.010 115.505 52.270 115.825 ;
        RECT 45.570 115.165 45.830 115.485 ;
        RECT 45.570 114.485 45.830 114.805 ;
        RECT 42.350 112.105 42.610 112.425 ;
        RECT 45.630 106.285 45.770 114.485 ;
        RECT 48.390 110.725 48.530 115.505 ;
        RECT 53.910 115.145 54.050 123.325 ;
        RECT 54.370 121.605 54.510 128.425 ;
        RECT 54.770 122.645 55.030 122.965 ;
        RECT 54.830 121.605 54.970 122.645 ;
        RECT 54.310 121.285 54.570 121.605 ;
        RECT 54.770 121.285 55.030 121.605 ;
        RECT 55.290 115.485 55.430 141.265 ;
        RECT 55.750 131.125 55.890 155.625 ;
        RECT 60.350 153.225 60.490 161.405 ;
        RECT 62.190 155.265 62.330 201.185 ;
        RECT 62.650 197.675 62.790 203.905 ;
        RECT 63.110 203.205 63.250 204.505 ;
        RECT 63.050 202.885 63.310 203.205 ;
        RECT 63.570 200.145 63.710 207.305 ;
        RECT 65.350 205.265 65.610 205.585 ;
        RECT 65.410 204.905 65.550 205.265 ;
        RECT 65.350 204.585 65.610 204.905 ;
        RECT 66.270 204.585 66.530 204.905 ;
        RECT 68.110 204.585 68.370 204.905 ;
        RECT 64.260 203.370 65.800 203.740 ;
        RECT 66.330 202.525 66.470 204.585 ;
        RECT 68.170 202.865 68.310 204.585 ;
        RECT 68.110 202.545 68.370 202.865 ;
        RECT 69.090 202.525 69.230 210.025 ;
        RECT 91.050 208.810 92.590 209.180 ;
        RECT 92.950 207.985 93.210 208.305 ;
        RECT 72.250 207.305 72.510 207.625 ;
        RECT 84.670 207.305 84.930 207.625 ;
        RECT 72.310 205.925 72.450 207.305 ;
        RECT 77.655 206.090 79.195 206.460 ;
        RECT 72.250 205.605 72.510 205.925 ;
        RECT 83.750 204.585 84.010 204.905 ;
        RECT 66.270 202.205 66.530 202.525 ;
        RECT 69.030 202.205 69.290 202.525 ;
        RECT 69.090 200.485 69.230 202.205 ;
        RECT 77.655 200.650 79.195 201.020 ;
        RECT 69.030 200.165 69.290 200.485 ;
        RECT 63.510 199.825 63.770 200.145 ;
        RECT 63.510 199.145 63.770 199.465 ;
        RECT 63.050 197.675 63.310 197.765 ;
        RECT 62.650 197.535 63.310 197.675 ;
        RECT 63.050 197.445 63.310 197.535 ;
        RECT 63.570 197.675 63.710 199.145 ;
        RECT 79.150 199.035 79.410 199.125 ;
        RECT 79.150 198.895 79.810 199.035 ;
        RECT 79.150 198.805 79.410 198.895 ;
        RECT 75.930 198.465 76.190 198.785 ;
        RECT 64.260 197.930 65.800 198.300 ;
        RECT 63.570 197.535 64.630 197.675 ;
        RECT 63.050 190.305 63.310 190.625 ;
        RECT 62.590 188.265 62.850 188.585 ;
        RECT 62.650 185.865 62.790 188.265 ;
        RECT 62.590 185.545 62.850 185.865 ;
        RECT 62.650 180.165 62.790 185.545 ;
        RECT 63.110 183.145 63.250 190.305 ;
        RECT 63.570 186.205 63.710 197.535 ;
        RECT 64.490 197.085 64.630 197.535 ;
        RECT 75.990 197.085 76.130 198.465 ;
        RECT 63.970 196.765 64.230 197.085 ;
        RECT 64.430 196.765 64.690 197.085 ;
        RECT 65.810 196.765 66.070 197.085 ;
        RECT 74.090 196.765 74.350 197.085 ;
        RECT 75.930 196.765 76.190 197.085 ;
        RECT 77.310 196.765 77.570 197.085 ;
        RECT 64.030 195.045 64.170 196.765 ;
        RECT 63.970 194.725 64.230 195.045 ;
        RECT 65.870 194.365 66.010 196.765 ;
        RECT 67.650 196.085 67.910 196.405 ;
        RECT 73.630 196.085 73.890 196.405 ;
        RECT 66.730 194.385 66.990 194.705 ;
        RECT 65.810 194.045 66.070 194.365 ;
        RECT 66.270 193.705 66.530 194.025 ;
        RECT 64.260 192.490 65.800 192.860 ;
        RECT 64.260 187.050 65.800 187.420 ;
        RECT 65.350 186.565 65.610 186.885 ;
        RECT 65.410 186.205 65.550 186.565 ;
        RECT 66.330 186.205 66.470 193.705 ;
        RECT 66.790 186.545 66.930 194.385 ;
        RECT 67.710 194.025 67.850 196.085 ;
        RECT 68.570 195.745 68.830 196.065 ;
        RECT 67.650 193.705 67.910 194.025 ;
        RECT 68.630 193.345 68.770 195.745 ;
        RECT 67.650 193.025 67.910 193.345 ;
        RECT 68.570 193.025 68.830 193.345 ;
        RECT 71.330 193.025 71.590 193.345 ;
        RECT 67.710 191.645 67.850 193.025 ;
        RECT 67.650 191.325 67.910 191.645 ;
        RECT 68.630 191.305 68.770 193.025 ;
        RECT 71.390 192.325 71.530 193.025 ;
        RECT 71.330 192.005 71.590 192.325 ;
        RECT 68.570 190.985 68.830 191.305 ;
        RECT 66.730 186.225 66.990 186.545 ;
        RECT 69.030 186.225 69.290 186.545 ;
        RECT 63.510 185.885 63.770 186.205 ;
        RECT 64.890 185.885 65.150 186.205 ;
        RECT 65.350 185.885 65.610 186.205 ;
        RECT 65.810 185.885 66.070 186.205 ;
        RECT 66.270 185.885 66.530 186.205 ;
        RECT 64.950 184.165 65.090 185.885 ;
        RECT 65.410 185.185 65.550 185.885 ;
        RECT 65.350 184.865 65.610 185.185 ;
        RECT 64.890 183.845 65.150 184.165 ;
        RECT 63.050 182.825 63.310 183.145 ;
        RECT 63.110 180.765 63.250 182.825 ;
        RECT 65.410 182.805 65.550 184.865 ;
        RECT 65.870 183.485 66.010 185.885 ;
        RECT 66.330 183.735 66.470 185.885 ;
        RECT 66.730 183.735 66.990 183.825 ;
        RECT 66.330 183.595 66.990 183.735 ;
        RECT 66.730 183.505 66.990 183.595 ;
        RECT 65.810 183.395 66.070 183.485 ;
        RECT 65.810 183.255 66.470 183.395 ;
        RECT 65.810 183.165 66.070 183.255 ;
        RECT 65.350 182.485 65.610 182.805 ;
        RECT 64.260 181.610 65.800 181.980 ;
        RECT 66.330 181.105 66.470 183.255 ;
        RECT 66.270 180.785 66.530 181.105 ;
        RECT 66.790 180.765 66.930 183.505 ;
        RECT 69.090 183.485 69.230 186.225 ;
        RECT 69.490 184.865 69.750 185.185 ;
        RECT 69.550 183.485 69.690 184.865 ;
        RECT 67.190 183.165 67.450 183.485 ;
        RECT 69.030 183.165 69.290 183.485 ;
        RECT 69.490 183.165 69.750 183.485 ;
        RECT 63.050 180.445 63.310 180.765 ;
        RECT 66.730 180.445 66.990 180.765 ;
        RECT 62.650 180.025 63.250 180.165 ;
        RECT 62.590 179.425 62.850 179.745 ;
        RECT 62.650 177.705 62.790 179.425 ;
        RECT 62.590 177.385 62.850 177.705 ;
        RECT 62.650 175.665 62.790 177.385 ;
        RECT 62.590 175.345 62.850 175.665 ;
        RECT 62.590 173.985 62.850 174.305 ;
        RECT 62.650 173.285 62.790 173.985 ;
        RECT 62.590 172.965 62.850 173.285 ;
        RECT 63.110 169.205 63.250 180.025 ;
        RECT 66.730 179.425 66.990 179.745 ;
        RECT 66.790 178.045 66.930 179.425 ;
        RECT 65.810 177.725 66.070 178.045 ;
        RECT 66.730 177.725 66.990 178.045 ;
        RECT 65.870 177.445 66.010 177.725 ;
        RECT 65.870 177.305 66.930 177.445 ;
        RECT 63.510 176.705 63.770 177.025 ;
        RECT 66.270 176.705 66.530 177.025 ;
        RECT 63.050 168.885 63.310 169.205 ;
        RECT 62.590 155.285 62.850 155.605 ;
        RECT 62.130 154.945 62.390 155.265 ;
        RECT 62.190 153.565 62.330 154.945 ;
        RECT 62.130 153.245 62.390 153.565 ;
        RECT 60.290 152.905 60.550 153.225 ;
        RECT 57.990 146.785 58.250 147.105 ;
        RECT 57.530 145.765 57.790 146.085 ;
        RECT 56.150 144.405 56.410 144.725 ;
        RECT 55.690 130.805 55.950 131.125 ;
        RECT 55.750 129.765 55.890 130.805 ;
        RECT 55.690 129.445 55.950 129.765 ;
        RECT 55.690 125.025 55.950 125.345 ;
        RECT 55.750 120.925 55.890 125.025 ;
        RECT 55.690 120.605 55.950 120.925 ;
        RECT 56.210 115.485 56.350 144.405 ;
        RECT 57.590 139.625 57.730 145.765 ;
        RECT 58.050 144.725 58.190 146.785 ;
        RECT 57.990 144.405 58.250 144.725 ;
        RECT 57.990 141.685 58.250 142.005 ;
        RECT 58.050 139.625 58.190 141.685 ;
        RECT 58.450 141.345 58.710 141.665 ;
        RECT 58.510 139.625 58.650 141.345 ;
        RECT 60.350 140.645 60.490 152.905 ;
        RECT 62.120 152.710 62.400 153.080 ;
        RECT 62.190 152.545 62.330 152.710 ;
        RECT 61.210 152.225 61.470 152.545 ;
        RECT 62.130 152.225 62.390 152.545 ;
        RECT 60.750 150.185 61.010 150.505 ;
        RECT 60.290 140.325 60.550 140.645 ;
        RECT 57.530 139.305 57.790 139.625 ;
        RECT 57.990 139.305 58.250 139.625 ;
        RECT 58.450 139.305 58.710 139.625 ;
        RECT 57.590 137.925 57.730 139.305 ;
        RECT 59.830 138.965 60.090 139.285 ;
        RECT 57.530 137.605 57.790 137.925 ;
        RECT 59.890 137.245 60.030 138.965 ;
        RECT 59.830 136.925 60.090 137.245 ;
        RECT 59.890 135.205 60.030 136.925 ;
        RECT 60.350 136.905 60.490 140.325 ;
        RECT 60.290 136.585 60.550 136.905 ;
        RECT 59.830 134.885 60.090 135.205 ;
        RECT 59.890 132.485 60.030 134.885 ;
        RECT 59.830 132.165 60.090 132.485 ;
        RECT 60.350 131.465 60.490 136.585 ;
        RECT 60.810 134.525 60.950 150.185 ;
        RECT 61.270 150.165 61.410 152.225 ;
        RECT 62.650 151.525 62.790 155.285 ;
        RECT 62.590 151.205 62.850 151.525 ;
        RECT 63.110 150.505 63.250 168.885 ;
        RECT 63.570 167.165 63.710 176.705 ;
        RECT 64.260 176.170 65.800 176.540 ;
        RECT 66.330 175.405 66.470 176.705 ;
        RECT 65.870 175.325 66.470 175.405 ;
        RECT 66.790 175.325 66.930 177.305 ;
        RECT 65.810 175.265 66.470 175.325 ;
        RECT 65.810 175.005 66.070 175.265 ;
        RECT 66.730 175.005 66.990 175.325 ;
        RECT 64.260 170.730 65.800 171.100 ;
        RECT 66.790 170.645 66.930 175.005 ;
        RECT 66.330 170.505 66.930 170.645 ;
        RECT 63.970 169.565 64.230 169.885 ;
        RECT 65.810 169.565 66.070 169.885 ;
        RECT 63.510 166.845 63.770 167.165 ;
        RECT 64.030 166.825 64.170 169.565 ;
        RECT 65.870 169.205 66.010 169.565 ;
        RECT 65.810 168.885 66.070 169.205 ;
        RECT 64.430 168.545 64.690 168.865 ;
        RECT 63.970 166.505 64.230 166.825 ;
        RECT 64.490 166.485 64.630 168.545 ;
        RECT 64.430 166.165 64.690 166.485 ;
        RECT 64.260 165.290 65.800 165.660 ;
        RECT 66.330 162.065 66.470 170.505 ;
        RECT 67.250 169.965 67.390 183.165 ;
        RECT 67.650 182.485 67.910 182.805 ;
        RECT 66.790 169.825 67.390 169.965 ;
        RECT 66.270 161.745 66.530 162.065 ;
        RECT 64.260 159.850 65.800 160.220 ;
        RECT 65.810 158.685 66.070 159.005 ;
        RECT 64.430 157.665 64.690 157.985 ;
        RECT 64.490 156.285 64.630 157.665 ;
        RECT 64.430 155.965 64.690 156.285 ;
        RECT 65.870 155.125 66.010 158.685 ;
        RECT 66.330 156.625 66.470 161.745 ;
        RECT 66.790 159.005 66.930 169.825 ;
        RECT 67.190 168.885 67.450 169.205 ;
        RECT 67.250 164.785 67.390 168.885 ;
        RECT 67.190 164.465 67.450 164.785 ;
        RECT 66.730 158.685 66.990 159.005 ;
        RECT 66.790 156.965 66.930 158.685 ;
        RECT 66.730 156.645 66.990 156.965 ;
        RECT 66.270 156.305 66.530 156.625 ;
        RECT 66.790 156.365 66.930 156.645 ;
        RECT 66.790 156.225 67.390 156.365 ;
        RECT 65.870 154.985 66.470 155.125 ;
        RECT 64.260 154.410 65.800 154.780 ;
        RECT 65.810 153.925 66.070 154.245 ;
        RECT 65.870 151.185 66.010 153.925 ;
        RECT 65.810 150.865 66.070 151.185 ;
        RECT 63.050 150.185 63.310 150.505 ;
        RECT 61.210 149.845 61.470 150.165 ;
        RECT 64.260 148.970 65.800 149.340 ;
        RECT 66.330 147.640 66.470 154.985 ;
        RECT 67.250 153.565 67.390 156.225 ;
        RECT 67.190 153.245 67.450 153.565 ;
        RECT 67.710 148.125 67.850 182.485 ;
        RECT 68.110 180.445 68.370 180.765 ;
        RECT 68.170 174.305 68.310 180.445 ;
        RECT 70.870 174.665 71.130 174.985 ;
        RECT 68.110 173.985 68.370 174.305 ;
        RECT 69.490 173.985 69.750 174.305 ;
        RECT 68.170 171.585 68.310 173.985 ;
        RECT 69.550 173.285 69.690 173.985 ;
        RECT 69.490 172.965 69.750 173.285 ;
        RECT 68.570 171.945 68.830 172.265 ;
        RECT 68.110 171.265 68.370 171.585 ;
        RECT 68.630 169.885 68.770 171.945 ;
        RECT 69.490 171.265 69.750 171.585 ;
        RECT 69.550 170.565 69.690 171.265 ;
        RECT 69.490 170.245 69.750 170.565 ;
        RECT 69.550 169.885 69.690 170.245 ;
        RECT 68.570 169.565 68.830 169.885 ;
        RECT 69.030 169.565 69.290 169.885 ;
        RECT 69.490 169.565 69.750 169.885 ;
        RECT 69.090 169.400 69.230 169.565 ;
        RECT 69.020 169.030 69.300 169.400 ;
        RECT 68.110 165.825 68.370 166.145 ;
        RECT 69.950 165.825 70.210 166.145 ;
        RECT 68.170 161.920 68.310 165.825 ;
        RECT 70.010 163.425 70.150 165.825 ;
        RECT 69.950 163.105 70.210 163.425 ;
        RECT 68.100 161.550 68.380 161.920 ;
        RECT 68.170 158.665 68.310 161.550 ;
        RECT 70.930 161.385 71.070 174.665 ;
        RECT 69.490 161.065 69.750 161.385 ;
        RECT 70.870 161.065 71.130 161.385 ;
        RECT 68.570 159.365 68.830 159.685 ;
        RECT 68.110 158.345 68.370 158.665 ;
        RECT 68.630 156.965 68.770 159.365 ;
        RECT 69.550 159.005 69.690 161.065 ;
        RECT 70.870 160.385 71.130 160.705 ;
        RECT 70.930 159.005 71.070 160.385 ;
        RECT 69.490 158.685 69.750 159.005 ;
        RECT 70.870 158.685 71.130 159.005 ;
        RECT 68.570 156.645 68.830 156.965 ;
        RECT 68.110 156.305 68.370 156.625 ;
        RECT 67.650 147.805 67.910 148.125 ;
        RECT 66.260 147.270 66.540 147.640 ;
        RECT 63.510 146.785 63.770 147.105 ;
        RECT 63.050 145.085 63.310 145.405 ;
        RECT 61.210 142.025 61.470 142.345 ;
        RECT 61.270 140.645 61.410 142.025 ;
        RECT 61.660 141.830 61.940 142.200 ;
        RECT 61.210 140.325 61.470 140.645 ;
        RECT 60.750 134.205 61.010 134.525 ;
        RECT 60.290 131.145 60.550 131.465 ;
        RECT 57.070 130.465 57.330 130.785 ;
        RECT 57.130 126.025 57.270 130.465 ;
        RECT 60.810 126.365 60.950 134.205 ;
        RECT 60.750 126.045 61.010 126.365 ;
        RECT 57.070 125.705 57.330 126.025 ;
        RECT 60.810 124.235 60.950 126.045 ;
        RECT 60.350 124.095 60.950 124.235 ;
        RECT 60.350 120.925 60.490 124.095 ;
        RECT 60.750 123.325 61.010 123.645 ;
        RECT 60.810 121.605 60.950 123.325 ;
        RECT 60.750 121.285 61.010 121.605 ;
        RECT 60.290 120.605 60.550 120.925 ;
        RECT 60.350 117.865 60.490 120.605 ;
        RECT 61.730 117.865 61.870 141.830 ;
        RECT 63.110 140.645 63.250 145.085 ;
        RECT 63.050 140.325 63.310 140.645 ;
        RECT 63.570 137.585 63.710 146.785 ;
        RECT 65.810 144.975 66.070 145.065 ;
        RECT 65.810 144.835 66.470 144.975 ;
        RECT 65.810 144.745 66.070 144.835 ;
        RECT 64.260 143.530 65.800 143.900 ;
        RECT 65.810 142.085 66.070 142.345 ;
        RECT 66.330 142.085 66.470 144.835 ;
        RECT 65.810 142.025 66.470 142.085 ;
        RECT 65.870 141.945 66.470 142.025 ;
        RECT 64.260 138.090 65.800 138.460 ;
        RECT 63.510 137.265 63.770 137.585 ;
        RECT 64.430 135.905 64.690 136.225 ;
        RECT 65.810 135.905 66.070 136.225 ;
        RECT 64.490 134.525 64.630 135.905 ;
        RECT 64.430 134.205 64.690 134.525 ;
        RECT 65.870 133.845 66.010 135.905 ;
        RECT 66.330 134.185 66.470 141.945 ;
        RECT 67.190 135.905 67.450 136.225 ;
        RECT 67.250 134.185 67.390 135.905 ;
        RECT 66.270 133.865 66.530 134.185 ;
        RECT 67.190 133.865 67.450 134.185 ;
        RECT 65.810 133.525 66.070 133.845 ;
        RECT 64.260 132.650 65.800 133.020 ;
        RECT 65.350 130.465 65.610 130.785 ;
        RECT 65.410 129.085 65.550 130.465 ;
        RECT 65.350 128.765 65.610 129.085 ;
        RECT 66.330 128.745 66.470 133.865 ;
        RECT 66.730 133.525 66.990 133.845 ;
        RECT 66.790 131.805 66.930 133.525 ;
        RECT 67.250 133.505 67.390 133.865 ;
        RECT 67.190 133.185 67.450 133.505 ;
        RECT 66.730 131.485 66.990 131.805 ;
        RECT 68.170 131.465 68.310 156.305 ;
        RECT 69.550 156.285 69.690 158.685 ;
        RECT 69.490 155.965 69.750 156.285 ;
        RECT 69.030 154.945 69.290 155.265 ;
        RECT 69.090 153.905 69.230 154.945 ;
        RECT 69.030 153.585 69.290 153.905 ;
        RECT 69.550 153.565 69.690 155.965 ;
        RECT 70.410 155.625 70.670 155.945 ;
        RECT 70.870 155.625 71.130 155.945 ;
        RECT 70.470 155.265 70.610 155.625 ;
        RECT 70.410 154.945 70.670 155.265 ;
        RECT 69.490 153.245 69.750 153.565 ;
        RECT 70.930 153.225 71.070 155.625 ;
        RECT 71.390 153.645 71.530 192.005 ;
        RECT 73.170 191.325 73.430 191.645 ;
        RECT 72.710 184.925 72.970 185.185 ;
        RECT 73.230 184.925 73.370 191.325 ;
        RECT 73.690 191.305 73.830 196.085 ;
        RECT 73.630 190.985 73.890 191.305 ;
        RECT 73.690 188.925 73.830 190.985 ;
        RECT 73.630 188.605 73.890 188.925 ;
        RECT 72.710 184.865 73.370 184.925 ;
        RECT 72.770 184.785 73.370 184.865 ;
        RECT 73.230 183.145 73.370 184.785 ;
        RECT 73.690 183.485 73.830 188.605 ;
        RECT 74.150 188.585 74.290 196.765 ;
        RECT 74.550 196.425 74.810 196.745 ;
        RECT 74.610 193.685 74.750 196.425 ;
        RECT 74.550 193.365 74.810 193.685 ;
        RECT 74.090 188.265 74.350 188.585 ;
        RECT 74.150 185.865 74.290 188.265 ;
        RECT 74.550 187.585 74.810 187.905 ;
        RECT 74.610 186.545 74.750 187.585 ;
        RECT 74.550 186.225 74.810 186.545 ;
        RECT 74.090 185.545 74.350 185.865 ;
        RECT 74.090 184.865 74.350 185.185 ;
        RECT 73.630 183.165 73.890 183.485 ;
        RECT 73.170 182.825 73.430 183.145 ;
        RECT 71.790 178.065 72.050 178.385 ;
        RECT 71.850 172.175 71.990 178.065 ;
        RECT 73.230 173.195 73.370 182.825 ;
        RECT 73.690 181.105 73.830 183.165 ;
        RECT 74.150 182.465 74.290 184.865 ;
        RECT 74.090 182.145 74.350 182.465 ;
        RECT 73.630 180.785 73.890 181.105 ;
        RECT 72.770 173.055 73.370 173.195 ;
        RECT 72.250 172.175 72.510 172.265 ;
        RECT 71.850 172.035 72.510 172.175 ;
        RECT 71.850 169.885 71.990 172.035 ;
        RECT 72.250 171.945 72.510 172.035 ;
        RECT 72.250 171.440 72.510 171.585 ;
        RECT 72.240 171.070 72.520 171.440 ;
        RECT 72.770 169.965 72.910 173.055 ;
        RECT 73.630 171.265 73.890 171.585 ;
        RECT 71.790 169.565 72.050 169.885 ;
        RECT 72.770 169.825 73.370 169.965 ;
        RECT 71.790 169.115 72.050 169.205 ;
        RECT 71.790 168.975 72.450 169.115 ;
        RECT 72.700 169.030 72.980 169.400 ;
        RECT 71.790 168.885 72.050 168.975 ;
        RECT 71.390 153.505 71.990 153.645 ;
        RECT 70.870 152.905 71.130 153.225 ;
        RECT 70.930 150.505 71.070 152.905 ;
        RECT 71.330 150.865 71.590 151.185 ;
        RECT 70.870 150.185 71.130 150.505 ;
        RECT 70.870 147.125 71.130 147.445 ;
        RECT 70.930 144.805 71.070 147.125 ;
        RECT 71.390 145.405 71.530 150.865 ;
        RECT 71.850 150.505 71.990 153.505 ;
        RECT 71.790 150.185 72.050 150.505 ;
        RECT 71.790 146.785 72.050 147.105 ;
        RECT 71.330 145.085 71.590 145.405 ;
        RECT 70.930 144.665 71.530 144.805 ;
        RECT 69.950 144.065 70.210 144.385 ;
        RECT 69.490 134.885 69.750 135.205 ;
        RECT 68.570 133.185 68.830 133.505 ;
        RECT 68.630 132.485 68.770 133.185 ;
        RECT 68.570 132.165 68.830 132.485 ;
        RECT 68.110 131.145 68.370 131.465 ;
        RECT 66.270 128.425 66.530 128.745 ;
        RECT 62.590 128.085 62.850 128.405 ;
        RECT 62.650 127.045 62.790 128.085 ;
        RECT 64.260 127.210 65.800 127.580 ;
        RECT 62.590 126.725 62.850 127.045 ;
        RECT 68.170 124.325 68.310 131.145 ;
        RECT 69.550 126.365 69.690 134.885 ;
        RECT 69.490 126.045 69.750 126.365 ;
        RECT 68.110 124.005 68.370 124.325 ;
        RECT 64.260 121.770 65.800 122.140 ;
        RECT 70.010 118.545 70.150 144.065 ;
        RECT 70.400 140.470 70.680 140.840 ;
        RECT 70.470 139.625 70.610 140.470 ;
        RECT 70.870 140.325 71.130 140.645 ;
        RECT 70.410 139.305 70.670 139.625 ;
        RECT 70.410 138.625 70.670 138.945 ;
        RECT 69.950 118.225 70.210 118.545 ;
        RECT 59.370 117.545 59.630 117.865 ;
        RECT 60.290 117.545 60.550 117.865 ;
        RECT 61.670 117.545 61.930 117.865 ;
        RECT 57.990 116.865 58.250 117.185 ;
        RECT 58.050 115.825 58.190 116.865 ;
        RECT 57.990 115.505 58.250 115.825 ;
        RECT 55.230 115.165 55.490 115.485 ;
        RECT 56.150 115.165 56.410 115.485 ;
        RECT 53.850 114.825 54.110 115.145 ;
        RECT 52.930 114.145 53.190 114.465 ;
        RECT 50.865 113.610 52.405 113.980 ;
        RECT 50.170 112.445 50.430 112.765 ;
        RECT 48.330 110.405 48.590 110.725 ;
        RECT 50.230 107.405 50.370 112.445 ;
        RECT 52.990 112.085 53.130 114.145 ;
        RECT 53.910 113.445 54.050 114.825 ;
        RECT 57.070 114.145 57.330 114.465 ;
        RECT 53.850 113.125 54.110 113.445 ;
        RECT 53.910 112.765 54.050 113.125 ;
        RECT 57.130 112.765 57.270 114.145 ;
        RECT 53.850 112.445 54.110 112.765 ;
        RECT 57.070 112.445 57.330 112.765 ;
        RECT 52.010 111.765 52.270 112.085 ;
        RECT 52.930 111.765 53.190 112.085 ;
        RECT 56.610 111.765 56.870 112.085 ;
        RECT 57.990 111.765 58.250 112.085 ;
        RECT 52.070 110.725 52.210 111.765 ;
        RECT 52.010 110.405 52.270 110.725 ;
        RECT 50.865 108.170 52.405 108.540 ;
        RECT 50.230 107.265 51.290 107.405 ;
        RECT 51.150 106.285 51.290 107.265 ;
        RECT 56.670 106.285 56.810 111.765 ;
        RECT 58.050 110.725 58.190 111.765 ;
        RECT 57.990 110.405 58.250 110.725 ;
        RECT 59.430 110.045 59.570 117.545 ;
        RECT 70.470 117.525 70.610 138.625 ;
        RECT 70.930 135.205 71.070 140.325 ;
        RECT 71.390 137.925 71.530 144.665 ;
        RECT 71.850 144.125 71.990 146.785 ;
        RECT 72.310 145.065 72.450 168.975 ;
        RECT 72.710 168.885 72.970 169.030 ;
        RECT 72.710 158.685 72.970 159.005 ;
        RECT 72.770 155.945 72.910 158.685 ;
        RECT 73.230 157.840 73.370 169.825 ;
        RECT 73.690 159.880 73.830 171.265 ;
        RECT 73.620 159.510 73.900 159.880 ;
        RECT 73.630 158.915 73.890 159.005 ;
        RECT 74.150 158.915 74.290 182.145 ;
        RECT 75.470 174.665 75.730 174.985 ;
        RECT 75.010 171.945 75.270 172.265 ;
        RECT 75.070 169.885 75.210 171.945 ;
        RECT 75.010 169.565 75.270 169.885 ;
        RECT 75.530 169.545 75.670 174.665 ;
        RECT 75.470 169.225 75.730 169.545 ;
        RECT 75.470 168.545 75.730 168.865 ;
        RECT 74.550 167.185 74.810 167.505 ;
        RECT 74.610 159.005 74.750 167.185 ;
        RECT 73.630 158.775 74.290 158.915 ;
        RECT 73.630 158.685 73.890 158.775 ;
        RECT 74.550 158.685 74.810 159.005 ;
        RECT 75.010 158.005 75.270 158.325 ;
        RECT 73.160 157.470 73.440 157.840 ;
        RECT 74.540 157.045 74.820 157.160 ;
        RECT 74.150 156.965 74.820 157.045 ;
        RECT 74.090 156.905 74.820 156.965 ;
        RECT 74.090 156.645 74.350 156.905 ;
        RECT 74.540 156.790 74.820 156.905 ;
        RECT 72.710 155.625 72.970 155.945 ;
        RECT 74.090 155.855 74.350 155.945 ;
        RECT 74.090 155.715 74.750 155.855 ;
        RECT 74.090 155.625 74.350 155.715 ;
        RECT 74.610 155.685 74.750 155.715 ;
        RECT 75.070 155.685 75.210 158.005 ;
        RECT 74.610 155.545 75.210 155.685 ;
        RECT 73.160 154.070 73.440 154.440 ;
        RECT 73.170 153.925 73.430 154.070 ;
        RECT 74.090 153.925 74.350 154.245 ;
        RECT 73.170 153.475 73.430 153.565 ;
        RECT 72.770 153.335 73.430 153.475 ;
        RECT 72.770 150.505 72.910 153.335 ;
        RECT 73.170 153.245 73.430 153.335 ;
        RECT 73.630 153.245 73.890 153.565 ;
        RECT 73.160 152.710 73.440 153.080 ;
        RECT 72.710 150.185 72.970 150.505 ;
        RECT 73.230 148.125 73.370 152.710 ;
        RECT 73.690 150.505 73.830 153.245 ;
        RECT 73.630 150.185 73.890 150.505 ;
        RECT 73.170 147.805 73.430 148.125 ;
        RECT 74.150 147.785 74.290 153.925 ;
        RECT 74.610 153.905 74.750 155.545 ;
        RECT 75.010 154.945 75.270 155.265 ;
        RECT 75.070 153.905 75.210 154.945 ;
        RECT 74.550 153.585 74.810 153.905 ;
        RECT 75.010 153.585 75.270 153.905 ;
        RECT 75.010 152.225 75.270 152.545 ;
        RECT 74.550 149.505 74.810 149.825 ;
        RECT 74.610 148.465 74.750 149.505 ;
        RECT 74.550 148.145 74.810 148.465 ;
        RECT 74.090 147.465 74.350 147.785 ;
        RECT 72.710 145.765 72.970 146.085 ;
        RECT 72.250 144.745 72.510 145.065 ;
        RECT 71.850 143.985 72.450 144.125 ;
        RECT 71.790 141.685 72.050 142.005 ;
        RECT 71.850 139.625 71.990 141.685 ;
        RECT 71.790 139.305 72.050 139.625 ;
        RECT 71.330 137.605 71.590 137.925 ;
        RECT 70.870 134.885 71.130 135.205 ;
        RECT 72.310 117.865 72.450 143.985 ;
        RECT 72.770 137.925 72.910 145.765 ;
        RECT 73.170 144.065 73.430 144.385 ;
        RECT 73.230 142.345 73.370 144.065 ;
        RECT 73.170 142.025 73.430 142.345 ;
        RECT 74.550 141.345 74.810 141.665 ;
        RECT 73.170 140.325 73.430 140.645 ;
        RECT 72.710 137.605 72.970 137.925 ;
        RECT 73.230 135.205 73.370 140.325 ;
        RECT 74.610 139.625 74.750 141.345 ;
        RECT 75.070 139.965 75.210 152.225 ;
        RECT 75.530 140.305 75.670 168.545 ;
        RECT 75.990 156.285 76.130 196.765 ;
        RECT 77.370 192.325 77.510 196.765 ;
        RECT 77.655 195.210 79.195 195.580 ;
        RECT 79.670 195.045 79.810 198.895 ;
        RECT 83.810 197.765 83.950 204.585 ;
        RECT 84.730 203.425 84.870 207.305 ;
        RECT 90.650 206.625 90.910 206.945 ;
        RECT 86.050 203.905 86.310 204.225 ;
        RECT 84.730 203.285 85.790 203.425 ;
        RECT 85.650 202.185 85.790 203.285 ;
        RECT 86.110 202.865 86.250 203.905 ;
        RECT 86.050 202.545 86.310 202.865 ;
        RECT 85.590 201.865 85.850 202.185 ;
        RECT 85.650 199.465 85.790 201.865 ;
        RECT 84.210 199.145 84.470 199.465 ;
        RECT 85.590 199.145 85.850 199.465 ;
        RECT 84.270 197.765 84.410 199.145 ;
        RECT 83.750 197.445 84.010 197.765 ;
        RECT 84.210 197.445 84.470 197.765 ;
        RECT 79.610 194.725 79.870 195.045 ;
        RECT 85.650 194.365 85.790 199.145 ;
        RECT 90.710 199.125 90.850 206.625 ;
        RECT 91.050 203.370 92.590 203.740 ;
        RECT 93.010 203.205 93.150 207.985 ;
        RECT 99.850 207.305 100.110 207.625 ;
        RECT 101.690 207.305 101.950 207.625 ;
        RECT 93.410 204.585 93.670 204.905 ;
        RECT 92.950 202.885 93.210 203.205 ;
        RECT 92.950 202.205 93.210 202.525 ;
        RECT 90.650 198.805 90.910 199.125 ;
        RECT 91.050 197.930 92.590 198.300 ;
        RECT 93.010 196.745 93.150 202.205 ;
        RECT 93.470 202.185 93.610 204.585 ;
        RECT 98.930 204.245 99.190 204.565 ;
        RECT 93.870 203.905 94.130 204.225 ;
        RECT 93.930 202.525 94.070 203.905 ;
        RECT 98.990 203.205 99.130 204.245 ;
        RECT 99.910 203.205 100.050 207.305 ;
        RECT 101.750 204.905 101.890 207.305 ;
        RECT 104.445 206.090 105.985 206.460 ;
        RECT 101.690 204.585 101.950 204.905 ;
        RECT 103.990 204.585 104.250 204.905 ;
        RECT 98.930 202.885 99.190 203.205 ;
        RECT 99.850 202.885 100.110 203.205 ;
        RECT 93.870 202.205 94.130 202.525 ;
        RECT 99.390 202.205 99.650 202.525 ;
        RECT 93.410 201.865 93.670 202.185 ;
        RECT 94.790 201.865 95.050 202.185 ;
        RECT 96.630 201.865 96.890 202.185 ;
        RECT 93.470 197.085 93.610 201.865 ;
        RECT 94.850 199.885 94.990 201.865 ;
        RECT 94.850 199.805 95.450 199.885 ;
        RECT 94.850 199.745 95.510 199.805 ;
        RECT 95.250 199.485 95.510 199.745 ;
        RECT 93.410 196.765 93.670 197.085 ;
        RECT 92.950 196.425 93.210 196.745 ;
        RECT 91.110 196.085 91.370 196.405 ;
        RECT 86.970 194.385 87.230 194.705 ;
        RECT 80.530 194.045 80.790 194.365 ;
        RECT 85.590 194.045 85.850 194.365 ;
        RECT 78.690 193.705 78.950 194.025 ;
        RECT 78.750 192.325 78.890 193.705 ;
        RECT 77.310 192.005 77.570 192.325 ;
        RECT 78.690 192.005 78.950 192.325 ;
        RECT 80.590 191.985 80.730 194.045 ;
        RECT 82.830 193.705 83.090 194.025 ;
        RECT 80.530 191.665 80.790 191.985 ;
        RECT 82.890 191.645 83.030 193.705 ;
        RECT 85.130 193.365 85.390 193.685 ;
        RECT 82.830 191.325 83.090 191.645 ;
        RECT 77.655 189.770 79.195 190.140 ;
        RECT 82.890 189.605 83.030 191.325 ;
        RECT 85.190 190.625 85.330 193.365 ;
        RECT 85.650 191.305 85.790 194.045 ;
        RECT 85.590 190.985 85.850 191.305 ;
        RECT 85.130 190.305 85.390 190.625 ;
        RECT 78.690 189.285 78.950 189.605 ;
        RECT 82.830 189.285 83.090 189.605 ;
        RECT 78.750 188.585 78.890 189.285 ;
        RECT 78.690 188.265 78.950 188.585 ;
        RECT 80.990 188.265 81.250 188.585 ;
        RECT 79.150 187.925 79.410 188.245 ;
        RECT 79.610 187.925 79.870 188.245 ;
        RECT 77.770 187.585 78.030 187.905 ;
        RECT 77.830 186.545 77.970 187.585 ;
        RECT 79.210 186.545 79.350 187.925 ;
        RECT 77.770 186.225 78.030 186.545 ;
        RECT 79.150 186.225 79.410 186.545 ;
        RECT 79.670 185.185 79.810 187.925 ;
        RECT 79.610 184.865 79.870 185.185 ;
        RECT 77.655 184.330 79.195 184.700 ;
        RECT 81.050 184.165 81.190 188.265 ;
        RECT 82.890 184.165 83.030 189.285 ;
        RECT 85.190 187.905 85.330 190.305 ;
        RECT 85.130 187.585 85.390 187.905 ;
        RECT 80.990 183.845 81.250 184.165 ;
        RECT 82.830 183.845 83.090 184.165 ;
        RECT 84.670 183.000 84.930 183.145 ;
        RECT 84.660 182.630 84.940 183.000 ;
        RECT 77.655 178.890 79.195 179.260 ;
        RECT 80.530 177.725 80.790 178.045 ;
        RECT 79.610 177.045 79.870 177.365 ;
        RECT 76.390 176.705 76.650 177.025 ;
        RECT 76.450 176.005 76.590 176.705 ;
        RECT 76.390 175.685 76.650 176.005 ;
        RECT 76.450 172.945 76.590 175.685 ;
        RECT 79.670 175.665 79.810 177.045 ;
        RECT 79.610 175.345 79.870 175.665 ;
        RECT 80.590 175.325 80.730 177.725 ;
        RECT 83.290 177.385 83.550 177.705 ;
        RECT 83.350 176.005 83.490 177.385 ;
        RECT 83.290 175.685 83.550 176.005 ;
        RECT 76.850 175.005 77.110 175.325 ;
        RECT 80.530 175.005 80.790 175.325 ;
        RECT 81.450 175.005 81.710 175.325 ;
        RECT 81.910 175.005 82.170 175.325 ;
        RECT 76.390 172.625 76.650 172.945 ;
        RECT 76.910 170.565 77.050 175.005 ;
        RECT 77.655 173.450 79.195 173.820 ;
        RECT 80.590 172.605 80.730 175.005 ;
        RECT 81.510 173.285 81.650 175.005 ;
        RECT 81.450 172.965 81.710 173.285 ;
        RECT 80.530 172.285 80.790 172.605 ;
        RECT 77.310 171.945 77.570 172.265 ;
        RECT 76.850 170.245 77.110 170.565 ;
        RECT 76.910 167.845 77.050 170.245 ;
        RECT 76.850 167.525 77.110 167.845 ;
        RECT 77.370 159.005 77.510 171.945 ;
        RECT 79.610 171.265 79.870 171.585 ;
        RECT 80.530 171.265 80.790 171.585 ;
        RECT 77.655 168.010 79.195 168.380 ;
        RECT 79.670 166.485 79.810 171.265 ;
        RECT 80.590 169.885 80.730 171.265 ;
        RECT 80.530 169.565 80.790 169.885 ;
        RECT 81.970 169.205 82.110 175.005 ;
        RECT 84.210 173.985 84.470 174.305 ;
        RECT 83.750 171.265 84.010 171.585 ;
        RECT 83.810 170.225 83.950 171.265 ;
        RECT 83.750 169.905 84.010 170.225 ;
        RECT 81.910 168.885 82.170 169.205 ;
        RECT 84.270 167.165 84.410 173.985 ;
        RECT 84.210 166.845 84.470 167.165 ;
        RECT 79.610 166.165 79.870 166.485 ;
        RECT 77.655 162.570 79.195 162.940 ;
        RECT 85.190 161.725 85.330 187.585 ;
        RECT 85.650 185.865 85.790 190.985 ;
        RECT 87.030 188.585 87.170 194.385 ;
        RECT 91.170 194.365 91.310 196.085 ;
        RECT 91.110 194.045 91.370 194.365 ;
        RECT 88.350 193.025 88.610 193.345 ;
        RECT 88.410 189.605 88.550 193.025 ;
        RECT 91.050 192.490 92.590 192.860 ;
        RECT 91.110 191.665 91.370 191.985 ;
        RECT 88.350 189.285 88.610 189.605 ;
        RECT 91.170 189.265 91.310 191.665 ;
        RECT 91.110 188.945 91.370 189.265 ;
        RECT 86.970 188.265 87.230 188.585 ;
        RECT 90.190 188.265 90.450 188.585 ;
        RECT 88.350 187.585 88.610 187.905 ;
        RECT 87.430 186.225 87.690 186.545 ;
        RECT 85.590 185.605 85.850 185.865 ;
        RECT 85.590 185.545 86.250 185.605 ;
        RECT 85.650 185.465 86.250 185.545 ;
        RECT 86.110 183.825 86.250 185.465 ;
        RECT 87.490 184.165 87.630 186.225 ;
        RECT 87.430 183.845 87.690 184.165 ;
        RECT 86.050 183.505 86.310 183.825 ;
        RECT 86.110 180.765 86.250 183.505 ;
        RECT 88.410 183.145 88.550 187.585 ;
        RECT 88.350 182.825 88.610 183.145 ;
        RECT 88.810 182.825 89.070 183.145 ;
        RECT 89.730 182.825 89.990 183.145 ;
        RECT 86.050 180.445 86.310 180.765 ;
        RECT 86.110 177.705 86.250 180.445 ;
        RECT 87.890 179.425 88.150 179.745 ;
        RECT 87.950 178.045 88.090 179.425 ;
        RECT 87.890 177.725 88.150 178.045 ;
        RECT 86.050 177.385 86.310 177.705 ;
        RECT 86.110 169.545 86.250 177.385 ;
        RECT 88.870 174.645 89.010 182.825 ;
        RECT 89.790 181.105 89.930 182.825 ;
        RECT 89.730 180.785 89.990 181.105 ;
        RECT 89.730 178.405 89.990 178.725 ;
        RECT 88.810 174.325 89.070 174.645 ;
        RECT 89.270 173.985 89.530 174.305 ;
        RECT 89.330 172.945 89.470 173.985 ;
        RECT 89.270 172.625 89.530 172.945 ;
        RECT 89.790 172.265 89.930 178.405 ;
        RECT 89.730 171.945 89.990 172.265 ;
        RECT 87.430 171.265 87.690 171.585 ;
        RECT 89.730 171.265 89.990 171.585 ;
        RECT 87.490 169.885 87.630 171.265 ;
        RECT 87.430 169.565 87.690 169.885 ;
        RECT 86.050 169.225 86.310 169.545 ;
        RECT 86.110 166.825 86.250 169.225 ;
        RECT 86.050 166.505 86.310 166.825 ;
        RECT 86.110 164.105 86.250 166.505 ;
        RECT 88.810 164.125 89.070 164.445 ;
        RECT 86.050 163.785 86.310 164.105 ;
        RECT 85.130 161.405 85.390 161.725 ;
        RECT 84.670 161.065 84.930 161.385 ;
        RECT 76.850 158.685 77.110 159.005 ;
        RECT 77.310 158.685 77.570 159.005 ;
        RECT 76.390 157.665 76.650 157.985 ;
        RECT 75.930 155.965 76.190 156.285 ;
        RECT 75.930 154.945 76.190 155.265 ;
        RECT 75.990 154.245 76.130 154.945 ;
        RECT 75.930 153.925 76.190 154.245 ;
        RECT 75.930 149.845 76.190 150.165 ;
        RECT 75.990 145.745 76.130 149.845 ;
        RECT 75.930 145.425 76.190 145.745 ;
        RECT 75.990 142.685 76.130 145.425 ;
        RECT 75.930 142.365 76.190 142.685 ;
        RECT 75.470 139.985 75.730 140.305 ;
        RECT 75.010 139.645 75.270 139.965 ;
        RECT 74.550 139.305 74.810 139.625 ;
        RECT 76.450 139.285 76.590 157.665 ;
        RECT 76.910 155.945 77.050 158.685 ;
        RECT 81.910 158.005 82.170 158.325 ;
        RECT 77.655 157.130 79.195 157.500 ;
        RECT 80.990 156.645 81.250 156.965 ;
        RECT 81.050 156.285 81.190 156.645 ;
        RECT 81.970 156.285 82.110 158.005 ;
        RECT 84.730 156.965 84.870 161.065 ;
        RECT 86.110 159.685 86.250 163.785 ;
        RECT 88.870 161.385 89.010 164.125 ;
        RECT 88.810 161.065 89.070 161.385 ;
        RECT 87.430 160.385 87.690 160.705 ;
        RECT 86.050 159.365 86.310 159.685 ;
        RECT 87.490 159.345 87.630 160.385 ;
        RECT 87.430 159.025 87.690 159.345 ;
        RECT 84.670 156.645 84.930 156.965 ;
        RECT 80.990 155.965 81.250 156.285 ;
        RECT 81.910 155.965 82.170 156.285 ;
        RECT 76.850 155.625 77.110 155.945 ;
        RECT 76.910 153.565 77.050 155.625 ;
        RECT 76.850 153.245 77.110 153.565 ;
        RECT 77.310 152.905 77.570 153.225 ;
        RECT 76.850 150.185 77.110 150.505 ;
        RECT 77.370 150.245 77.510 152.905 ;
        RECT 77.655 151.690 79.195 152.060 ;
        RECT 81.050 150.845 81.190 155.965 ;
        RECT 81.910 154.945 82.170 155.265 ;
        RECT 81.450 154.155 81.710 154.245 ;
        RECT 81.970 154.155 82.110 154.945 ;
        RECT 81.450 154.015 82.110 154.155 ;
        RECT 81.450 153.925 81.710 154.015 ;
        RECT 81.970 150.845 82.110 154.015 ;
        RECT 85.590 153.585 85.850 153.905 ;
        RECT 85.650 151.525 85.790 153.585 ;
        RECT 89.790 153.565 89.930 171.265 ;
        RECT 90.250 165.125 90.390 188.265 ;
        RECT 91.050 187.050 92.590 187.420 ;
        RECT 93.010 183.565 93.150 196.425 ;
        RECT 93.470 194.445 93.610 196.765 ;
        RECT 94.790 195.745 95.050 196.065 ;
        RECT 93.470 194.305 94.070 194.445 ;
        RECT 93.410 193.365 93.670 193.685 ;
        RECT 93.470 190.625 93.610 193.365 ;
        RECT 93.410 190.305 93.670 190.625 ;
        RECT 93.470 188.585 93.610 190.305 ;
        RECT 93.930 188.585 94.070 194.305 ;
        RECT 94.850 193.345 94.990 195.745 ;
        RECT 95.310 194.365 95.450 199.485 ;
        RECT 96.690 198.785 96.830 201.865 ;
        RECT 99.450 200.485 99.590 202.205 ;
        RECT 99.390 200.165 99.650 200.485 ;
        RECT 100.770 199.145 101.030 199.465 ;
        RECT 99.390 198.805 99.650 199.125 ;
        RECT 96.630 198.640 96.890 198.785 ;
        RECT 96.620 198.270 96.900 198.640 ;
        RECT 95.250 194.045 95.510 194.365 ;
        RECT 99.450 193.345 99.590 198.805 ;
        RECT 100.830 195.045 100.970 199.145 ;
        RECT 102.610 198.465 102.870 198.785 ;
        RECT 102.670 197.425 102.810 198.465 ;
        RECT 102.610 197.105 102.870 197.425 ;
        RECT 104.050 197.085 104.190 204.585 ;
        RECT 104.445 200.650 105.985 201.020 ;
        RECT 103.990 196.765 104.250 197.085 ;
        RECT 100.770 194.725 101.030 195.045 ;
        RECT 94.790 193.025 95.050 193.345 ;
        RECT 98.010 193.025 98.270 193.345 ;
        RECT 99.390 193.025 99.650 193.345 ;
        RECT 93.410 188.265 93.670 188.585 ;
        RECT 93.870 188.265 94.130 188.585 ;
        RECT 93.010 183.425 94.070 183.565 ;
        RECT 90.650 182.825 90.910 183.145 ;
        RECT 93.410 182.885 93.670 183.145 ;
        RECT 93.010 182.825 93.670 182.885 ;
        RECT 90.710 178.725 90.850 182.825 ;
        RECT 93.010 182.745 93.610 182.825 ;
        RECT 91.050 181.610 92.590 181.980 ;
        RECT 90.650 178.405 90.910 178.725 ;
        RECT 93.010 178.045 93.150 182.745 ;
        RECT 93.410 182.145 93.670 182.465 ;
        RECT 93.470 181.105 93.610 182.145 ;
        RECT 93.410 180.785 93.670 181.105 ;
        RECT 93.930 180.165 94.070 183.425 ;
        RECT 94.330 182.825 94.590 183.145 ;
        RECT 94.390 181.445 94.530 182.825 ;
        RECT 94.330 181.125 94.590 181.445 ;
        RECT 93.470 180.025 94.070 180.165 ;
        RECT 92.950 177.725 93.210 178.045 ;
        RECT 91.050 176.170 92.590 176.540 ;
        RECT 92.950 175.345 93.210 175.665 ;
        RECT 92.030 174.325 92.290 174.645 ;
        RECT 90.650 173.985 90.910 174.305 ;
        RECT 90.710 172.265 90.850 173.985 ;
        RECT 92.090 173.285 92.230 174.325 ;
        RECT 91.110 172.965 91.370 173.285 ;
        RECT 92.030 172.965 92.290 173.285 ;
        RECT 90.650 171.945 90.910 172.265 ;
        RECT 91.170 171.495 91.310 172.965 ;
        RECT 92.090 172.265 92.230 172.965 ;
        RECT 92.490 172.625 92.750 172.945 ;
        RECT 92.030 171.945 92.290 172.265 ;
        RECT 92.550 171.925 92.690 172.625 ;
        RECT 92.490 171.605 92.750 171.925 ;
        RECT 90.710 171.355 91.310 171.495 ;
        RECT 90.710 170.225 90.850 171.355 ;
        RECT 91.050 170.730 92.590 171.100 ;
        RECT 93.010 170.565 93.150 175.345 ;
        RECT 92.950 170.245 93.210 170.565 ;
        RECT 90.650 169.905 90.910 170.225 ;
        RECT 92.950 166.505 93.210 166.825 ;
        RECT 90.650 165.825 90.910 166.145 ;
        RECT 90.710 165.125 90.850 165.825 ;
        RECT 91.050 165.290 92.590 165.660 ;
        RECT 90.190 164.805 90.450 165.125 ;
        RECT 90.650 164.805 90.910 165.125 ;
        RECT 90.710 164.445 90.850 164.805 ;
        RECT 90.190 164.125 90.450 164.445 ;
        RECT 90.650 164.125 90.910 164.445 ;
        RECT 90.250 163.425 90.390 164.125 ;
        RECT 90.190 163.105 90.450 163.425 ;
        RECT 90.250 161.385 90.390 163.105 ;
        RECT 90.710 161.385 90.850 164.125 ;
        RECT 93.010 164.105 93.150 166.505 ;
        RECT 93.470 164.445 93.610 180.025 ;
        RECT 94.390 174.305 94.530 181.125 ;
        RECT 94.330 173.985 94.590 174.305 ;
        RECT 94.850 166.825 94.990 193.025 ;
        RECT 95.250 191.325 95.510 191.645 ;
        RECT 95.310 189.605 95.450 191.325 ;
        RECT 95.250 189.285 95.510 189.605 ;
        RECT 98.070 188.585 98.210 193.025 ;
        RECT 98.930 190.985 99.190 191.305 ;
        RECT 98.990 189.605 99.130 190.985 ;
        RECT 98.930 189.285 99.190 189.605 ;
        RECT 98.010 188.265 98.270 188.585 ;
        RECT 98.470 184.865 98.730 185.185 ;
        RECT 95.250 183.165 95.510 183.485 ;
        RECT 94.790 166.505 95.050 166.825 ;
        RECT 93.870 165.825 94.130 166.145 ;
        RECT 94.330 165.825 94.590 166.145 ;
        RECT 93.930 164.445 94.070 165.825 ;
        RECT 94.390 165.125 94.530 165.825 ;
        RECT 94.330 164.805 94.590 165.125 ;
        RECT 94.390 164.445 94.530 164.805 ;
        RECT 94.790 164.465 95.050 164.785 ;
        RECT 93.410 164.125 93.670 164.445 ;
        RECT 93.870 164.125 94.130 164.445 ;
        RECT 94.330 164.125 94.590 164.445 ;
        RECT 92.950 163.785 93.210 164.105 ;
        RECT 93.930 163.765 94.070 164.125 ;
        RECT 93.870 163.445 94.130 163.765 ;
        RECT 93.410 163.105 93.670 163.425 ;
        RECT 90.190 161.065 90.450 161.385 ;
        RECT 90.650 161.065 90.910 161.385 ;
        RECT 92.950 160.385 93.210 160.705 ;
        RECT 91.050 159.850 92.590 160.220 ;
        RECT 91.050 154.410 92.590 154.780 ;
        RECT 89.270 153.245 89.530 153.565 ;
        RECT 89.730 153.245 89.990 153.565 ;
        RECT 87.430 152.905 87.690 153.225 ;
        RECT 87.490 151.525 87.630 152.905 ;
        RECT 85.590 151.205 85.850 151.525 ;
        RECT 87.430 151.205 87.690 151.525 ;
        RECT 80.990 150.525 81.250 150.845 ;
        RECT 81.910 150.525 82.170 150.845 ;
        RECT 77.770 150.245 78.030 150.505 ;
        RECT 77.370 150.185 78.030 150.245 ;
        RECT 76.910 144.385 77.050 150.185 ;
        RECT 77.370 150.105 77.970 150.185 ;
        RECT 77.370 144.975 77.510 150.105 ;
        RECT 81.050 148.805 81.190 150.525 ;
        RECT 86.050 150.185 86.310 150.505 ;
        RECT 82.370 149.505 82.630 149.825 ;
        RECT 80.990 148.485 81.250 148.805 ;
        RECT 77.655 146.250 79.195 146.620 ;
        RECT 81.050 145.405 81.190 148.485 ;
        RECT 82.430 147.445 82.570 149.505 ;
        RECT 82.370 147.125 82.630 147.445 ;
        RECT 80.990 145.085 81.250 145.405 ;
        RECT 77.770 144.975 78.030 145.065 ;
        RECT 77.370 144.835 78.030 144.975 ;
        RECT 77.770 144.745 78.030 144.835 ;
        RECT 76.850 144.065 77.110 144.385 ;
        RECT 76.910 142.005 77.050 144.065 ;
        RECT 77.830 143.365 77.970 144.745 ;
        RECT 77.770 143.045 78.030 143.365 ;
        RECT 77.830 142.685 77.970 143.045 ;
        RECT 77.770 142.365 78.030 142.685 ;
        RECT 81.050 142.345 81.190 145.085 ;
        RECT 82.430 144.725 82.570 147.125 ;
        RECT 86.110 145.065 86.250 150.185 ;
        RECT 86.510 148.145 86.770 148.465 ;
        RECT 86.570 146.085 86.710 148.145 ;
        RECT 89.330 147.785 89.470 153.245 ;
        RECT 93.010 153.225 93.150 160.385 ;
        RECT 93.470 156.285 93.610 163.105 ;
        RECT 93.930 161.725 94.070 163.445 ;
        RECT 94.390 162.405 94.530 164.125 ;
        RECT 94.850 163.765 94.990 164.465 ;
        RECT 94.790 163.445 95.050 163.765 ;
        RECT 94.330 162.085 94.590 162.405 ;
        RECT 93.870 161.405 94.130 161.725 ;
        RECT 94.320 161.550 94.600 161.920 ;
        RECT 94.390 161.385 94.530 161.550 ;
        RECT 94.330 161.065 94.590 161.385 ;
        RECT 95.310 159.005 95.450 183.165 ;
        RECT 98.530 183.145 98.670 184.865 ;
        RECT 97.550 182.825 97.810 183.145 ;
        RECT 98.470 182.825 98.730 183.145 ;
        RECT 97.610 175.235 97.750 182.825 ;
        RECT 98.930 182.145 99.190 182.465 ;
        RECT 98.990 178.045 99.130 182.145 ;
        RECT 98.930 177.725 99.190 178.045 ;
        RECT 98.930 175.235 99.190 175.325 ;
        RECT 97.610 175.095 99.190 175.235 ;
        RECT 97.090 174.665 97.350 174.985 ;
        RECT 96.630 171.265 96.890 171.585 ;
        RECT 96.690 169.885 96.830 171.265 ;
        RECT 97.150 170.565 97.290 174.665 ;
        RECT 98.530 172.265 98.670 175.095 ;
        RECT 98.930 175.005 99.190 175.095 ;
        RECT 98.930 173.985 99.190 174.305 ;
        RECT 98.990 172.265 99.130 173.985 ;
        RECT 98.470 171.945 98.730 172.265 ;
        RECT 98.930 171.945 99.190 172.265 ;
        RECT 97.550 171.265 97.810 171.585 ;
        RECT 97.090 170.245 97.350 170.565 ;
        RECT 96.630 169.565 96.890 169.885 ;
        RECT 97.090 168.545 97.350 168.865 ;
        RECT 97.150 164.445 97.290 168.545 ;
        RECT 97.090 164.125 97.350 164.445 ;
        RECT 96.630 163.785 96.890 164.105 ;
        RECT 95.710 163.105 95.970 163.425 ;
        RECT 95.770 159.005 95.910 163.105 ;
        RECT 96.690 162.405 96.830 163.785 ;
        RECT 96.630 162.085 96.890 162.405 ;
        RECT 95.250 158.685 95.510 159.005 ;
        RECT 95.710 158.685 95.970 159.005 ;
        RECT 93.870 157.665 94.130 157.985 ;
        RECT 94.330 157.665 94.590 157.985 ;
        RECT 97.090 157.665 97.350 157.985 ;
        RECT 93.410 155.965 93.670 156.285 ;
        RECT 93.930 153.905 94.070 157.665 ;
        RECT 94.390 156.625 94.530 157.665 ;
        RECT 94.330 156.305 94.590 156.625 ;
        RECT 96.160 156.110 96.440 156.480 ;
        RECT 95.710 154.945 95.970 155.265 ;
        RECT 93.870 153.585 94.130 153.905 ;
        RECT 92.950 152.905 93.210 153.225 ;
        RECT 90.190 152.225 90.450 152.545 ;
        RECT 90.650 152.225 90.910 152.545 ;
        RECT 88.350 147.465 88.610 147.785 ;
        RECT 89.270 147.465 89.530 147.785 ;
        RECT 88.410 146.085 88.550 147.465 ;
        RECT 86.510 145.765 86.770 146.085 ;
        RECT 88.350 145.765 88.610 146.085 ;
        RECT 86.050 144.745 86.310 145.065 ;
        RECT 82.370 144.405 82.630 144.725 ;
        RECT 83.290 144.065 83.550 144.385 ;
        RECT 83.350 143.025 83.490 144.065 ;
        RECT 83.290 142.705 83.550 143.025 ;
        RECT 80.990 142.025 81.250 142.345 ;
        RECT 76.850 141.685 77.110 142.005 ;
        RECT 77.655 140.810 79.195 141.180 ;
        RECT 83.350 140.645 83.490 142.705 ;
        RECT 88.350 141.345 88.610 141.665 ;
        RECT 83.290 140.325 83.550 140.645 ;
        RECT 88.410 139.965 88.550 141.345 ;
        RECT 89.330 139.965 89.470 147.465 ;
        RECT 88.350 139.645 88.610 139.965 ;
        RECT 89.270 139.645 89.530 139.965 ;
        RECT 76.390 138.965 76.650 139.285 ;
        RECT 86.510 138.965 86.770 139.285 ;
        RECT 75.930 138.625 76.190 138.945 ;
        RECT 75.470 136.585 75.730 136.905 ;
        RECT 73.170 134.885 73.430 135.205 ;
        RECT 74.550 133.865 74.810 134.185 ;
        RECT 75.010 133.865 75.270 134.185 ;
        RECT 74.090 128.085 74.350 128.405 ;
        RECT 74.150 127.045 74.290 128.085 ;
        RECT 74.610 127.045 74.750 133.865 ;
        RECT 75.070 131.465 75.210 133.865 ;
        RECT 75.530 133.505 75.670 136.585 ;
        RECT 75.470 133.185 75.730 133.505 ;
        RECT 75.530 131.805 75.670 133.185 ;
        RECT 75.470 131.485 75.730 131.805 ;
        RECT 75.010 131.145 75.270 131.465 ;
        RECT 75.530 129.765 75.670 131.485 ;
        RECT 75.470 129.445 75.730 129.765 ;
        RECT 74.090 126.725 74.350 127.045 ;
        RECT 74.550 126.725 74.810 127.045 ;
        RECT 72.710 125.025 72.970 125.345 ;
        RECT 72.770 122.965 72.910 125.025 ;
        RECT 72.710 122.645 72.970 122.965 ;
        RECT 72.710 120.605 72.970 120.925 ;
        RECT 74.090 120.605 74.350 120.925 ;
        RECT 72.250 117.545 72.510 117.865 ;
        RECT 70.410 117.205 70.670 117.525 ;
        RECT 66.270 116.865 66.530 117.185 ;
        RECT 69.030 116.865 69.290 117.185 ;
        RECT 64.260 116.330 65.800 116.700 ;
        RECT 66.330 115.825 66.470 116.865 ;
        RECT 69.090 115.825 69.230 116.865 ;
        RECT 66.270 115.505 66.530 115.825 ;
        RECT 67.650 115.505 67.910 115.825 ;
        RECT 69.030 115.505 69.290 115.825 ;
        RECT 61.210 114.825 61.470 115.145 ;
        RECT 64.430 114.825 64.690 115.145 ;
        RECT 61.270 112.675 61.410 114.825 ;
        RECT 64.490 113.445 64.630 114.825 ;
        RECT 64.430 113.125 64.690 113.445 ;
        RECT 64.490 112.765 64.630 113.125 ;
        RECT 61.270 112.535 62.330 112.675 ;
        RECT 59.370 109.725 59.630 110.045 ;
        RECT 62.190 106.285 62.330 112.535 ;
        RECT 64.430 112.445 64.690 112.765 ;
        RECT 64.260 110.890 65.800 111.260 ;
        RECT 67.710 106.285 67.850 115.505 ;
        RECT 72.770 112.085 72.910 120.605 ;
        RECT 73.630 118.115 73.890 118.205 ;
        RECT 74.150 118.115 74.290 120.605 ;
        RECT 73.630 117.975 74.290 118.115 ;
        RECT 73.630 117.885 73.890 117.975 ;
        RECT 73.630 116.865 73.890 117.185 ;
        RECT 73.690 116.165 73.830 116.865 ;
        RECT 73.630 115.845 73.890 116.165 ;
        RECT 73.170 112.445 73.430 112.765 ;
        RECT 72.710 111.765 72.970 112.085 ;
        RECT 73.230 106.285 73.370 112.445 ;
        RECT 74.150 110.045 74.290 117.975 ;
        RECT 75.990 117.865 76.130 138.625 ;
        RECT 86.570 137.925 86.710 138.965 ;
        RECT 86.510 137.605 86.770 137.925 ;
        RECT 80.070 137.265 80.330 137.585 ;
        RECT 77.655 135.370 79.195 135.740 ;
        RECT 76.390 134.205 76.650 134.525 ;
        RECT 76.450 131.125 76.590 134.205 ;
        RECT 80.130 134.185 80.270 137.265 ;
        RECT 81.910 136.925 82.170 137.245 ;
        RECT 80.070 133.865 80.330 134.185 ;
        RECT 76.850 131.145 77.110 131.465 ;
        RECT 76.390 130.805 76.650 131.125 ;
        RECT 76.450 126.025 76.590 130.805 ;
        RECT 76.910 126.365 77.050 131.145 ;
        RECT 80.070 130.465 80.330 130.785 ;
        RECT 77.655 129.930 79.195 130.300 ;
        RECT 80.130 128.745 80.270 130.465 ;
        RECT 81.970 129.085 82.110 136.925 ;
        RECT 84.210 135.905 84.470 136.225 ;
        RECT 84.270 133.845 84.410 135.905 ;
        RECT 89.330 134.525 89.470 139.645 ;
        RECT 89.270 134.205 89.530 134.525 ;
        RECT 86.970 133.865 87.230 134.185 ;
        RECT 84.210 133.525 84.470 133.845 ;
        RECT 82.370 133.185 82.630 133.505 ;
        RECT 82.430 131.805 82.570 133.185 ;
        RECT 87.030 132.485 87.170 133.865 ;
        RECT 86.970 132.165 87.230 132.485 ;
        RECT 82.370 131.485 82.630 131.805 ;
        RECT 88.350 131.145 88.610 131.465 ;
        RECT 81.910 128.765 82.170 129.085 ;
        RECT 80.070 128.425 80.330 128.745 ;
        RECT 79.610 126.725 79.870 127.045 ;
        RECT 76.850 126.045 77.110 126.365 ;
        RECT 76.390 125.705 76.650 126.025 ;
        RECT 76.910 124.325 77.050 126.045 ;
        RECT 77.310 125.025 77.570 125.345 ;
        RECT 76.850 124.005 77.110 124.325 ;
        RECT 77.370 120.925 77.510 125.025 ;
        RECT 77.655 124.490 79.195 124.860 ;
        RECT 79.670 124.325 79.810 126.725 ;
        RECT 81.970 126.365 82.110 128.765 ;
        RECT 88.410 126.705 88.550 131.145 ;
        RECT 89.330 129.765 89.470 134.205 ;
        RECT 89.270 129.445 89.530 129.765 ;
        RECT 88.810 128.600 89.070 128.745 ;
        RECT 88.800 128.230 89.080 128.600 ;
        RECT 88.350 126.385 88.610 126.705 ;
        RECT 81.910 126.045 82.170 126.365 ;
        RECT 89.330 126.025 89.470 129.445 ;
        RECT 89.730 127.745 89.990 128.065 ;
        RECT 89.790 126.705 89.930 127.745 ;
        RECT 89.730 126.385 89.990 126.705 ;
        RECT 89.270 125.705 89.530 126.025 ;
        RECT 82.370 125.025 82.630 125.345 ;
        RECT 86.970 125.025 87.230 125.345 ;
        RECT 79.610 124.005 79.870 124.325 ;
        RECT 79.610 122.985 79.870 123.305 ;
        RECT 79.670 121.605 79.810 122.985 ;
        RECT 82.430 122.965 82.570 125.025 ;
        RECT 85.590 123.325 85.850 123.645 ;
        RECT 82.370 122.645 82.630 122.965 ;
        RECT 79.610 121.285 79.870 121.605 ;
        RECT 77.310 120.605 77.570 120.925 ;
        RECT 77.655 119.050 79.195 119.420 ;
        RECT 75.930 117.545 76.190 117.865 ;
        RECT 76.390 116.865 76.650 117.185 ;
        RECT 79.610 116.865 79.870 117.185 ;
        RECT 76.450 112.765 76.590 116.865 ;
        RECT 77.655 113.610 79.195 113.980 ;
        RECT 79.670 113.445 79.810 116.865 ;
        RECT 84.210 115.845 84.470 116.165 ;
        RECT 80.070 114.825 80.330 115.145 ;
        RECT 79.610 113.125 79.870 113.445 ;
        RECT 76.390 112.445 76.650 112.765 ;
        RECT 79.610 112.445 79.870 112.765 ;
        RECT 78.690 111.765 78.950 112.085 ;
        RECT 78.750 110.725 78.890 111.765 ;
        RECT 78.690 110.405 78.950 110.725 ;
        RECT 74.090 109.725 74.350 110.045 ;
        RECT 77.655 108.170 79.195 108.540 ;
        RECT 79.670 107.405 79.810 112.445 ;
        RECT 80.130 112.425 80.270 114.825 ;
        RECT 80.070 112.105 80.330 112.425 ;
        RECT 78.750 107.265 79.810 107.405 ;
        RECT 78.750 106.285 78.890 107.265 ;
        RECT 84.270 106.285 84.410 115.845 ;
        RECT 85.650 115.145 85.790 123.325 ;
        RECT 87.030 120.925 87.170 125.025 ;
        RECT 89.330 123.725 89.470 125.705 ;
        RECT 89.330 123.645 89.930 123.725 ;
        RECT 89.330 123.585 89.990 123.645 ;
        RECT 89.730 123.325 89.990 123.585 ;
        RECT 89.270 122.985 89.530 123.305 ;
        RECT 89.330 121.605 89.470 122.985 ;
        RECT 89.270 121.285 89.530 121.605 ;
        RECT 86.970 120.605 87.230 120.925 ;
        RECT 88.810 116.865 89.070 117.185 ;
        RECT 88.870 115.825 89.010 116.865 ;
        RECT 90.250 115.825 90.390 152.225 ;
        RECT 90.710 132.485 90.850 152.225 ;
        RECT 91.050 148.970 92.590 149.340 ;
        RECT 92.950 147.125 93.210 147.445 ;
        RECT 91.050 143.530 92.590 143.900 ;
        RECT 93.010 143.365 93.150 147.125 ;
        RECT 93.870 144.745 94.130 145.065 ;
        RECT 92.950 143.045 93.210 143.365 ;
        RECT 93.930 139.965 94.070 144.745 ;
        RECT 93.870 139.645 94.130 139.965 ;
        RECT 91.050 138.090 92.590 138.460 ;
        RECT 93.930 137.245 94.070 139.645 ;
        RECT 93.870 136.925 94.130 137.245 ;
        RECT 93.410 136.585 93.670 136.905 ;
        RECT 93.470 133.925 93.610 136.585 ;
        RECT 93.930 134.525 94.070 136.925 ;
        RECT 94.790 135.905 95.050 136.225 ;
        RECT 94.850 134.525 94.990 135.905 ;
        RECT 93.870 134.205 94.130 134.525 ;
        RECT 94.790 134.205 95.050 134.525 ;
        RECT 94.330 133.925 94.590 134.185 ;
        RECT 93.470 133.865 94.590 133.925 ;
        RECT 93.470 133.785 94.530 133.865 ;
        RECT 91.050 132.650 92.590 133.020 ;
        RECT 90.650 132.165 90.910 132.485 ;
        RECT 94.390 131.465 94.530 133.785 ;
        RECT 94.330 131.145 94.590 131.465 ;
        RECT 91.050 127.210 92.590 127.580 ;
        RECT 94.390 127.045 94.530 131.145 ;
        RECT 95.250 128.425 95.510 128.745 ;
        RECT 95.310 127.045 95.450 128.425 ;
        RECT 94.330 126.725 94.590 127.045 ;
        RECT 95.250 126.725 95.510 127.045 ;
        RECT 94.790 126.045 95.050 126.365 ;
        RECT 94.850 124.325 94.990 126.045 ;
        RECT 94.790 124.005 95.050 124.325 ;
        RECT 91.050 121.770 92.590 122.140 ;
        RECT 93.410 117.885 93.670 118.205 ;
        RECT 91.050 116.330 92.590 116.700 ;
        RECT 86.510 115.505 86.770 115.825 ;
        RECT 88.810 115.505 89.070 115.825 ;
        RECT 90.190 115.505 90.450 115.825 ;
        RECT 85.590 114.825 85.850 115.145 ;
        RECT 85.650 112.085 85.790 114.825 ;
        RECT 86.570 113.445 86.710 115.505 ;
        RECT 93.470 115.485 93.610 117.885 ;
        RECT 95.770 117.865 95.910 154.945 ;
        RECT 96.230 153.565 96.370 156.110 ;
        RECT 96.170 153.245 96.430 153.565 ;
        RECT 96.170 152.565 96.430 152.885 ;
        RECT 96.230 148.805 96.370 152.565 ;
        RECT 96.170 148.485 96.430 148.805 ;
        RECT 96.230 146.085 96.370 148.485 ;
        RECT 96.170 145.765 96.430 146.085 ;
        RECT 96.630 142.705 96.890 143.025 ;
        RECT 96.690 140.645 96.830 142.705 ;
        RECT 96.630 140.325 96.890 140.645 ;
        RECT 97.150 137.925 97.290 157.665 ;
        RECT 97.610 155.945 97.750 171.265 ;
        RECT 99.450 168.865 99.590 193.025 ;
        RECT 104.050 191.645 104.190 196.765 ;
        RECT 104.445 195.210 105.985 195.580 ;
        RECT 103.990 191.325 104.250 191.645 ;
        RECT 110.890 191.325 111.150 191.645 ;
        RECT 102.610 188.945 102.870 189.265 ;
        RECT 100.310 188.265 100.570 188.585 ;
        RECT 100.370 186.205 100.510 188.265 ;
        RECT 101.230 187.585 101.490 187.905 ;
        RECT 101.290 186.205 101.430 187.585 ;
        RECT 100.310 185.885 100.570 186.205 ;
        RECT 101.230 185.885 101.490 186.205 ;
        RECT 100.370 184.165 100.510 185.885 ;
        RECT 102.670 185.865 102.810 188.945 ;
        RECT 103.070 188.265 103.330 188.585 ;
        RECT 103.130 186.545 103.270 188.265 ;
        RECT 103.070 186.225 103.330 186.545 ;
        RECT 102.150 185.545 102.410 185.865 ;
        RECT 102.610 185.545 102.870 185.865 ;
        RECT 102.210 184.165 102.350 185.545 ;
        RECT 100.310 183.845 100.570 184.165 ;
        RECT 102.150 183.845 102.410 184.165 ;
        RECT 101.230 180.105 101.490 180.425 ;
        RECT 100.310 179.425 100.570 179.745 ;
        RECT 99.850 178.065 100.110 178.385 ;
        RECT 99.910 174.645 100.050 178.065 ;
        RECT 100.370 177.365 100.510 179.425 ;
        RECT 101.290 178.725 101.430 180.105 ;
        RECT 101.230 178.405 101.490 178.725 ;
        RECT 101.690 178.405 101.950 178.725 ;
        RECT 101.750 177.705 101.890 178.405 ;
        RECT 101.690 177.385 101.950 177.705 ;
        RECT 100.310 177.045 100.570 177.365 ;
        RECT 100.370 174.985 100.510 177.045 ;
        RECT 101.230 176.705 101.490 177.025 ;
        RECT 100.310 174.665 100.570 174.985 ;
        RECT 99.850 174.325 100.110 174.645 ;
        RECT 99.910 172.605 100.050 174.325 ;
        RECT 100.770 173.985 101.030 174.305 ;
        RECT 99.850 172.285 100.110 172.605 ;
        RECT 99.390 168.545 99.650 168.865 ;
        RECT 98.010 165.825 98.270 166.145 ;
        RECT 97.550 155.625 97.810 155.945 ;
        RECT 98.070 150.845 98.210 165.825 ;
        RECT 99.850 164.125 100.110 164.445 ;
        RECT 99.390 163.105 99.650 163.425 ;
        RECT 99.450 161.725 99.590 163.105 ;
        RECT 99.910 162.065 100.050 164.125 ;
        RECT 100.310 163.105 100.570 163.425 ;
        RECT 99.850 161.745 100.110 162.065 ;
        RECT 99.390 161.405 99.650 161.725 ;
        RECT 98.930 160.725 99.190 161.045 ;
        RECT 98.990 159.685 99.130 160.725 ;
        RECT 98.930 159.365 99.190 159.685 ;
        RECT 98.930 158.685 99.190 159.005 ;
        RECT 99.850 158.685 100.110 159.005 ;
        RECT 98.990 157.985 99.130 158.685 ;
        RECT 98.930 157.665 99.190 157.985 ;
        RECT 98.470 156.645 98.730 156.965 ;
        RECT 98.010 150.525 98.270 150.845 ;
        RECT 98.010 146.785 98.270 147.105 ;
        RECT 98.070 139.625 98.210 146.785 ;
        RECT 98.010 139.305 98.270 139.625 ;
        RECT 97.090 137.605 97.350 137.925 ;
        RECT 98.530 132.485 98.670 156.645 ;
        RECT 99.910 156.285 100.050 158.685 ;
        RECT 99.850 155.965 100.110 156.285 ;
        RECT 98.930 155.285 99.190 155.605 ;
        RECT 98.990 154.245 99.130 155.285 ;
        RECT 99.390 154.945 99.650 155.265 ;
        RECT 98.930 153.925 99.190 154.245 ;
        RECT 98.930 153.245 99.190 153.565 ;
        RECT 98.990 152.545 99.130 153.245 ;
        RECT 98.930 152.225 99.190 152.545 ;
        RECT 99.450 150.505 99.590 154.945 ;
        RECT 99.910 153.225 100.050 155.965 ;
        RECT 99.850 152.905 100.110 153.225 ;
        RECT 100.370 152.285 100.510 163.105 ;
        RECT 99.910 152.145 100.510 152.285 ;
        RECT 99.390 150.185 99.650 150.505 ;
        RECT 98.930 147.465 99.190 147.785 ;
        RECT 98.990 145.405 99.130 147.465 ;
        RECT 98.930 145.085 99.190 145.405 ;
        RECT 99.390 142.025 99.650 142.345 ;
        RECT 99.450 140.645 99.590 142.025 ;
        RECT 99.390 140.325 99.650 140.645 ;
        RECT 99.910 137.925 100.050 152.145 ;
        RECT 100.310 151.205 100.570 151.525 ;
        RECT 99.850 137.605 100.110 137.925 ;
        RECT 99.390 136.925 99.650 137.245 ;
        RECT 99.450 134.185 99.590 136.925 ;
        RECT 99.390 133.865 99.650 134.185 ;
        RECT 100.370 132.485 100.510 151.205 ;
        RECT 100.830 150.505 100.970 173.985 ;
        RECT 101.290 164.445 101.430 176.705 ;
        RECT 101.750 175.325 101.890 177.385 ;
        RECT 102.670 175.325 102.810 185.545 ;
        RECT 103.130 185.185 103.270 186.225 ;
        RECT 103.070 184.865 103.330 185.185 ;
        RECT 104.050 183.485 104.190 191.325 ;
        RECT 109.510 190.305 109.770 190.625 ;
        RECT 104.445 189.770 105.985 190.140 ;
        RECT 109.570 188.245 109.710 190.305 ;
        RECT 110.950 188.925 111.090 191.325 ;
        RECT 110.890 188.605 111.150 188.925 ;
        RECT 109.510 187.925 109.770 188.245 ;
        RECT 106.290 187.585 106.550 187.905 ;
        RECT 104.445 184.330 105.985 184.700 ;
        RECT 106.350 184.165 106.490 187.585 ;
        RECT 106.750 184.865 107.010 185.185 ;
        RECT 106.290 183.845 106.550 184.165 ;
        RECT 103.990 183.165 104.250 183.485 ;
        RECT 106.290 183.165 106.550 183.485 ;
        RECT 104.050 181.445 104.190 183.165 ;
        RECT 105.830 182.485 106.090 182.805 ;
        RECT 103.990 181.125 104.250 181.445 ;
        RECT 103.530 180.785 103.790 181.105 ;
        RECT 103.590 177.025 103.730 180.785 ;
        RECT 103.980 180.590 104.260 180.960 ;
        RECT 103.990 180.445 104.250 180.590 ;
        RECT 105.890 180.085 106.030 182.485 ;
        RECT 105.830 179.765 106.090 180.085 ;
        RECT 104.445 178.890 105.985 179.260 ;
        RECT 106.350 177.705 106.490 183.165 ;
        RECT 106.810 180.765 106.950 184.865 ;
        RECT 107.670 183.165 107.930 183.485 ;
        RECT 106.750 180.445 107.010 180.765 ;
        RECT 107.210 180.445 107.470 180.765 ;
        RECT 107.270 179.745 107.410 180.445 ;
        RECT 107.210 179.425 107.470 179.745 ;
        RECT 106.290 177.385 106.550 177.705 ;
        RECT 103.530 176.705 103.790 177.025 ;
        RECT 103.590 175.325 103.730 176.705 ;
        RECT 106.350 175.665 106.490 177.385 ;
        RECT 107.730 176.085 107.870 183.165 ;
        RECT 110.950 180.765 111.090 188.605 ;
        RECT 114.570 188.265 114.830 188.585 ;
        RECT 113.190 187.925 113.450 188.245 ;
        RECT 113.250 186.885 113.390 187.925 ;
        RECT 113.190 186.565 113.450 186.885 ;
        RECT 114.630 185.865 114.770 188.265 ;
        RECT 113.190 185.545 113.450 185.865 ;
        RECT 114.570 185.545 114.830 185.865 ;
        RECT 116.410 185.545 116.670 185.865 ;
        RECT 113.250 184.165 113.390 185.545 ;
        RECT 113.190 183.845 113.450 184.165 ;
        RECT 108.130 180.445 108.390 180.765 ;
        RECT 110.890 180.445 111.150 180.765 ;
        RECT 112.730 180.445 112.990 180.765 ;
        RECT 108.190 178.725 108.330 180.445 ;
        RECT 108.590 179.425 108.850 179.745 ;
        RECT 111.350 179.425 111.610 179.745 ;
        RECT 108.130 178.405 108.390 178.725 ;
        RECT 108.130 176.705 108.390 177.025 ;
        RECT 107.270 175.945 107.870 176.085 ;
        RECT 106.290 175.345 106.550 175.665 ;
        RECT 101.690 175.005 101.950 175.325 ;
        RECT 102.610 175.005 102.870 175.325 ;
        RECT 103.530 175.005 103.790 175.325 ;
        RECT 103.590 173.285 103.730 175.005 ;
        RECT 107.270 174.985 107.410 175.945 ;
        RECT 108.190 174.985 108.330 176.705 ;
        RECT 107.210 174.665 107.470 174.985 ;
        RECT 108.130 174.665 108.390 174.985 ;
        RECT 104.445 173.450 105.985 173.820 ;
        RECT 101.690 172.965 101.950 173.285 ;
        RECT 103.530 172.965 103.790 173.285 ;
        RECT 101.750 172.265 101.890 172.965 ;
        RECT 108.190 172.265 108.330 174.665 ;
        RECT 101.690 171.945 101.950 172.265 ;
        RECT 108.130 171.945 108.390 172.265 ;
        RECT 107.210 171.605 107.470 171.925 ;
        RECT 107.270 170.565 107.410 171.605 ;
        RECT 107.210 170.245 107.470 170.565 ;
        RECT 106.290 169.565 106.550 169.885 ;
        RECT 104.445 168.010 105.985 168.380 ;
        RECT 101.230 164.125 101.490 164.445 ;
        RECT 105.830 164.355 106.090 164.445 ;
        RECT 106.350 164.355 106.490 169.565 ;
        RECT 105.830 164.215 106.490 164.355 ;
        RECT 105.830 164.125 106.090 164.215 ;
        RECT 104.445 162.570 105.985 162.940 ;
        RECT 103.070 162.085 103.330 162.405 ;
        RECT 102.610 161.065 102.870 161.385 ;
        RECT 102.150 160.725 102.410 161.045 ;
        RECT 102.210 158.665 102.350 160.725 ;
        RECT 102.670 159.005 102.810 161.065 ;
        RECT 102.610 158.685 102.870 159.005 ;
        RECT 102.150 158.345 102.410 158.665 ;
        RECT 102.670 158.325 102.810 158.685 ;
        RECT 102.610 158.005 102.870 158.325 ;
        RECT 102.670 155.945 102.810 158.005 ;
        RECT 102.610 155.625 102.870 155.945 ;
        RECT 102.150 155.285 102.410 155.605 ;
        RECT 102.210 154.245 102.350 155.285 ;
        RECT 102.150 153.925 102.410 154.245 ;
        RECT 101.690 153.245 101.950 153.565 ;
        RECT 100.770 150.185 101.030 150.505 ;
        RECT 101.230 149.505 101.490 149.825 ;
        RECT 98.470 132.165 98.730 132.485 ;
        RECT 100.310 132.165 100.570 132.485 ;
        RECT 98.930 130.805 99.190 131.125 ;
        RECT 96.170 130.465 96.430 130.785 ;
        RECT 96.230 123.305 96.370 130.465 ;
        RECT 98.990 126.705 99.130 130.805 ;
        RECT 100.310 127.745 100.570 128.065 ;
        RECT 98.930 126.385 99.190 126.705 ;
        RECT 98.990 124.325 99.130 126.385 ;
        RECT 99.850 125.025 100.110 125.345 ;
        RECT 98.930 124.005 99.190 124.325 ;
        RECT 96.170 122.985 96.430 123.305 ;
        RECT 99.910 122.965 100.050 125.025 ;
        RECT 100.370 123.645 100.510 127.745 ;
        RECT 100.310 123.325 100.570 123.645 ;
        RECT 99.850 122.645 100.110 122.965 ;
        RECT 101.290 117.865 101.430 149.505 ;
        RECT 101.750 148.465 101.890 153.245 ;
        RECT 102.670 152.545 102.810 155.625 ;
        RECT 102.610 152.225 102.870 152.545 ;
        RECT 101.690 148.145 101.950 148.465 ;
        RECT 102.150 146.785 102.410 147.105 ;
        RECT 102.210 142.685 102.350 146.785 ;
        RECT 102.610 144.745 102.870 145.065 ;
        RECT 102.670 143.365 102.810 144.745 ;
        RECT 102.610 143.045 102.870 143.365 ;
        RECT 102.150 142.365 102.410 142.685 ;
        RECT 102.610 136.925 102.870 137.245 ;
        RECT 102.670 131.805 102.810 136.925 ;
        RECT 103.130 132.485 103.270 162.085 ;
        RECT 106.350 161.385 106.490 164.215 ;
        RECT 107.210 163.105 107.470 163.425 ;
        RECT 104.450 161.065 104.710 161.385 ;
        RECT 106.290 161.065 106.550 161.385 ;
        RECT 103.530 160.385 103.790 160.705 ;
        RECT 103.070 132.165 103.330 132.485 ;
        RECT 102.610 131.485 102.870 131.805 ;
        RECT 103.070 131.145 103.330 131.465 ;
        RECT 103.130 128.745 103.270 131.145 ;
        RECT 103.070 128.425 103.330 128.745 ;
        RECT 103.130 127.045 103.270 128.425 ;
        RECT 103.070 126.725 103.330 127.045 ;
        RECT 103.590 118.205 103.730 160.385 ;
        RECT 104.510 159.005 104.650 161.065 ;
        RECT 104.450 158.915 104.710 159.005 ;
        RECT 104.050 158.775 104.710 158.915 ;
        RECT 104.050 156.285 104.190 158.775 ;
        RECT 104.450 158.685 104.710 158.775 ;
        RECT 104.445 157.130 105.985 157.500 ;
        RECT 103.990 155.965 104.250 156.285 ;
        RECT 104.445 151.690 105.985 152.060 ;
        RECT 106.350 150.505 106.490 161.065 ;
        RECT 107.270 160.705 107.410 163.105 ;
        RECT 108.650 162.065 108.790 179.425 ;
        RECT 111.410 177.365 111.550 179.425 ;
        RECT 111.350 177.045 111.610 177.365 ;
        RECT 112.790 176.005 112.930 180.445 ;
        RECT 115.030 179.425 115.290 179.745 ;
        RECT 115.090 178.045 115.230 179.425 ;
        RECT 115.030 177.725 115.290 178.045 ;
        RECT 116.470 177.705 116.610 185.545 ;
        RECT 116.410 177.385 116.670 177.705 ;
        RECT 112.730 175.685 112.990 176.005 ;
        RECT 116.470 175.665 116.610 177.385 ;
        RECT 116.410 175.345 116.670 175.665 ;
        RECT 115.480 174.470 115.760 174.840 ;
        RECT 115.550 172.265 115.690 174.470 ;
        RECT 116.470 172.605 116.610 175.345 ;
        RECT 135.630 173.380 136.780 174.600 ;
        RECT 116.410 172.285 116.670 172.605 ;
        RECT 112.270 171.945 112.530 172.265 ;
        RECT 115.490 171.945 115.750 172.265 ;
        RECT 109.050 171.265 109.310 171.585 ;
        RECT 109.110 170.225 109.250 171.265 ;
        RECT 112.330 170.565 112.470 171.945 ;
        RECT 113.650 171.605 113.910 171.925 ;
        RECT 112.270 170.245 112.530 170.565 ;
        RECT 109.050 169.905 109.310 170.225 ;
        RECT 113.710 169.545 113.850 171.605 ;
        RECT 113.650 169.225 113.910 169.545 ;
        RECT 113.190 164.805 113.450 165.125 ;
        RECT 108.590 161.745 108.850 162.065 ;
        RECT 107.670 161.405 107.930 161.725 ;
        RECT 107.210 160.385 107.470 160.705 ;
        RECT 107.270 155.945 107.410 160.385 ;
        RECT 107.730 156.285 107.870 161.405 ;
        RECT 112.730 161.065 112.990 161.385 ;
        RECT 108.130 160.385 108.390 160.705 ;
        RECT 110.890 160.385 111.150 160.705 ;
        RECT 108.190 159.345 108.330 160.385 ;
        RECT 110.950 159.345 111.090 160.385 ;
        RECT 108.130 159.025 108.390 159.345 ;
        RECT 110.890 159.025 111.150 159.345 ;
        RECT 109.050 157.665 109.310 157.985 ;
        RECT 107.670 155.965 107.930 156.285 ;
        RECT 107.210 155.625 107.470 155.945 ;
        RECT 107.730 153.225 107.870 155.965 ;
        RECT 108.130 155.285 108.390 155.605 ;
        RECT 108.190 154.245 108.330 155.285 ;
        RECT 109.110 155.265 109.250 157.665 ;
        RECT 112.790 156.965 112.930 161.065 ;
        RECT 112.730 156.645 112.990 156.965 ;
        RECT 111.810 156.305 112.070 156.625 ;
        RECT 109.050 154.945 109.310 155.265 ;
        RECT 109.110 154.245 109.250 154.945 ;
        RECT 108.130 153.925 108.390 154.245 ;
        RECT 109.050 153.925 109.310 154.245 ;
        RECT 107.670 152.905 107.930 153.225 ;
        RECT 107.210 150.865 107.470 151.185 ;
        RECT 106.290 150.185 106.550 150.505 ;
        RECT 105.370 149.505 105.630 149.825 ;
        RECT 105.430 148.465 105.570 149.505 ;
        RECT 105.370 148.145 105.630 148.465 ;
        RECT 106.350 148.125 106.490 150.185 ;
        RECT 106.750 149.845 107.010 150.165 ;
        RECT 106.810 148.805 106.950 149.845 ;
        RECT 106.750 148.485 107.010 148.805 ;
        RECT 106.290 147.805 106.550 148.125 ;
        RECT 107.270 147.785 107.410 150.865 ;
        RECT 107.210 147.465 107.470 147.785 ;
        RECT 104.445 146.250 105.985 146.620 ;
        RECT 104.450 144.745 104.710 145.065 ;
        RECT 104.510 143.025 104.650 144.745 ;
        RECT 107.270 144.385 107.410 147.465 ;
        RECT 107.730 145.405 107.870 152.905 ;
        RECT 108.190 148.805 108.330 153.925 ;
        RECT 109.510 152.905 109.770 153.225 ;
        RECT 108.130 148.485 108.390 148.805 ;
        RECT 107.670 145.085 107.930 145.405 ;
        RECT 108.190 145.065 108.330 148.485 ;
        RECT 108.130 144.745 108.390 145.065 ;
        RECT 107.210 144.065 107.470 144.385 ;
        RECT 104.450 142.705 104.710 143.025 ;
        RECT 104.445 140.810 105.985 141.180 ;
        RECT 109.570 139.625 109.710 152.905 ;
        RECT 109.510 139.305 109.770 139.625 ;
        RECT 110.890 139.305 111.150 139.625 ;
        RECT 106.290 136.585 106.550 136.905 ;
        RECT 104.445 135.370 105.985 135.740 ;
        RECT 106.350 134.185 106.490 136.585 ;
        RECT 107.670 134.205 107.930 134.525 ;
        RECT 109.570 134.425 109.710 139.305 ;
        RECT 109.970 138.625 110.230 138.945 ;
        RECT 110.030 137.585 110.170 138.625 ;
        RECT 109.970 137.265 110.230 137.585 ;
        RECT 110.950 135.205 111.090 139.305 ;
        RECT 110.890 134.885 111.150 135.205 ;
        RECT 109.110 134.285 109.710 134.425 ;
        RECT 106.290 133.865 106.550 134.185 ;
        RECT 104.445 129.930 105.985 130.300 ;
        RECT 107.730 129.425 107.870 134.205 ;
        RECT 107.670 129.105 107.930 129.425 ;
        RECT 106.750 128.085 107.010 128.405 ;
        RECT 104.445 124.490 105.985 124.860 ;
        RECT 106.810 123.305 106.950 128.085 ;
        RECT 107.730 126.025 107.870 129.105 ;
        RECT 109.110 128.745 109.250 134.285 ;
        RECT 110.430 133.185 110.690 133.505 ;
        RECT 110.490 131.465 110.630 133.185 ;
        RECT 110.430 131.145 110.690 131.465 ;
        RECT 110.490 129.085 110.630 131.145 ;
        RECT 110.890 129.105 111.150 129.425 ;
        RECT 110.430 128.765 110.690 129.085 ;
        RECT 109.050 128.425 109.310 128.745 ;
        RECT 107.670 125.705 107.930 126.025 ;
        RECT 109.110 125.685 109.250 128.425 ;
        RECT 109.510 126.385 109.770 126.705 ;
        RECT 109.050 125.365 109.310 125.685 ;
        RECT 109.110 123.305 109.250 125.365 ;
        RECT 109.570 124.325 109.710 126.385 ;
        RECT 109.510 124.005 109.770 124.325 ;
        RECT 110.950 123.305 111.090 129.105 ;
        RECT 106.750 122.985 107.010 123.305 ;
        RECT 109.050 122.985 109.310 123.305 ;
        RECT 110.890 122.985 111.150 123.305 ;
        RECT 104.445 119.050 105.985 119.420 ;
        RECT 103.530 117.885 103.790 118.205 ;
        RECT 106.810 117.865 106.950 122.985 ;
        RECT 111.870 120.925 112.010 156.305 ;
        RECT 113.250 134.425 113.390 164.805 ;
        RECT 113.710 153.565 113.850 169.225 ;
        RECT 116.470 164.105 116.610 172.285 ;
        RECT 133.750 170.070 134.880 172.730 ;
        RECT 135.630 166.640 136.740 173.380 ;
        RECT 135.630 165.420 136.780 166.640 ;
        RECT 114.570 163.785 114.830 164.105 ;
        RECT 116.410 163.785 116.670 164.105 ;
        RECT 114.630 162.405 114.770 163.785 ;
        RECT 114.570 162.085 114.830 162.405 ;
        RECT 114.570 160.385 114.830 160.705 ;
        RECT 114.630 159.005 114.770 160.385 ;
        RECT 116.470 159.005 116.610 163.785 ;
        RECT 114.570 158.685 114.830 159.005 ;
        RECT 116.410 158.685 116.670 159.005 ;
        RECT 113.650 153.245 113.910 153.565 ;
        RECT 116.870 152.225 117.130 152.545 ;
        RECT 116.930 150.505 117.070 152.225 ;
        RECT 113.650 150.185 113.910 150.505 ;
        RECT 115.490 150.185 115.750 150.505 ;
        RECT 116.870 150.185 117.130 150.505 ;
        RECT 113.710 146.085 113.850 150.185 ;
        RECT 115.030 149.505 115.290 149.825 ;
        RECT 115.090 148.125 115.230 149.505 ;
        RECT 115.030 147.805 115.290 148.125 ;
        RECT 115.550 147.785 115.690 150.185 ;
        RECT 115.490 147.465 115.750 147.785 ;
        RECT 113.650 145.765 113.910 146.085 ;
        RECT 115.550 144.725 115.690 147.465 ;
        RECT 115.490 144.405 115.750 144.725 ;
        RECT 113.650 138.625 113.910 138.945 ;
        RECT 113.710 137.245 113.850 138.625 ;
        RECT 113.650 136.925 113.910 137.245 ;
        RECT 115.550 136.905 115.690 144.405 ;
        RECT 135.630 141.200 136.780 141.270 ;
        RECT 135.630 140.180 136.800 141.200 ;
        RECT 132.560 138.140 135.160 140.060 ;
        RECT 115.490 136.585 115.750 136.905 ;
        RECT 113.250 134.285 113.850 134.425 ;
        RECT 112.730 133.185 112.990 133.505 ;
        RECT 112.270 131.825 112.530 132.145 ;
        RECT 112.330 129.765 112.470 131.825 ;
        RECT 112.270 129.445 112.530 129.765 ;
        RECT 112.790 128.745 112.930 133.185 ;
        RECT 112.730 128.425 112.990 128.745 ;
        RECT 113.190 125.705 113.450 126.025 ;
        RECT 113.250 124.325 113.390 125.705 ;
        RECT 113.190 124.005 113.450 124.325 ;
        RECT 113.710 123.045 113.850 134.285 ;
        RECT 115.550 131.805 115.690 136.585 ;
        RECT 135.640 133.320 136.800 140.180 ;
        RECT 115.490 131.485 115.750 131.805 ;
        RECT 114.110 131.145 114.370 131.465 ;
        RECT 114.170 129.765 114.310 131.145 ;
        RECT 114.110 129.445 114.370 129.765 ;
        RECT 115.550 128.065 115.690 131.485 ;
        RECT 115.490 127.745 115.750 128.065 ;
        RECT 115.550 126.365 115.690 127.745 ;
        RECT 115.490 126.045 115.750 126.365 ;
        RECT 113.710 122.905 114.310 123.045 ;
        RECT 111.350 120.605 111.610 120.925 ;
        RECT 111.810 120.605 112.070 120.925 ;
        RECT 107.210 120.265 107.470 120.585 ;
        RECT 107.270 118.885 107.410 120.265 ;
        RECT 108.130 119.585 108.390 119.905 ;
        RECT 107.210 118.565 107.470 118.885 ;
        RECT 108.190 118.205 108.330 119.585 ;
        RECT 108.590 118.565 108.850 118.885 ;
        RECT 108.130 117.885 108.390 118.205 ;
        RECT 95.710 117.545 95.970 117.865 ;
        RECT 101.230 117.545 101.490 117.865 ;
        RECT 106.750 117.545 107.010 117.865 ;
        RECT 98.930 116.865 99.190 117.185 ;
        RECT 100.310 116.865 100.570 117.185 ;
        RECT 102.150 116.865 102.410 117.185 ;
        RECT 103.990 116.865 104.250 117.185 ;
        RECT 93.410 115.165 93.670 115.485 ;
        RECT 90.650 114.145 90.910 114.465 ;
        RECT 86.510 113.125 86.770 113.445 ;
        RECT 89.730 112.105 89.990 112.425 ;
        RECT 85.590 111.765 85.850 112.085 ;
        RECT 85.650 109.705 85.790 111.765 ;
        RECT 88.350 111.425 88.610 111.745 ;
        RECT 88.410 110.385 88.550 111.425 ;
        RECT 89.790 110.725 89.930 112.105 ;
        RECT 89.730 110.405 89.990 110.725 ;
        RECT 90.710 110.385 90.850 114.145 ;
        RECT 93.470 112.425 93.610 115.165 ;
        RECT 93.870 114.145 94.130 114.465 ;
        RECT 93.930 112.425 94.070 114.145 ;
        RECT 98.990 112.765 99.130 116.865 ;
        RECT 100.370 115.825 100.510 116.865 ;
        RECT 102.210 115.825 102.350 116.865 ;
        RECT 100.310 115.505 100.570 115.825 ;
        RECT 102.150 115.505 102.410 115.825 ;
        RECT 100.770 114.825 101.030 115.145 ;
        RECT 103.070 114.825 103.330 115.145 ;
        RECT 98.930 112.445 99.190 112.765 ;
        RECT 93.410 112.105 93.670 112.425 ;
        RECT 93.870 112.105 94.130 112.425 ;
        RECT 95.250 111.765 95.510 112.085 ;
        RECT 91.050 110.890 92.590 111.260 ;
        RECT 88.350 110.065 88.610 110.385 ;
        RECT 90.650 110.065 90.910 110.385 ;
        RECT 85.590 109.385 85.850 109.705 ;
        RECT 89.730 108.705 89.990 109.025 ;
        RECT 89.790 106.285 89.930 108.705 ;
        RECT 95.310 106.285 95.450 111.765 ;
        RECT 100.830 106.285 100.970 114.825 ;
        RECT 103.130 112.765 103.270 114.825 ;
        RECT 103.070 112.445 103.330 112.765 ;
        RECT 104.050 112.085 104.190 116.865 ;
        RECT 106.810 115.145 106.950 117.545 ;
        RECT 106.750 114.825 107.010 115.145 ;
        RECT 104.445 113.610 105.985 113.980 ;
        RECT 106.290 112.445 106.550 112.765 ;
        RECT 103.990 111.765 104.250 112.085 ;
        RECT 104.445 108.170 105.985 108.540 ;
        RECT 106.350 106.285 106.490 112.445 ;
        RECT 108.650 110.045 108.790 118.565 ;
        RECT 111.410 117.525 111.550 120.605 ;
        RECT 111.350 117.205 111.610 117.525 ;
        RECT 112.270 116.865 112.530 117.185 ;
        RECT 110.430 115.505 110.690 115.825 ;
        RECT 110.490 110.725 110.630 115.505 ;
        RECT 111.810 114.825 112.070 115.145 ;
        RECT 110.430 110.405 110.690 110.725 ;
        RECT 108.590 109.725 108.850 110.045 ;
        RECT 111.870 106.285 112.010 114.825 ;
        RECT 112.330 112.765 112.470 116.865 ;
        RECT 112.270 112.445 112.530 112.765 ;
        RECT 114.170 112.425 114.310 122.905 ;
        RECT 115.030 115.505 115.290 115.825 ;
        RECT 115.090 113.445 115.230 115.505 ;
        RECT 115.550 115.145 115.690 126.045 ;
        RECT 115.950 122.305 116.210 122.625 ;
        RECT 116.010 121.605 116.150 122.305 ;
        RECT 115.950 121.285 116.210 121.605 ;
        RECT 116.870 120.605 117.130 120.925 ;
        RECT 116.930 120.440 117.070 120.605 ;
        RECT 116.860 120.070 117.140 120.440 ;
        RECT 117.330 117.205 117.590 117.525 ;
        RECT 115.490 114.825 115.750 115.145 ;
        RECT 115.030 113.125 115.290 113.445 ;
        RECT 115.550 112.765 115.690 114.825 ;
        RECT 115.490 112.445 115.750 112.765 ;
        RECT 114.110 112.105 114.370 112.425 ;
        RECT 117.390 106.285 117.530 117.205 ;
        RECT 12.440 104.285 12.720 106.285 ;
        RECT 17.960 104.285 18.240 106.285 ;
        RECT 23.480 104.285 23.760 106.285 ;
        RECT 29.000 104.285 29.280 106.285 ;
        RECT 34.520 104.285 34.800 106.285 ;
        RECT 40.040 104.285 40.320 106.285 ;
        RECT 45.560 104.285 45.840 106.285 ;
        RECT 51.080 104.285 51.360 106.285 ;
        RECT 56.600 104.285 56.880 106.285 ;
        RECT 62.120 104.285 62.400 106.285 ;
        RECT 67.640 104.285 67.920 106.285 ;
        RECT 73.160 104.285 73.440 106.285 ;
        RECT 78.680 104.285 78.960 106.285 ;
        RECT 84.200 104.285 84.480 106.285 ;
        RECT 89.720 104.285 90.000 106.285 ;
        RECT 95.240 104.285 95.520 106.285 ;
        RECT 100.760 104.285 101.040 106.285 ;
        RECT 106.280 104.285 106.560 106.285 ;
        RECT 111.800 104.285 112.080 106.285 ;
        RECT 117.320 104.285 117.600 106.285 ;
        RECT 129.750 105.580 133.160 106.650 ;
        RECT 13.920 85.550 15.140 89.420 ;
        RECT 19.910 85.980 21.130 89.850 ;
        RECT 67.730 89.640 68.670 89.840 ;
        RECT 25.730 85.120 26.950 88.990 ;
        RECT 31.780 85.510 33.000 89.380 ;
        RECT 37.750 88.780 38.970 89.290 ;
        RECT 37.680 88.620 38.970 88.780 ;
        RECT 43.810 88.630 45.030 89.530 ;
        RECT 49.740 88.640 50.960 89.040 ;
        RECT 37.680 86.810 39.070 88.620 ;
        RECT 37.750 85.420 38.970 86.810 ;
        RECT 43.810 86.720 45.140 88.630 ;
        RECT 49.740 86.920 51.010 88.640 ;
        RECT 43.810 85.660 45.030 86.720 ;
        RECT 49.740 85.170 50.960 86.920 ;
        RECT 55.530 85.320 56.750 89.190 ;
        RECT 61.720 88.640 62.940 88.870 ;
        RECT 61.720 86.600 63.130 88.640 ;
        RECT 61.720 85.000 62.940 86.600 ;
        RECT 67.580 85.770 68.800 89.640 ;
        RECT 73.850 84.290 75.070 88.160 ;
        RECT 79.730 84.310 80.950 88.180 ;
        RECT 74.090 80.440 74.370 84.290 ;
        RECT 20.140 80.160 74.370 80.440 ;
        RECT 20.140 75.650 20.420 80.160 ;
        RECT 80.070 79.800 80.350 84.310 ;
        RECT 85.470 84.100 86.690 87.970 ;
        RECT 91.460 84.500 92.680 88.320 ;
        RECT 97.600 84.630 98.820 88.240 ;
        RECT 103.650 84.740 104.870 88.610 ;
        RECT 109.620 85.420 110.840 89.290 ;
        RECT 115.740 85.700 116.960 89.570 ;
        RECT 121.520 85.700 122.740 89.570 ;
        RECT 31.380 79.520 80.350 79.800 ;
        RECT 31.380 75.850 31.660 79.520 ;
        RECT 86.050 79.170 86.330 84.100 ;
        RECT 42.510 78.890 86.330 79.170 ;
        RECT 3.960 71.320 6.050 73.240 ;
        RECT 19.330 73.120 21.890 75.650 ;
        RECT 28.185 73.180 30.255 74.460 ;
        RECT 30.670 73.320 33.230 75.850 ;
        RECT 42.510 75.750 42.790 78.890 ;
        RECT 92.030 78.570 92.310 84.500 ;
        RECT 53.830 78.290 92.310 78.570 ;
        RECT 53.830 75.820 54.110 78.290 ;
        RECT 98.010 77.990 98.290 84.630 ;
        RECT 64.900 77.710 98.290 77.990 ;
        RECT 19.005 71.800 19.865 72.640 ;
        RECT 15.560 68.610 16.990 71.210 ;
        RECT 19.305 68.570 19.845 71.800 ;
        RECT 20.145 70.600 20.555 73.120 ;
        RECT 30.205 71.810 31.065 72.650 ;
        RECT 19.325 47.770 19.825 68.570 ;
        RECT 20.165 49.090 20.555 70.600 ;
        RECT 20.955 70.010 21.845 70.740 ;
        RECT 21.055 65.190 21.315 70.010 ;
        RECT 22.695 68.620 25.405 69.470 ;
        RECT 22.895 65.840 24.825 68.620 ;
        RECT 30.505 68.580 31.045 71.810 ;
        RECT 31.345 70.610 31.755 73.320 ;
        RECT 39.475 73.150 41.545 74.430 ;
        RECT 41.910 73.220 44.470 75.750 ;
        RECT 41.425 71.780 42.285 72.620 ;
        RECT 27.795 67.130 28.915 67.810 ;
        RECT 28.075 65.850 28.745 67.130 ;
        RECT 21.455 65.460 26.505 65.840 ;
        RECT 27.865 65.440 28.915 65.850 ;
        RECT 21.055 63.640 21.435 65.190 ;
        RECT 21.175 55.800 21.435 63.640 ;
        RECT 26.485 63.200 26.755 65.240 ;
        RECT 27.615 63.200 27.885 65.200 ;
        RECT 26.485 56.510 27.885 63.200 ;
        RECT 21.085 55.290 21.445 55.800 ;
        RECT 21.065 54.860 21.445 55.290 ;
        RECT 26.485 55.190 26.755 56.510 ;
        RECT 27.615 55.150 27.885 56.510 ;
        RECT 28.885 55.260 29.205 65.190 ;
        RECT 28.885 55.200 29.215 55.260 ;
        RECT 21.065 54.580 21.315 54.860 ;
        RECT 20.865 54.180 25.505 54.580 ;
        RECT 26.405 54.290 27.535 54.300 ;
        RECT 28.895 54.290 29.215 55.200 ;
        RECT 21.065 52.060 21.315 54.180 ;
        RECT 25.765 53.490 26.125 54.110 ;
        RECT 25.845 52.610 26.105 53.490 ;
        RECT 26.385 53.240 29.215 54.290 ;
        RECT 25.675 52.230 26.205 52.610 ;
        RECT 21.065 51.970 21.565 52.060 ;
        RECT 21.055 51.240 21.565 51.970 ;
        RECT 21.295 50.240 21.565 51.240 ;
        RECT 22.205 50.990 22.475 51.940 ;
        RECT 22.205 50.840 22.675 50.990 ;
        RECT 22.205 50.160 22.765 50.840 ;
        RECT 22.285 50.150 22.765 50.160 ;
        RECT 21.575 49.620 22.195 49.980 ;
        RECT 21.615 49.090 22.045 49.620 ;
        RECT 20.165 48.670 22.045 49.090 ;
        RECT 22.535 48.960 22.765 50.150 ;
        RECT 21.615 47.800 22.045 48.670 ;
        RECT 22.455 48.360 22.835 48.960 ;
        RECT 19.325 47.060 20.015 47.770 ;
        RECT 21.435 47.440 22.055 47.800 ;
        RECT 21.135 47.060 21.425 47.250 ;
        RECT 19.325 46.620 21.425 47.060 ;
        RECT 19.325 46.600 20.015 46.620 ;
        RECT 21.135 46.380 21.425 46.620 ;
        RECT 22.055 46.990 22.325 47.240 ;
        RECT 22.535 46.990 22.765 48.360 ;
        RECT 25.355 47.010 25.685 52.030 ;
        RECT 26.405 52.020 27.535 53.240 ;
        RECT 28.895 53.220 29.215 53.240 ;
        RECT 22.055 46.880 22.765 46.990 ;
        RECT 25.345 46.960 25.685 47.010 ;
        RECT 26.235 47.780 27.615 52.020 ;
        RECT 22.055 46.570 22.715 46.880 ;
        RECT 22.055 46.400 22.325 46.570 ;
        RECT 25.345 45.000 25.625 46.960 ;
        RECT 26.235 46.920 26.535 47.780 ;
        RECT 27.315 46.920 27.615 47.780 ;
        RECT 28.165 46.920 28.495 51.990 ;
        RECT 27.565 46.380 28.045 46.760 ;
        RECT 27.665 45.760 27.915 46.380 ;
        RECT 27.565 45.160 27.945 45.760 ;
        RECT 24.825 44.230 25.925 45.000 ;
        RECT 28.215 44.930 28.495 46.920 ;
        RECT 30.525 47.780 31.025 68.580 ;
        RECT 31.365 49.100 31.755 70.610 ;
        RECT 32.155 70.020 33.045 70.750 ;
        RECT 32.255 65.200 32.515 70.020 ;
        RECT 33.895 68.630 36.605 69.480 ;
        RECT 34.095 65.850 36.025 68.630 ;
        RECT 41.725 68.550 42.265 71.780 ;
        RECT 42.565 70.580 42.975 73.220 ;
        RECT 50.055 73.090 52.125 74.370 ;
        RECT 53.150 73.290 55.710 75.820 ;
        RECT 64.900 75.810 65.180 77.710 ;
        RECT 103.990 77.230 104.270 84.740 ;
        RECT 76.140 76.950 104.270 77.230 ;
        RECT 52.675 71.760 53.535 72.600 ;
        RECT 38.995 67.140 40.115 67.820 ;
        RECT 39.275 65.860 39.945 67.140 ;
        RECT 32.655 65.470 37.705 65.850 ;
        RECT 39.065 65.450 40.115 65.860 ;
        RECT 32.255 63.650 32.635 65.200 ;
        RECT 32.375 55.810 32.635 63.650 ;
        RECT 37.685 63.210 37.955 65.250 ;
        RECT 38.815 63.210 39.085 65.210 ;
        RECT 37.685 56.520 39.085 63.210 ;
        RECT 32.285 55.300 32.645 55.810 ;
        RECT 32.265 54.870 32.645 55.300 ;
        RECT 37.685 55.200 37.955 56.520 ;
        RECT 38.815 55.160 39.085 56.520 ;
        RECT 40.085 55.270 40.405 65.200 ;
        RECT 40.085 55.210 40.415 55.270 ;
        RECT 32.265 54.590 32.515 54.870 ;
        RECT 32.065 54.190 36.705 54.590 ;
        RECT 37.605 54.300 38.735 54.310 ;
        RECT 40.095 54.300 40.415 55.210 ;
        RECT 32.265 52.070 32.515 54.190 ;
        RECT 36.965 53.500 37.325 54.120 ;
        RECT 37.045 52.620 37.305 53.500 ;
        RECT 37.585 53.250 40.415 54.300 ;
        RECT 36.875 52.240 37.405 52.620 ;
        RECT 32.265 51.980 32.765 52.070 ;
        RECT 32.255 51.250 32.765 51.980 ;
        RECT 32.495 50.250 32.765 51.250 ;
        RECT 33.405 51.000 33.675 51.950 ;
        RECT 33.405 50.850 33.875 51.000 ;
        RECT 33.405 50.170 33.965 50.850 ;
        RECT 33.485 50.160 33.965 50.170 ;
        RECT 32.775 49.630 33.395 49.990 ;
        RECT 32.815 49.100 33.245 49.630 ;
        RECT 31.365 48.680 33.245 49.100 ;
        RECT 33.735 48.970 33.965 50.160 ;
        RECT 32.815 47.810 33.245 48.680 ;
        RECT 33.655 48.370 34.035 48.970 ;
        RECT 30.525 47.070 31.215 47.780 ;
        RECT 32.635 47.450 33.255 47.810 ;
        RECT 32.335 47.070 32.625 47.260 ;
        RECT 30.525 46.630 32.625 47.070 ;
        RECT 30.525 46.610 31.215 46.630 ;
        RECT 32.335 46.390 32.625 46.630 ;
        RECT 33.255 47.000 33.525 47.250 ;
        RECT 33.735 47.000 33.965 48.370 ;
        RECT 36.555 47.020 36.885 52.040 ;
        RECT 37.605 52.030 38.735 53.250 ;
        RECT 40.095 53.230 40.415 53.250 ;
        RECT 33.255 46.890 33.965 47.000 ;
        RECT 36.545 46.970 36.885 47.020 ;
        RECT 37.435 47.790 38.815 52.030 ;
        RECT 33.255 46.580 33.915 46.890 ;
        RECT 33.255 46.410 33.525 46.580 ;
        RECT 36.545 45.010 36.825 46.970 ;
        RECT 37.435 46.930 37.735 47.790 ;
        RECT 38.515 46.930 38.815 47.790 ;
        RECT 39.365 46.930 39.695 52.000 ;
        RECT 38.765 46.390 39.245 46.770 ;
        RECT 38.865 45.770 39.115 46.390 ;
        RECT 38.765 45.170 39.145 45.770 ;
        RECT 28.215 43.200 28.515 44.930 ;
        RECT 36.025 44.240 37.125 45.010 ;
        RECT 39.415 44.940 39.695 46.930 ;
        RECT 41.745 47.750 42.245 68.550 ;
        RECT 42.585 49.070 42.975 70.580 ;
        RECT 43.375 69.990 44.265 70.720 ;
        RECT 43.475 65.170 43.735 69.990 ;
        RECT 45.115 68.600 47.825 69.450 ;
        RECT 45.315 65.820 47.245 68.600 ;
        RECT 52.975 68.530 53.515 71.760 ;
        RECT 53.815 70.560 54.225 73.290 ;
        RECT 61.475 73.120 63.545 74.400 ;
        RECT 64.400 73.280 66.960 75.810 ;
        RECT 76.140 75.740 76.420 76.950 ;
        RECT 109.970 76.610 110.250 85.420 ;
        RECT 87.580 76.330 110.250 76.610 ;
        RECT 87.580 75.760 87.860 76.330 ;
        RECT 115.950 76.030 116.230 85.700 ;
        RECT 98.850 75.840 116.230 76.030 ;
        RECT 63.895 71.750 64.755 72.590 ;
        RECT 50.215 67.110 51.335 67.790 ;
        RECT 50.495 65.830 51.165 67.110 ;
        RECT 43.875 65.440 48.925 65.820 ;
        RECT 50.285 65.420 51.335 65.830 ;
        RECT 43.475 63.620 43.855 65.170 ;
        RECT 43.595 55.780 43.855 63.620 ;
        RECT 48.905 63.180 49.175 65.220 ;
        RECT 50.035 63.180 50.305 65.180 ;
        RECT 48.905 56.490 50.305 63.180 ;
        RECT 43.505 55.270 43.865 55.780 ;
        RECT 43.485 54.840 43.865 55.270 ;
        RECT 48.905 55.170 49.175 56.490 ;
        RECT 50.035 55.130 50.305 56.490 ;
        RECT 51.305 55.240 51.625 65.170 ;
        RECT 51.305 55.180 51.635 55.240 ;
        RECT 43.485 54.560 43.735 54.840 ;
        RECT 43.285 54.160 47.925 54.560 ;
        RECT 48.825 54.270 49.955 54.280 ;
        RECT 51.315 54.270 51.635 55.180 ;
        RECT 43.485 52.040 43.735 54.160 ;
        RECT 48.185 53.470 48.545 54.090 ;
        RECT 48.265 52.590 48.525 53.470 ;
        RECT 48.805 53.220 51.635 54.270 ;
        RECT 48.095 52.210 48.625 52.590 ;
        RECT 43.485 51.950 43.985 52.040 ;
        RECT 43.475 51.220 43.985 51.950 ;
        RECT 43.715 50.220 43.985 51.220 ;
        RECT 44.625 50.970 44.895 51.920 ;
        RECT 44.625 50.820 45.095 50.970 ;
        RECT 44.625 50.140 45.185 50.820 ;
        RECT 44.705 50.130 45.185 50.140 ;
        RECT 43.995 49.600 44.615 49.960 ;
        RECT 44.035 49.070 44.465 49.600 ;
        RECT 42.585 48.650 44.465 49.070 ;
        RECT 44.955 48.940 45.185 50.130 ;
        RECT 44.035 47.780 44.465 48.650 ;
        RECT 44.875 48.340 45.255 48.940 ;
        RECT 41.745 47.040 42.435 47.750 ;
        RECT 43.855 47.420 44.475 47.780 ;
        RECT 43.555 47.040 43.845 47.230 ;
        RECT 41.745 46.600 43.845 47.040 ;
        RECT 41.745 46.580 42.435 46.600 ;
        RECT 43.555 46.360 43.845 46.600 ;
        RECT 44.475 46.970 44.745 47.220 ;
        RECT 44.955 46.970 45.185 48.340 ;
        RECT 47.775 46.990 48.105 52.010 ;
        RECT 48.825 52.000 49.955 53.220 ;
        RECT 51.315 53.200 51.635 53.220 ;
        RECT 44.475 46.860 45.185 46.970 ;
        RECT 47.765 46.940 48.105 46.990 ;
        RECT 48.655 47.760 50.035 52.000 ;
        RECT 44.475 46.550 45.135 46.860 ;
        RECT 44.475 46.380 44.745 46.550 ;
        RECT 47.765 44.980 48.045 46.940 ;
        RECT 48.655 46.900 48.955 47.760 ;
        RECT 49.735 46.900 50.035 47.760 ;
        RECT 50.585 46.900 50.915 51.970 ;
        RECT 49.985 46.360 50.465 46.740 ;
        RECT 50.085 45.740 50.335 46.360 ;
        RECT 49.985 45.140 50.365 45.740 ;
        RECT 39.415 43.210 39.715 44.940 ;
        RECT 47.245 44.210 48.345 44.980 ;
        RECT 50.635 44.910 50.915 46.900 ;
        RECT 52.995 47.730 53.495 68.530 ;
        RECT 53.835 49.050 54.225 70.560 ;
        RECT 54.625 69.970 55.515 70.700 ;
        RECT 54.725 65.150 54.985 69.970 ;
        RECT 56.365 68.580 59.075 69.430 ;
        RECT 56.565 65.800 58.495 68.580 ;
        RECT 64.195 68.520 64.735 71.750 ;
        RECT 65.035 70.550 65.445 73.280 ;
        RECT 72.585 73.130 74.655 74.410 ;
        RECT 75.550 73.210 78.110 75.740 ;
        RECT 75.135 71.740 75.995 72.580 ;
        RECT 61.465 67.090 62.585 67.770 ;
        RECT 61.745 65.810 62.415 67.090 ;
        RECT 55.125 65.420 60.175 65.800 ;
        RECT 61.535 65.400 62.585 65.810 ;
        RECT 54.725 63.600 55.105 65.150 ;
        RECT 54.845 55.760 55.105 63.600 ;
        RECT 60.155 63.160 60.425 65.200 ;
        RECT 61.285 63.160 61.555 65.160 ;
        RECT 60.155 56.470 61.555 63.160 ;
        RECT 54.755 55.250 55.115 55.760 ;
        RECT 54.735 54.820 55.115 55.250 ;
        RECT 60.155 55.150 60.425 56.470 ;
        RECT 61.285 55.110 61.555 56.470 ;
        RECT 62.555 55.220 62.875 65.150 ;
        RECT 62.555 55.160 62.885 55.220 ;
        RECT 54.735 54.540 54.985 54.820 ;
        RECT 54.535 54.140 59.175 54.540 ;
        RECT 60.075 54.250 61.205 54.260 ;
        RECT 62.565 54.250 62.885 55.160 ;
        RECT 54.735 52.020 54.985 54.140 ;
        RECT 59.435 53.450 59.795 54.070 ;
        RECT 59.515 52.570 59.775 53.450 ;
        RECT 60.055 53.200 62.885 54.250 ;
        RECT 59.345 52.190 59.875 52.570 ;
        RECT 54.735 51.930 55.235 52.020 ;
        RECT 54.725 51.200 55.235 51.930 ;
        RECT 54.965 50.200 55.235 51.200 ;
        RECT 55.875 50.950 56.145 51.900 ;
        RECT 55.875 50.800 56.345 50.950 ;
        RECT 55.875 50.120 56.435 50.800 ;
        RECT 55.955 50.110 56.435 50.120 ;
        RECT 55.245 49.580 55.865 49.940 ;
        RECT 55.285 49.050 55.715 49.580 ;
        RECT 53.835 48.630 55.715 49.050 ;
        RECT 56.205 48.920 56.435 50.110 ;
        RECT 55.285 47.760 55.715 48.630 ;
        RECT 56.125 48.320 56.505 48.920 ;
        RECT 52.995 47.020 53.685 47.730 ;
        RECT 55.105 47.400 55.725 47.760 ;
        RECT 54.805 47.020 55.095 47.210 ;
        RECT 52.995 46.580 55.095 47.020 ;
        RECT 52.995 46.560 53.685 46.580 ;
        RECT 54.805 46.340 55.095 46.580 ;
        RECT 55.725 46.950 55.995 47.200 ;
        RECT 56.205 46.950 56.435 48.320 ;
        RECT 59.025 46.970 59.355 51.990 ;
        RECT 60.075 51.980 61.205 53.200 ;
        RECT 62.565 53.180 62.885 53.200 ;
        RECT 55.725 46.840 56.435 46.950 ;
        RECT 59.015 46.920 59.355 46.970 ;
        RECT 59.905 47.740 61.285 51.980 ;
        RECT 55.725 46.530 56.385 46.840 ;
        RECT 55.725 46.360 55.995 46.530 ;
        RECT 59.015 44.960 59.295 46.920 ;
        RECT 59.905 46.880 60.205 47.740 ;
        RECT 60.985 46.880 61.285 47.740 ;
        RECT 61.835 46.880 62.165 51.950 ;
        RECT 61.235 46.340 61.715 46.720 ;
        RECT 61.335 45.720 61.585 46.340 ;
        RECT 61.235 45.120 61.615 45.720 ;
        RECT 19.865 42.210 21.245 42.780 ;
        RECT 27.495 42.630 28.875 43.200 ;
        RECT 31.145 42.210 32.525 42.780 ;
        RECT 38.695 42.640 40.075 43.210 ;
        RECT 50.635 43.180 50.935 44.910 ;
        RECT 58.495 44.190 59.595 44.960 ;
        RECT 61.885 44.890 62.165 46.880 ;
        RECT 64.215 47.720 64.715 68.520 ;
        RECT 65.055 49.040 65.445 70.550 ;
        RECT 65.845 69.960 66.735 70.690 ;
        RECT 65.945 65.140 66.205 69.960 ;
        RECT 67.585 68.570 70.295 69.420 ;
        RECT 67.785 65.790 69.715 68.570 ;
        RECT 75.435 68.510 75.975 71.740 ;
        RECT 76.275 70.540 76.685 73.210 ;
        RECT 83.855 73.120 85.925 74.400 ;
        RECT 86.850 73.230 89.410 75.760 ;
        RECT 98.150 75.750 116.230 75.840 ;
        RECT 86.385 71.750 87.245 72.590 ;
        RECT 72.685 67.080 73.805 67.760 ;
        RECT 72.965 65.800 73.635 67.080 ;
        RECT 66.345 65.410 71.395 65.790 ;
        RECT 72.755 65.390 73.805 65.800 ;
        RECT 65.945 63.590 66.325 65.140 ;
        RECT 66.065 55.750 66.325 63.590 ;
        RECT 71.375 63.150 71.645 65.190 ;
        RECT 72.505 63.150 72.775 65.150 ;
        RECT 71.375 56.460 72.775 63.150 ;
        RECT 65.975 55.240 66.335 55.750 ;
        RECT 65.955 54.810 66.335 55.240 ;
        RECT 71.375 55.140 71.645 56.460 ;
        RECT 72.505 55.100 72.775 56.460 ;
        RECT 73.775 55.210 74.095 65.140 ;
        RECT 73.775 55.150 74.105 55.210 ;
        RECT 65.955 54.530 66.205 54.810 ;
        RECT 65.755 54.130 70.395 54.530 ;
        RECT 71.295 54.240 72.425 54.250 ;
        RECT 73.785 54.240 74.105 55.150 ;
        RECT 65.955 52.010 66.205 54.130 ;
        RECT 70.655 53.440 71.015 54.060 ;
        RECT 70.735 52.560 70.995 53.440 ;
        RECT 71.275 53.190 74.105 54.240 ;
        RECT 70.565 52.180 71.095 52.560 ;
        RECT 65.955 51.920 66.455 52.010 ;
        RECT 65.945 51.190 66.455 51.920 ;
        RECT 66.185 50.190 66.455 51.190 ;
        RECT 67.095 50.940 67.365 51.890 ;
        RECT 67.095 50.790 67.565 50.940 ;
        RECT 67.095 50.110 67.655 50.790 ;
        RECT 67.175 50.100 67.655 50.110 ;
        RECT 66.465 49.570 67.085 49.930 ;
        RECT 66.505 49.040 66.935 49.570 ;
        RECT 65.055 48.620 66.935 49.040 ;
        RECT 67.425 48.910 67.655 50.100 ;
        RECT 66.505 47.750 66.935 48.620 ;
        RECT 67.345 48.310 67.725 48.910 ;
        RECT 64.215 47.010 64.905 47.720 ;
        RECT 66.325 47.390 66.945 47.750 ;
        RECT 66.025 47.010 66.315 47.200 ;
        RECT 64.215 46.570 66.315 47.010 ;
        RECT 64.215 46.550 64.905 46.570 ;
        RECT 66.025 46.330 66.315 46.570 ;
        RECT 66.945 46.940 67.215 47.190 ;
        RECT 67.425 46.940 67.655 48.310 ;
        RECT 70.245 46.960 70.575 51.980 ;
        RECT 71.295 51.970 72.425 53.190 ;
        RECT 73.785 53.170 74.105 53.190 ;
        RECT 66.945 46.830 67.655 46.940 ;
        RECT 70.235 46.910 70.575 46.960 ;
        RECT 71.125 47.730 72.505 51.970 ;
        RECT 66.945 46.520 67.605 46.830 ;
        RECT 66.945 46.350 67.215 46.520 ;
        RECT 70.235 44.950 70.515 46.910 ;
        RECT 71.125 46.870 71.425 47.730 ;
        RECT 72.205 46.870 72.505 47.730 ;
        RECT 73.055 46.870 73.385 51.940 ;
        RECT 72.455 46.330 72.935 46.710 ;
        RECT 72.555 45.710 72.805 46.330 ;
        RECT 72.455 45.110 72.835 45.710 ;
        RECT 20.225 40.480 20.525 42.210 ;
        RECT 20.245 38.490 20.525 40.480 ;
        RECT 22.815 40.410 23.915 41.180 ;
        RECT 31.505 40.480 31.805 42.210 ;
        RECT 42.435 42.190 43.815 42.760 ;
        RECT 49.915 42.610 51.295 43.180 ;
        RECT 61.885 43.160 62.185 44.890 ;
        RECT 69.715 44.180 70.815 44.950 ;
        RECT 73.105 44.880 73.385 46.870 ;
        RECT 75.455 47.710 75.955 68.510 ;
        RECT 76.295 49.030 76.685 70.540 ;
        RECT 77.085 69.950 77.975 70.680 ;
        RECT 77.185 65.130 77.445 69.950 ;
        RECT 78.825 68.560 81.535 69.410 ;
        RECT 79.025 65.780 80.955 68.560 ;
        RECT 86.685 68.520 87.225 71.750 ;
        RECT 87.525 70.550 87.935 73.230 ;
        RECT 95.045 73.060 97.115 74.340 ;
        RECT 98.150 73.310 100.710 75.750 ;
        RECT 109.390 75.480 111.950 75.560 ;
        RECT 121.930 75.480 122.210 85.700 ;
        RECT 127.550 85.510 128.770 89.380 ;
        RECT 127.910 76.040 128.190 85.510 ;
        RECT 133.380 76.580 136.010 77.880 ;
        RECT 137.240 76.560 139.870 77.860 ;
        RECT 109.390 75.200 122.210 75.480 ;
        RECT 97.665 71.740 98.525 72.580 ;
        RECT 83.925 67.070 85.045 67.750 ;
        RECT 84.205 65.790 84.875 67.070 ;
        RECT 77.585 65.400 82.635 65.780 ;
        RECT 83.995 65.380 85.045 65.790 ;
        RECT 77.185 63.580 77.565 65.130 ;
        RECT 77.305 55.740 77.565 63.580 ;
        RECT 82.615 63.140 82.885 65.180 ;
        RECT 83.745 63.140 84.015 65.140 ;
        RECT 82.615 56.450 84.015 63.140 ;
        RECT 77.215 55.230 77.575 55.740 ;
        RECT 77.195 54.800 77.575 55.230 ;
        RECT 82.615 55.130 82.885 56.450 ;
        RECT 83.745 55.090 84.015 56.450 ;
        RECT 85.015 55.200 85.335 65.130 ;
        RECT 85.015 55.140 85.345 55.200 ;
        RECT 77.195 54.520 77.445 54.800 ;
        RECT 76.995 54.120 81.635 54.520 ;
        RECT 82.535 54.230 83.665 54.240 ;
        RECT 85.025 54.230 85.345 55.140 ;
        RECT 77.195 52.000 77.445 54.120 ;
        RECT 81.895 53.430 82.255 54.050 ;
        RECT 81.975 52.550 82.235 53.430 ;
        RECT 82.515 53.180 85.345 54.230 ;
        RECT 81.805 52.170 82.335 52.550 ;
        RECT 77.195 51.910 77.695 52.000 ;
        RECT 77.185 51.180 77.695 51.910 ;
        RECT 77.425 50.180 77.695 51.180 ;
        RECT 78.335 50.930 78.605 51.880 ;
        RECT 78.335 50.780 78.805 50.930 ;
        RECT 78.335 50.100 78.895 50.780 ;
        RECT 78.415 50.090 78.895 50.100 ;
        RECT 77.705 49.560 78.325 49.920 ;
        RECT 77.745 49.030 78.175 49.560 ;
        RECT 76.295 48.610 78.175 49.030 ;
        RECT 78.665 48.900 78.895 50.090 ;
        RECT 77.745 47.740 78.175 48.610 ;
        RECT 78.585 48.300 78.965 48.900 ;
        RECT 75.455 47.000 76.145 47.710 ;
        RECT 77.565 47.380 78.185 47.740 ;
        RECT 77.265 47.000 77.555 47.190 ;
        RECT 75.455 46.560 77.555 47.000 ;
        RECT 75.455 46.540 76.145 46.560 ;
        RECT 77.265 46.320 77.555 46.560 ;
        RECT 78.185 46.930 78.455 47.180 ;
        RECT 78.665 46.930 78.895 48.300 ;
        RECT 81.485 46.950 81.815 51.970 ;
        RECT 82.535 51.960 83.665 53.180 ;
        RECT 85.025 53.160 85.345 53.180 ;
        RECT 78.185 46.820 78.895 46.930 ;
        RECT 81.475 46.900 81.815 46.950 ;
        RECT 82.365 47.720 83.745 51.960 ;
        RECT 78.185 46.510 78.845 46.820 ;
        RECT 78.185 46.340 78.455 46.510 ;
        RECT 81.475 44.940 81.755 46.900 ;
        RECT 82.365 46.860 82.665 47.720 ;
        RECT 83.445 46.860 83.745 47.720 ;
        RECT 84.295 46.860 84.625 51.930 ;
        RECT 83.695 46.320 84.175 46.700 ;
        RECT 83.795 45.700 84.045 46.320 ;
        RECT 83.695 45.100 84.075 45.700 ;
        RECT 53.655 42.190 55.035 42.760 ;
        RECT 61.165 42.590 62.545 43.160 ;
        RECT 73.105 43.150 73.405 44.880 ;
        RECT 80.955 44.170 82.055 44.940 ;
        RECT 84.345 44.870 84.625 46.860 ;
        RECT 86.705 47.720 87.205 68.520 ;
        RECT 87.545 49.040 87.935 70.550 ;
        RECT 88.335 69.960 89.225 70.690 ;
        RECT 88.435 65.140 88.695 69.960 ;
        RECT 90.075 68.570 92.785 69.420 ;
        RECT 90.275 65.790 92.205 68.570 ;
        RECT 97.965 68.510 98.505 71.740 ;
        RECT 98.805 70.540 99.215 73.310 ;
        RECT 106.455 73.110 108.525 74.390 ;
        RECT 109.390 73.030 111.950 75.200 ;
        RECT 125.760 74.810 128.190 76.040 ;
        RECT 121.290 74.790 128.190 74.810 ;
        RECT 120.600 74.530 128.190 74.790 ;
        RECT 117.655 73.110 119.725 74.390 ;
        RECT 120.600 73.180 128.160 74.530 ;
        RECT 129.505 73.190 131.575 74.470 ;
        RECT 120.600 73.110 126.160 73.180 ;
        RECT 108.935 71.740 109.795 72.580 ;
        RECT 95.175 67.080 96.295 67.760 ;
        RECT 95.455 65.800 96.125 67.080 ;
        RECT 88.835 65.410 93.885 65.790 ;
        RECT 95.245 65.390 96.295 65.800 ;
        RECT 88.435 63.590 88.815 65.140 ;
        RECT 88.555 55.750 88.815 63.590 ;
        RECT 93.865 63.150 94.135 65.190 ;
        RECT 94.995 63.150 95.265 65.150 ;
        RECT 93.865 56.460 95.265 63.150 ;
        RECT 88.465 55.240 88.825 55.750 ;
        RECT 88.445 54.810 88.825 55.240 ;
        RECT 93.865 55.140 94.135 56.460 ;
        RECT 94.995 55.100 95.265 56.460 ;
        RECT 96.265 55.210 96.585 65.140 ;
        RECT 96.265 55.150 96.595 55.210 ;
        RECT 88.445 54.530 88.695 54.810 ;
        RECT 88.245 54.130 92.885 54.530 ;
        RECT 93.785 54.240 94.915 54.250 ;
        RECT 96.275 54.240 96.595 55.150 ;
        RECT 88.445 52.010 88.695 54.130 ;
        RECT 93.145 53.440 93.505 54.060 ;
        RECT 93.225 52.560 93.485 53.440 ;
        RECT 93.765 53.190 96.595 54.240 ;
        RECT 93.055 52.180 93.585 52.560 ;
        RECT 88.445 51.920 88.945 52.010 ;
        RECT 88.435 51.190 88.945 51.920 ;
        RECT 88.675 50.190 88.945 51.190 ;
        RECT 89.585 50.940 89.855 51.890 ;
        RECT 89.585 50.790 90.055 50.940 ;
        RECT 89.585 50.110 90.145 50.790 ;
        RECT 89.665 50.100 90.145 50.110 ;
        RECT 88.955 49.570 89.575 49.930 ;
        RECT 88.995 49.040 89.425 49.570 ;
        RECT 87.545 48.620 89.425 49.040 ;
        RECT 89.915 48.910 90.145 50.100 ;
        RECT 88.995 47.750 89.425 48.620 ;
        RECT 89.835 48.310 90.215 48.910 ;
        RECT 86.705 47.010 87.395 47.720 ;
        RECT 88.815 47.390 89.435 47.750 ;
        RECT 88.515 47.010 88.805 47.200 ;
        RECT 86.705 46.570 88.805 47.010 ;
        RECT 86.705 46.550 87.395 46.570 ;
        RECT 88.515 46.330 88.805 46.570 ;
        RECT 89.435 46.940 89.705 47.190 ;
        RECT 89.915 46.940 90.145 48.310 ;
        RECT 92.735 46.960 93.065 51.980 ;
        RECT 93.785 51.970 94.915 53.190 ;
        RECT 96.275 53.170 96.595 53.190 ;
        RECT 89.435 46.830 90.145 46.940 ;
        RECT 92.725 46.910 93.065 46.960 ;
        RECT 93.615 47.730 94.995 51.970 ;
        RECT 89.435 46.520 90.095 46.830 ;
        RECT 89.435 46.350 89.705 46.520 ;
        RECT 92.725 44.950 93.005 46.910 ;
        RECT 93.615 46.870 93.915 47.730 ;
        RECT 94.695 46.870 94.995 47.730 ;
        RECT 95.545 46.870 95.875 51.940 ;
        RECT 94.945 46.330 95.425 46.710 ;
        RECT 95.045 45.710 95.295 46.330 ;
        RECT 94.945 45.110 95.325 45.710 ;
        RECT 64.855 42.190 66.235 42.760 ;
        RECT 72.385 42.580 73.765 43.150 ;
        RECT 84.345 43.140 84.645 44.870 ;
        RECT 92.205 44.180 93.305 44.950 ;
        RECT 95.595 44.880 95.875 46.870 ;
        RECT 97.985 47.710 98.485 68.510 ;
        RECT 98.825 49.030 99.215 70.540 ;
        RECT 99.615 69.950 100.505 70.680 ;
        RECT 99.715 65.130 99.975 69.950 ;
        RECT 101.355 68.560 104.065 69.410 ;
        RECT 101.555 65.780 103.485 68.560 ;
        RECT 109.235 68.510 109.775 71.740 ;
        RECT 110.075 70.540 110.485 73.030 ;
        RECT 120.185 71.740 121.045 72.580 ;
        RECT 106.455 67.070 107.575 67.750 ;
        RECT 106.735 65.790 107.405 67.070 ;
        RECT 100.115 65.400 105.165 65.780 ;
        RECT 106.525 65.380 107.575 65.790 ;
        RECT 99.715 63.580 100.095 65.130 ;
        RECT 99.835 55.740 100.095 63.580 ;
        RECT 105.145 63.140 105.415 65.180 ;
        RECT 106.275 63.140 106.545 65.140 ;
        RECT 105.145 56.450 106.545 63.140 ;
        RECT 99.745 55.230 100.105 55.740 ;
        RECT 99.725 54.800 100.105 55.230 ;
        RECT 105.145 55.130 105.415 56.450 ;
        RECT 106.275 55.090 106.545 56.450 ;
        RECT 107.545 55.200 107.865 65.130 ;
        RECT 107.545 55.140 107.875 55.200 ;
        RECT 99.725 54.520 99.975 54.800 ;
        RECT 99.525 54.120 104.165 54.520 ;
        RECT 105.065 54.230 106.195 54.240 ;
        RECT 107.555 54.230 107.875 55.140 ;
        RECT 99.725 52.000 99.975 54.120 ;
        RECT 104.425 53.430 104.785 54.050 ;
        RECT 104.505 52.550 104.765 53.430 ;
        RECT 105.045 53.180 107.875 54.230 ;
        RECT 104.335 52.170 104.865 52.550 ;
        RECT 99.725 51.910 100.225 52.000 ;
        RECT 99.715 51.180 100.225 51.910 ;
        RECT 99.955 50.180 100.225 51.180 ;
        RECT 100.865 50.930 101.135 51.880 ;
        RECT 100.865 50.780 101.335 50.930 ;
        RECT 100.865 50.100 101.425 50.780 ;
        RECT 100.945 50.090 101.425 50.100 ;
        RECT 100.235 49.560 100.855 49.920 ;
        RECT 100.275 49.030 100.705 49.560 ;
        RECT 98.825 48.610 100.705 49.030 ;
        RECT 101.195 48.900 101.425 50.090 ;
        RECT 100.275 47.740 100.705 48.610 ;
        RECT 101.115 48.300 101.495 48.900 ;
        RECT 97.985 47.000 98.675 47.710 ;
        RECT 100.095 47.380 100.715 47.740 ;
        RECT 99.795 47.000 100.085 47.190 ;
        RECT 97.985 46.560 100.085 47.000 ;
        RECT 97.985 46.540 98.675 46.560 ;
        RECT 99.795 46.320 100.085 46.560 ;
        RECT 100.715 46.930 100.985 47.180 ;
        RECT 101.195 46.930 101.425 48.300 ;
        RECT 104.015 46.950 104.345 51.970 ;
        RECT 105.065 51.960 106.195 53.180 ;
        RECT 107.555 53.160 107.875 53.180 ;
        RECT 100.715 46.820 101.425 46.930 ;
        RECT 104.005 46.900 104.345 46.950 ;
        RECT 104.895 47.720 106.275 51.960 ;
        RECT 100.715 46.510 101.375 46.820 ;
        RECT 100.715 46.340 100.985 46.510 ;
        RECT 104.005 44.940 104.285 46.900 ;
        RECT 104.895 46.860 105.195 47.720 ;
        RECT 105.975 46.860 106.275 47.720 ;
        RECT 106.825 46.860 107.155 51.930 ;
        RECT 106.225 46.320 106.705 46.700 ;
        RECT 106.325 45.700 106.575 46.320 ;
        RECT 106.225 45.100 106.605 45.700 ;
        RECT 95.595 43.150 95.895 44.880 ;
        RECT 103.485 44.170 104.585 44.940 ;
        RECT 106.875 44.870 107.155 46.860 ;
        RECT 109.255 47.710 109.755 68.510 ;
        RECT 110.095 49.030 110.485 70.540 ;
        RECT 110.885 69.950 111.775 70.680 ;
        RECT 110.985 65.130 111.245 69.950 ;
        RECT 112.625 68.560 115.335 69.410 ;
        RECT 112.825 65.780 114.755 68.560 ;
        RECT 120.485 68.510 121.025 71.740 ;
        RECT 121.325 70.540 121.735 73.110 ;
        RECT 132.925 70.810 133.225 70.900 ;
        RECT 117.725 67.070 118.845 67.750 ;
        RECT 118.005 65.790 118.675 67.070 ;
        RECT 111.385 65.400 116.435 65.780 ;
        RECT 117.795 65.380 118.845 65.790 ;
        RECT 110.985 63.580 111.365 65.130 ;
        RECT 111.105 55.740 111.365 63.580 ;
        RECT 116.415 63.140 116.685 65.180 ;
        RECT 117.545 63.140 117.815 65.140 ;
        RECT 116.415 56.450 117.815 63.140 ;
        RECT 111.015 55.230 111.375 55.740 ;
        RECT 110.995 54.800 111.375 55.230 ;
        RECT 116.415 55.130 116.685 56.450 ;
        RECT 117.545 55.090 117.815 56.450 ;
        RECT 118.815 55.200 119.135 65.130 ;
        RECT 118.815 55.140 119.145 55.200 ;
        RECT 110.995 54.520 111.245 54.800 ;
        RECT 110.795 54.120 115.435 54.520 ;
        RECT 116.335 54.230 117.465 54.240 ;
        RECT 118.825 54.230 119.145 55.140 ;
        RECT 110.995 52.000 111.245 54.120 ;
        RECT 115.695 53.430 116.055 54.050 ;
        RECT 115.775 52.550 116.035 53.430 ;
        RECT 116.315 53.180 119.145 54.230 ;
        RECT 115.605 52.170 116.135 52.550 ;
        RECT 110.995 51.910 111.495 52.000 ;
        RECT 110.985 51.180 111.495 51.910 ;
        RECT 111.225 50.180 111.495 51.180 ;
        RECT 112.135 50.930 112.405 51.880 ;
        RECT 112.135 50.780 112.605 50.930 ;
        RECT 112.135 50.100 112.695 50.780 ;
        RECT 112.215 50.090 112.695 50.100 ;
        RECT 111.505 49.560 112.125 49.920 ;
        RECT 111.545 49.030 111.975 49.560 ;
        RECT 110.095 48.610 111.975 49.030 ;
        RECT 112.465 48.900 112.695 50.090 ;
        RECT 111.545 47.740 111.975 48.610 ;
        RECT 112.385 48.300 112.765 48.900 ;
        RECT 109.255 47.000 109.945 47.710 ;
        RECT 111.365 47.380 111.985 47.740 ;
        RECT 111.065 47.000 111.355 47.190 ;
        RECT 109.255 46.560 111.355 47.000 ;
        RECT 109.255 46.540 109.945 46.560 ;
        RECT 111.065 46.320 111.355 46.560 ;
        RECT 111.985 46.930 112.255 47.180 ;
        RECT 112.465 46.930 112.695 48.300 ;
        RECT 115.285 46.950 115.615 51.970 ;
        RECT 116.335 51.960 117.465 53.180 ;
        RECT 118.825 53.160 119.145 53.180 ;
        RECT 111.985 46.820 112.695 46.930 ;
        RECT 115.275 46.900 115.615 46.950 ;
        RECT 116.165 47.720 117.545 51.960 ;
        RECT 111.985 46.510 112.645 46.820 ;
        RECT 111.985 46.340 112.255 46.510 ;
        RECT 115.275 44.940 115.555 46.900 ;
        RECT 116.165 46.860 116.465 47.720 ;
        RECT 117.245 46.860 117.545 47.720 ;
        RECT 118.095 46.860 118.425 51.930 ;
        RECT 117.495 46.320 117.975 46.700 ;
        RECT 117.595 45.700 117.845 46.320 ;
        RECT 117.495 45.100 117.875 45.700 ;
        RECT 20.795 39.650 21.175 40.250 ;
        RECT 20.825 39.030 21.075 39.650 ;
        RECT 20.695 38.650 21.175 39.030 ;
        RECT 20.245 33.420 20.575 38.490 ;
        RECT 21.125 37.630 21.425 38.490 ;
        RECT 22.205 37.630 22.505 38.490 ;
        RECT 23.115 38.450 23.395 40.410 ;
        RECT 26.415 38.840 26.685 39.010 ;
        RECT 26.025 38.530 26.685 38.840 ;
        RECT 21.125 33.390 22.505 37.630 ;
        RECT 23.055 38.400 23.395 38.450 ;
        RECT 25.975 38.420 26.685 38.530 ;
        RECT 19.525 32.170 19.845 32.190 ;
        RECT 21.205 32.170 22.335 33.390 ;
        RECT 23.055 33.380 23.385 38.400 ;
        RECT 25.975 37.050 26.205 38.420 ;
        RECT 26.415 38.170 26.685 38.420 ;
        RECT 27.315 38.790 27.605 39.030 ;
        RECT 28.725 38.790 29.415 38.810 ;
        RECT 27.315 38.350 29.415 38.790 ;
        RECT 27.315 38.160 27.605 38.350 ;
        RECT 26.685 37.610 27.305 37.970 ;
        RECT 28.725 37.640 29.415 38.350 ;
        RECT 25.905 36.450 26.285 37.050 ;
        RECT 26.695 36.740 27.125 37.610 ;
        RECT 25.975 35.260 26.205 36.450 ;
        RECT 26.695 36.320 28.575 36.740 ;
        RECT 26.695 35.790 27.125 36.320 ;
        RECT 26.545 35.430 27.165 35.790 ;
        RECT 25.975 35.250 26.455 35.260 ;
        RECT 25.975 34.570 26.535 35.250 ;
        RECT 26.065 34.420 26.535 34.570 ;
        RECT 26.265 33.470 26.535 34.420 ;
        RECT 27.175 34.170 27.445 35.170 ;
        RECT 27.175 33.440 27.685 34.170 ;
        RECT 27.175 33.350 27.675 33.440 ;
        RECT 22.535 32.800 23.065 33.180 ;
        RECT 19.525 31.120 22.355 32.170 ;
        RECT 22.635 31.920 22.895 32.800 ;
        RECT 22.615 31.300 22.975 31.920 ;
        RECT 27.425 31.230 27.675 33.350 ;
        RECT 19.525 30.210 19.845 31.120 ;
        RECT 21.205 31.110 22.335 31.120 ;
        RECT 23.235 30.830 27.875 31.230 ;
        RECT 27.425 30.550 27.675 30.830 ;
        RECT 19.525 30.150 19.855 30.210 ;
        RECT 19.535 20.220 19.855 30.150 ;
        RECT 20.855 28.900 21.125 30.260 ;
        RECT 21.985 28.900 22.255 30.220 ;
        RECT 27.295 30.120 27.675 30.550 ;
        RECT 27.295 29.610 27.655 30.120 ;
        RECT 20.855 22.210 22.255 28.900 ;
        RECT 20.855 20.210 21.125 22.210 ;
        RECT 21.985 20.170 22.255 22.210 ;
        RECT 27.305 21.770 27.565 29.610 ;
        RECT 27.305 20.220 27.685 21.770 ;
        RECT 19.825 19.560 20.875 19.970 ;
        RECT 22.235 19.570 27.285 19.950 ;
        RECT 19.995 18.280 20.665 19.560 ;
        RECT 19.825 17.600 20.945 18.280 ;
        RECT 23.915 16.790 25.845 19.570 ;
        RECT 23.335 15.940 26.045 16.790 ;
        RECT 27.425 15.400 27.685 20.220 ;
        RECT 26.895 14.670 27.785 15.400 ;
        RECT 28.185 14.810 28.575 36.320 ;
        RECT 28.915 16.840 29.415 37.640 ;
        RECT 31.525 38.490 31.805 40.480 ;
        RECT 34.095 40.410 35.195 41.180 ;
        RECT 42.795 40.460 43.095 42.190 ;
        RECT 32.075 39.650 32.455 40.250 ;
        RECT 32.105 39.030 32.355 39.650 ;
        RECT 31.975 38.650 32.455 39.030 ;
        RECT 31.525 33.420 31.855 38.490 ;
        RECT 32.405 37.630 32.705 38.490 ;
        RECT 33.485 37.630 33.785 38.490 ;
        RECT 34.395 38.450 34.675 40.410 ;
        RECT 37.695 38.840 37.965 39.010 ;
        RECT 37.305 38.530 37.965 38.840 ;
        RECT 32.405 33.390 33.785 37.630 ;
        RECT 34.335 38.400 34.675 38.450 ;
        RECT 37.255 38.420 37.965 38.530 ;
        RECT 30.805 32.170 31.125 32.190 ;
        RECT 32.485 32.170 33.615 33.390 ;
        RECT 34.335 33.380 34.665 38.400 ;
        RECT 37.255 37.050 37.485 38.420 ;
        RECT 37.695 38.170 37.965 38.420 ;
        RECT 38.595 38.790 38.885 39.030 ;
        RECT 40.005 38.790 40.695 38.810 ;
        RECT 38.595 38.350 40.695 38.790 ;
        RECT 38.595 38.160 38.885 38.350 ;
        RECT 37.965 37.610 38.585 37.970 ;
        RECT 40.005 37.640 40.695 38.350 ;
        RECT 37.185 36.450 37.565 37.050 ;
        RECT 37.975 36.740 38.405 37.610 ;
        RECT 37.255 35.260 37.485 36.450 ;
        RECT 37.975 36.320 39.855 36.740 ;
        RECT 37.975 35.790 38.405 36.320 ;
        RECT 37.825 35.430 38.445 35.790 ;
        RECT 37.255 35.250 37.735 35.260 ;
        RECT 37.255 34.570 37.815 35.250 ;
        RECT 37.345 34.420 37.815 34.570 ;
        RECT 37.545 33.470 37.815 34.420 ;
        RECT 38.455 34.170 38.725 35.170 ;
        RECT 38.455 33.440 38.965 34.170 ;
        RECT 38.455 33.350 38.955 33.440 ;
        RECT 33.815 32.800 34.345 33.180 ;
        RECT 30.805 31.120 33.635 32.170 ;
        RECT 33.915 31.920 34.175 32.800 ;
        RECT 33.895 31.300 34.255 31.920 ;
        RECT 38.705 31.230 38.955 33.350 ;
        RECT 30.805 30.210 31.125 31.120 ;
        RECT 32.485 31.110 33.615 31.120 ;
        RECT 34.515 30.830 39.155 31.230 ;
        RECT 38.705 30.550 38.955 30.830 ;
        RECT 30.805 30.150 31.135 30.210 ;
        RECT 30.815 20.220 31.135 30.150 ;
        RECT 32.135 28.900 32.405 30.260 ;
        RECT 33.265 28.900 33.535 30.220 ;
        RECT 38.575 30.120 38.955 30.550 ;
        RECT 38.575 29.610 38.935 30.120 ;
        RECT 32.135 22.210 33.535 28.900 ;
        RECT 32.135 20.210 32.405 22.210 ;
        RECT 33.265 20.170 33.535 22.210 ;
        RECT 38.585 21.770 38.845 29.610 ;
        RECT 38.585 20.220 38.965 21.770 ;
        RECT 31.105 19.560 32.155 19.970 ;
        RECT 33.515 19.570 38.565 19.950 ;
        RECT 31.275 18.280 31.945 19.560 ;
        RECT 31.105 17.600 32.225 18.280 ;
        RECT 28.185 12.290 28.595 14.810 ;
        RECT 28.895 13.610 29.435 16.840 ;
        RECT 35.195 16.790 37.125 19.570 ;
        RECT 34.615 15.940 37.325 16.790 ;
        RECT 38.705 15.400 38.965 20.220 ;
        RECT 38.175 14.670 39.065 15.400 ;
        RECT 39.465 14.810 39.855 36.320 ;
        RECT 40.195 16.840 40.695 37.640 ;
        RECT 42.815 38.470 43.095 40.460 ;
        RECT 45.385 40.390 46.485 41.160 ;
        RECT 54.015 40.460 54.315 42.190 ;
        RECT 43.365 39.630 43.745 40.230 ;
        RECT 43.395 39.010 43.645 39.630 ;
        RECT 43.265 38.630 43.745 39.010 ;
        RECT 42.815 33.400 43.145 38.470 ;
        RECT 43.695 37.610 43.995 38.470 ;
        RECT 44.775 37.610 45.075 38.470 ;
        RECT 45.685 38.430 45.965 40.390 ;
        RECT 48.985 38.820 49.255 38.990 ;
        RECT 48.595 38.510 49.255 38.820 ;
        RECT 43.695 33.370 45.075 37.610 ;
        RECT 45.625 38.380 45.965 38.430 ;
        RECT 48.545 38.400 49.255 38.510 ;
        RECT 42.095 32.150 42.415 32.170 ;
        RECT 43.775 32.150 44.905 33.370 ;
        RECT 45.625 33.360 45.955 38.380 ;
        RECT 48.545 37.030 48.775 38.400 ;
        RECT 48.985 38.150 49.255 38.400 ;
        RECT 49.885 38.770 50.175 39.010 ;
        RECT 51.295 38.770 51.985 38.790 ;
        RECT 49.885 38.330 51.985 38.770 ;
        RECT 49.885 38.140 50.175 38.330 ;
        RECT 49.255 37.590 49.875 37.950 ;
        RECT 51.295 37.620 51.985 38.330 ;
        RECT 48.475 36.430 48.855 37.030 ;
        RECT 49.265 36.720 49.695 37.590 ;
        RECT 48.545 35.240 48.775 36.430 ;
        RECT 49.265 36.300 51.145 36.720 ;
        RECT 49.265 35.770 49.695 36.300 ;
        RECT 49.115 35.410 49.735 35.770 ;
        RECT 48.545 35.230 49.025 35.240 ;
        RECT 48.545 34.550 49.105 35.230 ;
        RECT 48.635 34.400 49.105 34.550 ;
        RECT 48.835 33.450 49.105 34.400 ;
        RECT 49.745 34.150 50.015 35.150 ;
        RECT 49.745 33.420 50.255 34.150 ;
        RECT 49.745 33.330 50.245 33.420 ;
        RECT 45.105 32.780 45.635 33.160 ;
        RECT 42.095 31.100 44.925 32.150 ;
        RECT 45.205 31.900 45.465 32.780 ;
        RECT 45.185 31.280 45.545 31.900 ;
        RECT 49.995 31.210 50.245 33.330 ;
        RECT 42.095 30.190 42.415 31.100 ;
        RECT 43.775 31.090 44.905 31.100 ;
        RECT 45.805 30.810 50.445 31.210 ;
        RECT 49.995 30.530 50.245 30.810 ;
        RECT 42.095 30.130 42.425 30.190 ;
        RECT 42.105 20.200 42.425 30.130 ;
        RECT 43.425 28.880 43.695 30.240 ;
        RECT 44.555 28.880 44.825 30.200 ;
        RECT 49.865 30.100 50.245 30.530 ;
        RECT 49.865 29.590 50.225 30.100 ;
        RECT 43.425 22.190 44.825 28.880 ;
        RECT 43.425 20.190 43.695 22.190 ;
        RECT 44.555 20.150 44.825 22.190 ;
        RECT 49.875 21.750 50.135 29.590 ;
        RECT 49.875 20.200 50.255 21.750 ;
        RECT 42.395 19.540 43.445 19.950 ;
        RECT 44.805 19.550 49.855 19.930 ;
        RECT 42.565 18.260 43.235 19.540 ;
        RECT 42.395 17.580 43.515 18.260 ;
        RECT 28.875 12.770 29.735 13.610 ;
        RECT 28.185 11.950 30.415 12.290 ;
        RECT 39.465 11.990 39.875 14.810 ;
        RECT 40.175 13.610 40.715 16.840 ;
        RECT 46.485 16.770 48.415 19.550 ;
        RECT 45.905 15.920 48.615 16.770 ;
        RECT 49.995 15.380 50.255 20.200 ;
        RECT 49.465 14.650 50.355 15.380 ;
        RECT 50.755 14.790 51.145 36.300 ;
        RECT 51.485 16.820 51.985 37.620 ;
        RECT 54.035 38.470 54.315 40.460 ;
        RECT 56.605 40.390 57.705 41.160 ;
        RECT 65.215 40.460 65.515 42.190 ;
        RECT 76.145 42.180 77.525 42.750 ;
        RECT 83.625 42.570 85.005 43.140 ;
        RECT 87.385 42.200 88.765 42.770 ;
        RECT 94.875 42.580 96.255 43.150 ;
        RECT 106.875 43.140 107.175 44.870 ;
        RECT 114.755 44.170 115.855 44.940 ;
        RECT 118.145 44.870 118.425 46.860 ;
        RECT 120.505 47.710 121.005 68.510 ;
        RECT 121.345 49.030 121.735 70.540 ;
        RECT 122.135 69.950 123.025 70.680 ;
        RECT 132.615 70.040 134.265 70.810 ;
        RECT 122.235 65.130 122.495 69.950 ;
        RECT 123.875 68.560 126.585 69.410 ;
        RECT 124.075 65.780 126.005 68.560 ;
        RECT 128.975 67.070 130.095 67.750 ;
        RECT 129.255 65.790 129.925 67.070 ;
        RECT 122.635 65.400 127.685 65.780 ;
        RECT 129.045 65.380 130.095 65.790 ;
        RECT 132.925 65.180 133.225 70.040 ;
        RECT 137.675 68.690 139.075 69.460 ;
        RECT 138.385 65.740 138.645 68.690 ;
        RECT 149.410 68.420 150.690 69.620 ;
        RECT 149.480 65.810 150.640 68.420 ;
        RECT 133.365 65.380 138.645 65.740 ;
        RECT 122.235 63.580 122.615 65.130 ;
        RECT 122.355 55.740 122.615 63.580 ;
        RECT 127.665 63.140 127.935 65.180 ;
        RECT 128.795 63.140 129.065 65.140 ;
        RECT 127.665 56.450 129.065 63.140 ;
        RECT 122.265 55.230 122.625 55.740 ;
        RECT 122.245 54.800 122.625 55.230 ;
        RECT 127.665 55.130 127.935 56.450 ;
        RECT 128.795 55.090 129.065 56.450 ;
        RECT 130.065 55.200 130.385 65.130 ;
        RECT 132.925 61.010 133.355 65.180 ;
        RECT 138.385 65.150 138.645 65.380 ;
        RECT 138.385 64.770 138.675 65.150 ;
        RECT 130.065 55.140 130.395 55.200 ;
        RECT 133.055 55.190 133.355 61.010 ;
        RECT 122.245 54.520 122.495 54.800 ;
        RECT 122.045 54.120 126.685 54.520 ;
        RECT 127.585 54.230 128.715 54.240 ;
        RECT 130.075 54.230 130.395 55.140 ;
        RECT 138.395 55.080 138.675 64.770 ;
        RECT 149.390 64.610 150.670 65.810 ;
        RECT 122.245 52.000 122.495 54.120 ;
        RECT 126.945 53.430 127.305 54.050 ;
        RECT 127.025 52.550 127.285 53.430 ;
        RECT 127.565 53.180 130.395 54.230 ;
        RECT 126.855 52.170 127.385 52.550 ;
        RECT 122.245 51.910 122.745 52.000 ;
        RECT 122.235 51.180 122.745 51.910 ;
        RECT 122.475 50.180 122.745 51.180 ;
        RECT 123.385 50.930 123.655 51.880 ;
        RECT 123.385 50.780 123.855 50.930 ;
        RECT 123.385 50.100 123.945 50.780 ;
        RECT 123.465 50.090 123.945 50.100 ;
        RECT 122.755 49.560 123.375 49.920 ;
        RECT 122.795 49.030 123.225 49.560 ;
        RECT 121.345 48.610 123.225 49.030 ;
        RECT 123.715 48.900 123.945 50.090 ;
        RECT 122.795 47.740 123.225 48.610 ;
        RECT 123.635 48.300 124.015 48.900 ;
        RECT 120.505 47.000 121.195 47.710 ;
        RECT 122.615 47.380 123.235 47.740 ;
        RECT 122.315 47.000 122.605 47.190 ;
        RECT 120.505 46.560 122.605 47.000 ;
        RECT 120.505 46.540 121.195 46.560 ;
        RECT 122.315 46.320 122.605 46.560 ;
        RECT 123.235 46.930 123.505 47.180 ;
        RECT 123.715 46.930 123.945 48.300 ;
        RECT 126.535 46.950 126.865 51.970 ;
        RECT 127.585 51.960 128.715 53.180 ;
        RECT 130.075 53.160 130.395 53.180 ;
        RECT 123.235 46.820 123.945 46.930 ;
        RECT 126.525 46.900 126.865 46.950 ;
        RECT 127.415 47.720 128.795 51.960 ;
        RECT 123.235 46.510 123.895 46.820 ;
        RECT 123.235 46.340 123.505 46.510 ;
        RECT 126.525 44.940 126.805 46.900 ;
        RECT 127.415 46.860 127.715 47.720 ;
        RECT 128.495 46.860 128.795 47.720 ;
        RECT 129.345 46.860 129.675 51.930 ;
        RECT 128.745 46.320 129.225 46.700 ;
        RECT 128.845 45.700 129.095 46.320 ;
        RECT 128.745 45.100 129.125 45.700 ;
        RECT 118.145 43.140 118.445 44.870 ;
        RECT 126.005 44.170 127.105 44.940 ;
        RECT 129.395 44.870 129.675 46.860 ;
        RECT 129.395 43.140 129.695 44.870 ;
        RECT 98.595 42.220 99.975 42.790 ;
        RECT 106.155 42.570 107.535 43.140 ;
        RECT 109.795 42.260 111.175 42.830 ;
        RECT 117.425 42.570 118.805 43.140 ;
        RECT 121.005 42.280 122.385 42.850 ;
        RECT 128.675 42.570 130.055 43.140 ;
        RECT 54.585 39.630 54.965 40.230 ;
        RECT 54.615 39.010 54.865 39.630 ;
        RECT 54.485 38.630 54.965 39.010 ;
        RECT 54.035 33.400 54.365 38.470 ;
        RECT 54.915 37.610 55.215 38.470 ;
        RECT 55.995 37.610 56.295 38.470 ;
        RECT 56.905 38.430 57.185 40.390 ;
        RECT 60.205 38.820 60.475 38.990 ;
        RECT 59.815 38.510 60.475 38.820 ;
        RECT 54.915 33.370 56.295 37.610 ;
        RECT 56.845 38.380 57.185 38.430 ;
        RECT 59.765 38.400 60.475 38.510 ;
        RECT 53.315 32.150 53.635 32.170 ;
        RECT 54.995 32.150 56.125 33.370 ;
        RECT 56.845 33.360 57.175 38.380 ;
        RECT 59.765 37.030 59.995 38.400 ;
        RECT 60.205 38.150 60.475 38.400 ;
        RECT 61.105 38.770 61.395 39.010 ;
        RECT 62.515 38.770 63.205 38.790 ;
        RECT 61.105 38.330 63.205 38.770 ;
        RECT 61.105 38.140 61.395 38.330 ;
        RECT 60.475 37.590 61.095 37.950 ;
        RECT 62.515 37.620 63.205 38.330 ;
        RECT 59.695 36.430 60.075 37.030 ;
        RECT 60.485 36.720 60.915 37.590 ;
        RECT 59.765 35.240 59.995 36.430 ;
        RECT 60.485 36.300 62.365 36.720 ;
        RECT 60.485 35.770 60.915 36.300 ;
        RECT 60.335 35.410 60.955 35.770 ;
        RECT 59.765 35.230 60.245 35.240 ;
        RECT 59.765 34.550 60.325 35.230 ;
        RECT 59.855 34.400 60.325 34.550 ;
        RECT 60.055 33.450 60.325 34.400 ;
        RECT 60.965 34.150 61.235 35.150 ;
        RECT 60.965 33.420 61.475 34.150 ;
        RECT 60.965 33.330 61.465 33.420 ;
        RECT 56.325 32.780 56.855 33.160 ;
        RECT 53.315 31.100 56.145 32.150 ;
        RECT 56.425 31.900 56.685 32.780 ;
        RECT 56.405 31.280 56.765 31.900 ;
        RECT 61.215 31.210 61.465 33.330 ;
        RECT 53.315 30.190 53.635 31.100 ;
        RECT 54.995 31.090 56.125 31.100 ;
        RECT 57.025 30.810 61.665 31.210 ;
        RECT 61.215 30.530 61.465 30.810 ;
        RECT 53.315 30.130 53.645 30.190 ;
        RECT 53.325 20.200 53.645 30.130 ;
        RECT 54.645 28.880 54.915 30.240 ;
        RECT 55.775 28.880 56.045 30.200 ;
        RECT 61.085 30.100 61.465 30.530 ;
        RECT 61.085 29.590 61.445 30.100 ;
        RECT 54.645 22.190 56.045 28.880 ;
        RECT 54.645 20.190 54.915 22.190 ;
        RECT 55.775 20.150 56.045 22.190 ;
        RECT 61.095 21.750 61.355 29.590 ;
        RECT 61.095 20.200 61.475 21.750 ;
        RECT 53.615 19.540 54.665 19.950 ;
        RECT 56.025 19.550 61.075 19.930 ;
        RECT 53.785 18.260 54.455 19.540 ;
        RECT 53.615 17.580 54.735 18.260 ;
        RECT 40.155 12.770 41.015 13.610 ;
        RECT 50.755 12.170 51.165 14.790 ;
        RECT 51.465 13.590 52.005 16.820 ;
        RECT 57.705 16.770 59.635 19.550 ;
        RECT 57.125 15.920 59.835 16.770 ;
        RECT 61.215 15.380 61.475 20.200 ;
        RECT 60.685 14.650 61.575 15.380 ;
        RECT 61.975 14.790 62.365 36.300 ;
        RECT 62.705 16.820 63.205 37.620 ;
        RECT 65.235 38.470 65.515 40.460 ;
        RECT 67.805 40.390 68.905 41.160 ;
        RECT 76.505 40.450 76.805 42.180 ;
        RECT 65.785 39.630 66.165 40.230 ;
        RECT 65.815 39.010 66.065 39.630 ;
        RECT 65.685 38.630 66.165 39.010 ;
        RECT 65.235 33.400 65.565 38.470 ;
        RECT 66.115 37.610 66.415 38.470 ;
        RECT 67.195 37.610 67.495 38.470 ;
        RECT 68.105 38.430 68.385 40.390 ;
        RECT 71.405 38.820 71.675 38.990 ;
        RECT 71.015 38.510 71.675 38.820 ;
        RECT 66.115 33.370 67.495 37.610 ;
        RECT 68.045 38.380 68.385 38.430 ;
        RECT 70.965 38.400 71.675 38.510 ;
        RECT 64.515 32.150 64.835 32.170 ;
        RECT 66.195 32.150 67.325 33.370 ;
        RECT 68.045 33.360 68.375 38.380 ;
        RECT 70.965 37.030 71.195 38.400 ;
        RECT 71.405 38.150 71.675 38.400 ;
        RECT 72.305 38.770 72.595 39.010 ;
        RECT 73.715 38.770 74.405 38.790 ;
        RECT 72.305 38.330 74.405 38.770 ;
        RECT 72.305 38.140 72.595 38.330 ;
        RECT 71.675 37.590 72.295 37.950 ;
        RECT 73.715 37.620 74.405 38.330 ;
        RECT 70.895 36.430 71.275 37.030 ;
        RECT 71.685 36.720 72.115 37.590 ;
        RECT 70.965 35.240 71.195 36.430 ;
        RECT 71.685 36.300 73.565 36.720 ;
        RECT 71.685 35.770 72.115 36.300 ;
        RECT 71.535 35.410 72.155 35.770 ;
        RECT 70.965 35.230 71.445 35.240 ;
        RECT 70.965 34.550 71.525 35.230 ;
        RECT 71.055 34.400 71.525 34.550 ;
        RECT 71.255 33.450 71.525 34.400 ;
        RECT 72.165 34.150 72.435 35.150 ;
        RECT 72.165 33.420 72.675 34.150 ;
        RECT 72.165 33.330 72.665 33.420 ;
        RECT 67.525 32.780 68.055 33.160 ;
        RECT 64.515 31.100 67.345 32.150 ;
        RECT 67.625 31.900 67.885 32.780 ;
        RECT 67.605 31.280 67.965 31.900 ;
        RECT 72.415 31.210 72.665 33.330 ;
        RECT 64.515 30.190 64.835 31.100 ;
        RECT 66.195 31.090 67.325 31.100 ;
        RECT 68.225 30.810 72.865 31.210 ;
        RECT 72.415 30.530 72.665 30.810 ;
        RECT 64.515 30.130 64.845 30.190 ;
        RECT 64.525 20.200 64.845 30.130 ;
        RECT 65.845 28.880 66.115 30.240 ;
        RECT 66.975 28.880 67.245 30.200 ;
        RECT 72.285 30.100 72.665 30.530 ;
        RECT 72.285 29.590 72.645 30.100 ;
        RECT 65.845 22.190 67.245 28.880 ;
        RECT 65.845 20.190 66.115 22.190 ;
        RECT 66.975 20.150 67.245 22.190 ;
        RECT 72.295 21.750 72.555 29.590 ;
        RECT 72.295 20.200 72.675 21.750 ;
        RECT 64.815 19.540 65.865 19.950 ;
        RECT 67.225 19.550 72.275 19.930 ;
        RECT 64.985 18.260 65.655 19.540 ;
        RECT 64.815 17.580 65.935 18.260 ;
        RECT 51.445 12.750 52.305 13.590 ;
        RECT 27.865 11.130 30.415 11.950 ;
        RECT 28.395 11.090 30.415 11.130 ;
        RECT 39.115 10.980 41.565 11.990 ;
        RECT 50.335 10.970 52.355 12.170 ;
        RECT 61.975 12.160 62.385 14.790 ;
        RECT 62.685 13.590 63.225 16.820 ;
        RECT 68.905 16.770 70.835 19.550 ;
        RECT 68.325 15.920 71.035 16.770 ;
        RECT 72.415 15.380 72.675 20.200 ;
        RECT 71.885 14.650 72.775 15.380 ;
        RECT 73.175 14.790 73.565 36.300 ;
        RECT 73.905 16.820 74.405 37.620 ;
        RECT 76.525 38.460 76.805 40.450 ;
        RECT 79.095 40.380 80.195 41.150 ;
        RECT 87.745 40.470 88.045 42.200 ;
        RECT 77.075 39.620 77.455 40.220 ;
        RECT 77.105 39.000 77.355 39.620 ;
        RECT 76.975 38.620 77.455 39.000 ;
        RECT 76.525 33.390 76.855 38.460 ;
        RECT 77.405 37.600 77.705 38.460 ;
        RECT 78.485 37.600 78.785 38.460 ;
        RECT 79.395 38.420 79.675 40.380 ;
        RECT 82.695 38.810 82.965 38.980 ;
        RECT 82.305 38.500 82.965 38.810 ;
        RECT 77.405 33.360 78.785 37.600 ;
        RECT 79.335 38.370 79.675 38.420 ;
        RECT 82.255 38.390 82.965 38.500 ;
        RECT 75.805 32.140 76.125 32.160 ;
        RECT 77.485 32.140 78.615 33.360 ;
        RECT 79.335 33.350 79.665 38.370 ;
        RECT 82.255 37.020 82.485 38.390 ;
        RECT 82.695 38.140 82.965 38.390 ;
        RECT 83.595 38.760 83.885 39.000 ;
        RECT 85.005 38.760 85.695 38.780 ;
        RECT 83.595 38.320 85.695 38.760 ;
        RECT 83.595 38.130 83.885 38.320 ;
        RECT 82.965 37.580 83.585 37.940 ;
        RECT 85.005 37.610 85.695 38.320 ;
        RECT 82.185 36.420 82.565 37.020 ;
        RECT 82.975 36.710 83.405 37.580 ;
        RECT 82.255 35.230 82.485 36.420 ;
        RECT 82.975 36.290 84.855 36.710 ;
        RECT 82.975 35.760 83.405 36.290 ;
        RECT 82.825 35.400 83.445 35.760 ;
        RECT 82.255 35.220 82.735 35.230 ;
        RECT 82.255 34.540 82.815 35.220 ;
        RECT 82.345 34.390 82.815 34.540 ;
        RECT 82.545 33.440 82.815 34.390 ;
        RECT 83.455 34.140 83.725 35.140 ;
        RECT 83.455 33.410 83.965 34.140 ;
        RECT 83.455 33.320 83.955 33.410 ;
        RECT 78.815 32.770 79.345 33.150 ;
        RECT 75.805 31.090 78.635 32.140 ;
        RECT 78.915 31.890 79.175 32.770 ;
        RECT 78.895 31.270 79.255 31.890 ;
        RECT 83.705 31.200 83.955 33.320 ;
        RECT 75.805 30.180 76.125 31.090 ;
        RECT 77.485 31.080 78.615 31.090 ;
        RECT 79.515 30.800 84.155 31.200 ;
        RECT 83.705 30.520 83.955 30.800 ;
        RECT 75.805 30.120 76.135 30.180 ;
        RECT 75.815 20.190 76.135 30.120 ;
        RECT 77.135 28.870 77.405 30.230 ;
        RECT 78.265 28.870 78.535 30.190 ;
        RECT 83.575 30.090 83.955 30.520 ;
        RECT 83.575 29.580 83.935 30.090 ;
        RECT 77.135 22.180 78.535 28.870 ;
        RECT 77.135 20.180 77.405 22.180 ;
        RECT 78.265 20.140 78.535 22.180 ;
        RECT 83.585 21.740 83.845 29.580 ;
        RECT 83.585 20.190 83.965 21.740 ;
        RECT 76.105 19.530 77.155 19.940 ;
        RECT 78.515 19.540 83.565 19.920 ;
        RECT 76.275 18.250 76.945 19.530 ;
        RECT 76.105 17.570 77.225 18.250 ;
        RECT 62.665 12.750 63.525 13.590 ;
        RECT 73.175 12.190 73.585 14.790 ;
        RECT 73.885 13.590 74.425 16.820 ;
        RECT 80.195 16.760 82.125 19.540 ;
        RECT 79.615 15.910 82.325 16.760 ;
        RECT 83.705 15.370 83.965 20.190 ;
        RECT 83.175 14.640 84.065 15.370 ;
        RECT 84.465 14.780 84.855 36.290 ;
        RECT 85.195 16.810 85.695 37.610 ;
        RECT 87.765 38.480 88.045 40.470 ;
        RECT 90.335 40.400 91.435 41.170 ;
        RECT 98.955 40.490 99.255 42.220 ;
        RECT 88.315 39.640 88.695 40.240 ;
        RECT 88.345 39.020 88.595 39.640 ;
        RECT 88.215 38.640 88.695 39.020 ;
        RECT 87.765 33.410 88.095 38.480 ;
        RECT 88.645 37.620 88.945 38.480 ;
        RECT 89.725 37.620 90.025 38.480 ;
        RECT 90.635 38.440 90.915 40.400 ;
        RECT 93.935 38.830 94.205 39.000 ;
        RECT 93.545 38.520 94.205 38.830 ;
        RECT 88.645 33.380 90.025 37.620 ;
        RECT 90.575 38.390 90.915 38.440 ;
        RECT 93.495 38.410 94.205 38.520 ;
        RECT 87.045 32.160 87.365 32.180 ;
        RECT 88.725 32.160 89.855 33.380 ;
        RECT 90.575 33.370 90.905 38.390 ;
        RECT 93.495 37.040 93.725 38.410 ;
        RECT 93.935 38.160 94.205 38.410 ;
        RECT 94.835 38.780 95.125 39.020 ;
        RECT 96.245 38.780 96.935 38.800 ;
        RECT 94.835 38.340 96.935 38.780 ;
        RECT 94.835 38.150 95.125 38.340 ;
        RECT 94.205 37.600 94.825 37.960 ;
        RECT 96.245 37.630 96.935 38.340 ;
        RECT 93.425 36.440 93.805 37.040 ;
        RECT 94.215 36.730 94.645 37.600 ;
        RECT 93.495 35.250 93.725 36.440 ;
        RECT 94.215 36.310 96.095 36.730 ;
        RECT 94.215 35.780 94.645 36.310 ;
        RECT 94.065 35.420 94.685 35.780 ;
        RECT 93.495 35.240 93.975 35.250 ;
        RECT 93.495 34.560 94.055 35.240 ;
        RECT 93.585 34.410 94.055 34.560 ;
        RECT 93.785 33.460 94.055 34.410 ;
        RECT 94.695 34.160 94.965 35.160 ;
        RECT 94.695 33.430 95.205 34.160 ;
        RECT 94.695 33.340 95.195 33.430 ;
        RECT 90.055 32.790 90.585 33.170 ;
        RECT 87.045 31.110 89.875 32.160 ;
        RECT 90.155 31.910 90.415 32.790 ;
        RECT 90.135 31.290 90.495 31.910 ;
        RECT 94.945 31.220 95.195 33.340 ;
        RECT 87.045 30.200 87.365 31.110 ;
        RECT 88.725 31.100 89.855 31.110 ;
        RECT 90.755 30.820 95.395 31.220 ;
        RECT 94.945 30.540 95.195 30.820 ;
        RECT 87.045 30.140 87.375 30.200 ;
        RECT 87.055 20.210 87.375 30.140 ;
        RECT 88.375 28.890 88.645 30.250 ;
        RECT 89.505 28.890 89.775 30.210 ;
        RECT 94.815 30.110 95.195 30.540 ;
        RECT 94.815 29.600 95.175 30.110 ;
        RECT 88.375 22.200 89.775 28.890 ;
        RECT 88.375 20.200 88.645 22.200 ;
        RECT 89.505 20.160 89.775 22.200 ;
        RECT 94.825 21.760 95.085 29.600 ;
        RECT 94.825 20.210 95.205 21.760 ;
        RECT 87.345 19.550 88.395 19.960 ;
        RECT 89.755 19.560 94.805 19.940 ;
        RECT 87.515 18.270 88.185 19.550 ;
        RECT 87.345 17.590 88.465 18.270 ;
        RECT 73.865 12.750 74.725 13.590 ;
        RECT 61.415 10.960 63.435 12.160 ;
        RECT 72.725 10.990 74.745 12.190 ;
        RECT 84.465 12.180 84.875 14.780 ;
        RECT 85.175 13.580 85.715 16.810 ;
        RECT 91.435 16.780 93.365 19.560 ;
        RECT 90.855 15.930 93.565 16.780 ;
        RECT 94.945 15.390 95.205 20.210 ;
        RECT 94.415 14.660 95.305 15.390 ;
        RECT 95.705 14.800 96.095 36.310 ;
        RECT 96.435 16.830 96.935 37.630 ;
        RECT 98.975 38.500 99.255 40.490 ;
        RECT 101.545 40.420 102.645 41.190 ;
        RECT 110.155 40.530 110.455 42.260 ;
        RECT 99.525 39.660 99.905 40.260 ;
        RECT 99.555 39.040 99.805 39.660 ;
        RECT 99.425 38.660 99.905 39.040 ;
        RECT 98.975 33.430 99.305 38.500 ;
        RECT 99.855 37.640 100.155 38.500 ;
        RECT 100.935 37.640 101.235 38.500 ;
        RECT 101.845 38.460 102.125 40.420 ;
        RECT 105.145 38.850 105.415 39.020 ;
        RECT 104.755 38.540 105.415 38.850 ;
        RECT 99.855 33.400 101.235 37.640 ;
        RECT 101.785 38.410 102.125 38.460 ;
        RECT 104.705 38.430 105.415 38.540 ;
        RECT 98.255 32.180 98.575 32.200 ;
        RECT 99.935 32.180 101.065 33.400 ;
        RECT 101.785 33.390 102.115 38.410 ;
        RECT 104.705 37.060 104.935 38.430 ;
        RECT 105.145 38.180 105.415 38.430 ;
        RECT 106.045 38.800 106.335 39.040 ;
        RECT 107.455 38.800 108.145 38.820 ;
        RECT 106.045 38.360 108.145 38.800 ;
        RECT 106.045 38.170 106.335 38.360 ;
        RECT 105.415 37.620 106.035 37.980 ;
        RECT 107.455 37.650 108.145 38.360 ;
        RECT 104.635 36.460 105.015 37.060 ;
        RECT 105.425 36.750 105.855 37.620 ;
        RECT 104.705 35.270 104.935 36.460 ;
        RECT 105.425 36.330 107.305 36.750 ;
        RECT 105.425 35.800 105.855 36.330 ;
        RECT 105.275 35.440 105.895 35.800 ;
        RECT 104.705 35.260 105.185 35.270 ;
        RECT 104.705 34.580 105.265 35.260 ;
        RECT 104.795 34.430 105.265 34.580 ;
        RECT 104.995 33.480 105.265 34.430 ;
        RECT 105.905 34.180 106.175 35.180 ;
        RECT 105.905 33.450 106.415 34.180 ;
        RECT 105.905 33.360 106.405 33.450 ;
        RECT 101.265 32.810 101.795 33.190 ;
        RECT 98.255 31.130 101.085 32.180 ;
        RECT 101.365 31.930 101.625 32.810 ;
        RECT 101.345 31.310 101.705 31.930 ;
        RECT 106.155 31.240 106.405 33.360 ;
        RECT 98.255 30.220 98.575 31.130 ;
        RECT 99.935 31.120 101.065 31.130 ;
        RECT 101.965 30.840 106.605 31.240 ;
        RECT 106.155 30.560 106.405 30.840 ;
        RECT 98.255 30.160 98.585 30.220 ;
        RECT 98.265 20.230 98.585 30.160 ;
        RECT 99.585 28.910 99.855 30.270 ;
        RECT 100.715 28.910 100.985 30.230 ;
        RECT 106.025 30.130 106.405 30.560 ;
        RECT 106.025 29.620 106.385 30.130 ;
        RECT 99.585 22.220 100.985 28.910 ;
        RECT 99.585 20.220 99.855 22.220 ;
        RECT 100.715 20.180 100.985 22.220 ;
        RECT 106.035 21.780 106.295 29.620 ;
        RECT 106.035 20.230 106.415 21.780 ;
        RECT 98.555 19.570 99.605 19.980 ;
        RECT 100.965 19.580 106.015 19.960 ;
        RECT 98.725 18.290 99.395 19.570 ;
        RECT 98.555 17.610 99.675 18.290 ;
        RECT 85.155 12.740 86.015 13.580 ;
        RECT 95.705 12.180 96.115 14.800 ;
        RECT 96.415 13.600 96.955 16.830 ;
        RECT 102.645 16.800 104.575 19.580 ;
        RECT 102.065 15.950 104.775 16.800 ;
        RECT 106.155 15.410 106.415 20.230 ;
        RECT 105.625 14.680 106.515 15.410 ;
        RECT 106.915 14.820 107.305 36.330 ;
        RECT 107.645 16.850 108.145 37.650 ;
        RECT 110.175 38.540 110.455 40.530 ;
        RECT 112.745 40.460 113.845 41.230 ;
        RECT 121.365 40.550 121.665 42.280 ;
        RECT 142.880 42.020 144.100 43.390 ;
        RECT 110.725 39.700 111.105 40.300 ;
        RECT 110.755 39.080 111.005 39.700 ;
        RECT 110.625 38.700 111.105 39.080 ;
        RECT 110.175 33.470 110.505 38.540 ;
        RECT 111.055 37.680 111.355 38.540 ;
        RECT 112.135 37.680 112.435 38.540 ;
        RECT 113.045 38.500 113.325 40.460 ;
        RECT 116.345 38.890 116.615 39.060 ;
        RECT 115.955 38.580 116.615 38.890 ;
        RECT 111.055 33.440 112.435 37.680 ;
        RECT 112.985 38.450 113.325 38.500 ;
        RECT 115.905 38.470 116.615 38.580 ;
        RECT 109.455 32.220 109.775 32.240 ;
        RECT 111.135 32.220 112.265 33.440 ;
        RECT 112.985 33.430 113.315 38.450 ;
        RECT 115.905 37.100 116.135 38.470 ;
        RECT 116.345 38.220 116.615 38.470 ;
        RECT 117.245 38.840 117.535 39.080 ;
        RECT 118.655 38.840 119.345 38.860 ;
        RECT 117.245 38.400 119.345 38.840 ;
        RECT 117.245 38.210 117.535 38.400 ;
        RECT 116.615 37.660 117.235 38.020 ;
        RECT 118.655 37.690 119.345 38.400 ;
        RECT 115.835 36.500 116.215 37.100 ;
        RECT 116.625 36.790 117.055 37.660 ;
        RECT 115.905 35.310 116.135 36.500 ;
        RECT 116.625 36.370 118.505 36.790 ;
        RECT 116.625 35.840 117.055 36.370 ;
        RECT 116.475 35.480 117.095 35.840 ;
        RECT 115.905 35.300 116.385 35.310 ;
        RECT 115.905 34.620 116.465 35.300 ;
        RECT 115.995 34.470 116.465 34.620 ;
        RECT 116.195 33.520 116.465 34.470 ;
        RECT 117.105 34.220 117.375 35.220 ;
        RECT 117.105 33.490 117.615 34.220 ;
        RECT 117.105 33.400 117.605 33.490 ;
        RECT 112.465 32.850 112.995 33.230 ;
        RECT 109.455 31.170 112.285 32.220 ;
        RECT 112.565 31.970 112.825 32.850 ;
        RECT 112.545 31.350 112.905 31.970 ;
        RECT 117.355 31.280 117.605 33.400 ;
        RECT 109.455 30.260 109.775 31.170 ;
        RECT 111.135 31.160 112.265 31.170 ;
        RECT 113.165 30.880 117.805 31.280 ;
        RECT 117.355 30.600 117.605 30.880 ;
        RECT 109.455 30.200 109.785 30.260 ;
        RECT 109.465 20.270 109.785 30.200 ;
        RECT 110.785 28.950 111.055 30.310 ;
        RECT 111.915 28.950 112.185 30.270 ;
        RECT 117.225 30.170 117.605 30.600 ;
        RECT 117.225 29.660 117.585 30.170 ;
        RECT 110.785 22.260 112.185 28.950 ;
        RECT 110.785 20.260 111.055 22.260 ;
        RECT 111.915 20.220 112.185 22.260 ;
        RECT 117.235 21.820 117.495 29.660 ;
        RECT 117.235 20.270 117.615 21.820 ;
        RECT 109.755 19.610 110.805 20.020 ;
        RECT 112.165 19.620 117.215 20.000 ;
        RECT 109.925 18.330 110.595 19.610 ;
        RECT 109.755 17.650 110.875 18.330 ;
        RECT 96.395 12.760 97.255 13.600 ;
        RECT 106.915 12.230 107.325 14.820 ;
        RECT 107.625 13.620 108.165 16.850 ;
        RECT 113.845 16.840 115.775 19.620 ;
        RECT 113.265 15.990 115.975 16.840 ;
        RECT 117.355 15.450 117.615 20.270 ;
        RECT 116.825 14.720 117.715 15.450 ;
        RECT 118.115 14.860 118.505 36.370 ;
        RECT 118.845 16.890 119.345 37.690 ;
        RECT 121.385 38.560 121.665 40.550 ;
        RECT 123.955 40.480 125.055 41.250 ;
        RECT 121.935 39.720 122.315 40.320 ;
        RECT 121.965 39.100 122.215 39.720 ;
        RECT 121.835 38.720 122.315 39.100 ;
        RECT 121.385 33.490 121.715 38.560 ;
        RECT 122.265 37.700 122.565 38.560 ;
        RECT 123.345 37.700 123.645 38.560 ;
        RECT 124.255 38.520 124.535 40.480 ;
        RECT 127.555 38.910 127.825 39.080 ;
        RECT 127.165 38.600 127.825 38.910 ;
        RECT 122.265 33.460 123.645 37.700 ;
        RECT 124.195 38.470 124.535 38.520 ;
        RECT 127.115 38.490 127.825 38.600 ;
        RECT 120.665 32.240 120.985 32.260 ;
        RECT 122.345 32.240 123.475 33.460 ;
        RECT 124.195 33.450 124.525 38.470 ;
        RECT 127.115 37.120 127.345 38.490 ;
        RECT 127.555 38.240 127.825 38.490 ;
        RECT 128.455 38.860 128.745 39.100 ;
        RECT 142.940 38.950 144.100 42.020 ;
        RECT 129.865 38.860 130.555 38.880 ;
        RECT 128.455 38.420 130.555 38.860 ;
        RECT 128.455 38.230 128.745 38.420 ;
        RECT 127.825 37.680 128.445 38.040 ;
        RECT 129.865 37.710 130.555 38.420 ;
        RECT 127.045 36.520 127.425 37.120 ;
        RECT 127.835 36.810 128.265 37.680 ;
        RECT 127.115 35.330 127.345 36.520 ;
        RECT 127.835 36.390 129.715 36.810 ;
        RECT 127.835 35.860 128.265 36.390 ;
        RECT 127.685 35.500 128.305 35.860 ;
        RECT 127.115 35.320 127.595 35.330 ;
        RECT 127.115 34.640 127.675 35.320 ;
        RECT 127.205 34.490 127.675 34.640 ;
        RECT 127.405 33.540 127.675 34.490 ;
        RECT 128.315 34.240 128.585 35.240 ;
        RECT 128.315 33.510 128.825 34.240 ;
        RECT 128.315 33.420 128.815 33.510 ;
        RECT 123.675 32.870 124.205 33.250 ;
        RECT 120.665 31.190 123.495 32.240 ;
        RECT 123.775 31.990 124.035 32.870 ;
        RECT 123.755 31.370 124.115 31.990 ;
        RECT 128.565 31.300 128.815 33.420 ;
        RECT 120.665 30.280 120.985 31.190 ;
        RECT 122.345 31.180 123.475 31.190 ;
        RECT 124.375 30.900 129.015 31.300 ;
        RECT 128.565 30.620 128.815 30.900 ;
        RECT 120.665 30.220 120.995 30.280 ;
        RECT 120.675 20.290 120.995 30.220 ;
        RECT 121.995 28.970 122.265 30.330 ;
        RECT 123.125 28.970 123.395 30.290 ;
        RECT 128.435 30.190 128.815 30.620 ;
        RECT 128.435 29.680 128.795 30.190 ;
        RECT 121.995 22.280 123.395 28.970 ;
        RECT 121.995 20.280 122.265 22.280 ;
        RECT 123.125 20.240 123.395 22.280 ;
        RECT 128.445 21.840 128.705 29.680 ;
        RECT 128.445 20.290 128.825 21.840 ;
        RECT 120.965 19.630 122.015 20.040 ;
        RECT 123.375 19.640 128.425 20.020 ;
        RECT 121.135 18.350 121.805 19.630 ;
        RECT 120.965 17.670 122.085 18.350 ;
        RECT 107.605 12.780 108.465 13.620 ;
        RECT 118.115 12.230 118.525 14.860 ;
        RECT 118.825 13.660 119.365 16.890 ;
        RECT 125.055 16.860 126.985 19.640 ;
        RECT 124.475 16.010 127.185 16.860 ;
        RECT 128.565 15.470 128.825 20.290 ;
        RECT 128.035 14.740 128.925 15.470 ;
        RECT 129.325 14.880 129.715 36.390 ;
        RECT 130.055 16.910 130.555 37.710 ;
        RECT 142.900 37.580 144.120 38.950 ;
        RECT 132.395 24.340 132.705 30.230 ;
        RECT 132.195 20.120 132.705 24.340 ;
        RECT 118.805 12.820 119.665 13.660 ;
        RECT 129.325 12.260 129.735 14.880 ;
        RECT 130.035 13.680 130.575 16.910 ;
        RECT 132.195 15.510 132.505 20.120 ;
        RECT 137.715 19.980 138.005 30.170 ;
        RECT 132.685 19.590 138.005 19.980 ;
        RECT 137.715 16.940 138.005 19.590 ;
        RECT 142.940 17.940 144.090 19.160 ;
        RECT 145.080 18.760 146.200 18.930 ;
        RECT 137.395 15.890 138.295 16.940 ;
        RECT 137.715 15.720 138.005 15.890 ;
        RECT 131.975 14.270 132.735 15.510 ;
        RECT 142.940 15.090 144.050 17.940 ;
        RECT 142.900 13.870 144.050 15.090 ;
        RECT 145.070 14.920 146.200 18.760 ;
        RECT 145.030 13.970 146.200 14.920 ;
        RECT 145.030 13.900 146.150 13.970 ;
        RECT 130.015 12.840 130.875 13.680 ;
        RECT 83.845 10.980 85.865 12.180 ;
        RECT 95.145 10.980 97.165 12.180 ;
        RECT 106.335 11.030 108.355 12.230 ;
        RECT 117.565 11.030 119.585 12.230 ;
        RECT 128.865 11.060 130.885 12.260 ;
        RECT 74.340 0.110 75.630 1.460 ;
        RECT 93.550 0.180 94.840 1.530 ;
        RECT 112.950 0.310 114.240 1.660 ;
        RECT 131.850 0.380 133.490 1.930 ;
        RECT 151.650 0.250 152.920 1.470 ;
      LAYER met3 ;
        RECT 135.340 223.855 136.790 225.205 ;
        RECT 138.130 223.785 139.580 225.135 ;
        RECT 143.180 223.815 144.630 225.165 ;
        RECT 10.660 214.270 12.240 214.600 ;
        RECT 37.450 214.270 39.030 214.600 ;
        RECT 64.240 214.270 65.820 214.600 ;
        RECT 91.030 214.270 92.610 214.600 ;
        RECT 24.055 211.550 25.635 211.880 ;
        RECT 50.845 211.550 52.425 211.880 ;
        RECT 77.635 211.550 79.215 211.880 ;
        RECT 104.425 211.550 106.005 211.880 ;
        RECT 10.660 208.830 12.240 209.160 ;
        RECT 37.450 208.830 39.030 209.160 ;
        RECT 64.240 208.830 65.820 209.160 ;
        RECT 91.030 208.830 92.610 209.160 ;
        RECT 24.055 206.110 25.635 206.440 ;
        RECT 50.845 206.110 52.425 206.440 ;
        RECT 77.635 206.110 79.215 206.440 ;
        RECT 104.425 206.110 106.005 206.440 ;
        RECT 10.660 203.390 12.240 203.720 ;
        RECT 37.450 203.390 39.030 203.720 ;
        RECT 64.240 203.390 65.820 203.720 ;
        RECT 91.030 203.390 92.610 203.720 ;
        RECT 24.055 200.670 25.635 201.000 ;
        RECT 50.845 200.670 52.425 201.000 ;
        RECT 77.635 200.670 79.215 201.000 ;
        RECT 104.425 200.670 106.005 201.000 ;
        RECT 95.880 198.605 96.260 198.615 ;
        RECT 96.595 198.605 96.925 198.620 ;
        RECT 95.880 198.305 96.925 198.605 ;
        RECT 95.880 198.295 96.260 198.305 ;
        RECT 96.595 198.290 96.925 198.305 ;
        RECT 10.660 197.950 12.240 198.280 ;
        RECT 37.450 197.950 39.030 198.280 ;
        RECT 64.240 197.950 65.820 198.280 ;
        RECT 91.030 197.950 92.610 198.280 ;
        RECT 24.055 195.230 25.635 195.560 ;
        RECT 50.845 195.230 52.425 195.560 ;
        RECT 77.635 195.230 79.215 195.560 ;
        RECT 104.425 195.230 106.005 195.560 ;
        RECT 10.660 192.510 12.240 192.840 ;
        RECT 37.450 192.510 39.030 192.840 ;
        RECT 64.240 192.510 65.820 192.840 ;
        RECT 91.030 192.510 92.610 192.840 ;
        RECT 24.055 189.790 25.635 190.120 ;
        RECT 50.845 189.790 52.425 190.120 ;
        RECT 77.635 189.790 79.215 190.120 ;
        RECT 104.425 189.790 106.005 190.120 ;
        RECT 10.660 187.070 12.240 187.400 ;
        RECT 37.450 187.070 39.030 187.400 ;
        RECT 64.240 187.070 65.820 187.400 ;
        RECT 91.030 187.070 92.610 187.400 ;
        RECT 24.055 184.350 25.635 184.680 ;
        RECT 50.845 184.350 52.425 184.680 ;
        RECT 77.635 184.350 79.215 184.680 ;
        RECT 104.425 184.350 106.005 184.680 ;
        RECT 83.920 182.965 84.300 182.975 ;
        RECT 84.635 182.965 84.965 182.980 ;
        RECT 83.920 182.665 84.965 182.965 ;
        RECT 83.920 182.655 84.300 182.665 ;
        RECT 84.635 182.650 84.965 182.665 ;
        RECT 10.660 181.630 12.240 181.960 ;
        RECT 37.450 181.630 39.030 181.960 ;
        RECT 64.240 181.630 65.820 181.960 ;
        RECT 91.030 181.630 92.610 181.960 ;
        RECT 83.920 180.925 84.300 180.935 ;
        RECT 103.955 180.925 104.285 180.940 ;
        RECT 83.920 180.625 104.285 180.925 ;
        RECT 83.920 180.615 84.300 180.625 ;
        RECT 103.955 180.610 104.285 180.625 ;
        RECT 24.055 178.910 25.635 179.240 ;
        RECT 50.845 178.910 52.425 179.240 ;
        RECT 77.635 178.910 79.215 179.240 ;
        RECT 104.425 178.910 106.005 179.240 ;
        RECT 10.660 176.190 12.240 176.520 ;
        RECT 37.450 176.190 39.030 176.520 ;
        RECT 64.240 176.190 65.820 176.520 ;
        RECT 91.030 176.190 92.610 176.520 ;
        RECT 83.920 176.165 84.300 176.175 ;
        RECT 66.480 175.865 84.300 176.165 ;
        RECT 27.595 175.485 27.925 175.500 ;
        RECT 39.095 175.485 39.425 175.500 ;
        RECT 58.415 175.485 58.745 175.500 ;
        RECT 66.480 175.485 66.780 175.865 ;
        RECT 83.920 175.855 84.300 175.865 ;
        RECT 27.595 175.185 66.780 175.485 ;
        RECT 27.595 175.170 27.925 175.185 ;
        RECT 39.095 175.170 39.425 175.185 ;
        RECT 58.415 175.170 58.745 175.185 ;
        RECT 34.240 174.805 34.620 174.815 ;
        RECT 36.335 174.805 36.665 174.820 ;
        RECT 34.240 174.505 36.665 174.805 ;
        RECT 34.240 174.495 34.620 174.505 ;
        RECT 36.335 174.490 36.665 174.505 ;
        RECT 39.555 174.805 39.885 174.820 ;
        RECT 49.675 174.805 50.005 174.820 ;
        RECT 39.555 174.505 50.005 174.805 ;
        RECT 39.555 174.490 39.885 174.505 ;
        RECT 49.675 174.490 50.005 174.505 ;
        RECT 115.455 174.805 115.785 174.820 ;
        RECT 119.370 174.805 121.370 174.955 ;
        RECT 115.455 174.505 121.370 174.805 ;
        RECT 115.455 174.490 115.785 174.505 ;
        RECT 119.370 174.355 121.370 174.505 ;
        RECT 24.055 173.470 25.635 173.800 ;
        RECT 50.845 173.470 52.425 173.800 ;
        RECT 77.635 173.470 79.215 173.800 ;
        RECT 104.425 173.470 106.005 173.800 ;
        RECT 133.700 172.500 134.930 172.705 ;
        RECT 72.215 171.415 72.545 171.420 ;
        RECT 71.960 171.405 72.545 171.415 ;
        RECT 71.960 171.105 72.770 171.405 ;
        RECT 71.960 171.095 72.545 171.105 ;
        RECT 72.215 171.090 72.545 171.095 ;
        RECT 10.660 170.750 12.240 171.080 ;
        RECT 37.450 170.750 39.030 171.080 ;
        RECT 64.240 170.750 65.820 171.080 ;
        RECT 91.030 170.750 92.610 171.080 ;
        RECT 129.030 170.130 134.930 172.500 ;
        RECT 133.700 170.095 134.930 170.130 ;
        RECT 68.995 169.365 69.325 169.380 ;
        RECT 72.675 169.365 73.005 169.380 ;
        RECT 68.995 169.065 73.005 169.365 ;
        RECT 68.995 169.050 69.325 169.065 ;
        RECT 72.675 169.050 73.005 169.065 ;
        RECT 24.055 168.030 25.635 168.360 ;
        RECT 50.845 168.030 52.425 168.360 ;
        RECT 77.635 168.030 79.215 168.360 ;
        RECT 104.425 168.030 106.005 168.360 ;
        RECT 10.660 165.310 12.240 165.640 ;
        RECT 37.450 165.310 39.030 165.640 ;
        RECT 64.240 165.310 65.820 165.640 ;
        RECT 91.030 165.310 92.610 165.640 ;
        RECT 41.855 164.605 42.185 164.620 ;
        RECT 46.455 164.605 46.785 164.620 ;
        RECT 41.855 164.305 46.785 164.605 ;
        RECT 41.855 164.290 42.185 164.305 ;
        RECT 46.455 164.290 46.785 164.305 ;
        RECT 24.055 162.590 25.635 162.920 ;
        RECT 50.845 162.590 52.425 162.920 ;
        RECT 77.635 162.590 79.215 162.920 ;
        RECT 104.425 162.590 106.005 162.920 ;
        RECT 42.315 161.885 42.645 161.900 ;
        RECT 50.135 161.885 50.465 161.900 ;
        RECT 68.075 161.885 68.405 161.900 ;
        RECT 42.315 161.585 50.465 161.885 ;
        RECT 42.315 161.570 42.645 161.585 ;
        RECT 50.135 161.570 50.465 161.585 ;
        RECT 50.840 161.585 68.405 161.885 ;
        RECT 36.795 161.205 37.125 161.220 ;
        RECT 38.635 161.205 38.965 161.220 ;
        RECT 50.840 161.205 51.140 161.585 ;
        RECT 68.075 161.570 68.405 161.585 ;
        RECT 94.295 161.885 94.625 161.900 ;
        RECT 95.880 161.885 96.260 161.895 ;
        RECT 94.295 161.585 96.260 161.885 ;
        RECT 94.295 161.570 94.625 161.585 ;
        RECT 95.880 161.575 96.260 161.585 ;
        RECT 36.795 160.905 51.140 161.205 ;
        RECT 51.975 161.205 52.305 161.220 ;
        RECT 54.735 161.205 55.065 161.220 ;
        RECT 51.975 160.905 55.065 161.205 ;
        RECT 36.795 160.890 37.125 160.905 ;
        RECT 38.635 160.890 38.965 160.905 ;
        RECT 51.975 160.890 52.305 160.905 ;
        RECT 54.735 160.890 55.065 160.905 ;
        RECT 10.660 159.870 12.240 160.200 ;
        RECT 37.450 159.870 39.030 160.200 ;
        RECT 64.240 159.870 65.820 160.200 ;
        RECT 91.030 159.870 92.610 160.200 ;
        RECT 73.595 159.855 73.925 159.860 ;
        RECT 73.595 159.845 74.180 159.855 ;
        RECT 73.370 159.545 74.180 159.845 ;
        RECT 73.595 159.535 74.180 159.545 ;
        RECT 73.595 159.530 73.925 159.535 ;
        RECT 32.400 157.805 32.780 157.815 ;
        RECT 46.915 157.805 47.245 157.820 ;
        RECT 32.400 157.505 47.245 157.805 ;
        RECT 32.400 157.495 32.780 157.505 ;
        RECT 46.915 157.490 47.245 157.505 ;
        RECT 58.415 157.805 58.745 157.820 ;
        RECT 59.335 157.815 59.665 157.820 ;
        RECT 59.080 157.805 59.665 157.815 ;
        RECT 73.135 157.805 73.465 157.820 ;
        RECT 58.415 157.505 59.665 157.805 ;
        RECT 58.415 157.490 58.745 157.505 ;
        RECT 59.080 157.495 59.665 157.505 ;
        RECT 59.335 157.490 59.665 157.495 ;
        RECT 72.920 157.490 73.465 157.805 ;
        RECT 24.055 157.150 25.635 157.480 ;
        RECT 50.845 157.150 52.425 157.480 ;
        RECT 10.660 154.430 12.240 154.760 ;
        RECT 37.450 154.430 39.030 154.760 ;
        RECT 64.240 154.430 65.820 154.760 ;
        RECT 72.920 154.420 73.220 157.490 ;
        RECT 77.635 157.150 79.215 157.480 ;
        RECT 104.425 157.150 106.005 157.480 ;
        RECT 74.515 157.125 74.845 157.140 ;
        RECT 74.515 156.825 76.900 157.125 ;
        RECT 74.515 156.810 74.845 156.825 ;
        RECT 76.600 156.445 76.900 156.825 ;
        RECT 96.135 156.445 96.465 156.460 ;
        RECT 76.600 156.145 96.465 156.445 ;
        RECT 96.135 156.130 96.465 156.145 ;
        RECT 91.030 154.430 92.610 154.760 ;
        RECT 72.920 154.105 73.465 154.420 ;
        RECT 73.135 154.090 73.465 154.105 ;
        RECT 54.735 153.045 55.065 153.060 ;
        RECT 62.095 153.045 62.425 153.060 ;
        RECT 54.735 152.745 62.425 153.045 ;
        RECT 54.735 152.730 55.065 152.745 ;
        RECT 62.095 152.730 62.425 152.745 ;
        RECT 73.135 153.045 73.465 153.060 ;
        RECT 73.800 153.045 74.180 153.055 ;
        RECT 73.135 152.745 74.180 153.045 ;
        RECT 73.135 152.730 73.465 152.745 ;
        RECT 73.800 152.735 74.180 152.745 ;
        RECT 24.055 151.710 25.635 152.040 ;
        RECT 50.845 151.710 52.425 152.040 ;
        RECT 77.635 151.710 79.215 152.040 ;
        RECT 104.425 151.710 106.005 152.040 ;
        RECT 10.660 148.990 12.240 149.320 ;
        RECT 37.450 148.990 39.030 149.320 ;
        RECT 64.240 148.990 65.820 149.320 ;
        RECT 91.030 148.990 92.610 149.320 ;
        RECT 66.235 147.605 66.565 147.620 ;
        RECT 119.370 147.605 121.370 147.755 ;
        RECT 66.235 147.305 121.370 147.605 ;
        RECT 66.235 147.290 66.565 147.305 ;
        RECT 119.370 147.155 121.370 147.305 ;
        RECT 31.275 146.925 31.605 146.940 ;
        RECT 37.255 146.925 37.585 146.940 ;
        RECT 31.275 146.625 37.585 146.925 ;
        RECT 31.275 146.610 31.605 146.625 ;
        RECT 37.255 146.610 37.585 146.625 ;
        RECT 24.055 146.270 25.635 146.600 ;
        RECT 50.845 146.270 52.425 146.600 ;
        RECT 77.635 146.270 79.215 146.600 ;
        RECT 104.425 146.270 106.005 146.600 ;
        RECT 10.660 143.550 12.240 143.880 ;
        RECT 37.450 143.550 39.030 143.880 ;
        RECT 64.240 143.550 65.820 143.880 ;
        RECT 91.030 143.550 92.610 143.880 ;
        RECT 32.655 142.165 32.985 142.180 ;
        RECT 61.635 142.165 61.965 142.180 ;
        RECT 32.655 141.865 61.965 142.165 ;
        RECT 32.655 141.850 32.985 141.865 ;
        RECT 61.635 141.850 61.965 141.865 ;
        RECT 24.055 140.830 25.635 141.160 ;
        RECT 50.845 140.830 52.425 141.160 ;
        RECT 77.635 140.830 79.215 141.160 ;
        RECT 104.425 140.830 106.005 141.160 ;
        RECT 33.575 140.805 33.905 140.820 ;
        RECT 34.240 140.805 34.620 140.815 ;
        RECT 33.575 140.505 34.620 140.805 ;
        RECT 33.575 140.490 33.905 140.505 ;
        RECT 34.240 140.495 34.620 140.505 ;
        RECT 70.375 140.805 70.705 140.820 ;
        RECT 71.960 140.805 72.340 140.815 ;
        RECT 70.375 140.505 72.340 140.805 ;
        RECT 70.375 140.490 70.705 140.505 ;
        RECT 71.960 140.495 72.340 140.505 ;
        RECT 47.375 139.445 47.705 139.460 ;
        RECT 51.055 139.445 51.385 139.460 ;
        RECT 47.375 139.145 51.385 139.445 ;
        RECT 47.375 139.130 47.705 139.145 ;
        RECT 51.055 139.130 51.385 139.145 ;
        RECT 10.660 138.110 12.240 138.440 ;
        RECT 37.450 138.110 39.030 138.440 ;
        RECT 64.240 138.110 65.820 138.440 ;
        RECT 91.030 138.110 92.610 138.440 ;
        RECT 132.510 138.165 135.210 140.035 ;
        RECT 24.055 135.390 25.635 135.720 ;
        RECT 50.845 135.390 52.425 135.720 ;
        RECT 77.635 135.390 79.215 135.720 ;
        RECT 104.425 135.390 106.005 135.720 ;
        RECT 10.660 132.670 12.240 133.000 ;
        RECT 37.450 132.670 39.030 133.000 ;
        RECT 64.240 132.670 65.820 133.000 ;
        RECT 91.030 132.670 92.610 133.000 ;
        RECT 24.055 129.950 25.635 130.280 ;
        RECT 50.845 129.950 52.425 130.280 ;
        RECT 77.635 129.950 79.215 130.280 ;
        RECT 104.425 129.950 106.005 130.280 ;
        RECT 58.160 128.565 58.540 128.575 ;
        RECT 88.775 128.565 89.105 128.580 ;
        RECT 58.160 128.265 89.105 128.565 ;
        RECT 58.160 128.255 58.540 128.265 ;
        RECT 10.660 127.230 12.240 127.560 ;
        RECT 37.450 127.230 39.030 127.560 ;
        RECT 52.895 127.205 53.225 127.220 ;
        RECT 58.200 127.205 58.500 128.255 ;
        RECT 88.775 128.250 89.105 128.265 ;
        RECT 64.240 127.230 65.820 127.560 ;
        RECT 91.030 127.230 92.610 127.560 ;
        RECT 52.895 126.905 58.500 127.205 ;
        RECT 52.895 126.890 53.225 126.905 ;
        RECT 24.055 124.510 25.635 124.840 ;
        RECT 50.845 124.510 52.425 124.840 ;
        RECT 77.635 124.510 79.215 124.840 ;
        RECT 104.425 124.510 106.005 124.840 ;
        RECT 27.595 123.125 27.925 123.140 ;
        RECT 52.895 123.125 53.225 123.140 ;
        RECT 27.595 122.825 53.225 123.125 ;
        RECT 27.595 122.810 27.925 122.825 ;
        RECT 52.895 122.810 53.225 122.825 ;
        RECT 10.660 121.790 12.240 122.120 ;
        RECT 37.450 121.790 39.030 122.120 ;
        RECT 64.240 121.790 65.820 122.120 ;
        RECT 91.030 121.790 92.610 122.120 ;
        RECT 32.195 120.415 32.525 120.420 ;
        RECT 32.195 120.405 32.780 120.415 ;
        RECT 116.835 120.405 117.165 120.420 ;
        RECT 119.370 120.405 121.370 120.555 ;
        RECT 32.195 120.105 32.980 120.405 ;
        RECT 116.835 120.105 121.370 120.405 ;
        RECT 32.195 120.095 32.780 120.105 ;
        RECT 32.195 120.090 32.525 120.095 ;
        RECT 116.835 120.090 117.165 120.105 ;
        RECT 119.370 119.955 121.370 120.105 ;
        RECT 24.055 119.070 25.635 119.400 ;
        RECT 50.845 119.070 52.425 119.400 ;
        RECT 77.635 119.070 79.215 119.400 ;
        RECT 104.425 119.070 106.005 119.400 ;
        RECT 10.660 116.350 12.240 116.680 ;
        RECT 37.450 116.350 39.030 116.680 ;
        RECT 64.240 116.350 65.820 116.680 ;
        RECT 91.030 116.350 92.610 116.680 ;
        RECT 24.055 113.630 25.635 113.960 ;
        RECT 50.845 113.630 52.425 113.960 ;
        RECT 77.635 113.630 79.215 113.960 ;
        RECT 104.425 113.630 106.005 113.960 ;
        RECT 10.660 110.910 12.240 111.240 ;
        RECT 37.450 110.910 39.030 111.240 ;
        RECT 64.240 110.910 65.820 111.240 ;
        RECT 91.030 110.910 92.610 111.240 ;
        RECT 24.055 108.190 25.635 108.520 ;
        RECT 50.845 108.190 52.425 108.520 ;
        RECT 77.635 108.190 79.215 108.520 ;
        RECT 104.425 108.190 106.005 108.520 ;
        RECT 129.700 105.605 133.210 106.625 ;
        RECT 37.630 88.620 38.970 88.755 ;
        RECT 13.950 87.980 14.980 88.515 ;
        RECT 13.950 87.500 14.990 87.980 ;
        RECT 13.950 87.175 14.980 87.500 ;
        RECT 14.070 86.570 14.810 87.175 ;
        RECT 20.050 87.105 20.920 88.515 ;
        RECT 14.070 75.715 14.700 86.570 ;
        RECT 20.170 77.115 20.800 87.105 ;
        RECT 25.910 87.055 26.860 88.515 ;
        RECT 26.070 78.385 26.700 87.055 ;
        RECT 31.730 86.965 32.910 88.585 ;
        RECT 32.005 79.615 32.635 86.965 ;
        RECT 37.630 86.835 39.120 88.620 ;
        RECT 38.060 81.125 38.690 86.835 ;
        RECT 43.790 86.745 45.190 88.605 ;
        RECT 49.710 86.945 51.060 88.615 ;
        RECT 44.175 82.625 44.805 86.745 ;
        RECT 50.070 83.875 50.700 86.945 ;
        RECT 55.530 86.785 56.750 88.545 ;
        RECT 55.825 85.115 56.455 86.785 ;
        RECT 61.670 86.625 63.180 88.615 ;
        RECT 67.680 88.305 68.720 89.815 ;
        RECT 67.885 87.225 68.515 88.305 ;
        RECT 62.110 86.175 62.740 86.625 ;
        RECT 67.885 86.595 130.605 87.225 ;
        RECT 62.110 85.545 118.855 86.175 ;
        RECT 55.825 84.485 107.605 85.115 ;
        RECT 50.070 83.245 96.285 83.875 ;
        RECT 44.175 81.995 85.055 82.625 ;
        RECT 38.060 80.495 73.765 81.125 ;
        RECT 32.005 78.985 62.635 79.615 ;
        RECT 26.070 77.755 51.245 78.385 ;
        RECT 20.170 76.485 40.645 77.115 ;
        RECT 14.070 75.660 29.295 75.715 ;
        RECT 40.015 75.710 40.645 76.485 ;
        RECT 14.070 75.085 30.410 75.660 ;
        RECT 27.850 74.670 30.410 75.085 ;
        RECT 3.910 71.345 6.100 73.215 ;
        RECT 27.850 73.120 30.450 74.670 ;
        RECT 39.060 74.510 41.620 75.710 ;
        RECT 50.615 75.580 51.245 77.755 ;
        RECT 62.005 75.690 62.635 78.985 ;
        RECT 49.930 74.650 52.490 75.580 ;
        RECT 0.970 70.330 3.070 70.430 ;
        RECT 15.510 70.330 17.040 71.185 ;
        RECT 0.960 68.750 17.040 70.330 ;
        RECT 0.970 68.710 3.070 68.750 ;
        RECT 15.510 68.635 17.040 68.750 ;
        RECT 20.145 54.060 20.605 54.135 ;
        RECT 25.715 54.060 26.175 54.085 ;
        RECT 20.145 53.620 26.175 54.060 ;
        RECT 20.145 53.565 20.605 53.620 ;
        RECT 25.715 53.515 26.175 53.620 ;
        RECT 22.405 48.870 22.885 48.935 ;
        RECT 22.405 48.550 24.205 48.870 ;
        RECT 22.405 48.385 22.885 48.550 ;
        RECT 23.635 45.710 24.195 48.550 ;
        RECT 27.515 45.710 27.995 45.735 ;
        RECT 23.635 45.290 27.995 45.710 ;
        RECT 23.635 45.280 24.195 45.290 ;
        RECT 27.515 45.185 27.995 45.290 ;
        RECT 20.745 40.120 21.225 40.225 ;
        RECT 24.545 40.120 25.105 40.130 ;
        RECT 20.745 39.700 25.105 40.120 ;
        RECT 20.745 39.675 21.225 39.700 ;
        RECT 24.545 36.860 25.105 39.700 ;
        RECT 25.855 36.860 26.335 37.025 ;
        RECT 24.535 36.540 26.335 36.860 ;
        RECT 25.855 36.475 26.335 36.540 ;
        RECT 22.565 31.790 23.025 31.895 ;
        RECT 28.135 31.790 28.595 31.845 ;
        RECT 22.565 31.350 28.595 31.790 ;
        RECT 22.565 31.325 23.025 31.350 ;
        RECT 28.135 31.275 28.595 31.350 ;
        RECT 29.765 12.265 30.255 73.120 ;
        RECT 38.960 73.080 41.730 74.510 ;
        RECT 31.345 54.070 31.805 54.145 ;
        RECT 36.915 54.070 37.375 54.095 ;
        RECT 31.345 53.630 37.375 54.070 ;
        RECT 31.345 53.575 31.805 53.630 ;
        RECT 36.915 53.525 37.375 53.630 ;
        RECT 33.605 48.880 34.085 48.945 ;
        RECT 33.605 48.560 35.405 48.880 ;
        RECT 33.605 48.395 34.085 48.560 ;
        RECT 34.835 45.720 35.395 48.560 ;
        RECT 38.715 45.720 39.195 45.745 ;
        RECT 34.835 45.300 39.195 45.720 ;
        RECT 34.835 45.290 35.395 45.300 ;
        RECT 38.715 45.195 39.195 45.300 ;
        RECT 32.025 40.120 32.505 40.225 ;
        RECT 35.825 40.120 36.385 40.130 ;
        RECT 32.025 39.700 36.385 40.120 ;
        RECT 32.025 39.675 32.505 39.700 ;
        RECT 35.825 36.860 36.385 39.700 ;
        RECT 37.135 36.860 37.615 37.025 ;
        RECT 35.815 36.540 37.615 36.860 ;
        RECT 37.135 36.475 37.615 36.540 ;
        RECT 33.845 31.790 34.305 31.895 ;
        RECT 39.415 31.790 39.875 31.845 ;
        RECT 33.845 31.350 39.875 31.790 ;
        RECT 33.845 31.325 34.305 31.350 ;
        RECT 39.415 31.275 39.875 31.350 ;
        RECT 41.055 12.360 41.545 73.080 ;
        RECT 49.930 73.030 52.530 74.650 ;
        RECT 61.330 74.530 63.890 75.690 ;
        RECT 73.135 75.580 73.765 80.495 ;
        RECT 84.425 75.690 85.055 81.995 ;
        RECT 72.340 74.980 74.900 75.580 ;
        RECT 42.565 54.040 43.025 54.115 ;
        RECT 48.135 54.040 48.595 54.065 ;
        RECT 42.565 53.600 48.595 54.040 ;
        RECT 42.565 53.545 43.025 53.600 ;
        RECT 48.135 53.495 48.595 53.600 ;
        RECT 44.825 48.850 45.305 48.915 ;
        RECT 44.825 48.530 46.625 48.850 ;
        RECT 44.825 48.365 45.305 48.530 ;
        RECT 46.055 45.690 46.615 48.530 ;
        RECT 49.935 45.690 50.415 45.715 ;
        RECT 46.055 45.270 50.415 45.690 ;
        RECT 46.055 45.260 46.615 45.270 ;
        RECT 49.935 45.165 50.415 45.270 ;
        RECT 43.315 40.100 43.795 40.205 ;
        RECT 47.115 40.100 47.675 40.110 ;
        RECT 43.315 39.680 47.675 40.100 ;
        RECT 43.315 39.655 43.795 39.680 ;
        RECT 47.115 36.840 47.675 39.680 ;
        RECT 48.425 36.840 48.905 37.005 ;
        RECT 47.105 36.520 48.905 36.840 ;
        RECT 48.425 36.455 48.905 36.520 ;
        RECT 45.135 31.770 45.595 31.875 ;
        RECT 50.705 31.770 51.165 31.825 ;
        RECT 45.135 31.330 51.165 31.770 ;
        RECT 45.135 31.305 45.595 31.330 ;
        RECT 50.705 31.255 51.165 31.330 ;
        RECT 41.055 12.350 41.555 12.360 ;
        RECT 28.345 11.115 30.465 12.265 ;
        RECT 41.065 11.965 41.555 12.350 ;
        RECT 51.635 12.145 52.125 73.030 ;
        RECT 61.260 73.010 64.060 74.530 ;
        RECT 72.340 73.050 75.020 74.980 ;
        RECT 83.730 74.540 86.290 75.690 ;
        RECT 95.655 75.580 96.285 83.245 ;
        RECT 106.975 75.640 107.605 84.485 ;
        RECT 118.225 75.650 118.855 85.545 ;
        RECT 129.975 75.650 130.605 86.595 ;
        RECT 133.330 76.605 136.060 77.855 ;
        RECT 137.190 76.585 139.920 77.835 ;
        RECT 53.815 54.020 54.275 54.095 ;
        RECT 59.385 54.020 59.845 54.045 ;
        RECT 53.815 53.580 59.845 54.020 ;
        RECT 53.815 53.525 54.275 53.580 ;
        RECT 59.385 53.475 59.845 53.580 ;
        RECT 56.075 48.830 56.555 48.895 ;
        RECT 56.075 48.510 57.875 48.830 ;
        RECT 56.075 48.345 56.555 48.510 ;
        RECT 57.305 45.670 57.865 48.510 ;
        RECT 61.185 45.670 61.665 45.695 ;
        RECT 57.305 45.250 61.665 45.670 ;
        RECT 57.305 45.240 57.865 45.250 ;
        RECT 61.185 45.145 61.665 45.250 ;
        RECT 54.535 40.100 55.015 40.205 ;
        RECT 58.335 40.100 58.895 40.110 ;
        RECT 54.535 39.680 58.895 40.100 ;
        RECT 54.535 39.655 55.015 39.680 ;
        RECT 58.335 36.840 58.895 39.680 ;
        RECT 59.645 36.840 60.125 37.005 ;
        RECT 58.325 36.520 60.125 36.840 ;
        RECT 59.645 36.455 60.125 36.520 ;
        RECT 56.355 31.770 56.815 31.875 ;
        RECT 61.925 31.770 62.385 31.825 ;
        RECT 56.355 31.330 62.385 31.770 ;
        RECT 56.355 31.305 56.815 31.330 ;
        RECT 61.925 31.255 62.385 31.330 ;
        RECT 29.765 11.100 30.255 11.115 ;
        RECT 39.065 11.005 41.615 11.965 ;
        RECT 50.285 10.995 52.405 12.145 ;
        RECT 62.915 12.135 63.405 73.010 ;
        RECT 65.035 54.010 65.495 54.085 ;
        RECT 70.605 54.010 71.065 54.035 ;
        RECT 65.035 53.570 71.065 54.010 ;
        RECT 65.035 53.515 65.495 53.570 ;
        RECT 70.605 53.465 71.065 53.570 ;
        RECT 67.295 48.820 67.775 48.885 ;
        RECT 67.295 48.500 69.095 48.820 ;
        RECT 67.295 48.335 67.775 48.500 ;
        RECT 68.525 45.660 69.085 48.500 ;
        RECT 72.405 45.660 72.885 45.685 ;
        RECT 68.525 45.240 72.885 45.660 ;
        RECT 68.525 45.230 69.085 45.240 ;
        RECT 72.405 45.135 72.885 45.240 ;
        RECT 65.735 40.100 66.215 40.205 ;
        RECT 69.535 40.100 70.095 40.110 ;
        RECT 65.735 39.680 70.095 40.100 ;
        RECT 65.735 39.655 66.215 39.680 ;
        RECT 69.535 36.840 70.095 39.680 ;
        RECT 70.845 36.840 71.325 37.005 ;
        RECT 69.525 36.520 71.325 36.840 ;
        RECT 70.845 36.455 71.325 36.520 ;
        RECT 67.555 31.770 68.015 31.875 ;
        RECT 73.125 31.770 73.585 31.825 ;
        RECT 67.555 31.330 73.585 31.770 ;
        RECT 67.555 31.305 68.015 31.330 ;
        RECT 73.125 31.255 73.585 31.330 ;
        RECT 74.055 12.165 74.545 73.050 ;
        RECT 83.690 73.000 86.290 74.540 ;
        RECT 94.960 74.710 97.520 75.580 ;
        RECT 94.960 73.020 97.570 74.710 ;
        RECT 106.340 74.460 108.900 75.640 ;
        RECT 117.470 74.720 120.030 75.650 ;
        RECT 76.275 54.000 76.735 54.075 ;
        RECT 81.845 54.000 82.305 54.025 ;
        RECT 76.275 53.560 82.305 54.000 ;
        RECT 76.275 53.505 76.735 53.560 ;
        RECT 81.845 53.455 82.305 53.560 ;
        RECT 78.535 48.810 79.015 48.875 ;
        RECT 78.535 48.490 80.335 48.810 ;
        RECT 78.535 48.325 79.015 48.490 ;
        RECT 79.765 45.650 80.325 48.490 ;
        RECT 83.645 45.650 84.125 45.675 ;
        RECT 79.765 45.230 84.125 45.650 ;
        RECT 79.765 45.220 80.325 45.230 ;
        RECT 83.645 45.125 84.125 45.230 ;
        RECT 77.025 40.090 77.505 40.195 ;
        RECT 80.825 40.090 81.385 40.100 ;
        RECT 77.025 39.670 81.385 40.090 ;
        RECT 77.025 39.645 77.505 39.670 ;
        RECT 80.825 36.830 81.385 39.670 ;
        RECT 82.135 36.830 82.615 36.995 ;
        RECT 80.815 36.510 82.615 36.830 ;
        RECT 82.135 36.445 82.615 36.510 ;
        RECT 78.845 31.760 79.305 31.865 ;
        RECT 84.415 31.760 84.875 31.815 ;
        RECT 78.845 31.320 84.875 31.760 ;
        RECT 78.845 31.295 79.305 31.320 ;
        RECT 84.415 31.245 84.875 31.320 ;
        RECT 61.365 10.985 63.485 12.135 ;
        RECT 72.675 11.015 74.795 12.165 ;
        RECT 85.375 12.155 85.865 73.000 ;
        RECT 87.525 54.010 87.985 54.085 ;
        RECT 93.095 54.010 93.555 54.035 ;
        RECT 87.525 53.570 93.555 54.010 ;
        RECT 87.525 53.515 87.985 53.570 ;
        RECT 93.095 53.465 93.555 53.570 ;
        RECT 89.785 48.820 90.265 48.885 ;
        RECT 89.785 48.500 91.585 48.820 ;
        RECT 89.785 48.335 90.265 48.500 ;
        RECT 91.015 45.660 91.575 48.500 ;
        RECT 94.895 45.660 95.375 45.685 ;
        RECT 91.015 45.240 95.375 45.660 ;
        RECT 91.015 45.230 91.575 45.240 ;
        RECT 94.895 45.135 95.375 45.240 ;
        RECT 88.265 40.110 88.745 40.215 ;
        RECT 92.065 40.110 92.625 40.120 ;
        RECT 88.265 39.690 92.625 40.110 ;
        RECT 88.265 39.665 88.745 39.690 ;
        RECT 92.065 36.850 92.625 39.690 ;
        RECT 93.375 36.850 93.855 37.015 ;
        RECT 92.055 36.530 93.855 36.850 ;
        RECT 93.375 36.465 93.855 36.530 ;
        RECT 90.085 31.780 90.545 31.885 ;
        RECT 95.655 31.780 96.115 31.835 ;
        RECT 90.085 31.340 96.115 31.780 ;
        RECT 90.085 31.315 90.545 31.340 ;
        RECT 95.655 31.265 96.115 31.340 ;
        RECT 96.605 12.155 97.095 73.020 ;
        RECT 106.150 73.000 109.060 74.460 ;
        RECT 117.470 73.070 120.000 74.720 ;
        RECT 129.290 74.650 131.850 75.650 ;
        RECT 129.300 73.140 131.820 74.650 ;
        RECT 98.805 54.000 99.265 54.075 ;
        RECT 104.375 54.000 104.835 54.025 ;
        RECT 98.805 53.560 104.835 54.000 ;
        RECT 98.805 53.505 99.265 53.560 ;
        RECT 104.375 53.455 104.835 53.560 ;
        RECT 101.065 48.810 101.545 48.875 ;
        RECT 101.065 48.490 102.865 48.810 ;
        RECT 101.065 48.325 101.545 48.490 ;
        RECT 102.295 45.650 102.855 48.490 ;
        RECT 106.175 45.650 106.655 45.675 ;
        RECT 102.295 45.230 106.655 45.650 ;
        RECT 102.295 45.220 102.855 45.230 ;
        RECT 106.175 45.125 106.655 45.230 ;
        RECT 99.475 40.130 99.955 40.235 ;
        RECT 103.275 40.130 103.835 40.140 ;
        RECT 99.475 39.710 103.835 40.130 ;
        RECT 99.475 39.685 99.955 39.710 ;
        RECT 103.275 36.870 103.835 39.710 ;
        RECT 104.585 36.870 105.065 37.035 ;
        RECT 103.265 36.550 105.065 36.870 ;
        RECT 104.585 36.485 105.065 36.550 ;
        RECT 101.295 31.800 101.755 31.905 ;
        RECT 106.865 31.800 107.325 31.855 ;
        RECT 101.295 31.360 107.325 31.800 ;
        RECT 101.295 31.335 101.755 31.360 ;
        RECT 106.865 31.285 107.325 31.360 ;
        RECT 107.865 12.205 108.355 73.000 ;
        RECT 110.075 54.000 110.535 54.075 ;
        RECT 115.645 54.000 116.105 54.025 ;
        RECT 110.075 53.560 116.105 54.000 ;
        RECT 110.075 53.505 110.535 53.560 ;
        RECT 115.645 53.455 116.105 53.560 ;
        RECT 112.335 48.810 112.815 48.875 ;
        RECT 112.335 48.490 114.135 48.810 ;
        RECT 112.335 48.325 112.815 48.490 ;
        RECT 113.565 45.650 114.125 48.490 ;
        RECT 117.445 45.650 117.925 45.675 ;
        RECT 113.565 45.230 117.925 45.650 ;
        RECT 113.565 45.220 114.125 45.230 ;
        RECT 117.445 45.125 117.925 45.230 ;
        RECT 110.675 40.170 111.155 40.275 ;
        RECT 114.475 40.170 115.035 40.180 ;
        RECT 110.675 39.750 115.035 40.170 ;
        RECT 110.675 39.725 111.155 39.750 ;
        RECT 114.475 36.910 115.035 39.750 ;
        RECT 115.785 36.910 116.265 37.075 ;
        RECT 114.465 36.590 116.265 36.910 ;
        RECT 115.785 36.525 116.265 36.590 ;
        RECT 112.495 31.840 112.955 31.945 ;
        RECT 118.065 31.840 118.525 31.895 ;
        RECT 112.495 31.400 118.525 31.840 ;
        RECT 112.495 31.375 112.955 31.400 ;
        RECT 118.065 31.325 118.525 31.400 ;
        RECT 119.085 12.205 119.575 73.070 ;
        RECT 121.325 54.000 121.785 54.075 ;
        RECT 126.895 54.000 127.355 54.025 ;
        RECT 121.325 53.560 127.355 54.000 ;
        RECT 121.325 53.505 121.785 53.560 ;
        RECT 126.895 53.455 127.355 53.560 ;
        RECT 123.585 48.810 124.065 48.875 ;
        RECT 123.585 48.490 125.385 48.810 ;
        RECT 123.585 48.325 124.065 48.490 ;
        RECT 124.815 45.650 125.375 48.490 ;
        RECT 128.695 45.650 129.175 45.675 ;
        RECT 124.815 45.230 129.175 45.650 ;
        RECT 124.815 45.220 125.375 45.230 ;
        RECT 128.695 45.125 129.175 45.230 ;
        RECT 121.885 40.190 122.365 40.295 ;
        RECT 125.685 40.190 126.245 40.200 ;
        RECT 121.885 39.770 126.245 40.190 ;
        RECT 121.885 39.745 122.365 39.770 ;
        RECT 125.685 36.930 126.245 39.770 ;
        RECT 126.995 36.930 127.475 37.095 ;
        RECT 125.675 36.610 127.475 36.930 ;
        RECT 126.995 36.545 127.475 36.610 ;
        RECT 123.705 31.860 124.165 31.965 ;
        RECT 129.275 31.860 129.735 31.915 ;
        RECT 123.705 31.420 129.735 31.860 ;
        RECT 123.705 31.395 124.165 31.420 ;
        RECT 129.275 31.345 129.735 31.420 ;
        RECT 130.335 12.235 130.825 73.140 ;
        RECT 74.055 11.010 74.545 11.015 ;
        RECT 83.795 11.005 85.915 12.155 ;
        RECT 95.095 11.005 97.215 12.155 ;
        RECT 106.285 11.055 108.405 12.205 ;
        RECT 117.515 11.055 119.635 12.205 ;
        RECT 128.815 11.085 130.935 12.235 ;
        RECT 107.865 11.010 108.355 11.055 ;
        RECT 119.085 11.050 119.575 11.055 ;
        RECT 85.375 11.000 85.865 11.005 ;
        RECT 96.605 10.980 97.095 11.005 ;
        RECT 74.290 0.135 75.680 1.435 ;
        RECT 93.500 0.205 94.890 1.505 ;
        RECT 112.900 0.335 114.290 1.635 ;
        RECT 131.800 0.405 133.540 1.905 ;
        RECT 151.600 0.275 152.970 1.445 ;
      LAYER met4 ;
        RECT 30.420 225.130 30.670 225.140 ;
        RECT 30.300 224.760 30.670 225.130 ;
        RECT 30.970 224.760 33.430 225.140 ;
        RECT 33.730 224.760 36.190 225.140 ;
        RECT 36.490 224.760 38.950 225.140 ;
        RECT 39.250 224.760 41.710 225.140 ;
        RECT 42.010 224.760 44.470 225.140 ;
        RECT 44.770 224.760 47.230 225.140 ;
        RECT 47.530 224.760 49.990 225.140 ;
        RECT 50.290 224.760 52.750 225.140 ;
        RECT 53.050 224.760 55.510 225.140 ;
        RECT 55.810 224.760 58.270 225.140 ;
        RECT 58.570 224.760 61.030 225.140 ;
        RECT 61.330 224.760 63.790 225.140 ;
        RECT 64.090 224.760 66.550 225.140 ;
        RECT 66.850 224.760 69.310 225.140 ;
        RECT 69.610 224.760 72.070 225.140 ;
        RECT 72.370 224.760 74.830 225.140 ;
        RECT 75.130 224.760 77.590 225.140 ;
        RECT 77.890 224.760 80.350 225.140 ;
        RECT 80.650 224.760 83.110 225.140 ;
        RECT 83.410 224.760 85.870 225.140 ;
        RECT 86.170 224.760 88.630 225.140 ;
        RECT 88.930 224.760 91.390 225.140 ;
        RECT 91.690 224.760 94.150 225.140 ;
        RECT 94.450 224.760 96.910 225.140 ;
        RECT 97.210 224.760 99.670 225.140 ;
        RECT 99.970 224.760 102.430 225.140 ;
        RECT 102.730 224.760 105.190 225.140 ;
        RECT 105.490 224.760 107.950 225.140 ;
        RECT 108.250 224.760 110.710 225.140 ;
        RECT 111.010 224.760 113.470 225.140 ;
        RECT 113.770 224.760 116.230 225.140 ;
        RECT 116.530 224.760 118.990 225.140 ;
        RECT 119.290 224.760 121.750 225.140 ;
        RECT 122.050 224.760 124.510 225.140 ;
        RECT 124.810 224.760 127.270 225.140 ;
        RECT 127.570 224.760 130.030 225.140 ;
        RECT 130.330 224.760 132.790 225.140 ;
        RECT 133.090 224.760 133.520 225.140 ;
        RECT 30.300 224.240 133.520 224.760 ;
        RECT 135.385 224.760 135.550 225.185 ;
        RECT 135.850 224.760 136.745 225.185 ;
        RECT 30.300 219.100 31.660 224.240 ;
        RECT 135.385 223.875 136.745 224.760 ;
        RECT 138.175 224.760 138.310 225.115 ;
        RECT 138.610 224.760 139.535 225.115 ;
        RECT 138.175 223.805 139.535 224.760 ;
        RECT 143.225 224.760 143.830 225.145 ;
        RECT 144.130 224.760 144.585 225.145 ;
        RECT 143.225 223.835 144.585 224.760 ;
        RECT 6.000 218.040 31.660 219.100 ;
        RECT 30.300 217.960 31.660 218.040 ;
        RECT 10.650 108.115 12.250 214.675 ;
        RECT 24.045 108.115 25.645 214.675 ;
        RECT 34.265 174.490 34.595 174.820 ;
        RECT 32.425 157.490 32.755 157.820 ;
        RECT 32.440 120.420 32.740 157.490 ;
        RECT 34.280 140.820 34.580 174.490 ;
        RECT 34.265 140.490 34.595 140.820 ;
        RECT 32.425 120.090 32.755 120.420 ;
        RECT 37.440 108.115 39.040 214.675 ;
        RECT 50.835 108.115 52.435 214.675 ;
        RECT 59.105 157.805 59.435 157.820 ;
        RECT 58.200 157.505 59.435 157.805 ;
        RECT 58.200 128.580 58.500 157.505 ;
        RECT 59.105 157.490 59.435 157.505 ;
        RECT 58.185 128.250 58.515 128.580 ;
        RECT 64.230 108.115 65.830 214.675 ;
        RECT 71.985 171.090 72.315 171.420 ;
        RECT 72.000 140.820 72.300 171.090 ;
        RECT 73.825 159.530 74.155 159.860 ;
        RECT 73.840 153.060 74.140 159.530 ;
        RECT 73.825 152.730 74.155 153.060 ;
        RECT 71.985 140.490 72.315 140.820 ;
        RECT 77.625 108.115 79.225 214.675 ;
        RECT 83.945 182.650 84.275 182.980 ;
        RECT 83.960 180.940 84.260 182.650 ;
        RECT 83.945 180.610 84.275 180.940 ;
        RECT 83.960 176.180 84.260 180.610 ;
        RECT 83.945 175.850 84.275 176.180 ;
        RECT 91.020 108.115 92.620 214.675 ;
        RECT 95.905 198.290 96.235 198.620 ;
        RECT 95.920 161.900 96.220 198.290 ;
        RECT 95.905 161.570 96.235 161.900 ;
        RECT 104.415 108.115 106.015 214.675 ;
        RECT 118.110 97.700 120.130 99.670 ;
        RECT 121.810 97.750 123.830 99.720 ;
        RECT 118.130 93.980 120.130 97.700 ;
        RECT 121.820 96.830 123.820 97.750 ;
        RECT 121.820 94.830 139.410 96.830 ;
        RECT 118.130 91.980 135.580 93.980 ;
        RECT 133.580 77.835 135.580 91.980 ;
        RECT 133.375 76.625 136.015 77.835 ;
        RECT 137.410 77.815 139.410 94.830 ;
        RECT 137.235 76.605 139.875 77.815 ;
        RECT 3.955 71.365 4.000 73.195 ;
        RECT 6.000 71.365 6.055 73.195 ;
        RECT 3.000 68.705 3.025 70.435 ;
        RECT 15.555 68.655 16.995 71.165 ;
        RECT 74.335 1.000 75.635 1.415 ;
        RECT 74.335 0.155 74.530 1.000 ;
        RECT 75.430 0.155 75.635 1.000 ;
        RECT 93.545 1.000 94.845 1.485 ;
        RECT 93.545 0.225 93.850 1.000 ;
        RECT 94.750 0.225 94.845 1.000 ;
        RECT 112.945 1.000 114.245 1.615 ;
        RECT 112.945 0.355 113.170 1.000 ;
        RECT 114.070 0.355 114.245 1.000 ;
        RECT 131.845 1.000 133.495 1.885 ;
        RECT 131.845 0.425 132.490 1.000 ;
        RECT 133.390 0.425 133.495 1.000 ;
        RECT 151.645 1.000 152.925 1.425 ;
        RECT 151.645 0.295 151.810 1.000 ;
        RECT 152.710 0.295 152.925 1.000 ;
  END
END tt_um_08_sws
END LIBRARY

