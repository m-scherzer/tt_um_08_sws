VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_08_sws
  CLASS BLOCK ;
  FOREIGN tt_um_08_sws ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    ANTENNAGATEAREA 200.000000 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    ANTENNAGATEAREA 550.000000 ;
    ANTENNADIFFAREA 2.900000 ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    ANTENNAGATEAREA 550.000000 ;
    ANTENNADIFFAREA 2.900000 ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    ANTENNADIFFAREA 29.000000 ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    ANTENNADIFFAREA 29.000000 ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    ANTENNADIFFAREA 394.109192 ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 22.975 203.925 23.145 204.115 ;
        RECT 24.410 203.975 24.530 204.085 ;
        RECT 29.875 203.925 30.045 204.115 ;
        RECT 35.395 203.925 35.565 204.115 ;
        RECT 37.235 203.925 37.405 204.115 ;
        RECT 42.755 203.925 42.925 204.115 ;
        RECT 48.275 203.925 48.445 204.115 ;
        RECT 49.250 203.975 49.370 204.085 ;
        RECT 52.875 203.925 53.045 204.115 ;
        RECT 58.395 203.925 58.565 204.115 ;
        RECT 59.775 203.925 59.945 204.115 ;
        RECT 61.155 203.925 61.325 204.115 ;
        RECT 62.130 203.975 62.250 204.085 ;
        RECT 64.375 203.925 64.545 204.115 ;
        RECT 64.840 203.925 65.010 204.115 ;
        RECT 22.835 203.115 24.205 203.925 ;
        RECT 24.675 203.115 30.185 203.925 ;
        RECT 30.195 203.115 35.705 203.925 ;
        RECT 35.725 203.055 36.155 203.840 ;
        RECT 36.175 203.115 37.545 203.925 ;
        RECT 37.555 203.115 43.065 203.925 ;
        RECT 43.075 203.115 48.585 203.925 ;
        RECT 48.605 203.055 49.035 203.840 ;
        RECT 49.515 203.115 53.185 203.925 ;
        RECT 53.195 203.115 58.705 203.925 ;
        RECT 58.725 203.015 60.075 203.925 ;
        RECT 60.095 203.145 61.465 203.925 ;
        RECT 61.485 203.055 61.915 203.840 ;
        RECT 62.395 203.245 64.685 203.925 ;
        RECT 62.395 203.015 63.315 203.245 ;
        RECT 64.695 203.015 67.615 203.925 ;
        RECT 67.915 203.895 68.860 203.925 ;
        RECT 70.815 203.895 70.985 204.115 ;
        RECT 71.280 203.925 71.450 204.115 ;
        RECT 74.035 203.970 74.195 204.080 ;
        RECT 75.875 203.925 76.045 204.115 ;
        RECT 77.255 203.925 77.425 204.115 ;
        RECT 77.715 203.925 77.885 204.115 ;
        RECT 81.395 203.925 81.565 204.115 ;
        RECT 86.915 203.925 87.085 204.115 ;
        RECT 89.215 203.925 89.385 204.115 ;
        RECT 94.735 203.925 94.905 204.115 ;
        RECT 96.115 203.925 96.285 204.115 ;
        RECT 97.035 203.970 97.195 204.080 ;
        RECT 97.495 203.925 97.665 204.115 ;
        RECT 98.875 203.925 99.045 204.115 ;
        RECT 101.635 203.925 101.805 204.115 ;
        RECT 102.150 203.975 102.270 204.085 ;
        RECT 102.555 203.925 102.725 204.115 ;
        RECT 106.290 203.975 106.410 204.085 ;
        RECT 111.755 203.925 111.925 204.115 ;
        RECT 113.135 203.925 113.305 204.115 ;
        RECT 67.915 203.695 70.985 203.895 ;
        RECT 67.915 203.215 71.125 203.695 ;
        RECT 67.915 203.015 68.860 203.215 ;
        RECT 70.195 203.015 71.125 203.215 ;
        RECT 71.135 203.015 73.425 203.925 ;
        RECT 74.365 203.055 74.795 203.840 ;
        RECT 74.825 203.015 76.175 203.925 ;
        RECT 76.205 203.015 77.555 203.925 ;
        RECT 77.575 203.145 78.945 203.925 ;
        RECT 78.955 203.115 81.705 203.925 ;
        RECT 81.715 203.115 87.225 203.925 ;
        RECT 87.245 203.055 87.675 203.840 ;
        RECT 87.695 203.115 89.525 203.925 ;
        RECT 89.535 203.115 95.045 203.925 ;
        RECT 95.065 203.015 96.415 203.925 ;
        RECT 97.355 203.145 98.725 203.925 ;
        RECT 98.745 203.015 100.095 203.925 ;
        RECT 100.125 203.055 100.555 203.840 ;
        RECT 100.585 203.015 101.935 203.925 ;
        RECT 102.525 203.245 105.990 203.925 ;
        RECT 105.070 203.015 105.990 203.245 ;
        RECT 106.555 203.115 112.065 203.925 ;
        RECT 112.075 203.115 113.445 203.925 ;
      LAYER nwell ;
        RECT 22.640 199.895 113.640 202.725 ;
      LAYER pwell ;
        RECT 22.835 198.695 24.205 199.505 ;
        RECT 24.675 198.695 30.185 199.505 ;
        RECT 30.195 198.695 35.705 199.505 ;
        RECT 35.725 198.780 36.155 199.565 ;
        RECT 36.175 198.695 37.545 199.505 ;
        RECT 37.555 198.695 41.225 199.505 ;
        RECT 41.235 198.695 46.745 199.505 ;
        RECT 46.755 198.695 52.265 199.505 ;
        RECT 56.785 199.375 57.715 199.595 ;
        RECT 60.545 199.375 61.465 199.605 ;
        RECT 52.275 198.695 61.465 199.375 ;
        RECT 61.485 198.780 61.915 199.565 ;
        RECT 61.935 198.695 63.765 199.505 ;
        RECT 63.775 198.695 66.885 199.605 ;
        RECT 69.735 199.375 70.665 199.605 ;
        RECT 66.995 198.695 70.665 199.375 ;
        RECT 70.675 199.375 71.595 199.605 ;
        RECT 74.425 199.375 75.355 199.595 ;
        RECT 70.675 198.695 79.865 199.375 ;
        RECT 79.875 198.695 82.985 199.605 ;
        RECT 83.095 198.695 85.845 199.505 ;
        RECT 85.865 198.695 87.215 199.605 ;
        RECT 87.245 198.780 87.675 199.565 ;
        RECT 88.625 198.695 89.975 199.605 ;
        RECT 92.650 199.375 93.570 199.605 ;
        RECT 96.330 199.375 97.250 199.605 ;
        RECT 90.105 198.695 93.570 199.375 ;
        RECT 93.785 198.695 97.250 199.375 ;
        RECT 97.355 199.375 98.275 199.605 ;
        RECT 101.105 199.375 102.035 199.595 ;
        RECT 97.355 198.695 106.545 199.375 ;
        RECT 107.015 198.695 108.385 199.475 ;
        RECT 108.395 198.695 112.065 199.505 ;
        RECT 112.075 198.695 113.445 199.505 ;
        RECT 22.975 198.485 23.145 198.695 ;
        RECT 24.410 198.535 24.530 198.645 ;
        RECT 26.195 198.485 26.365 198.675 ;
        RECT 29.875 198.505 30.045 198.695 ;
        RECT 31.715 198.485 31.885 198.675 ;
        RECT 35.395 198.505 35.565 198.695 ;
        RECT 37.235 198.485 37.405 198.695 ;
        RECT 40.915 198.505 41.085 198.695 ;
        RECT 42.755 198.485 42.925 198.675 ;
        RECT 46.435 198.505 46.605 198.695 ;
        RECT 48.275 198.485 48.445 198.675 ;
        RECT 50.115 198.485 50.285 198.675 ;
        RECT 50.630 198.535 50.750 198.645 ;
        RECT 51.955 198.505 52.125 198.695 ;
        RECT 52.415 198.505 52.585 198.695 ;
        RECT 54.255 198.485 54.425 198.675 ;
        RECT 54.715 198.485 54.885 198.675 ;
        RECT 63.455 198.505 63.625 198.695 ;
        RECT 65.295 198.485 65.465 198.675 ;
        RECT 66.675 198.505 66.845 198.695 ;
        RECT 67.135 198.505 67.305 198.695 ;
        RECT 70.355 198.485 70.525 198.675 ;
        RECT 70.815 198.485 70.985 198.675 ;
        RECT 75.010 198.535 75.130 198.645 ;
        RECT 77.255 198.485 77.425 198.675 ;
        RECT 79.555 198.505 79.725 198.695 ;
        RECT 82.775 198.505 82.945 198.695 ;
        RECT 85.535 198.505 85.705 198.695 ;
        RECT 85.995 198.505 86.165 198.695 ;
        RECT 86.455 198.485 86.625 198.675 ;
        RECT 86.970 198.535 87.090 198.645 ;
        RECT 87.375 198.485 87.545 198.675 ;
        RECT 88.295 198.540 88.455 198.650 ;
        RECT 88.755 198.505 88.925 198.695 ;
        RECT 90.135 198.505 90.305 198.695 ;
        RECT 93.815 198.505 93.985 198.695 ;
        RECT 99.795 198.485 99.965 198.675 ;
        RECT 104.120 198.485 104.290 198.675 ;
        RECT 104.855 198.485 105.025 198.675 ;
        RECT 106.235 198.505 106.405 198.695 ;
        RECT 106.750 198.535 106.870 198.645 ;
        RECT 108.075 198.505 108.245 198.695 ;
        RECT 109.455 198.485 109.625 198.675 ;
        RECT 110.835 198.485 111.005 198.675 ;
        RECT 111.755 198.505 111.925 198.695 ;
        RECT 113.135 198.485 113.305 198.695 ;
        RECT 22.835 197.675 24.205 198.485 ;
        RECT 24.675 197.675 26.505 198.485 ;
        RECT 26.515 197.675 32.025 198.485 ;
        RECT 32.035 197.675 37.545 198.485 ;
        RECT 37.555 197.675 43.065 198.485 ;
        RECT 43.075 197.675 48.585 198.485 ;
        RECT 48.605 197.615 49.035 198.400 ;
        RECT 49.055 197.705 50.425 198.485 ;
        RECT 50.895 197.675 54.565 198.485 ;
        RECT 54.575 197.805 64.945 198.485 ;
        RECT 65.265 197.805 68.730 198.485 ;
        RECT 59.085 197.585 60.015 197.805 ;
        RECT 62.735 197.575 64.945 197.805 ;
        RECT 67.810 197.575 68.730 197.805 ;
        RECT 68.835 197.805 70.665 198.485 ;
        RECT 70.785 197.805 74.250 198.485 ;
        RECT 68.835 197.575 70.180 197.805 ;
        RECT 73.330 197.575 74.250 197.805 ;
        RECT 74.365 197.615 74.795 198.400 ;
        RECT 75.275 197.805 77.565 198.485 ;
        RECT 77.575 197.805 86.765 198.485 ;
        RECT 87.345 197.805 90.810 198.485 ;
        RECT 75.275 197.575 76.195 197.805 ;
        RECT 77.575 197.575 78.495 197.805 ;
        RECT 81.325 197.585 82.255 197.805 ;
        RECT 89.890 197.575 90.810 197.805 ;
        RECT 90.915 197.805 100.105 198.485 ;
        RECT 90.915 197.575 91.835 197.805 ;
        RECT 94.665 197.585 95.595 197.805 ;
        RECT 100.125 197.615 100.555 198.400 ;
        RECT 100.805 197.805 104.705 198.485 ;
        RECT 104.825 197.805 108.290 198.485 ;
        RECT 103.775 197.575 104.705 197.805 ;
        RECT 107.370 197.575 108.290 197.805 ;
        RECT 108.395 197.705 109.765 198.485 ;
        RECT 109.775 197.705 111.145 198.485 ;
        RECT 112.075 197.675 113.445 198.485 ;
      LAYER nwell ;
        RECT 22.640 194.455 113.640 197.285 ;
      LAYER pwell ;
        RECT 22.835 193.255 24.205 194.065 ;
        RECT 25.135 193.255 30.645 194.065 ;
        RECT 30.665 193.255 32.015 194.165 ;
        RECT 32.230 193.255 35.705 194.165 ;
        RECT 35.725 193.340 36.155 194.125 ;
        RECT 36.175 193.255 37.545 194.065 ;
        RECT 40.210 193.935 41.130 194.165 ;
        RECT 37.665 193.255 41.130 193.935 ;
        RECT 41.235 193.255 43.065 194.065 ;
        RECT 45.730 193.935 46.650 194.165 ;
        RECT 49.410 193.935 50.330 194.165 ;
        RECT 43.185 193.255 46.650 193.935 ;
        RECT 46.865 193.255 50.330 193.935 ;
        RECT 50.905 193.255 52.255 194.165 ;
        RECT 53.195 193.255 58.705 194.065 ;
        RECT 58.725 193.255 60.075 194.165 ;
        RECT 60.095 193.255 61.465 194.065 ;
        RECT 61.485 193.340 61.915 194.125 ;
        RECT 62.855 193.965 63.785 194.165 ;
        RECT 65.120 193.965 66.065 194.165 ;
        RECT 62.855 193.485 66.065 193.965 ;
        RECT 67.655 193.935 70.655 194.165 ;
        RECT 62.995 193.285 66.065 193.485 ;
        RECT 22.975 193.045 23.145 193.255 ;
        RECT 24.815 193.100 24.975 193.210 ;
        RECT 25.275 193.045 25.445 193.235 ;
        RECT 28.955 193.045 29.125 193.235 ;
        RECT 30.335 193.045 30.505 193.255 ;
        RECT 30.795 193.045 30.965 193.255 ;
        RECT 32.175 193.045 32.345 193.235 ;
        RECT 35.390 193.065 35.560 193.255 ;
        RECT 35.860 193.045 36.030 193.235 ;
        RECT 37.235 193.065 37.405 193.255 ;
        RECT 37.695 193.065 37.865 193.255 ;
        RECT 42.755 193.065 42.925 193.255 ;
        RECT 43.215 193.065 43.385 193.255 ;
        RECT 46.895 193.065 47.065 193.255 ;
        RECT 48.275 193.045 48.445 193.235 ;
        RECT 49.655 193.090 49.815 193.200 ;
        RECT 50.630 193.095 50.750 193.205 ;
        RECT 51.035 193.045 51.205 193.235 ;
        RECT 51.495 193.045 51.665 193.235 ;
        RECT 51.955 193.065 52.125 193.255 ;
        RECT 52.875 193.100 53.035 193.210 ;
        RECT 56.095 193.045 56.265 193.235 ;
        RECT 57.015 193.090 57.175 193.200 ;
        RECT 58.395 193.065 58.565 193.255 ;
        RECT 59.775 193.065 59.945 193.255 ;
        RECT 61.155 193.065 61.325 193.255 ;
        RECT 62.535 193.045 62.705 193.235 ;
        RECT 62.995 193.065 63.165 193.285 ;
        RECT 65.120 193.255 66.065 193.285 ;
        RECT 66.075 193.845 70.655 193.935 ;
        RECT 70.675 193.935 71.595 194.165 ;
        RECT 74.425 193.935 75.355 194.155 ;
        RECT 66.075 193.485 70.665 193.845 ;
        RECT 66.075 193.255 67.645 193.485 ;
        RECT 69.735 193.295 70.665 193.485 ;
        RECT 69.735 193.255 70.655 193.295 ;
        RECT 70.675 193.255 79.865 193.935 ;
        RECT 79.875 193.255 81.225 194.165 ;
        RECT 81.265 193.255 82.615 194.165 ;
        RECT 86.210 193.935 87.130 194.165 ;
        RECT 83.665 193.255 87.130 193.935 ;
        RECT 87.245 193.340 87.675 194.125 ;
        RECT 87.695 193.935 88.615 194.165 ;
        RECT 91.445 193.935 92.375 194.155 ;
        RECT 99.550 193.935 100.470 194.165 ;
        RECT 105.085 193.935 106.015 194.155 ;
        RECT 108.845 193.935 109.765 194.165 ;
        RECT 87.695 193.255 96.885 193.935 ;
        RECT 97.005 193.255 100.470 193.935 ;
        RECT 100.575 193.255 109.765 193.935 ;
        RECT 109.785 193.255 111.135 194.165 ;
        RECT 112.075 193.255 113.445 194.065 ;
        RECT 66.215 193.065 66.385 193.255 ;
        RECT 68.055 193.045 68.225 193.235 ;
        RECT 69.895 193.045 70.065 193.235 ;
        RECT 70.410 193.095 70.530 193.205 ;
        RECT 72.195 193.045 72.365 193.235 ;
        RECT 72.655 193.045 72.825 193.235 ;
        RECT 74.960 193.045 75.130 193.235 ;
        RECT 79.555 193.065 79.725 193.255 ;
        RECT 80.475 193.090 80.635 193.200 ;
        RECT 80.940 193.065 81.110 193.255 ;
        RECT 82.315 193.065 82.485 193.255 ;
        RECT 83.235 193.100 83.395 193.210 ;
        RECT 83.695 193.065 83.865 193.255 ;
        RECT 79.555 193.045 79.720 193.065 ;
        RECT 84.340 193.045 84.510 193.235 ;
        RECT 85.130 193.095 85.250 193.205 ;
        RECT 86.455 193.045 86.625 193.235 ;
        RECT 87.835 193.045 88.005 193.235 ;
        RECT 91.700 193.045 91.870 193.235 ;
        RECT 92.435 193.045 92.605 193.235 ;
        RECT 96.575 193.065 96.745 193.255 ;
        RECT 97.035 193.065 97.205 193.255 ;
        RECT 97.220 193.045 97.390 193.235 ;
        RECT 98.415 193.090 98.575 193.200 ;
        RECT 98.875 193.045 99.045 193.235 ;
        RECT 100.715 193.065 100.885 193.255 ;
        RECT 104.120 193.045 104.290 193.235 ;
        RECT 108.075 193.045 108.245 193.235 ;
        RECT 109.915 193.065 110.085 193.255 ;
        RECT 111.755 193.045 111.925 193.235 ;
        RECT 113.135 193.045 113.305 193.255 ;
        RECT 22.835 192.235 24.205 193.045 ;
        RECT 24.215 192.235 25.585 193.045 ;
        RECT 25.595 192.235 29.265 193.045 ;
        RECT 29.285 192.135 30.635 193.045 ;
        RECT 30.655 192.265 32.025 193.045 ;
        RECT 32.145 192.365 35.610 193.045 ;
        RECT 34.690 192.135 35.610 192.365 ;
        RECT 35.715 192.135 39.190 193.045 ;
        RECT 39.395 192.365 48.585 193.045 ;
        RECT 39.395 192.135 40.315 192.365 ;
        RECT 43.145 192.145 44.075 192.365 ;
        RECT 48.605 192.175 49.035 192.960 ;
        RECT 49.975 192.265 51.345 193.045 ;
        RECT 51.465 192.365 54.930 193.045 ;
        RECT 54.010 192.135 54.930 192.365 ;
        RECT 55.045 192.135 56.395 193.045 ;
        RECT 57.335 192.235 62.845 193.045 ;
        RECT 62.855 192.235 68.365 193.045 ;
        RECT 68.375 192.365 70.205 193.045 ;
        RECT 70.675 192.235 72.505 193.045 ;
        RECT 72.515 192.365 74.345 193.045 ;
        RECT 74.365 192.175 74.795 192.960 ;
        RECT 74.815 192.135 77.425 193.045 ;
        RECT 77.885 192.365 79.720 193.045 ;
        RECT 81.025 192.365 84.925 193.045 ;
        RECT 77.885 192.135 78.815 192.365 ;
        RECT 83.995 192.135 84.925 192.365 ;
        RECT 85.395 192.265 86.765 193.045 ;
        RECT 86.785 192.135 88.135 193.045 ;
        RECT 88.385 192.365 92.285 193.045 ;
        RECT 91.355 192.135 92.285 192.365 ;
        RECT 92.295 192.265 93.665 193.045 ;
        RECT 93.905 192.365 97.805 193.045 ;
        RECT 96.875 192.135 97.805 192.365 ;
        RECT 98.735 192.265 100.105 193.045 ;
        RECT 100.125 192.175 100.555 192.960 ;
        RECT 100.805 192.365 104.705 193.045 ;
        RECT 103.775 192.135 104.705 192.365 ;
        RECT 104.810 192.365 108.275 193.045 ;
        RECT 108.490 192.365 111.955 193.045 ;
        RECT 104.810 192.135 105.730 192.365 ;
        RECT 108.490 192.135 109.410 192.365 ;
        RECT 112.075 192.235 113.445 193.045 ;
      LAYER nwell ;
        RECT 22.640 189.015 113.640 191.845 ;
      LAYER pwell ;
        RECT 22.835 187.815 24.205 188.625 ;
        RECT 26.870 188.495 27.790 188.725 ;
        RECT 24.325 187.815 27.790 188.495 ;
        RECT 28.450 188.495 29.370 188.725 ;
        RECT 28.450 187.815 31.915 188.495 ;
        RECT 32.035 187.815 35.510 188.725 ;
        RECT 35.725 187.900 36.155 188.685 ;
        RECT 36.175 188.495 37.105 188.725 ;
        RECT 36.175 187.815 40.075 188.495 ;
        RECT 40.315 187.815 41.685 188.595 ;
        RECT 41.705 187.815 43.055 188.725 ;
        RECT 47.585 188.495 48.515 188.715 ;
        RECT 51.345 188.495 52.265 188.725 ;
        RECT 43.075 187.815 52.265 188.495 ;
        RECT 52.275 188.495 53.195 188.725 ;
        RECT 56.025 188.495 56.955 188.715 ;
        RECT 52.275 187.815 61.465 188.495 ;
        RECT 61.485 187.900 61.915 188.685 ;
        RECT 61.935 187.815 67.445 188.625 ;
        RECT 67.695 188.045 70.450 188.725 ;
        RECT 70.890 188.045 73.645 188.725 ;
        RECT 67.695 187.815 69.965 188.045 ;
        RECT 71.375 187.815 73.645 188.045 ;
        RECT 73.895 187.815 76.505 188.725 ;
        RECT 77.945 188.615 78.865 188.725 ;
        RECT 77.945 188.495 80.280 188.615 ;
        RECT 84.945 188.495 85.865 188.715 ;
        RECT 77.945 187.815 87.225 188.495 ;
        RECT 87.245 187.900 87.675 188.685 ;
        RECT 90.350 188.495 91.270 188.725 ;
        RECT 95.035 188.495 95.965 188.725 ;
        RECT 100.095 188.495 101.025 188.725 ;
        RECT 87.805 187.815 91.270 188.495 ;
        RECT 92.065 187.815 95.965 188.495 ;
        RECT 97.125 187.815 101.025 188.495 ;
        RECT 101.035 188.495 101.955 188.725 ;
        RECT 104.785 188.495 105.715 188.715 ;
        RECT 101.035 187.815 110.225 188.495 ;
        RECT 110.235 187.815 111.605 188.595 ;
        RECT 112.075 187.815 113.445 188.625 ;
        RECT 22.975 187.605 23.145 187.815 ;
        RECT 24.355 187.765 24.525 187.815 ;
        RECT 24.355 187.655 24.530 187.765 ;
        RECT 24.355 187.625 24.525 187.655 ;
        RECT 26.195 187.605 26.365 187.795 ;
        RECT 28.090 187.655 28.210 187.765 ;
        RECT 31.715 187.625 31.885 187.815 ;
        RECT 32.180 187.625 32.350 187.815 ;
        RECT 35.395 187.605 35.565 187.795 ;
        RECT 36.590 187.625 36.760 187.815 ;
        RECT 40.455 187.625 40.625 187.815 ;
        RECT 41.835 187.625 42.005 187.815 ;
        RECT 43.215 187.625 43.385 187.815 ;
        RECT 44.595 187.605 44.765 187.795 ;
        RECT 48.270 187.605 48.440 187.795 ;
        RECT 49.655 187.650 49.815 187.760 ;
        RECT 50.115 187.605 50.285 187.795 ;
        RECT 51.770 187.605 51.940 187.795 ;
        RECT 55.910 187.605 56.080 187.795 ;
        RECT 60.695 187.605 60.865 187.795 ;
        RECT 61.155 187.625 61.325 187.815 ;
        RECT 61.615 187.650 61.775 187.760 ;
        RECT 62.995 187.605 63.165 187.795 ;
        RECT 63.510 187.655 63.630 187.765 ;
        RECT 63.915 187.625 64.085 187.795 ;
        RECT 64.015 187.605 64.085 187.625 ;
        RECT 67.135 187.605 67.305 187.815 ;
        RECT 67.695 187.795 67.765 187.815 ;
        RECT 73.575 187.795 73.645 187.815 ;
        RECT 67.595 187.625 67.765 187.795 ;
        RECT 71.735 187.605 71.905 187.795 ;
        RECT 73.575 187.625 73.745 187.795 ;
        RECT 74.040 187.625 74.210 187.815 ;
        RECT 75.415 187.650 75.575 187.760 ;
        RECT 75.875 187.605 76.045 187.795 ;
        RECT 77.255 187.660 77.415 187.770 ;
        RECT 86.455 187.605 86.625 187.795 ;
        RECT 86.915 187.605 87.085 187.815 ;
        RECT 87.835 187.625 88.005 187.815 ;
        RECT 91.570 187.655 91.690 187.765 ;
        RECT 95.380 187.625 95.550 187.815 ;
        RECT 96.575 187.660 96.735 187.770 ;
        RECT 97.035 187.605 97.205 187.795 ;
        RECT 97.495 187.605 97.665 187.795 ;
        RECT 98.875 187.605 99.045 187.795 ;
        RECT 100.440 187.625 100.610 187.815 ;
        RECT 101.175 187.650 101.335 187.760 ;
        RECT 109.915 187.625 110.085 187.815 ;
        RECT 110.375 187.605 110.545 187.795 ;
        RECT 110.835 187.605 111.005 187.795 ;
        RECT 111.295 187.625 111.465 187.815 ;
        RECT 111.810 187.655 111.930 187.765 ;
        RECT 113.135 187.605 113.305 187.815 ;
        RECT 22.835 186.795 24.205 187.605 ;
        RECT 24.675 186.795 26.505 187.605 ;
        RECT 26.515 186.925 35.705 187.605 ;
        RECT 35.715 186.925 44.905 187.605 ;
        RECT 26.515 186.695 27.435 186.925 ;
        RECT 30.265 186.705 31.195 186.925 ;
        RECT 35.715 186.695 36.635 186.925 ;
        RECT 39.465 186.705 40.395 186.925 ;
        RECT 45.110 186.695 48.585 187.605 ;
        RECT 48.605 186.735 49.035 187.520 ;
        RECT 49.975 186.825 51.345 187.605 ;
        RECT 51.355 186.925 55.255 187.605 ;
        RECT 55.495 186.925 59.395 187.605 ;
        RECT 51.355 186.695 52.285 186.925 ;
        RECT 55.495 186.695 56.425 186.925 ;
        RECT 59.645 186.695 60.995 187.605 ;
        RECT 61.935 186.825 63.305 187.605 ;
        RECT 64.015 187.375 66.285 187.605 ;
        RECT 66.995 187.375 68.565 187.605 ;
        RECT 70.655 187.565 71.575 187.605 ;
        RECT 70.655 187.375 71.585 187.565 ;
        RECT 64.015 186.695 66.770 187.375 ;
        RECT 66.995 187.015 71.585 187.375 ;
        RECT 66.995 186.925 71.575 187.015 ;
        RECT 71.595 186.925 74.335 187.605 ;
        RECT 68.575 186.695 71.575 186.925 ;
        RECT 74.365 186.735 74.795 187.520 ;
        RECT 75.745 186.695 77.095 187.605 ;
        RECT 77.485 186.925 86.765 187.605 ;
        RECT 77.485 186.805 79.820 186.925 ;
        RECT 77.485 186.695 78.405 186.805 ;
        RECT 84.485 186.705 85.405 186.925 ;
        RECT 86.785 186.695 88.135 187.605 ;
        RECT 88.155 186.925 97.345 187.605 ;
        RECT 88.155 186.695 89.075 186.925 ;
        RECT 91.905 186.705 92.835 186.925 ;
        RECT 97.365 186.695 98.715 187.605 ;
        RECT 98.745 186.695 100.095 187.605 ;
        RECT 100.125 186.735 100.555 187.520 ;
        RECT 101.495 186.925 110.685 187.605 ;
        RECT 101.495 186.695 102.415 186.925 ;
        RECT 105.245 186.705 106.175 186.925 ;
        RECT 110.705 186.695 112.055 187.605 ;
        RECT 112.075 186.795 113.445 187.605 ;
      LAYER nwell ;
        RECT 22.640 183.575 113.640 186.405 ;
      LAYER pwell ;
        RECT 22.835 182.375 24.205 183.185 ;
        RECT 25.145 182.375 26.495 183.285 ;
        RECT 26.515 183.055 27.435 183.285 ;
        RECT 30.265 183.055 31.195 183.275 ;
        RECT 26.515 182.375 35.705 183.055 ;
        RECT 35.725 182.460 36.155 183.245 ;
        RECT 36.830 182.375 40.305 183.285 ;
        RECT 40.315 183.055 41.245 183.285 ;
        RECT 40.315 182.375 44.215 183.055 ;
        RECT 44.915 182.375 46.745 183.185 ;
        RECT 46.755 183.055 47.685 183.285 ;
        RECT 46.755 182.375 50.655 183.055 ;
        RECT 50.895 182.375 52.265 183.185 ;
        RECT 52.275 183.055 53.195 183.285 ;
        RECT 56.025 183.055 56.955 183.275 ;
        RECT 52.275 182.375 61.465 183.055 ;
        RECT 61.485 182.460 61.915 183.245 ;
        RECT 61.945 182.375 64.685 183.055 ;
        RECT 64.705 182.375 66.055 183.285 ;
        RECT 66.075 183.055 67.420 183.285 ;
        RECT 67.915 183.055 69.260 183.285 ;
        RECT 66.075 182.375 67.905 183.055 ;
        RECT 67.915 182.375 69.745 183.055 ;
        RECT 69.995 182.605 72.750 183.285 ;
        RECT 69.995 182.375 72.265 182.605 ;
        RECT 73.435 182.375 76.155 183.285 ;
        RECT 79.395 183.055 80.325 183.285 ;
        RECT 83.535 183.055 84.465 183.285 ;
        RECT 76.425 182.375 80.325 183.055 ;
        RECT 80.565 182.375 84.465 183.055 ;
        RECT 84.475 182.375 85.845 183.155 ;
        RECT 85.855 182.375 87.225 183.155 ;
        RECT 87.245 182.460 87.675 183.245 ;
        RECT 87.695 182.375 91.170 183.285 ;
        RECT 91.570 182.375 95.045 183.285 ;
        RECT 97.710 183.055 98.630 183.285 ;
        RECT 95.165 182.375 98.630 183.055 ;
        RECT 99.195 182.375 100.565 183.155 ;
        RECT 103.775 183.055 104.705 183.285 ;
        RECT 100.805 182.375 104.705 183.055 ;
        RECT 104.715 182.375 108.190 183.285 ;
        RECT 108.395 182.375 111.870 183.285 ;
        RECT 112.075 182.375 113.445 183.185 ;
        RECT 22.975 182.165 23.145 182.375 ;
        RECT 24.815 182.210 24.975 182.330 ;
        RECT 25.275 182.165 25.445 182.355 ;
        RECT 26.195 182.185 26.365 182.375 ;
        RECT 26.930 182.165 27.100 182.355 ;
        RECT 30.795 182.165 30.965 182.355 ;
        RECT 35.395 182.185 35.565 182.375 ;
        RECT 36.370 182.215 36.490 182.325 ;
        RECT 39.990 182.185 40.160 182.375 ;
        RECT 40.730 182.185 40.900 182.375 ;
        RECT 44.590 182.325 44.760 182.355 ;
        RECT 40.915 182.210 41.075 182.320 ;
        RECT 44.590 182.215 44.770 182.325 ;
        RECT 44.590 182.165 44.760 182.215 ;
        RECT 45.055 182.165 45.225 182.355 ;
        RECT 46.435 182.185 46.605 182.375 ;
        RECT 47.170 182.185 47.340 182.375 ;
        RECT 49.655 182.210 49.815 182.320 ;
        RECT 50.115 182.165 50.285 182.355 ;
        RECT 51.955 182.185 52.125 182.375 ;
        RECT 54.710 182.165 54.880 182.355 ;
        RECT 58.580 182.165 58.750 182.355 ;
        RECT 61.155 182.185 61.325 182.375 ;
        RECT 64.375 182.185 64.545 182.375 ;
        RECT 64.835 182.185 65.005 182.375 ;
        RECT 67.595 182.185 67.765 182.375 ;
        RECT 68.055 182.165 68.225 182.355 ;
        RECT 68.570 182.215 68.690 182.325 ;
        RECT 68.975 182.165 69.145 182.355 ;
        RECT 69.435 182.185 69.605 182.375 ;
        RECT 69.995 182.355 70.065 182.375 ;
        RECT 69.895 182.185 70.065 182.355 ;
        RECT 73.170 182.215 73.290 182.325 ;
        RECT 73.575 182.185 73.745 182.375 ;
        RECT 74.030 182.165 74.200 182.355 ;
        RECT 74.955 182.165 75.125 182.355 ;
        RECT 79.740 182.185 79.910 182.375 ;
        RECT 83.880 182.185 84.050 182.375 ;
        RECT 84.615 182.185 84.785 182.375 ;
        RECT 86.915 182.185 87.085 182.375 ;
        RECT 87.375 182.165 87.545 182.355 ;
        RECT 87.840 182.185 88.010 182.375 ;
        RECT 91.510 182.165 91.680 182.355 ;
        RECT 92.030 182.215 92.150 182.325 ;
        RECT 92.435 182.165 92.605 182.355 ;
        RECT 94.730 182.185 94.900 182.375 ;
        RECT 95.195 182.185 95.365 182.375 ;
        RECT 98.930 182.215 99.050 182.325 ;
        RECT 99.520 182.165 99.690 182.355 ;
        RECT 100.255 182.185 100.425 182.375 ;
        RECT 103.935 182.165 104.105 182.355 ;
        RECT 104.120 182.185 104.290 182.375 ;
        RECT 104.400 182.165 104.570 182.355 ;
        RECT 104.860 182.185 105.030 182.375 ;
        RECT 108.075 182.165 108.245 182.355 ;
        RECT 108.540 182.185 108.710 182.375 ;
        RECT 111.810 182.215 111.930 182.325 ;
        RECT 113.135 182.165 113.305 182.375 ;
        RECT 22.835 181.355 24.205 182.165 ;
        RECT 25.135 181.385 26.505 182.165 ;
        RECT 26.515 181.485 30.415 182.165 ;
        RECT 30.655 181.485 39.935 182.165 ;
        RECT 26.515 181.255 27.445 181.485 ;
        RECT 32.015 181.265 32.935 181.485 ;
        RECT 37.600 181.365 39.935 181.485 ;
        RECT 39.015 181.255 39.935 181.365 ;
        RECT 41.430 181.255 44.905 182.165 ;
        RECT 45.025 181.485 48.490 182.165 ;
        RECT 47.570 181.255 48.490 181.485 ;
        RECT 48.605 181.295 49.035 182.080 ;
        RECT 49.975 181.385 51.345 182.165 ;
        RECT 51.550 181.255 55.025 182.165 ;
        RECT 55.265 181.485 59.165 182.165 ;
        RECT 58.235 181.255 59.165 181.485 ;
        RECT 59.175 181.485 68.365 182.165 ;
        RECT 68.835 181.485 70.665 182.165 ;
        RECT 59.175 181.255 60.095 181.485 ;
        RECT 62.925 181.265 63.855 181.485 ;
        RECT 69.320 181.255 70.665 181.485 ;
        RECT 70.870 181.255 74.345 182.165 ;
        RECT 74.365 181.295 74.795 182.080 ;
        RECT 74.925 181.485 78.390 182.165 ;
        RECT 77.470 181.255 78.390 181.485 ;
        RECT 78.495 181.485 87.685 182.165 ;
        RECT 78.495 181.255 79.415 181.485 ;
        RECT 82.245 181.265 83.175 181.485 ;
        RECT 88.350 181.255 91.825 182.165 ;
        RECT 92.405 181.485 95.870 182.165 ;
        RECT 96.205 181.485 100.105 182.165 ;
        RECT 94.950 181.255 95.870 181.485 ;
        RECT 99.175 181.255 100.105 181.485 ;
        RECT 100.125 181.295 100.555 182.080 ;
        RECT 100.670 181.485 104.135 182.165 ;
        RECT 100.670 181.255 101.590 181.485 ;
        RECT 104.255 181.255 107.730 182.165 ;
        RECT 108.045 181.485 111.510 182.165 ;
        RECT 110.590 181.255 111.510 181.485 ;
        RECT 112.075 181.355 113.445 182.165 ;
      LAYER nwell ;
        RECT 22.640 178.135 113.640 180.965 ;
      LAYER pwell ;
        RECT 22.835 176.935 24.205 177.745 ;
        RECT 26.870 177.615 27.790 177.845 ;
        RECT 24.325 176.935 27.790 177.615 ;
        RECT 28.090 176.935 31.565 177.845 ;
        RECT 31.575 177.615 32.505 177.845 ;
        RECT 31.575 176.935 35.475 177.615 ;
        RECT 35.725 177.020 36.155 177.805 ;
        RECT 39.290 177.615 40.210 177.845 ;
        RECT 43.515 177.615 44.445 177.845 ;
        RECT 36.745 176.935 40.210 177.615 ;
        RECT 40.545 176.935 44.445 177.615 ;
        RECT 44.455 177.615 45.375 177.845 ;
        RECT 48.205 177.615 49.135 177.835 ;
        RECT 56.310 177.615 57.230 177.845 ;
        RECT 60.535 177.615 61.465 177.845 ;
        RECT 44.455 176.935 53.645 177.615 ;
        RECT 53.765 176.935 57.230 177.615 ;
        RECT 57.565 176.935 61.465 177.615 ;
        RECT 61.485 177.020 61.915 177.805 ;
        RECT 61.945 176.935 63.295 177.845 ;
        RECT 63.775 176.935 65.145 177.715 ;
        RECT 65.155 176.935 66.525 177.745 ;
        RECT 66.535 177.615 67.880 177.845 ;
        RECT 68.375 177.615 69.720 177.845 ;
        RECT 66.535 176.935 68.365 177.615 ;
        RECT 68.375 176.935 70.205 177.615 ;
        RECT 70.215 176.935 73.690 177.845 ;
        RECT 73.895 176.935 77.370 177.845 ;
        RECT 77.575 176.935 81.050 177.845 ;
        RECT 83.910 177.615 84.830 177.845 ;
        RECT 81.365 176.935 84.830 177.615 ;
        RECT 84.945 176.935 86.295 177.845 ;
        RECT 87.245 177.020 87.675 177.805 ;
        RECT 87.705 176.935 89.055 177.845 ;
        RECT 92.650 177.615 93.570 177.845 ;
        RECT 90.105 176.935 93.570 177.615 ;
        RECT 93.675 176.935 95.045 177.715 ;
        RECT 95.515 177.615 96.445 177.845 ;
        RECT 95.515 176.935 99.415 177.615 ;
        RECT 100.115 176.935 101.485 177.715 ;
        RECT 101.505 176.935 102.855 177.845 ;
        RECT 102.875 177.615 103.795 177.845 ;
        RECT 106.625 177.615 107.555 177.835 ;
        RECT 102.875 176.935 112.065 177.615 ;
        RECT 112.075 176.935 113.445 177.745 ;
        RECT 22.975 176.725 23.145 176.935 ;
        RECT 24.355 176.885 24.525 176.935 ;
        RECT 24.355 176.775 24.530 176.885 ;
        RECT 24.355 176.745 24.525 176.775 ;
        RECT 26.195 176.725 26.365 176.915 ;
        RECT 26.655 176.725 26.825 176.915 ;
        RECT 28.035 176.725 28.205 176.915 ;
        RECT 29.420 176.725 29.590 176.915 ;
        RECT 31.250 176.745 31.420 176.935 ;
        RECT 31.990 176.745 32.160 176.935 ;
        RECT 36.370 176.775 36.490 176.885 ;
        RECT 36.775 176.745 36.945 176.935 ;
        RECT 41.835 176.725 42.005 176.915 ;
        RECT 43.215 176.725 43.385 176.915 ;
        RECT 43.860 176.745 44.030 176.935 ;
        RECT 44.595 176.725 44.765 176.915 ;
        RECT 48.270 176.725 48.440 176.915 ;
        RECT 50.115 176.725 50.285 176.915 ;
        RECT 50.575 176.725 50.745 176.915 ;
        RECT 53.335 176.745 53.505 176.935 ;
        RECT 53.795 176.745 53.965 176.935 ;
        RECT 55.635 176.745 55.805 176.915 ;
        RECT 55.635 176.725 55.780 176.745 ;
        RECT 57.475 176.725 57.645 176.915 ;
        RECT 57.940 176.725 58.110 176.915 ;
        RECT 60.880 176.745 61.050 176.935 ;
        RECT 61.615 176.725 61.785 176.915 ;
        RECT 62.995 176.745 63.165 176.935 ;
        RECT 63.510 176.775 63.630 176.885 ;
        RECT 63.915 176.745 64.085 176.935 ;
        RECT 66.215 176.745 66.385 176.935 ;
        RECT 67.595 176.725 67.765 176.915 ;
        RECT 68.055 176.745 68.225 176.935 ;
        RECT 69.435 176.725 69.605 176.915 ;
        RECT 69.895 176.725 70.065 176.935 ;
        RECT 70.360 176.745 70.530 176.935 ;
        RECT 74.040 176.915 74.210 176.935 ;
        RECT 74.035 176.745 74.210 176.915 ;
        RECT 74.035 176.725 74.205 176.745 ;
        RECT 75.875 176.725 76.045 176.915 ;
        RECT 77.255 176.725 77.425 176.915 ;
        RECT 77.720 176.745 77.890 176.935 ;
        RECT 78.635 176.725 78.805 176.915 ;
        RECT 80.015 176.725 80.185 176.915 ;
        RECT 80.475 176.725 80.645 176.915 ;
        RECT 81.395 176.745 81.565 176.935 ;
        RECT 85.995 176.745 86.165 176.935 ;
        RECT 86.915 176.780 87.075 176.890 ;
        RECT 87.835 176.745 88.005 176.935 ;
        RECT 89.675 176.780 89.835 176.890 ;
        RECT 90.135 176.745 90.305 176.935 ;
        RECT 93.815 176.745 93.985 176.935 ;
        RECT 95.250 176.775 95.370 176.885 ;
        RECT 95.930 176.745 96.100 176.935 ;
        RECT 98.415 176.725 98.585 176.915 ;
        RECT 99.795 176.885 99.965 176.915 ;
        RECT 99.795 176.775 99.970 176.885 ;
        RECT 99.795 176.725 99.965 176.775 ;
        RECT 100.255 176.745 100.425 176.935 ;
        RECT 101.175 176.770 101.335 176.880 ;
        RECT 101.635 176.725 101.805 176.935 ;
        RECT 103.015 176.725 103.185 176.915 ;
        RECT 111.755 176.745 111.925 176.935 ;
        RECT 113.135 176.725 113.305 176.935 ;
        RECT 22.835 175.915 24.205 176.725 ;
        RECT 24.675 175.915 26.505 176.725 ;
        RECT 26.515 175.945 27.885 176.725 ;
        RECT 27.905 175.815 29.255 176.725 ;
        RECT 29.275 175.815 32.750 176.725 ;
        RECT 32.955 176.045 42.145 176.725 ;
        RECT 32.955 175.815 33.875 176.045 ;
        RECT 36.705 175.825 37.635 176.045 ;
        RECT 42.155 175.945 43.525 176.725 ;
        RECT 43.545 175.815 44.895 176.725 ;
        RECT 45.110 175.815 48.585 176.725 ;
        RECT 48.605 175.855 49.035 176.640 ;
        RECT 49.055 175.945 50.425 176.725 ;
        RECT 50.445 175.815 51.795 176.725 ;
        RECT 51.910 175.815 55.780 176.725 ;
        RECT 55.955 175.915 57.785 176.725 ;
        RECT 57.795 175.815 61.270 176.725 ;
        RECT 61.585 176.045 65.050 176.725 ;
        RECT 64.130 175.815 65.050 176.045 ;
        RECT 65.155 175.915 67.905 176.725 ;
        RECT 67.915 176.045 69.745 176.725 ;
        RECT 67.915 175.815 69.260 176.045 ;
        RECT 69.755 175.815 72.475 176.725 ;
        RECT 72.515 175.915 74.345 176.725 ;
        RECT 74.365 175.855 74.795 176.640 ;
        RECT 74.815 175.915 76.185 176.725 ;
        RECT 76.195 175.945 77.565 176.725 ;
        RECT 77.585 175.815 78.935 176.725 ;
        RECT 78.965 175.815 80.315 176.725 ;
        RECT 80.335 176.045 89.440 176.725 ;
        RECT 89.535 176.045 98.725 176.725 ;
        RECT 89.535 175.815 90.455 176.045 ;
        RECT 93.285 175.825 94.215 176.045 ;
        RECT 98.735 175.945 100.105 176.725 ;
        RECT 100.125 175.855 100.555 176.640 ;
        RECT 101.495 175.945 102.865 176.725 ;
        RECT 102.875 176.045 112.065 176.725 ;
        RECT 107.385 175.825 108.315 176.045 ;
        RECT 111.145 175.815 112.065 176.045 ;
        RECT 112.075 175.915 113.445 176.725 ;
      LAYER nwell ;
        RECT 22.640 172.695 113.640 175.525 ;
      LAYER pwell ;
        RECT 22.835 171.495 24.205 172.305 ;
        RECT 24.225 171.495 25.575 172.405 ;
        RECT 25.595 171.495 26.965 172.275 ;
        RECT 26.985 171.495 28.335 172.405 ;
        RECT 31.010 172.175 31.930 172.405 ;
        RECT 28.465 171.495 31.930 172.175 ;
        RECT 32.230 171.495 35.705 172.405 ;
        RECT 35.725 171.580 36.155 172.365 ;
        RECT 36.260 171.495 45.365 172.175 ;
        RECT 45.385 171.495 46.735 172.405 ;
        RECT 46.755 171.495 55.860 172.175 ;
        RECT 56.415 171.495 60.085 172.305 ;
        RECT 60.105 171.495 61.455 172.405 ;
        RECT 61.485 171.580 61.915 172.365 ;
        RECT 61.935 172.175 63.280 172.405 ;
        RECT 66.905 172.295 67.825 172.405 ;
        RECT 66.905 172.175 69.240 172.295 ;
        RECT 73.905 172.175 74.825 172.395 ;
        RECT 61.935 171.495 63.765 172.175 ;
        RECT 63.785 171.495 66.525 172.175 ;
        RECT 66.905 171.495 76.185 172.175 ;
        RECT 76.215 171.495 87.225 172.405 ;
        RECT 87.245 171.580 87.675 172.365 ;
        RECT 87.705 171.495 89.055 172.405 ;
        RECT 89.085 171.495 90.435 172.405 ;
        RECT 90.915 172.175 91.835 172.405 ;
        RECT 94.665 172.175 95.595 172.395 ;
        RECT 100.115 172.175 101.035 172.405 ;
        RECT 103.865 172.175 104.795 172.395 ;
        RECT 90.915 171.495 100.105 172.175 ;
        RECT 100.115 171.495 109.305 172.175 ;
        RECT 109.455 171.495 112.065 172.405 ;
        RECT 112.075 171.495 113.445 172.305 ;
        RECT 22.975 171.285 23.145 171.495 ;
        RECT 24.815 171.330 24.975 171.440 ;
        RECT 25.275 171.305 25.445 171.495 ;
        RECT 25.735 171.305 25.905 171.495 ;
        RECT 27.115 171.305 27.285 171.495 ;
        RECT 28.495 171.305 28.665 171.495 ;
        RECT 34.475 171.285 34.645 171.475 ;
        RECT 35.390 171.305 35.560 171.495 ;
        RECT 39.070 171.285 39.240 171.475 ;
        RECT 45.055 171.305 45.225 171.495 ;
        RECT 46.435 171.305 46.605 171.495 ;
        RECT 46.895 171.305 47.065 171.495 ;
        RECT 48.275 171.285 48.445 171.475 ;
        RECT 56.150 171.335 56.270 171.445 ;
        RECT 57.935 171.285 58.105 171.475 ;
        RECT 58.855 171.330 59.015 171.440 ;
        RECT 59.315 171.285 59.485 171.475 ;
        RECT 59.775 171.305 59.945 171.495 ;
        RECT 60.235 171.305 60.405 171.495 ;
        RECT 62.995 171.285 63.165 171.475 ;
        RECT 63.455 171.305 63.625 171.495 ;
        RECT 65.750 171.285 65.920 171.475 ;
        RECT 66.215 171.305 66.385 171.495 ;
        RECT 66.675 171.330 66.835 171.440 ;
        RECT 69.430 171.285 69.600 171.475 ;
        RECT 69.950 171.335 70.070 171.445 ;
        RECT 73.760 171.285 73.930 171.475 ;
        RECT 75.875 171.305 76.045 171.495 ;
        RECT 84.155 171.285 84.325 171.475 ;
        RECT 84.670 171.335 84.790 171.445 ;
        RECT 86.910 171.305 87.080 171.495 ;
        RECT 87.835 171.305 88.005 171.495 ;
        RECT 89.215 171.305 89.385 171.495 ;
        RECT 90.650 171.335 90.770 171.445 ;
        RECT 93.815 171.285 93.985 171.475 ;
        RECT 97.680 171.285 97.850 171.475 ;
        RECT 99.795 171.285 99.965 171.495 ;
        RECT 100.990 171.285 101.160 171.475 ;
        RECT 108.075 171.285 108.245 171.475 ;
        RECT 108.995 171.305 109.165 171.495 ;
        RECT 111.295 171.285 111.465 171.475 ;
        RECT 111.750 171.445 111.920 171.495 ;
        RECT 111.750 171.335 111.930 171.445 ;
        RECT 111.750 171.305 111.920 171.335 ;
        RECT 113.135 171.285 113.305 171.495 ;
        RECT 22.835 170.475 24.205 171.285 ;
        RECT 25.505 170.605 34.785 171.285 ;
        RECT 25.505 170.485 27.840 170.605 ;
        RECT 25.505 170.375 26.425 170.485 ;
        RECT 32.505 170.385 33.425 170.605 ;
        RECT 35.910 170.375 39.385 171.285 ;
        RECT 39.395 170.605 48.585 171.285 ;
        RECT 39.395 170.375 40.315 170.605 ;
        RECT 43.145 170.385 44.075 170.605 ;
        RECT 48.605 170.415 49.035 171.200 ;
        RECT 49.055 170.605 58.245 171.285 ;
        RECT 49.055 170.375 49.975 170.605 ;
        RECT 52.805 170.385 53.735 170.605 ;
        RECT 59.175 170.505 60.545 171.285 ;
        RECT 60.565 170.605 63.305 171.285 ;
        RECT 63.455 170.375 66.065 171.285 ;
        RECT 67.135 170.375 69.745 171.285 ;
        RECT 70.445 170.605 74.345 171.285 ;
        RECT 73.415 170.375 74.345 170.605 ;
        RECT 74.365 170.415 74.795 171.200 ;
        RECT 75.185 170.605 84.465 171.285 ;
        RECT 85.020 170.605 94.125 171.285 ;
        RECT 94.365 170.605 98.265 171.285 ;
        RECT 98.275 170.605 100.105 171.285 ;
        RECT 75.185 170.485 77.520 170.605 ;
        RECT 75.185 170.375 76.105 170.485 ;
        RECT 82.185 170.385 83.105 170.605 ;
        RECT 97.335 170.375 98.265 170.605 ;
        RECT 100.125 170.415 100.555 171.200 ;
        RECT 100.575 170.605 104.475 171.285 ;
        RECT 104.810 170.605 108.275 171.285 ;
        RECT 100.575 170.375 101.505 170.605 ;
        RECT 104.810 170.375 105.730 170.605 ;
        RECT 108.395 170.375 111.555 171.285 ;
        RECT 112.075 170.475 113.445 171.285 ;
      LAYER nwell ;
        RECT 22.640 167.255 113.640 170.085 ;
      LAYER pwell ;
        RECT 22.835 166.055 24.205 166.865 ;
        RECT 24.215 166.735 25.145 166.965 ;
        RECT 31.555 166.735 32.485 166.965 ;
        RECT 24.215 166.055 28.115 166.735 ;
        RECT 28.585 166.055 32.485 166.735 ;
        RECT 32.875 166.055 35.300 166.735 ;
        RECT 35.725 166.140 36.155 166.925 ;
        RECT 39.375 166.735 40.305 166.965 ;
        RECT 36.405 166.055 40.305 166.735 ;
        RECT 40.325 166.055 41.675 166.965 ;
        RECT 44.350 166.735 45.270 166.965 ;
        RECT 48.575 166.735 49.505 166.965 ;
        RECT 41.805 166.055 45.270 166.735 ;
        RECT 45.605 166.055 49.505 166.735 ;
        RECT 49.515 166.055 50.885 166.835 ;
        RECT 50.905 166.055 52.255 166.965 ;
        RECT 52.275 166.735 53.195 166.965 ;
        RECT 56.025 166.735 56.955 166.955 ;
        RECT 52.275 166.055 61.465 166.735 ;
        RECT 61.485 166.140 61.915 166.925 ;
        RECT 62.855 166.735 64.200 166.965 ;
        RECT 62.855 166.055 64.685 166.735 ;
        RECT 64.835 166.055 67.445 166.965 ;
        RECT 67.455 166.735 68.800 166.965 ;
        RECT 72.540 166.735 73.885 166.965 ;
        RECT 67.455 166.055 69.285 166.735 ;
        RECT 69.295 166.055 72.035 166.735 ;
        RECT 72.055 166.055 73.885 166.735 ;
        RECT 74.355 166.735 75.285 166.965 ;
        RECT 82.155 166.735 83.085 166.965 ;
        RECT 86.295 166.735 87.225 166.965 ;
        RECT 74.355 166.055 78.255 166.735 ;
        RECT 79.185 166.055 83.085 166.735 ;
        RECT 83.325 166.055 87.225 166.735 ;
        RECT 87.245 166.140 87.675 166.925 ;
        RECT 88.065 166.855 88.985 166.965 ;
        RECT 88.065 166.735 90.400 166.855 ;
        RECT 95.065 166.735 95.985 166.955 ;
        RECT 100.470 166.735 101.390 166.965 ;
        RECT 104.695 166.735 105.625 166.965 ;
        RECT 88.065 166.055 97.345 166.735 ;
        RECT 97.925 166.055 101.390 166.735 ;
        RECT 101.725 166.055 105.625 166.735 ;
        RECT 105.730 166.735 106.650 166.965 ;
        RECT 105.730 166.055 109.195 166.735 ;
        RECT 109.455 166.055 112.065 166.965 ;
        RECT 112.075 166.055 113.445 166.865 ;
        RECT 22.975 165.845 23.145 166.055 ;
        RECT 24.630 165.865 24.800 166.055 ;
        RECT 31.900 165.865 32.070 166.055 ;
        RECT 33.555 165.845 33.725 166.035 ;
        RECT 34.015 165.845 34.185 166.035 ;
        RECT 35.395 165.865 35.565 166.035 ;
        RECT 37.695 165.845 37.865 166.035 ;
        RECT 39.720 165.865 39.890 166.055 ;
        RECT 40.455 165.865 40.625 166.055 ;
        RECT 41.375 165.845 41.545 166.035 ;
        RECT 41.835 165.865 42.005 166.055 ;
        RECT 45.055 165.845 45.225 166.035 ;
        RECT 48.920 165.865 49.090 166.055 ;
        RECT 49.250 165.895 49.370 166.005 ;
        RECT 49.655 165.865 49.825 166.055 ;
        RECT 51.035 165.845 51.205 166.055 ;
        RECT 51.770 165.845 51.940 166.035 ;
        RECT 59.040 165.845 59.210 166.035 ;
        RECT 61.155 165.865 61.325 166.055 ;
        RECT 62.535 165.900 62.695 166.010 ;
        RECT 64.375 165.865 64.545 166.055 ;
        RECT 67.130 165.865 67.300 166.055 ;
        RECT 68.515 165.845 68.685 166.035 ;
        RECT 68.975 165.845 69.145 166.055 ;
        RECT 69.435 165.865 69.605 166.055 ;
        RECT 72.195 165.865 72.365 166.055 ;
        RECT 74.030 166.005 74.200 166.035 ;
        RECT 74.030 165.895 74.210 166.005 ;
        RECT 74.030 165.845 74.200 165.895 ;
        RECT 74.770 165.865 74.940 166.055 ;
        RECT 74.955 165.845 75.125 166.035 ;
        RECT 78.690 165.895 78.810 166.005 ;
        RECT 79.740 165.845 79.910 166.035 ;
        RECT 82.500 165.865 82.670 166.055 ;
        RECT 86.640 165.865 86.810 166.055 ;
        RECT 97.035 166.035 97.205 166.055 ;
        RECT 89.675 165.845 89.845 166.035 ;
        RECT 93.350 165.845 93.520 166.035 ;
        RECT 97.030 165.865 97.205 166.035 ;
        RECT 97.550 165.895 97.670 166.005 ;
        RECT 97.955 165.865 98.125 166.055 ;
        RECT 97.030 165.845 97.200 165.865 ;
        RECT 98.415 165.845 98.585 166.035 ;
        RECT 98.875 165.845 99.045 166.035 ;
        RECT 100.770 165.895 100.890 166.005 ;
        RECT 101.175 165.845 101.345 166.035 ;
        RECT 105.040 165.865 105.210 166.055 ;
        RECT 108.995 165.865 109.165 166.055 ;
        RECT 111.295 165.845 111.465 166.035 ;
        RECT 111.750 166.005 111.920 166.055 ;
        RECT 111.750 165.895 111.930 166.005 ;
        RECT 111.750 165.865 111.920 165.895 ;
        RECT 113.135 165.845 113.305 166.055 ;
        RECT 22.835 165.035 24.205 165.845 ;
        RECT 24.585 165.165 33.865 165.845 ;
        RECT 33.985 165.165 37.450 165.845 ;
        RECT 37.665 165.165 41.130 165.845 ;
        RECT 41.345 165.165 44.810 165.845 ;
        RECT 45.025 165.165 48.490 165.845 ;
        RECT 24.585 165.045 26.920 165.165 ;
        RECT 24.585 164.935 25.505 165.045 ;
        RECT 31.585 164.945 32.505 165.165 ;
        RECT 36.530 164.935 37.450 165.165 ;
        RECT 40.210 164.935 41.130 165.165 ;
        RECT 43.890 164.935 44.810 165.165 ;
        RECT 47.570 164.935 48.490 165.165 ;
        RECT 48.605 164.975 49.035 165.760 ;
        RECT 49.515 165.035 51.345 165.845 ;
        RECT 51.355 165.165 55.255 165.845 ;
        RECT 55.725 165.165 59.625 165.845 ;
        RECT 51.355 164.935 52.285 165.165 ;
        RECT 58.695 164.935 59.625 165.165 ;
        RECT 59.635 165.165 68.825 165.845 ;
        RECT 68.835 165.165 70.665 165.845 ;
        RECT 59.635 164.935 60.555 165.165 ;
        RECT 63.385 164.945 64.315 165.165 ;
        RECT 69.320 164.935 70.665 165.165 ;
        RECT 70.870 164.935 74.345 165.845 ;
        RECT 74.365 164.975 74.795 165.760 ;
        RECT 74.815 165.065 76.185 165.845 ;
        RECT 76.425 165.165 80.325 165.845 ;
        RECT 79.395 164.935 80.325 165.165 ;
        RECT 80.705 165.165 89.985 165.845 ;
        RECT 80.705 165.045 83.040 165.165 ;
        RECT 80.705 164.935 81.625 165.045 ;
        RECT 87.705 164.945 88.625 165.165 ;
        RECT 90.190 164.935 93.665 165.845 ;
        RECT 93.870 164.935 97.345 165.845 ;
        RECT 97.355 165.065 98.725 165.845 ;
        RECT 98.735 165.065 100.105 165.845 ;
        RECT 100.125 164.975 100.555 165.760 ;
        RECT 101.045 164.935 102.395 165.845 ;
        RECT 102.415 165.165 111.605 165.845 ;
        RECT 102.415 164.935 103.335 165.165 ;
        RECT 106.165 164.945 107.095 165.165 ;
        RECT 112.075 165.035 113.445 165.845 ;
      LAYER nwell ;
        RECT 22.640 161.815 113.640 164.645 ;
      LAYER pwell ;
        RECT 22.835 160.615 24.205 161.425 ;
        RECT 24.585 161.415 25.505 161.525 ;
        RECT 24.585 161.295 26.920 161.415 ;
        RECT 31.585 161.295 32.505 161.515 ;
        RECT 24.585 160.615 33.865 161.295 ;
        RECT 33.875 160.615 35.245 161.395 ;
        RECT 35.725 160.700 36.155 161.485 ;
        RECT 36.185 160.615 37.535 161.525 ;
        RECT 39.305 161.415 40.225 161.525 ;
        RECT 37.555 160.615 38.925 161.395 ;
        RECT 39.305 161.295 41.640 161.415 ;
        RECT 46.305 161.295 47.225 161.515 ;
        RECT 48.595 161.295 49.525 161.525 ;
        RECT 56.310 161.295 57.230 161.525 ;
        RECT 39.305 160.615 48.585 161.295 ;
        RECT 48.595 160.615 52.495 161.295 ;
        RECT 53.765 160.615 57.230 161.295 ;
        RECT 57.335 161.295 58.265 161.525 ;
        RECT 57.335 160.615 61.235 161.295 ;
        RECT 61.485 160.700 61.915 161.485 ;
        RECT 61.935 160.615 65.410 161.525 ;
        RECT 65.615 160.615 66.985 161.395 ;
        RECT 67.190 160.615 70.665 161.525 ;
        RECT 70.675 160.615 74.150 161.525 ;
        RECT 74.725 161.415 75.645 161.525 ;
        RECT 74.725 161.295 77.060 161.415 ;
        RECT 81.725 161.295 82.645 161.515 ;
        RECT 74.725 160.615 84.005 161.295 ;
        RECT 84.025 160.615 85.375 161.525 ;
        RECT 85.855 160.615 87.225 161.395 ;
        RECT 87.245 160.700 87.675 161.485 ;
        RECT 87.695 160.615 89.065 161.425 ;
        RECT 89.075 160.615 92.550 161.525 ;
        RECT 92.755 160.615 96.230 161.525 ;
        RECT 96.435 160.615 99.910 161.525 ;
        RECT 101.045 160.615 102.395 161.525 ;
        RECT 103.775 161.295 104.695 161.515 ;
        RECT 110.775 161.415 111.695 161.525 ;
        RECT 109.360 161.295 111.695 161.415 ;
        RECT 102.415 160.615 111.695 161.295 ;
        RECT 112.075 160.615 113.445 161.425 ;
        RECT 22.975 160.405 23.145 160.615 ;
        RECT 24.815 160.450 24.975 160.560 ;
        RECT 28.680 160.405 28.850 160.595 ;
        RECT 33.555 160.425 33.725 160.615 ;
        RECT 34.935 160.425 35.105 160.615 ;
        RECT 35.450 160.455 35.570 160.565 ;
        RECT 37.235 160.425 37.405 160.615 ;
        RECT 38.615 160.405 38.785 160.615 ;
        RECT 48.275 160.595 48.445 160.615 ;
        RECT 39.350 160.405 39.520 160.595 ;
        RECT 43.270 160.455 43.390 160.565 ;
        RECT 43.675 160.405 43.845 160.595 ;
        RECT 48.270 160.425 48.445 160.595 ;
        RECT 49.010 160.425 49.180 160.615 ;
        RECT 48.270 160.405 48.440 160.425 ;
        RECT 50.115 160.405 50.285 160.595 ;
        RECT 50.575 160.405 50.745 160.595 ;
        RECT 51.960 160.405 52.130 160.595 ;
        RECT 53.335 160.460 53.495 160.570 ;
        RECT 53.795 160.425 53.965 160.615 ;
        RECT 57.750 160.425 57.920 160.615 ;
        RECT 58.850 160.405 59.020 160.595 ;
        RECT 62.080 160.425 62.250 160.615 ;
        RECT 65.755 160.425 65.925 160.615 ;
        RECT 68.055 160.405 68.225 160.595 ;
        RECT 68.515 160.405 68.685 160.595 ;
        RECT 70.350 160.565 70.520 160.615 ;
        RECT 70.350 160.455 70.530 160.565 ;
        RECT 70.350 160.425 70.520 160.455 ;
        RECT 70.820 160.405 70.990 160.615 ;
        RECT 74.955 160.405 75.125 160.595 ;
        RECT 76.850 160.455 76.970 160.565 ;
        RECT 78.175 160.405 78.345 160.595 ;
        RECT 79.555 160.405 79.725 160.595 ;
        RECT 80.015 160.405 80.185 160.595 ;
        RECT 81.395 160.405 81.565 160.595 ;
        RECT 83.695 160.425 83.865 160.615 ;
        RECT 85.075 160.425 85.245 160.615 ;
        RECT 85.590 160.455 85.710 160.565 ;
        RECT 85.995 160.425 86.165 160.615 ;
        RECT 88.755 160.425 88.925 160.615 ;
        RECT 89.220 160.425 89.390 160.615 ;
        RECT 91.515 160.405 91.685 160.595 ;
        RECT 92.435 160.450 92.595 160.560 ;
        RECT 92.900 160.405 93.070 160.615 ;
        RECT 96.580 160.405 96.750 160.615 ;
        RECT 100.715 160.460 100.875 160.570 ;
        RECT 101.175 160.425 101.345 160.615 ;
        RECT 102.555 160.425 102.725 160.615 ;
        RECT 105.040 160.405 105.210 160.595 ;
        RECT 106.050 160.405 106.220 160.595 ;
        RECT 110.835 160.405 111.005 160.595 ;
        RECT 111.755 160.450 111.915 160.560 ;
        RECT 113.135 160.405 113.305 160.615 ;
        RECT 22.835 159.595 24.205 160.405 ;
        RECT 25.365 159.725 29.265 160.405 ;
        RECT 28.335 159.495 29.265 159.725 ;
        RECT 29.645 159.725 38.925 160.405 ;
        RECT 38.935 159.725 42.835 160.405 ;
        RECT 29.645 159.605 31.980 159.725 ;
        RECT 29.645 159.495 30.565 159.605 ;
        RECT 36.645 159.505 37.565 159.725 ;
        RECT 38.935 159.495 39.865 159.725 ;
        RECT 43.535 159.625 44.905 160.405 ;
        RECT 45.110 159.495 48.585 160.405 ;
        RECT 48.605 159.535 49.035 160.320 ;
        RECT 49.055 159.595 50.425 160.405 ;
        RECT 50.435 159.625 51.805 160.405 ;
        RECT 51.815 159.495 55.290 160.405 ;
        RECT 55.690 159.495 59.165 160.405 ;
        RECT 59.260 159.725 68.365 160.405 ;
        RECT 68.375 159.725 70.205 160.405 ;
        RECT 68.860 159.495 70.205 159.725 ;
        RECT 70.675 159.495 74.150 160.405 ;
        RECT 74.365 159.535 74.795 160.320 ;
        RECT 74.815 159.725 76.645 160.405 ;
        RECT 75.300 159.495 76.645 159.725 ;
        RECT 77.125 159.495 78.475 160.405 ;
        RECT 78.505 159.495 79.855 160.405 ;
        RECT 79.875 159.625 81.245 160.405 ;
        RECT 81.255 159.625 82.625 160.405 ;
        RECT 82.635 159.725 91.825 160.405 ;
        RECT 82.635 159.495 83.555 159.725 ;
        RECT 86.385 159.505 87.315 159.725 ;
        RECT 92.755 159.495 96.230 160.405 ;
        RECT 96.435 159.495 99.910 160.405 ;
        RECT 100.125 159.535 100.555 160.320 ;
        RECT 101.725 159.725 105.625 160.405 ;
        RECT 104.695 159.495 105.625 159.725 ;
        RECT 105.635 159.725 109.535 160.405 ;
        RECT 105.635 159.495 106.565 159.725 ;
        RECT 109.775 159.625 111.145 160.405 ;
        RECT 112.075 159.595 113.445 160.405 ;
      LAYER nwell ;
        RECT 22.640 156.375 113.640 159.205 ;
      LAYER pwell ;
        RECT 22.835 155.175 24.205 155.985 ;
        RECT 24.215 155.175 27.885 155.985 ;
        RECT 27.905 155.175 29.255 156.085 ;
        RECT 29.275 155.175 30.645 155.955 ;
        RECT 30.665 155.175 32.015 156.085 ;
        RECT 32.230 155.175 35.705 156.085 ;
        RECT 35.725 155.260 36.155 156.045 ;
        RECT 36.635 155.175 38.465 155.985 ;
        RECT 38.475 155.175 41.950 156.085 ;
        RECT 42.615 155.175 46.090 156.085 ;
        RECT 46.665 155.975 47.585 156.085 ;
        RECT 46.665 155.855 49.000 155.975 ;
        RECT 53.665 155.855 54.585 156.075 ;
        RECT 46.665 155.175 55.945 155.855 ;
        RECT 55.965 155.175 57.315 156.085 ;
        RECT 59.990 155.855 60.910 156.085 ;
        RECT 57.445 155.175 60.910 155.855 ;
        RECT 61.485 155.260 61.915 156.045 ;
        RECT 61.945 155.175 63.295 156.085 ;
        RECT 63.315 155.855 64.660 156.085 ;
        RECT 65.640 155.855 66.985 156.085 ;
        RECT 67.480 155.855 68.825 156.085 ;
        RECT 69.320 155.855 70.665 156.085 ;
        RECT 63.315 155.175 65.145 155.855 ;
        RECT 65.155 155.175 66.985 155.855 ;
        RECT 66.995 155.175 68.825 155.855 ;
        RECT 68.835 155.175 70.665 155.855 ;
        RECT 70.675 155.175 73.395 156.085 ;
        RECT 73.920 155.855 75.265 156.085 ;
        RECT 73.435 155.175 75.265 155.855 ;
        RECT 75.735 155.175 77.565 155.985 ;
        RECT 77.585 155.175 78.935 156.085 ;
        RECT 81.610 155.855 82.530 156.085 ;
        RECT 85.835 155.855 86.765 156.085 ;
        RECT 79.065 155.175 82.530 155.855 ;
        RECT 82.865 155.175 86.765 155.855 ;
        RECT 87.245 155.260 87.675 156.045 ;
        RECT 89.960 155.885 90.905 156.085 ;
        RECT 92.720 155.885 93.665 156.085 ;
        RECT 88.155 155.205 90.905 155.885 ;
        RECT 90.915 155.205 93.665 155.885 ;
        RECT 22.975 154.965 23.145 155.175 ;
        RECT 24.410 155.015 24.530 155.125 ;
        RECT 26.195 154.965 26.365 155.155 ;
        RECT 26.655 154.965 26.825 155.155 ;
        RECT 27.575 154.985 27.745 155.175 ;
        RECT 28.955 154.985 29.125 155.175 ;
        RECT 29.415 154.985 29.585 155.175 ;
        RECT 30.795 154.985 30.965 155.175 ;
        RECT 31.440 154.965 31.610 155.155 ;
        RECT 32.230 155.015 32.350 155.125 ;
        RECT 34.935 154.965 35.105 155.155 ;
        RECT 35.390 154.985 35.560 155.175 ;
        RECT 38.155 155.155 38.325 155.175 ;
        RECT 36.370 155.015 36.490 155.125 ;
        RECT 22.835 154.155 24.205 154.965 ;
        RECT 24.675 154.155 26.505 154.965 ;
        RECT 26.525 154.055 27.875 154.965 ;
        RECT 28.125 154.285 32.025 154.965 ;
        RECT 31.095 154.055 32.025 154.285 ;
        RECT 32.495 154.155 35.245 154.965 ;
        RECT 35.255 154.935 36.200 154.965 ;
        RECT 37.690 154.935 37.860 155.155 ;
        RECT 38.155 154.985 38.330 155.155 ;
        RECT 38.620 154.985 38.790 155.175 ;
        RECT 38.160 154.965 38.330 154.985 ;
        RECT 35.255 154.255 38.005 154.935 ;
        RECT 35.255 154.055 36.200 154.255 ;
        RECT 38.015 154.055 41.490 154.965 ;
        RECT 41.840 154.935 42.010 155.155 ;
        RECT 42.350 155.015 42.470 155.125 ;
        RECT 42.760 154.985 42.930 155.175 ;
        RECT 48.000 154.965 48.170 155.155 ;
        RECT 49.200 154.965 49.370 155.155 ;
        RECT 52.930 155.015 53.050 155.125 ;
        RECT 53.335 154.965 53.505 155.155 ;
        RECT 55.635 154.985 55.805 155.175 ;
        RECT 56.095 154.985 56.265 155.175 ;
        RECT 57.475 154.985 57.645 155.175 ;
        RECT 61.210 155.015 61.330 155.125 ;
        RECT 62.995 154.985 63.165 155.175 ;
        RECT 63.915 154.965 64.085 155.155 ;
        RECT 64.835 154.985 65.005 155.175 ;
        RECT 65.295 154.985 65.465 155.175 ;
        RECT 67.135 154.965 67.305 155.175 ;
        RECT 68.975 154.985 69.145 155.175 ;
        RECT 69.895 154.965 70.065 155.155 ;
        RECT 70.815 154.985 70.985 155.175 ;
        RECT 71.275 154.965 71.445 155.155 ;
        RECT 71.735 154.965 71.905 155.155 ;
        RECT 73.575 154.985 73.745 155.175 ;
        RECT 75.010 155.015 75.130 155.125 ;
        RECT 75.470 155.015 75.590 155.125 ;
        RECT 76.795 154.965 76.965 155.155 ;
        RECT 77.255 154.985 77.425 155.175 ;
        RECT 77.715 154.985 77.885 155.175 ;
        RECT 79.095 154.985 79.265 155.175 ;
        RECT 86.180 154.985 86.350 155.175 ;
        RECT 86.455 154.965 86.625 155.155 ;
        RECT 87.835 155.125 88.005 155.155 ;
        RECT 86.970 155.015 87.090 155.125 ;
        RECT 87.375 155.010 87.535 155.120 ;
        RECT 87.835 155.015 88.010 155.125 ;
        RECT 87.835 154.965 88.005 155.015 ;
        RECT 88.300 154.985 88.470 155.205 ;
        RECT 89.960 155.175 90.905 155.205 ;
        RECT 91.060 154.985 91.230 155.205 ;
        RECT 92.720 155.175 93.665 155.205 ;
        RECT 93.675 155.175 97.150 156.085 ;
        RECT 97.815 155.175 101.290 156.085 ;
        RECT 101.495 155.175 102.865 155.985 ;
        RECT 106.075 155.855 107.005 156.085 ;
        RECT 109.670 155.855 110.590 156.085 ;
        RECT 103.105 155.175 107.005 155.855 ;
        RECT 107.125 155.175 110.590 155.855 ;
        RECT 110.695 155.175 112.065 155.955 ;
        RECT 112.075 155.175 113.445 155.985 ;
        RECT 92.435 154.965 92.605 155.155 ;
        RECT 93.820 154.985 93.990 155.175 ;
        RECT 97.960 155.155 98.130 155.175 ;
        RECT 43.500 154.935 44.445 154.965 ;
        RECT 41.695 154.255 44.445 154.935 ;
        RECT 44.685 154.285 48.585 154.965 ;
        RECT 43.500 154.055 44.445 154.255 ;
        RECT 47.655 154.055 48.585 154.285 ;
        RECT 48.605 154.095 49.035 154.880 ;
        RECT 49.055 154.055 52.530 154.965 ;
        RECT 53.195 154.185 54.565 154.965 ;
        RECT 54.945 154.285 64.225 154.965 ;
        RECT 54.945 154.165 57.280 154.285 ;
        RECT 54.945 154.055 55.865 154.165 ;
        RECT 61.945 154.065 62.865 154.285 ;
        RECT 64.235 154.055 67.445 154.965 ;
        RECT 67.465 154.285 70.205 154.965 ;
        RECT 70.215 154.155 71.585 154.965 ;
        RECT 71.595 154.285 74.335 154.965 ;
        RECT 74.365 154.095 74.795 154.880 ;
        RECT 75.275 154.155 77.105 154.965 ;
        RECT 77.485 154.285 86.765 154.965 ;
        RECT 77.485 154.165 79.820 154.285 ;
        RECT 77.485 154.055 78.405 154.165 ;
        RECT 84.485 154.065 85.405 154.285 ;
        RECT 87.695 154.185 89.065 154.965 ;
        RECT 89.075 154.155 92.745 154.965 ;
        RECT 92.755 154.935 93.700 154.965 ;
        RECT 95.190 154.935 95.360 155.155 ;
        RECT 97.550 155.015 97.670 155.125 ;
        RECT 97.950 154.985 98.130 155.155 ;
        RECT 95.515 154.935 96.460 154.965 ;
        RECT 97.950 154.935 98.120 154.985 ;
        RECT 99.795 154.965 99.965 155.155 ;
        RECT 100.770 155.015 100.890 155.125 ;
        RECT 101.175 154.965 101.345 155.155 ;
        RECT 102.555 154.985 102.725 155.175 ;
        RECT 106.420 154.985 106.590 155.175 ;
        RECT 107.155 154.985 107.325 155.175 ;
        RECT 111.755 154.965 111.925 155.175 ;
        RECT 113.135 154.965 113.305 155.175 ;
        RECT 92.755 154.255 95.505 154.935 ;
        RECT 95.515 154.255 98.265 154.935 ;
        RECT 92.755 154.055 93.700 154.255 ;
        RECT 95.515 154.055 96.460 154.255 ;
        RECT 98.275 154.155 100.105 154.965 ;
        RECT 100.125 154.095 100.555 154.880 ;
        RECT 101.045 154.055 102.395 154.965 ;
        RECT 102.785 154.285 112.065 154.965 ;
        RECT 102.785 154.165 105.120 154.285 ;
        RECT 102.785 154.055 103.705 154.165 ;
        RECT 109.785 154.065 110.705 154.285 ;
        RECT 112.075 154.155 113.445 154.965 ;
      LAYER nwell ;
        RECT 22.640 150.935 113.640 153.765 ;
      LAYER pwell ;
        RECT 22.835 149.735 24.205 150.545 ;
        RECT 25.045 150.535 25.965 150.645 ;
        RECT 25.045 150.415 27.380 150.535 ;
        RECT 32.045 150.415 32.965 150.635 ;
        RECT 25.045 149.735 34.325 150.415 ;
        RECT 34.335 149.735 35.705 150.515 ;
        RECT 35.725 149.820 36.155 150.605 ;
        RECT 36.175 150.445 37.120 150.645 ;
        RECT 38.935 150.445 39.880 150.645 ;
        RECT 36.175 149.765 38.925 150.445 ;
        RECT 38.935 149.765 41.685 150.445 ;
        RECT 36.175 149.735 37.120 149.765 ;
        RECT 22.975 149.525 23.145 149.735 ;
        RECT 24.410 149.575 24.530 149.685 ;
        RECT 33.555 149.525 33.725 149.715 ;
        RECT 34.015 149.545 34.185 149.735 ;
        RECT 34.290 149.525 34.460 149.715 ;
        RECT 35.395 149.545 35.565 149.735 ;
        RECT 38.610 149.715 38.780 149.765 ;
        RECT 38.935 149.735 39.880 149.765 ;
        RECT 38.210 149.575 38.330 149.685 ;
        RECT 38.610 149.545 38.785 149.715 ;
        RECT 40.915 149.545 41.085 149.715 ;
        RECT 41.370 149.545 41.540 149.765 ;
        RECT 41.695 149.735 45.170 150.645 ;
        RECT 45.375 149.735 48.850 150.645 ;
        RECT 52.715 150.415 53.645 150.645 ;
        RECT 49.745 149.735 53.645 150.415 ;
        RECT 54.115 149.735 57.590 150.645 ;
        RECT 60.450 150.415 61.370 150.645 ;
        RECT 57.905 149.735 61.370 150.415 ;
        RECT 61.485 149.820 61.915 150.605 ;
        RECT 61.935 150.415 62.855 150.645 ;
        RECT 65.685 150.415 66.615 150.635 ;
        RECT 71.135 150.445 72.080 150.645 ;
        RECT 61.935 149.735 71.125 150.415 ;
        RECT 71.135 149.765 73.885 150.445 ;
        RECT 71.135 149.735 72.080 149.765 ;
        RECT 41.840 149.545 42.010 149.735 ;
        RECT 45.055 149.545 45.225 149.715 ;
        RECT 45.520 149.545 45.690 149.735 ;
        RECT 38.635 149.525 38.785 149.545 ;
        RECT 40.935 149.525 41.085 149.545 ;
        RECT 45.055 149.525 45.205 149.545 ;
        RECT 46.895 149.525 47.065 149.715 ;
        RECT 47.355 149.525 47.525 149.715 ;
        RECT 49.250 149.575 49.370 149.685 ;
        RECT 53.060 149.545 53.230 149.735 ;
        RECT 53.850 149.575 53.970 149.685 ;
        RECT 54.260 149.545 54.430 149.735 ;
        RECT 57.935 149.545 58.105 149.735 ;
        RECT 70.815 149.715 70.985 149.735 ;
        RECT 58.395 149.525 58.565 149.715 ;
        RECT 60.235 149.525 60.405 149.715 ;
        RECT 60.695 149.525 60.865 149.715 ;
        RECT 65.480 149.525 65.650 149.715 ;
        RECT 66.215 149.525 66.385 149.715 ;
        RECT 67.650 149.575 67.770 149.685 ;
        RECT 22.835 148.715 24.205 149.525 ;
        RECT 24.585 148.845 33.865 149.525 ;
        RECT 33.875 148.845 37.775 149.525 ;
        RECT 24.585 148.725 26.920 148.845 ;
        RECT 24.585 148.615 25.505 148.725 ;
        RECT 31.585 148.625 32.505 148.845 ;
        RECT 33.875 148.615 34.805 148.845 ;
        RECT 38.635 148.705 40.565 149.525 ;
        RECT 40.935 148.705 42.865 149.525 ;
        RECT 39.615 148.615 40.565 148.705 ;
        RECT 41.915 148.615 42.865 148.705 ;
        RECT 43.275 148.705 45.205 149.525 ;
        RECT 45.375 148.715 47.205 149.525 ;
        RECT 43.275 148.615 44.225 148.705 ;
        RECT 47.225 148.615 48.575 149.525 ;
        RECT 48.605 148.655 49.035 149.440 ;
        RECT 49.425 148.845 58.705 149.525 ;
        RECT 49.425 148.725 51.760 148.845 ;
        RECT 49.425 148.615 50.345 148.725 ;
        RECT 56.425 148.625 57.345 148.845 ;
        RECT 58.715 148.715 60.545 149.525 ;
        RECT 60.565 148.615 61.915 149.525 ;
        RECT 62.165 148.845 66.065 149.525 ;
        RECT 65.135 148.615 66.065 148.845 ;
        RECT 66.075 148.745 67.445 149.525 ;
        RECT 68.060 149.495 68.230 149.715 ;
        RECT 70.815 149.545 70.990 149.715 ;
        RECT 73.570 149.545 73.740 149.765 ;
        RECT 73.895 149.735 77.370 150.645 ;
        RECT 81.235 150.415 82.165 150.645 ;
        RECT 78.265 149.735 82.165 150.415 ;
        RECT 82.175 150.415 83.105 150.645 ;
        RECT 82.175 149.735 86.075 150.415 ;
        RECT 87.245 149.820 87.675 150.605 ;
        RECT 88.155 149.735 93.665 150.545 ;
        RECT 93.870 149.735 97.345 150.645 ;
        RECT 97.355 149.735 100.830 150.645 ;
        RECT 101.505 149.735 102.855 150.645 ;
        RECT 106.075 150.415 107.005 150.645 ;
        RECT 103.105 149.735 107.005 150.415 ;
        RECT 107.935 149.735 109.305 150.515 ;
        RECT 109.315 149.735 112.065 150.545 ;
        RECT 112.075 149.735 113.445 150.545 ;
        RECT 74.040 149.545 74.210 149.735 ;
        RECT 75.415 149.570 75.575 149.680 ;
        RECT 70.820 149.525 70.990 149.545 ;
        RECT 76.795 149.525 76.965 149.715 ;
        RECT 77.770 149.575 77.890 149.685 ;
        RECT 81.580 149.545 81.750 149.735 ;
        RECT 82.590 149.545 82.760 149.735 ;
        RECT 86.455 149.525 86.625 149.715 ;
        RECT 86.915 149.580 87.075 149.690 ;
        RECT 87.835 149.685 88.005 149.715 ;
        RECT 87.835 149.575 88.010 149.685 ;
        RECT 87.835 149.525 88.005 149.575 ;
        RECT 88.755 149.570 88.915 149.680 ;
        RECT 69.720 149.495 70.665 149.525 ;
        RECT 67.915 148.815 70.665 149.495 ;
        RECT 69.720 148.615 70.665 148.815 ;
        RECT 70.675 148.615 74.150 149.525 ;
        RECT 74.365 148.655 74.795 149.440 ;
        RECT 75.745 148.615 77.095 149.525 ;
        RECT 77.485 148.845 86.765 149.525 ;
        RECT 77.485 148.725 79.820 148.845 ;
        RECT 77.485 148.615 78.405 148.725 ;
        RECT 84.485 148.625 85.405 148.845 ;
        RECT 86.775 148.745 88.145 149.525 ;
        RECT 89.220 149.495 89.390 149.715 ;
        RECT 91.980 149.525 92.150 149.715 ;
        RECT 93.355 149.545 93.525 149.735 ;
        RECT 90.880 149.495 91.825 149.525 ;
        RECT 89.075 148.815 91.825 149.495 ;
        RECT 90.880 148.615 91.825 148.815 ;
        RECT 91.835 148.615 95.310 149.525 ;
        RECT 95.660 149.495 95.830 149.715 ;
        RECT 97.030 149.545 97.200 149.735 ;
        RECT 97.500 149.545 97.670 149.735 ;
        RECT 99.795 149.525 99.965 149.715 ;
        RECT 101.230 149.575 101.350 149.685 ;
        RECT 101.635 149.545 101.805 149.735 ;
        RECT 102.095 149.525 102.265 149.715 ;
        RECT 106.420 149.545 106.590 149.735 ;
        RECT 107.615 149.580 107.775 149.690 ;
        RECT 108.075 149.545 108.245 149.735 ;
        RECT 111.755 149.525 111.925 149.735 ;
        RECT 113.135 149.525 113.305 149.735 ;
        RECT 97.320 149.495 98.265 149.525 ;
        RECT 95.515 148.815 98.265 149.495 ;
        RECT 97.320 148.615 98.265 148.815 ;
        RECT 98.275 148.715 100.105 149.525 ;
        RECT 100.125 148.655 100.555 149.440 ;
        RECT 100.575 148.715 102.405 149.525 ;
        RECT 102.785 148.845 112.065 149.525 ;
        RECT 102.785 148.725 105.120 148.845 ;
        RECT 102.785 148.615 103.705 148.725 ;
        RECT 109.785 148.625 110.705 148.845 ;
        RECT 112.075 148.715 113.445 149.525 ;
      LAYER nwell ;
        RECT 22.640 145.495 113.640 148.325 ;
      LAYER pwell ;
        RECT 22.835 144.295 24.205 145.105 ;
        RECT 24.685 144.295 26.035 145.205 ;
        RECT 27.415 144.975 28.335 145.195 ;
        RECT 34.415 145.095 35.335 145.205 ;
        RECT 33.000 144.975 35.335 145.095 ;
        RECT 26.055 144.295 35.335 144.975 ;
        RECT 35.725 144.380 36.155 145.165 ;
        RECT 37.775 145.115 38.725 145.205 ;
        RECT 36.795 144.295 38.725 145.115 ;
        RECT 38.935 144.975 39.865 145.205 ;
        RECT 45.135 145.115 46.085 145.205 ;
        RECT 47.435 145.115 48.385 145.205 ;
        RECT 38.935 144.295 42.835 144.975 ;
        RECT 44.155 144.295 46.085 145.115 ;
        RECT 46.455 144.295 48.385 145.115 ;
        RECT 49.055 144.295 51.805 145.105 ;
        RECT 53.620 145.005 54.565 145.205 ;
        RECT 51.815 144.325 54.565 145.005 ;
        RECT 22.975 144.085 23.145 144.295 ;
        RECT 24.410 144.135 24.530 144.245 ;
        RECT 25.735 144.105 25.905 144.295 ;
        RECT 26.195 144.085 26.365 144.295 ;
        RECT 36.795 144.275 36.945 144.295 ;
        RECT 26.655 144.085 26.825 144.275 ;
        RECT 28.035 144.085 28.205 144.275 ;
        RECT 30.335 144.085 30.505 144.275 ;
        RECT 30.795 144.085 30.965 144.275 ;
        RECT 32.450 144.085 32.620 144.275 ;
        RECT 36.315 144.245 36.485 144.275 ;
        RECT 36.315 144.135 36.490 144.245 ;
        RECT 36.315 144.085 36.485 144.135 ;
        RECT 36.775 144.105 36.945 144.275 ;
        RECT 39.350 144.105 39.520 144.295 ;
        RECT 44.155 144.275 44.305 144.295 ;
        RECT 46.455 144.275 46.605 144.295 ;
        RECT 43.675 144.140 43.835 144.250 ;
        RECT 44.135 144.105 44.305 144.275 ;
        RECT 46.435 144.105 46.605 144.275 ;
        RECT 22.835 143.275 24.205 144.085 ;
        RECT 24.675 143.275 26.505 144.085 ;
        RECT 26.525 143.175 27.875 144.085 ;
        RECT 27.895 143.305 29.265 144.085 ;
        RECT 29.275 143.305 30.645 144.085 ;
        RECT 30.665 143.175 32.015 144.085 ;
        RECT 32.035 143.405 35.935 144.085 ;
        RECT 36.175 143.405 45.455 144.085 ;
        RECT 32.035 143.175 32.965 143.405 ;
        RECT 37.535 143.185 38.455 143.405 ;
        RECT 43.120 143.285 45.455 143.405 ;
        RECT 44.535 143.175 45.455 143.285 ;
        RECT 45.835 144.055 46.780 144.085 ;
        RECT 48.270 144.055 48.440 144.275 ;
        RECT 48.790 144.135 48.910 144.245 ;
        RECT 49.195 144.085 49.365 144.275 ;
        RECT 50.850 144.085 51.020 144.275 ;
        RECT 51.495 144.105 51.665 144.295 ;
        RECT 51.960 144.105 52.130 144.325 ;
        RECT 53.620 144.295 54.565 144.325 ;
        RECT 54.575 144.295 57.325 145.105 ;
        RECT 59.140 145.005 60.085 145.205 ;
        RECT 57.335 144.325 60.085 145.005 ;
        RECT 57.015 144.275 57.185 144.295 ;
        RECT 54.770 144.135 54.890 144.245 ;
        RECT 56.555 144.085 56.725 144.275 ;
        RECT 57.015 144.105 57.190 144.275 ;
        RECT 57.480 144.105 57.650 144.325 ;
        RECT 59.140 144.295 60.085 144.325 ;
        RECT 60.095 144.295 61.465 145.105 ;
        RECT 61.485 144.380 61.915 145.165 ;
        RECT 65.135 144.975 66.065 145.205 ;
        RECT 62.165 144.295 66.065 144.975 ;
        RECT 66.075 144.295 67.905 144.975 ;
        RECT 67.915 144.295 69.285 145.075 ;
        RECT 69.295 144.295 70.665 145.105 ;
        RECT 70.675 144.295 74.345 145.105 ;
        RECT 74.550 144.295 78.025 145.205 ;
        RECT 78.035 144.295 79.405 145.105 ;
        RECT 82.615 144.975 83.545 145.205 ;
        RECT 79.645 144.295 83.545 144.975 ;
        RECT 83.555 144.295 84.925 145.075 ;
        RECT 85.395 144.295 87.225 145.105 ;
        RECT 87.245 144.380 87.675 145.165 ;
        RECT 88.835 145.115 89.785 145.205 ;
        RECT 87.855 144.295 89.785 145.115 ;
        RECT 93.195 144.975 94.125 145.205 ;
        RECT 90.225 144.295 94.125 144.975 ;
        RECT 94.335 145.115 95.285 145.205 ;
        RECT 97.095 145.115 98.045 145.205 ;
        RECT 94.335 144.295 96.265 145.115 ;
        RECT 97.095 144.295 99.025 145.115 ;
        RECT 99.195 144.295 101.945 145.105 ;
        RECT 105.155 144.975 106.085 145.205 ;
        RECT 102.185 144.295 106.085 144.975 ;
        RECT 106.095 144.295 107.465 145.105 ;
        RECT 107.475 144.295 108.845 145.075 ;
        RECT 109.315 144.295 112.065 145.105 ;
        RECT 112.075 144.295 113.445 145.105 ;
        RECT 61.155 144.105 61.325 144.295 ;
        RECT 65.480 144.105 65.650 144.295 ;
        RECT 66.215 144.105 66.385 144.295 ;
        RECT 68.055 144.105 68.225 144.295 ;
        RECT 57.020 144.085 57.190 144.105 ;
        RECT 69.895 144.085 70.065 144.275 ;
        RECT 70.355 144.245 70.525 144.295 ;
        RECT 74.035 144.275 74.205 144.295 ;
        RECT 70.355 144.135 70.530 144.245 ;
        RECT 70.355 144.105 70.525 144.135 ;
        RECT 74.030 144.105 74.205 144.275 ;
        RECT 74.030 144.085 74.200 144.105 ;
        RECT 45.835 143.375 48.585 144.055 ;
        RECT 45.835 143.175 46.780 143.375 ;
        RECT 48.605 143.215 49.035 144.000 ;
        RECT 49.065 143.175 50.415 144.085 ;
        RECT 50.435 143.405 54.335 144.085 ;
        RECT 50.435 143.175 51.365 143.405 ;
        RECT 55.035 143.275 56.865 144.085 ;
        RECT 56.875 143.175 60.350 144.085 ;
        RECT 60.925 143.405 70.205 144.085 ;
        RECT 60.925 143.285 63.260 143.405 ;
        RECT 60.925 143.175 61.845 143.285 ;
        RECT 67.925 143.185 68.845 143.405 ;
        RECT 70.870 143.175 74.345 144.085 ;
        RECT 74.960 144.055 75.130 144.275 ;
        RECT 77.710 144.105 77.880 144.295 ;
        RECT 79.095 144.105 79.265 144.295 ;
        RECT 82.960 144.105 83.130 144.295 ;
        RECT 83.695 144.105 83.865 144.295 ;
        RECT 85.130 144.135 85.250 144.245 ;
        RECT 86.915 144.085 87.085 144.295 ;
        RECT 87.855 144.275 88.005 144.295 ;
        RECT 87.835 144.105 88.005 144.275 ;
        RECT 93.540 144.105 93.710 144.295 ;
        RECT 96.115 144.275 96.265 144.295 ;
        RECT 98.875 144.275 99.025 144.295 ;
        RECT 96.115 144.105 96.285 144.275 ;
        RECT 96.575 144.245 96.745 144.275 ;
        RECT 96.575 144.135 96.750 144.245 ;
        RECT 96.575 144.085 96.745 144.135 ;
        RECT 98.875 144.105 99.045 144.275 ;
        RECT 99.795 144.130 99.955 144.240 ;
        RECT 98.875 144.085 99.025 144.105 ;
        RECT 100.715 144.085 100.885 144.275 ;
        RECT 101.635 144.105 101.805 144.295 ;
        RECT 105.500 144.105 105.670 144.295 ;
        RECT 107.155 144.105 107.325 144.295 ;
        RECT 107.615 144.105 107.785 144.295 ;
        RECT 109.050 144.135 109.170 144.245 ;
        RECT 111.295 144.085 111.465 144.275 ;
        RECT 111.755 144.245 111.925 144.295 ;
        RECT 111.755 144.135 111.930 144.245 ;
        RECT 111.755 144.105 111.925 144.135 ;
        RECT 113.135 144.085 113.305 144.295 ;
        RECT 76.620 144.055 77.565 144.085 ;
        RECT 74.365 143.215 74.795 144.000 ;
        RECT 74.815 143.375 77.565 144.055 ;
        RECT 76.620 143.175 77.565 143.375 ;
        RECT 77.945 143.405 87.225 144.085 ;
        RECT 87.605 143.405 96.885 144.085 ;
        RECT 77.945 143.285 80.280 143.405 ;
        RECT 77.945 143.175 78.865 143.285 ;
        RECT 84.945 143.185 85.865 143.405 ;
        RECT 87.605 143.285 89.940 143.405 ;
        RECT 87.605 143.175 88.525 143.285 ;
        RECT 94.605 143.185 95.525 143.405 ;
        RECT 97.095 143.265 99.025 144.085 ;
        RECT 97.095 143.175 98.045 143.265 ;
        RECT 100.125 143.215 100.555 144.000 ;
        RECT 100.585 143.175 101.935 144.085 ;
        RECT 102.325 143.405 111.605 144.085 ;
        RECT 102.325 143.285 104.660 143.405 ;
        RECT 102.325 143.175 103.245 143.285 ;
        RECT 109.325 143.185 110.245 143.405 ;
        RECT 112.075 143.275 113.445 144.085 ;
      LAYER nwell ;
        RECT 22.640 140.055 113.640 142.885 ;
      LAYER pwell ;
        RECT 22.835 138.855 24.205 139.665 ;
        RECT 24.215 138.855 26.045 139.665 ;
        RECT 26.065 138.855 27.415 139.765 ;
        RECT 27.435 138.855 28.805 139.635 ;
        RECT 28.815 139.535 29.745 139.765 ;
        RECT 28.815 138.855 32.715 139.535 ;
        RECT 32.965 138.855 35.705 139.535 ;
        RECT 35.725 138.940 36.155 139.725 ;
        RECT 36.195 138.855 47.205 139.765 ;
        RECT 47.585 139.655 48.505 139.765 ;
        RECT 47.585 139.535 49.920 139.655 ;
        RECT 54.585 139.535 55.505 139.755 ;
        RECT 58.680 139.565 59.625 139.765 ;
        RECT 47.585 138.855 56.865 139.535 ;
        RECT 56.875 138.885 59.625 139.565 ;
        RECT 22.975 138.645 23.145 138.855 ;
        RECT 24.410 138.695 24.530 138.805 ;
        RECT 24.815 138.645 24.985 138.835 ;
        RECT 25.735 138.665 25.905 138.855 ;
        RECT 26.195 138.665 26.365 138.855 ;
        RECT 28.495 138.665 28.665 138.855 ;
        RECT 29.230 138.665 29.400 138.855 ;
        RECT 34.475 138.645 34.645 138.835 ;
        RECT 35.395 138.665 35.565 138.855 ;
        RECT 44.595 138.645 44.765 138.835 ;
        RECT 45.060 138.645 45.230 138.835 ;
        RECT 46.890 138.665 47.060 138.855 ;
        RECT 49.195 138.645 49.365 138.835 ;
        RECT 56.555 138.665 56.725 138.855 ;
        RECT 57.020 138.665 57.190 138.885 ;
        RECT 58.680 138.855 59.625 138.885 ;
        RECT 59.635 138.855 61.465 139.665 ;
        RECT 61.485 138.940 61.915 139.725 ;
        RECT 62.865 138.855 64.215 139.765 ;
        RECT 66.275 139.675 67.225 139.765 ;
        RECT 81.455 139.675 82.405 139.765 ;
        RECT 64.235 138.855 66.065 139.535 ;
        RECT 66.275 138.855 68.205 139.675 ;
        RECT 68.375 138.855 71.115 139.535 ;
        RECT 72.140 138.855 81.245 139.535 ;
        RECT 81.455 138.855 83.385 139.675 ;
        RECT 83.565 138.855 84.915 139.765 ;
        RECT 86.075 139.675 87.025 139.765 ;
        RECT 85.095 138.855 87.025 139.675 ;
        RECT 87.245 138.940 87.675 139.725 ;
        RECT 97.095 139.675 98.045 139.765 ;
        RECT 87.695 138.855 96.800 139.535 ;
        RECT 97.095 138.855 99.025 139.675 ;
        RECT 99.195 138.855 100.565 139.665 ;
        RECT 100.945 139.655 101.865 139.765 ;
        RECT 100.945 139.535 103.280 139.655 ;
        RECT 107.945 139.535 108.865 139.755 ;
        RECT 100.945 138.855 110.225 139.535 ;
        RECT 110.235 138.855 112.065 139.665 ;
        RECT 112.075 138.855 113.445 139.665 ;
        RECT 58.450 138.695 58.570 138.805 ;
        RECT 58.860 138.645 59.030 138.835 ;
        RECT 61.155 138.665 61.325 138.855 ;
        RECT 62.535 138.700 62.695 138.810 ;
        RECT 62.995 138.665 63.165 138.855 ;
        RECT 65.755 138.665 65.925 138.855 ;
        RECT 68.055 138.835 68.205 138.855 ;
        RECT 65.940 138.645 66.110 138.835 ;
        RECT 66.730 138.695 66.850 138.805 ;
        RECT 68.055 138.665 68.225 138.835 ;
        RECT 68.515 138.665 68.685 138.855 ;
        RECT 68.975 138.665 69.145 138.835 ;
        RECT 69.435 138.665 69.605 138.835 ;
        RECT 71.735 138.700 71.895 138.810 ;
        RECT 68.975 138.645 69.125 138.665 ;
        RECT 22.835 137.835 24.205 138.645 ;
        RECT 24.675 137.965 33.955 138.645 ;
        RECT 26.035 137.745 26.955 137.965 ;
        RECT 31.620 137.845 33.955 137.965 ;
        RECT 34.335 137.865 35.705 138.645 ;
        RECT 35.800 137.965 44.905 138.645 ;
        RECT 33.035 137.735 33.955 137.845 ;
        RECT 44.915 137.735 48.390 138.645 ;
        RECT 48.605 137.775 49.035 138.560 ;
        RECT 49.055 137.965 58.160 138.645 ;
        RECT 58.715 137.735 62.190 138.645 ;
        RECT 62.625 137.965 66.525 138.645 ;
        RECT 65.595 137.735 66.525 137.965 ;
        RECT 67.195 137.825 69.125 138.645 ;
        RECT 69.455 138.645 69.605 138.665 ;
        RECT 69.455 137.825 71.385 138.645 ;
        RECT 67.195 137.735 68.145 137.825 ;
        RECT 70.435 137.735 71.385 137.825 ;
        RECT 71.595 138.615 72.540 138.645 ;
        RECT 74.030 138.615 74.200 138.835 ;
        RECT 75.415 138.690 75.575 138.800 ;
        RECT 79.280 138.645 79.450 138.835 ;
        RECT 80.475 138.690 80.635 138.800 ;
        RECT 80.935 138.665 81.105 138.855 ;
        RECT 83.235 138.835 83.385 138.855 ;
        RECT 83.235 138.665 83.405 138.835 ;
        RECT 84.340 138.645 84.510 138.835 ;
        RECT 84.615 138.665 84.785 138.855 ;
        RECT 85.095 138.835 85.245 138.855 ;
        RECT 85.075 138.645 85.245 138.835 ;
        RECT 87.835 138.665 88.005 138.855 ;
        RECT 98.875 138.835 99.025 138.855 ;
        RECT 94.735 138.645 94.905 138.835 ;
        RECT 98.875 138.665 99.045 138.835 ;
        RECT 99.520 138.645 99.690 138.835 ;
        RECT 100.255 138.665 100.425 138.855 ;
        RECT 104.120 138.645 104.290 138.835 ;
        RECT 105.775 138.645 105.945 138.835 ;
        RECT 106.235 138.645 106.405 138.835 ;
        RECT 107.615 138.645 107.785 138.835 ;
        RECT 109.050 138.695 109.170 138.805 ;
        RECT 109.915 138.665 110.085 138.855 ;
        RECT 111.755 138.645 111.925 138.855 ;
        RECT 113.135 138.645 113.305 138.855 ;
        RECT 71.595 137.935 74.345 138.615 ;
        RECT 71.595 137.735 72.540 137.935 ;
        RECT 74.365 137.775 74.795 138.560 ;
        RECT 75.965 137.965 79.865 138.645 ;
        RECT 81.025 137.965 84.925 138.645 ;
        RECT 84.935 137.965 94.215 138.645 ;
        RECT 78.935 137.735 79.865 137.965 ;
        RECT 83.995 137.735 84.925 137.965 ;
        RECT 86.295 137.745 87.215 137.965 ;
        RECT 91.880 137.845 94.215 137.965 ;
        RECT 94.595 137.865 95.965 138.645 ;
        RECT 96.205 137.965 100.105 138.645 ;
        RECT 93.295 137.735 94.215 137.845 ;
        RECT 99.175 137.735 100.105 137.965 ;
        RECT 100.125 137.775 100.555 138.560 ;
        RECT 100.805 137.965 104.705 138.645 ;
        RECT 103.775 137.735 104.705 137.965 ;
        RECT 104.725 137.735 106.075 138.645 ;
        RECT 106.095 137.865 107.465 138.645 ;
        RECT 107.475 137.865 108.845 138.645 ;
        RECT 109.315 137.835 112.065 138.645 ;
        RECT 112.075 137.835 113.445 138.645 ;
      LAYER nwell ;
        RECT 22.640 134.615 113.640 137.445 ;
      LAYER pwell ;
        RECT 22.835 133.415 24.205 134.225 ;
        RECT 24.225 133.415 25.575 134.325 ;
        RECT 25.595 133.415 26.965 134.195 ;
        RECT 26.985 133.415 28.335 134.325 ;
        RECT 28.355 134.095 29.285 134.325 ;
        RECT 34.555 134.235 35.505 134.325 ;
        RECT 28.355 133.415 32.255 134.095 ;
        RECT 33.575 133.415 35.505 134.235 ;
        RECT 35.725 133.500 36.155 134.285 ;
        RECT 37.535 134.095 38.455 134.315 ;
        RECT 44.535 134.215 45.455 134.325 ;
        RECT 43.120 134.095 45.455 134.215 ;
        RECT 47.640 134.125 48.585 134.325 ;
        RECT 36.175 133.415 45.455 134.095 ;
        RECT 45.835 133.445 48.585 134.125 ;
        RECT 22.975 133.205 23.145 133.415 ;
        RECT 25.275 133.225 25.445 133.415 ;
        RECT 25.735 133.225 25.905 133.415 ;
        RECT 27.115 133.225 27.285 133.415 ;
        RECT 28.770 133.225 28.940 133.415 ;
        RECT 33.575 133.395 33.725 133.415 ;
        RECT 33.095 133.260 33.255 133.370 ;
        RECT 33.555 133.205 33.725 133.395 ;
        RECT 34.070 133.255 34.190 133.365 ;
        RECT 36.315 133.225 36.485 133.415 ;
        RECT 37.880 133.205 38.050 133.395 ;
        RECT 38.890 133.205 39.060 133.395 ;
        RECT 43.030 133.205 43.200 133.395 ;
        RECT 45.980 133.225 46.150 133.445 ;
        RECT 47.640 133.415 48.585 133.445 ;
        RECT 48.790 133.415 52.265 134.325 ;
        RECT 52.370 133.415 56.240 134.325 ;
        RECT 56.415 133.415 59.890 134.325 ;
        RECT 60.105 133.415 61.455 134.325 ;
        RECT 61.485 133.500 61.915 134.285 ;
        RECT 62.305 134.215 63.225 134.325 ;
        RECT 62.305 134.095 64.640 134.215 ;
        RECT 69.305 134.095 70.225 134.315 ;
        RECT 75.645 134.215 76.565 134.325 ;
        RECT 75.645 134.095 77.980 134.215 ;
        RECT 82.645 134.095 83.565 134.315 ;
        RECT 62.305 133.415 71.585 134.095 ;
        RECT 72.435 133.415 74.860 134.095 ;
        RECT 75.645 133.415 84.925 134.095 ;
        RECT 85.865 133.415 87.215 134.325 ;
        RECT 87.245 133.500 87.675 134.285 ;
        RECT 88.625 133.415 89.975 134.325 ;
        RECT 92.205 134.215 93.125 134.325 ;
        RECT 89.995 133.415 91.365 134.195 ;
        RECT 92.205 134.095 94.540 134.215 ;
        RECT 99.205 134.095 100.125 134.315 ;
        RECT 102.325 134.215 103.245 134.325 ;
        RECT 102.325 134.095 104.660 134.215 ;
        RECT 109.325 134.095 110.245 134.315 ;
        RECT 92.205 133.415 101.485 134.095 ;
        RECT 102.325 133.415 111.605 134.095 ;
        RECT 112.075 133.415 113.445 134.225 ;
        RECT 51.950 133.395 52.120 133.415 ;
        RECT 56.095 133.395 56.240 133.415 ;
        RECT 46.895 133.205 47.065 133.395 ;
        RECT 48.330 133.255 48.450 133.365 ;
        RECT 22.835 132.395 24.205 133.205 ;
        RECT 24.585 132.525 33.865 133.205 ;
        RECT 34.565 132.525 38.465 133.205 ;
        RECT 24.585 132.405 26.920 132.525 ;
        RECT 24.585 132.295 25.505 132.405 ;
        RECT 31.585 132.305 32.505 132.525 ;
        RECT 37.535 132.295 38.465 132.525 ;
        RECT 38.475 132.525 42.375 133.205 ;
        RECT 42.615 132.525 46.515 133.205 ;
        RECT 38.475 132.295 39.405 132.525 ;
        RECT 42.615 132.295 43.545 132.525 ;
        RECT 46.765 132.295 48.115 133.205 ;
        RECT 49.055 133.175 50.000 133.205 ;
        RECT 51.490 133.175 51.660 133.395 ;
        RECT 51.950 133.225 52.125 133.395 ;
        RECT 56.095 133.225 56.265 133.395 ;
        RECT 56.560 133.225 56.730 133.415 ;
        RECT 51.955 133.205 52.125 133.225 ;
        RECT 56.740 133.205 56.910 133.395 ;
        RECT 60.235 133.225 60.405 133.415 ;
        RECT 60.880 133.205 61.050 133.395 ;
        RECT 61.670 133.255 61.790 133.365 ;
        RECT 65.480 133.205 65.650 133.395 ;
        RECT 66.270 133.255 66.390 133.365 ;
        RECT 66.675 133.205 66.845 133.395 ;
        RECT 68.055 133.225 68.225 133.395 ;
        RECT 71.275 133.225 71.445 133.415 ;
        RECT 71.790 133.255 71.910 133.365 ;
        RECT 68.075 133.205 68.225 133.225 ;
        RECT 73.760 133.205 73.930 133.395 ;
        RECT 74.955 133.365 75.125 133.395 ;
        RECT 74.955 133.255 75.130 133.365 ;
        RECT 74.955 133.225 75.125 133.255 ;
        RECT 78.820 133.205 78.990 133.395 ;
        RECT 80.475 133.205 80.645 133.395 ;
        RECT 80.935 133.205 81.105 133.395 ;
        RECT 83.235 133.205 83.405 133.395 ;
        RECT 83.695 133.205 83.865 133.395 ;
        RECT 84.615 133.225 84.785 133.415 ;
        RECT 85.535 133.260 85.695 133.370 ;
        RECT 85.995 133.225 86.165 133.415 ;
        RECT 88.295 133.260 88.455 133.370 ;
        RECT 88.755 133.225 88.925 133.415 ;
        RECT 91.055 133.225 91.225 133.415 ;
        RECT 91.570 133.255 91.690 133.365 ;
        RECT 94.275 133.205 94.445 133.395 ;
        RECT 94.735 133.205 94.905 133.395 ;
        RECT 99.520 133.205 99.690 133.395 ;
        RECT 101.175 133.225 101.345 133.415 ;
        RECT 101.690 133.255 101.810 133.365 ;
        RECT 109.915 133.205 110.085 133.395 ;
        RECT 111.295 133.225 111.465 133.415 ;
        RECT 111.755 133.365 111.925 133.395 ;
        RECT 111.755 133.255 111.930 133.365 ;
        RECT 111.755 133.205 111.925 133.255 ;
        RECT 113.135 133.205 113.305 133.415 ;
        RECT 48.605 132.335 49.035 133.120 ;
        RECT 49.055 132.495 51.805 133.175 ;
        RECT 49.055 132.295 50.000 132.495 ;
        RECT 51.815 132.425 53.185 133.205 ;
        RECT 53.425 132.525 57.325 133.205 ;
        RECT 57.565 132.525 61.465 133.205 ;
        RECT 62.165 132.525 66.065 133.205 ;
        RECT 56.395 132.295 57.325 132.525 ;
        RECT 60.535 132.295 61.465 132.525 ;
        RECT 65.135 132.295 66.065 132.525 ;
        RECT 66.535 132.425 67.905 133.205 ;
        RECT 68.075 132.385 70.005 133.205 ;
        RECT 70.445 132.525 74.345 133.205 ;
        RECT 69.055 132.295 70.005 132.385 ;
        RECT 73.415 132.295 74.345 132.525 ;
        RECT 74.365 132.335 74.795 133.120 ;
        RECT 75.505 132.525 79.405 133.205 ;
        RECT 78.475 132.295 79.405 132.525 ;
        RECT 79.415 132.425 80.785 133.205 ;
        RECT 80.795 132.425 82.165 133.205 ;
        RECT 82.175 132.395 83.545 133.205 ;
        RECT 83.565 132.295 84.915 133.205 ;
        RECT 85.305 132.525 94.585 133.205 ;
        RECT 85.305 132.405 87.640 132.525 ;
        RECT 85.305 132.295 86.225 132.405 ;
        RECT 92.305 132.305 93.225 132.525 ;
        RECT 94.605 132.295 95.955 133.205 ;
        RECT 96.205 132.525 100.105 133.205 ;
        RECT 99.175 132.295 100.105 132.525 ;
        RECT 100.125 132.335 100.555 133.120 ;
        RECT 100.945 132.525 110.225 133.205 ;
        RECT 100.945 132.405 103.280 132.525 ;
        RECT 100.945 132.295 101.865 132.405 ;
        RECT 107.945 132.305 108.865 132.525 ;
        RECT 110.235 132.395 112.065 133.205 ;
        RECT 112.075 132.395 113.445 133.205 ;
      LAYER nwell ;
        RECT 22.640 129.175 113.640 132.005 ;
      LAYER pwell ;
        RECT 22.835 127.975 24.205 128.785 ;
        RECT 26.495 128.655 27.415 128.875 ;
        RECT 33.495 128.775 34.415 128.885 ;
        RECT 32.080 128.655 34.415 128.775 ;
        RECT 25.135 127.975 34.415 128.655 ;
        RECT 35.725 128.060 36.155 128.845 ;
        RECT 37.095 127.975 38.465 128.755 ;
        RECT 40.295 128.655 41.215 128.875 ;
        RECT 47.295 128.775 48.215 128.885 ;
        RECT 45.880 128.655 48.215 128.775 ;
        RECT 38.935 127.975 48.215 128.655 ;
        RECT 49.255 128.795 50.205 128.885 ;
        RECT 49.255 127.975 51.185 128.795 ;
        RECT 52.185 128.775 53.105 128.885 ;
        RECT 52.185 128.655 54.520 128.775 ;
        RECT 59.185 128.655 60.105 128.875 ;
        RECT 52.185 127.975 61.465 128.655 ;
        RECT 61.485 128.060 61.915 128.845 ;
        RECT 62.305 128.775 63.225 128.885 ;
        RECT 62.305 128.655 64.640 128.775 ;
        RECT 69.305 128.655 70.225 128.875 ;
        RECT 71.965 128.775 72.885 128.885 ;
        RECT 71.965 128.655 74.300 128.775 ;
        RECT 78.965 128.655 79.885 128.875 ;
        RECT 62.305 127.975 71.585 128.655 ;
        RECT 71.965 127.975 81.245 128.655 ;
        RECT 81.265 127.975 82.615 128.885 ;
        RECT 86.295 128.655 87.225 128.885 ;
        RECT 83.325 127.975 87.225 128.655 ;
        RECT 87.245 128.060 87.675 128.845 ;
        RECT 87.705 127.975 89.055 128.885 ;
        RECT 89.075 127.975 90.445 128.755 ;
        RECT 94.115 128.655 95.045 128.885 ;
        RECT 91.145 127.975 95.045 128.655 ;
        RECT 95.055 127.975 96.425 128.755 ;
        RECT 96.435 127.975 98.265 128.785 ;
        RECT 98.275 127.975 99.645 128.755 ;
        RECT 102.855 128.655 103.785 128.885 ;
        RECT 99.885 127.975 103.785 128.655 ;
        RECT 103.805 127.975 105.155 128.885 ;
        RECT 105.185 127.975 106.535 128.885 ;
        RECT 106.555 127.975 107.925 128.755 ;
        RECT 108.395 127.975 112.065 128.785 ;
        RECT 112.075 127.975 113.445 128.785 ;
        RECT 22.975 127.765 23.145 127.975 ;
        RECT 24.815 127.820 24.975 127.930 ;
        RECT 25.275 127.765 25.445 127.975 ;
        RECT 25.735 127.765 25.905 127.955 ;
        RECT 27.115 127.765 27.285 127.955 ;
        RECT 28.770 127.765 28.940 127.955 ;
        RECT 35.395 127.820 35.555 127.930 ;
        RECT 36.775 127.820 36.935 127.930 ;
        RECT 38.155 127.785 38.325 127.975 ;
        RECT 38.670 127.815 38.790 127.925 ;
        RECT 39.075 127.785 39.245 127.975 ;
        RECT 51.035 127.955 51.185 127.975 ;
        RECT 41.835 127.765 42.005 127.955 ;
        RECT 42.295 127.785 42.465 127.955 ;
        RECT 42.315 127.765 42.465 127.785 ;
        RECT 46.890 127.765 47.060 127.955 ;
        RECT 47.355 127.765 47.525 127.955 ;
        RECT 48.790 127.815 48.910 127.925 ;
        RECT 51.035 127.785 51.205 127.955 ;
        RECT 51.550 127.815 51.670 127.925 ;
        RECT 58.395 127.765 58.565 127.955 ;
        RECT 59.775 127.765 59.945 127.955 ;
        RECT 60.290 127.815 60.410 127.925 ;
        RECT 61.155 127.785 61.325 127.975 ;
        RECT 61.615 127.765 61.785 127.955 ;
        RECT 63.455 127.765 63.625 127.955 ;
        RECT 63.915 127.765 64.085 127.955 ;
        RECT 65.755 127.810 65.915 127.920 ;
        RECT 66.215 127.765 66.385 127.955 ;
        RECT 69.895 127.765 70.065 127.955 ;
        RECT 70.355 127.765 70.525 127.955 ;
        RECT 71.275 127.785 71.445 127.975 ;
        RECT 71.735 127.765 71.905 127.955 ;
        RECT 74.035 127.765 74.205 127.955 ;
        RECT 80.935 127.785 81.105 127.975 ;
        RECT 82.315 127.785 82.485 127.975 ;
        RECT 82.830 127.815 82.950 127.925 ;
        RECT 84.155 127.765 84.325 127.955 ;
        RECT 86.640 127.785 86.810 127.975 ;
        RECT 87.835 127.785 88.005 127.975 ;
        RECT 89.215 127.785 89.385 127.975 ;
        RECT 90.650 127.815 90.770 127.925 ;
        RECT 93.815 127.765 93.985 127.955 ;
        RECT 94.330 127.815 94.450 127.925 ;
        RECT 94.460 127.785 94.630 127.975 ;
        RECT 96.115 127.785 96.285 127.975 ;
        RECT 97.955 127.785 98.125 127.975 ;
        RECT 98.415 127.785 98.585 127.975 ;
        RECT 99.795 127.765 99.965 127.955 ;
        RECT 103.200 127.785 103.370 127.975 ;
        RECT 103.935 127.785 104.105 127.975 ;
        RECT 105.315 127.785 105.485 127.975 ;
        RECT 105.775 127.765 105.945 127.955 ;
        RECT 106.235 127.765 106.405 127.955 ;
        RECT 106.695 127.785 106.865 127.975 ;
        RECT 111.755 127.955 111.925 127.975 ;
        RECT 108.130 127.815 108.250 127.925 ;
        RECT 108.535 127.765 108.705 127.955 ;
        RECT 109.915 127.765 110.085 127.955 ;
        RECT 110.430 127.815 110.550 127.925 ;
        RECT 111.745 127.785 111.925 127.955 ;
        RECT 111.745 127.765 111.915 127.785 ;
        RECT 113.135 127.765 113.305 127.975 ;
        RECT 22.835 126.955 24.205 127.765 ;
        RECT 24.225 126.855 25.575 127.765 ;
        RECT 25.605 126.855 26.955 127.765 ;
        RECT 26.975 126.985 28.345 127.765 ;
        RECT 28.355 127.085 32.255 127.765 ;
        RECT 32.865 127.085 42.145 127.765 ;
        RECT 28.355 126.855 29.285 127.085 ;
        RECT 32.865 126.965 35.200 127.085 ;
        RECT 32.865 126.855 33.785 126.965 ;
        RECT 39.865 126.865 40.785 127.085 ;
        RECT 42.315 126.945 44.245 127.765 ;
        RECT 43.295 126.855 44.245 126.945 ;
        RECT 44.595 126.855 47.205 127.765 ;
        RECT 47.225 126.855 48.575 127.765 ;
        RECT 48.605 126.895 49.035 127.680 ;
        RECT 49.425 127.085 58.705 127.765 ;
        RECT 49.425 126.965 51.760 127.085 ;
        RECT 49.425 126.855 50.345 126.965 ;
        RECT 56.425 126.865 57.345 127.085 ;
        RECT 58.725 126.855 60.075 127.765 ;
        RECT 60.555 126.985 61.925 127.765 ;
        RECT 61.935 126.955 63.765 127.765 ;
        RECT 63.785 126.855 65.135 127.765 ;
        RECT 66.075 126.985 67.445 127.765 ;
        RECT 67.455 126.955 70.205 127.765 ;
        RECT 70.225 126.855 71.575 127.765 ;
        RECT 71.605 126.855 72.955 127.765 ;
        RECT 72.975 126.955 74.345 127.765 ;
        RECT 74.365 126.895 74.795 127.680 ;
        RECT 75.185 127.085 84.465 127.765 ;
        RECT 84.845 127.085 94.125 127.765 ;
        RECT 75.185 126.965 77.520 127.085 ;
        RECT 75.185 126.855 76.105 126.965 ;
        RECT 82.185 126.865 83.105 127.085 ;
        RECT 84.845 126.965 87.180 127.085 ;
        RECT 84.845 126.855 85.765 126.965 ;
        RECT 91.845 126.865 92.765 127.085 ;
        RECT 94.595 126.955 100.105 127.765 ;
        RECT 100.125 126.895 100.555 127.680 ;
        RECT 100.575 126.955 106.085 127.765 ;
        RECT 106.105 126.855 107.455 127.765 ;
        RECT 107.475 126.955 108.845 127.765 ;
        RECT 108.855 126.985 110.225 127.765 ;
        RECT 110.695 126.985 112.065 127.765 ;
        RECT 112.075 126.955 113.445 127.765 ;
      LAYER nwell ;
        RECT 22.640 123.735 113.640 126.565 ;
      LAYER pwell ;
        RECT 22.835 122.535 24.205 123.345 ;
        RECT 24.415 123.215 26.625 123.445 ;
        RECT 29.345 123.215 30.275 123.435 ;
        RECT 24.415 122.535 34.785 123.215 ;
        RECT 35.725 122.620 36.155 123.405 ;
        RECT 41.455 123.355 42.405 123.445 ;
        RECT 37.095 122.535 38.465 123.315 ;
        RECT 38.475 122.535 39.845 123.315 ;
        RECT 40.475 122.535 42.405 123.355 ;
        RECT 42.815 123.215 45.025 123.445 ;
        RECT 47.745 123.215 48.675 123.435 ;
        RECT 42.815 122.535 53.185 123.215 ;
        RECT 53.195 122.535 55.945 123.345 ;
        RECT 55.955 122.535 57.325 123.315 ;
        RECT 57.335 122.535 58.705 123.345 ;
        RECT 58.715 122.535 60.085 123.315 ;
        RECT 60.095 122.535 61.465 123.345 ;
        RECT 61.485 122.620 61.915 123.405 ;
        RECT 61.935 122.535 63.765 123.345 ;
        RECT 63.775 122.535 65.145 123.315 ;
        RECT 65.615 122.535 69.285 123.345 ;
        RECT 69.295 122.535 74.805 123.345 ;
        RECT 74.815 122.535 76.185 123.315 ;
        RECT 76.195 122.535 78.805 123.445 ;
        RECT 78.955 122.535 80.325 123.315 ;
        RECT 80.335 122.535 81.705 123.345 ;
        RECT 81.715 122.535 87.225 123.345 ;
        RECT 87.245 122.620 87.675 123.405 ;
        RECT 87.695 122.535 89.065 123.345 ;
        RECT 89.075 122.535 92.745 123.345 ;
        RECT 92.755 122.535 94.125 123.315 ;
        RECT 95.055 122.535 96.425 123.315 ;
        RECT 96.435 122.535 97.805 123.315 ;
        RECT 97.815 122.535 99.185 123.315 ;
        RECT 100.125 122.535 101.475 123.445 ;
        RECT 106.005 123.215 106.935 123.435 ;
        RECT 109.655 123.215 111.865 123.445 ;
        RECT 101.495 122.535 111.865 123.215 ;
        RECT 112.075 122.535 113.445 123.345 ;
        RECT 22.975 122.325 23.145 122.535 ;
        RECT 24.355 122.325 24.525 122.515 ;
        RECT 26.655 122.325 26.825 122.515 ;
        RECT 27.170 122.375 27.290 122.485 ;
        RECT 34.475 122.345 34.645 122.535 ;
        RECT 35.395 122.380 35.555 122.490 ;
        RECT 36.775 122.380 36.935 122.490 ;
        RECT 37.235 122.345 37.405 122.535 ;
        RECT 37.695 122.325 37.865 122.515 ;
        RECT 38.615 122.345 38.785 122.535 ;
        RECT 40.475 122.515 40.625 122.535 ;
        RECT 40.050 122.375 40.170 122.485 ;
        RECT 40.455 122.345 40.625 122.515 ;
        RECT 48.275 122.325 48.445 122.515 ;
        RECT 49.655 122.370 49.815 122.480 ;
        RECT 50.115 122.325 50.285 122.515 ;
        RECT 51.550 122.375 51.670 122.485 ;
        RECT 52.875 122.325 53.045 122.535 ;
        RECT 55.635 122.515 55.805 122.535 ;
        RECT 53.795 122.370 53.955 122.480 ;
        RECT 55.175 122.325 55.345 122.515 ;
        RECT 55.635 122.345 55.810 122.515 ;
        RECT 57.015 122.345 57.185 122.535 ;
        RECT 58.395 122.345 58.565 122.535 ;
        RECT 58.855 122.345 59.025 122.535 ;
        RECT 61.155 122.345 61.325 122.535 ;
        RECT 63.455 122.345 63.625 122.535 ;
        RECT 63.915 122.345 64.085 122.535 ;
        RECT 65.350 122.375 65.470 122.485 ;
        RECT 55.640 122.325 55.810 122.345 ;
        RECT 68.515 122.325 68.685 122.515 ;
        RECT 68.975 122.325 69.145 122.535 ;
        RECT 70.355 122.325 70.525 122.515 ;
        RECT 71.735 122.325 71.905 122.515 ;
        RECT 74.035 122.325 74.205 122.515 ;
        RECT 74.495 122.345 74.665 122.535 ;
        RECT 74.955 122.345 75.125 122.535 ;
        RECT 76.340 122.345 76.510 122.535 ;
        RECT 79.095 122.345 79.265 122.535 ;
        RECT 81.395 122.345 81.565 122.535 ;
        RECT 85.075 122.325 85.245 122.515 ;
        RECT 85.995 122.370 86.155 122.480 ;
        RECT 86.455 122.325 86.625 122.515 ;
        RECT 86.915 122.345 87.085 122.535 ;
        RECT 88.755 122.345 88.925 122.535 ;
        RECT 92.435 122.345 92.605 122.535 ;
        RECT 92.895 122.345 93.065 122.535 ;
        RECT 94.735 122.380 94.895 122.490 ;
        RECT 95.195 122.345 95.365 122.535 ;
        RECT 96.575 122.345 96.745 122.535 ;
        RECT 97.955 122.325 98.125 122.535 ;
        RECT 99.335 122.325 99.505 122.515 ;
        RECT 99.795 122.485 99.955 122.490 ;
        RECT 99.795 122.380 99.970 122.485 ;
        RECT 99.850 122.375 99.970 122.380 ;
        RECT 100.255 122.345 100.425 122.535 ;
        RECT 101.175 122.370 101.335 122.480 ;
        RECT 101.635 122.325 101.805 122.535 ;
        RECT 113.135 122.325 113.305 122.535 ;
        RECT 22.835 121.515 24.205 122.325 ;
        RECT 24.215 121.545 25.585 122.325 ;
        RECT 25.605 121.415 26.955 122.325 ;
        RECT 27.635 121.645 38.005 122.325 ;
        RECT 38.215 121.645 48.585 122.325 ;
        RECT 27.635 121.415 29.845 121.645 ;
        RECT 32.565 121.425 33.495 121.645 ;
        RECT 38.215 121.415 40.425 121.645 ;
        RECT 43.145 121.425 44.075 121.645 ;
        RECT 48.605 121.455 49.035 122.240 ;
        RECT 49.975 121.545 51.345 122.325 ;
        RECT 51.825 121.415 53.175 122.325 ;
        RECT 54.115 121.545 55.485 122.325 ;
        RECT 55.495 121.415 58.105 122.325 ;
        RECT 58.455 121.645 68.825 122.325 ;
        RECT 58.455 121.415 60.665 121.645 ;
        RECT 63.385 121.425 64.315 121.645 ;
        RECT 68.835 121.545 70.205 122.325 ;
        RECT 70.215 121.545 71.585 122.325 ;
        RECT 71.595 121.545 72.965 122.325 ;
        RECT 72.985 121.415 74.335 122.325 ;
        RECT 74.365 121.455 74.795 122.240 ;
        RECT 75.015 121.645 85.385 122.325 ;
        RECT 75.015 121.415 77.225 121.645 ;
        RECT 79.945 121.425 80.875 121.645 ;
        RECT 86.315 121.545 87.685 122.325 ;
        RECT 87.895 121.645 98.265 122.325 ;
        RECT 87.895 121.415 90.105 121.645 ;
        RECT 92.825 121.425 93.755 121.645 ;
        RECT 98.275 121.545 99.645 122.325 ;
        RECT 100.125 121.455 100.555 122.240 ;
        RECT 101.495 121.645 111.865 122.325 ;
        RECT 106.005 121.425 106.935 121.645 ;
        RECT 109.655 121.415 111.865 121.645 ;
        RECT 112.075 121.515 113.445 122.325 ;
      LAYER nwell ;
        RECT 22.640 118.295 113.640 121.125 ;
      LAYER pwell ;
        RECT 22.835 117.095 24.205 117.905 ;
        RECT 29.645 117.775 30.575 117.995 ;
        RECT 33.295 117.775 35.505 118.005 ;
        RECT 25.135 117.095 35.505 117.775 ;
        RECT 35.725 117.180 36.155 117.965 ;
        RECT 36.185 117.095 37.535 118.005 ;
        RECT 37.555 117.095 38.925 117.875 ;
        RECT 38.935 117.095 40.305 117.875 ;
        RECT 44.825 117.775 45.755 117.995 ;
        RECT 48.475 117.775 50.685 118.005 ;
        RECT 40.315 117.095 50.685 117.775 ;
        RECT 51.095 117.775 53.305 118.005 ;
        RECT 56.025 117.775 56.955 117.995 ;
        RECT 51.095 117.095 61.465 117.775 ;
        RECT 61.485 117.180 61.915 117.965 ;
        RECT 62.135 117.775 64.345 118.005 ;
        RECT 67.065 117.775 67.995 117.995 ;
        RECT 72.715 117.775 74.925 118.005 ;
        RECT 77.645 117.775 78.575 117.995 ;
        RECT 62.135 117.095 72.505 117.775 ;
        RECT 72.715 117.095 83.085 117.775 ;
        RECT 83.105 117.095 84.455 118.005 ;
        RECT 84.485 117.095 85.835 118.005 ;
        RECT 85.865 117.095 87.215 118.005 ;
        RECT 87.245 117.180 87.675 117.965 ;
        RECT 87.895 117.775 90.105 118.005 ;
        RECT 92.825 117.775 93.755 117.995 ;
        RECT 102.785 117.775 103.715 117.995 ;
        RECT 106.435 117.775 108.645 118.005 ;
        RECT 87.895 117.095 98.265 117.775 ;
        RECT 98.275 117.095 108.645 117.775 ;
        RECT 108.865 117.095 110.215 118.005 ;
        RECT 110.245 117.095 111.595 118.005 ;
        RECT 112.075 117.095 113.445 117.905 ;
        RECT 22.975 116.885 23.145 117.095 ;
        RECT 24.815 116.940 24.975 117.050 ;
        RECT 25.275 116.905 25.445 117.095 ;
        RECT 34.475 116.885 34.645 117.075 ;
        RECT 35.395 116.930 35.555 117.040 ;
        RECT 36.315 116.905 36.485 117.095 ;
        RECT 37.235 116.885 37.405 117.075 ;
        RECT 38.615 116.885 38.785 117.095 ;
        RECT 39.995 116.885 40.165 117.095 ;
        RECT 40.455 116.905 40.625 117.095 ;
        RECT 41.375 116.885 41.545 117.075 ;
        RECT 44.135 116.885 44.305 117.075 ;
        RECT 44.595 116.885 44.765 117.075 ;
        RECT 45.975 116.885 46.145 117.075 ;
        RECT 48.275 116.885 48.445 117.075 ;
        RECT 51.495 116.885 51.665 117.075 ;
        RECT 57.015 116.885 57.185 117.075 ;
        RECT 58.395 116.885 58.565 117.075 ;
        RECT 61.155 116.885 61.325 117.095 ;
        RECT 62.075 116.885 62.245 117.075 ;
        RECT 63.510 116.935 63.630 117.045 ;
        RECT 63.915 116.885 64.085 117.075 ;
        RECT 65.350 116.935 65.470 117.045 ;
        RECT 67.135 116.885 67.305 117.075 ;
        RECT 72.195 116.905 72.365 117.095 ;
        RECT 72.655 116.885 72.825 117.075 ;
        RECT 74.035 116.885 74.205 117.075 ;
        RECT 75.010 116.935 75.130 117.045 ;
        RECT 75.415 116.885 75.585 117.075 ;
        RECT 76.795 116.885 76.965 117.075 ;
        RECT 82.775 116.905 82.945 117.095 ;
        RECT 84.155 116.905 84.325 117.095 ;
        RECT 84.615 116.905 84.785 117.095 ;
        RECT 85.995 116.905 86.165 117.095 ;
        RECT 87.890 116.935 88.010 117.045 ;
        RECT 88.295 116.885 88.465 117.075 ;
        RECT 97.955 116.905 98.125 117.095 ;
        RECT 98.415 116.905 98.585 117.095 ;
        RECT 99.795 116.885 99.965 117.075 ;
        RECT 101.175 116.930 101.335 117.040 ;
        RECT 101.635 116.885 101.805 117.075 ;
        RECT 109.915 116.905 110.085 117.095 ;
        RECT 110.375 116.905 110.545 117.095 ;
        RECT 111.810 116.935 111.930 117.045 ;
        RECT 113.135 116.885 113.305 117.095 ;
        RECT 22.835 116.075 24.205 116.885 ;
        RECT 24.415 116.205 34.785 116.885 ;
        RECT 24.415 115.975 26.625 116.205 ;
        RECT 29.345 115.985 30.275 116.205 ;
        RECT 35.725 116.015 36.155 116.800 ;
        RECT 36.185 115.975 37.535 116.885 ;
        RECT 37.555 116.105 38.925 116.885 ;
        RECT 38.945 115.975 40.295 116.885 ;
        RECT 40.325 115.975 41.675 116.885 ;
        RECT 41.695 116.075 44.445 116.885 ;
        RECT 44.465 115.975 45.815 116.885 ;
        RECT 45.835 116.105 47.205 116.885 ;
        RECT 47.215 116.075 48.585 116.885 ;
        RECT 48.605 116.015 49.035 116.800 ;
        RECT 49.055 116.075 51.805 116.885 ;
        RECT 51.815 116.075 57.325 116.885 ;
        RECT 57.345 115.975 58.695 116.885 ;
        RECT 58.715 116.075 61.465 116.885 ;
        RECT 61.485 116.015 61.915 116.800 ;
        RECT 61.945 115.975 63.295 116.885 ;
        RECT 63.785 115.975 65.135 116.885 ;
        RECT 65.615 116.075 67.445 116.885 ;
        RECT 67.455 116.075 72.965 116.885 ;
        RECT 72.985 115.975 74.335 116.885 ;
        RECT 74.365 116.015 74.795 116.800 ;
        RECT 75.285 115.975 76.635 116.885 ;
        RECT 76.655 116.205 87.025 116.885 ;
        RECT 81.165 115.985 82.095 116.205 ;
        RECT 84.815 115.975 87.025 116.205 ;
        RECT 87.245 116.015 87.675 116.800 ;
        RECT 88.165 115.975 89.515 116.885 ;
        RECT 89.735 116.205 100.105 116.885 ;
        RECT 89.735 115.975 91.945 116.205 ;
        RECT 94.665 115.985 95.595 116.205 ;
        RECT 100.125 116.015 100.555 116.800 ;
        RECT 101.495 116.205 111.865 116.885 ;
        RECT 106.005 115.985 106.935 116.205 ;
        RECT 109.655 115.975 111.865 116.205 ;
        RECT 112.075 116.075 113.445 116.885 ;
      LAYER nwell ;
        RECT 22.640 114.080 113.640 115.685 ;
        RECT 20.485 54.580 29.875 66.420 ;
        RECT 31.685 54.590 41.075 66.430 ;
        RECT 42.905 54.560 52.295 66.400 ;
        RECT 54.155 54.540 63.545 66.380 ;
        RECT 65.375 54.530 74.765 66.370 ;
        RECT 76.615 54.520 86.005 66.360 ;
        RECT 87.865 54.530 97.255 66.370 ;
        RECT 99.145 54.520 108.535 66.360 ;
        RECT 110.415 54.520 119.805 66.360 ;
        RECT 121.665 54.520 131.055 66.360 ;
        RECT 132.415 54.490 139.375 66.330 ;
        RECT 20.655 49.020 23.115 53.210 ;
      LAYER pwell ;
        RECT 20.555 45.340 22.915 48.340 ;
      LAYER nwell ;
        RECT 24.735 45.940 29.125 53.130 ;
        RECT 31.855 49.030 34.315 53.220 ;
      LAYER pwell ;
        RECT 31.755 45.350 34.115 48.350 ;
      LAYER nwell ;
        RECT 35.935 45.950 40.325 53.140 ;
        RECT 43.075 49.000 45.535 53.190 ;
      LAYER pwell ;
        RECT 42.975 45.320 45.335 48.320 ;
      LAYER nwell ;
        RECT 47.155 45.920 51.545 53.110 ;
        RECT 54.325 48.980 56.785 53.170 ;
      LAYER pwell ;
        RECT 54.225 45.300 56.585 48.300 ;
      LAYER nwell ;
        RECT 58.405 45.900 62.795 53.090 ;
        RECT 65.545 48.970 68.005 53.160 ;
      LAYER pwell ;
        RECT 65.445 45.290 67.805 48.290 ;
      LAYER nwell ;
        RECT 69.625 45.890 74.015 53.080 ;
        RECT 76.785 48.960 79.245 53.150 ;
      LAYER pwell ;
        RECT 76.685 45.280 79.045 48.280 ;
      LAYER nwell ;
        RECT 80.865 45.880 85.255 53.070 ;
        RECT 88.035 48.970 90.495 53.160 ;
      LAYER pwell ;
        RECT 87.935 45.290 90.295 48.290 ;
      LAYER nwell ;
        RECT 92.115 45.890 96.505 53.080 ;
        RECT 99.315 48.960 101.775 53.150 ;
      LAYER pwell ;
        RECT 99.215 45.280 101.575 48.280 ;
      LAYER nwell ;
        RECT 103.395 45.880 107.785 53.070 ;
        RECT 110.585 48.960 113.045 53.150 ;
      LAYER pwell ;
        RECT 110.485 45.280 112.845 48.280 ;
      LAYER nwell ;
        RECT 114.665 45.880 119.055 53.070 ;
        RECT 121.835 48.960 124.295 53.150 ;
      LAYER pwell ;
        RECT 121.735 45.280 124.095 48.280 ;
      LAYER nwell ;
        RECT 125.915 45.880 130.305 53.070 ;
        RECT 19.615 32.280 24.005 39.470 ;
      LAYER pwell ;
        RECT 25.825 37.070 28.185 40.070 ;
      LAYER nwell ;
        RECT 25.625 32.200 28.085 36.390 ;
        RECT 30.895 32.280 35.285 39.470 ;
      LAYER pwell ;
        RECT 37.105 37.070 39.465 40.070 ;
      LAYER nwell ;
        RECT 36.905 32.200 39.365 36.390 ;
        RECT 42.185 32.260 46.575 39.450 ;
      LAYER pwell ;
        RECT 48.395 37.050 50.755 40.050 ;
      LAYER nwell ;
        RECT 48.195 32.180 50.655 36.370 ;
        RECT 53.405 32.260 57.795 39.450 ;
      LAYER pwell ;
        RECT 59.615 37.050 61.975 40.050 ;
      LAYER nwell ;
        RECT 59.415 32.180 61.875 36.370 ;
        RECT 64.605 32.260 68.995 39.450 ;
      LAYER pwell ;
        RECT 70.815 37.050 73.175 40.050 ;
      LAYER nwell ;
        RECT 70.615 32.180 73.075 36.370 ;
        RECT 75.895 32.250 80.285 39.440 ;
      LAYER pwell ;
        RECT 82.105 37.040 84.465 40.040 ;
      LAYER nwell ;
        RECT 81.905 32.170 84.365 36.360 ;
        RECT 87.135 32.270 91.525 39.460 ;
      LAYER pwell ;
        RECT 93.345 37.060 95.705 40.060 ;
      LAYER nwell ;
        RECT 93.145 32.190 95.605 36.380 ;
        RECT 98.345 32.290 102.735 39.480 ;
      LAYER pwell ;
        RECT 104.555 37.080 106.915 40.080 ;
      LAYER nwell ;
        RECT 104.355 32.210 106.815 36.400 ;
        RECT 109.545 32.330 113.935 39.520 ;
      LAYER pwell ;
        RECT 115.755 37.120 118.115 40.120 ;
      LAYER nwell ;
        RECT 115.555 32.250 118.015 36.440 ;
        RECT 120.755 32.350 125.145 39.540 ;
      LAYER pwell ;
        RECT 126.965 37.140 129.325 40.140 ;
      LAYER nwell ;
        RECT 126.765 32.270 129.225 36.460 ;
        RECT 18.865 18.990 28.255 30.830 ;
        RECT 30.145 18.990 39.535 30.830 ;
        RECT 41.435 18.970 50.825 30.810 ;
        RECT 52.655 18.970 62.045 30.810 ;
        RECT 63.855 18.970 73.245 30.810 ;
        RECT 75.145 18.960 84.535 30.800 ;
        RECT 86.385 18.980 95.775 30.820 ;
        RECT 97.595 19.000 106.985 30.840 ;
        RECT 108.795 19.040 118.185 30.880 ;
        RECT 120.005 19.060 129.395 30.900 ;
        RECT 131.725 19.030 138.685 30.870 ;
      LAYER li1 ;
        RECT 22.830 203.945 113.450 204.115 ;
        RECT 22.915 203.195 24.125 203.945 ;
        RECT 24.760 203.400 30.105 203.945 ;
        RECT 30.280 203.400 35.625 203.945 ;
        RECT 22.915 202.655 23.435 203.195 ;
        RECT 23.605 202.485 24.125 203.025 ;
        RECT 22.915 201.395 24.125 202.485 ;
        RECT 26.350 201.830 26.700 203.080 ;
        RECT 28.180 202.570 28.520 203.400 ;
        RECT 31.870 201.830 32.220 203.080 ;
        RECT 33.700 202.570 34.040 203.400 ;
        RECT 35.795 203.220 36.085 203.945 ;
        RECT 36.255 203.195 37.465 203.945 ;
        RECT 37.640 203.400 42.985 203.945 ;
        RECT 43.160 203.400 48.505 203.945 ;
        RECT 24.760 201.395 30.105 201.830 ;
        RECT 30.280 201.395 35.625 201.830 ;
        RECT 35.795 201.395 36.085 202.560 ;
        RECT 36.255 202.485 36.775 203.025 ;
        RECT 36.945 202.655 37.465 203.195 ;
        RECT 36.255 201.395 37.465 202.485 ;
        RECT 39.230 201.830 39.580 203.080 ;
        RECT 41.060 202.570 41.400 203.400 ;
        RECT 44.750 201.830 45.100 203.080 ;
        RECT 46.580 202.570 46.920 203.400 ;
        RECT 48.675 203.220 48.965 203.945 ;
        RECT 49.595 203.175 53.105 203.945 ;
        RECT 53.280 203.400 58.625 203.945 ;
        RECT 37.640 201.395 42.985 201.830 ;
        RECT 43.160 201.395 48.505 201.830 ;
        RECT 48.675 201.395 48.965 202.560 ;
        RECT 49.595 202.485 51.285 203.005 ;
        RECT 51.455 202.655 53.105 203.175 ;
        RECT 49.595 201.395 53.105 202.485 ;
        RECT 54.870 201.830 55.220 203.080 ;
        RECT 56.700 202.570 57.040 203.400 ;
        RECT 58.855 203.125 59.065 203.945 ;
        RECT 59.235 203.145 59.565 203.775 ;
        RECT 59.235 202.545 59.485 203.145 ;
        RECT 59.735 203.125 59.965 203.945 ;
        RECT 60.175 203.270 60.435 203.775 ;
        RECT 60.615 203.565 60.945 203.945 ;
        RECT 61.125 203.395 61.295 203.775 ;
        RECT 59.655 202.705 59.985 202.955 ;
        RECT 53.280 201.395 58.625 201.830 ;
        RECT 58.855 201.395 59.065 202.535 ;
        RECT 59.235 201.565 59.565 202.545 ;
        RECT 59.735 201.395 59.965 202.535 ;
        RECT 60.175 202.470 60.345 203.270 ;
        RECT 60.630 203.225 61.295 203.395 ;
        RECT 60.630 202.970 60.800 203.225 ;
        RECT 61.555 203.220 61.845 203.945 ;
        RECT 62.475 203.295 62.735 203.775 ;
        RECT 62.905 203.405 63.155 203.945 ;
        RECT 60.515 202.640 60.800 202.970 ;
        RECT 61.035 202.675 61.365 203.045 ;
        RECT 60.630 202.495 60.800 202.640 ;
        RECT 60.175 201.565 60.445 202.470 ;
        RECT 60.630 202.325 61.295 202.495 ;
        RECT 60.615 201.395 60.945 202.155 ;
        RECT 61.125 201.565 61.295 202.325 ;
        RECT 61.555 201.395 61.845 202.560 ;
        RECT 62.475 202.265 62.645 203.295 ;
        RECT 63.325 203.240 63.545 203.725 ;
        RECT 62.815 202.645 63.045 203.040 ;
        RECT 63.215 202.815 63.545 203.240 ;
        RECT 63.715 203.565 64.605 203.735 ;
        RECT 63.715 202.840 63.885 203.565 ;
        RECT 64.055 203.010 64.605 203.395 ;
        RECT 64.785 203.220 65.115 203.730 ;
        RECT 65.285 203.545 65.615 203.945 ;
        RECT 66.665 203.375 66.995 203.715 ;
        RECT 67.165 203.545 67.495 203.945 ;
        RECT 63.715 202.770 64.605 202.840 ;
        RECT 63.710 202.745 64.605 202.770 ;
        RECT 63.700 202.730 64.605 202.745 ;
        RECT 63.695 202.715 64.605 202.730 ;
        RECT 63.685 202.710 64.605 202.715 ;
        RECT 63.680 202.700 64.605 202.710 ;
        RECT 63.675 202.690 64.605 202.700 ;
        RECT 63.665 202.685 64.605 202.690 ;
        RECT 63.655 202.675 64.605 202.685 ;
        RECT 63.645 202.670 64.605 202.675 ;
        RECT 63.645 202.665 63.980 202.670 ;
        RECT 63.630 202.660 63.980 202.665 ;
        RECT 63.615 202.650 63.980 202.660 ;
        RECT 63.590 202.645 63.980 202.650 ;
        RECT 62.815 202.640 63.980 202.645 ;
        RECT 62.815 202.605 63.950 202.640 ;
        RECT 62.815 202.580 63.915 202.605 ;
        RECT 62.815 202.550 63.885 202.580 ;
        RECT 62.815 202.520 63.865 202.550 ;
        RECT 62.815 202.490 63.845 202.520 ;
        RECT 62.815 202.480 63.775 202.490 ;
        RECT 62.815 202.470 63.750 202.480 ;
        RECT 62.815 202.455 63.730 202.470 ;
        RECT 62.815 202.440 63.710 202.455 ;
        RECT 62.920 202.430 63.705 202.440 ;
        RECT 62.920 202.395 63.690 202.430 ;
        RECT 62.475 201.565 62.750 202.265 ;
        RECT 62.920 202.145 63.675 202.395 ;
        RECT 63.845 202.075 64.175 202.320 ;
        RECT 64.345 202.220 64.605 202.670 ;
        RECT 64.785 202.455 64.975 203.220 ;
        RECT 65.285 203.205 67.650 203.375 ;
        RECT 65.285 203.035 65.455 203.205 ;
        RECT 65.145 202.705 65.455 203.035 ;
        RECT 65.625 202.705 65.930 203.035 ;
        RECT 63.990 202.050 64.175 202.075 ;
        RECT 63.990 201.950 64.605 202.050 ;
        RECT 62.920 201.395 63.175 201.940 ;
        RECT 63.345 201.565 63.825 201.905 ;
        RECT 64.000 201.395 64.605 201.950 ;
        RECT 64.785 201.605 65.115 202.455 ;
        RECT 65.285 201.395 65.535 202.535 ;
        RECT 65.715 202.375 65.930 202.705 ;
        RECT 66.105 202.375 66.390 203.035 ;
        RECT 66.585 202.375 66.850 203.035 ;
        RECT 67.065 202.375 67.310 203.035 ;
        RECT 67.480 202.205 67.650 203.205 ;
        RECT 65.725 202.035 67.015 202.205 ;
        RECT 65.725 201.615 65.975 202.035 ;
        RECT 66.205 201.395 66.535 201.865 ;
        RECT 66.765 201.615 67.015 202.035 ;
        RECT 67.195 202.035 67.650 202.205 ;
        RECT 67.995 203.270 68.270 203.615 ;
        RECT 68.460 203.545 68.835 203.945 ;
        RECT 69.005 203.375 69.175 203.725 ;
        RECT 69.345 203.545 69.675 203.945 ;
        RECT 69.845 203.375 70.105 203.775 ;
        RECT 67.995 202.535 68.165 203.270 ;
        RECT 68.440 203.205 70.105 203.375 ;
        RECT 68.440 203.035 68.610 203.205 ;
        RECT 70.285 203.125 70.615 203.545 ;
        RECT 70.785 203.125 71.045 203.945 ;
        RECT 71.220 203.205 71.555 203.945 ;
        RECT 70.285 203.035 70.535 203.125 ;
        RECT 71.725 203.035 71.940 203.730 ;
        RECT 72.130 203.205 72.480 203.730 ;
        RECT 72.650 203.205 73.345 203.775 ;
        RECT 74.435 203.220 74.725 203.945 ;
        RECT 72.275 203.035 72.480 203.205 ;
        RECT 68.335 202.705 68.610 203.035 ;
        RECT 68.780 202.705 69.605 203.035 ;
        RECT 69.820 202.705 70.535 203.035 ;
        RECT 70.705 202.705 71.040 202.955 ;
        RECT 71.240 202.705 71.525 203.035 ;
        RECT 71.725 202.705 72.105 203.035 ;
        RECT 72.275 202.705 72.585 203.035 ;
        RECT 68.440 202.535 68.610 202.705 ;
        RECT 67.195 201.605 67.525 202.035 ;
        RECT 67.995 201.565 68.270 202.535 ;
        RECT 68.440 202.365 69.100 202.535 ;
        RECT 69.360 202.415 69.605 202.705 ;
        RECT 68.930 202.245 69.100 202.365 ;
        RECT 69.775 202.245 70.105 202.535 ;
        RECT 68.480 201.395 68.760 202.195 ;
        RECT 68.930 202.075 70.105 202.245 ;
        RECT 70.365 202.145 70.535 202.705 ;
        RECT 72.755 202.535 72.925 203.205 ;
        RECT 74.955 203.125 75.165 203.945 ;
        RECT 75.335 203.145 75.665 203.775 ;
        RECT 68.930 201.575 70.545 201.905 ;
        RECT 70.785 201.395 71.045 202.535 ;
        RECT 71.215 201.395 71.475 202.535 ;
        RECT 71.645 202.365 72.925 202.535 ;
        RECT 73.105 202.365 73.345 203.035 ;
        RECT 71.645 201.565 71.975 202.365 ;
        RECT 72.145 201.395 72.315 202.195 ;
        RECT 72.515 201.565 72.845 202.365 ;
        RECT 73.045 201.395 73.325 202.195 ;
        RECT 74.435 201.395 74.725 202.560 ;
        RECT 75.335 202.545 75.585 203.145 ;
        RECT 75.835 203.125 76.065 203.945 ;
        RECT 76.335 203.125 76.545 203.945 ;
        RECT 76.715 203.145 77.045 203.775 ;
        RECT 75.755 202.705 76.085 202.955 ;
        RECT 76.715 202.545 76.965 203.145 ;
        RECT 77.215 203.125 77.445 203.945 ;
        RECT 77.745 203.395 77.915 203.775 ;
        RECT 78.095 203.565 78.425 203.945 ;
        RECT 77.745 203.225 78.410 203.395 ;
        RECT 78.605 203.270 78.865 203.775 ;
        RECT 77.135 202.705 77.465 202.955 ;
        RECT 77.675 202.675 78.005 203.045 ;
        RECT 78.240 202.970 78.410 203.225 ;
        RECT 78.240 202.640 78.525 202.970 ;
        RECT 74.955 201.395 75.165 202.535 ;
        RECT 75.335 201.565 75.665 202.545 ;
        RECT 75.835 201.395 76.065 202.535 ;
        RECT 76.335 201.395 76.545 202.535 ;
        RECT 76.715 201.565 77.045 202.545 ;
        RECT 77.215 201.395 77.445 202.535 ;
        RECT 78.240 202.495 78.410 202.640 ;
        RECT 77.745 202.325 78.410 202.495 ;
        RECT 78.695 202.470 78.865 203.270 ;
        RECT 79.035 203.175 81.625 203.945 ;
        RECT 81.800 203.400 87.145 203.945 ;
        RECT 77.745 201.565 77.915 202.325 ;
        RECT 78.095 201.395 78.425 202.155 ;
        RECT 78.595 201.565 78.865 202.470 ;
        RECT 79.035 202.485 80.245 203.005 ;
        RECT 80.415 202.655 81.625 203.175 ;
        RECT 79.035 201.395 81.625 202.485 ;
        RECT 83.390 201.830 83.740 203.080 ;
        RECT 85.220 202.570 85.560 203.400 ;
        RECT 87.315 203.220 87.605 203.945 ;
        RECT 87.775 203.175 89.445 203.945 ;
        RECT 89.620 203.400 94.965 203.945 ;
        RECT 81.800 201.395 87.145 201.830 ;
        RECT 87.315 201.395 87.605 202.560 ;
        RECT 87.775 202.485 88.525 203.005 ;
        RECT 88.695 202.655 89.445 203.175 ;
        RECT 87.775 201.395 89.445 202.485 ;
        RECT 91.210 201.830 91.560 203.080 ;
        RECT 93.040 202.570 93.380 203.400 ;
        RECT 95.195 203.125 95.405 203.945 ;
        RECT 95.575 203.145 95.905 203.775 ;
        RECT 95.575 202.545 95.825 203.145 ;
        RECT 96.075 203.125 96.305 203.945 ;
        RECT 97.525 203.395 97.695 203.775 ;
        RECT 97.875 203.565 98.205 203.945 ;
        RECT 97.525 203.225 98.190 203.395 ;
        RECT 98.385 203.270 98.645 203.775 ;
        RECT 95.995 202.705 96.325 202.955 ;
        RECT 97.455 202.675 97.785 203.045 ;
        RECT 98.020 202.970 98.190 203.225 ;
        RECT 98.020 202.640 98.305 202.970 ;
        RECT 89.620 201.395 94.965 201.830 ;
        RECT 95.195 201.395 95.405 202.535 ;
        RECT 95.575 201.565 95.905 202.545 ;
        RECT 96.075 201.395 96.305 202.535 ;
        RECT 98.020 202.495 98.190 202.640 ;
        RECT 97.525 202.325 98.190 202.495 ;
        RECT 98.475 202.470 98.645 203.270 ;
        RECT 98.855 203.125 99.085 203.945 ;
        RECT 99.255 203.145 99.585 203.775 ;
        RECT 98.835 202.705 99.165 202.955 ;
        RECT 99.335 202.545 99.585 203.145 ;
        RECT 99.755 203.125 99.965 203.945 ;
        RECT 100.195 203.220 100.485 203.945 ;
        RECT 100.715 203.125 100.925 203.945 ;
        RECT 101.095 203.145 101.425 203.775 ;
        RECT 97.525 201.565 97.695 202.325 ;
        RECT 97.875 201.395 98.205 202.155 ;
        RECT 98.375 201.565 98.645 202.470 ;
        RECT 98.855 201.395 99.085 202.535 ;
        RECT 99.255 201.565 99.585 202.545 ;
        RECT 99.755 201.395 99.965 202.535 ;
        RECT 100.195 201.395 100.485 202.560 ;
        RECT 101.095 202.545 101.345 203.145 ;
        RECT 101.595 203.125 101.825 203.945 ;
        RECT 102.610 203.315 102.895 203.775 ;
        RECT 103.065 203.485 103.335 203.945 ;
        RECT 102.610 203.145 103.565 203.315 ;
        RECT 101.515 202.705 101.845 202.955 ;
        RECT 100.715 201.395 100.925 202.535 ;
        RECT 101.095 201.565 101.425 202.545 ;
        RECT 101.595 201.395 101.825 202.535 ;
        RECT 102.495 202.415 103.185 202.975 ;
        RECT 103.355 202.245 103.565 203.145 ;
        RECT 102.610 202.025 103.565 202.245 ;
        RECT 103.735 202.975 104.135 203.775 ;
        RECT 104.325 203.315 104.605 203.775 ;
        RECT 105.125 203.485 105.450 203.945 ;
        RECT 104.325 203.145 105.450 203.315 ;
        RECT 105.620 203.205 106.005 203.775 ;
        RECT 106.640 203.400 111.985 203.945 ;
        RECT 105.000 203.035 105.450 203.145 ;
        RECT 103.735 202.415 104.830 202.975 ;
        RECT 105.000 202.705 105.555 203.035 ;
        RECT 102.610 201.565 102.895 202.025 ;
        RECT 103.065 201.395 103.335 201.855 ;
        RECT 103.735 201.565 104.135 202.415 ;
        RECT 105.000 202.245 105.450 202.705 ;
        RECT 105.725 202.535 106.005 203.205 ;
        RECT 104.325 202.025 105.450 202.245 ;
        RECT 104.325 201.565 104.605 202.025 ;
        RECT 105.125 201.395 105.450 201.855 ;
        RECT 105.620 201.565 106.005 202.535 ;
        RECT 108.230 201.830 108.580 203.080 ;
        RECT 110.060 202.570 110.400 203.400 ;
        RECT 112.155 203.195 113.365 203.945 ;
        RECT 112.155 202.485 112.675 203.025 ;
        RECT 112.845 202.655 113.365 203.195 ;
        RECT 106.640 201.395 111.985 201.830 ;
        RECT 112.155 201.395 113.365 202.485 ;
        RECT 22.830 201.225 113.450 201.395 ;
        RECT 22.915 200.135 24.125 201.225 ;
        RECT 24.760 200.790 30.105 201.225 ;
        RECT 30.280 200.790 35.625 201.225 ;
        RECT 22.915 199.425 23.435 199.965 ;
        RECT 23.605 199.595 24.125 200.135 ;
        RECT 26.350 199.540 26.700 200.790 ;
        RECT 22.915 198.675 24.125 199.425 ;
        RECT 28.180 199.220 28.520 200.050 ;
        RECT 31.870 199.540 32.220 200.790 ;
        RECT 35.795 200.060 36.085 201.225 ;
        RECT 36.255 200.135 37.465 201.225 ;
        RECT 37.635 200.135 41.145 201.225 ;
        RECT 41.320 200.790 46.665 201.225 ;
        RECT 46.840 200.790 52.185 201.225 ;
        RECT 33.700 199.220 34.040 200.050 ;
        RECT 36.255 199.595 36.775 200.135 ;
        RECT 36.945 199.425 37.465 199.965 ;
        RECT 37.635 199.615 39.325 200.135 ;
        RECT 39.495 199.445 41.145 199.965 ;
        RECT 42.910 199.540 43.260 200.790 ;
        RECT 24.760 198.675 30.105 199.220 ;
        RECT 30.280 198.675 35.625 199.220 ;
        RECT 35.795 198.675 36.085 199.400 ;
        RECT 36.255 198.675 37.465 199.425 ;
        RECT 37.635 198.675 41.145 199.445 ;
        RECT 44.740 199.220 45.080 200.050 ;
        RECT 48.430 199.540 48.780 200.790 ;
        RECT 52.360 200.555 52.615 201.055 ;
        RECT 52.785 200.725 53.115 201.225 ;
        RECT 52.360 200.385 53.110 200.555 ;
        RECT 50.260 199.220 50.600 200.050 ;
        RECT 52.360 199.565 52.710 200.215 ;
        RECT 52.880 199.395 53.110 200.385 ;
        RECT 52.360 199.225 53.110 199.395 ;
        RECT 41.320 198.675 46.665 199.220 ;
        RECT 46.840 198.675 52.185 199.220 ;
        RECT 52.360 198.935 52.615 199.225 ;
        RECT 52.785 198.675 53.115 199.055 ;
        RECT 53.285 198.935 53.455 201.055 ;
        RECT 53.625 200.255 53.950 201.040 ;
        RECT 54.120 200.765 54.370 201.225 ;
        RECT 54.540 200.725 54.790 201.055 ;
        RECT 55.005 200.725 55.685 201.055 ;
        RECT 54.540 200.595 54.710 200.725 ;
        RECT 54.315 200.425 54.710 200.595 ;
        RECT 53.685 199.205 54.145 200.255 ;
        RECT 54.315 199.065 54.485 200.425 ;
        RECT 54.880 200.165 55.345 200.555 ;
        RECT 54.655 199.355 55.005 199.975 ;
        RECT 55.175 199.575 55.345 200.165 ;
        RECT 55.515 199.945 55.685 200.725 ;
        RECT 55.855 200.625 56.025 200.965 ;
        RECT 56.260 200.795 56.590 201.225 ;
        RECT 56.760 200.625 56.930 200.965 ;
        RECT 57.225 200.765 57.595 201.225 ;
        RECT 55.855 200.455 56.930 200.625 ;
        RECT 57.765 200.595 57.935 201.055 ;
        RECT 58.170 200.715 59.040 201.055 ;
        RECT 59.210 200.765 59.460 201.225 ;
        RECT 57.375 200.425 57.935 200.595 ;
        RECT 57.375 200.285 57.545 200.425 ;
        RECT 56.045 200.115 57.545 200.285 ;
        RECT 58.240 200.255 58.700 200.545 ;
        RECT 55.515 199.775 57.205 199.945 ;
        RECT 55.175 199.355 55.530 199.575 ;
        RECT 55.700 199.065 55.870 199.775 ;
        RECT 56.075 199.355 56.865 199.605 ;
        RECT 57.035 199.595 57.205 199.775 ;
        RECT 57.375 199.425 57.545 200.115 ;
        RECT 53.815 198.675 54.145 199.035 ;
        RECT 54.315 198.895 54.810 199.065 ;
        RECT 55.015 198.895 55.870 199.065 ;
        RECT 56.745 198.675 57.075 199.135 ;
        RECT 57.285 199.035 57.545 199.425 ;
        RECT 57.735 200.245 58.700 200.255 ;
        RECT 58.870 200.335 59.040 200.715 ;
        RECT 59.630 200.675 59.800 200.965 ;
        RECT 59.980 200.845 60.310 201.225 ;
        RECT 59.630 200.505 60.430 200.675 ;
        RECT 57.735 200.085 58.410 200.245 ;
        RECT 58.870 200.165 60.090 200.335 ;
        RECT 57.735 199.295 57.945 200.085 ;
        RECT 58.870 200.075 59.040 200.165 ;
        RECT 58.115 199.295 58.465 199.915 ;
        RECT 58.635 199.905 59.040 200.075 ;
        RECT 58.635 199.125 58.805 199.905 ;
        RECT 58.975 199.455 59.195 199.735 ;
        RECT 59.375 199.625 59.915 199.995 ;
        RECT 60.260 199.915 60.430 200.505 ;
        RECT 60.650 200.085 60.955 201.225 ;
        RECT 61.125 200.035 61.380 200.915 ;
        RECT 61.555 200.060 61.845 201.225 ;
        RECT 62.015 200.135 63.685 201.225 ;
        RECT 63.875 200.715 64.175 201.225 ;
        RECT 64.345 200.715 64.725 200.885 ;
        RECT 65.305 200.715 65.935 201.225 ;
        RECT 64.345 200.545 64.515 200.715 ;
        RECT 66.105 200.545 66.435 201.055 ;
        RECT 66.605 200.715 66.905 201.225 ;
        RECT 67.160 200.605 67.335 201.055 ;
        RECT 67.505 200.785 67.835 201.225 ;
        RECT 68.140 200.635 68.310 201.055 ;
        RECT 68.545 200.815 69.215 201.225 ;
        RECT 69.430 200.635 69.600 201.055 ;
        RECT 69.800 200.815 70.130 201.225 ;
        RECT 63.855 200.345 64.515 200.545 ;
        RECT 64.685 200.375 66.905 200.545 ;
        RECT 67.160 200.435 67.790 200.605 ;
        RECT 60.260 199.885 61.000 199.915 ;
        RECT 58.975 199.285 59.505 199.455 ;
        RECT 57.285 198.865 57.635 199.035 ;
        RECT 57.855 198.845 58.805 199.125 ;
        RECT 58.975 198.675 59.165 199.115 ;
        RECT 59.335 199.055 59.505 199.285 ;
        RECT 59.675 199.225 59.915 199.625 ;
        RECT 60.085 199.585 61.000 199.885 ;
        RECT 60.085 199.410 60.410 199.585 ;
        RECT 60.085 199.055 60.405 199.410 ;
        RECT 61.170 199.385 61.380 200.035 ;
        RECT 62.015 199.615 62.765 200.135 ;
        RECT 62.935 199.445 63.685 199.965 ;
        RECT 59.335 198.885 60.405 199.055 ;
        RECT 60.650 198.675 60.955 199.135 ;
        RECT 61.125 198.855 61.380 199.385 ;
        RECT 61.555 198.675 61.845 199.400 ;
        RECT 62.015 198.675 63.685 199.445 ;
        RECT 63.855 199.415 64.025 200.345 ;
        RECT 64.685 200.175 64.855 200.375 ;
        RECT 64.195 200.005 64.855 200.175 ;
        RECT 65.025 200.035 66.565 200.205 ;
        RECT 64.195 199.585 64.365 200.005 ;
        RECT 65.025 199.835 65.195 200.035 ;
        RECT 64.595 199.665 65.195 199.835 ;
        RECT 65.365 199.665 66.060 199.865 ;
        RECT 66.320 199.585 66.565 200.035 ;
        RECT 64.685 199.415 65.595 199.495 ;
        RECT 63.855 198.935 64.175 199.415 ;
        RECT 64.345 199.325 65.595 199.415 ;
        RECT 64.345 199.245 64.855 199.325 ;
        RECT 64.345 198.845 64.575 199.245 ;
        RECT 64.745 198.675 65.095 199.065 ;
        RECT 65.265 198.845 65.595 199.325 ;
        RECT 65.765 198.675 65.935 199.495 ;
        RECT 66.735 199.415 66.905 200.375 ;
        RECT 67.075 199.585 67.440 200.265 ;
        RECT 67.620 199.915 67.790 200.435 ;
        RECT 68.140 200.465 70.155 200.635 ;
        RECT 67.620 199.585 67.970 199.915 ;
        RECT 67.620 199.415 67.790 199.585 ;
        RECT 66.440 198.870 66.905 199.415 ;
        RECT 67.160 199.245 67.790 199.415 ;
        RECT 67.160 198.845 67.335 199.245 ;
        RECT 68.140 199.175 68.310 200.465 ;
        RECT 67.505 198.675 67.835 199.055 ;
        RECT 68.080 198.845 68.310 199.175 ;
        RECT 68.510 199.010 68.790 200.285 ;
        RECT 69.015 199.865 69.285 200.285 ;
        RECT 68.975 199.695 69.285 199.865 ;
        RECT 69.015 199.010 69.285 199.695 ;
        RECT 69.475 199.255 69.815 200.285 ;
        RECT 69.985 199.915 70.155 200.465 ;
        RECT 70.325 200.085 70.585 201.055 ;
        RECT 69.985 199.585 70.245 199.915 ;
        RECT 70.415 199.395 70.585 200.085 ;
        RECT 69.745 198.675 70.075 199.055 ;
        RECT 70.245 198.930 70.585 199.395 ;
        RECT 70.760 200.035 71.015 200.915 ;
        RECT 71.185 200.085 71.490 201.225 ;
        RECT 71.830 200.845 72.160 201.225 ;
        RECT 72.340 200.675 72.510 200.965 ;
        RECT 72.680 200.765 72.930 201.225 ;
        RECT 71.710 200.505 72.510 200.675 ;
        RECT 73.100 200.715 73.970 201.055 ;
        RECT 70.760 199.385 70.970 200.035 ;
        RECT 71.710 199.915 71.880 200.505 ;
        RECT 73.100 200.335 73.270 200.715 ;
        RECT 74.205 200.595 74.375 201.055 ;
        RECT 74.545 200.765 74.915 201.225 ;
        RECT 75.210 200.625 75.380 200.965 ;
        RECT 75.550 200.795 75.880 201.225 ;
        RECT 76.115 200.625 76.285 200.965 ;
        RECT 72.050 200.165 73.270 200.335 ;
        RECT 73.440 200.255 73.900 200.545 ;
        RECT 74.205 200.425 74.765 200.595 ;
        RECT 75.210 200.455 76.285 200.625 ;
        RECT 76.455 200.725 77.135 201.055 ;
        RECT 77.350 200.725 77.600 201.055 ;
        RECT 77.770 200.765 78.020 201.225 ;
        RECT 74.595 200.285 74.765 200.425 ;
        RECT 73.440 200.245 74.405 200.255 ;
        RECT 73.100 200.075 73.270 200.165 ;
        RECT 73.730 200.085 74.405 200.245 ;
        RECT 71.140 199.885 71.880 199.915 ;
        RECT 71.140 199.585 72.055 199.885 ;
        RECT 71.730 199.410 72.055 199.585 ;
        RECT 70.245 198.885 70.580 198.930 ;
        RECT 70.760 198.855 71.015 199.385 ;
        RECT 71.185 198.675 71.490 199.135 ;
        RECT 71.735 199.055 72.055 199.410 ;
        RECT 72.225 199.625 72.765 199.995 ;
        RECT 73.100 199.905 73.505 200.075 ;
        RECT 72.225 199.225 72.465 199.625 ;
        RECT 72.945 199.455 73.165 199.735 ;
        RECT 72.635 199.285 73.165 199.455 ;
        RECT 72.635 199.055 72.805 199.285 ;
        RECT 73.335 199.125 73.505 199.905 ;
        RECT 73.675 199.295 74.025 199.915 ;
        RECT 74.195 199.295 74.405 200.085 ;
        RECT 74.595 200.115 76.095 200.285 ;
        RECT 74.595 199.425 74.765 200.115 ;
        RECT 76.455 199.945 76.625 200.725 ;
        RECT 77.430 200.595 77.600 200.725 ;
        RECT 74.935 199.775 76.625 199.945 ;
        RECT 76.795 200.165 77.260 200.555 ;
        RECT 77.430 200.425 77.825 200.595 ;
        RECT 74.935 199.595 75.105 199.775 ;
        RECT 71.735 198.885 72.805 199.055 ;
        RECT 72.975 198.675 73.165 199.115 ;
        RECT 73.335 198.845 74.285 199.125 ;
        RECT 74.595 199.035 74.855 199.425 ;
        RECT 75.275 199.355 76.065 199.605 ;
        RECT 74.505 198.865 74.855 199.035 ;
        RECT 75.065 198.675 75.395 199.135 ;
        RECT 76.270 199.065 76.440 199.775 ;
        RECT 76.795 199.575 76.965 200.165 ;
        RECT 76.610 199.355 76.965 199.575 ;
        RECT 77.135 199.355 77.485 199.975 ;
        RECT 77.655 199.065 77.825 200.425 ;
        RECT 78.190 200.255 78.515 201.040 ;
        RECT 77.995 199.205 78.455 200.255 ;
        RECT 76.270 198.895 77.125 199.065 ;
        RECT 77.330 198.895 77.825 199.065 ;
        RECT 77.995 198.675 78.325 199.035 ;
        RECT 78.685 198.935 78.855 201.055 ;
        RECT 79.025 200.725 79.355 201.225 ;
        RECT 79.525 200.555 79.780 201.055 ;
        RECT 79.975 200.715 80.275 201.225 ;
        RECT 80.445 200.715 80.825 200.885 ;
        RECT 81.405 200.715 82.035 201.225 ;
        RECT 79.030 200.385 79.780 200.555 ;
        RECT 80.445 200.545 80.615 200.715 ;
        RECT 82.205 200.545 82.535 201.055 ;
        RECT 82.705 200.715 83.005 201.225 ;
        RECT 79.030 199.395 79.260 200.385 ;
        RECT 79.955 200.345 80.615 200.545 ;
        RECT 80.785 200.375 83.005 200.545 ;
        RECT 79.430 199.565 79.780 200.215 ;
        RECT 79.955 199.415 80.125 200.345 ;
        RECT 80.785 200.175 80.955 200.375 ;
        RECT 80.295 200.005 80.955 200.175 ;
        RECT 81.125 200.035 82.665 200.205 ;
        RECT 80.295 199.585 80.465 200.005 ;
        RECT 81.125 199.835 81.295 200.035 ;
        RECT 80.695 199.665 81.295 199.835 ;
        RECT 81.465 199.665 82.160 199.865 ;
        RECT 82.420 199.585 82.665 200.035 ;
        RECT 80.785 199.415 81.695 199.495 ;
        RECT 79.030 199.225 79.780 199.395 ;
        RECT 79.025 198.675 79.355 199.055 ;
        RECT 79.525 198.935 79.780 199.225 ;
        RECT 79.955 198.935 80.275 199.415 ;
        RECT 80.445 199.325 81.695 199.415 ;
        RECT 80.445 199.245 80.955 199.325 ;
        RECT 80.445 198.845 80.675 199.245 ;
        RECT 80.845 198.675 81.195 199.065 ;
        RECT 81.365 198.845 81.695 199.325 ;
        RECT 81.865 198.675 82.035 199.495 ;
        RECT 82.835 199.415 83.005 200.375 ;
        RECT 83.175 200.135 85.765 201.225 ;
        RECT 83.175 199.615 84.385 200.135 ;
        RECT 85.975 200.085 86.205 201.225 ;
        RECT 86.375 200.075 86.705 201.055 ;
        RECT 86.875 200.085 87.085 201.225 ;
        RECT 84.555 199.445 85.765 199.965 ;
        RECT 85.955 199.665 86.285 199.915 ;
        RECT 82.540 198.870 83.005 199.415 ;
        RECT 83.175 198.675 85.765 199.445 ;
        RECT 85.975 198.675 86.205 199.495 ;
        RECT 86.455 199.475 86.705 200.075 ;
        RECT 87.315 200.060 87.605 201.225 ;
        RECT 88.735 200.085 88.965 201.225 ;
        RECT 89.135 200.075 89.465 201.055 ;
        RECT 89.635 200.085 89.845 201.225 ;
        RECT 90.190 200.595 90.475 201.055 ;
        RECT 90.645 200.765 90.915 201.225 ;
        RECT 90.190 200.375 91.145 200.595 ;
        RECT 88.715 199.665 89.045 199.915 ;
        RECT 86.375 198.845 86.705 199.475 ;
        RECT 86.875 198.675 87.085 199.495 ;
        RECT 87.315 198.675 87.605 199.400 ;
        RECT 88.735 198.675 88.965 199.495 ;
        RECT 89.215 199.475 89.465 200.075 ;
        RECT 90.075 199.645 90.765 200.205 ;
        RECT 89.135 198.845 89.465 199.475 ;
        RECT 89.635 198.675 89.845 199.495 ;
        RECT 90.935 199.475 91.145 200.375 ;
        RECT 90.190 199.305 91.145 199.475 ;
        RECT 91.315 200.205 91.715 201.055 ;
        RECT 91.905 200.595 92.185 201.055 ;
        RECT 92.705 200.765 93.030 201.225 ;
        RECT 91.905 200.375 93.030 200.595 ;
        RECT 91.315 199.645 92.410 200.205 ;
        RECT 92.580 199.915 93.030 200.375 ;
        RECT 93.200 200.085 93.585 201.055 ;
        RECT 93.870 200.595 94.155 201.055 ;
        RECT 94.325 200.765 94.595 201.225 ;
        RECT 93.870 200.375 94.825 200.595 ;
        RECT 90.190 198.845 90.475 199.305 ;
        RECT 90.645 198.675 90.915 199.135 ;
        RECT 91.315 198.845 91.715 199.645 ;
        RECT 92.580 199.585 93.135 199.915 ;
        RECT 92.580 199.475 93.030 199.585 ;
        RECT 91.905 199.305 93.030 199.475 ;
        RECT 93.305 199.415 93.585 200.085 ;
        RECT 93.755 199.645 94.445 200.205 ;
        RECT 94.615 199.475 94.825 200.375 ;
        RECT 91.905 198.845 92.185 199.305 ;
        RECT 92.705 198.675 93.030 199.135 ;
        RECT 93.200 198.845 93.585 199.415 ;
        RECT 93.870 199.305 94.825 199.475 ;
        RECT 94.995 200.205 95.395 201.055 ;
        RECT 95.585 200.595 95.865 201.055 ;
        RECT 96.385 200.765 96.710 201.225 ;
        RECT 95.585 200.375 96.710 200.595 ;
        RECT 94.995 199.645 96.090 200.205 ;
        RECT 96.260 199.915 96.710 200.375 ;
        RECT 96.880 200.085 97.265 201.055 ;
        RECT 93.870 198.845 94.155 199.305 ;
        RECT 94.325 198.675 94.595 199.135 ;
        RECT 94.995 198.845 95.395 199.645 ;
        RECT 96.260 199.585 96.815 199.915 ;
        RECT 96.260 199.475 96.710 199.585 ;
        RECT 95.585 199.305 96.710 199.475 ;
        RECT 96.985 199.415 97.265 200.085 ;
        RECT 95.585 198.845 95.865 199.305 ;
        RECT 96.385 198.675 96.710 199.135 ;
        RECT 96.880 198.845 97.265 199.415 ;
        RECT 97.440 200.035 97.695 200.915 ;
        RECT 97.865 200.085 98.170 201.225 ;
        RECT 98.510 200.845 98.840 201.225 ;
        RECT 99.020 200.675 99.190 200.965 ;
        RECT 99.360 200.765 99.610 201.225 ;
        RECT 98.390 200.505 99.190 200.675 ;
        RECT 99.780 200.715 100.650 201.055 ;
        RECT 97.440 199.385 97.650 200.035 ;
        RECT 98.390 199.915 98.560 200.505 ;
        RECT 99.780 200.335 99.950 200.715 ;
        RECT 100.885 200.595 101.055 201.055 ;
        RECT 101.225 200.765 101.595 201.225 ;
        RECT 101.890 200.625 102.060 200.965 ;
        RECT 102.230 200.795 102.560 201.225 ;
        RECT 102.795 200.625 102.965 200.965 ;
        RECT 98.730 200.165 99.950 200.335 ;
        RECT 100.120 200.255 100.580 200.545 ;
        RECT 100.885 200.425 101.445 200.595 ;
        RECT 101.890 200.455 102.965 200.625 ;
        RECT 103.135 200.725 103.815 201.055 ;
        RECT 104.030 200.725 104.280 201.055 ;
        RECT 104.450 200.765 104.700 201.225 ;
        RECT 101.275 200.285 101.445 200.425 ;
        RECT 100.120 200.245 101.085 200.255 ;
        RECT 99.780 200.075 99.950 200.165 ;
        RECT 100.410 200.085 101.085 200.245 ;
        RECT 97.820 199.885 98.560 199.915 ;
        RECT 97.820 199.585 98.735 199.885 ;
        RECT 98.410 199.410 98.735 199.585 ;
        RECT 97.440 198.855 97.695 199.385 ;
        RECT 97.865 198.675 98.170 199.135 ;
        RECT 98.415 199.055 98.735 199.410 ;
        RECT 98.905 199.625 99.445 199.995 ;
        RECT 99.780 199.905 100.185 200.075 ;
        RECT 98.905 199.225 99.145 199.625 ;
        RECT 99.625 199.455 99.845 199.735 ;
        RECT 99.315 199.285 99.845 199.455 ;
        RECT 99.315 199.055 99.485 199.285 ;
        RECT 100.015 199.125 100.185 199.905 ;
        RECT 100.355 199.295 100.705 199.915 ;
        RECT 100.875 199.295 101.085 200.085 ;
        RECT 101.275 200.115 102.775 200.285 ;
        RECT 101.275 199.425 101.445 200.115 ;
        RECT 103.135 199.945 103.305 200.725 ;
        RECT 104.110 200.595 104.280 200.725 ;
        RECT 101.615 199.775 103.305 199.945 ;
        RECT 103.475 200.165 103.940 200.555 ;
        RECT 104.110 200.425 104.505 200.595 ;
        RECT 101.615 199.595 101.785 199.775 ;
        RECT 98.415 198.885 99.485 199.055 ;
        RECT 99.655 198.675 99.845 199.115 ;
        RECT 100.015 198.845 100.965 199.125 ;
        RECT 101.275 199.035 101.535 199.425 ;
        RECT 101.955 199.355 102.745 199.605 ;
        RECT 101.185 198.865 101.535 199.035 ;
        RECT 101.745 198.675 102.075 199.135 ;
        RECT 102.950 199.065 103.120 199.775 ;
        RECT 103.475 199.575 103.645 200.165 ;
        RECT 103.290 199.355 103.645 199.575 ;
        RECT 103.815 199.355 104.165 199.975 ;
        RECT 104.335 199.065 104.505 200.425 ;
        RECT 104.870 200.255 105.195 201.040 ;
        RECT 104.675 199.205 105.135 200.255 ;
        RECT 102.950 198.895 103.805 199.065 ;
        RECT 104.010 198.895 104.505 199.065 ;
        RECT 104.675 198.675 105.005 199.035 ;
        RECT 105.365 198.935 105.535 201.055 ;
        RECT 105.705 200.725 106.035 201.225 ;
        RECT 106.205 200.555 106.460 201.055 ;
        RECT 105.710 200.385 106.460 200.555 ;
        RECT 105.710 199.395 105.940 200.385 ;
        RECT 106.110 199.565 106.460 200.215 ;
        RECT 107.095 200.150 107.365 201.055 ;
        RECT 107.535 200.465 107.865 201.225 ;
        RECT 108.045 200.295 108.215 201.055 ;
        RECT 105.710 199.225 106.460 199.395 ;
        RECT 105.705 198.675 106.035 199.055 ;
        RECT 106.205 198.935 106.460 199.225 ;
        RECT 107.095 199.350 107.265 200.150 ;
        RECT 107.550 200.125 108.215 200.295 ;
        RECT 108.475 200.135 111.985 201.225 ;
        RECT 112.155 200.135 113.365 201.225 ;
        RECT 107.550 199.980 107.720 200.125 ;
        RECT 107.435 199.650 107.720 199.980 ;
        RECT 107.550 199.395 107.720 199.650 ;
        RECT 107.955 199.575 108.285 199.945 ;
        RECT 108.475 199.615 110.165 200.135 ;
        RECT 110.335 199.445 111.985 199.965 ;
        RECT 112.155 199.595 112.675 200.135 ;
        RECT 107.095 198.845 107.355 199.350 ;
        RECT 107.550 199.225 108.215 199.395 ;
        RECT 107.535 198.675 107.865 199.055 ;
        RECT 108.045 198.845 108.215 199.225 ;
        RECT 108.475 198.675 111.985 199.445 ;
        RECT 112.845 199.425 113.365 199.965 ;
        RECT 112.155 198.675 113.365 199.425 ;
        RECT 22.830 198.505 113.450 198.675 ;
        RECT 22.915 197.755 24.125 198.505 ;
        RECT 22.915 197.215 23.435 197.755 ;
        RECT 24.755 197.735 26.425 198.505 ;
        RECT 26.600 197.960 31.945 198.505 ;
        RECT 32.120 197.960 37.465 198.505 ;
        RECT 37.640 197.960 42.985 198.505 ;
        RECT 43.160 197.960 48.505 198.505 ;
        RECT 23.605 197.045 24.125 197.585 ;
        RECT 22.915 195.955 24.125 197.045 ;
        RECT 24.755 197.045 25.505 197.565 ;
        RECT 25.675 197.215 26.425 197.735 ;
        RECT 24.755 195.955 26.425 197.045 ;
        RECT 28.190 196.390 28.540 197.640 ;
        RECT 30.020 197.130 30.360 197.960 ;
        RECT 33.710 196.390 34.060 197.640 ;
        RECT 35.540 197.130 35.880 197.960 ;
        RECT 39.230 196.390 39.580 197.640 ;
        RECT 41.060 197.130 41.400 197.960 ;
        RECT 44.750 196.390 45.100 197.640 ;
        RECT 46.580 197.130 46.920 197.960 ;
        RECT 48.675 197.780 48.965 198.505 ;
        RECT 49.135 197.830 49.395 198.335 ;
        RECT 49.575 198.125 49.905 198.505 ;
        RECT 50.085 197.955 50.255 198.335 ;
        RECT 26.600 195.955 31.945 196.390 ;
        RECT 32.120 195.955 37.465 196.390 ;
        RECT 37.640 195.955 42.985 196.390 ;
        RECT 43.160 195.955 48.505 196.390 ;
        RECT 48.675 195.955 48.965 197.120 ;
        RECT 49.135 197.030 49.305 197.830 ;
        RECT 49.590 197.785 50.255 197.955 ;
        RECT 49.590 197.530 49.760 197.785 ;
        RECT 50.975 197.735 54.485 198.505 ;
        RECT 54.660 197.955 54.915 198.245 ;
        RECT 55.085 198.125 55.415 198.505 ;
        RECT 54.660 197.785 55.410 197.955 ;
        RECT 49.475 197.200 49.760 197.530 ;
        RECT 49.995 197.235 50.325 197.605 ;
        RECT 49.590 197.055 49.760 197.200 ;
        RECT 49.135 196.125 49.405 197.030 ;
        RECT 49.590 196.885 50.255 197.055 ;
        RECT 49.575 195.955 49.905 196.715 ;
        RECT 50.085 196.125 50.255 196.885 ;
        RECT 50.975 197.045 52.665 197.565 ;
        RECT 52.835 197.215 54.485 197.735 ;
        RECT 50.975 195.955 54.485 197.045 ;
        RECT 54.660 196.965 55.010 197.615 ;
        RECT 55.180 196.795 55.410 197.785 ;
        RECT 54.660 196.625 55.410 196.795 ;
        RECT 54.660 196.125 54.915 196.625 ;
        RECT 55.085 195.955 55.415 196.455 ;
        RECT 55.585 196.125 55.755 198.245 ;
        RECT 56.115 198.145 56.445 198.505 ;
        RECT 56.615 198.115 57.110 198.285 ;
        RECT 57.315 198.115 58.170 198.285 ;
        RECT 55.985 196.925 56.445 197.975 ;
        RECT 55.925 196.140 56.250 196.925 ;
        RECT 56.615 196.755 56.785 198.115 ;
        RECT 56.955 197.205 57.305 197.825 ;
        RECT 57.475 197.605 57.830 197.825 ;
        RECT 57.475 197.015 57.645 197.605 ;
        RECT 58.000 197.405 58.170 198.115 ;
        RECT 59.045 198.045 59.375 198.505 ;
        RECT 59.585 198.145 59.935 198.315 ;
        RECT 58.375 197.575 59.165 197.825 ;
        RECT 59.585 197.755 59.845 198.145 ;
        RECT 60.155 198.055 61.105 198.335 ;
        RECT 61.275 198.065 61.465 198.505 ;
        RECT 61.635 198.125 62.705 198.295 ;
        RECT 59.335 197.405 59.505 197.585 ;
        RECT 56.615 196.585 57.010 196.755 ;
        RECT 57.180 196.625 57.645 197.015 ;
        RECT 57.815 197.235 59.505 197.405 ;
        RECT 56.840 196.455 57.010 196.585 ;
        RECT 57.815 196.455 57.985 197.235 ;
        RECT 59.675 197.065 59.845 197.755 ;
        RECT 58.345 196.895 59.845 197.065 ;
        RECT 60.035 197.095 60.245 197.885 ;
        RECT 60.415 197.265 60.765 197.885 ;
        RECT 60.935 197.275 61.105 198.055 ;
        RECT 61.635 197.895 61.805 198.125 ;
        RECT 61.275 197.725 61.805 197.895 ;
        RECT 61.275 197.445 61.495 197.725 ;
        RECT 61.975 197.555 62.215 197.955 ;
        RECT 60.935 197.105 61.340 197.275 ;
        RECT 61.675 197.185 62.215 197.555 ;
        RECT 62.385 197.770 62.705 198.125 ;
        RECT 62.385 197.515 62.710 197.770 ;
        RECT 62.905 197.695 63.075 198.505 ;
        RECT 63.245 197.855 63.575 198.335 ;
        RECT 63.745 198.035 63.915 198.505 ;
        RECT 64.085 197.855 64.415 198.335 ;
        RECT 64.585 198.035 64.755 198.505 ;
        RECT 65.350 197.875 65.635 198.335 ;
        RECT 65.805 198.045 66.075 198.505 ;
        RECT 63.245 197.685 65.010 197.855 ;
        RECT 65.350 197.705 66.305 197.875 ;
        RECT 62.385 197.305 64.415 197.515 ;
        RECT 62.385 197.295 62.730 197.305 ;
        RECT 60.035 196.935 60.710 197.095 ;
        RECT 61.170 197.015 61.340 197.105 ;
        RECT 60.035 196.925 61.000 196.935 ;
        RECT 59.675 196.755 59.845 196.895 ;
        RECT 56.420 195.955 56.670 196.415 ;
        RECT 56.840 196.125 57.090 196.455 ;
        RECT 57.305 196.125 57.985 196.455 ;
        RECT 58.155 196.555 59.230 196.725 ;
        RECT 59.675 196.585 60.235 196.755 ;
        RECT 60.540 196.635 61.000 196.925 ;
        RECT 61.170 196.845 62.390 197.015 ;
        RECT 58.155 196.215 58.325 196.555 ;
        RECT 58.560 195.955 58.890 196.385 ;
        RECT 59.060 196.215 59.230 196.555 ;
        RECT 59.525 195.955 59.895 196.415 ;
        RECT 60.065 196.125 60.235 196.585 ;
        RECT 61.170 196.465 61.340 196.845 ;
        RECT 62.560 196.675 62.730 197.295 ;
        RECT 64.600 197.135 65.010 197.685 ;
        RECT 60.470 196.125 61.340 196.465 ;
        RECT 61.930 196.505 62.730 196.675 ;
        RECT 61.510 195.955 61.760 196.415 ;
        RECT 61.930 196.215 62.100 196.505 ;
        RECT 62.280 195.955 62.610 196.335 ;
        RECT 62.905 195.955 63.075 197.015 ;
        RECT 63.285 196.965 65.010 197.135 ;
        RECT 65.235 196.975 65.925 197.535 ;
        RECT 63.285 196.125 63.575 196.965 ;
        RECT 63.745 195.955 63.915 196.795 ;
        RECT 64.125 196.125 64.375 196.965 ;
        RECT 66.095 196.805 66.305 197.705 ;
        RECT 64.585 195.955 64.755 196.795 ;
        RECT 65.350 196.585 66.305 196.805 ;
        RECT 66.475 197.535 66.875 198.335 ;
        RECT 67.065 197.875 67.345 198.335 ;
        RECT 67.865 198.045 68.190 198.505 ;
        RECT 67.065 197.705 68.190 197.875 ;
        RECT 68.360 197.765 68.745 198.335 ;
        RECT 67.740 197.595 68.190 197.705 ;
        RECT 66.475 196.975 67.570 197.535 ;
        RECT 67.740 197.265 68.295 197.595 ;
        RECT 65.350 196.125 65.635 196.585 ;
        RECT 65.805 195.955 66.075 196.415 ;
        RECT 66.475 196.125 66.875 196.975 ;
        RECT 67.740 196.805 68.190 197.265 ;
        RECT 68.465 197.095 68.745 197.765 ;
        RECT 68.920 197.665 69.180 198.505 ;
        RECT 69.355 197.760 69.610 198.335 ;
        RECT 69.780 198.125 70.110 198.505 ;
        RECT 70.325 197.955 70.495 198.335 ;
        RECT 69.780 197.785 70.495 197.955 ;
        RECT 70.870 197.875 71.155 198.335 ;
        RECT 71.325 198.045 71.595 198.505 ;
        RECT 67.065 196.585 68.190 196.805 ;
        RECT 67.065 196.125 67.345 196.585 ;
        RECT 67.865 195.955 68.190 196.415 ;
        RECT 68.360 196.125 68.745 197.095 ;
        RECT 68.920 195.955 69.180 197.105 ;
        RECT 69.355 197.030 69.525 197.760 ;
        RECT 69.780 197.595 69.950 197.785 ;
        RECT 70.870 197.705 71.825 197.875 ;
        RECT 69.695 197.265 69.950 197.595 ;
        RECT 69.780 197.055 69.950 197.265 ;
        RECT 70.230 197.235 70.585 197.605 ;
        RECT 69.355 196.125 69.610 197.030 ;
        RECT 69.780 196.885 70.495 197.055 ;
        RECT 70.755 196.975 71.445 197.535 ;
        RECT 69.780 195.955 70.110 196.715 ;
        RECT 70.325 196.125 70.495 196.885 ;
        RECT 71.615 196.805 71.825 197.705 ;
        RECT 70.870 196.585 71.825 196.805 ;
        RECT 71.995 197.535 72.395 198.335 ;
        RECT 72.585 197.875 72.865 198.335 ;
        RECT 73.385 198.045 73.710 198.505 ;
        RECT 72.585 197.705 73.710 197.875 ;
        RECT 73.880 197.765 74.265 198.335 ;
        RECT 74.435 197.780 74.725 198.505 ;
        RECT 75.355 197.855 75.615 198.335 ;
        RECT 75.785 197.965 76.035 198.505 ;
        RECT 73.260 197.595 73.710 197.705 ;
        RECT 71.995 196.975 73.090 197.535 ;
        RECT 73.260 197.265 73.815 197.595 ;
        RECT 70.870 196.125 71.155 196.585 ;
        RECT 71.325 195.955 71.595 196.415 ;
        RECT 71.995 196.125 72.395 196.975 ;
        RECT 73.260 196.805 73.710 197.265 ;
        RECT 73.985 197.095 74.265 197.765 ;
        RECT 72.585 196.585 73.710 196.805 ;
        RECT 72.585 196.125 72.865 196.585 ;
        RECT 73.385 195.955 73.710 196.415 ;
        RECT 73.880 196.125 74.265 197.095 ;
        RECT 74.435 195.955 74.725 197.120 ;
        RECT 75.355 196.825 75.525 197.855 ;
        RECT 76.205 197.825 76.425 198.285 ;
        RECT 76.175 197.800 76.425 197.825 ;
        RECT 75.695 197.205 75.925 197.600 ;
        RECT 76.095 197.375 76.425 197.800 ;
        RECT 76.595 198.125 77.485 198.295 ;
        RECT 76.595 197.400 76.765 198.125 ;
        RECT 76.935 197.570 77.485 197.955 ;
        RECT 77.660 197.795 77.915 198.325 ;
        RECT 78.085 198.045 78.390 198.505 ;
        RECT 78.635 198.125 79.705 198.295 ;
        RECT 76.595 197.330 77.485 197.400 ;
        RECT 76.590 197.305 77.485 197.330 ;
        RECT 76.580 197.290 77.485 197.305 ;
        RECT 76.575 197.275 77.485 197.290 ;
        RECT 76.565 197.270 77.485 197.275 ;
        RECT 76.560 197.260 77.485 197.270 ;
        RECT 76.555 197.250 77.485 197.260 ;
        RECT 76.545 197.245 77.485 197.250 ;
        RECT 76.535 197.235 77.485 197.245 ;
        RECT 76.525 197.230 77.485 197.235 ;
        RECT 76.525 197.225 76.860 197.230 ;
        RECT 76.510 197.220 76.860 197.225 ;
        RECT 76.495 197.210 76.860 197.220 ;
        RECT 76.470 197.205 76.860 197.210 ;
        RECT 75.695 197.200 76.860 197.205 ;
        RECT 75.695 197.165 76.830 197.200 ;
        RECT 75.695 197.140 76.795 197.165 ;
        RECT 75.695 197.110 76.765 197.140 ;
        RECT 75.695 197.080 76.745 197.110 ;
        RECT 75.695 197.050 76.725 197.080 ;
        RECT 75.695 197.040 76.655 197.050 ;
        RECT 75.695 197.030 76.630 197.040 ;
        RECT 75.695 197.015 76.610 197.030 ;
        RECT 75.695 197.000 76.590 197.015 ;
        RECT 75.800 196.990 76.585 197.000 ;
        RECT 75.800 196.955 76.570 196.990 ;
        RECT 75.355 196.125 75.630 196.825 ;
        RECT 75.800 196.705 76.555 196.955 ;
        RECT 76.725 196.635 77.055 196.880 ;
        RECT 77.225 196.780 77.485 197.230 ;
        RECT 77.660 197.145 77.870 197.795 ;
        RECT 78.635 197.770 78.955 198.125 ;
        RECT 78.630 197.595 78.955 197.770 ;
        RECT 78.040 197.295 78.955 197.595 ;
        RECT 79.125 197.555 79.365 197.955 ;
        RECT 79.535 197.895 79.705 198.125 ;
        RECT 79.875 198.065 80.065 198.505 ;
        RECT 80.235 198.055 81.185 198.335 ;
        RECT 81.405 198.145 81.755 198.315 ;
        RECT 79.535 197.725 80.065 197.895 ;
        RECT 78.040 197.265 78.780 197.295 ;
        RECT 76.870 196.610 77.055 196.635 ;
        RECT 76.870 196.510 77.485 196.610 ;
        RECT 75.800 195.955 76.055 196.500 ;
        RECT 76.225 196.125 76.705 196.465 ;
        RECT 76.880 195.955 77.485 196.510 ;
        RECT 77.660 196.265 77.915 197.145 ;
        RECT 78.085 195.955 78.390 197.095 ;
        RECT 78.610 196.675 78.780 197.265 ;
        RECT 79.125 197.185 79.665 197.555 ;
        RECT 79.845 197.445 80.065 197.725 ;
        RECT 80.235 197.275 80.405 198.055 ;
        RECT 80.000 197.105 80.405 197.275 ;
        RECT 80.575 197.265 80.925 197.885 ;
        RECT 80.000 197.015 80.170 197.105 ;
        RECT 81.095 197.095 81.305 197.885 ;
        RECT 78.950 196.845 80.170 197.015 ;
        RECT 80.630 196.935 81.305 197.095 ;
        RECT 78.610 196.505 79.410 196.675 ;
        RECT 78.730 195.955 79.060 196.335 ;
        RECT 79.240 196.215 79.410 196.505 ;
        RECT 80.000 196.465 80.170 196.845 ;
        RECT 80.340 196.925 81.305 196.935 ;
        RECT 81.495 197.755 81.755 198.145 ;
        RECT 81.965 198.045 82.295 198.505 ;
        RECT 83.170 198.115 84.025 198.285 ;
        RECT 84.230 198.115 84.725 198.285 ;
        RECT 84.895 198.145 85.225 198.505 ;
        RECT 81.495 197.065 81.665 197.755 ;
        RECT 81.835 197.405 82.005 197.585 ;
        RECT 82.175 197.575 82.965 197.825 ;
        RECT 83.170 197.405 83.340 198.115 ;
        RECT 83.510 197.605 83.865 197.825 ;
        RECT 81.835 197.235 83.525 197.405 ;
        RECT 80.340 196.635 80.800 196.925 ;
        RECT 81.495 196.895 82.995 197.065 ;
        RECT 81.495 196.755 81.665 196.895 ;
        RECT 81.105 196.585 81.665 196.755 ;
        RECT 79.580 195.955 79.830 196.415 ;
        RECT 80.000 196.125 80.870 196.465 ;
        RECT 81.105 196.125 81.275 196.585 ;
        RECT 82.110 196.555 83.185 196.725 ;
        RECT 81.445 195.955 81.815 196.415 ;
        RECT 82.110 196.215 82.280 196.555 ;
        RECT 82.450 195.955 82.780 196.385 ;
        RECT 83.015 196.215 83.185 196.555 ;
        RECT 83.355 196.455 83.525 197.235 ;
        RECT 83.695 197.015 83.865 197.605 ;
        RECT 84.035 197.205 84.385 197.825 ;
        RECT 83.695 196.625 84.160 197.015 ;
        RECT 84.555 196.755 84.725 198.115 ;
        RECT 84.895 196.925 85.355 197.975 ;
        RECT 84.330 196.585 84.725 196.755 ;
        RECT 84.330 196.455 84.500 196.585 ;
        RECT 83.355 196.125 84.035 196.455 ;
        RECT 84.250 196.125 84.500 196.455 ;
        RECT 84.670 195.955 84.920 196.415 ;
        RECT 85.090 196.140 85.415 196.925 ;
        RECT 85.585 196.125 85.755 198.245 ;
        RECT 85.925 198.125 86.255 198.505 ;
        RECT 86.425 197.955 86.680 198.245 ;
        RECT 85.930 197.785 86.680 197.955 ;
        RECT 87.430 197.875 87.715 198.335 ;
        RECT 87.885 198.045 88.155 198.505 ;
        RECT 85.930 196.795 86.160 197.785 ;
        RECT 87.430 197.705 88.385 197.875 ;
        RECT 86.330 196.965 86.680 197.615 ;
        RECT 87.315 196.975 88.005 197.535 ;
        RECT 88.175 196.805 88.385 197.705 ;
        RECT 85.930 196.625 86.680 196.795 ;
        RECT 85.925 195.955 86.255 196.455 ;
        RECT 86.425 196.125 86.680 196.625 ;
        RECT 87.430 196.585 88.385 196.805 ;
        RECT 88.555 197.535 88.955 198.335 ;
        RECT 89.145 197.875 89.425 198.335 ;
        RECT 89.945 198.045 90.270 198.505 ;
        RECT 89.145 197.705 90.270 197.875 ;
        RECT 90.440 197.765 90.825 198.335 ;
        RECT 89.820 197.595 90.270 197.705 ;
        RECT 88.555 196.975 89.650 197.535 ;
        RECT 89.820 197.265 90.375 197.595 ;
        RECT 87.430 196.125 87.715 196.585 ;
        RECT 87.885 195.955 88.155 196.415 ;
        RECT 88.555 196.125 88.955 196.975 ;
        RECT 89.820 196.805 90.270 197.265 ;
        RECT 90.545 197.095 90.825 197.765 ;
        RECT 89.145 196.585 90.270 196.805 ;
        RECT 89.145 196.125 89.425 196.585 ;
        RECT 89.945 195.955 90.270 196.415 ;
        RECT 90.440 196.125 90.825 197.095 ;
        RECT 91.000 197.795 91.255 198.325 ;
        RECT 91.425 198.045 91.730 198.505 ;
        RECT 91.975 198.125 93.045 198.295 ;
        RECT 91.000 197.145 91.210 197.795 ;
        RECT 91.975 197.770 92.295 198.125 ;
        RECT 91.970 197.595 92.295 197.770 ;
        RECT 91.380 197.295 92.295 197.595 ;
        RECT 92.465 197.555 92.705 197.955 ;
        RECT 92.875 197.895 93.045 198.125 ;
        RECT 93.215 198.065 93.405 198.505 ;
        RECT 93.575 198.055 94.525 198.335 ;
        RECT 94.745 198.145 95.095 198.315 ;
        RECT 92.875 197.725 93.405 197.895 ;
        RECT 91.380 197.265 92.120 197.295 ;
        RECT 91.000 196.265 91.255 197.145 ;
        RECT 91.425 195.955 91.730 197.095 ;
        RECT 91.950 196.675 92.120 197.265 ;
        RECT 92.465 197.185 93.005 197.555 ;
        RECT 93.185 197.445 93.405 197.725 ;
        RECT 93.575 197.275 93.745 198.055 ;
        RECT 93.340 197.105 93.745 197.275 ;
        RECT 93.915 197.265 94.265 197.885 ;
        RECT 93.340 197.015 93.510 197.105 ;
        RECT 94.435 197.095 94.645 197.885 ;
        RECT 92.290 196.845 93.510 197.015 ;
        RECT 93.970 196.935 94.645 197.095 ;
        RECT 91.950 196.505 92.750 196.675 ;
        RECT 92.070 195.955 92.400 196.335 ;
        RECT 92.580 196.215 92.750 196.505 ;
        RECT 93.340 196.465 93.510 196.845 ;
        RECT 93.680 196.925 94.645 196.935 ;
        RECT 94.835 197.755 95.095 198.145 ;
        RECT 95.305 198.045 95.635 198.505 ;
        RECT 96.510 198.115 97.365 198.285 ;
        RECT 97.570 198.115 98.065 198.285 ;
        RECT 98.235 198.145 98.565 198.505 ;
        RECT 94.835 197.065 95.005 197.755 ;
        RECT 95.175 197.405 95.345 197.585 ;
        RECT 95.515 197.575 96.305 197.825 ;
        RECT 96.510 197.405 96.680 198.115 ;
        RECT 96.850 197.605 97.205 197.825 ;
        RECT 95.175 197.235 96.865 197.405 ;
        RECT 93.680 196.635 94.140 196.925 ;
        RECT 94.835 196.895 96.335 197.065 ;
        RECT 94.835 196.755 95.005 196.895 ;
        RECT 94.445 196.585 95.005 196.755 ;
        RECT 92.920 195.955 93.170 196.415 ;
        RECT 93.340 196.125 94.210 196.465 ;
        RECT 94.445 196.125 94.615 196.585 ;
        RECT 95.450 196.555 96.525 196.725 ;
        RECT 94.785 195.955 95.155 196.415 ;
        RECT 95.450 196.215 95.620 196.555 ;
        RECT 95.790 195.955 96.120 196.385 ;
        RECT 96.355 196.215 96.525 196.555 ;
        RECT 96.695 196.455 96.865 197.235 ;
        RECT 97.035 197.015 97.205 197.605 ;
        RECT 97.375 197.205 97.725 197.825 ;
        RECT 97.035 196.625 97.500 197.015 ;
        RECT 97.895 196.755 98.065 198.115 ;
        RECT 98.235 196.925 98.695 197.975 ;
        RECT 97.670 196.585 98.065 196.755 ;
        RECT 97.670 196.455 97.840 196.585 ;
        RECT 96.695 196.125 97.375 196.455 ;
        RECT 97.590 196.125 97.840 196.455 ;
        RECT 98.010 195.955 98.260 196.415 ;
        RECT 98.430 196.140 98.755 196.925 ;
        RECT 98.925 196.125 99.095 198.245 ;
        RECT 99.265 198.125 99.595 198.505 ;
        RECT 99.765 197.955 100.020 198.245 ;
        RECT 99.270 197.785 100.020 197.955 ;
        RECT 99.270 196.795 99.500 197.785 ;
        RECT 100.195 197.780 100.485 198.505 ;
        RECT 100.930 197.695 101.175 198.300 ;
        RECT 101.395 197.970 101.905 198.505 ;
        RECT 99.670 196.965 100.020 197.615 ;
        RECT 100.655 197.525 101.885 197.695 ;
        RECT 99.270 196.625 100.020 196.795 ;
        RECT 99.265 195.955 99.595 196.455 ;
        RECT 99.765 196.125 100.020 196.625 ;
        RECT 100.195 195.955 100.485 197.120 ;
        RECT 100.655 196.715 100.995 197.525 ;
        RECT 101.165 196.960 101.915 197.150 ;
        RECT 100.655 196.305 101.170 196.715 ;
        RECT 101.405 195.955 101.575 196.715 ;
        RECT 101.745 196.295 101.915 196.960 ;
        RECT 102.085 196.975 102.275 198.335 ;
        RECT 102.445 197.825 102.720 198.335 ;
        RECT 102.910 197.970 103.440 198.335 ;
        RECT 103.865 198.105 104.195 198.505 ;
        RECT 103.265 197.935 103.440 197.970 ;
        RECT 102.445 197.655 102.725 197.825 ;
        RECT 102.445 197.175 102.720 197.655 ;
        RECT 102.925 196.975 103.095 197.775 ;
        RECT 102.085 196.805 103.095 196.975 ;
        RECT 103.265 197.765 104.195 197.935 ;
        RECT 104.365 197.765 104.620 198.335 ;
        RECT 103.265 196.635 103.435 197.765 ;
        RECT 104.025 197.595 104.195 197.765 ;
        RECT 102.310 196.465 103.435 196.635 ;
        RECT 103.605 197.265 103.800 197.595 ;
        RECT 104.025 197.265 104.280 197.595 ;
        RECT 103.605 196.295 103.775 197.265 ;
        RECT 104.450 197.095 104.620 197.765 ;
        RECT 104.910 197.875 105.195 198.335 ;
        RECT 105.365 198.045 105.635 198.505 ;
        RECT 104.910 197.705 105.865 197.875 ;
        RECT 101.745 196.125 103.775 196.295 ;
        RECT 103.945 195.955 104.115 197.095 ;
        RECT 104.285 196.125 104.620 197.095 ;
        RECT 104.795 196.975 105.485 197.535 ;
        RECT 105.655 196.805 105.865 197.705 ;
        RECT 104.910 196.585 105.865 196.805 ;
        RECT 106.035 197.535 106.435 198.335 ;
        RECT 106.625 197.875 106.905 198.335 ;
        RECT 107.425 198.045 107.750 198.505 ;
        RECT 106.625 197.705 107.750 197.875 ;
        RECT 107.920 197.765 108.305 198.335 ;
        RECT 107.300 197.595 107.750 197.705 ;
        RECT 106.035 196.975 107.130 197.535 ;
        RECT 107.300 197.265 107.855 197.595 ;
        RECT 104.910 196.125 105.195 196.585 ;
        RECT 105.365 195.955 105.635 196.415 ;
        RECT 106.035 196.125 106.435 196.975 ;
        RECT 107.300 196.805 107.750 197.265 ;
        RECT 108.025 197.095 108.305 197.765 ;
        RECT 106.625 196.585 107.750 196.805 ;
        RECT 106.625 196.125 106.905 196.585 ;
        RECT 107.425 195.955 107.750 196.415 ;
        RECT 107.920 196.125 108.305 197.095 ;
        RECT 108.475 197.830 108.735 198.335 ;
        RECT 108.915 198.125 109.245 198.505 ;
        RECT 109.425 197.955 109.595 198.335 ;
        RECT 108.475 197.030 108.645 197.830 ;
        RECT 108.930 197.785 109.595 197.955 ;
        RECT 109.855 197.830 110.115 198.335 ;
        RECT 110.295 198.125 110.625 198.505 ;
        RECT 110.805 197.955 110.975 198.335 ;
        RECT 108.930 197.530 109.100 197.785 ;
        RECT 108.815 197.200 109.100 197.530 ;
        RECT 109.335 197.235 109.665 197.605 ;
        RECT 108.930 197.055 109.100 197.200 ;
        RECT 108.475 196.125 108.745 197.030 ;
        RECT 108.930 196.885 109.595 197.055 ;
        RECT 108.915 195.955 109.245 196.715 ;
        RECT 109.425 196.125 109.595 196.885 ;
        RECT 109.855 197.030 110.025 197.830 ;
        RECT 110.310 197.785 110.975 197.955 ;
        RECT 110.310 197.530 110.480 197.785 ;
        RECT 112.155 197.755 113.365 198.505 ;
        RECT 110.195 197.200 110.480 197.530 ;
        RECT 110.715 197.235 111.045 197.605 ;
        RECT 110.310 197.055 110.480 197.200 ;
        RECT 109.855 196.125 110.125 197.030 ;
        RECT 110.310 196.885 110.975 197.055 ;
        RECT 110.295 195.955 110.625 196.715 ;
        RECT 110.805 196.125 110.975 196.885 ;
        RECT 112.155 197.045 112.675 197.585 ;
        RECT 112.845 197.215 113.365 197.755 ;
        RECT 112.155 195.955 113.365 197.045 ;
        RECT 22.830 195.785 113.450 195.955 ;
        RECT 22.915 194.695 24.125 195.785 ;
        RECT 25.220 195.350 30.565 195.785 ;
        RECT 22.915 193.985 23.435 194.525 ;
        RECT 23.605 194.155 24.125 194.695 ;
        RECT 26.810 194.100 27.160 195.350 ;
        RECT 30.775 194.645 31.005 195.785 ;
        RECT 31.175 194.635 31.505 195.615 ;
        RECT 31.675 194.645 31.885 195.785 ;
        RECT 32.320 194.815 32.650 195.615 ;
        RECT 32.820 194.985 33.150 195.785 ;
        RECT 33.450 194.815 33.780 195.615 ;
        RECT 34.425 194.985 34.675 195.785 ;
        RECT 32.320 194.645 34.755 194.815 ;
        RECT 34.945 194.645 35.115 195.785 ;
        RECT 35.285 194.645 35.625 195.615 ;
        RECT 22.915 193.235 24.125 193.985 ;
        RECT 28.640 193.780 28.980 194.610 ;
        RECT 30.755 194.225 31.085 194.475 ;
        RECT 25.220 193.235 30.565 193.780 ;
        RECT 30.775 193.235 31.005 194.055 ;
        RECT 31.255 194.035 31.505 194.635 ;
        RECT 32.115 194.225 32.465 194.475 ;
        RECT 31.175 193.405 31.505 194.035 ;
        RECT 31.675 193.235 31.885 194.055 ;
        RECT 32.650 194.015 32.820 194.645 ;
        RECT 32.990 194.225 33.320 194.425 ;
        RECT 33.490 194.225 33.820 194.425 ;
        RECT 33.990 194.225 34.410 194.425 ;
        RECT 34.585 194.395 34.755 194.645 ;
        RECT 34.585 194.225 35.280 194.395 ;
        RECT 32.320 193.405 32.820 194.015 ;
        RECT 33.450 193.885 34.675 194.055 ;
        RECT 35.450 194.035 35.625 194.645 ;
        RECT 35.795 194.620 36.085 195.785 ;
        RECT 36.255 194.695 37.465 195.785 ;
        RECT 37.750 195.155 38.035 195.615 ;
        RECT 38.205 195.325 38.475 195.785 ;
        RECT 37.750 194.935 38.705 195.155 ;
        RECT 36.255 194.155 36.775 194.695 ;
        RECT 33.450 193.405 33.780 193.885 ;
        RECT 33.950 193.235 34.175 193.695 ;
        RECT 34.345 193.405 34.675 193.885 ;
        RECT 34.865 193.235 35.115 194.035 ;
        RECT 35.285 193.405 35.625 194.035 ;
        RECT 36.945 193.985 37.465 194.525 ;
        RECT 37.635 194.205 38.325 194.765 ;
        RECT 38.495 194.035 38.705 194.935 ;
        RECT 35.795 193.235 36.085 193.960 ;
        RECT 36.255 193.235 37.465 193.985 ;
        RECT 37.750 193.865 38.705 194.035 ;
        RECT 38.875 194.765 39.275 195.615 ;
        RECT 39.465 195.155 39.745 195.615 ;
        RECT 40.265 195.325 40.590 195.785 ;
        RECT 39.465 194.935 40.590 195.155 ;
        RECT 38.875 194.205 39.970 194.765 ;
        RECT 40.140 194.475 40.590 194.935 ;
        RECT 40.760 194.645 41.145 195.615 ;
        RECT 37.750 193.405 38.035 193.865 ;
        RECT 38.205 193.235 38.475 193.695 ;
        RECT 38.875 193.405 39.275 194.205 ;
        RECT 40.140 194.145 40.695 194.475 ;
        RECT 40.140 194.035 40.590 194.145 ;
        RECT 39.465 193.865 40.590 194.035 ;
        RECT 40.865 193.975 41.145 194.645 ;
        RECT 41.315 194.695 42.985 195.785 ;
        RECT 43.270 195.155 43.555 195.615 ;
        RECT 43.725 195.325 43.995 195.785 ;
        RECT 43.270 194.935 44.225 195.155 ;
        RECT 41.315 194.175 42.065 194.695 ;
        RECT 42.235 194.005 42.985 194.525 ;
        RECT 43.155 194.205 43.845 194.765 ;
        RECT 44.015 194.035 44.225 194.935 ;
        RECT 39.465 193.405 39.745 193.865 ;
        RECT 40.265 193.235 40.590 193.695 ;
        RECT 40.760 193.405 41.145 193.975 ;
        RECT 41.315 193.235 42.985 194.005 ;
        RECT 43.270 193.865 44.225 194.035 ;
        RECT 44.395 194.765 44.795 195.615 ;
        RECT 44.985 195.155 45.265 195.615 ;
        RECT 45.785 195.325 46.110 195.785 ;
        RECT 44.985 194.935 46.110 195.155 ;
        RECT 44.395 194.205 45.490 194.765 ;
        RECT 45.660 194.475 46.110 194.935 ;
        RECT 46.280 194.645 46.665 195.615 ;
        RECT 46.950 195.155 47.235 195.615 ;
        RECT 47.405 195.325 47.675 195.785 ;
        RECT 46.950 194.935 47.905 195.155 ;
        RECT 43.270 193.405 43.555 193.865 ;
        RECT 43.725 193.235 43.995 193.695 ;
        RECT 44.395 193.405 44.795 194.205 ;
        RECT 45.660 194.145 46.215 194.475 ;
        RECT 45.660 194.035 46.110 194.145 ;
        RECT 44.985 193.865 46.110 194.035 ;
        RECT 46.385 193.975 46.665 194.645 ;
        RECT 46.835 194.205 47.525 194.765 ;
        RECT 47.695 194.035 47.905 194.935 ;
        RECT 44.985 193.405 45.265 193.865 ;
        RECT 45.785 193.235 46.110 193.695 ;
        RECT 46.280 193.405 46.665 193.975 ;
        RECT 46.950 193.865 47.905 194.035 ;
        RECT 48.075 194.765 48.475 195.615 ;
        RECT 48.665 195.155 48.945 195.615 ;
        RECT 49.465 195.325 49.790 195.785 ;
        RECT 48.665 194.935 49.790 195.155 ;
        RECT 48.075 194.205 49.170 194.765 ;
        RECT 49.340 194.475 49.790 194.935 ;
        RECT 49.960 194.645 50.345 195.615 ;
        RECT 51.035 194.645 51.245 195.785 ;
        RECT 46.950 193.405 47.235 193.865 ;
        RECT 47.405 193.235 47.675 193.695 ;
        RECT 48.075 193.405 48.475 194.205 ;
        RECT 49.340 194.145 49.895 194.475 ;
        RECT 49.340 194.035 49.790 194.145 ;
        RECT 48.665 193.865 49.790 194.035 ;
        RECT 50.065 193.975 50.345 194.645 ;
        RECT 51.415 194.635 51.745 195.615 ;
        RECT 51.915 194.645 52.145 195.785 ;
        RECT 53.280 195.350 58.625 195.785 ;
        RECT 48.665 193.405 48.945 193.865 ;
        RECT 49.465 193.235 49.790 193.695 ;
        RECT 49.960 193.405 50.345 193.975 ;
        RECT 51.035 193.235 51.245 194.055 ;
        RECT 51.415 194.035 51.665 194.635 ;
        RECT 51.835 194.225 52.165 194.475 ;
        RECT 54.870 194.100 55.220 195.350 ;
        RECT 58.855 194.645 59.065 195.785 ;
        RECT 59.235 194.635 59.565 195.615 ;
        RECT 59.735 194.645 59.965 195.785 ;
        RECT 60.175 194.695 61.385 195.785 ;
        RECT 51.415 193.405 51.745 194.035 ;
        RECT 51.915 193.235 52.145 194.055 ;
        RECT 56.700 193.780 57.040 194.610 ;
        RECT 53.280 193.235 58.625 193.780 ;
        RECT 58.855 193.235 59.065 194.055 ;
        RECT 59.235 194.035 59.485 194.635 ;
        RECT 59.655 194.225 59.985 194.475 ;
        RECT 60.175 194.155 60.695 194.695 ;
        RECT 61.555 194.620 61.845 195.785 ;
        RECT 62.935 194.645 63.195 195.785 ;
        RECT 63.435 195.275 65.050 195.605 ;
        RECT 59.235 193.405 59.565 194.035 ;
        RECT 59.735 193.235 59.965 194.055 ;
        RECT 60.865 193.985 61.385 194.525 ;
        RECT 63.445 194.475 63.615 195.035 ;
        RECT 63.875 194.935 65.050 195.105 ;
        RECT 65.220 194.985 65.500 195.785 ;
        RECT 63.875 194.645 64.205 194.935 ;
        RECT 64.880 194.815 65.050 194.935 ;
        RECT 64.375 194.475 64.620 194.765 ;
        RECT 64.880 194.645 65.540 194.815 ;
        RECT 65.710 194.645 65.985 195.615 ;
        RECT 65.370 194.475 65.540 194.645 ;
        RECT 62.940 194.225 63.275 194.475 ;
        RECT 63.445 194.145 64.160 194.475 ;
        RECT 64.375 194.145 65.200 194.475 ;
        RECT 65.370 194.145 65.645 194.475 ;
        RECT 63.445 194.055 63.695 194.145 ;
        RECT 60.175 193.235 61.385 193.985 ;
        RECT 61.555 193.235 61.845 193.960 ;
        RECT 62.935 193.235 63.195 194.055 ;
        RECT 63.365 193.635 63.695 194.055 ;
        RECT 65.370 193.975 65.540 194.145 ;
        RECT 63.875 193.805 65.540 193.975 ;
        RECT 65.815 193.910 65.985 194.645 ;
        RECT 63.875 193.405 64.135 193.805 ;
        RECT 64.305 193.235 64.635 193.635 ;
        RECT 64.805 193.455 64.975 193.805 ;
        RECT 65.145 193.235 65.520 193.635 ;
        RECT 65.710 193.565 65.985 193.910 ;
        RECT 66.155 195.285 66.415 195.615 ;
        RECT 66.725 195.405 67.055 195.785 ;
        RECT 66.155 194.605 66.325 195.285 ;
        RECT 67.295 195.235 67.485 195.615 ;
        RECT 67.735 195.405 68.065 195.785 ;
        RECT 68.275 195.235 68.445 195.615 ;
        RECT 68.640 195.405 68.970 195.785 ;
        RECT 69.230 195.235 69.400 195.615 ;
        RECT 69.825 195.405 70.155 195.785 ;
        RECT 66.495 194.775 66.845 195.105 ;
        RECT 67.295 195.065 68.035 195.235 ;
        RECT 67.115 194.725 67.695 194.895 ;
        RECT 67.115 194.605 67.285 194.725 ;
        RECT 66.155 194.435 67.285 194.605 ;
        RECT 67.865 194.555 68.035 195.065 ;
        RECT 66.155 193.735 66.325 194.435 ;
        RECT 67.465 194.385 68.035 194.555 ;
        RECT 68.205 195.065 70.155 195.235 ;
        RECT 66.675 194.095 67.295 194.265 ;
        RECT 66.675 193.915 66.885 194.095 ;
        RECT 67.465 193.905 67.635 194.385 ;
        RECT 68.205 194.075 68.375 195.065 ;
        RECT 68.965 194.475 69.150 194.785 ;
        RECT 69.420 194.475 69.615 194.785 ;
        RECT 66.155 193.405 66.415 193.735 ;
        RECT 66.725 193.235 67.055 193.615 ;
        RECT 67.235 193.575 67.635 193.905 ;
        RECT 67.825 193.745 68.375 194.075 ;
        RECT 68.545 193.575 68.715 194.475 ;
        RECT 67.235 193.405 68.715 193.575 ;
        RECT 68.965 194.145 69.195 194.475 ;
        RECT 69.420 194.145 69.675 194.475 ;
        RECT 69.985 194.145 70.155 195.065 ;
        RECT 68.965 193.565 69.150 194.145 ;
        RECT 69.420 193.570 69.615 194.145 ;
        RECT 69.825 193.235 70.155 193.615 ;
        RECT 70.325 193.405 70.585 195.615 ;
        RECT 70.760 194.595 71.015 195.475 ;
        RECT 71.185 194.645 71.490 195.785 ;
        RECT 71.830 195.405 72.160 195.785 ;
        RECT 72.340 195.235 72.510 195.525 ;
        RECT 72.680 195.325 72.930 195.785 ;
        RECT 71.710 195.065 72.510 195.235 ;
        RECT 73.100 195.275 73.970 195.615 ;
        RECT 70.760 193.945 70.970 194.595 ;
        RECT 71.710 194.475 71.880 195.065 ;
        RECT 73.100 194.895 73.270 195.275 ;
        RECT 74.205 195.155 74.375 195.615 ;
        RECT 74.545 195.325 74.915 195.785 ;
        RECT 75.210 195.185 75.380 195.525 ;
        RECT 75.550 195.355 75.880 195.785 ;
        RECT 76.115 195.185 76.285 195.525 ;
        RECT 72.050 194.725 73.270 194.895 ;
        RECT 73.440 194.815 73.900 195.105 ;
        RECT 74.205 194.985 74.765 195.155 ;
        RECT 75.210 195.015 76.285 195.185 ;
        RECT 76.455 195.285 77.135 195.615 ;
        RECT 77.350 195.285 77.600 195.615 ;
        RECT 77.770 195.325 78.020 195.785 ;
        RECT 74.595 194.845 74.765 194.985 ;
        RECT 73.440 194.805 74.405 194.815 ;
        RECT 73.100 194.635 73.270 194.725 ;
        RECT 73.730 194.645 74.405 194.805 ;
        RECT 71.140 194.445 71.880 194.475 ;
        RECT 71.140 194.145 72.055 194.445 ;
        RECT 71.730 193.970 72.055 194.145 ;
        RECT 70.760 193.415 71.015 193.945 ;
        RECT 71.185 193.235 71.490 193.695 ;
        RECT 71.735 193.615 72.055 193.970 ;
        RECT 72.225 194.185 72.765 194.555 ;
        RECT 73.100 194.465 73.505 194.635 ;
        RECT 72.225 193.785 72.465 194.185 ;
        RECT 72.945 194.015 73.165 194.295 ;
        RECT 72.635 193.845 73.165 194.015 ;
        RECT 72.635 193.615 72.805 193.845 ;
        RECT 73.335 193.685 73.505 194.465 ;
        RECT 73.675 193.855 74.025 194.475 ;
        RECT 74.195 193.855 74.405 194.645 ;
        RECT 74.595 194.675 76.095 194.845 ;
        RECT 74.595 193.985 74.765 194.675 ;
        RECT 76.455 194.505 76.625 195.285 ;
        RECT 77.430 195.155 77.600 195.285 ;
        RECT 74.935 194.335 76.625 194.505 ;
        RECT 76.795 194.725 77.260 195.115 ;
        RECT 77.430 194.985 77.825 195.155 ;
        RECT 74.935 194.155 75.105 194.335 ;
        RECT 71.735 193.445 72.805 193.615 ;
        RECT 72.975 193.235 73.165 193.675 ;
        RECT 73.335 193.405 74.285 193.685 ;
        RECT 74.595 193.595 74.855 193.985 ;
        RECT 75.275 193.915 76.065 194.165 ;
        RECT 74.505 193.425 74.855 193.595 ;
        RECT 75.065 193.235 75.395 193.695 ;
        RECT 76.270 193.625 76.440 194.335 ;
        RECT 76.795 194.135 76.965 194.725 ;
        RECT 76.610 193.915 76.965 194.135 ;
        RECT 77.135 193.915 77.485 194.535 ;
        RECT 77.655 193.625 77.825 194.985 ;
        RECT 78.190 194.815 78.515 195.600 ;
        RECT 77.995 193.765 78.455 194.815 ;
        RECT 76.270 193.455 77.125 193.625 ;
        RECT 77.330 193.455 77.825 193.625 ;
        RECT 77.995 193.235 78.325 193.595 ;
        RECT 78.685 193.495 78.855 195.615 ;
        RECT 79.025 195.285 79.355 195.785 ;
        RECT 79.525 195.115 79.780 195.615 ;
        RECT 79.030 194.945 79.780 195.115 ;
        RECT 79.030 193.955 79.260 194.945 ;
        RECT 79.430 194.125 79.780 194.775 ;
        RECT 79.955 194.645 80.215 195.785 ;
        RECT 80.385 194.635 80.715 195.615 ;
        RECT 80.885 194.645 81.165 195.785 ;
        RECT 81.395 194.645 81.605 195.785 ;
        RECT 81.775 194.635 82.105 195.615 ;
        RECT 82.275 194.645 82.505 195.785 ;
        RECT 83.750 195.155 84.035 195.615 ;
        RECT 84.205 195.325 84.475 195.785 ;
        RECT 83.750 194.935 84.705 195.155 ;
        RECT 79.975 194.225 80.310 194.475 ;
        RECT 80.480 194.035 80.650 194.635 ;
        RECT 80.820 194.205 81.155 194.475 ;
        RECT 79.030 193.785 79.780 193.955 ;
        RECT 79.025 193.235 79.355 193.615 ;
        RECT 79.525 193.495 79.780 193.785 ;
        RECT 79.955 193.405 80.650 194.035 ;
        RECT 80.855 193.235 81.165 194.035 ;
        RECT 81.395 193.235 81.605 194.055 ;
        RECT 81.775 194.035 82.025 194.635 ;
        RECT 82.195 194.225 82.525 194.475 ;
        RECT 83.635 194.205 84.325 194.765 ;
        RECT 81.775 193.405 82.105 194.035 ;
        RECT 82.275 193.235 82.505 194.055 ;
        RECT 84.495 194.035 84.705 194.935 ;
        RECT 83.750 193.865 84.705 194.035 ;
        RECT 84.875 194.765 85.275 195.615 ;
        RECT 85.465 195.155 85.745 195.615 ;
        RECT 86.265 195.325 86.590 195.785 ;
        RECT 85.465 194.935 86.590 195.155 ;
        RECT 84.875 194.205 85.970 194.765 ;
        RECT 86.140 194.475 86.590 194.935 ;
        RECT 86.760 194.645 87.145 195.615 ;
        RECT 83.750 193.405 84.035 193.865 ;
        RECT 84.205 193.235 84.475 193.695 ;
        RECT 84.875 193.405 85.275 194.205 ;
        RECT 86.140 194.145 86.695 194.475 ;
        RECT 86.140 194.035 86.590 194.145 ;
        RECT 85.465 193.865 86.590 194.035 ;
        RECT 86.865 193.975 87.145 194.645 ;
        RECT 87.315 194.620 87.605 195.785 ;
        RECT 85.465 193.405 85.745 193.865 ;
        RECT 86.265 193.235 86.590 193.695 ;
        RECT 86.760 193.405 87.145 193.975 ;
        RECT 87.780 194.595 88.035 195.475 ;
        RECT 88.205 194.645 88.510 195.785 ;
        RECT 88.850 195.405 89.180 195.785 ;
        RECT 89.360 195.235 89.530 195.525 ;
        RECT 89.700 195.325 89.950 195.785 ;
        RECT 88.730 195.065 89.530 195.235 ;
        RECT 90.120 195.275 90.990 195.615 ;
        RECT 87.315 193.235 87.605 193.960 ;
        RECT 87.780 193.945 87.990 194.595 ;
        RECT 88.730 194.475 88.900 195.065 ;
        RECT 90.120 194.895 90.290 195.275 ;
        RECT 91.225 195.155 91.395 195.615 ;
        RECT 91.565 195.325 91.935 195.785 ;
        RECT 92.230 195.185 92.400 195.525 ;
        RECT 92.570 195.355 92.900 195.785 ;
        RECT 93.135 195.185 93.305 195.525 ;
        RECT 89.070 194.725 90.290 194.895 ;
        RECT 90.460 194.815 90.920 195.105 ;
        RECT 91.225 194.985 91.785 195.155 ;
        RECT 92.230 195.015 93.305 195.185 ;
        RECT 93.475 195.285 94.155 195.615 ;
        RECT 94.370 195.285 94.620 195.615 ;
        RECT 94.790 195.325 95.040 195.785 ;
        RECT 91.615 194.845 91.785 194.985 ;
        RECT 90.460 194.805 91.425 194.815 ;
        RECT 90.120 194.635 90.290 194.725 ;
        RECT 90.750 194.645 91.425 194.805 ;
        RECT 88.160 194.445 88.900 194.475 ;
        RECT 88.160 194.145 89.075 194.445 ;
        RECT 88.750 193.970 89.075 194.145 ;
        RECT 87.780 193.415 88.035 193.945 ;
        RECT 88.205 193.235 88.510 193.695 ;
        RECT 88.755 193.615 89.075 193.970 ;
        RECT 89.245 194.185 89.785 194.555 ;
        RECT 90.120 194.465 90.525 194.635 ;
        RECT 89.245 193.785 89.485 194.185 ;
        RECT 89.965 194.015 90.185 194.295 ;
        RECT 89.655 193.845 90.185 194.015 ;
        RECT 89.655 193.615 89.825 193.845 ;
        RECT 90.355 193.685 90.525 194.465 ;
        RECT 90.695 193.855 91.045 194.475 ;
        RECT 91.215 193.855 91.425 194.645 ;
        RECT 91.615 194.675 93.115 194.845 ;
        RECT 91.615 193.985 91.785 194.675 ;
        RECT 93.475 194.505 93.645 195.285 ;
        RECT 94.450 195.155 94.620 195.285 ;
        RECT 91.955 194.335 93.645 194.505 ;
        RECT 93.815 194.725 94.280 195.115 ;
        RECT 94.450 194.985 94.845 195.155 ;
        RECT 91.955 194.155 92.125 194.335 ;
        RECT 88.755 193.445 89.825 193.615 ;
        RECT 89.995 193.235 90.185 193.675 ;
        RECT 90.355 193.405 91.305 193.685 ;
        RECT 91.615 193.595 91.875 193.985 ;
        RECT 92.295 193.915 93.085 194.165 ;
        RECT 91.525 193.425 91.875 193.595 ;
        RECT 92.085 193.235 92.415 193.695 ;
        RECT 93.290 193.625 93.460 194.335 ;
        RECT 93.815 194.135 93.985 194.725 ;
        RECT 93.630 193.915 93.985 194.135 ;
        RECT 94.155 193.915 94.505 194.535 ;
        RECT 94.675 193.625 94.845 194.985 ;
        RECT 95.210 194.815 95.535 195.600 ;
        RECT 95.015 193.765 95.475 194.815 ;
        RECT 93.290 193.455 94.145 193.625 ;
        RECT 94.350 193.455 94.845 193.625 ;
        RECT 95.015 193.235 95.345 193.595 ;
        RECT 95.705 193.495 95.875 195.615 ;
        RECT 96.045 195.285 96.375 195.785 ;
        RECT 96.545 195.115 96.800 195.615 ;
        RECT 96.050 194.945 96.800 195.115 ;
        RECT 97.090 195.155 97.375 195.615 ;
        RECT 97.545 195.325 97.815 195.785 ;
        RECT 96.050 193.955 96.280 194.945 ;
        RECT 97.090 194.935 98.045 195.155 ;
        RECT 96.450 194.125 96.800 194.775 ;
        RECT 96.975 194.205 97.665 194.765 ;
        RECT 97.835 194.035 98.045 194.935 ;
        RECT 96.050 193.785 96.800 193.955 ;
        RECT 96.045 193.235 96.375 193.615 ;
        RECT 96.545 193.495 96.800 193.785 ;
        RECT 97.090 193.865 98.045 194.035 ;
        RECT 98.215 194.765 98.615 195.615 ;
        RECT 98.805 195.155 99.085 195.615 ;
        RECT 99.605 195.325 99.930 195.785 ;
        RECT 98.805 194.935 99.930 195.155 ;
        RECT 98.215 194.205 99.310 194.765 ;
        RECT 99.480 194.475 99.930 194.935 ;
        RECT 100.100 194.645 100.485 195.615 ;
        RECT 100.660 195.115 100.915 195.615 ;
        RECT 101.085 195.285 101.415 195.785 ;
        RECT 100.660 194.945 101.410 195.115 ;
        RECT 97.090 193.405 97.375 193.865 ;
        RECT 97.545 193.235 97.815 193.695 ;
        RECT 98.215 193.405 98.615 194.205 ;
        RECT 99.480 194.145 100.035 194.475 ;
        RECT 99.480 194.035 99.930 194.145 ;
        RECT 98.805 193.865 99.930 194.035 ;
        RECT 100.205 193.975 100.485 194.645 ;
        RECT 100.660 194.125 101.010 194.775 ;
        RECT 98.805 193.405 99.085 193.865 ;
        RECT 99.605 193.235 99.930 193.695 ;
        RECT 100.100 193.405 100.485 193.975 ;
        RECT 101.180 193.955 101.410 194.945 ;
        RECT 100.660 193.785 101.410 193.955 ;
        RECT 100.660 193.495 100.915 193.785 ;
        RECT 101.085 193.235 101.415 193.615 ;
        RECT 101.585 193.495 101.755 195.615 ;
        RECT 101.925 194.815 102.250 195.600 ;
        RECT 102.420 195.325 102.670 195.785 ;
        RECT 102.840 195.285 103.090 195.615 ;
        RECT 103.305 195.285 103.985 195.615 ;
        RECT 102.840 195.155 103.010 195.285 ;
        RECT 102.615 194.985 103.010 195.155 ;
        RECT 101.985 193.765 102.445 194.815 ;
        RECT 102.615 193.625 102.785 194.985 ;
        RECT 103.180 194.725 103.645 195.115 ;
        RECT 102.955 193.915 103.305 194.535 ;
        RECT 103.475 194.135 103.645 194.725 ;
        RECT 103.815 194.505 103.985 195.285 ;
        RECT 104.155 195.185 104.325 195.525 ;
        RECT 104.560 195.355 104.890 195.785 ;
        RECT 105.060 195.185 105.230 195.525 ;
        RECT 105.525 195.325 105.895 195.785 ;
        RECT 104.155 195.015 105.230 195.185 ;
        RECT 106.065 195.155 106.235 195.615 ;
        RECT 106.470 195.275 107.340 195.615 ;
        RECT 107.510 195.325 107.760 195.785 ;
        RECT 105.675 194.985 106.235 195.155 ;
        RECT 105.675 194.845 105.845 194.985 ;
        RECT 104.345 194.675 105.845 194.845 ;
        RECT 106.540 194.815 107.000 195.105 ;
        RECT 103.815 194.335 105.505 194.505 ;
        RECT 103.475 193.915 103.830 194.135 ;
        RECT 104.000 193.625 104.170 194.335 ;
        RECT 104.375 193.915 105.165 194.165 ;
        RECT 105.335 194.155 105.505 194.335 ;
        RECT 105.675 193.985 105.845 194.675 ;
        RECT 102.115 193.235 102.445 193.595 ;
        RECT 102.615 193.455 103.110 193.625 ;
        RECT 103.315 193.455 104.170 193.625 ;
        RECT 105.045 193.235 105.375 193.695 ;
        RECT 105.585 193.595 105.845 193.985 ;
        RECT 106.035 194.805 107.000 194.815 ;
        RECT 107.170 194.895 107.340 195.275 ;
        RECT 107.930 195.235 108.100 195.525 ;
        RECT 108.280 195.405 108.610 195.785 ;
        RECT 107.930 195.065 108.730 195.235 ;
        RECT 106.035 194.645 106.710 194.805 ;
        RECT 107.170 194.725 108.390 194.895 ;
        RECT 106.035 193.855 106.245 194.645 ;
        RECT 107.170 194.635 107.340 194.725 ;
        RECT 106.415 193.855 106.765 194.475 ;
        RECT 106.935 194.465 107.340 194.635 ;
        RECT 106.935 193.685 107.105 194.465 ;
        RECT 107.275 194.015 107.495 194.295 ;
        RECT 107.675 194.185 108.215 194.555 ;
        RECT 108.560 194.475 108.730 195.065 ;
        RECT 108.950 194.645 109.255 195.785 ;
        RECT 109.425 194.595 109.680 195.475 ;
        RECT 109.895 194.645 110.125 195.785 ;
        RECT 110.295 194.635 110.625 195.615 ;
        RECT 110.795 194.645 111.005 195.785 ;
        RECT 112.155 194.695 113.365 195.785 ;
        RECT 108.560 194.445 109.300 194.475 ;
        RECT 107.275 193.845 107.805 194.015 ;
        RECT 105.585 193.425 105.935 193.595 ;
        RECT 106.155 193.405 107.105 193.685 ;
        RECT 107.275 193.235 107.465 193.675 ;
        RECT 107.635 193.615 107.805 193.845 ;
        RECT 107.975 193.785 108.215 194.185 ;
        RECT 108.385 194.145 109.300 194.445 ;
        RECT 108.385 193.970 108.710 194.145 ;
        RECT 108.385 193.615 108.705 193.970 ;
        RECT 109.470 193.945 109.680 194.595 ;
        RECT 109.875 194.225 110.205 194.475 ;
        RECT 107.635 193.445 108.705 193.615 ;
        RECT 108.950 193.235 109.255 193.695 ;
        RECT 109.425 193.415 109.680 193.945 ;
        RECT 109.895 193.235 110.125 194.055 ;
        RECT 110.375 194.035 110.625 194.635 ;
        RECT 112.155 194.155 112.675 194.695 ;
        RECT 110.295 193.405 110.625 194.035 ;
        RECT 110.795 193.235 111.005 194.055 ;
        RECT 112.845 193.985 113.365 194.525 ;
        RECT 112.155 193.235 113.365 193.985 ;
        RECT 22.830 193.065 113.450 193.235 ;
        RECT 22.915 192.315 24.125 193.065 ;
        RECT 24.295 192.315 25.505 193.065 ;
        RECT 22.915 191.775 23.435 192.315 ;
        RECT 23.605 191.605 24.125 192.145 ;
        RECT 22.915 190.515 24.125 191.605 ;
        RECT 24.295 191.605 24.815 192.145 ;
        RECT 24.985 191.775 25.505 192.315 ;
        RECT 25.675 192.295 29.185 193.065 ;
        RECT 25.675 191.605 27.365 192.125 ;
        RECT 27.535 191.775 29.185 192.295 ;
        RECT 29.415 192.245 29.625 193.065 ;
        RECT 29.795 192.265 30.125 192.895 ;
        RECT 29.795 191.665 30.045 192.265 ;
        RECT 30.295 192.245 30.525 193.065 ;
        RECT 30.825 192.515 30.995 192.895 ;
        RECT 31.175 192.685 31.505 193.065 ;
        RECT 30.825 192.345 31.490 192.515 ;
        RECT 31.685 192.390 31.945 192.895 ;
        RECT 30.215 191.825 30.545 192.075 ;
        RECT 30.755 191.795 31.085 192.165 ;
        RECT 31.320 192.090 31.490 192.345 ;
        RECT 31.320 191.760 31.605 192.090 ;
        RECT 24.295 190.515 25.505 191.605 ;
        RECT 25.675 190.515 29.185 191.605 ;
        RECT 29.415 190.515 29.625 191.655 ;
        RECT 29.795 190.685 30.125 191.665 ;
        RECT 30.295 190.515 30.525 191.655 ;
        RECT 31.320 191.615 31.490 191.760 ;
        RECT 30.825 191.445 31.490 191.615 ;
        RECT 31.775 191.590 31.945 192.390 ;
        RECT 32.230 192.435 32.515 192.895 ;
        RECT 32.685 192.605 32.955 193.065 ;
        RECT 32.230 192.265 33.185 192.435 ;
        RECT 30.825 190.685 30.995 191.445 ;
        RECT 31.175 190.515 31.505 191.275 ;
        RECT 31.675 190.685 31.945 191.590 ;
        RECT 32.115 191.535 32.805 192.095 ;
        RECT 32.975 191.365 33.185 192.265 ;
        RECT 32.230 191.145 33.185 191.365 ;
        RECT 33.355 192.095 33.755 192.895 ;
        RECT 33.945 192.435 34.225 192.895 ;
        RECT 34.745 192.605 35.070 193.065 ;
        RECT 33.945 192.265 35.070 192.435 ;
        RECT 35.240 192.325 35.625 192.895 ;
        RECT 34.620 192.155 35.070 192.265 ;
        RECT 33.355 191.535 34.450 192.095 ;
        RECT 34.620 191.825 35.175 192.155 ;
        RECT 32.230 190.685 32.515 191.145 ;
        RECT 32.685 190.515 32.955 190.975 ;
        RECT 33.355 190.685 33.755 191.535 ;
        RECT 34.620 191.365 35.070 191.825 ;
        RECT 35.345 191.655 35.625 192.325 ;
        RECT 33.945 191.145 35.070 191.365 ;
        RECT 33.945 190.685 34.225 191.145 ;
        RECT 34.745 190.515 35.070 190.975 ;
        RECT 35.240 190.685 35.625 191.655 ;
        RECT 35.795 192.265 36.135 192.895 ;
        RECT 36.305 192.265 36.555 193.065 ;
        RECT 36.745 192.415 37.075 192.895 ;
        RECT 37.245 192.605 37.470 193.065 ;
        RECT 37.640 192.415 37.970 192.895 ;
        RECT 35.795 191.655 35.970 192.265 ;
        RECT 36.745 192.245 37.970 192.415 ;
        RECT 38.600 192.285 39.100 192.895 ;
        RECT 39.480 192.355 39.735 192.885 ;
        RECT 39.905 192.605 40.210 193.065 ;
        RECT 40.455 192.685 41.525 192.855 ;
        RECT 36.140 191.905 36.835 192.075 ;
        RECT 36.665 191.655 36.835 191.905 ;
        RECT 37.010 191.875 37.430 192.075 ;
        RECT 37.600 191.875 37.930 192.075 ;
        RECT 38.100 191.875 38.430 192.075 ;
        RECT 38.600 191.655 38.770 192.285 ;
        RECT 38.955 191.825 39.305 192.075 ;
        RECT 39.480 191.705 39.690 192.355 ;
        RECT 40.455 192.330 40.775 192.685 ;
        RECT 40.450 192.155 40.775 192.330 ;
        RECT 39.860 191.855 40.775 192.155 ;
        RECT 40.945 192.115 41.185 192.515 ;
        RECT 41.355 192.455 41.525 192.685 ;
        RECT 41.695 192.625 41.885 193.065 ;
        RECT 42.055 192.615 43.005 192.895 ;
        RECT 43.225 192.705 43.575 192.875 ;
        RECT 41.355 192.285 41.885 192.455 ;
        RECT 39.860 191.825 40.600 191.855 ;
        RECT 35.795 190.685 36.135 191.655 ;
        RECT 36.305 190.515 36.475 191.655 ;
        RECT 36.665 191.485 39.100 191.655 ;
        RECT 36.745 190.515 36.995 191.315 ;
        RECT 37.640 190.685 37.970 191.485 ;
        RECT 38.270 190.515 38.600 191.315 ;
        RECT 38.770 190.685 39.100 191.485 ;
        RECT 39.480 190.825 39.735 191.705 ;
        RECT 39.905 190.515 40.210 191.655 ;
        RECT 40.430 191.235 40.600 191.825 ;
        RECT 40.945 191.745 41.485 192.115 ;
        RECT 41.665 192.005 41.885 192.285 ;
        RECT 42.055 191.835 42.225 192.615 ;
        RECT 41.820 191.665 42.225 191.835 ;
        RECT 42.395 191.825 42.745 192.445 ;
        RECT 41.820 191.575 41.990 191.665 ;
        RECT 42.915 191.655 43.125 192.445 ;
        RECT 40.770 191.405 41.990 191.575 ;
        RECT 42.450 191.495 43.125 191.655 ;
        RECT 40.430 191.065 41.230 191.235 ;
        RECT 40.550 190.515 40.880 190.895 ;
        RECT 41.060 190.775 41.230 191.065 ;
        RECT 41.820 191.025 41.990 191.405 ;
        RECT 42.160 191.485 43.125 191.495 ;
        RECT 43.315 192.315 43.575 192.705 ;
        RECT 43.785 192.605 44.115 193.065 ;
        RECT 44.990 192.675 45.845 192.845 ;
        RECT 46.050 192.675 46.545 192.845 ;
        RECT 46.715 192.705 47.045 193.065 ;
        RECT 43.315 191.625 43.485 192.315 ;
        RECT 43.655 191.965 43.825 192.145 ;
        RECT 43.995 192.135 44.785 192.385 ;
        RECT 44.990 191.965 45.160 192.675 ;
        RECT 45.330 192.165 45.685 192.385 ;
        RECT 43.655 191.795 45.345 191.965 ;
        RECT 42.160 191.195 42.620 191.485 ;
        RECT 43.315 191.455 44.815 191.625 ;
        RECT 43.315 191.315 43.485 191.455 ;
        RECT 42.925 191.145 43.485 191.315 ;
        RECT 41.400 190.515 41.650 190.975 ;
        RECT 41.820 190.685 42.690 191.025 ;
        RECT 42.925 190.685 43.095 191.145 ;
        RECT 43.930 191.115 45.005 191.285 ;
        RECT 43.265 190.515 43.635 190.975 ;
        RECT 43.930 190.775 44.100 191.115 ;
        RECT 44.270 190.515 44.600 190.945 ;
        RECT 44.835 190.775 45.005 191.115 ;
        RECT 45.175 191.015 45.345 191.795 ;
        RECT 45.515 191.575 45.685 192.165 ;
        RECT 45.855 191.765 46.205 192.385 ;
        RECT 45.515 191.185 45.980 191.575 ;
        RECT 46.375 191.315 46.545 192.675 ;
        RECT 46.715 191.485 47.175 192.535 ;
        RECT 46.150 191.145 46.545 191.315 ;
        RECT 46.150 191.015 46.320 191.145 ;
        RECT 45.175 190.685 45.855 191.015 ;
        RECT 46.070 190.685 46.320 191.015 ;
        RECT 46.490 190.515 46.740 190.975 ;
        RECT 46.910 190.700 47.235 191.485 ;
        RECT 47.405 190.685 47.575 192.805 ;
        RECT 47.745 192.685 48.075 193.065 ;
        RECT 48.245 192.515 48.500 192.805 ;
        RECT 47.750 192.345 48.500 192.515 ;
        RECT 47.750 191.355 47.980 192.345 ;
        RECT 48.675 192.340 48.965 193.065 ;
        RECT 50.055 192.390 50.315 192.895 ;
        RECT 50.495 192.685 50.825 193.065 ;
        RECT 51.005 192.515 51.175 192.895 ;
        RECT 48.150 191.525 48.500 192.175 ;
        RECT 47.750 191.185 48.500 191.355 ;
        RECT 47.745 190.515 48.075 191.015 ;
        RECT 48.245 190.685 48.500 191.185 ;
        RECT 48.675 190.515 48.965 191.680 ;
        RECT 50.055 191.590 50.225 192.390 ;
        RECT 50.510 192.345 51.175 192.515 ;
        RECT 51.550 192.435 51.835 192.895 ;
        RECT 52.005 192.605 52.275 193.065 ;
        RECT 50.510 192.090 50.680 192.345 ;
        RECT 51.550 192.265 52.505 192.435 ;
        RECT 50.395 191.760 50.680 192.090 ;
        RECT 50.915 191.795 51.245 192.165 ;
        RECT 50.510 191.615 50.680 191.760 ;
        RECT 50.055 190.685 50.325 191.590 ;
        RECT 50.510 191.445 51.175 191.615 ;
        RECT 51.435 191.535 52.125 192.095 ;
        RECT 50.495 190.515 50.825 191.275 ;
        RECT 51.005 190.685 51.175 191.445 ;
        RECT 52.295 191.365 52.505 192.265 ;
        RECT 51.550 191.145 52.505 191.365 ;
        RECT 52.675 192.095 53.075 192.895 ;
        RECT 53.265 192.435 53.545 192.895 ;
        RECT 54.065 192.605 54.390 193.065 ;
        RECT 53.265 192.265 54.390 192.435 ;
        RECT 54.560 192.325 54.945 192.895 ;
        RECT 53.940 192.155 54.390 192.265 ;
        RECT 52.675 191.535 53.770 192.095 ;
        RECT 53.940 191.825 54.495 192.155 ;
        RECT 51.550 190.685 51.835 191.145 ;
        RECT 52.005 190.515 52.275 190.975 ;
        RECT 52.675 190.685 53.075 191.535 ;
        RECT 53.940 191.365 54.390 191.825 ;
        RECT 54.665 191.655 54.945 192.325 ;
        RECT 55.175 192.245 55.385 193.065 ;
        RECT 55.555 192.265 55.885 192.895 ;
        RECT 55.555 191.665 55.805 192.265 ;
        RECT 56.055 192.245 56.285 193.065 ;
        RECT 57.420 192.520 62.765 193.065 ;
        RECT 62.940 192.520 68.285 193.065 ;
        RECT 68.460 192.665 68.795 193.065 ;
        RECT 55.975 191.825 56.305 192.075 ;
        RECT 53.265 191.145 54.390 191.365 ;
        RECT 53.265 190.685 53.545 191.145 ;
        RECT 54.065 190.515 54.390 190.975 ;
        RECT 54.560 190.685 54.945 191.655 ;
        RECT 55.175 190.515 55.385 191.655 ;
        RECT 55.555 190.685 55.885 191.665 ;
        RECT 56.055 190.515 56.285 191.655 ;
        RECT 59.010 190.950 59.360 192.200 ;
        RECT 60.840 191.690 61.180 192.520 ;
        RECT 64.530 190.950 64.880 192.200 ;
        RECT 66.360 191.690 66.700 192.520 ;
        RECT 68.965 192.495 69.170 192.895 ;
        RECT 69.380 192.585 69.655 193.065 ;
        RECT 69.865 192.565 70.125 192.895 ;
        RECT 68.485 192.325 69.170 192.495 ;
        RECT 68.485 191.295 68.825 192.325 ;
        RECT 68.995 191.655 69.245 192.155 ;
        RECT 69.425 191.825 69.785 192.405 ;
        RECT 69.955 191.655 70.125 192.565 ;
        RECT 70.755 192.295 72.425 193.065 ;
        RECT 68.995 191.485 70.125 191.655 ;
        RECT 68.485 191.120 69.150 191.295 ;
        RECT 57.420 190.515 62.765 190.950 ;
        RECT 62.940 190.515 68.285 190.950 ;
        RECT 68.460 190.515 68.795 190.940 ;
        RECT 68.965 190.715 69.150 191.120 ;
        RECT 69.355 190.515 69.685 191.295 ;
        RECT 69.855 190.715 70.125 191.485 ;
        RECT 70.755 191.605 71.505 192.125 ;
        RECT 71.675 191.775 72.425 192.295 ;
        RECT 72.595 192.565 72.855 192.895 ;
        RECT 73.065 192.585 73.340 193.065 ;
        RECT 72.595 191.655 72.765 192.565 ;
        RECT 73.550 192.495 73.755 192.895 ;
        RECT 73.925 192.665 74.260 193.065 ;
        RECT 72.935 191.825 73.295 192.405 ;
        RECT 73.550 192.325 74.235 192.495 ;
        RECT 74.435 192.340 74.725 193.065 ;
        RECT 74.985 192.415 75.155 192.895 ;
        RECT 75.335 192.585 75.575 193.065 ;
        RECT 75.825 192.415 75.995 192.895 ;
        RECT 76.165 192.585 76.495 193.065 ;
        RECT 76.665 192.415 76.835 192.895 ;
        RECT 73.475 191.655 73.725 192.155 ;
        RECT 70.755 190.515 72.425 191.605 ;
        RECT 72.595 191.485 73.725 191.655 ;
        RECT 72.595 190.715 72.865 191.485 ;
        RECT 73.895 191.295 74.235 192.325 ;
        RECT 74.985 192.245 75.620 192.415 ;
        RECT 75.825 192.245 76.835 192.415 ;
        RECT 77.005 192.265 77.335 193.065 ;
        RECT 77.690 192.325 78.305 192.895 ;
        RECT 78.475 192.555 78.690 193.065 ;
        RECT 78.920 192.555 79.200 192.885 ;
        RECT 79.380 192.555 79.620 193.065 ;
        RECT 75.450 192.075 75.620 192.245 ;
        RECT 76.335 192.215 76.835 192.245 ;
        RECT 74.900 191.835 75.280 192.075 ;
        RECT 75.450 191.905 75.950 192.075 ;
        RECT 73.035 190.515 73.365 191.295 ;
        RECT 73.570 191.120 74.235 191.295 ;
        RECT 73.570 190.715 73.755 191.120 ;
        RECT 73.925 190.515 74.260 190.940 ;
        RECT 74.435 190.515 74.725 191.680 ;
        RECT 75.450 191.665 75.620 191.905 ;
        RECT 76.340 191.705 76.835 192.215 ;
        RECT 74.905 191.495 75.620 191.665 ;
        RECT 75.825 191.535 76.835 191.705 ;
        RECT 74.905 190.685 75.235 191.495 ;
        RECT 75.405 190.515 75.645 191.315 ;
        RECT 75.825 190.685 75.995 191.535 ;
        RECT 76.165 190.515 76.495 191.315 ;
        RECT 76.665 190.685 76.835 191.535 ;
        RECT 77.005 190.515 77.335 191.665 ;
        RECT 77.690 191.305 78.005 192.325 ;
        RECT 78.175 191.655 78.345 192.155 ;
        RECT 78.595 191.825 78.860 192.385 ;
        RECT 79.030 191.655 79.200 192.555 ;
        RECT 79.370 191.825 79.725 192.385 ;
        RECT 81.150 192.255 81.395 192.860 ;
        RECT 81.615 192.530 82.125 193.065 ;
        RECT 80.875 192.085 82.105 192.255 ;
        RECT 78.175 191.485 79.600 191.655 ;
        RECT 77.690 190.685 78.225 191.305 ;
        RECT 78.395 190.515 78.725 191.315 ;
        RECT 79.210 191.310 79.600 191.485 ;
        RECT 80.875 191.275 81.215 192.085 ;
        RECT 81.385 191.520 82.135 191.710 ;
        RECT 80.875 190.865 81.390 191.275 ;
        RECT 81.625 190.515 81.795 191.275 ;
        RECT 81.965 190.855 82.135 191.520 ;
        RECT 82.305 191.535 82.495 192.895 ;
        RECT 82.665 192.045 82.940 192.895 ;
        RECT 83.130 192.530 83.660 192.895 ;
        RECT 84.085 192.665 84.415 193.065 ;
        RECT 83.485 192.495 83.660 192.530 ;
        RECT 82.665 191.875 82.945 192.045 ;
        RECT 82.665 191.735 82.940 191.875 ;
        RECT 83.145 191.535 83.315 192.335 ;
        RECT 82.305 191.365 83.315 191.535 ;
        RECT 83.485 192.325 84.415 192.495 ;
        RECT 84.585 192.325 84.840 192.895 ;
        RECT 83.485 191.195 83.655 192.325 ;
        RECT 84.245 192.155 84.415 192.325 ;
        RECT 82.530 191.025 83.655 191.195 ;
        RECT 83.825 191.825 84.020 192.155 ;
        RECT 84.245 191.825 84.500 192.155 ;
        RECT 83.825 190.855 83.995 191.825 ;
        RECT 84.670 191.655 84.840 192.325 ;
        RECT 81.965 190.685 83.995 190.855 ;
        RECT 84.165 190.515 84.335 191.655 ;
        RECT 84.505 190.685 84.840 191.655 ;
        RECT 85.475 192.390 85.735 192.895 ;
        RECT 85.915 192.685 86.245 193.065 ;
        RECT 86.425 192.515 86.595 192.895 ;
        RECT 85.475 191.590 85.645 192.390 ;
        RECT 85.930 192.345 86.595 192.515 ;
        RECT 85.930 192.090 86.100 192.345 ;
        RECT 86.915 192.245 87.125 193.065 ;
        RECT 87.295 192.265 87.625 192.895 ;
        RECT 85.815 191.760 86.100 192.090 ;
        RECT 86.335 191.795 86.665 192.165 ;
        RECT 85.930 191.615 86.100 191.760 ;
        RECT 87.295 191.665 87.545 192.265 ;
        RECT 87.795 192.245 88.025 193.065 ;
        RECT 88.510 192.255 88.755 192.860 ;
        RECT 88.975 192.530 89.485 193.065 ;
        RECT 88.235 192.085 89.465 192.255 ;
        RECT 87.715 191.825 88.045 192.075 ;
        RECT 85.475 190.685 85.745 191.590 ;
        RECT 85.930 191.445 86.595 191.615 ;
        RECT 85.915 190.515 86.245 191.275 ;
        RECT 86.425 190.685 86.595 191.445 ;
        RECT 86.915 190.515 87.125 191.655 ;
        RECT 87.295 190.685 87.625 191.665 ;
        RECT 87.795 190.515 88.025 191.655 ;
        RECT 88.235 191.275 88.575 192.085 ;
        RECT 88.745 191.520 89.495 191.710 ;
        RECT 88.235 190.865 88.750 191.275 ;
        RECT 88.985 190.515 89.155 191.275 ;
        RECT 89.325 190.855 89.495 191.520 ;
        RECT 89.665 191.535 89.855 192.895 ;
        RECT 90.025 192.725 90.300 192.895 ;
        RECT 90.025 192.555 90.305 192.725 ;
        RECT 90.025 191.735 90.300 192.555 ;
        RECT 90.490 192.530 91.020 192.895 ;
        RECT 91.445 192.665 91.775 193.065 ;
        RECT 90.845 192.495 91.020 192.530 ;
        RECT 90.505 191.535 90.675 192.335 ;
        RECT 89.665 191.365 90.675 191.535 ;
        RECT 90.845 192.325 91.775 192.495 ;
        RECT 91.945 192.325 92.200 192.895 ;
        RECT 92.465 192.515 92.635 192.895 ;
        RECT 92.815 192.685 93.145 193.065 ;
        RECT 92.465 192.345 93.130 192.515 ;
        RECT 93.325 192.390 93.585 192.895 ;
        RECT 90.845 191.195 91.015 192.325 ;
        RECT 91.605 192.155 91.775 192.325 ;
        RECT 89.890 191.025 91.015 191.195 ;
        RECT 91.185 191.825 91.380 192.155 ;
        RECT 91.605 191.825 91.860 192.155 ;
        RECT 91.185 190.855 91.355 191.825 ;
        RECT 92.030 191.655 92.200 192.325 ;
        RECT 92.395 191.795 92.725 192.165 ;
        RECT 92.960 192.090 93.130 192.345 ;
        RECT 89.325 190.685 91.355 190.855 ;
        RECT 91.525 190.515 91.695 191.655 ;
        RECT 91.865 190.685 92.200 191.655 ;
        RECT 92.960 191.760 93.245 192.090 ;
        RECT 92.960 191.615 93.130 191.760 ;
        RECT 92.465 191.445 93.130 191.615 ;
        RECT 93.415 191.590 93.585 192.390 ;
        RECT 94.030 192.255 94.275 192.860 ;
        RECT 94.495 192.530 95.005 193.065 ;
        RECT 92.465 190.685 92.635 191.445 ;
        RECT 92.815 190.515 93.145 191.275 ;
        RECT 93.315 190.685 93.585 191.590 ;
        RECT 93.755 192.085 94.985 192.255 ;
        RECT 93.755 191.275 94.095 192.085 ;
        RECT 94.265 191.520 95.015 191.710 ;
        RECT 93.755 190.865 94.270 191.275 ;
        RECT 94.505 190.515 94.675 191.275 ;
        RECT 94.845 190.855 95.015 191.520 ;
        RECT 95.185 191.535 95.375 192.895 ;
        RECT 95.545 192.045 95.820 192.895 ;
        RECT 96.010 192.530 96.540 192.895 ;
        RECT 96.965 192.665 97.295 193.065 ;
        RECT 96.365 192.495 96.540 192.530 ;
        RECT 95.545 191.875 95.825 192.045 ;
        RECT 95.545 191.735 95.820 191.875 ;
        RECT 96.025 191.535 96.195 192.335 ;
        RECT 95.185 191.365 96.195 191.535 ;
        RECT 96.365 192.325 97.295 192.495 ;
        RECT 97.465 192.325 97.720 192.895 ;
        RECT 98.905 192.515 99.075 192.895 ;
        RECT 99.255 192.685 99.585 193.065 ;
        RECT 98.905 192.345 99.570 192.515 ;
        RECT 99.765 192.390 100.025 192.895 ;
        RECT 96.365 191.195 96.535 192.325 ;
        RECT 97.125 192.155 97.295 192.325 ;
        RECT 95.410 191.025 96.535 191.195 ;
        RECT 96.705 191.825 96.900 192.155 ;
        RECT 97.125 191.825 97.380 192.155 ;
        RECT 96.705 190.855 96.875 191.825 ;
        RECT 97.550 191.655 97.720 192.325 ;
        RECT 98.835 191.795 99.165 192.165 ;
        RECT 99.400 192.090 99.570 192.345 ;
        RECT 94.845 190.685 96.875 190.855 ;
        RECT 97.045 190.515 97.215 191.655 ;
        RECT 97.385 190.685 97.720 191.655 ;
        RECT 99.400 191.760 99.685 192.090 ;
        RECT 99.400 191.615 99.570 191.760 ;
        RECT 98.905 191.445 99.570 191.615 ;
        RECT 99.855 191.590 100.025 192.390 ;
        RECT 100.195 192.340 100.485 193.065 ;
        RECT 100.930 192.255 101.175 192.860 ;
        RECT 101.395 192.530 101.905 193.065 ;
        RECT 100.655 192.085 101.885 192.255 ;
        RECT 98.905 190.685 99.075 191.445 ;
        RECT 99.255 190.515 99.585 191.275 ;
        RECT 99.755 190.685 100.025 191.590 ;
        RECT 100.195 190.515 100.485 191.680 ;
        RECT 100.655 191.275 100.995 192.085 ;
        RECT 101.165 191.520 101.915 191.710 ;
        RECT 100.655 190.865 101.170 191.275 ;
        RECT 101.405 190.515 101.575 191.275 ;
        RECT 101.745 190.855 101.915 191.520 ;
        RECT 102.085 191.535 102.275 192.895 ;
        RECT 102.445 192.725 102.720 192.895 ;
        RECT 102.445 192.555 102.725 192.725 ;
        RECT 102.445 191.735 102.720 192.555 ;
        RECT 102.910 192.530 103.440 192.895 ;
        RECT 103.865 192.665 104.195 193.065 ;
        RECT 103.265 192.495 103.440 192.530 ;
        RECT 102.925 191.535 103.095 192.335 ;
        RECT 102.085 191.365 103.095 191.535 ;
        RECT 103.265 192.325 104.195 192.495 ;
        RECT 104.365 192.325 104.620 192.895 ;
        RECT 103.265 191.195 103.435 192.325 ;
        RECT 104.025 192.155 104.195 192.325 ;
        RECT 102.310 191.025 103.435 191.195 ;
        RECT 103.605 191.825 103.800 192.155 ;
        RECT 104.025 191.825 104.280 192.155 ;
        RECT 103.605 190.855 103.775 191.825 ;
        RECT 104.450 191.655 104.620 192.325 ;
        RECT 101.745 190.685 103.775 190.855 ;
        RECT 103.945 190.515 104.115 191.655 ;
        RECT 104.285 190.685 104.620 191.655 ;
        RECT 104.795 192.325 105.180 192.895 ;
        RECT 105.350 192.605 105.675 193.065 ;
        RECT 106.195 192.435 106.475 192.895 ;
        RECT 104.795 191.655 105.075 192.325 ;
        RECT 105.350 192.265 106.475 192.435 ;
        RECT 105.350 192.155 105.800 192.265 ;
        RECT 105.245 191.825 105.800 192.155 ;
        RECT 106.665 192.095 107.065 192.895 ;
        RECT 107.465 192.605 107.735 193.065 ;
        RECT 107.905 192.435 108.190 192.895 ;
        RECT 104.795 190.685 105.180 191.655 ;
        RECT 105.350 191.365 105.800 191.825 ;
        RECT 105.970 191.535 107.065 192.095 ;
        RECT 105.350 191.145 106.475 191.365 ;
        RECT 105.350 190.515 105.675 190.975 ;
        RECT 106.195 190.685 106.475 191.145 ;
        RECT 106.665 190.685 107.065 191.535 ;
        RECT 107.235 192.265 108.190 192.435 ;
        RECT 108.475 192.325 108.860 192.895 ;
        RECT 109.030 192.605 109.355 193.065 ;
        RECT 109.875 192.435 110.155 192.895 ;
        RECT 107.235 191.365 107.445 192.265 ;
        RECT 107.615 191.535 108.305 192.095 ;
        RECT 108.475 191.655 108.755 192.325 ;
        RECT 109.030 192.265 110.155 192.435 ;
        RECT 109.030 192.155 109.480 192.265 ;
        RECT 108.925 191.825 109.480 192.155 ;
        RECT 110.345 192.095 110.745 192.895 ;
        RECT 111.145 192.605 111.415 193.065 ;
        RECT 111.585 192.435 111.870 192.895 ;
        RECT 107.235 191.145 108.190 191.365 ;
        RECT 107.465 190.515 107.735 190.975 ;
        RECT 107.905 190.685 108.190 191.145 ;
        RECT 108.475 190.685 108.860 191.655 ;
        RECT 109.030 191.365 109.480 191.825 ;
        RECT 109.650 191.535 110.745 192.095 ;
        RECT 109.030 191.145 110.155 191.365 ;
        RECT 109.030 190.515 109.355 190.975 ;
        RECT 109.875 190.685 110.155 191.145 ;
        RECT 110.345 190.685 110.745 191.535 ;
        RECT 110.915 192.265 111.870 192.435 ;
        RECT 112.155 192.315 113.365 193.065 ;
        RECT 110.915 191.365 111.125 192.265 ;
        RECT 111.295 191.535 111.985 192.095 ;
        RECT 112.155 191.605 112.675 192.145 ;
        RECT 112.845 191.775 113.365 192.315 ;
        RECT 110.915 191.145 111.870 191.365 ;
        RECT 111.145 190.515 111.415 190.975 ;
        RECT 111.585 190.685 111.870 191.145 ;
        RECT 112.155 190.515 113.365 191.605 ;
        RECT 22.830 190.345 113.450 190.515 ;
        RECT 22.915 189.255 24.125 190.345 ;
        RECT 24.410 189.715 24.695 190.175 ;
        RECT 24.865 189.885 25.135 190.345 ;
        RECT 24.410 189.495 25.365 189.715 ;
        RECT 22.915 188.545 23.435 189.085 ;
        RECT 23.605 188.715 24.125 189.255 ;
        RECT 24.295 188.765 24.985 189.325 ;
        RECT 25.155 188.595 25.365 189.495 ;
        RECT 22.915 187.795 24.125 188.545 ;
        RECT 24.410 188.425 25.365 188.595 ;
        RECT 25.535 189.325 25.935 190.175 ;
        RECT 26.125 189.715 26.405 190.175 ;
        RECT 26.925 189.885 27.250 190.345 ;
        RECT 26.125 189.495 27.250 189.715 ;
        RECT 25.535 188.765 26.630 189.325 ;
        RECT 26.800 189.035 27.250 189.495 ;
        RECT 27.420 189.205 27.805 190.175 ;
        RECT 24.410 187.965 24.695 188.425 ;
        RECT 24.865 187.795 25.135 188.255 ;
        RECT 25.535 187.965 25.935 188.765 ;
        RECT 26.800 188.705 27.355 189.035 ;
        RECT 26.800 188.595 27.250 188.705 ;
        RECT 26.125 188.425 27.250 188.595 ;
        RECT 27.525 188.535 27.805 189.205 ;
        RECT 26.125 187.965 26.405 188.425 ;
        RECT 26.925 187.795 27.250 188.255 ;
        RECT 27.420 187.965 27.805 188.535 ;
        RECT 28.435 189.205 28.820 190.175 ;
        RECT 28.990 189.885 29.315 190.345 ;
        RECT 29.835 189.715 30.115 190.175 ;
        RECT 28.990 189.495 30.115 189.715 ;
        RECT 28.435 188.535 28.715 189.205 ;
        RECT 28.990 189.035 29.440 189.495 ;
        RECT 30.305 189.325 30.705 190.175 ;
        RECT 31.105 189.885 31.375 190.345 ;
        RECT 31.545 189.715 31.830 190.175 ;
        RECT 28.885 188.705 29.440 189.035 ;
        RECT 29.610 188.765 30.705 189.325 ;
        RECT 28.990 188.595 29.440 188.705 ;
        RECT 28.435 187.965 28.820 188.535 ;
        RECT 28.990 188.425 30.115 188.595 ;
        RECT 28.990 187.795 29.315 188.255 ;
        RECT 29.835 187.965 30.115 188.425 ;
        RECT 30.305 187.965 30.705 188.765 ;
        RECT 30.875 189.495 31.830 189.715 ;
        RECT 30.875 188.595 31.085 189.495 ;
        RECT 31.255 188.765 31.945 189.325 ;
        RECT 32.115 189.205 32.455 190.175 ;
        RECT 32.625 189.205 32.795 190.345 ;
        RECT 33.065 189.545 33.315 190.345 ;
        RECT 33.960 189.375 34.290 190.175 ;
        RECT 34.590 189.545 34.920 190.345 ;
        RECT 35.090 189.375 35.420 190.175 ;
        RECT 32.985 189.205 35.420 189.375 ;
        RECT 32.115 189.155 32.345 189.205 ;
        RECT 32.115 188.595 32.290 189.155 ;
        RECT 32.985 188.955 33.155 189.205 ;
        RECT 32.460 188.785 33.155 188.955 ;
        RECT 33.330 188.785 33.750 188.985 ;
        RECT 33.920 188.785 34.250 188.985 ;
        RECT 34.420 188.785 34.750 188.985 ;
        RECT 30.875 188.425 31.830 188.595 ;
        RECT 31.105 187.795 31.375 188.255 ;
        RECT 31.545 187.965 31.830 188.425 ;
        RECT 32.115 187.965 32.455 188.595 ;
        RECT 32.625 187.795 32.875 188.595 ;
        RECT 33.065 188.445 34.290 188.615 ;
        RECT 33.065 187.965 33.395 188.445 ;
        RECT 33.565 187.795 33.790 188.255 ;
        RECT 33.960 187.965 34.290 188.445 ;
        RECT 34.920 188.575 35.090 189.205 ;
        RECT 35.795 189.180 36.085 190.345 ;
        RECT 36.260 189.205 36.595 190.175 ;
        RECT 36.765 189.205 36.935 190.345 ;
        RECT 37.105 190.005 39.135 190.175 ;
        RECT 35.275 188.785 35.625 189.035 ;
        RECT 34.920 187.965 35.420 188.575 ;
        RECT 36.260 188.535 36.430 189.205 ;
        RECT 37.105 189.035 37.275 190.005 ;
        RECT 36.600 188.705 36.855 189.035 ;
        RECT 37.080 188.705 37.275 189.035 ;
        RECT 37.445 189.665 38.570 189.835 ;
        RECT 36.685 188.535 36.855 188.705 ;
        RECT 37.445 188.535 37.615 189.665 ;
        RECT 35.795 187.795 36.085 188.520 ;
        RECT 36.260 187.965 36.515 188.535 ;
        RECT 36.685 188.365 37.615 188.535 ;
        RECT 37.785 189.325 38.795 189.495 ;
        RECT 37.785 188.525 37.955 189.325 ;
        RECT 37.440 188.330 37.615 188.365 ;
        RECT 36.685 187.795 37.015 188.195 ;
        RECT 37.440 187.965 37.970 188.330 ;
        RECT 38.160 188.305 38.435 189.125 ;
        RECT 38.155 188.135 38.435 188.305 ;
        RECT 38.160 187.965 38.435 188.135 ;
        RECT 38.605 187.965 38.795 189.325 ;
        RECT 38.965 189.340 39.135 190.005 ;
        RECT 39.305 189.585 39.475 190.345 ;
        RECT 39.710 189.585 40.225 189.995 ;
        RECT 38.965 189.150 39.715 189.340 ;
        RECT 39.885 188.775 40.225 189.585 ;
        RECT 40.485 189.415 40.655 190.175 ;
        RECT 40.835 189.585 41.165 190.345 ;
        RECT 40.485 189.245 41.150 189.415 ;
        RECT 41.335 189.270 41.605 190.175 ;
        RECT 40.980 189.100 41.150 189.245 ;
        RECT 38.995 188.605 40.225 188.775 ;
        RECT 40.415 188.695 40.745 189.065 ;
        RECT 40.980 188.770 41.265 189.100 ;
        RECT 38.975 187.795 39.485 188.330 ;
        RECT 39.705 188.000 39.950 188.605 ;
        RECT 40.980 188.515 41.150 188.770 ;
        RECT 40.485 188.345 41.150 188.515 ;
        RECT 41.435 188.470 41.605 189.270 ;
        RECT 41.815 189.205 42.045 190.345 ;
        RECT 42.215 189.195 42.545 190.175 ;
        RECT 42.715 189.205 42.925 190.345 ;
        RECT 43.160 189.675 43.415 190.175 ;
        RECT 43.585 189.845 43.915 190.345 ;
        RECT 43.160 189.505 43.910 189.675 ;
        RECT 41.795 188.785 42.125 189.035 ;
        RECT 40.485 187.965 40.655 188.345 ;
        RECT 40.835 187.795 41.165 188.175 ;
        RECT 41.345 187.965 41.605 188.470 ;
        RECT 41.815 187.795 42.045 188.615 ;
        RECT 42.295 188.595 42.545 189.195 ;
        RECT 43.160 188.685 43.510 189.335 ;
        RECT 42.215 187.965 42.545 188.595 ;
        RECT 42.715 187.795 42.925 188.615 ;
        RECT 43.680 188.515 43.910 189.505 ;
        RECT 43.160 188.345 43.910 188.515 ;
        RECT 43.160 188.055 43.415 188.345 ;
        RECT 43.585 187.795 43.915 188.175 ;
        RECT 44.085 188.055 44.255 190.175 ;
        RECT 44.425 189.375 44.750 190.160 ;
        RECT 44.920 189.885 45.170 190.345 ;
        RECT 45.340 189.845 45.590 190.175 ;
        RECT 45.805 189.845 46.485 190.175 ;
        RECT 45.340 189.715 45.510 189.845 ;
        RECT 45.115 189.545 45.510 189.715 ;
        RECT 44.485 188.325 44.945 189.375 ;
        RECT 45.115 188.185 45.285 189.545 ;
        RECT 45.680 189.285 46.145 189.675 ;
        RECT 45.455 188.475 45.805 189.095 ;
        RECT 45.975 188.695 46.145 189.285 ;
        RECT 46.315 189.065 46.485 189.845 ;
        RECT 46.655 189.745 46.825 190.085 ;
        RECT 47.060 189.915 47.390 190.345 ;
        RECT 47.560 189.745 47.730 190.085 ;
        RECT 48.025 189.885 48.395 190.345 ;
        RECT 46.655 189.575 47.730 189.745 ;
        RECT 48.565 189.715 48.735 190.175 ;
        RECT 48.970 189.835 49.840 190.175 ;
        RECT 50.010 189.885 50.260 190.345 ;
        RECT 48.175 189.545 48.735 189.715 ;
        RECT 48.175 189.405 48.345 189.545 ;
        RECT 46.845 189.235 48.345 189.405 ;
        RECT 49.040 189.375 49.500 189.665 ;
        RECT 46.315 188.895 48.005 189.065 ;
        RECT 45.975 188.475 46.330 188.695 ;
        RECT 46.500 188.185 46.670 188.895 ;
        RECT 46.875 188.475 47.665 188.725 ;
        RECT 47.835 188.715 48.005 188.895 ;
        RECT 48.175 188.545 48.345 189.235 ;
        RECT 44.615 187.795 44.945 188.155 ;
        RECT 45.115 188.015 45.610 188.185 ;
        RECT 45.815 188.015 46.670 188.185 ;
        RECT 47.545 187.795 47.875 188.255 ;
        RECT 48.085 188.155 48.345 188.545 ;
        RECT 48.535 189.365 49.500 189.375 ;
        RECT 49.670 189.455 49.840 189.835 ;
        RECT 50.430 189.795 50.600 190.085 ;
        RECT 50.780 189.965 51.110 190.345 ;
        RECT 50.430 189.625 51.230 189.795 ;
        RECT 48.535 189.205 49.210 189.365 ;
        RECT 49.670 189.285 50.890 189.455 ;
        RECT 48.535 188.415 48.745 189.205 ;
        RECT 49.670 189.195 49.840 189.285 ;
        RECT 48.915 188.415 49.265 189.035 ;
        RECT 49.435 189.025 49.840 189.195 ;
        RECT 49.435 188.245 49.605 189.025 ;
        RECT 49.775 188.575 49.995 188.855 ;
        RECT 50.175 188.745 50.715 189.115 ;
        RECT 51.060 189.035 51.230 189.625 ;
        RECT 51.450 189.205 51.755 190.345 ;
        RECT 51.925 189.155 52.180 190.035 ;
        RECT 51.060 189.005 51.800 189.035 ;
        RECT 49.775 188.405 50.305 188.575 ;
        RECT 48.085 187.985 48.435 188.155 ;
        RECT 48.655 187.965 49.605 188.245 ;
        RECT 49.775 187.795 49.965 188.235 ;
        RECT 50.135 188.175 50.305 188.405 ;
        RECT 50.475 188.345 50.715 188.745 ;
        RECT 50.885 188.705 51.800 189.005 ;
        RECT 50.885 188.530 51.210 188.705 ;
        RECT 50.885 188.175 51.205 188.530 ;
        RECT 51.970 188.505 52.180 189.155 ;
        RECT 50.135 188.005 51.205 188.175 ;
        RECT 51.450 187.795 51.755 188.255 ;
        RECT 51.925 187.975 52.180 188.505 ;
        RECT 52.360 189.155 52.615 190.035 ;
        RECT 52.785 189.205 53.090 190.345 ;
        RECT 53.430 189.965 53.760 190.345 ;
        RECT 53.940 189.795 54.110 190.085 ;
        RECT 54.280 189.885 54.530 190.345 ;
        RECT 53.310 189.625 54.110 189.795 ;
        RECT 54.700 189.835 55.570 190.175 ;
        RECT 52.360 188.505 52.570 189.155 ;
        RECT 53.310 189.035 53.480 189.625 ;
        RECT 54.700 189.455 54.870 189.835 ;
        RECT 55.805 189.715 55.975 190.175 ;
        RECT 56.145 189.885 56.515 190.345 ;
        RECT 56.810 189.745 56.980 190.085 ;
        RECT 57.150 189.915 57.480 190.345 ;
        RECT 57.715 189.745 57.885 190.085 ;
        RECT 53.650 189.285 54.870 189.455 ;
        RECT 55.040 189.375 55.500 189.665 ;
        RECT 55.805 189.545 56.365 189.715 ;
        RECT 56.810 189.575 57.885 189.745 ;
        RECT 58.055 189.845 58.735 190.175 ;
        RECT 58.950 189.845 59.200 190.175 ;
        RECT 59.370 189.885 59.620 190.345 ;
        RECT 56.195 189.405 56.365 189.545 ;
        RECT 55.040 189.365 56.005 189.375 ;
        RECT 54.700 189.195 54.870 189.285 ;
        RECT 55.330 189.205 56.005 189.365 ;
        RECT 52.740 189.005 53.480 189.035 ;
        RECT 52.740 188.705 53.655 189.005 ;
        RECT 53.330 188.530 53.655 188.705 ;
        RECT 52.360 187.975 52.615 188.505 ;
        RECT 52.785 187.795 53.090 188.255 ;
        RECT 53.335 188.175 53.655 188.530 ;
        RECT 53.825 188.745 54.365 189.115 ;
        RECT 54.700 189.025 55.105 189.195 ;
        RECT 53.825 188.345 54.065 188.745 ;
        RECT 54.545 188.575 54.765 188.855 ;
        RECT 54.235 188.405 54.765 188.575 ;
        RECT 54.235 188.175 54.405 188.405 ;
        RECT 54.935 188.245 55.105 189.025 ;
        RECT 55.275 188.415 55.625 189.035 ;
        RECT 55.795 188.415 56.005 189.205 ;
        RECT 56.195 189.235 57.695 189.405 ;
        RECT 56.195 188.545 56.365 189.235 ;
        RECT 58.055 189.065 58.225 189.845 ;
        RECT 59.030 189.715 59.200 189.845 ;
        RECT 56.535 188.895 58.225 189.065 ;
        RECT 58.395 189.285 58.860 189.675 ;
        RECT 59.030 189.545 59.425 189.715 ;
        RECT 56.535 188.715 56.705 188.895 ;
        RECT 53.335 188.005 54.405 188.175 ;
        RECT 54.575 187.795 54.765 188.235 ;
        RECT 54.935 187.965 55.885 188.245 ;
        RECT 56.195 188.155 56.455 188.545 ;
        RECT 56.875 188.475 57.665 188.725 ;
        RECT 56.105 187.985 56.455 188.155 ;
        RECT 56.665 187.795 56.995 188.255 ;
        RECT 57.870 188.185 58.040 188.895 ;
        RECT 58.395 188.695 58.565 189.285 ;
        RECT 58.210 188.475 58.565 188.695 ;
        RECT 58.735 188.475 59.085 189.095 ;
        RECT 59.255 188.185 59.425 189.545 ;
        RECT 59.790 189.375 60.115 190.160 ;
        RECT 59.595 188.325 60.055 189.375 ;
        RECT 57.870 188.015 58.725 188.185 ;
        RECT 58.930 188.015 59.425 188.185 ;
        RECT 59.595 187.795 59.925 188.155 ;
        RECT 60.285 188.055 60.455 190.175 ;
        RECT 60.625 189.845 60.955 190.345 ;
        RECT 61.125 189.675 61.380 190.175 ;
        RECT 60.630 189.505 61.380 189.675 ;
        RECT 60.630 188.515 60.860 189.505 ;
        RECT 61.030 188.685 61.380 189.335 ;
        RECT 61.555 189.180 61.845 190.345 ;
        RECT 62.020 189.910 67.365 190.345 ;
        RECT 63.610 188.660 63.960 189.910 ;
        RECT 60.630 188.345 61.380 188.515 ;
        RECT 60.625 187.795 60.955 188.175 ;
        RECT 61.125 188.055 61.380 188.345 ;
        RECT 61.555 187.795 61.845 188.520 ;
        RECT 65.440 188.340 65.780 189.170 ;
        RECT 67.535 188.535 67.795 190.160 ;
        RECT 69.545 189.895 69.875 190.345 ;
        RECT 71.465 189.895 71.795 190.345 ;
        RECT 67.975 189.505 70.585 189.715 ;
        RECT 67.975 188.705 68.195 189.505 ;
        RECT 68.435 188.705 68.735 189.325 ;
        RECT 68.905 188.705 69.235 189.325 ;
        RECT 69.405 188.705 69.725 189.325 ;
        RECT 69.895 188.705 70.245 189.325 ;
        RECT 70.415 188.535 70.585 189.505 ;
        RECT 67.535 188.365 69.375 188.535 ;
        RECT 62.020 187.795 67.365 188.340 ;
        RECT 67.805 187.795 68.135 188.190 ;
        RECT 68.305 188.010 68.505 188.365 ;
        RECT 68.675 187.795 69.005 188.195 ;
        RECT 69.175 188.020 69.375 188.365 ;
        RECT 69.545 187.795 69.875 188.535 ;
        RECT 70.110 188.365 70.585 188.535 ;
        RECT 70.755 189.505 73.365 189.715 ;
        RECT 70.755 188.535 70.925 189.505 ;
        RECT 71.095 188.705 71.445 189.325 ;
        RECT 71.615 188.705 71.935 189.325 ;
        RECT 72.105 188.705 72.435 189.325 ;
        RECT 72.605 188.705 72.905 189.325 ;
        RECT 73.145 188.705 73.365 189.505 ;
        RECT 73.545 188.535 73.805 190.160 ;
        RECT 73.985 189.365 74.315 190.175 ;
        RECT 74.485 189.545 74.725 190.345 ;
        RECT 73.985 189.195 74.700 189.365 ;
        RECT 73.980 188.785 74.360 189.025 ;
        RECT 74.530 188.955 74.700 189.195 ;
        RECT 74.905 189.325 75.075 190.175 ;
        RECT 75.245 189.545 75.575 190.345 ;
        RECT 75.745 189.325 75.915 190.175 ;
        RECT 74.905 189.155 75.915 189.325 ;
        RECT 76.085 189.195 76.415 190.345 ;
        RECT 78.030 189.365 78.285 190.035 ;
        RECT 78.465 189.545 78.750 190.345 ;
        RECT 78.930 189.625 79.260 190.135 ;
        RECT 74.530 188.785 75.030 188.955 ;
        RECT 74.530 188.615 74.700 188.785 ;
        RECT 75.420 188.645 75.915 189.155 ;
        RECT 75.415 188.615 75.915 188.645 ;
        RECT 70.755 188.365 71.230 188.535 ;
        RECT 70.110 188.115 70.280 188.365 ;
        RECT 71.060 188.115 71.230 188.365 ;
        RECT 71.465 187.795 71.795 188.535 ;
        RECT 71.965 188.365 73.805 188.535 ;
        RECT 74.065 188.445 74.700 188.615 ;
        RECT 74.905 188.445 75.915 188.615 ;
        RECT 71.965 188.020 72.165 188.365 ;
        RECT 72.335 187.795 72.665 188.195 ;
        RECT 72.835 188.010 73.035 188.365 ;
        RECT 73.205 187.795 73.535 188.190 ;
        RECT 74.065 187.965 74.235 188.445 ;
        RECT 74.415 187.795 74.655 188.275 ;
        RECT 74.905 187.965 75.075 188.445 ;
        RECT 75.245 187.795 75.575 188.275 ;
        RECT 75.745 187.965 75.915 188.445 ;
        RECT 76.085 187.795 76.415 188.595 ;
        RECT 78.030 188.505 78.210 189.365 ;
        RECT 78.930 189.035 79.180 189.625 ;
        RECT 79.530 189.475 79.700 190.085 ;
        RECT 79.870 189.655 80.200 190.345 ;
        RECT 80.430 189.795 80.670 190.085 ;
        RECT 80.870 189.965 81.290 190.345 ;
        RECT 81.470 189.875 82.100 190.125 ;
        RECT 82.570 189.965 82.900 190.345 ;
        RECT 81.470 189.795 81.640 189.875 ;
        RECT 83.070 189.795 83.240 190.085 ;
        RECT 83.420 189.965 83.800 190.345 ;
        RECT 84.040 189.960 84.870 190.130 ;
        RECT 80.430 189.625 81.640 189.795 ;
        RECT 78.380 188.705 79.180 189.035 ;
        RECT 78.030 188.305 78.285 188.505 ;
        RECT 77.945 188.135 78.285 188.305 ;
        RECT 78.030 187.975 78.285 188.135 ;
        RECT 78.465 187.795 78.750 188.255 ;
        RECT 78.930 188.055 79.180 188.705 ;
        RECT 79.380 189.455 79.700 189.475 ;
        RECT 79.380 189.285 81.300 189.455 ;
        RECT 79.380 188.390 79.570 189.285 ;
        RECT 81.470 189.115 81.640 189.625 ;
        RECT 81.810 189.365 82.330 189.675 ;
        RECT 79.740 188.945 81.640 189.115 ;
        RECT 79.740 188.885 80.070 188.945 ;
        RECT 80.220 188.715 80.550 188.775 ;
        RECT 79.890 188.445 80.550 188.715 ;
        RECT 79.380 188.060 79.700 188.390 ;
        RECT 79.880 187.795 80.540 188.275 ;
        RECT 80.740 188.185 80.910 188.945 ;
        RECT 81.810 188.775 81.990 189.185 ;
        RECT 81.080 188.605 81.410 188.725 ;
        RECT 82.160 188.605 82.330 189.365 ;
        RECT 81.080 188.435 82.330 188.605 ;
        RECT 82.500 189.545 83.870 189.795 ;
        RECT 82.500 188.775 82.690 189.545 ;
        RECT 83.620 189.285 83.870 189.545 ;
        RECT 82.860 189.115 83.110 189.275 ;
        RECT 84.040 189.115 84.210 189.960 ;
        RECT 85.105 189.675 85.275 190.175 ;
        RECT 85.445 189.845 85.775 190.345 ;
        RECT 84.380 189.285 84.880 189.665 ;
        RECT 85.105 189.505 85.800 189.675 ;
        RECT 82.860 188.945 84.210 189.115 ;
        RECT 83.790 188.905 84.210 188.945 ;
        RECT 82.500 188.435 82.920 188.775 ;
        RECT 83.210 188.445 83.620 188.775 ;
        RECT 80.740 188.015 81.590 188.185 ;
        RECT 82.150 187.795 82.470 188.255 ;
        RECT 82.670 188.005 82.920 188.435 ;
        RECT 83.210 187.795 83.620 188.235 ;
        RECT 83.790 188.175 83.960 188.905 ;
        RECT 84.130 188.355 84.480 188.725 ;
        RECT 84.660 188.415 84.880 189.285 ;
        RECT 85.050 188.715 85.460 189.335 ;
        RECT 85.630 188.535 85.800 189.505 ;
        RECT 85.105 188.345 85.800 188.535 ;
        RECT 83.790 187.975 84.805 188.175 ;
        RECT 85.105 188.015 85.275 188.345 ;
        RECT 85.445 187.795 85.775 188.175 ;
        RECT 85.990 188.055 86.215 190.175 ;
        RECT 86.385 189.845 86.715 190.345 ;
        RECT 86.885 189.675 87.055 190.175 ;
        RECT 86.390 189.505 87.055 189.675 ;
        RECT 86.390 188.515 86.620 189.505 ;
        RECT 86.790 188.685 87.140 189.335 ;
        RECT 87.315 189.180 87.605 190.345 ;
        RECT 87.890 189.715 88.175 190.175 ;
        RECT 88.345 189.885 88.615 190.345 ;
        RECT 87.890 189.495 88.845 189.715 ;
        RECT 87.775 188.765 88.465 189.325 ;
        RECT 88.635 188.595 88.845 189.495 ;
        RECT 86.390 188.345 87.055 188.515 ;
        RECT 86.385 187.795 86.715 188.175 ;
        RECT 86.885 188.055 87.055 188.345 ;
        RECT 87.315 187.795 87.605 188.520 ;
        RECT 87.890 188.425 88.845 188.595 ;
        RECT 89.015 189.325 89.415 190.175 ;
        RECT 89.605 189.715 89.885 190.175 ;
        RECT 90.405 189.885 90.730 190.345 ;
        RECT 89.605 189.495 90.730 189.715 ;
        RECT 89.015 188.765 90.110 189.325 ;
        RECT 90.280 189.035 90.730 189.495 ;
        RECT 90.900 189.205 91.285 190.175 ;
        RECT 87.890 187.965 88.175 188.425 ;
        RECT 88.345 187.795 88.615 188.255 ;
        RECT 89.015 187.965 89.415 188.765 ;
        RECT 90.280 188.705 90.835 189.035 ;
        RECT 90.280 188.595 90.730 188.705 ;
        RECT 89.605 188.425 90.730 188.595 ;
        RECT 91.005 188.535 91.285 189.205 ;
        RECT 91.915 189.585 92.430 189.995 ;
        RECT 92.665 189.585 92.835 190.345 ;
        RECT 93.005 190.005 95.035 190.175 ;
        RECT 91.915 188.775 92.255 189.585 ;
        RECT 93.005 189.340 93.175 190.005 ;
        RECT 93.570 189.665 94.695 189.835 ;
        RECT 92.425 189.150 93.175 189.340 ;
        RECT 93.345 189.325 94.355 189.495 ;
        RECT 91.915 188.605 93.145 188.775 ;
        RECT 89.605 187.965 89.885 188.425 ;
        RECT 90.405 187.795 90.730 188.255 ;
        RECT 90.900 187.965 91.285 188.535 ;
        RECT 92.190 188.000 92.435 188.605 ;
        RECT 92.655 187.795 93.165 188.330 ;
        RECT 93.345 187.965 93.535 189.325 ;
        RECT 93.705 188.985 93.980 189.125 ;
        RECT 93.705 188.815 93.985 188.985 ;
        RECT 93.705 187.965 93.980 188.815 ;
        RECT 94.185 188.525 94.355 189.325 ;
        RECT 94.525 188.535 94.695 189.665 ;
        RECT 94.865 189.035 95.035 190.005 ;
        RECT 95.205 189.205 95.375 190.345 ;
        RECT 95.545 189.205 95.880 190.175 ;
        RECT 94.865 188.705 95.060 189.035 ;
        RECT 95.285 188.705 95.540 189.035 ;
        RECT 95.285 188.535 95.455 188.705 ;
        RECT 95.710 188.535 95.880 189.205 ;
        RECT 96.975 189.585 97.490 189.995 ;
        RECT 97.725 189.585 97.895 190.345 ;
        RECT 98.065 190.005 100.095 190.175 ;
        RECT 96.975 188.775 97.315 189.585 ;
        RECT 98.065 189.340 98.235 190.005 ;
        RECT 98.630 189.665 99.755 189.835 ;
        RECT 97.485 189.150 98.235 189.340 ;
        RECT 98.405 189.325 99.415 189.495 ;
        RECT 96.975 188.605 98.205 188.775 ;
        RECT 94.525 188.365 95.455 188.535 ;
        RECT 94.525 188.330 94.700 188.365 ;
        RECT 94.170 187.965 94.700 188.330 ;
        RECT 95.125 187.795 95.455 188.195 ;
        RECT 95.625 187.965 95.880 188.535 ;
        RECT 97.250 188.000 97.495 188.605 ;
        RECT 97.715 187.795 98.225 188.330 ;
        RECT 98.405 187.965 98.595 189.325 ;
        RECT 98.765 188.985 99.040 189.125 ;
        RECT 98.765 188.815 99.045 188.985 ;
        RECT 98.765 187.965 99.040 188.815 ;
        RECT 99.245 188.525 99.415 189.325 ;
        RECT 99.585 188.535 99.755 189.665 ;
        RECT 99.925 189.035 100.095 190.005 ;
        RECT 100.265 189.205 100.435 190.345 ;
        RECT 100.605 189.205 100.940 190.175 ;
        RECT 99.925 188.705 100.120 189.035 ;
        RECT 100.345 188.705 100.600 189.035 ;
        RECT 100.345 188.535 100.515 188.705 ;
        RECT 100.770 188.535 100.940 189.205 ;
        RECT 99.585 188.365 100.515 188.535 ;
        RECT 99.585 188.330 99.760 188.365 ;
        RECT 99.230 187.965 99.760 188.330 ;
        RECT 100.185 187.795 100.515 188.195 ;
        RECT 100.685 187.965 100.940 188.535 ;
        RECT 101.120 189.155 101.375 190.035 ;
        RECT 101.545 189.205 101.850 190.345 ;
        RECT 102.190 189.965 102.520 190.345 ;
        RECT 102.700 189.795 102.870 190.085 ;
        RECT 103.040 189.885 103.290 190.345 ;
        RECT 102.070 189.625 102.870 189.795 ;
        RECT 103.460 189.835 104.330 190.175 ;
        RECT 101.120 188.505 101.330 189.155 ;
        RECT 102.070 189.035 102.240 189.625 ;
        RECT 103.460 189.455 103.630 189.835 ;
        RECT 104.565 189.715 104.735 190.175 ;
        RECT 104.905 189.885 105.275 190.345 ;
        RECT 105.570 189.745 105.740 190.085 ;
        RECT 105.910 189.915 106.240 190.345 ;
        RECT 106.475 189.745 106.645 190.085 ;
        RECT 102.410 189.285 103.630 189.455 ;
        RECT 103.800 189.375 104.260 189.665 ;
        RECT 104.565 189.545 105.125 189.715 ;
        RECT 105.570 189.575 106.645 189.745 ;
        RECT 106.815 189.845 107.495 190.175 ;
        RECT 107.710 189.845 107.960 190.175 ;
        RECT 108.130 189.885 108.380 190.345 ;
        RECT 104.955 189.405 105.125 189.545 ;
        RECT 103.800 189.365 104.765 189.375 ;
        RECT 103.460 189.195 103.630 189.285 ;
        RECT 104.090 189.205 104.765 189.365 ;
        RECT 101.500 189.005 102.240 189.035 ;
        RECT 101.500 188.705 102.415 189.005 ;
        RECT 102.090 188.530 102.415 188.705 ;
        RECT 101.120 187.975 101.375 188.505 ;
        RECT 101.545 187.795 101.850 188.255 ;
        RECT 102.095 188.175 102.415 188.530 ;
        RECT 102.585 188.745 103.125 189.115 ;
        RECT 103.460 189.025 103.865 189.195 ;
        RECT 102.585 188.345 102.825 188.745 ;
        RECT 103.305 188.575 103.525 188.855 ;
        RECT 102.995 188.405 103.525 188.575 ;
        RECT 102.995 188.175 103.165 188.405 ;
        RECT 103.695 188.245 103.865 189.025 ;
        RECT 104.035 188.415 104.385 189.035 ;
        RECT 104.555 188.415 104.765 189.205 ;
        RECT 104.955 189.235 106.455 189.405 ;
        RECT 104.955 188.545 105.125 189.235 ;
        RECT 106.815 189.065 106.985 189.845 ;
        RECT 107.790 189.715 107.960 189.845 ;
        RECT 105.295 188.895 106.985 189.065 ;
        RECT 107.155 189.285 107.620 189.675 ;
        RECT 107.790 189.545 108.185 189.715 ;
        RECT 105.295 188.715 105.465 188.895 ;
        RECT 102.095 188.005 103.165 188.175 ;
        RECT 103.335 187.795 103.525 188.235 ;
        RECT 103.695 187.965 104.645 188.245 ;
        RECT 104.955 188.155 105.215 188.545 ;
        RECT 105.635 188.475 106.425 188.725 ;
        RECT 104.865 187.985 105.215 188.155 ;
        RECT 105.425 187.795 105.755 188.255 ;
        RECT 106.630 188.185 106.800 188.895 ;
        RECT 107.155 188.695 107.325 189.285 ;
        RECT 106.970 188.475 107.325 188.695 ;
        RECT 107.495 188.475 107.845 189.095 ;
        RECT 108.015 188.185 108.185 189.545 ;
        RECT 108.550 189.375 108.875 190.160 ;
        RECT 108.355 188.325 108.815 189.375 ;
        RECT 106.630 188.015 107.485 188.185 ;
        RECT 107.690 188.015 108.185 188.185 ;
        RECT 108.355 187.795 108.685 188.155 ;
        RECT 109.045 188.055 109.215 190.175 ;
        RECT 109.385 189.845 109.715 190.345 ;
        RECT 109.885 189.675 110.140 190.175 ;
        RECT 109.390 189.505 110.140 189.675 ;
        RECT 109.390 188.515 109.620 189.505 ;
        RECT 109.790 188.685 110.140 189.335 ;
        RECT 110.315 189.270 110.585 190.175 ;
        RECT 110.755 189.585 111.085 190.345 ;
        RECT 111.265 189.415 111.435 190.175 ;
        RECT 109.390 188.345 110.140 188.515 ;
        RECT 109.385 187.795 109.715 188.175 ;
        RECT 109.885 188.055 110.140 188.345 ;
        RECT 110.315 188.470 110.485 189.270 ;
        RECT 110.770 189.245 111.435 189.415 ;
        RECT 112.155 189.255 113.365 190.345 ;
        RECT 110.770 189.100 110.940 189.245 ;
        RECT 110.655 188.770 110.940 189.100 ;
        RECT 110.770 188.515 110.940 188.770 ;
        RECT 111.175 188.695 111.505 189.065 ;
        RECT 112.155 188.715 112.675 189.255 ;
        RECT 112.845 188.545 113.365 189.085 ;
        RECT 110.315 187.965 110.575 188.470 ;
        RECT 110.770 188.345 111.435 188.515 ;
        RECT 110.755 187.795 111.085 188.175 ;
        RECT 111.265 187.965 111.435 188.345 ;
        RECT 112.155 187.795 113.365 188.545 ;
        RECT 22.830 187.625 113.450 187.795 ;
        RECT 22.915 186.875 24.125 187.625 ;
        RECT 22.915 186.335 23.435 186.875 ;
        RECT 24.755 186.855 26.425 187.625 ;
        RECT 23.605 186.165 24.125 186.705 ;
        RECT 22.915 185.075 24.125 186.165 ;
        RECT 24.755 186.165 25.505 186.685 ;
        RECT 25.675 186.335 26.425 186.855 ;
        RECT 26.600 186.915 26.855 187.445 ;
        RECT 27.025 187.165 27.330 187.625 ;
        RECT 27.575 187.245 28.645 187.415 ;
        RECT 26.600 186.265 26.810 186.915 ;
        RECT 27.575 186.890 27.895 187.245 ;
        RECT 27.570 186.715 27.895 186.890 ;
        RECT 26.980 186.415 27.895 186.715 ;
        RECT 28.065 186.675 28.305 187.075 ;
        RECT 28.475 187.015 28.645 187.245 ;
        RECT 28.815 187.185 29.005 187.625 ;
        RECT 29.175 187.175 30.125 187.455 ;
        RECT 30.345 187.265 30.695 187.435 ;
        RECT 28.475 186.845 29.005 187.015 ;
        RECT 26.980 186.385 27.720 186.415 ;
        RECT 24.755 185.075 26.425 186.165 ;
        RECT 26.600 185.385 26.855 186.265 ;
        RECT 27.025 185.075 27.330 186.215 ;
        RECT 27.550 185.795 27.720 186.385 ;
        RECT 28.065 186.305 28.605 186.675 ;
        RECT 28.785 186.565 29.005 186.845 ;
        RECT 29.175 186.395 29.345 187.175 ;
        RECT 28.940 186.225 29.345 186.395 ;
        RECT 29.515 186.385 29.865 187.005 ;
        RECT 28.940 186.135 29.110 186.225 ;
        RECT 30.035 186.215 30.245 187.005 ;
        RECT 27.890 185.965 29.110 186.135 ;
        RECT 29.570 186.055 30.245 186.215 ;
        RECT 27.550 185.625 28.350 185.795 ;
        RECT 27.670 185.075 28.000 185.455 ;
        RECT 28.180 185.335 28.350 185.625 ;
        RECT 28.940 185.585 29.110 185.965 ;
        RECT 29.280 186.045 30.245 186.055 ;
        RECT 30.435 186.875 30.695 187.265 ;
        RECT 30.905 187.165 31.235 187.625 ;
        RECT 32.110 187.235 32.965 187.405 ;
        RECT 33.170 187.235 33.665 187.405 ;
        RECT 33.835 187.265 34.165 187.625 ;
        RECT 30.435 186.185 30.605 186.875 ;
        RECT 30.775 186.525 30.945 186.705 ;
        RECT 31.115 186.695 31.905 186.945 ;
        RECT 32.110 186.525 32.280 187.235 ;
        RECT 32.450 186.725 32.805 186.945 ;
        RECT 30.775 186.355 32.465 186.525 ;
        RECT 29.280 185.755 29.740 186.045 ;
        RECT 30.435 186.015 31.935 186.185 ;
        RECT 30.435 185.875 30.605 186.015 ;
        RECT 30.045 185.705 30.605 185.875 ;
        RECT 28.520 185.075 28.770 185.535 ;
        RECT 28.940 185.245 29.810 185.585 ;
        RECT 30.045 185.245 30.215 185.705 ;
        RECT 31.050 185.675 32.125 185.845 ;
        RECT 30.385 185.075 30.755 185.535 ;
        RECT 31.050 185.335 31.220 185.675 ;
        RECT 31.390 185.075 31.720 185.505 ;
        RECT 31.955 185.335 32.125 185.675 ;
        RECT 32.295 185.575 32.465 186.355 ;
        RECT 32.635 186.135 32.805 186.725 ;
        RECT 32.975 186.325 33.325 186.945 ;
        RECT 32.635 185.745 33.100 186.135 ;
        RECT 33.495 185.875 33.665 187.235 ;
        RECT 33.835 186.045 34.295 187.095 ;
        RECT 33.270 185.705 33.665 185.875 ;
        RECT 33.270 185.575 33.440 185.705 ;
        RECT 32.295 185.245 32.975 185.575 ;
        RECT 33.190 185.245 33.440 185.575 ;
        RECT 33.610 185.075 33.860 185.535 ;
        RECT 34.030 185.260 34.355 186.045 ;
        RECT 34.525 185.245 34.695 187.365 ;
        RECT 34.865 187.245 35.195 187.625 ;
        RECT 35.365 187.075 35.620 187.365 ;
        RECT 34.870 186.905 35.620 187.075 ;
        RECT 35.800 186.915 36.055 187.445 ;
        RECT 36.225 187.165 36.530 187.625 ;
        RECT 36.775 187.245 37.845 187.415 ;
        RECT 34.870 185.915 35.100 186.905 ;
        RECT 35.270 186.085 35.620 186.735 ;
        RECT 35.800 186.265 36.010 186.915 ;
        RECT 36.775 186.890 37.095 187.245 ;
        RECT 36.770 186.715 37.095 186.890 ;
        RECT 36.180 186.415 37.095 186.715 ;
        RECT 37.265 186.675 37.505 187.075 ;
        RECT 37.675 187.015 37.845 187.245 ;
        RECT 38.015 187.185 38.205 187.625 ;
        RECT 38.375 187.175 39.325 187.455 ;
        RECT 39.545 187.265 39.895 187.435 ;
        RECT 37.675 186.845 38.205 187.015 ;
        RECT 36.180 186.385 36.920 186.415 ;
        RECT 34.870 185.745 35.620 185.915 ;
        RECT 34.865 185.075 35.195 185.575 ;
        RECT 35.365 185.245 35.620 185.745 ;
        RECT 35.800 185.385 36.055 186.265 ;
        RECT 36.225 185.075 36.530 186.215 ;
        RECT 36.750 185.795 36.920 186.385 ;
        RECT 37.265 186.305 37.805 186.675 ;
        RECT 37.985 186.565 38.205 186.845 ;
        RECT 38.375 186.395 38.545 187.175 ;
        RECT 38.140 186.225 38.545 186.395 ;
        RECT 38.715 186.385 39.065 187.005 ;
        RECT 38.140 186.135 38.310 186.225 ;
        RECT 39.235 186.215 39.445 187.005 ;
        RECT 37.090 185.965 38.310 186.135 ;
        RECT 38.770 186.055 39.445 186.215 ;
        RECT 36.750 185.625 37.550 185.795 ;
        RECT 36.870 185.075 37.200 185.455 ;
        RECT 37.380 185.335 37.550 185.625 ;
        RECT 38.140 185.585 38.310 185.965 ;
        RECT 38.480 186.045 39.445 186.055 ;
        RECT 39.635 186.875 39.895 187.265 ;
        RECT 40.105 187.165 40.435 187.625 ;
        RECT 41.310 187.235 42.165 187.405 ;
        RECT 42.370 187.235 42.865 187.405 ;
        RECT 43.035 187.265 43.365 187.625 ;
        RECT 39.635 186.185 39.805 186.875 ;
        RECT 39.975 186.525 40.145 186.705 ;
        RECT 40.315 186.695 41.105 186.945 ;
        RECT 41.310 186.525 41.480 187.235 ;
        RECT 41.650 186.725 42.005 186.945 ;
        RECT 39.975 186.355 41.665 186.525 ;
        RECT 38.480 185.755 38.940 186.045 ;
        RECT 39.635 186.015 41.135 186.185 ;
        RECT 39.635 185.875 39.805 186.015 ;
        RECT 39.245 185.705 39.805 185.875 ;
        RECT 37.720 185.075 37.970 185.535 ;
        RECT 38.140 185.245 39.010 185.585 ;
        RECT 39.245 185.245 39.415 185.705 ;
        RECT 40.250 185.675 41.325 185.845 ;
        RECT 39.585 185.075 39.955 185.535 ;
        RECT 40.250 185.335 40.420 185.675 ;
        RECT 40.590 185.075 40.920 185.505 ;
        RECT 41.155 185.335 41.325 185.675 ;
        RECT 41.495 185.575 41.665 186.355 ;
        RECT 41.835 186.135 42.005 186.725 ;
        RECT 42.175 186.325 42.525 186.945 ;
        RECT 41.835 185.745 42.300 186.135 ;
        RECT 42.695 185.875 42.865 187.235 ;
        RECT 43.035 186.045 43.495 187.095 ;
        RECT 42.470 185.705 42.865 185.875 ;
        RECT 42.470 185.575 42.640 185.705 ;
        RECT 41.495 185.245 42.175 185.575 ;
        RECT 42.390 185.245 42.640 185.575 ;
        RECT 42.810 185.075 43.060 185.535 ;
        RECT 43.230 185.260 43.555 186.045 ;
        RECT 43.725 185.245 43.895 187.365 ;
        RECT 44.065 187.245 44.395 187.625 ;
        RECT 44.565 187.075 44.820 187.365 ;
        RECT 44.070 186.905 44.820 187.075 ;
        RECT 44.070 185.915 44.300 186.905 ;
        RECT 45.200 186.845 45.700 187.455 ;
        RECT 44.470 186.085 44.820 186.735 ;
        RECT 44.995 186.385 45.345 186.635 ;
        RECT 45.530 186.215 45.700 186.845 ;
        RECT 46.330 186.975 46.660 187.455 ;
        RECT 46.830 187.165 47.055 187.625 ;
        RECT 47.225 186.975 47.555 187.455 ;
        RECT 46.330 186.805 47.555 186.975 ;
        RECT 47.745 186.825 47.995 187.625 ;
        RECT 48.165 186.825 48.505 187.455 ;
        RECT 48.675 186.900 48.965 187.625 ;
        RECT 50.145 187.075 50.315 187.455 ;
        RECT 50.495 187.245 50.825 187.625 ;
        RECT 50.145 186.905 50.810 187.075 ;
        RECT 51.005 186.950 51.265 187.455 ;
        RECT 45.870 186.435 46.200 186.635 ;
        RECT 46.370 186.435 46.700 186.635 ;
        RECT 46.870 186.435 47.290 186.635 ;
        RECT 47.465 186.465 48.160 186.635 ;
        RECT 47.465 186.215 47.635 186.465 ;
        RECT 48.330 186.215 48.505 186.825 ;
        RECT 50.075 186.355 50.405 186.725 ;
        RECT 50.640 186.650 50.810 186.905 ;
        RECT 50.640 186.320 50.925 186.650 ;
        RECT 45.200 186.045 47.635 186.215 ;
        RECT 44.070 185.745 44.820 185.915 ;
        RECT 44.065 185.075 44.395 185.575 ;
        RECT 44.565 185.245 44.820 185.745 ;
        RECT 45.200 185.245 45.530 186.045 ;
        RECT 45.700 185.075 46.030 185.875 ;
        RECT 46.330 185.245 46.660 186.045 ;
        RECT 47.305 185.075 47.555 185.875 ;
        RECT 47.825 185.075 47.995 186.215 ;
        RECT 48.165 185.245 48.505 186.215 ;
        RECT 48.675 185.075 48.965 186.240 ;
        RECT 50.640 186.175 50.810 186.320 ;
        RECT 50.145 186.005 50.810 186.175 ;
        RECT 51.095 186.150 51.265 186.950 ;
        RECT 50.145 185.245 50.315 186.005 ;
        RECT 50.495 185.075 50.825 185.835 ;
        RECT 50.995 185.245 51.265 186.150 ;
        RECT 51.440 186.885 51.695 187.455 ;
        RECT 51.865 187.225 52.195 187.625 ;
        RECT 52.620 187.090 53.150 187.455 ;
        RECT 52.620 187.055 52.795 187.090 ;
        RECT 51.865 186.885 52.795 187.055 ;
        RECT 53.340 186.945 53.615 187.455 ;
        RECT 51.440 186.215 51.610 186.885 ;
        RECT 51.865 186.715 52.035 186.885 ;
        RECT 51.780 186.385 52.035 186.715 ;
        RECT 52.260 186.385 52.455 186.715 ;
        RECT 51.440 185.245 51.775 186.215 ;
        RECT 51.945 185.075 52.115 186.215 ;
        RECT 52.285 185.415 52.455 186.385 ;
        RECT 52.625 185.755 52.795 186.885 ;
        RECT 52.965 186.095 53.135 186.895 ;
        RECT 53.335 186.775 53.615 186.945 ;
        RECT 53.340 186.295 53.615 186.775 ;
        RECT 53.785 186.095 53.975 187.455 ;
        RECT 54.155 187.090 54.665 187.625 ;
        RECT 54.885 186.815 55.130 187.420 ;
        RECT 55.580 186.885 55.835 187.455 ;
        RECT 56.005 187.225 56.335 187.625 ;
        RECT 56.760 187.090 57.290 187.455 ;
        RECT 56.760 187.055 56.935 187.090 ;
        RECT 56.005 186.885 56.935 187.055 ;
        RECT 54.175 186.645 55.405 186.815 ;
        RECT 52.965 185.925 53.975 186.095 ;
        RECT 54.145 186.080 54.895 186.270 ;
        RECT 52.625 185.585 53.750 185.755 ;
        RECT 54.145 185.415 54.315 186.080 ;
        RECT 55.065 185.835 55.405 186.645 ;
        RECT 52.285 185.245 54.315 185.415 ;
        RECT 54.485 185.075 54.655 185.835 ;
        RECT 54.890 185.425 55.405 185.835 ;
        RECT 55.580 186.215 55.750 186.885 ;
        RECT 56.005 186.715 56.175 186.885 ;
        RECT 55.920 186.385 56.175 186.715 ;
        RECT 56.400 186.385 56.595 186.715 ;
        RECT 55.580 185.245 55.915 186.215 ;
        RECT 56.085 185.075 56.255 186.215 ;
        RECT 56.425 185.415 56.595 186.385 ;
        RECT 56.765 185.755 56.935 186.885 ;
        RECT 57.105 186.095 57.275 186.895 ;
        RECT 57.480 186.605 57.755 187.455 ;
        RECT 57.475 186.435 57.755 186.605 ;
        RECT 57.480 186.295 57.755 186.435 ;
        RECT 57.925 186.095 58.115 187.455 ;
        RECT 58.295 187.090 58.805 187.625 ;
        RECT 59.025 186.815 59.270 187.420 ;
        RECT 58.315 186.645 59.545 186.815 ;
        RECT 59.775 186.805 59.985 187.625 ;
        RECT 60.155 186.825 60.485 187.455 ;
        RECT 57.105 185.925 58.115 186.095 ;
        RECT 58.285 186.080 59.035 186.270 ;
        RECT 56.765 185.585 57.890 185.755 ;
        RECT 58.285 185.415 58.455 186.080 ;
        RECT 59.205 185.835 59.545 186.645 ;
        RECT 60.155 186.225 60.405 186.825 ;
        RECT 60.655 186.805 60.885 187.625 ;
        RECT 62.015 186.950 62.275 187.455 ;
        RECT 62.455 187.245 62.785 187.625 ;
        RECT 62.965 187.075 63.135 187.455 ;
        RECT 64.125 187.230 64.455 187.625 ;
        RECT 60.575 186.385 60.905 186.635 ;
        RECT 56.425 185.245 58.455 185.415 ;
        RECT 58.625 185.075 58.795 185.835 ;
        RECT 59.030 185.425 59.545 185.835 ;
        RECT 59.775 185.075 59.985 186.215 ;
        RECT 60.155 185.245 60.485 186.225 ;
        RECT 60.655 185.075 60.885 186.215 ;
        RECT 62.015 186.150 62.185 186.950 ;
        RECT 62.470 186.905 63.135 187.075 ;
        RECT 64.625 187.055 64.825 187.410 ;
        RECT 64.995 187.225 65.325 187.625 ;
        RECT 65.495 187.055 65.695 187.400 ;
        RECT 62.470 186.650 62.640 186.905 ;
        RECT 63.855 186.885 65.695 187.055 ;
        RECT 65.865 186.885 66.195 187.625 ;
        RECT 66.430 187.055 66.600 187.305 ;
        RECT 67.075 187.125 67.335 187.455 ;
        RECT 67.645 187.245 67.975 187.625 ;
        RECT 68.155 187.285 69.635 187.455 ;
        RECT 66.430 186.885 66.905 187.055 ;
        RECT 62.355 186.320 62.640 186.650 ;
        RECT 62.875 186.355 63.205 186.725 ;
        RECT 62.470 186.175 62.640 186.320 ;
        RECT 62.015 185.245 62.285 186.150 ;
        RECT 62.470 186.005 63.135 186.175 ;
        RECT 62.455 185.075 62.785 185.835 ;
        RECT 62.965 185.245 63.135 186.005 ;
        RECT 63.855 185.260 64.115 186.885 ;
        RECT 64.295 185.915 64.515 186.715 ;
        RECT 64.755 186.095 65.055 186.715 ;
        RECT 65.225 186.095 65.555 186.715 ;
        RECT 65.725 186.095 66.045 186.715 ;
        RECT 66.215 186.095 66.565 186.715 ;
        RECT 66.735 185.915 66.905 186.885 ;
        RECT 64.295 185.705 66.905 185.915 ;
        RECT 67.075 186.425 67.245 187.125 ;
        RECT 68.155 186.955 68.555 187.285 ;
        RECT 67.595 186.765 67.805 186.945 ;
        RECT 67.595 186.595 68.215 186.765 ;
        RECT 68.385 186.475 68.555 186.955 ;
        RECT 68.745 186.785 69.295 187.115 ;
        RECT 67.075 186.255 68.205 186.425 ;
        RECT 68.385 186.305 68.955 186.475 ;
        RECT 67.075 185.575 67.245 186.255 ;
        RECT 68.035 186.135 68.205 186.255 ;
        RECT 67.415 185.755 67.765 186.085 ;
        RECT 68.035 185.965 68.615 186.135 ;
        RECT 68.785 185.795 68.955 186.305 ;
        RECT 68.215 185.625 68.955 185.795 ;
        RECT 69.125 185.795 69.295 186.785 ;
        RECT 69.465 186.385 69.635 187.285 ;
        RECT 69.885 186.715 70.070 187.295 ;
        RECT 70.340 186.715 70.535 187.290 ;
        RECT 70.745 187.245 71.075 187.625 ;
        RECT 69.885 186.385 70.115 186.715 ;
        RECT 70.340 186.385 70.595 186.715 ;
        RECT 69.885 186.075 70.070 186.385 ;
        RECT 70.340 186.075 70.535 186.385 ;
        RECT 70.905 185.795 71.075 186.715 ;
        RECT 69.125 185.625 71.075 185.795 ;
        RECT 65.865 185.075 66.195 185.525 ;
        RECT 67.075 185.245 67.335 185.575 ;
        RECT 67.645 185.075 67.975 185.455 ;
        RECT 68.215 185.245 68.405 185.625 ;
        RECT 68.655 185.075 68.985 185.455 ;
        RECT 69.195 185.245 69.365 185.625 ;
        RECT 69.560 185.075 69.890 185.455 ;
        RECT 70.150 185.245 70.320 185.625 ;
        RECT 70.745 185.075 71.075 185.455 ;
        RECT 71.245 185.245 71.505 187.455 ;
        RECT 71.675 187.125 71.975 187.455 ;
        RECT 72.145 187.145 72.420 187.625 ;
        RECT 71.675 186.215 71.845 187.125 ;
        RECT 72.600 186.975 72.895 187.365 ;
        RECT 73.065 187.145 73.320 187.625 ;
        RECT 73.495 186.975 73.755 187.365 ;
        RECT 73.925 187.145 74.205 187.625 ;
        RECT 72.015 186.385 72.365 186.955 ;
        RECT 72.600 186.805 74.250 186.975 ;
        RECT 74.435 186.900 74.725 187.625 ;
        RECT 75.855 186.805 76.085 187.625 ;
        RECT 76.255 186.825 76.585 187.455 ;
        RECT 72.535 186.465 73.675 186.635 ;
        RECT 72.535 186.215 72.705 186.465 ;
        RECT 73.845 186.295 74.250 186.805 ;
        RECT 75.835 186.385 76.165 186.635 ;
        RECT 71.675 186.045 72.705 186.215 ;
        RECT 73.495 186.125 74.250 186.295 ;
        RECT 71.675 185.245 71.985 186.045 ;
        RECT 73.495 185.875 73.755 186.125 ;
        RECT 72.155 185.075 72.465 185.875 ;
        RECT 72.635 185.705 73.755 185.875 ;
        RECT 72.635 185.245 72.895 185.705 ;
        RECT 73.065 185.075 73.320 185.535 ;
        RECT 73.495 185.245 73.755 185.705 ;
        RECT 73.925 185.075 74.210 185.945 ;
        RECT 74.435 185.075 74.725 186.240 ;
        RECT 76.335 186.225 76.585 186.825 ;
        RECT 76.755 186.805 76.965 187.625 ;
        RECT 77.570 186.915 77.825 187.445 ;
        RECT 78.005 187.165 78.290 187.625 ;
        RECT 75.855 185.075 76.085 186.215 ;
        RECT 76.255 185.245 76.585 186.225 ;
        RECT 76.755 185.075 76.965 186.215 ;
        RECT 77.570 186.055 77.750 186.915 ;
        RECT 78.470 186.715 78.720 187.365 ;
        RECT 77.920 186.385 78.720 186.715 ;
        RECT 77.570 185.585 77.825 186.055 ;
        RECT 77.485 185.415 77.825 185.585 ;
        RECT 77.570 185.385 77.825 185.415 ;
        RECT 78.005 185.075 78.290 185.875 ;
        RECT 78.470 185.795 78.720 186.385 ;
        RECT 78.920 187.030 79.240 187.360 ;
        RECT 79.420 187.145 80.080 187.625 ;
        RECT 80.280 187.235 81.130 187.405 ;
        RECT 78.920 186.135 79.110 187.030 ;
        RECT 79.430 186.705 80.090 186.975 ;
        RECT 79.760 186.645 80.090 186.705 ;
        RECT 79.280 186.475 79.610 186.535 ;
        RECT 80.280 186.475 80.450 187.235 ;
        RECT 81.690 187.165 82.010 187.625 ;
        RECT 82.210 186.985 82.460 187.415 ;
        RECT 82.750 187.185 83.160 187.625 ;
        RECT 83.330 187.245 84.345 187.445 ;
        RECT 80.620 186.815 81.870 186.985 ;
        RECT 80.620 186.695 80.950 186.815 ;
        RECT 79.280 186.305 81.180 186.475 ;
        RECT 78.920 185.965 80.840 186.135 ;
        RECT 78.920 185.945 79.240 185.965 ;
        RECT 78.470 185.285 78.800 185.795 ;
        RECT 79.070 185.335 79.240 185.945 ;
        RECT 81.010 185.795 81.180 186.305 ;
        RECT 81.350 186.235 81.530 186.645 ;
        RECT 81.700 186.055 81.870 186.815 ;
        RECT 79.410 185.075 79.740 185.765 ;
        RECT 79.970 185.625 81.180 185.795 ;
        RECT 81.350 185.745 81.870 186.055 ;
        RECT 82.040 186.645 82.460 186.985 ;
        RECT 82.750 186.645 83.160 186.975 ;
        RECT 82.040 185.875 82.230 186.645 ;
        RECT 83.330 186.515 83.500 187.245 ;
        RECT 84.645 187.075 84.815 187.405 ;
        RECT 84.985 187.245 85.315 187.625 ;
        RECT 83.670 186.695 84.020 187.065 ;
        RECT 83.330 186.475 83.750 186.515 ;
        RECT 82.400 186.305 83.750 186.475 ;
        RECT 82.400 186.145 82.650 186.305 ;
        RECT 83.160 185.875 83.410 186.135 ;
        RECT 82.040 185.625 83.410 185.875 ;
        RECT 79.970 185.335 80.210 185.625 ;
        RECT 81.010 185.545 81.180 185.625 ;
        RECT 80.410 185.075 80.830 185.455 ;
        RECT 81.010 185.295 81.640 185.545 ;
        RECT 82.110 185.075 82.440 185.455 ;
        RECT 82.610 185.335 82.780 185.625 ;
        RECT 83.580 185.460 83.750 186.305 ;
        RECT 84.200 186.135 84.420 187.005 ;
        RECT 84.645 186.885 85.340 187.075 ;
        RECT 83.920 185.755 84.420 186.135 ;
        RECT 84.590 186.085 85.000 186.705 ;
        RECT 85.170 185.915 85.340 186.885 ;
        RECT 84.645 185.745 85.340 185.915 ;
        RECT 82.960 185.075 83.340 185.455 ;
        RECT 83.580 185.290 84.410 185.460 ;
        RECT 84.645 185.245 84.815 185.745 ;
        RECT 84.985 185.075 85.315 185.575 ;
        RECT 85.530 185.245 85.755 187.365 ;
        RECT 85.925 187.245 86.255 187.625 ;
        RECT 86.425 187.075 86.595 187.365 ;
        RECT 85.930 186.905 86.595 187.075 ;
        RECT 85.930 185.915 86.160 186.905 ;
        RECT 86.895 186.805 87.125 187.625 ;
        RECT 87.295 186.825 87.625 187.455 ;
        RECT 86.330 186.085 86.680 186.735 ;
        RECT 86.875 186.385 87.205 186.635 ;
        RECT 87.375 186.225 87.625 186.825 ;
        RECT 87.795 186.805 88.005 187.625 ;
        RECT 88.240 186.915 88.495 187.445 ;
        RECT 88.665 187.165 88.970 187.625 ;
        RECT 89.215 187.245 90.285 187.415 ;
        RECT 85.930 185.745 86.595 185.915 ;
        RECT 85.925 185.075 86.255 185.575 ;
        RECT 86.425 185.245 86.595 185.745 ;
        RECT 86.895 185.075 87.125 186.215 ;
        RECT 87.295 185.245 87.625 186.225 ;
        RECT 88.240 186.265 88.450 186.915 ;
        RECT 89.215 186.890 89.535 187.245 ;
        RECT 89.210 186.715 89.535 186.890 ;
        RECT 88.620 186.415 89.535 186.715 ;
        RECT 89.705 186.675 89.945 187.075 ;
        RECT 90.115 187.015 90.285 187.245 ;
        RECT 90.455 187.185 90.645 187.625 ;
        RECT 90.815 187.175 91.765 187.455 ;
        RECT 91.985 187.265 92.335 187.435 ;
        RECT 90.115 186.845 90.645 187.015 ;
        RECT 88.620 186.385 89.360 186.415 ;
        RECT 87.795 185.075 88.005 186.215 ;
        RECT 88.240 185.385 88.495 186.265 ;
        RECT 88.665 185.075 88.970 186.215 ;
        RECT 89.190 185.795 89.360 186.385 ;
        RECT 89.705 186.305 90.245 186.675 ;
        RECT 90.425 186.565 90.645 186.845 ;
        RECT 90.815 186.395 90.985 187.175 ;
        RECT 90.580 186.225 90.985 186.395 ;
        RECT 91.155 186.385 91.505 187.005 ;
        RECT 90.580 186.135 90.750 186.225 ;
        RECT 91.675 186.215 91.885 187.005 ;
        RECT 89.530 185.965 90.750 186.135 ;
        RECT 91.210 186.055 91.885 186.215 ;
        RECT 89.190 185.625 89.990 185.795 ;
        RECT 89.310 185.075 89.640 185.455 ;
        RECT 89.820 185.335 89.990 185.625 ;
        RECT 90.580 185.585 90.750 185.965 ;
        RECT 90.920 186.045 91.885 186.055 ;
        RECT 92.075 186.875 92.335 187.265 ;
        RECT 92.545 187.165 92.875 187.625 ;
        RECT 93.750 187.235 94.605 187.405 ;
        RECT 94.810 187.235 95.305 187.405 ;
        RECT 95.475 187.265 95.805 187.625 ;
        RECT 92.075 186.185 92.245 186.875 ;
        RECT 92.415 186.525 92.585 186.705 ;
        RECT 92.755 186.695 93.545 186.945 ;
        RECT 93.750 186.525 93.920 187.235 ;
        RECT 94.090 186.725 94.445 186.945 ;
        RECT 92.415 186.355 94.105 186.525 ;
        RECT 90.920 185.755 91.380 186.045 ;
        RECT 92.075 186.015 93.575 186.185 ;
        RECT 92.075 185.875 92.245 186.015 ;
        RECT 91.685 185.705 92.245 185.875 ;
        RECT 90.160 185.075 90.410 185.535 ;
        RECT 90.580 185.245 91.450 185.585 ;
        RECT 91.685 185.245 91.855 185.705 ;
        RECT 92.690 185.675 93.765 185.845 ;
        RECT 92.025 185.075 92.395 185.535 ;
        RECT 92.690 185.335 92.860 185.675 ;
        RECT 93.030 185.075 93.360 185.505 ;
        RECT 93.595 185.335 93.765 185.675 ;
        RECT 93.935 185.575 94.105 186.355 ;
        RECT 94.275 186.135 94.445 186.725 ;
        RECT 94.615 186.325 94.965 186.945 ;
        RECT 94.275 185.745 94.740 186.135 ;
        RECT 95.135 185.875 95.305 187.235 ;
        RECT 95.475 186.045 95.935 187.095 ;
        RECT 94.910 185.705 95.305 185.875 ;
        RECT 94.910 185.575 95.080 185.705 ;
        RECT 93.935 185.245 94.615 185.575 ;
        RECT 94.830 185.245 95.080 185.575 ;
        RECT 95.250 185.075 95.500 185.535 ;
        RECT 95.670 185.260 95.995 186.045 ;
        RECT 96.165 185.245 96.335 187.365 ;
        RECT 96.505 187.245 96.835 187.625 ;
        RECT 97.005 187.075 97.260 187.365 ;
        RECT 96.510 186.905 97.260 187.075 ;
        RECT 96.510 185.915 96.740 186.905 ;
        RECT 97.475 186.805 97.705 187.625 ;
        RECT 97.875 186.825 98.205 187.455 ;
        RECT 96.910 186.085 97.260 186.735 ;
        RECT 97.455 186.385 97.785 186.635 ;
        RECT 97.955 186.225 98.205 186.825 ;
        RECT 98.375 186.805 98.585 187.625 ;
        RECT 98.855 186.805 99.085 187.625 ;
        RECT 99.255 186.825 99.585 187.455 ;
        RECT 98.835 186.385 99.165 186.635 ;
        RECT 99.335 186.225 99.585 186.825 ;
        RECT 99.755 186.805 99.965 187.625 ;
        RECT 100.195 186.900 100.485 187.625 ;
        RECT 101.580 186.915 101.835 187.445 ;
        RECT 102.005 187.165 102.310 187.625 ;
        RECT 102.555 187.245 103.625 187.415 ;
        RECT 101.580 186.265 101.790 186.915 ;
        RECT 102.555 186.890 102.875 187.245 ;
        RECT 102.550 186.715 102.875 186.890 ;
        RECT 101.960 186.415 102.875 186.715 ;
        RECT 103.045 186.675 103.285 187.075 ;
        RECT 103.455 187.015 103.625 187.245 ;
        RECT 103.795 187.185 103.985 187.625 ;
        RECT 104.155 187.175 105.105 187.455 ;
        RECT 105.325 187.265 105.675 187.435 ;
        RECT 103.455 186.845 103.985 187.015 ;
        RECT 101.960 186.385 102.700 186.415 ;
        RECT 96.510 185.745 97.260 185.915 ;
        RECT 96.505 185.075 96.835 185.575 ;
        RECT 97.005 185.245 97.260 185.745 ;
        RECT 97.475 185.075 97.705 186.215 ;
        RECT 97.875 185.245 98.205 186.225 ;
        RECT 98.375 185.075 98.585 186.215 ;
        RECT 98.855 185.075 99.085 186.215 ;
        RECT 99.255 185.245 99.585 186.225 ;
        RECT 99.755 185.075 99.965 186.215 ;
        RECT 100.195 185.075 100.485 186.240 ;
        RECT 101.580 185.385 101.835 186.265 ;
        RECT 102.005 185.075 102.310 186.215 ;
        RECT 102.530 185.795 102.700 186.385 ;
        RECT 103.045 186.305 103.585 186.675 ;
        RECT 103.765 186.565 103.985 186.845 ;
        RECT 104.155 186.395 104.325 187.175 ;
        RECT 103.920 186.225 104.325 186.395 ;
        RECT 104.495 186.385 104.845 187.005 ;
        RECT 103.920 186.135 104.090 186.225 ;
        RECT 105.015 186.215 105.225 187.005 ;
        RECT 102.870 185.965 104.090 186.135 ;
        RECT 104.550 186.055 105.225 186.215 ;
        RECT 102.530 185.625 103.330 185.795 ;
        RECT 102.650 185.075 102.980 185.455 ;
        RECT 103.160 185.335 103.330 185.625 ;
        RECT 103.920 185.585 104.090 185.965 ;
        RECT 104.260 186.045 105.225 186.055 ;
        RECT 105.415 186.875 105.675 187.265 ;
        RECT 105.885 187.165 106.215 187.625 ;
        RECT 107.090 187.235 107.945 187.405 ;
        RECT 108.150 187.235 108.645 187.405 ;
        RECT 108.815 187.265 109.145 187.625 ;
        RECT 105.415 186.185 105.585 186.875 ;
        RECT 105.755 186.525 105.925 186.705 ;
        RECT 106.095 186.695 106.885 186.945 ;
        RECT 107.090 186.525 107.260 187.235 ;
        RECT 107.430 186.725 107.785 186.945 ;
        RECT 105.755 186.355 107.445 186.525 ;
        RECT 104.260 185.755 104.720 186.045 ;
        RECT 105.415 186.015 106.915 186.185 ;
        RECT 105.415 185.875 105.585 186.015 ;
        RECT 105.025 185.705 105.585 185.875 ;
        RECT 103.500 185.075 103.750 185.535 ;
        RECT 103.920 185.245 104.790 185.585 ;
        RECT 105.025 185.245 105.195 185.705 ;
        RECT 106.030 185.675 107.105 185.845 ;
        RECT 105.365 185.075 105.735 185.535 ;
        RECT 106.030 185.335 106.200 185.675 ;
        RECT 106.370 185.075 106.700 185.505 ;
        RECT 106.935 185.335 107.105 185.675 ;
        RECT 107.275 185.575 107.445 186.355 ;
        RECT 107.615 186.135 107.785 186.725 ;
        RECT 107.955 186.325 108.305 186.945 ;
        RECT 107.615 185.745 108.080 186.135 ;
        RECT 108.475 185.875 108.645 187.235 ;
        RECT 108.815 186.045 109.275 187.095 ;
        RECT 108.250 185.705 108.645 185.875 ;
        RECT 108.250 185.575 108.420 185.705 ;
        RECT 107.275 185.245 107.955 185.575 ;
        RECT 108.170 185.245 108.420 185.575 ;
        RECT 108.590 185.075 108.840 185.535 ;
        RECT 109.010 185.260 109.335 186.045 ;
        RECT 109.505 185.245 109.675 187.365 ;
        RECT 109.845 187.245 110.175 187.625 ;
        RECT 110.345 187.075 110.600 187.365 ;
        RECT 109.850 186.905 110.600 187.075 ;
        RECT 109.850 185.915 110.080 186.905 ;
        RECT 110.815 186.805 111.045 187.625 ;
        RECT 111.215 186.825 111.545 187.455 ;
        RECT 110.250 186.085 110.600 186.735 ;
        RECT 110.795 186.385 111.125 186.635 ;
        RECT 111.295 186.225 111.545 186.825 ;
        RECT 111.715 186.805 111.925 187.625 ;
        RECT 112.155 186.875 113.365 187.625 ;
        RECT 109.850 185.745 110.600 185.915 ;
        RECT 109.845 185.075 110.175 185.575 ;
        RECT 110.345 185.245 110.600 185.745 ;
        RECT 110.815 185.075 111.045 186.215 ;
        RECT 111.215 185.245 111.545 186.225 ;
        RECT 111.715 185.075 111.925 186.215 ;
        RECT 112.155 186.165 112.675 186.705 ;
        RECT 112.845 186.335 113.365 186.875 ;
        RECT 112.155 185.075 113.365 186.165 ;
        RECT 22.830 184.905 113.450 185.075 ;
        RECT 22.915 183.815 24.125 184.905 ;
        RECT 22.915 183.105 23.435 183.645 ;
        RECT 23.605 183.275 24.125 183.815 ;
        RECT 25.275 183.765 25.485 184.905 ;
        RECT 25.655 183.755 25.985 184.735 ;
        RECT 26.155 183.765 26.385 184.905 ;
        RECT 22.915 182.355 24.125 183.105 ;
        RECT 25.275 182.355 25.485 183.175 ;
        RECT 25.655 183.155 25.905 183.755 ;
        RECT 26.600 183.715 26.855 184.595 ;
        RECT 27.025 183.765 27.330 184.905 ;
        RECT 27.670 184.525 28.000 184.905 ;
        RECT 28.180 184.355 28.350 184.645 ;
        RECT 28.520 184.445 28.770 184.905 ;
        RECT 27.550 184.185 28.350 184.355 ;
        RECT 28.940 184.395 29.810 184.735 ;
        RECT 26.075 183.345 26.405 183.595 ;
        RECT 25.655 182.525 25.985 183.155 ;
        RECT 26.155 182.355 26.385 183.175 ;
        RECT 26.600 183.065 26.810 183.715 ;
        RECT 27.550 183.595 27.720 184.185 ;
        RECT 28.940 184.015 29.110 184.395 ;
        RECT 30.045 184.275 30.215 184.735 ;
        RECT 30.385 184.445 30.755 184.905 ;
        RECT 31.050 184.305 31.220 184.645 ;
        RECT 31.390 184.475 31.720 184.905 ;
        RECT 31.955 184.305 32.125 184.645 ;
        RECT 27.890 183.845 29.110 184.015 ;
        RECT 29.280 183.935 29.740 184.225 ;
        RECT 30.045 184.105 30.605 184.275 ;
        RECT 31.050 184.135 32.125 184.305 ;
        RECT 32.295 184.405 32.975 184.735 ;
        RECT 33.190 184.405 33.440 184.735 ;
        RECT 33.610 184.445 33.860 184.905 ;
        RECT 30.435 183.965 30.605 184.105 ;
        RECT 29.280 183.925 30.245 183.935 ;
        RECT 28.940 183.755 29.110 183.845 ;
        RECT 29.570 183.765 30.245 183.925 ;
        RECT 26.980 183.565 27.720 183.595 ;
        RECT 26.980 183.265 27.895 183.565 ;
        RECT 27.570 183.090 27.895 183.265 ;
        RECT 26.600 182.535 26.855 183.065 ;
        RECT 27.025 182.355 27.330 182.815 ;
        RECT 27.575 182.735 27.895 183.090 ;
        RECT 28.065 183.305 28.605 183.675 ;
        RECT 28.940 183.585 29.345 183.755 ;
        RECT 28.065 182.905 28.305 183.305 ;
        RECT 28.785 183.135 29.005 183.415 ;
        RECT 28.475 182.965 29.005 183.135 ;
        RECT 28.475 182.735 28.645 182.965 ;
        RECT 29.175 182.805 29.345 183.585 ;
        RECT 29.515 182.975 29.865 183.595 ;
        RECT 30.035 182.975 30.245 183.765 ;
        RECT 30.435 183.795 31.935 183.965 ;
        RECT 30.435 183.105 30.605 183.795 ;
        RECT 32.295 183.625 32.465 184.405 ;
        RECT 33.270 184.275 33.440 184.405 ;
        RECT 30.775 183.455 32.465 183.625 ;
        RECT 32.635 183.845 33.100 184.235 ;
        RECT 33.270 184.105 33.665 184.275 ;
        RECT 30.775 183.275 30.945 183.455 ;
        RECT 27.575 182.565 28.645 182.735 ;
        RECT 28.815 182.355 29.005 182.795 ;
        RECT 29.175 182.525 30.125 182.805 ;
        RECT 30.435 182.715 30.695 183.105 ;
        RECT 31.115 183.035 31.905 183.285 ;
        RECT 30.345 182.545 30.695 182.715 ;
        RECT 30.905 182.355 31.235 182.815 ;
        RECT 32.110 182.745 32.280 183.455 ;
        RECT 32.635 183.255 32.805 183.845 ;
        RECT 32.450 183.035 32.805 183.255 ;
        RECT 32.975 183.035 33.325 183.655 ;
        RECT 33.495 182.745 33.665 184.105 ;
        RECT 34.030 183.935 34.355 184.720 ;
        RECT 33.835 182.885 34.295 183.935 ;
        RECT 32.110 182.575 32.965 182.745 ;
        RECT 33.170 182.575 33.665 182.745 ;
        RECT 33.835 182.355 34.165 182.715 ;
        RECT 34.525 182.615 34.695 184.735 ;
        RECT 34.865 184.405 35.195 184.905 ;
        RECT 35.365 184.235 35.620 184.735 ;
        RECT 34.870 184.065 35.620 184.235 ;
        RECT 34.870 183.075 35.100 184.065 ;
        RECT 35.270 183.245 35.620 183.895 ;
        RECT 35.795 183.740 36.085 184.905 ;
        RECT 36.920 183.935 37.250 184.735 ;
        RECT 37.420 184.105 37.750 184.905 ;
        RECT 38.050 183.935 38.380 184.735 ;
        RECT 39.025 184.105 39.275 184.905 ;
        RECT 36.920 183.765 39.355 183.935 ;
        RECT 39.545 183.765 39.715 184.905 ;
        RECT 39.885 183.765 40.225 184.735 ;
        RECT 36.715 183.345 37.065 183.595 ;
        RECT 37.250 183.135 37.420 183.765 ;
        RECT 37.590 183.345 37.920 183.545 ;
        RECT 38.090 183.345 38.420 183.545 ;
        RECT 38.590 183.345 39.010 183.545 ;
        RECT 39.185 183.515 39.355 183.765 ;
        RECT 39.185 183.345 39.880 183.515 ;
        RECT 34.870 182.905 35.620 183.075 ;
        RECT 34.865 182.355 35.195 182.735 ;
        RECT 35.365 182.615 35.620 182.905 ;
        RECT 35.795 182.355 36.085 183.080 ;
        RECT 36.920 182.525 37.420 183.135 ;
        RECT 38.050 183.005 39.275 183.175 ;
        RECT 40.050 183.155 40.225 183.765 ;
        RECT 38.050 182.525 38.380 183.005 ;
        RECT 38.550 182.355 38.775 182.815 ;
        RECT 38.945 182.525 39.275 183.005 ;
        RECT 39.465 182.355 39.715 183.155 ;
        RECT 39.885 182.525 40.225 183.155 ;
        RECT 40.400 183.765 40.735 184.735 ;
        RECT 40.905 183.765 41.075 184.905 ;
        RECT 41.245 184.565 43.275 184.735 ;
        RECT 40.400 183.095 40.570 183.765 ;
        RECT 41.245 183.595 41.415 184.565 ;
        RECT 40.740 183.265 40.995 183.595 ;
        RECT 41.220 183.265 41.415 183.595 ;
        RECT 41.585 184.225 42.710 184.395 ;
        RECT 40.825 183.095 40.995 183.265 ;
        RECT 41.585 183.095 41.755 184.225 ;
        RECT 40.400 182.525 40.655 183.095 ;
        RECT 40.825 182.925 41.755 183.095 ;
        RECT 41.925 183.885 42.935 184.055 ;
        RECT 41.925 183.085 42.095 183.885 ;
        RECT 42.300 183.545 42.575 183.685 ;
        RECT 42.295 183.375 42.575 183.545 ;
        RECT 41.580 182.890 41.755 182.925 ;
        RECT 40.825 182.355 41.155 182.755 ;
        RECT 41.580 182.525 42.110 182.890 ;
        RECT 42.300 182.525 42.575 183.375 ;
        RECT 42.745 182.525 42.935 183.885 ;
        RECT 43.105 183.900 43.275 184.565 ;
        RECT 43.445 184.145 43.615 184.905 ;
        RECT 43.850 184.145 44.365 184.555 ;
        RECT 43.105 183.710 43.855 183.900 ;
        RECT 44.025 183.335 44.365 184.145 ;
        RECT 43.135 183.165 44.365 183.335 ;
        RECT 44.995 183.815 46.665 184.905 ;
        RECT 44.995 183.295 45.745 183.815 ;
        RECT 46.840 183.765 47.175 184.735 ;
        RECT 47.345 183.765 47.515 184.905 ;
        RECT 47.685 184.565 49.715 184.735 ;
        RECT 43.115 182.355 43.625 182.890 ;
        RECT 43.845 182.560 44.090 183.165 ;
        RECT 45.915 183.125 46.665 183.645 ;
        RECT 44.995 182.355 46.665 183.125 ;
        RECT 46.840 183.095 47.010 183.765 ;
        RECT 47.685 183.595 47.855 184.565 ;
        RECT 47.180 183.265 47.435 183.595 ;
        RECT 47.660 183.265 47.855 183.595 ;
        RECT 48.025 184.225 49.150 184.395 ;
        RECT 47.265 183.095 47.435 183.265 ;
        RECT 48.025 183.095 48.195 184.225 ;
        RECT 46.840 182.525 47.095 183.095 ;
        RECT 47.265 182.925 48.195 183.095 ;
        RECT 48.365 183.885 49.375 184.055 ;
        RECT 48.365 183.085 48.535 183.885 ;
        RECT 48.740 183.545 49.015 183.685 ;
        RECT 48.735 183.375 49.015 183.545 ;
        RECT 48.020 182.890 48.195 182.925 ;
        RECT 47.265 182.355 47.595 182.755 ;
        RECT 48.020 182.525 48.550 182.890 ;
        RECT 48.740 182.525 49.015 183.375 ;
        RECT 49.185 182.525 49.375 183.885 ;
        RECT 49.545 183.900 49.715 184.565 ;
        RECT 49.885 184.145 50.055 184.905 ;
        RECT 50.290 184.145 50.805 184.555 ;
        RECT 49.545 183.710 50.295 183.900 ;
        RECT 50.465 183.335 50.805 184.145 ;
        RECT 49.575 183.165 50.805 183.335 ;
        RECT 50.975 183.815 52.185 184.905 ;
        RECT 50.975 183.275 51.495 183.815 ;
        RECT 52.360 183.715 52.615 184.595 ;
        RECT 52.785 183.765 53.090 184.905 ;
        RECT 53.430 184.525 53.760 184.905 ;
        RECT 53.940 184.355 54.110 184.645 ;
        RECT 54.280 184.445 54.530 184.905 ;
        RECT 53.310 184.185 54.110 184.355 ;
        RECT 54.700 184.395 55.570 184.735 ;
        RECT 49.555 182.355 50.065 182.890 ;
        RECT 50.285 182.560 50.530 183.165 ;
        RECT 51.665 183.105 52.185 183.645 ;
        RECT 50.975 182.355 52.185 183.105 ;
        RECT 52.360 183.065 52.570 183.715 ;
        RECT 53.310 183.595 53.480 184.185 ;
        RECT 54.700 184.015 54.870 184.395 ;
        RECT 55.805 184.275 55.975 184.735 ;
        RECT 56.145 184.445 56.515 184.905 ;
        RECT 56.810 184.305 56.980 184.645 ;
        RECT 57.150 184.475 57.480 184.905 ;
        RECT 57.715 184.305 57.885 184.645 ;
        RECT 53.650 183.845 54.870 184.015 ;
        RECT 55.040 183.935 55.500 184.225 ;
        RECT 55.805 184.105 56.365 184.275 ;
        RECT 56.810 184.135 57.885 184.305 ;
        RECT 58.055 184.405 58.735 184.735 ;
        RECT 58.950 184.405 59.200 184.735 ;
        RECT 59.370 184.445 59.620 184.905 ;
        RECT 56.195 183.965 56.365 184.105 ;
        RECT 55.040 183.925 56.005 183.935 ;
        RECT 54.700 183.755 54.870 183.845 ;
        RECT 55.330 183.765 56.005 183.925 ;
        RECT 52.740 183.565 53.480 183.595 ;
        RECT 52.740 183.265 53.655 183.565 ;
        RECT 53.330 183.090 53.655 183.265 ;
        RECT 52.360 182.535 52.615 183.065 ;
        RECT 52.785 182.355 53.090 182.815 ;
        RECT 53.335 182.735 53.655 183.090 ;
        RECT 53.825 183.305 54.365 183.675 ;
        RECT 54.700 183.585 55.105 183.755 ;
        RECT 53.825 182.905 54.065 183.305 ;
        RECT 54.545 183.135 54.765 183.415 ;
        RECT 54.235 182.965 54.765 183.135 ;
        RECT 54.235 182.735 54.405 182.965 ;
        RECT 54.935 182.805 55.105 183.585 ;
        RECT 55.275 182.975 55.625 183.595 ;
        RECT 55.795 182.975 56.005 183.765 ;
        RECT 56.195 183.795 57.695 183.965 ;
        RECT 56.195 183.105 56.365 183.795 ;
        RECT 58.055 183.625 58.225 184.405 ;
        RECT 59.030 184.275 59.200 184.405 ;
        RECT 56.535 183.455 58.225 183.625 ;
        RECT 58.395 183.845 58.860 184.235 ;
        RECT 59.030 184.105 59.425 184.275 ;
        RECT 56.535 183.275 56.705 183.455 ;
        RECT 53.335 182.565 54.405 182.735 ;
        RECT 54.575 182.355 54.765 182.795 ;
        RECT 54.935 182.525 55.885 182.805 ;
        RECT 56.195 182.715 56.455 183.105 ;
        RECT 56.875 183.035 57.665 183.285 ;
        RECT 56.105 182.545 56.455 182.715 ;
        RECT 56.665 182.355 56.995 182.815 ;
        RECT 57.870 182.745 58.040 183.455 ;
        RECT 58.395 183.255 58.565 183.845 ;
        RECT 58.210 183.035 58.565 183.255 ;
        RECT 58.735 183.035 59.085 183.655 ;
        RECT 59.255 182.745 59.425 184.105 ;
        RECT 59.790 183.935 60.115 184.720 ;
        RECT 59.595 182.885 60.055 183.935 ;
        RECT 57.870 182.575 58.725 182.745 ;
        RECT 58.930 182.575 59.425 182.745 ;
        RECT 59.595 182.355 59.925 182.715 ;
        RECT 60.285 182.615 60.455 184.735 ;
        RECT 60.625 184.405 60.955 184.905 ;
        RECT 61.125 184.235 61.380 184.735 ;
        RECT 60.630 184.065 61.380 184.235 ;
        RECT 60.630 183.075 60.860 184.065 ;
        RECT 61.030 183.245 61.380 183.895 ;
        RECT 61.555 183.740 61.845 184.905 ;
        RECT 62.070 184.035 62.355 184.905 ;
        RECT 62.525 184.275 62.785 184.735 ;
        RECT 62.960 184.445 63.215 184.905 ;
        RECT 63.385 184.275 63.645 184.735 ;
        RECT 62.525 184.105 63.645 184.275 ;
        RECT 63.815 184.105 64.125 184.905 ;
        RECT 62.525 183.855 62.785 184.105 ;
        RECT 64.295 183.935 64.605 184.735 ;
        RECT 62.030 183.685 62.785 183.855 ;
        RECT 63.575 183.765 64.605 183.935 ;
        RECT 64.815 183.765 65.045 184.905 ;
        RECT 62.030 183.175 62.435 183.685 ;
        RECT 63.575 183.515 63.745 183.765 ;
        RECT 62.605 183.345 63.745 183.515 ;
        RECT 60.630 182.905 61.380 183.075 ;
        RECT 60.625 182.355 60.955 182.735 ;
        RECT 61.125 182.615 61.380 182.905 ;
        RECT 61.555 182.355 61.845 183.080 ;
        RECT 62.030 183.005 63.680 183.175 ;
        RECT 63.915 183.025 64.265 183.595 ;
        RECT 62.075 182.355 62.355 182.835 ;
        RECT 62.525 182.615 62.785 183.005 ;
        RECT 62.960 182.355 63.215 182.835 ;
        RECT 63.385 182.615 63.680 183.005 ;
        RECT 64.435 182.855 64.605 183.765 ;
        RECT 65.215 183.755 65.545 184.735 ;
        RECT 65.715 183.765 65.925 184.905 ;
        RECT 66.160 183.755 66.420 184.905 ;
        RECT 66.595 183.830 66.850 184.735 ;
        RECT 67.020 184.145 67.350 184.905 ;
        RECT 67.565 183.975 67.735 184.735 ;
        RECT 64.795 183.345 65.125 183.595 ;
        RECT 63.860 182.355 64.135 182.835 ;
        RECT 64.305 182.525 64.605 182.855 ;
        RECT 64.815 182.355 65.045 183.175 ;
        RECT 65.295 183.155 65.545 183.755 ;
        RECT 65.215 182.525 65.545 183.155 ;
        RECT 65.715 182.355 65.925 183.175 ;
        RECT 66.160 182.355 66.420 183.195 ;
        RECT 66.595 183.100 66.765 183.830 ;
        RECT 67.020 183.805 67.735 183.975 ;
        RECT 67.020 183.595 67.190 183.805 ;
        RECT 68.000 183.755 68.260 184.905 ;
        RECT 68.435 183.830 68.690 184.735 ;
        RECT 68.860 184.145 69.190 184.905 ;
        RECT 69.405 183.975 69.575 184.735 ;
        RECT 66.935 183.265 67.190 183.595 ;
        RECT 66.595 182.525 66.850 183.100 ;
        RECT 67.020 183.075 67.190 183.265 ;
        RECT 67.470 183.255 67.825 183.625 ;
        RECT 67.020 182.905 67.735 183.075 ;
        RECT 67.020 182.355 67.350 182.735 ;
        RECT 67.565 182.525 67.735 182.905 ;
        RECT 68.000 182.355 68.260 183.195 ;
        RECT 68.435 183.100 68.605 183.830 ;
        RECT 68.860 183.805 69.575 183.975 ;
        RECT 68.860 183.595 69.030 183.805 ;
        RECT 68.775 183.265 69.030 183.595 ;
        RECT 68.435 182.525 68.690 183.100 ;
        RECT 68.860 183.075 69.030 183.265 ;
        RECT 69.310 183.255 69.665 183.625 ;
        RECT 69.835 183.095 70.095 184.720 ;
        RECT 71.845 184.455 72.175 184.905 ;
        RECT 70.275 184.065 72.885 184.275 ;
        RECT 70.275 183.265 70.495 184.065 ;
        RECT 70.735 183.265 71.035 183.885 ;
        RECT 71.205 183.265 71.535 183.885 ;
        RECT 71.705 183.265 72.025 183.885 ;
        RECT 72.195 183.265 72.545 183.885 ;
        RECT 72.715 183.095 72.885 184.065 ;
        RECT 73.525 183.845 73.855 184.905 ;
        RECT 74.035 183.595 74.205 184.520 ;
        RECT 74.375 184.315 74.705 184.715 ;
        RECT 74.875 184.545 75.205 184.905 ;
        RECT 75.405 184.315 76.105 184.735 ;
        RECT 74.375 184.085 76.105 184.315 ;
        RECT 74.375 183.865 74.705 184.085 ;
        RECT 74.900 183.595 75.225 183.885 ;
        RECT 73.515 183.265 73.825 183.595 ;
        RECT 74.035 183.265 74.410 183.595 ;
        RECT 74.730 183.265 75.225 183.595 ;
        RECT 75.400 183.345 75.730 183.885 ;
        RECT 75.900 183.115 76.105 184.085 ;
        RECT 76.275 184.145 76.790 184.555 ;
        RECT 77.025 184.145 77.195 184.905 ;
        RECT 77.365 184.565 79.395 184.735 ;
        RECT 76.275 183.335 76.615 184.145 ;
        RECT 77.365 183.900 77.535 184.565 ;
        RECT 77.930 184.225 79.055 184.395 ;
        RECT 76.785 183.710 77.535 183.900 ;
        RECT 77.705 183.885 78.715 184.055 ;
        RECT 76.275 183.165 77.505 183.335 ;
        RECT 68.860 182.905 69.575 183.075 ;
        RECT 69.835 182.925 71.675 183.095 ;
        RECT 68.860 182.355 69.190 182.735 ;
        RECT 69.405 182.525 69.575 182.905 ;
        RECT 70.105 182.355 70.435 182.750 ;
        RECT 70.605 182.570 70.805 182.925 ;
        RECT 70.975 182.355 71.305 182.755 ;
        RECT 71.475 182.580 71.675 182.925 ;
        RECT 71.845 182.355 72.175 183.095 ;
        RECT 72.410 182.925 72.885 183.095 ;
        RECT 72.410 182.675 72.580 182.925 ;
        RECT 73.525 182.885 74.885 183.095 ;
        RECT 73.525 182.525 73.855 182.885 ;
        RECT 74.025 182.355 74.355 182.715 ;
        RECT 74.555 182.525 74.885 182.885 ;
        RECT 75.395 182.525 76.105 183.115 ;
        RECT 76.550 182.560 76.795 183.165 ;
        RECT 77.015 182.355 77.525 182.890 ;
        RECT 77.705 182.525 77.895 183.885 ;
        RECT 78.065 182.865 78.340 183.685 ;
        RECT 78.545 183.085 78.715 183.885 ;
        RECT 78.885 183.095 79.055 184.225 ;
        RECT 79.225 183.595 79.395 184.565 ;
        RECT 79.565 183.765 79.735 184.905 ;
        RECT 79.905 183.765 80.240 184.735 ;
        RECT 79.225 183.265 79.420 183.595 ;
        RECT 79.645 183.265 79.900 183.595 ;
        RECT 79.645 183.095 79.815 183.265 ;
        RECT 80.070 183.095 80.240 183.765 ;
        RECT 80.415 184.145 80.930 184.555 ;
        RECT 81.165 184.145 81.335 184.905 ;
        RECT 81.505 184.565 83.535 184.735 ;
        RECT 80.415 183.335 80.755 184.145 ;
        RECT 81.505 183.900 81.675 184.565 ;
        RECT 82.070 184.225 83.195 184.395 ;
        RECT 80.925 183.710 81.675 183.900 ;
        RECT 81.845 183.885 82.855 184.055 ;
        RECT 80.415 183.165 81.645 183.335 ;
        RECT 78.885 182.925 79.815 183.095 ;
        RECT 78.885 182.890 79.060 182.925 ;
        RECT 78.065 182.695 78.345 182.865 ;
        RECT 78.065 182.525 78.340 182.695 ;
        RECT 78.530 182.525 79.060 182.890 ;
        RECT 79.485 182.355 79.815 182.755 ;
        RECT 79.985 182.525 80.240 183.095 ;
        RECT 80.690 182.560 80.935 183.165 ;
        RECT 81.155 182.355 81.665 182.890 ;
        RECT 81.845 182.525 82.035 183.885 ;
        RECT 82.205 183.545 82.480 183.685 ;
        RECT 82.205 183.375 82.485 183.545 ;
        RECT 82.205 182.525 82.480 183.375 ;
        RECT 82.685 183.085 82.855 183.885 ;
        RECT 83.025 183.095 83.195 184.225 ;
        RECT 83.365 183.595 83.535 184.565 ;
        RECT 83.705 183.765 83.875 184.905 ;
        RECT 84.045 183.765 84.380 184.735 ;
        RECT 84.645 183.975 84.815 184.735 ;
        RECT 84.995 184.145 85.325 184.905 ;
        RECT 84.645 183.805 85.310 183.975 ;
        RECT 85.495 183.830 85.765 184.735 ;
        RECT 83.365 183.265 83.560 183.595 ;
        RECT 83.785 183.265 84.040 183.595 ;
        RECT 83.785 183.095 83.955 183.265 ;
        RECT 84.210 183.095 84.380 183.765 ;
        RECT 85.140 183.660 85.310 183.805 ;
        RECT 84.575 183.255 84.905 183.625 ;
        RECT 85.140 183.330 85.425 183.660 ;
        RECT 83.025 182.925 83.955 183.095 ;
        RECT 83.025 182.890 83.200 182.925 ;
        RECT 82.670 182.525 83.200 182.890 ;
        RECT 83.625 182.355 83.955 182.755 ;
        RECT 84.125 182.525 84.380 183.095 ;
        RECT 85.140 183.075 85.310 183.330 ;
        RECT 84.645 182.905 85.310 183.075 ;
        RECT 85.595 183.030 85.765 183.830 ;
        RECT 84.645 182.525 84.815 182.905 ;
        RECT 84.995 182.355 85.325 182.735 ;
        RECT 85.505 182.525 85.765 183.030 ;
        RECT 85.935 183.830 86.205 184.735 ;
        RECT 86.375 184.145 86.705 184.905 ;
        RECT 86.885 183.975 87.055 184.735 ;
        RECT 85.935 183.030 86.105 183.830 ;
        RECT 86.390 183.805 87.055 183.975 ;
        RECT 86.390 183.660 86.560 183.805 ;
        RECT 87.315 183.740 87.605 184.905 ;
        RECT 87.775 183.765 88.115 184.735 ;
        RECT 88.285 183.765 88.455 184.905 ;
        RECT 88.725 184.105 88.975 184.905 ;
        RECT 89.620 183.935 89.950 184.735 ;
        RECT 90.250 184.105 90.580 184.905 ;
        RECT 90.750 183.935 91.080 184.735 ;
        RECT 88.645 183.765 91.080 183.935 ;
        RECT 91.660 183.935 91.990 184.735 ;
        RECT 92.160 184.105 92.490 184.905 ;
        RECT 92.790 183.935 93.120 184.735 ;
        RECT 93.765 184.105 94.015 184.905 ;
        RECT 91.660 183.765 94.095 183.935 ;
        RECT 94.285 183.765 94.455 184.905 ;
        RECT 94.625 183.765 94.965 184.735 ;
        RECT 95.250 184.275 95.535 184.735 ;
        RECT 95.705 184.445 95.975 184.905 ;
        RECT 95.250 184.055 96.205 184.275 ;
        RECT 86.275 183.330 86.560 183.660 ;
        RECT 86.390 183.075 86.560 183.330 ;
        RECT 86.795 183.255 87.125 183.625 ;
        RECT 87.775 183.155 87.950 183.765 ;
        RECT 88.645 183.515 88.815 183.765 ;
        RECT 88.120 183.345 88.815 183.515 ;
        RECT 88.990 183.345 89.410 183.545 ;
        RECT 89.580 183.345 89.910 183.545 ;
        RECT 90.080 183.345 90.410 183.545 ;
        RECT 85.935 182.525 86.195 183.030 ;
        RECT 86.390 182.905 87.055 183.075 ;
        RECT 86.375 182.355 86.705 182.735 ;
        RECT 86.885 182.525 87.055 182.905 ;
        RECT 87.315 182.355 87.605 183.080 ;
        RECT 87.775 182.525 88.115 183.155 ;
        RECT 88.285 182.355 88.535 183.155 ;
        RECT 88.725 183.005 89.950 183.175 ;
        RECT 88.725 182.525 89.055 183.005 ;
        RECT 89.225 182.355 89.450 182.815 ;
        RECT 89.620 182.525 89.950 183.005 ;
        RECT 90.580 183.135 90.750 183.765 ;
        RECT 90.935 183.345 91.285 183.595 ;
        RECT 91.455 183.345 91.805 183.595 ;
        RECT 91.990 183.135 92.160 183.765 ;
        RECT 92.330 183.345 92.660 183.545 ;
        RECT 92.830 183.345 93.160 183.545 ;
        RECT 93.330 183.345 93.750 183.545 ;
        RECT 93.925 183.515 94.095 183.765 ;
        RECT 93.925 183.345 94.620 183.515 ;
        RECT 90.580 182.525 91.080 183.135 ;
        RECT 91.660 182.525 92.160 183.135 ;
        RECT 92.790 183.005 94.015 183.175 ;
        RECT 94.790 183.155 94.965 183.765 ;
        RECT 95.135 183.325 95.825 183.885 ;
        RECT 95.995 183.155 96.205 184.055 ;
        RECT 92.790 182.525 93.120 183.005 ;
        RECT 93.290 182.355 93.515 182.815 ;
        RECT 93.685 182.525 94.015 183.005 ;
        RECT 94.205 182.355 94.455 183.155 ;
        RECT 94.625 182.525 94.965 183.155 ;
        RECT 95.250 182.985 96.205 183.155 ;
        RECT 96.375 183.885 96.775 184.735 ;
        RECT 96.965 184.275 97.245 184.735 ;
        RECT 97.765 184.445 98.090 184.905 ;
        RECT 96.965 184.055 98.090 184.275 ;
        RECT 96.375 183.325 97.470 183.885 ;
        RECT 97.640 183.595 98.090 184.055 ;
        RECT 98.260 183.765 98.645 184.735 ;
        RECT 95.250 182.525 95.535 182.985 ;
        RECT 95.705 182.355 95.975 182.815 ;
        RECT 96.375 182.525 96.775 183.325 ;
        RECT 97.640 183.265 98.195 183.595 ;
        RECT 97.640 183.155 98.090 183.265 ;
        RECT 96.965 182.985 98.090 183.155 ;
        RECT 98.365 183.095 98.645 183.765 ;
        RECT 96.965 182.525 97.245 182.985 ;
        RECT 97.765 182.355 98.090 182.815 ;
        RECT 98.260 182.525 98.645 183.095 ;
        RECT 99.275 183.830 99.545 184.735 ;
        RECT 99.715 184.145 100.045 184.905 ;
        RECT 100.225 183.975 100.395 184.735 ;
        RECT 99.275 183.030 99.445 183.830 ;
        RECT 99.730 183.805 100.395 183.975 ;
        RECT 100.655 184.145 101.170 184.555 ;
        RECT 101.405 184.145 101.575 184.905 ;
        RECT 101.745 184.565 103.775 184.735 ;
        RECT 99.730 183.660 99.900 183.805 ;
        RECT 99.615 183.330 99.900 183.660 ;
        RECT 99.730 183.075 99.900 183.330 ;
        RECT 100.135 183.255 100.465 183.625 ;
        RECT 100.655 183.335 100.995 184.145 ;
        RECT 101.745 183.900 101.915 184.565 ;
        RECT 102.310 184.225 103.435 184.395 ;
        RECT 101.165 183.710 101.915 183.900 ;
        RECT 102.085 183.885 103.095 184.055 ;
        RECT 100.655 183.165 101.885 183.335 ;
        RECT 99.275 182.525 99.535 183.030 ;
        RECT 99.730 182.905 100.395 183.075 ;
        RECT 99.715 182.355 100.045 182.735 ;
        RECT 100.225 182.525 100.395 182.905 ;
        RECT 100.930 182.560 101.175 183.165 ;
        RECT 101.395 182.355 101.905 182.890 ;
        RECT 102.085 182.525 102.275 183.885 ;
        RECT 102.445 183.205 102.720 183.685 ;
        RECT 102.445 183.035 102.725 183.205 ;
        RECT 102.925 183.085 103.095 183.885 ;
        RECT 103.265 183.095 103.435 184.225 ;
        RECT 103.605 183.595 103.775 184.565 ;
        RECT 103.945 183.765 104.115 184.905 ;
        RECT 104.285 183.765 104.620 184.735 ;
        RECT 103.605 183.265 103.800 183.595 ;
        RECT 104.025 183.265 104.280 183.595 ;
        RECT 104.025 183.095 104.195 183.265 ;
        RECT 104.450 183.095 104.620 183.765 ;
        RECT 102.445 182.525 102.720 183.035 ;
        RECT 103.265 182.925 104.195 183.095 ;
        RECT 103.265 182.890 103.440 182.925 ;
        RECT 102.910 182.525 103.440 182.890 ;
        RECT 103.865 182.355 104.195 182.755 ;
        RECT 104.365 182.525 104.620 183.095 ;
        RECT 104.795 183.765 105.135 184.735 ;
        RECT 105.305 183.765 105.475 184.905 ;
        RECT 105.745 184.105 105.995 184.905 ;
        RECT 106.640 183.935 106.970 184.735 ;
        RECT 107.270 184.105 107.600 184.905 ;
        RECT 107.770 183.935 108.100 184.735 ;
        RECT 105.665 183.765 108.100 183.935 ;
        RECT 108.475 183.765 108.815 184.735 ;
        RECT 108.985 183.765 109.155 184.905 ;
        RECT 109.425 184.105 109.675 184.905 ;
        RECT 110.320 183.935 110.650 184.735 ;
        RECT 110.950 184.105 111.280 184.905 ;
        RECT 111.450 183.935 111.780 184.735 ;
        RECT 109.345 183.765 111.780 183.935 ;
        RECT 112.155 183.815 113.365 184.905 ;
        RECT 104.795 183.155 104.970 183.765 ;
        RECT 105.665 183.515 105.835 183.765 ;
        RECT 105.140 183.345 105.835 183.515 ;
        RECT 106.010 183.345 106.430 183.545 ;
        RECT 106.600 183.345 106.930 183.545 ;
        RECT 107.100 183.345 107.430 183.545 ;
        RECT 104.795 182.525 105.135 183.155 ;
        RECT 105.305 182.355 105.555 183.155 ;
        RECT 105.745 183.005 106.970 183.175 ;
        RECT 105.745 182.525 106.075 183.005 ;
        RECT 106.245 182.355 106.470 182.815 ;
        RECT 106.640 182.525 106.970 183.005 ;
        RECT 107.600 183.135 107.770 183.765 ;
        RECT 107.955 183.345 108.305 183.595 ;
        RECT 108.475 183.155 108.650 183.765 ;
        RECT 109.345 183.515 109.515 183.765 ;
        RECT 108.820 183.345 109.515 183.515 ;
        RECT 109.690 183.345 110.110 183.545 ;
        RECT 110.280 183.345 110.610 183.545 ;
        RECT 110.780 183.345 111.110 183.545 ;
        RECT 107.600 182.525 108.100 183.135 ;
        RECT 108.475 182.525 108.815 183.155 ;
        RECT 108.985 182.355 109.235 183.155 ;
        RECT 109.425 183.005 110.650 183.175 ;
        RECT 109.425 182.525 109.755 183.005 ;
        RECT 109.925 182.355 110.150 182.815 ;
        RECT 110.320 182.525 110.650 183.005 ;
        RECT 111.280 183.135 111.450 183.765 ;
        RECT 111.635 183.345 111.985 183.595 ;
        RECT 112.155 183.275 112.675 183.815 ;
        RECT 111.280 182.525 111.780 183.135 ;
        RECT 112.845 183.105 113.365 183.645 ;
        RECT 112.155 182.355 113.365 183.105 ;
        RECT 22.830 182.185 113.450 182.355 ;
        RECT 22.915 181.435 24.125 182.185 ;
        RECT 25.305 181.635 25.475 182.015 ;
        RECT 25.655 181.805 25.985 182.185 ;
        RECT 25.305 181.465 25.970 181.635 ;
        RECT 26.165 181.510 26.425 182.015 ;
        RECT 22.915 180.895 23.435 181.435 ;
        RECT 23.605 180.725 24.125 181.265 ;
        RECT 25.235 180.915 25.565 181.285 ;
        RECT 25.800 181.210 25.970 181.465 ;
        RECT 25.800 180.880 26.085 181.210 ;
        RECT 25.800 180.735 25.970 180.880 ;
        RECT 22.915 179.635 24.125 180.725 ;
        RECT 25.305 180.565 25.970 180.735 ;
        RECT 26.255 180.710 26.425 181.510 ;
        RECT 25.305 179.805 25.475 180.565 ;
        RECT 25.655 179.635 25.985 180.395 ;
        RECT 26.155 179.805 26.425 180.710 ;
        RECT 26.600 181.445 26.855 182.015 ;
        RECT 27.025 181.785 27.355 182.185 ;
        RECT 27.780 181.650 28.310 182.015 ;
        RECT 28.500 181.845 28.775 182.015 ;
        RECT 28.495 181.675 28.775 181.845 ;
        RECT 27.780 181.615 27.955 181.650 ;
        RECT 27.025 181.445 27.955 181.615 ;
        RECT 26.600 180.775 26.770 181.445 ;
        RECT 27.025 181.275 27.195 181.445 ;
        RECT 26.940 180.945 27.195 181.275 ;
        RECT 27.420 180.945 27.615 181.275 ;
        RECT 26.600 179.805 26.935 180.775 ;
        RECT 27.105 179.635 27.275 180.775 ;
        RECT 27.445 179.975 27.615 180.945 ;
        RECT 27.785 180.315 27.955 181.445 ;
        RECT 28.125 180.655 28.295 181.455 ;
        RECT 28.500 180.855 28.775 181.675 ;
        RECT 28.945 180.655 29.135 182.015 ;
        RECT 29.315 181.650 29.825 182.185 ;
        RECT 30.045 181.375 30.290 181.980 ;
        RECT 30.825 181.635 30.995 181.925 ;
        RECT 31.165 181.805 31.495 182.185 ;
        RECT 30.825 181.465 31.490 181.635 ;
        RECT 29.335 181.205 30.565 181.375 ;
        RECT 28.125 180.485 29.135 180.655 ;
        RECT 29.305 180.640 30.055 180.830 ;
        RECT 27.785 180.145 28.910 180.315 ;
        RECT 29.305 179.975 29.475 180.640 ;
        RECT 30.225 180.395 30.565 181.205 ;
        RECT 30.740 180.645 31.090 181.295 ;
        RECT 31.260 180.475 31.490 181.465 ;
        RECT 27.445 179.805 29.475 179.975 ;
        RECT 29.645 179.635 29.815 180.395 ;
        RECT 30.050 179.985 30.565 180.395 ;
        RECT 30.825 180.305 31.490 180.475 ;
        RECT 30.825 179.805 30.995 180.305 ;
        RECT 31.165 179.635 31.495 180.135 ;
        RECT 31.665 179.805 31.890 181.925 ;
        RECT 32.105 181.805 32.435 182.185 ;
        RECT 32.605 181.635 32.775 181.965 ;
        RECT 33.075 181.805 34.090 182.005 ;
        RECT 32.080 181.445 32.775 181.635 ;
        RECT 32.080 180.475 32.250 181.445 ;
        RECT 32.420 180.645 32.830 181.265 ;
        RECT 33.000 180.695 33.220 181.565 ;
        RECT 33.400 181.255 33.750 181.625 ;
        RECT 33.920 181.075 34.090 181.805 ;
        RECT 34.260 181.745 34.670 182.185 ;
        RECT 34.960 181.545 35.210 181.975 ;
        RECT 35.410 181.725 35.730 182.185 ;
        RECT 36.290 181.795 37.140 181.965 ;
        RECT 34.260 181.205 34.670 181.535 ;
        RECT 34.960 181.205 35.380 181.545 ;
        RECT 33.670 181.035 34.090 181.075 ;
        RECT 33.670 180.865 35.020 181.035 ;
        RECT 32.080 180.305 32.775 180.475 ;
        RECT 33.000 180.315 33.500 180.695 ;
        RECT 32.105 179.635 32.435 180.135 ;
        RECT 32.605 179.805 32.775 180.305 ;
        RECT 33.670 180.020 33.840 180.865 ;
        RECT 34.770 180.705 35.020 180.865 ;
        RECT 34.010 180.435 34.260 180.695 ;
        RECT 35.190 180.435 35.380 181.205 ;
        RECT 34.010 180.185 35.380 180.435 ;
        RECT 35.550 181.375 36.800 181.545 ;
        RECT 35.550 180.615 35.720 181.375 ;
        RECT 36.470 181.255 36.800 181.375 ;
        RECT 35.890 180.795 36.070 181.205 ;
        RECT 36.970 181.035 37.140 181.795 ;
        RECT 37.340 181.705 38.000 182.185 ;
        RECT 38.180 181.590 38.500 181.920 ;
        RECT 37.330 181.265 37.990 181.535 ;
        RECT 37.330 181.205 37.660 181.265 ;
        RECT 37.810 181.035 38.140 181.095 ;
        RECT 36.240 180.865 38.140 181.035 ;
        RECT 35.550 180.305 36.070 180.615 ;
        RECT 36.240 180.355 36.410 180.865 ;
        RECT 38.310 180.695 38.500 181.590 ;
        RECT 36.580 180.525 38.500 180.695 ;
        RECT 38.180 180.505 38.500 180.525 ;
        RECT 38.700 181.275 38.950 181.925 ;
        RECT 39.130 181.725 39.415 182.185 ;
        RECT 39.595 181.475 39.850 182.005 ;
        RECT 38.700 180.945 39.500 181.275 ;
        RECT 36.240 180.185 37.450 180.355 ;
        RECT 33.010 179.850 33.840 180.020 ;
        RECT 34.080 179.635 34.460 180.015 ;
        RECT 34.640 179.895 34.810 180.185 ;
        RECT 36.240 180.105 36.410 180.185 ;
        RECT 34.980 179.635 35.310 180.015 ;
        RECT 35.780 179.855 36.410 180.105 ;
        RECT 36.590 179.635 37.010 180.015 ;
        RECT 37.210 179.895 37.450 180.185 ;
        RECT 37.680 179.635 38.010 180.325 ;
        RECT 38.180 179.895 38.350 180.505 ;
        RECT 38.700 180.355 38.950 180.945 ;
        RECT 39.670 180.615 39.850 181.475 ;
        RECT 41.520 181.405 42.020 182.015 ;
        RECT 41.315 180.945 41.665 181.195 ;
        RECT 41.850 180.775 42.020 181.405 ;
        RECT 42.650 181.535 42.980 182.015 ;
        RECT 43.150 181.725 43.375 182.185 ;
        RECT 43.545 181.535 43.875 182.015 ;
        RECT 42.650 181.365 43.875 181.535 ;
        RECT 44.065 181.385 44.315 182.185 ;
        RECT 44.485 181.385 44.825 182.015 ;
        RECT 45.110 181.555 45.395 182.015 ;
        RECT 45.565 181.725 45.835 182.185 ;
        RECT 45.110 181.385 46.065 181.555 ;
        RECT 42.190 180.995 42.520 181.195 ;
        RECT 42.690 180.995 43.020 181.195 ;
        RECT 43.190 180.995 43.610 181.195 ;
        RECT 43.785 181.025 44.480 181.195 ;
        RECT 43.785 180.775 43.955 181.025 ;
        RECT 44.650 180.825 44.825 181.385 ;
        RECT 44.595 180.775 44.825 180.825 ;
        RECT 38.620 179.845 38.950 180.355 ;
        RECT 39.130 179.635 39.415 180.435 ;
        RECT 39.595 180.145 39.850 180.615 ;
        RECT 41.520 180.605 43.955 180.775 ;
        RECT 39.595 179.975 39.935 180.145 ;
        RECT 39.595 179.945 39.850 179.975 ;
        RECT 41.520 179.805 41.850 180.605 ;
        RECT 42.020 179.635 42.350 180.435 ;
        RECT 42.650 179.805 42.980 180.605 ;
        RECT 43.625 179.635 43.875 180.435 ;
        RECT 44.145 179.635 44.315 180.775 ;
        RECT 44.485 179.805 44.825 180.775 ;
        RECT 44.995 180.655 45.685 181.215 ;
        RECT 45.855 180.485 46.065 181.385 ;
        RECT 45.110 180.265 46.065 180.485 ;
        RECT 46.235 181.215 46.635 182.015 ;
        RECT 46.825 181.555 47.105 182.015 ;
        RECT 47.625 181.725 47.950 182.185 ;
        RECT 46.825 181.385 47.950 181.555 ;
        RECT 48.120 181.445 48.505 182.015 ;
        RECT 48.675 181.460 48.965 182.185 ;
        RECT 50.145 181.635 50.315 182.015 ;
        RECT 50.495 181.805 50.825 182.185 ;
        RECT 50.145 181.465 50.810 181.635 ;
        RECT 51.005 181.510 51.265 182.015 ;
        RECT 47.500 181.275 47.950 181.385 ;
        RECT 46.235 180.655 47.330 181.215 ;
        RECT 47.500 180.945 48.055 181.275 ;
        RECT 45.110 179.805 45.395 180.265 ;
        RECT 45.565 179.635 45.835 180.095 ;
        RECT 46.235 179.805 46.635 180.655 ;
        RECT 47.500 180.485 47.950 180.945 ;
        RECT 48.225 180.775 48.505 181.445 ;
        RECT 50.075 180.915 50.405 181.285 ;
        RECT 50.640 181.210 50.810 181.465 ;
        RECT 50.640 180.880 50.925 181.210 ;
        RECT 46.825 180.265 47.950 180.485 ;
        RECT 46.825 179.805 47.105 180.265 ;
        RECT 47.625 179.635 47.950 180.095 ;
        RECT 48.120 179.805 48.505 180.775 ;
        RECT 48.675 179.635 48.965 180.800 ;
        RECT 50.640 180.735 50.810 180.880 ;
        RECT 50.145 180.565 50.810 180.735 ;
        RECT 51.095 180.710 51.265 181.510 ;
        RECT 51.640 181.405 52.140 182.015 ;
        RECT 51.435 180.945 51.785 181.195 ;
        RECT 51.970 180.775 52.140 181.405 ;
        RECT 52.770 181.535 53.100 182.015 ;
        RECT 53.270 181.725 53.495 182.185 ;
        RECT 53.665 181.535 53.995 182.015 ;
        RECT 52.770 181.365 53.995 181.535 ;
        RECT 54.185 181.385 54.435 182.185 ;
        RECT 54.605 181.385 54.945 182.015 ;
        RECT 52.310 180.995 52.640 181.195 ;
        RECT 52.810 180.995 53.140 181.195 ;
        RECT 53.310 180.995 53.730 181.195 ;
        RECT 53.905 181.025 54.600 181.195 ;
        RECT 53.905 180.775 54.075 181.025 ;
        RECT 54.770 180.825 54.945 181.385 ;
        RECT 55.390 181.375 55.635 181.980 ;
        RECT 55.855 181.650 56.365 182.185 ;
        RECT 54.715 180.775 54.945 180.825 ;
        RECT 50.145 179.805 50.315 180.565 ;
        RECT 50.495 179.635 50.825 180.395 ;
        RECT 50.995 179.805 51.265 180.710 ;
        RECT 51.640 180.605 54.075 180.775 ;
        RECT 51.640 179.805 51.970 180.605 ;
        RECT 52.140 179.635 52.470 180.435 ;
        RECT 52.770 179.805 53.100 180.605 ;
        RECT 53.745 179.635 53.995 180.435 ;
        RECT 54.265 179.635 54.435 180.775 ;
        RECT 54.605 179.805 54.945 180.775 ;
        RECT 55.115 181.205 56.345 181.375 ;
        RECT 55.115 180.395 55.455 181.205 ;
        RECT 55.625 180.640 56.375 180.830 ;
        RECT 55.115 179.985 55.630 180.395 ;
        RECT 55.865 179.635 56.035 180.395 ;
        RECT 56.205 179.975 56.375 180.640 ;
        RECT 56.545 180.655 56.735 182.015 ;
        RECT 56.905 181.165 57.180 182.015 ;
        RECT 57.370 181.650 57.900 182.015 ;
        RECT 58.325 181.785 58.655 182.185 ;
        RECT 57.725 181.615 57.900 181.650 ;
        RECT 56.905 180.995 57.185 181.165 ;
        RECT 56.905 180.855 57.180 180.995 ;
        RECT 57.385 180.655 57.555 181.455 ;
        RECT 56.545 180.485 57.555 180.655 ;
        RECT 57.725 181.445 58.655 181.615 ;
        RECT 58.825 181.445 59.080 182.015 ;
        RECT 57.725 180.315 57.895 181.445 ;
        RECT 58.485 181.275 58.655 181.445 ;
        RECT 56.770 180.145 57.895 180.315 ;
        RECT 58.065 180.945 58.260 181.275 ;
        RECT 58.485 180.945 58.740 181.275 ;
        RECT 58.065 179.975 58.235 180.945 ;
        RECT 58.910 180.775 59.080 181.445 ;
        RECT 56.205 179.805 58.235 179.975 ;
        RECT 58.405 179.635 58.575 180.775 ;
        RECT 58.745 179.805 59.080 180.775 ;
        RECT 59.260 181.475 59.515 182.005 ;
        RECT 59.685 181.725 59.990 182.185 ;
        RECT 60.235 181.805 61.305 181.975 ;
        RECT 59.260 180.825 59.470 181.475 ;
        RECT 60.235 181.450 60.555 181.805 ;
        RECT 60.230 181.275 60.555 181.450 ;
        RECT 59.640 180.975 60.555 181.275 ;
        RECT 60.725 181.235 60.965 181.635 ;
        RECT 61.135 181.575 61.305 181.805 ;
        RECT 61.475 181.745 61.665 182.185 ;
        RECT 61.835 181.735 62.785 182.015 ;
        RECT 63.005 181.825 63.355 181.995 ;
        RECT 61.135 181.405 61.665 181.575 ;
        RECT 59.640 180.945 60.380 180.975 ;
        RECT 59.260 179.945 59.515 180.825 ;
        RECT 59.685 179.635 59.990 180.775 ;
        RECT 60.210 180.355 60.380 180.945 ;
        RECT 60.725 180.865 61.265 181.235 ;
        RECT 61.445 181.125 61.665 181.405 ;
        RECT 61.835 180.955 62.005 181.735 ;
        RECT 61.600 180.785 62.005 180.955 ;
        RECT 62.175 180.945 62.525 181.565 ;
        RECT 61.600 180.695 61.770 180.785 ;
        RECT 62.695 180.775 62.905 181.565 ;
        RECT 60.550 180.525 61.770 180.695 ;
        RECT 62.230 180.615 62.905 180.775 ;
        RECT 60.210 180.185 61.010 180.355 ;
        RECT 60.330 179.635 60.660 180.015 ;
        RECT 60.840 179.895 61.010 180.185 ;
        RECT 61.600 180.145 61.770 180.525 ;
        RECT 61.940 180.605 62.905 180.615 ;
        RECT 63.095 181.435 63.355 181.825 ;
        RECT 63.565 181.725 63.895 182.185 ;
        RECT 64.770 181.795 65.625 181.965 ;
        RECT 65.830 181.795 66.325 181.965 ;
        RECT 66.495 181.825 66.825 182.185 ;
        RECT 63.095 180.745 63.265 181.435 ;
        RECT 63.435 181.085 63.605 181.265 ;
        RECT 63.775 181.255 64.565 181.505 ;
        RECT 64.770 181.085 64.940 181.795 ;
        RECT 65.110 181.285 65.465 181.505 ;
        RECT 63.435 180.915 65.125 181.085 ;
        RECT 61.940 180.315 62.400 180.605 ;
        RECT 63.095 180.575 64.595 180.745 ;
        RECT 63.095 180.435 63.265 180.575 ;
        RECT 62.705 180.265 63.265 180.435 ;
        RECT 61.180 179.635 61.430 180.095 ;
        RECT 61.600 179.805 62.470 180.145 ;
        RECT 62.705 179.805 62.875 180.265 ;
        RECT 63.710 180.235 64.785 180.405 ;
        RECT 63.045 179.635 63.415 180.095 ;
        RECT 63.710 179.895 63.880 180.235 ;
        RECT 64.050 179.635 64.380 180.065 ;
        RECT 64.615 179.895 64.785 180.235 ;
        RECT 64.955 180.135 65.125 180.915 ;
        RECT 65.295 180.695 65.465 181.285 ;
        RECT 65.635 180.885 65.985 181.505 ;
        RECT 65.295 180.305 65.760 180.695 ;
        RECT 66.155 180.435 66.325 181.795 ;
        RECT 66.495 180.605 66.955 181.655 ;
        RECT 65.930 180.265 66.325 180.435 ;
        RECT 65.930 180.135 66.100 180.265 ;
        RECT 64.955 179.805 65.635 180.135 ;
        RECT 65.850 179.805 66.100 180.135 ;
        RECT 66.270 179.635 66.520 180.095 ;
        RECT 66.690 179.820 67.015 180.605 ;
        RECT 67.185 179.805 67.355 181.925 ;
        RECT 67.525 181.805 67.855 182.185 ;
        RECT 68.025 181.635 68.280 181.925 ;
        RECT 67.530 181.465 68.280 181.635 ;
        RECT 69.005 181.635 69.175 182.015 ;
        RECT 69.390 181.805 69.720 182.185 ;
        RECT 69.005 181.465 69.720 181.635 ;
        RECT 67.530 180.475 67.760 181.465 ;
        RECT 67.930 180.645 68.280 181.295 ;
        RECT 68.915 180.915 69.270 181.285 ;
        RECT 69.550 181.275 69.720 181.465 ;
        RECT 69.890 181.440 70.145 182.015 ;
        RECT 69.550 180.945 69.805 181.275 ;
        RECT 69.550 180.735 69.720 180.945 ;
        RECT 69.005 180.565 69.720 180.735 ;
        RECT 69.975 180.710 70.145 181.440 ;
        RECT 70.320 181.345 70.580 182.185 ;
        RECT 70.960 181.405 71.460 182.015 ;
        RECT 70.755 180.945 71.105 181.195 ;
        RECT 67.530 180.305 68.280 180.475 ;
        RECT 67.525 179.635 67.855 180.135 ;
        RECT 68.025 179.805 68.280 180.305 ;
        RECT 69.005 179.805 69.175 180.565 ;
        RECT 69.390 179.635 69.720 180.395 ;
        RECT 69.890 179.805 70.145 180.710 ;
        RECT 70.320 179.635 70.580 180.785 ;
        RECT 71.290 180.775 71.460 181.405 ;
        RECT 72.090 181.535 72.420 182.015 ;
        RECT 72.590 181.725 72.815 182.185 ;
        RECT 72.985 181.535 73.315 182.015 ;
        RECT 72.090 181.365 73.315 181.535 ;
        RECT 73.505 181.385 73.755 182.185 ;
        RECT 73.925 181.385 74.265 182.015 ;
        RECT 74.435 181.460 74.725 182.185 ;
        RECT 75.010 181.555 75.295 182.015 ;
        RECT 75.465 181.725 75.735 182.185 ;
        RECT 75.010 181.385 75.965 181.555 ;
        RECT 74.035 181.335 74.265 181.385 ;
        RECT 71.630 180.995 71.960 181.195 ;
        RECT 72.130 180.995 72.460 181.195 ;
        RECT 72.630 180.995 73.050 181.195 ;
        RECT 73.225 181.025 73.920 181.195 ;
        RECT 73.225 180.775 73.395 181.025 ;
        RECT 74.090 180.775 74.265 181.335 ;
        RECT 70.960 180.605 73.395 180.775 ;
        RECT 70.960 179.805 71.290 180.605 ;
        RECT 71.460 179.635 71.790 180.435 ;
        RECT 72.090 179.805 72.420 180.605 ;
        RECT 73.065 179.635 73.315 180.435 ;
        RECT 73.585 179.635 73.755 180.775 ;
        RECT 73.925 179.805 74.265 180.775 ;
        RECT 74.435 179.635 74.725 180.800 ;
        RECT 74.895 180.655 75.585 181.215 ;
        RECT 75.755 180.485 75.965 181.385 ;
        RECT 75.010 180.265 75.965 180.485 ;
        RECT 76.135 181.215 76.535 182.015 ;
        RECT 76.725 181.555 77.005 182.015 ;
        RECT 77.525 181.725 77.850 182.185 ;
        RECT 76.725 181.385 77.850 181.555 ;
        RECT 78.020 181.445 78.405 182.015 ;
        RECT 77.400 181.275 77.850 181.385 ;
        RECT 76.135 180.655 77.230 181.215 ;
        RECT 77.400 180.945 77.955 181.275 ;
        RECT 75.010 179.805 75.295 180.265 ;
        RECT 75.465 179.635 75.735 180.095 ;
        RECT 76.135 179.805 76.535 180.655 ;
        RECT 77.400 180.485 77.850 180.945 ;
        RECT 78.125 180.775 78.405 181.445 ;
        RECT 76.725 180.265 77.850 180.485 ;
        RECT 76.725 179.805 77.005 180.265 ;
        RECT 77.525 179.635 77.850 180.095 ;
        RECT 78.020 179.805 78.405 180.775 ;
        RECT 78.580 181.475 78.835 182.005 ;
        RECT 79.005 181.725 79.310 182.185 ;
        RECT 79.555 181.805 80.625 181.975 ;
        RECT 78.580 180.825 78.790 181.475 ;
        RECT 79.555 181.450 79.875 181.805 ;
        RECT 79.550 181.275 79.875 181.450 ;
        RECT 78.960 180.975 79.875 181.275 ;
        RECT 80.045 181.235 80.285 181.635 ;
        RECT 80.455 181.575 80.625 181.805 ;
        RECT 80.795 181.745 80.985 182.185 ;
        RECT 81.155 181.735 82.105 182.015 ;
        RECT 82.325 181.825 82.675 181.995 ;
        RECT 80.455 181.405 80.985 181.575 ;
        RECT 78.960 180.945 79.700 180.975 ;
        RECT 78.580 179.945 78.835 180.825 ;
        RECT 79.005 179.635 79.310 180.775 ;
        RECT 79.530 180.355 79.700 180.945 ;
        RECT 80.045 180.865 80.585 181.235 ;
        RECT 80.765 181.125 80.985 181.405 ;
        RECT 81.155 180.955 81.325 181.735 ;
        RECT 80.920 180.785 81.325 180.955 ;
        RECT 81.495 180.945 81.845 181.565 ;
        RECT 80.920 180.695 81.090 180.785 ;
        RECT 82.015 180.775 82.225 181.565 ;
        RECT 79.870 180.525 81.090 180.695 ;
        RECT 81.550 180.615 82.225 180.775 ;
        RECT 79.530 180.185 80.330 180.355 ;
        RECT 79.650 179.635 79.980 180.015 ;
        RECT 80.160 179.895 80.330 180.185 ;
        RECT 80.920 180.145 81.090 180.525 ;
        RECT 81.260 180.605 82.225 180.615 ;
        RECT 82.415 181.435 82.675 181.825 ;
        RECT 82.885 181.725 83.215 182.185 ;
        RECT 84.090 181.795 84.945 181.965 ;
        RECT 85.150 181.795 85.645 181.965 ;
        RECT 85.815 181.825 86.145 182.185 ;
        RECT 82.415 180.745 82.585 181.435 ;
        RECT 82.755 181.085 82.925 181.265 ;
        RECT 83.095 181.255 83.885 181.505 ;
        RECT 84.090 181.085 84.260 181.795 ;
        RECT 84.430 181.285 84.785 181.505 ;
        RECT 82.755 180.915 84.445 181.085 ;
        RECT 81.260 180.315 81.720 180.605 ;
        RECT 82.415 180.575 83.915 180.745 ;
        RECT 82.415 180.435 82.585 180.575 ;
        RECT 82.025 180.265 82.585 180.435 ;
        RECT 80.500 179.635 80.750 180.095 ;
        RECT 80.920 179.805 81.790 180.145 ;
        RECT 82.025 179.805 82.195 180.265 ;
        RECT 83.030 180.235 84.105 180.405 ;
        RECT 82.365 179.635 82.735 180.095 ;
        RECT 83.030 179.895 83.200 180.235 ;
        RECT 83.370 179.635 83.700 180.065 ;
        RECT 83.935 179.895 84.105 180.235 ;
        RECT 84.275 180.135 84.445 180.915 ;
        RECT 84.615 180.695 84.785 181.285 ;
        RECT 84.955 180.885 85.305 181.505 ;
        RECT 84.615 180.305 85.080 180.695 ;
        RECT 85.475 180.435 85.645 181.795 ;
        RECT 85.815 180.605 86.275 181.655 ;
        RECT 85.250 180.265 85.645 180.435 ;
        RECT 85.250 180.135 85.420 180.265 ;
        RECT 84.275 179.805 84.955 180.135 ;
        RECT 85.170 179.805 85.420 180.135 ;
        RECT 85.590 179.635 85.840 180.095 ;
        RECT 86.010 179.820 86.335 180.605 ;
        RECT 86.505 179.805 86.675 181.925 ;
        RECT 86.845 181.805 87.175 182.185 ;
        RECT 87.345 181.635 87.600 181.925 ;
        RECT 86.850 181.465 87.600 181.635 ;
        RECT 86.850 180.475 87.080 181.465 ;
        RECT 88.440 181.405 88.940 182.015 ;
        RECT 87.250 180.645 87.600 181.295 ;
        RECT 88.235 180.945 88.585 181.195 ;
        RECT 88.770 180.775 88.940 181.405 ;
        RECT 89.570 181.535 89.900 182.015 ;
        RECT 90.070 181.725 90.295 182.185 ;
        RECT 90.465 181.535 90.795 182.015 ;
        RECT 89.570 181.365 90.795 181.535 ;
        RECT 90.985 181.385 91.235 182.185 ;
        RECT 91.405 181.385 91.745 182.015 ;
        RECT 92.490 181.555 92.775 182.015 ;
        RECT 92.945 181.725 93.215 182.185 ;
        RECT 92.490 181.385 93.445 181.555 ;
        RECT 89.110 180.995 89.440 181.195 ;
        RECT 89.610 180.995 89.940 181.195 ;
        RECT 90.110 180.995 90.530 181.195 ;
        RECT 90.705 181.025 91.400 181.195 ;
        RECT 90.705 180.775 90.875 181.025 ;
        RECT 91.570 180.825 91.745 181.385 ;
        RECT 91.515 180.775 91.745 180.825 ;
        RECT 88.440 180.605 90.875 180.775 ;
        RECT 86.850 180.305 87.600 180.475 ;
        RECT 86.845 179.635 87.175 180.135 ;
        RECT 87.345 179.805 87.600 180.305 ;
        RECT 88.440 179.805 88.770 180.605 ;
        RECT 88.940 179.635 89.270 180.435 ;
        RECT 89.570 179.805 89.900 180.605 ;
        RECT 90.545 179.635 90.795 180.435 ;
        RECT 91.065 179.635 91.235 180.775 ;
        RECT 91.405 179.805 91.745 180.775 ;
        RECT 92.375 180.655 93.065 181.215 ;
        RECT 93.235 180.485 93.445 181.385 ;
        RECT 92.490 180.265 93.445 180.485 ;
        RECT 93.615 181.215 94.015 182.015 ;
        RECT 94.205 181.555 94.485 182.015 ;
        RECT 95.005 181.725 95.330 182.185 ;
        RECT 94.205 181.385 95.330 181.555 ;
        RECT 95.500 181.445 95.885 182.015 ;
        RECT 94.880 181.275 95.330 181.385 ;
        RECT 93.615 180.655 94.710 181.215 ;
        RECT 94.880 180.945 95.435 181.275 ;
        RECT 92.490 179.805 92.775 180.265 ;
        RECT 92.945 179.635 93.215 180.095 ;
        RECT 93.615 179.805 94.015 180.655 ;
        RECT 94.880 180.485 95.330 180.945 ;
        RECT 95.605 180.775 95.885 181.445 ;
        RECT 96.330 181.375 96.575 181.980 ;
        RECT 96.795 181.650 97.305 182.185 ;
        RECT 94.205 180.265 95.330 180.485 ;
        RECT 94.205 179.805 94.485 180.265 ;
        RECT 95.005 179.635 95.330 180.095 ;
        RECT 95.500 179.805 95.885 180.775 ;
        RECT 96.055 181.205 97.285 181.375 ;
        RECT 96.055 180.395 96.395 181.205 ;
        RECT 96.565 180.640 97.315 180.830 ;
        RECT 96.055 179.985 96.570 180.395 ;
        RECT 96.805 179.635 96.975 180.395 ;
        RECT 97.145 179.975 97.315 180.640 ;
        RECT 97.485 180.655 97.675 182.015 ;
        RECT 97.845 181.845 98.120 182.015 ;
        RECT 97.845 181.675 98.125 181.845 ;
        RECT 97.845 180.855 98.120 181.675 ;
        RECT 98.310 181.650 98.840 182.015 ;
        RECT 99.265 181.785 99.595 182.185 ;
        RECT 98.665 181.615 98.840 181.650 ;
        RECT 98.325 180.655 98.495 181.455 ;
        RECT 97.485 180.485 98.495 180.655 ;
        RECT 98.665 181.445 99.595 181.615 ;
        RECT 99.765 181.445 100.020 182.015 ;
        RECT 100.195 181.460 100.485 182.185 ;
        RECT 98.665 180.315 98.835 181.445 ;
        RECT 99.425 181.275 99.595 181.445 ;
        RECT 97.710 180.145 98.835 180.315 ;
        RECT 99.005 180.945 99.200 181.275 ;
        RECT 99.425 180.945 99.680 181.275 ;
        RECT 99.005 179.975 99.175 180.945 ;
        RECT 99.850 180.775 100.020 181.445 ;
        RECT 100.655 181.445 101.040 182.015 ;
        RECT 101.210 181.725 101.535 182.185 ;
        RECT 102.055 181.555 102.335 182.015 ;
        RECT 97.145 179.805 99.175 179.975 ;
        RECT 99.345 179.635 99.515 180.775 ;
        RECT 99.685 179.805 100.020 180.775 ;
        RECT 100.195 179.635 100.485 180.800 ;
        RECT 100.655 180.775 100.935 181.445 ;
        RECT 101.210 181.385 102.335 181.555 ;
        RECT 101.210 181.275 101.660 181.385 ;
        RECT 101.105 180.945 101.660 181.275 ;
        RECT 102.525 181.215 102.925 182.015 ;
        RECT 103.325 181.725 103.595 182.185 ;
        RECT 103.765 181.555 104.050 182.015 ;
        RECT 100.655 179.805 101.040 180.775 ;
        RECT 101.210 180.485 101.660 180.945 ;
        RECT 101.830 180.655 102.925 181.215 ;
        RECT 101.210 180.265 102.335 180.485 ;
        RECT 101.210 179.635 101.535 180.095 ;
        RECT 102.055 179.805 102.335 180.265 ;
        RECT 102.525 179.805 102.925 180.655 ;
        RECT 103.095 181.385 104.050 181.555 ;
        RECT 104.335 181.385 104.675 182.015 ;
        RECT 104.845 181.385 105.095 182.185 ;
        RECT 105.285 181.535 105.615 182.015 ;
        RECT 105.785 181.725 106.010 182.185 ;
        RECT 106.180 181.535 106.510 182.015 ;
        RECT 103.095 180.485 103.305 181.385 ;
        RECT 104.335 181.335 104.565 181.385 ;
        RECT 105.285 181.365 106.510 181.535 ;
        RECT 107.140 181.405 107.640 182.015 ;
        RECT 108.130 181.555 108.415 182.015 ;
        RECT 108.585 181.725 108.855 182.185 ;
        RECT 103.475 180.655 104.165 181.215 ;
        RECT 104.335 180.775 104.510 181.335 ;
        RECT 104.680 181.025 105.375 181.195 ;
        RECT 105.205 180.775 105.375 181.025 ;
        RECT 105.550 180.995 105.970 181.195 ;
        RECT 106.140 180.995 106.470 181.195 ;
        RECT 106.640 180.995 106.970 181.195 ;
        RECT 107.140 180.775 107.310 181.405 ;
        RECT 108.130 181.385 109.085 181.555 ;
        RECT 107.495 180.945 107.845 181.195 ;
        RECT 103.095 180.265 104.050 180.485 ;
        RECT 103.325 179.635 103.595 180.095 ;
        RECT 103.765 179.805 104.050 180.265 ;
        RECT 104.335 179.805 104.675 180.775 ;
        RECT 104.845 179.635 105.015 180.775 ;
        RECT 105.205 180.605 107.640 180.775 ;
        RECT 108.015 180.655 108.705 181.215 ;
        RECT 105.285 179.635 105.535 180.435 ;
        RECT 106.180 179.805 106.510 180.605 ;
        RECT 106.810 179.635 107.140 180.435 ;
        RECT 107.310 179.805 107.640 180.605 ;
        RECT 108.875 180.485 109.085 181.385 ;
        RECT 108.130 180.265 109.085 180.485 ;
        RECT 109.255 181.215 109.655 182.015 ;
        RECT 109.845 181.555 110.125 182.015 ;
        RECT 110.645 181.725 110.970 182.185 ;
        RECT 109.845 181.385 110.970 181.555 ;
        RECT 111.140 181.445 111.525 182.015 ;
        RECT 110.520 181.275 110.970 181.385 ;
        RECT 109.255 180.655 110.350 181.215 ;
        RECT 110.520 180.945 111.075 181.275 ;
        RECT 108.130 179.805 108.415 180.265 ;
        RECT 108.585 179.635 108.855 180.095 ;
        RECT 109.255 179.805 109.655 180.655 ;
        RECT 110.520 180.485 110.970 180.945 ;
        RECT 111.245 180.775 111.525 181.445 ;
        RECT 112.155 181.435 113.365 182.185 ;
        RECT 109.845 180.265 110.970 180.485 ;
        RECT 109.845 179.805 110.125 180.265 ;
        RECT 110.645 179.635 110.970 180.095 ;
        RECT 111.140 179.805 111.525 180.775 ;
        RECT 112.155 180.725 112.675 181.265 ;
        RECT 112.845 180.895 113.365 181.435 ;
        RECT 112.155 179.635 113.365 180.725 ;
        RECT 22.830 179.465 113.450 179.635 ;
        RECT 22.915 178.375 24.125 179.465 ;
        RECT 24.410 178.835 24.695 179.295 ;
        RECT 24.865 179.005 25.135 179.465 ;
        RECT 24.410 178.615 25.365 178.835 ;
        RECT 22.915 177.665 23.435 178.205 ;
        RECT 23.605 177.835 24.125 178.375 ;
        RECT 24.295 177.885 24.985 178.445 ;
        RECT 25.155 177.715 25.365 178.615 ;
        RECT 22.915 176.915 24.125 177.665 ;
        RECT 24.410 177.545 25.365 177.715 ;
        RECT 25.535 178.445 25.935 179.295 ;
        RECT 26.125 178.835 26.405 179.295 ;
        RECT 26.925 179.005 27.250 179.465 ;
        RECT 26.125 178.615 27.250 178.835 ;
        RECT 25.535 177.885 26.630 178.445 ;
        RECT 26.800 178.155 27.250 178.615 ;
        RECT 27.420 178.325 27.805 179.295 ;
        RECT 28.180 178.495 28.510 179.295 ;
        RECT 28.680 178.665 29.010 179.465 ;
        RECT 29.310 178.495 29.640 179.295 ;
        RECT 30.285 178.665 30.535 179.465 ;
        RECT 28.180 178.325 30.615 178.495 ;
        RECT 30.805 178.325 30.975 179.465 ;
        RECT 31.145 178.325 31.485 179.295 ;
        RECT 24.410 177.085 24.695 177.545 ;
        RECT 24.865 176.915 25.135 177.375 ;
        RECT 25.535 177.085 25.935 177.885 ;
        RECT 26.800 177.825 27.355 178.155 ;
        RECT 26.800 177.715 27.250 177.825 ;
        RECT 26.125 177.545 27.250 177.715 ;
        RECT 27.525 177.655 27.805 178.325 ;
        RECT 27.975 177.905 28.325 178.155 ;
        RECT 28.510 177.695 28.680 178.325 ;
        RECT 28.850 177.905 29.180 178.105 ;
        RECT 29.350 177.905 29.680 178.105 ;
        RECT 29.850 177.905 30.270 178.105 ;
        RECT 30.445 178.075 30.615 178.325 ;
        RECT 30.445 177.905 31.140 178.075 ;
        RECT 26.125 177.085 26.405 177.545 ;
        RECT 26.925 176.915 27.250 177.375 ;
        RECT 27.420 177.085 27.805 177.655 ;
        RECT 28.180 177.085 28.680 177.695 ;
        RECT 29.310 177.565 30.535 177.735 ;
        RECT 31.310 177.715 31.485 178.325 ;
        RECT 29.310 177.085 29.640 177.565 ;
        RECT 29.810 176.915 30.035 177.375 ;
        RECT 30.205 177.085 30.535 177.565 ;
        RECT 30.725 176.915 30.975 177.715 ;
        RECT 31.145 177.085 31.485 177.715 ;
        RECT 31.660 178.325 31.995 179.295 ;
        RECT 32.165 178.325 32.335 179.465 ;
        RECT 32.505 179.125 34.535 179.295 ;
        RECT 31.660 177.655 31.830 178.325 ;
        RECT 32.505 178.155 32.675 179.125 ;
        RECT 32.000 177.825 32.255 178.155 ;
        RECT 32.480 177.825 32.675 178.155 ;
        RECT 32.845 178.785 33.970 178.955 ;
        RECT 32.085 177.655 32.255 177.825 ;
        RECT 32.845 177.655 33.015 178.785 ;
        RECT 31.660 177.085 31.915 177.655 ;
        RECT 32.085 177.485 33.015 177.655 ;
        RECT 33.185 178.445 34.195 178.615 ;
        RECT 33.185 177.645 33.355 178.445 ;
        RECT 33.560 177.765 33.835 178.245 ;
        RECT 33.555 177.595 33.835 177.765 ;
        RECT 32.840 177.450 33.015 177.485 ;
        RECT 32.085 176.915 32.415 177.315 ;
        RECT 32.840 177.085 33.370 177.450 ;
        RECT 33.560 177.085 33.835 177.595 ;
        RECT 34.005 177.085 34.195 178.445 ;
        RECT 34.365 178.460 34.535 179.125 ;
        RECT 34.705 178.705 34.875 179.465 ;
        RECT 35.110 178.705 35.625 179.115 ;
        RECT 34.365 178.270 35.115 178.460 ;
        RECT 35.285 177.895 35.625 178.705 ;
        RECT 35.795 178.300 36.085 179.465 ;
        RECT 36.830 178.835 37.115 179.295 ;
        RECT 37.285 179.005 37.555 179.465 ;
        RECT 36.830 178.615 37.785 178.835 ;
        RECT 34.395 177.725 35.625 177.895 ;
        RECT 36.715 177.885 37.405 178.445 ;
        RECT 34.375 176.915 34.885 177.450 ;
        RECT 35.105 177.120 35.350 177.725 ;
        RECT 37.575 177.715 37.785 178.615 ;
        RECT 35.795 176.915 36.085 177.640 ;
        RECT 36.830 177.545 37.785 177.715 ;
        RECT 37.955 178.445 38.355 179.295 ;
        RECT 38.545 178.835 38.825 179.295 ;
        RECT 39.345 179.005 39.670 179.465 ;
        RECT 38.545 178.615 39.670 178.835 ;
        RECT 37.955 177.885 39.050 178.445 ;
        RECT 39.220 178.155 39.670 178.615 ;
        RECT 39.840 178.325 40.225 179.295 ;
        RECT 36.830 177.085 37.115 177.545 ;
        RECT 37.285 176.915 37.555 177.375 ;
        RECT 37.955 177.085 38.355 177.885 ;
        RECT 39.220 177.825 39.775 178.155 ;
        RECT 39.220 177.715 39.670 177.825 ;
        RECT 38.545 177.545 39.670 177.715 ;
        RECT 39.945 177.655 40.225 178.325 ;
        RECT 40.395 178.705 40.910 179.115 ;
        RECT 41.145 178.705 41.315 179.465 ;
        RECT 41.485 179.125 43.515 179.295 ;
        RECT 40.395 177.895 40.735 178.705 ;
        RECT 41.485 178.460 41.655 179.125 ;
        RECT 42.050 178.785 43.175 178.955 ;
        RECT 40.905 178.270 41.655 178.460 ;
        RECT 41.825 178.445 42.835 178.615 ;
        RECT 40.395 177.725 41.625 177.895 ;
        RECT 38.545 177.085 38.825 177.545 ;
        RECT 39.345 176.915 39.670 177.375 ;
        RECT 39.840 177.085 40.225 177.655 ;
        RECT 40.670 177.120 40.915 177.725 ;
        RECT 41.135 176.915 41.645 177.450 ;
        RECT 41.825 177.085 42.015 178.445 ;
        RECT 42.185 177.765 42.460 178.245 ;
        RECT 42.185 177.595 42.465 177.765 ;
        RECT 42.665 177.645 42.835 178.445 ;
        RECT 43.005 177.655 43.175 178.785 ;
        RECT 43.345 178.155 43.515 179.125 ;
        RECT 43.685 178.325 43.855 179.465 ;
        RECT 44.025 178.325 44.360 179.295 ;
        RECT 43.345 177.825 43.540 178.155 ;
        RECT 43.765 177.825 44.020 178.155 ;
        RECT 43.765 177.655 43.935 177.825 ;
        RECT 44.190 177.655 44.360 178.325 ;
        RECT 42.185 177.085 42.460 177.595 ;
        RECT 43.005 177.485 43.935 177.655 ;
        RECT 43.005 177.450 43.180 177.485 ;
        RECT 42.650 177.085 43.180 177.450 ;
        RECT 43.605 176.915 43.935 177.315 ;
        RECT 44.105 177.085 44.360 177.655 ;
        RECT 44.540 178.275 44.795 179.155 ;
        RECT 44.965 178.325 45.270 179.465 ;
        RECT 45.610 179.085 45.940 179.465 ;
        RECT 46.120 178.915 46.290 179.205 ;
        RECT 46.460 179.005 46.710 179.465 ;
        RECT 45.490 178.745 46.290 178.915 ;
        RECT 46.880 178.955 47.750 179.295 ;
        RECT 44.540 177.625 44.750 178.275 ;
        RECT 45.490 178.155 45.660 178.745 ;
        RECT 46.880 178.575 47.050 178.955 ;
        RECT 47.985 178.835 48.155 179.295 ;
        RECT 48.325 179.005 48.695 179.465 ;
        RECT 48.990 178.865 49.160 179.205 ;
        RECT 49.330 179.035 49.660 179.465 ;
        RECT 49.895 178.865 50.065 179.205 ;
        RECT 45.830 178.405 47.050 178.575 ;
        RECT 47.220 178.495 47.680 178.785 ;
        RECT 47.985 178.665 48.545 178.835 ;
        RECT 48.990 178.695 50.065 178.865 ;
        RECT 50.235 178.965 50.915 179.295 ;
        RECT 51.130 178.965 51.380 179.295 ;
        RECT 51.550 179.005 51.800 179.465 ;
        RECT 48.375 178.525 48.545 178.665 ;
        RECT 47.220 178.485 48.185 178.495 ;
        RECT 46.880 178.315 47.050 178.405 ;
        RECT 47.510 178.325 48.185 178.485 ;
        RECT 44.920 178.125 45.660 178.155 ;
        RECT 44.920 177.825 45.835 178.125 ;
        RECT 45.510 177.650 45.835 177.825 ;
        RECT 44.540 177.095 44.795 177.625 ;
        RECT 44.965 176.915 45.270 177.375 ;
        RECT 45.515 177.295 45.835 177.650 ;
        RECT 46.005 177.865 46.545 178.235 ;
        RECT 46.880 178.145 47.285 178.315 ;
        RECT 46.005 177.465 46.245 177.865 ;
        RECT 46.725 177.695 46.945 177.975 ;
        RECT 46.415 177.525 46.945 177.695 ;
        RECT 46.415 177.295 46.585 177.525 ;
        RECT 47.115 177.365 47.285 178.145 ;
        RECT 47.455 177.535 47.805 178.155 ;
        RECT 47.975 177.535 48.185 178.325 ;
        RECT 48.375 178.355 49.875 178.525 ;
        RECT 48.375 177.665 48.545 178.355 ;
        RECT 50.235 178.185 50.405 178.965 ;
        RECT 51.210 178.835 51.380 178.965 ;
        RECT 48.715 178.015 50.405 178.185 ;
        RECT 50.575 178.405 51.040 178.795 ;
        RECT 51.210 178.665 51.605 178.835 ;
        RECT 48.715 177.835 48.885 178.015 ;
        RECT 45.515 177.125 46.585 177.295 ;
        RECT 46.755 176.915 46.945 177.355 ;
        RECT 47.115 177.085 48.065 177.365 ;
        RECT 48.375 177.275 48.635 177.665 ;
        RECT 49.055 177.595 49.845 177.845 ;
        RECT 48.285 177.105 48.635 177.275 ;
        RECT 48.845 176.915 49.175 177.375 ;
        RECT 50.050 177.305 50.220 178.015 ;
        RECT 50.575 177.815 50.745 178.405 ;
        RECT 50.390 177.595 50.745 177.815 ;
        RECT 50.915 177.595 51.265 178.215 ;
        RECT 51.435 177.305 51.605 178.665 ;
        RECT 51.970 178.495 52.295 179.280 ;
        RECT 51.775 177.445 52.235 178.495 ;
        RECT 50.050 177.135 50.905 177.305 ;
        RECT 51.110 177.135 51.605 177.305 ;
        RECT 51.775 176.915 52.105 177.275 ;
        RECT 52.465 177.175 52.635 179.295 ;
        RECT 52.805 178.965 53.135 179.465 ;
        RECT 53.305 178.795 53.560 179.295 ;
        RECT 52.810 178.625 53.560 178.795 ;
        RECT 53.850 178.835 54.135 179.295 ;
        RECT 54.305 179.005 54.575 179.465 ;
        RECT 52.810 177.635 53.040 178.625 ;
        RECT 53.850 178.615 54.805 178.835 ;
        RECT 53.210 177.805 53.560 178.455 ;
        RECT 53.735 177.885 54.425 178.445 ;
        RECT 54.595 177.715 54.805 178.615 ;
        RECT 52.810 177.465 53.560 177.635 ;
        RECT 52.805 176.915 53.135 177.295 ;
        RECT 53.305 177.175 53.560 177.465 ;
        RECT 53.850 177.545 54.805 177.715 ;
        RECT 54.975 178.445 55.375 179.295 ;
        RECT 55.565 178.835 55.845 179.295 ;
        RECT 56.365 179.005 56.690 179.465 ;
        RECT 55.565 178.615 56.690 178.835 ;
        RECT 54.975 177.885 56.070 178.445 ;
        RECT 56.240 178.155 56.690 178.615 ;
        RECT 56.860 178.325 57.245 179.295 ;
        RECT 53.850 177.085 54.135 177.545 ;
        RECT 54.305 176.915 54.575 177.375 ;
        RECT 54.975 177.085 55.375 177.885 ;
        RECT 56.240 177.825 56.795 178.155 ;
        RECT 56.240 177.715 56.690 177.825 ;
        RECT 55.565 177.545 56.690 177.715 ;
        RECT 56.965 177.655 57.245 178.325 ;
        RECT 57.415 178.705 57.930 179.115 ;
        RECT 58.165 178.705 58.335 179.465 ;
        RECT 58.505 179.125 60.535 179.295 ;
        RECT 57.415 177.895 57.755 178.705 ;
        RECT 58.505 178.460 58.675 179.125 ;
        RECT 59.070 178.785 60.195 178.955 ;
        RECT 57.925 178.270 58.675 178.460 ;
        RECT 58.845 178.445 59.855 178.615 ;
        RECT 57.415 177.725 58.645 177.895 ;
        RECT 55.565 177.085 55.845 177.545 ;
        RECT 56.365 176.915 56.690 177.375 ;
        RECT 56.860 177.085 57.245 177.655 ;
        RECT 57.690 177.120 57.935 177.725 ;
        RECT 58.155 176.915 58.665 177.450 ;
        RECT 58.845 177.085 59.035 178.445 ;
        RECT 59.205 177.425 59.480 178.245 ;
        RECT 59.685 177.645 59.855 178.445 ;
        RECT 60.025 177.655 60.195 178.785 ;
        RECT 60.365 178.155 60.535 179.125 ;
        RECT 60.705 178.325 60.875 179.465 ;
        RECT 61.045 178.325 61.380 179.295 ;
        RECT 60.365 177.825 60.560 178.155 ;
        RECT 60.785 177.825 61.040 178.155 ;
        RECT 60.785 177.655 60.955 177.825 ;
        RECT 61.210 177.655 61.380 178.325 ;
        RECT 61.555 178.300 61.845 179.465 ;
        RECT 62.075 178.325 62.285 179.465 ;
        RECT 62.455 178.315 62.785 179.295 ;
        RECT 62.955 178.325 63.185 179.465 ;
        RECT 63.945 178.535 64.115 179.295 ;
        RECT 64.295 178.705 64.625 179.465 ;
        RECT 63.945 178.365 64.610 178.535 ;
        RECT 64.795 178.390 65.065 179.295 ;
        RECT 60.025 177.485 60.955 177.655 ;
        RECT 60.025 177.450 60.200 177.485 ;
        RECT 59.205 177.255 59.485 177.425 ;
        RECT 59.205 177.085 59.480 177.255 ;
        RECT 59.670 177.085 60.200 177.450 ;
        RECT 60.625 176.915 60.955 177.315 ;
        RECT 61.125 177.085 61.380 177.655 ;
        RECT 61.555 176.915 61.845 177.640 ;
        RECT 62.075 176.915 62.285 177.735 ;
        RECT 62.455 177.715 62.705 178.315 ;
        RECT 64.440 178.220 64.610 178.365 ;
        RECT 62.875 177.905 63.205 178.155 ;
        RECT 63.875 177.815 64.205 178.185 ;
        RECT 64.440 177.890 64.725 178.220 ;
        RECT 62.455 177.085 62.785 177.715 ;
        RECT 62.955 176.915 63.185 177.735 ;
        RECT 64.440 177.635 64.610 177.890 ;
        RECT 63.945 177.465 64.610 177.635 ;
        RECT 64.895 177.590 65.065 178.390 ;
        RECT 65.235 178.375 66.445 179.465 ;
        RECT 65.235 177.835 65.755 178.375 ;
        RECT 66.620 178.315 66.880 179.465 ;
        RECT 67.055 178.390 67.310 179.295 ;
        RECT 67.480 178.705 67.810 179.465 ;
        RECT 68.025 178.535 68.195 179.295 ;
        RECT 65.925 177.665 66.445 178.205 ;
        RECT 63.945 177.085 64.115 177.465 ;
        RECT 64.295 176.915 64.625 177.295 ;
        RECT 64.805 177.085 65.065 177.590 ;
        RECT 65.235 176.915 66.445 177.665 ;
        RECT 66.620 176.915 66.880 177.755 ;
        RECT 67.055 177.660 67.225 178.390 ;
        RECT 67.480 178.365 68.195 178.535 ;
        RECT 67.480 178.155 67.650 178.365 ;
        RECT 68.460 178.315 68.720 179.465 ;
        RECT 68.895 178.390 69.150 179.295 ;
        RECT 69.320 178.705 69.650 179.465 ;
        RECT 69.865 178.535 70.035 179.295 ;
        RECT 67.395 177.825 67.650 178.155 ;
        RECT 67.055 177.085 67.310 177.660 ;
        RECT 67.480 177.635 67.650 177.825 ;
        RECT 67.930 177.815 68.285 178.185 ;
        RECT 67.480 177.465 68.195 177.635 ;
        RECT 67.480 176.915 67.810 177.295 ;
        RECT 68.025 177.085 68.195 177.465 ;
        RECT 68.460 176.915 68.720 177.755 ;
        RECT 68.895 177.660 69.065 178.390 ;
        RECT 69.320 178.365 70.035 178.535 ;
        RECT 69.320 178.155 69.490 178.365 ;
        RECT 70.295 178.325 70.635 179.295 ;
        RECT 70.805 178.325 70.975 179.465 ;
        RECT 71.245 178.665 71.495 179.465 ;
        RECT 72.140 178.495 72.470 179.295 ;
        RECT 72.770 178.665 73.100 179.465 ;
        RECT 73.270 178.495 73.600 179.295 ;
        RECT 71.165 178.325 73.600 178.495 ;
        RECT 73.975 178.325 74.315 179.295 ;
        RECT 74.485 178.325 74.655 179.465 ;
        RECT 74.925 178.665 75.175 179.465 ;
        RECT 75.820 178.495 76.150 179.295 ;
        RECT 76.450 178.665 76.780 179.465 ;
        RECT 76.950 178.495 77.280 179.295 ;
        RECT 74.845 178.325 77.280 178.495 ;
        RECT 77.655 178.325 77.995 179.295 ;
        RECT 78.165 178.325 78.335 179.465 ;
        RECT 78.605 178.665 78.855 179.465 ;
        RECT 79.500 178.495 79.830 179.295 ;
        RECT 80.130 178.665 80.460 179.465 ;
        RECT 80.630 178.495 80.960 179.295 ;
        RECT 81.450 178.835 81.735 179.295 ;
        RECT 81.905 179.005 82.175 179.465 ;
        RECT 81.450 178.615 82.405 178.835 ;
        RECT 78.525 178.325 80.960 178.495 ;
        RECT 69.235 177.825 69.490 178.155 ;
        RECT 68.895 177.085 69.150 177.660 ;
        RECT 69.320 177.635 69.490 177.825 ;
        RECT 69.770 177.815 70.125 178.185 ;
        RECT 70.295 177.715 70.470 178.325 ;
        RECT 71.165 178.075 71.335 178.325 ;
        RECT 70.640 177.905 71.335 178.075 ;
        RECT 71.510 177.905 71.930 178.105 ;
        RECT 72.100 177.905 72.430 178.105 ;
        RECT 72.600 177.905 72.930 178.105 ;
        RECT 69.320 177.465 70.035 177.635 ;
        RECT 69.320 176.915 69.650 177.295 ;
        RECT 69.865 177.085 70.035 177.465 ;
        RECT 70.295 177.085 70.635 177.715 ;
        RECT 70.805 176.915 71.055 177.715 ;
        RECT 71.245 177.565 72.470 177.735 ;
        RECT 71.245 177.085 71.575 177.565 ;
        RECT 71.745 176.915 71.970 177.375 ;
        RECT 72.140 177.085 72.470 177.565 ;
        RECT 73.100 177.695 73.270 178.325 ;
        RECT 73.455 177.905 73.805 178.155 ;
        RECT 73.975 177.715 74.150 178.325 ;
        RECT 74.845 178.075 75.015 178.325 ;
        RECT 74.320 177.905 75.015 178.075 ;
        RECT 75.190 177.905 75.610 178.105 ;
        RECT 75.780 177.905 76.110 178.105 ;
        RECT 76.280 177.905 76.610 178.105 ;
        RECT 73.100 177.085 73.600 177.695 ;
        RECT 73.975 177.085 74.315 177.715 ;
        RECT 74.485 176.915 74.735 177.715 ;
        RECT 74.925 177.565 76.150 177.735 ;
        RECT 74.925 177.085 75.255 177.565 ;
        RECT 75.425 176.915 75.650 177.375 ;
        RECT 75.820 177.085 76.150 177.565 ;
        RECT 76.780 177.695 76.950 178.325 ;
        RECT 77.135 177.905 77.485 178.155 ;
        RECT 77.655 177.715 77.830 178.325 ;
        RECT 78.525 178.075 78.695 178.325 ;
        RECT 78.000 177.905 78.695 178.075 ;
        RECT 78.870 177.905 79.290 178.105 ;
        RECT 79.460 177.905 79.790 178.105 ;
        RECT 79.960 177.905 80.290 178.105 ;
        RECT 76.780 177.085 77.280 177.695 ;
        RECT 77.655 177.085 77.995 177.715 ;
        RECT 78.165 176.915 78.415 177.715 ;
        RECT 78.605 177.565 79.830 177.735 ;
        RECT 78.605 177.085 78.935 177.565 ;
        RECT 79.105 176.915 79.330 177.375 ;
        RECT 79.500 177.085 79.830 177.565 ;
        RECT 80.460 177.695 80.630 178.325 ;
        RECT 80.815 177.905 81.165 178.155 ;
        RECT 81.335 177.885 82.025 178.445 ;
        RECT 82.195 177.715 82.405 178.615 ;
        RECT 80.460 177.085 80.960 177.695 ;
        RECT 81.450 177.545 82.405 177.715 ;
        RECT 82.575 178.445 82.975 179.295 ;
        RECT 83.165 178.835 83.445 179.295 ;
        RECT 83.965 179.005 84.290 179.465 ;
        RECT 83.165 178.615 84.290 178.835 ;
        RECT 82.575 177.885 83.670 178.445 ;
        RECT 83.840 178.155 84.290 178.615 ;
        RECT 84.460 178.325 84.845 179.295 ;
        RECT 85.075 178.325 85.285 179.465 ;
        RECT 81.450 177.085 81.735 177.545 ;
        RECT 81.905 176.915 82.175 177.375 ;
        RECT 82.575 177.085 82.975 177.885 ;
        RECT 83.840 177.825 84.395 178.155 ;
        RECT 83.840 177.715 84.290 177.825 ;
        RECT 83.165 177.545 84.290 177.715 ;
        RECT 84.565 177.655 84.845 178.325 ;
        RECT 85.455 178.315 85.785 179.295 ;
        RECT 85.955 178.325 86.185 179.465 ;
        RECT 83.165 177.085 83.445 177.545 ;
        RECT 83.965 176.915 84.290 177.375 ;
        RECT 84.460 177.085 84.845 177.655 ;
        RECT 85.075 176.915 85.285 177.735 ;
        RECT 85.455 177.715 85.705 178.315 ;
        RECT 87.315 178.300 87.605 179.465 ;
        RECT 87.815 178.325 88.045 179.465 ;
        RECT 88.215 178.315 88.545 179.295 ;
        RECT 88.715 178.325 88.925 179.465 ;
        RECT 90.190 178.835 90.475 179.295 ;
        RECT 90.645 179.005 90.915 179.465 ;
        RECT 90.190 178.615 91.145 178.835 ;
        RECT 85.875 177.905 86.205 178.155 ;
        RECT 87.795 177.905 88.125 178.155 ;
        RECT 85.455 177.085 85.785 177.715 ;
        RECT 85.955 176.915 86.185 177.735 ;
        RECT 87.315 176.915 87.605 177.640 ;
        RECT 87.815 176.915 88.045 177.735 ;
        RECT 88.295 177.715 88.545 178.315 ;
        RECT 90.075 177.885 90.765 178.445 ;
        RECT 88.215 177.085 88.545 177.715 ;
        RECT 88.715 176.915 88.925 177.735 ;
        RECT 90.935 177.715 91.145 178.615 ;
        RECT 90.190 177.545 91.145 177.715 ;
        RECT 91.315 178.445 91.715 179.295 ;
        RECT 91.905 178.835 92.185 179.295 ;
        RECT 92.705 179.005 93.030 179.465 ;
        RECT 91.905 178.615 93.030 178.835 ;
        RECT 91.315 177.885 92.410 178.445 ;
        RECT 92.580 178.155 93.030 178.615 ;
        RECT 93.200 178.325 93.585 179.295 ;
        RECT 93.845 178.535 94.015 179.295 ;
        RECT 94.195 178.705 94.525 179.465 ;
        RECT 93.845 178.365 94.510 178.535 ;
        RECT 94.695 178.390 94.965 179.295 ;
        RECT 90.190 177.085 90.475 177.545 ;
        RECT 90.645 176.915 90.915 177.375 ;
        RECT 91.315 177.085 91.715 177.885 ;
        RECT 92.580 177.825 93.135 178.155 ;
        RECT 92.580 177.715 93.030 177.825 ;
        RECT 91.905 177.545 93.030 177.715 ;
        RECT 93.305 177.655 93.585 178.325 ;
        RECT 94.340 178.220 94.510 178.365 ;
        RECT 93.775 177.815 94.105 178.185 ;
        RECT 94.340 177.890 94.625 178.220 ;
        RECT 91.905 177.085 92.185 177.545 ;
        RECT 92.705 176.915 93.030 177.375 ;
        RECT 93.200 177.085 93.585 177.655 ;
        RECT 94.340 177.635 94.510 177.890 ;
        RECT 93.845 177.465 94.510 177.635 ;
        RECT 94.795 177.590 94.965 178.390 ;
        RECT 93.845 177.085 94.015 177.465 ;
        RECT 94.195 176.915 94.525 177.295 ;
        RECT 94.705 177.085 94.965 177.590 ;
        RECT 95.600 178.325 95.935 179.295 ;
        RECT 96.105 178.325 96.275 179.465 ;
        RECT 96.445 179.125 98.475 179.295 ;
        RECT 95.600 177.655 95.770 178.325 ;
        RECT 96.445 178.155 96.615 179.125 ;
        RECT 95.940 177.825 96.195 178.155 ;
        RECT 96.420 177.825 96.615 178.155 ;
        RECT 96.785 178.785 97.910 178.955 ;
        RECT 96.025 177.655 96.195 177.825 ;
        RECT 96.785 177.655 96.955 178.785 ;
        RECT 95.600 177.085 95.855 177.655 ;
        RECT 96.025 177.485 96.955 177.655 ;
        RECT 97.125 178.445 98.135 178.615 ;
        RECT 97.125 177.645 97.295 178.445 ;
        RECT 96.780 177.450 96.955 177.485 ;
        RECT 96.025 176.915 96.355 177.315 ;
        RECT 96.780 177.085 97.310 177.450 ;
        RECT 97.500 177.425 97.775 178.245 ;
        RECT 97.495 177.255 97.775 177.425 ;
        RECT 97.500 177.085 97.775 177.255 ;
        RECT 97.945 177.085 98.135 178.445 ;
        RECT 98.305 178.460 98.475 179.125 ;
        RECT 98.645 178.705 98.815 179.465 ;
        RECT 99.050 178.705 99.565 179.115 ;
        RECT 98.305 178.270 99.055 178.460 ;
        RECT 99.225 177.895 99.565 178.705 ;
        RECT 100.285 178.535 100.455 179.295 ;
        RECT 100.635 178.705 100.965 179.465 ;
        RECT 100.285 178.365 100.950 178.535 ;
        RECT 101.135 178.390 101.405 179.295 ;
        RECT 100.780 178.220 100.950 178.365 ;
        RECT 98.335 177.725 99.565 177.895 ;
        RECT 100.215 177.815 100.545 178.185 ;
        RECT 100.780 177.890 101.065 178.220 ;
        RECT 98.315 176.915 98.825 177.450 ;
        RECT 99.045 177.120 99.290 177.725 ;
        RECT 100.780 177.635 100.950 177.890 ;
        RECT 100.285 177.465 100.950 177.635 ;
        RECT 101.235 177.590 101.405 178.390 ;
        RECT 101.615 178.325 101.845 179.465 ;
        RECT 102.015 178.315 102.345 179.295 ;
        RECT 102.515 178.325 102.725 179.465 ;
        RECT 101.595 177.905 101.925 178.155 ;
        RECT 100.285 177.085 100.455 177.465 ;
        RECT 100.635 176.915 100.965 177.295 ;
        RECT 101.145 177.085 101.405 177.590 ;
        RECT 101.615 176.915 101.845 177.735 ;
        RECT 102.095 177.715 102.345 178.315 ;
        RECT 102.960 178.275 103.215 179.155 ;
        RECT 103.385 178.325 103.690 179.465 ;
        RECT 104.030 179.085 104.360 179.465 ;
        RECT 104.540 178.915 104.710 179.205 ;
        RECT 104.880 179.005 105.130 179.465 ;
        RECT 103.910 178.745 104.710 178.915 ;
        RECT 105.300 178.955 106.170 179.295 ;
        RECT 102.015 177.085 102.345 177.715 ;
        RECT 102.515 176.915 102.725 177.735 ;
        RECT 102.960 177.625 103.170 178.275 ;
        RECT 103.910 178.155 104.080 178.745 ;
        RECT 105.300 178.575 105.470 178.955 ;
        RECT 106.405 178.835 106.575 179.295 ;
        RECT 106.745 179.005 107.115 179.465 ;
        RECT 107.410 178.865 107.580 179.205 ;
        RECT 107.750 179.035 108.080 179.465 ;
        RECT 108.315 178.865 108.485 179.205 ;
        RECT 104.250 178.405 105.470 178.575 ;
        RECT 105.640 178.495 106.100 178.785 ;
        RECT 106.405 178.665 106.965 178.835 ;
        RECT 107.410 178.695 108.485 178.865 ;
        RECT 108.655 178.965 109.335 179.295 ;
        RECT 109.550 178.965 109.800 179.295 ;
        RECT 109.970 179.005 110.220 179.465 ;
        RECT 106.795 178.525 106.965 178.665 ;
        RECT 105.640 178.485 106.605 178.495 ;
        RECT 105.300 178.315 105.470 178.405 ;
        RECT 105.930 178.325 106.605 178.485 ;
        RECT 103.340 178.125 104.080 178.155 ;
        RECT 103.340 177.825 104.255 178.125 ;
        RECT 103.930 177.650 104.255 177.825 ;
        RECT 102.960 177.095 103.215 177.625 ;
        RECT 103.385 176.915 103.690 177.375 ;
        RECT 103.935 177.295 104.255 177.650 ;
        RECT 104.425 177.865 104.965 178.235 ;
        RECT 105.300 178.145 105.705 178.315 ;
        RECT 104.425 177.465 104.665 177.865 ;
        RECT 105.145 177.695 105.365 177.975 ;
        RECT 104.835 177.525 105.365 177.695 ;
        RECT 104.835 177.295 105.005 177.525 ;
        RECT 105.535 177.365 105.705 178.145 ;
        RECT 105.875 177.535 106.225 178.155 ;
        RECT 106.395 177.535 106.605 178.325 ;
        RECT 106.795 178.355 108.295 178.525 ;
        RECT 106.795 177.665 106.965 178.355 ;
        RECT 108.655 178.185 108.825 178.965 ;
        RECT 109.630 178.835 109.800 178.965 ;
        RECT 107.135 178.015 108.825 178.185 ;
        RECT 108.995 178.405 109.460 178.795 ;
        RECT 109.630 178.665 110.025 178.835 ;
        RECT 107.135 177.835 107.305 178.015 ;
        RECT 103.935 177.125 105.005 177.295 ;
        RECT 105.175 176.915 105.365 177.355 ;
        RECT 105.535 177.085 106.485 177.365 ;
        RECT 106.795 177.275 107.055 177.665 ;
        RECT 107.475 177.595 108.265 177.845 ;
        RECT 106.705 177.105 107.055 177.275 ;
        RECT 107.265 176.915 107.595 177.375 ;
        RECT 108.470 177.305 108.640 178.015 ;
        RECT 108.995 177.815 109.165 178.405 ;
        RECT 108.810 177.595 109.165 177.815 ;
        RECT 109.335 177.595 109.685 178.215 ;
        RECT 109.855 177.305 110.025 178.665 ;
        RECT 110.390 178.495 110.715 179.280 ;
        RECT 110.195 177.445 110.655 178.495 ;
        RECT 108.470 177.135 109.325 177.305 ;
        RECT 109.530 177.135 110.025 177.305 ;
        RECT 110.195 176.915 110.525 177.275 ;
        RECT 110.885 177.175 111.055 179.295 ;
        RECT 111.225 178.965 111.555 179.465 ;
        RECT 111.725 178.795 111.980 179.295 ;
        RECT 111.230 178.625 111.980 178.795 ;
        RECT 111.230 177.635 111.460 178.625 ;
        RECT 111.630 177.805 111.980 178.455 ;
        RECT 112.155 178.375 113.365 179.465 ;
        RECT 112.155 177.835 112.675 178.375 ;
        RECT 112.845 177.665 113.365 178.205 ;
        RECT 111.230 177.465 111.980 177.635 ;
        RECT 111.225 176.915 111.555 177.295 ;
        RECT 111.725 177.175 111.980 177.465 ;
        RECT 112.155 176.915 113.365 177.665 ;
        RECT 22.830 176.745 113.450 176.915 ;
        RECT 22.915 175.995 24.125 176.745 ;
        RECT 22.915 175.455 23.435 175.995 ;
        RECT 24.755 175.975 26.425 176.745 ;
        RECT 26.685 176.195 26.855 176.575 ;
        RECT 27.035 176.365 27.365 176.745 ;
        RECT 26.685 176.025 27.350 176.195 ;
        RECT 27.545 176.070 27.805 176.575 ;
        RECT 23.605 175.285 24.125 175.825 ;
        RECT 22.915 174.195 24.125 175.285 ;
        RECT 24.755 175.285 25.505 175.805 ;
        RECT 25.675 175.455 26.425 175.975 ;
        RECT 26.615 175.475 26.945 175.845 ;
        RECT 27.180 175.770 27.350 176.025 ;
        RECT 27.180 175.440 27.465 175.770 ;
        RECT 27.180 175.295 27.350 175.440 ;
        RECT 24.755 174.195 26.425 175.285 ;
        RECT 26.685 175.125 27.350 175.295 ;
        RECT 27.635 175.270 27.805 176.070 ;
        RECT 28.015 175.925 28.245 176.745 ;
        RECT 28.415 175.945 28.745 176.575 ;
        RECT 27.995 175.505 28.325 175.755 ;
        RECT 28.495 175.345 28.745 175.945 ;
        RECT 28.915 175.925 29.125 176.745 ;
        RECT 29.355 175.945 29.695 176.575 ;
        RECT 29.865 175.945 30.115 176.745 ;
        RECT 30.305 176.095 30.635 176.575 ;
        RECT 30.805 176.285 31.030 176.745 ;
        RECT 31.200 176.095 31.530 176.575 ;
        RECT 26.685 174.365 26.855 175.125 ;
        RECT 27.035 174.195 27.365 174.955 ;
        RECT 27.535 174.365 27.805 175.270 ;
        RECT 28.015 174.195 28.245 175.335 ;
        RECT 28.415 174.365 28.745 175.345 ;
        RECT 29.355 175.335 29.530 175.945 ;
        RECT 30.305 175.925 31.530 176.095 ;
        RECT 32.160 175.965 32.660 176.575 ;
        RECT 33.040 176.035 33.295 176.565 ;
        RECT 33.465 176.285 33.770 176.745 ;
        RECT 34.015 176.365 35.085 176.535 ;
        RECT 29.700 175.585 30.395 175.755 ;
        RECT 30.225 175.335 30.395 175.585 ;
        RECT 30.570 175.555 30.990 175.755 ;
        RECT 31.160 175.555 31.490 175.755 ;
        RECT 31.660 175.555 31.990 175.755 ;
        RECT 32.160 175.335 32.330 175.965 ;
        RECT 32.515 175.505 32.865 175.755 ;
        RECT 33.040 175.385 33.250 176.035 ;
        RECT 34.015 176.010 34.335 176.365 ;
        RECT 34.010 175.835 34.335 176.010 ;
        RECT 33.420 175.535 34.335 175.835 ;
        RECT 34.505 175.795 34.745 176.195 ;
        RECT 34.915 176.135 35.085 176.365 ;
        RECT 35.255 176.305 35.445 176.745 ;
        RECT 35.615 176.295 36.565 176.575 ;
        RECT 36.785 176.385 37.135 176.555 ;
        RECT 34.915 175.965 35.445 176.135 ;
        RECT 33.420 175.505 34.160 175.535 ;
        RECT 28.915 174.195 29.125 175.335 ;
        RECT 29.355 174.365 29.695 175.335 ;
        RECT 29.865 174.195 30.035 175.335 ;
        RECT 30.225 175.165 32.660 175.335 ;
        RECT 30.305 174.195 30.555 174.995 ;
        RECT 31.200 174.365 31.530 175.165 ;
        RECT 31.830 174.195 32.160 174.995 ;
        RECT 32.330 174.365 32.660 175.165 ;
        RECT 33.040 174.505 33.295 175.385 ;
        RECT 33.465 174.195 33.770 175.335 ;
        RECT 33.990 174.915 34.160 175.505 ;
        RECT 34.505 175.425 35.045 175.795 ;
        RECT 35.225 175.685 35.445 175.965 ;
        RECT 35.615 175.515 35.785 176.295 ;
        RECT 35.380 175.345 35.785 175.515 ;
        RECT 35.955 175.505 36.305 176.125 ;
        RECT 35.380 175.255 35.550 175.345 ;
        RECT 36.475 175.335 36.685 176.125 ;
        RECT 34.330 175.085 35.550 175.255 ;
        RECT 36.010 175.175 36.685 175.335 ;
        RECT 33.990 174.745 34.790 174.915 ;
        RECT 34.110 174.195 34.440 174.575 ;
        RECT 34.620 174.455 34.790 174.745 ;
        RECT 35.380 174.705 35.550 175.085 ;
        RECT 35.720 175.165 36.685 175.175 ;
        RECT 36.875 175.995 37.135 176.385 ;
        RECT 37.345 176.285 37.675 176.745 ;
        RECT 38.550 176.355 39.405 176.525 ;
        RECT 39.610 176.355 40.105 176.525 ;
        RECT 40.275 176.385 40.605 176.745 ;
        RECT 36.875 175.305 37.045 175.995 ;
        RECT 37.215 175.645 37.385 175.825 ;
        RECT 37.555 175.815 38.345 176.065 ;
        RECT 38.550 175.645 38.720 176.355 ;
        RECT 38.890 175.845 39.245 176.065 ;
        RECT 37.215 175.475 38.905 175.645 ;
        RECT 35.720 174.875 36.180 175.165 ;
        RECT 36.875 175.135 38.375 175.305 ;
        RECT 36.875 174.995 37.045 175.135 ;
        RECT 36.485 174.825 37.045 174.995 ;
        RECT 34.960 174.195 35.210 174.655 ;
        RECT 35.380 174.365 36.250 174.705 ;
        RECT 36.485 174.365 36.655 174.825 ;
        RECT 37.490 174.795 38.565 174.965 ;
        RECT 36.825 174.195 37.195 174.655 ;
        RECT 37.490 174.455 37.660 174.795 ;
        RECT 37.830 174.195 38.160 174.625 ;
        RECT 38.395 174.455 38.565 174.795 ;
        RECT 38.735 174.695 38.905 175.475 ;
        RECT 39.075 175.255 39.245 175.845 ;
        RECT 39.415 175.445 39.765 176.065 ;
        RECT 39.075 174.865 39.540 175.255 ;
        RECT 39.935 174.995 40.105 176.355 ;
        RECT 40.275 175.165 40.735 176.215 ;
        RECT 39.710 174.825 40.105 174.995 ;
        RECT 39.710 174.695 39.880 174.825 ;
        RECT 38.735 174.365 39.415 174.695 ;
        RECT 39.630 174.365 39.880 174.695 ;
        RECT 40.050 174.195 40.300 174.655 ;
        RECT 40.470 174.380 40.795 175.165 ;
        RECT 40.965 174.365 41.135 176.485 ;
        RECT 41.305 176.365 41.635 176.745 ;
        RECT 41.805 176.195 42.060 176.485 ;
        RECT 41.310 176.025 42.060 176.195 ;
        RECT 42.235 176.070 42.495 176.575 ;
        RECT 42.675 176.365 43.005 176.745 ;
        RECT 43.185 176.195 43.355 176.575 ;
        RECT 41.310 175.035 41.540 176.025 ;
        RECT 41.710 175.205 42.060 175.855 ;
        RECT 42.235 175.270 42.405 176.070 ;
        RECT 42.690 176.025 43.355 176.195 ;
        RECT 42.690 175.770 42.860 176.025 ;
        RECT 43.675 175.925 43.885 176.745 ;
        RECT 44.055 175.945 44.385 176.575 ;
        RECT 42.575 175.440 42.860 175.770 ;
        RECT 43.095 175.475 43.425 175.845 ;
        RECT 42.690 175.295 42.860 175.440 ;
        RECT 44.055 175.345 44.305 175.945 ;
        RECT 44.555 175.925 44.785 176.745 ;
        RECT 45.200 175.965 45.700 176.575 ;
        RECT 44.475 175.505 44.805 175.755 ;
        RECT 44.995 175.505 45.345 175.755 ;
        RECT 41.310 174.865 42.060 175.035 ;
        RECT 41.305 174.195 41.635 174.695 ;
        RECT 41.805 174.365 42.060 174.865 ;
        RECT 42.235 174.365 42.505 175.270 ;
        RECT 42.690 175.125 43.355 175.295 ;
        RECT 42.675 174.195 43.005 174.955 ;
        RECT 43.185 174.365 43.355 175.125 ;
        RECT 43.675 174.195 43.885 175.335 ;
        RECT 44.055 174.365 44.385 175.345 ;
        RECT 45.530 175.335 45.700 175.965 ;
        RECT 46.330 176.095 46.660 176.575 ;
        RECT 46.830 176.285 47.055 176.745 ;
        RECT 47.225 176.095 47.555 176.575 ;
        RECT 46.330 175.925 47.555 176.095 ;
        RECT 47.745 175.945 47.995 176.745 ;
        RECT 48.165 175.945 48.505 176.575 ;
        RECT 48.675 176.020 48.965 176.745 ;
        RECT 49.135 176.070 49.395 176.575 ;
        RECT 49.575 176.365 49.905 176.745 ;
        RECT 50.085 176.195 50.255 176.575 ;
        RECT 45.870 175.555 46.200 175.755 ;
        RECT 46.370 175.555 46.700 175.755 ;
        RECT 46.870 175.555 47.290 175.755 ;
        RECT 47.465 175.585 48.160 175.755 ;
        RECT 47.465 175.335 47.635 175.585 ;
        RECT 48.330 175.335 48.505 175.945 ;
        RECT 44.555 174.195 44.785 175.335 ;
        RECT 45.200 175.165 47.635 175.335 ;
        RECT 45.200 174.365 45.530 175.165 ;
        RECT 45.700 174.195 46.030 174.995 ;
        RECT 46.330 174.365 46.660 175.165 ;
        RECT 47.305 174.195 47.555 174.995 ;
        RECT 47.825 174.195 47.995 175.335 ;
        RECT 48.165 174.365 48.505 175.335 ;
        RECT 48.675 174.195 48.965 175.360 ;
        RECT 49.135 175.270 49.305 176.070 ;
        RECT 49.590 176.025 50.255 176.195 ;
        RECT 49.590 175.770 49.760 176.025 ;
        RECT 50.555 175.925 50.785 176.745 ;
        RECT 50.955 175.945 51.285 176.575 ;
        RECT 49.475 175.440 49.760 175.770 ;
        RECT 49.995 175.475 50.325 175.845 ;
        RECT 50.535 175.505 50.865 175.755 ;
        RECT 49.590 175.295 49.760 175.440 ;
        RECT 51.035 175.345 51.285 175.945 ;
        RECT 51.455 175.925 51.665 176.745 ;
        RECT 51.945 176.285 52.250 176.745 ;
        RECT 52.420 176.115 52.750 176.575 ;
        RECT 52.920 176.285 53.090 176.745 ;
        RECT 53.260 176.115 53.590 176.575 ;
        RECT 53.760 176.285 53.930 176.745 ;
        RECT 54.100 176.115 54.430 176.575 ;
        RECT 54.600 176.285 54.770 176.745 ;
        RECT 54.940 176.115 55.270 176.575 ;
        RECT 55.440 176.285 55.695 176.745 ;
        RECT 51.895 175.925 55.865 176.115 ;
        RECT 56.035 175.975 57.705 176.745 ;
        RECT 49.135 174.365 49.405 175.270 ;
        RECT 49.590 175.125 50.255 175.295 ;
        RECT 49.575 174.195 49.905 174.955 ;
        RECT 50.085 174.365 50.255 175.125 ;
        RECT 50.555 174.195 50.785 175.335 ;
        RECT 50.955 174.365 51.285 175.345 ;
        RECT 51.895 175.335 52.215 175.925 ;
        RECT 52.415 175.725 55.270 175.755 ;
        RECT 52.415 175.555 55.345 175.725 ;
        RECT 52.415 175.505 55.270 175.555 ;
        RECT 55.520 175.335 55.865 175.925 ;
        RECT 51.455 174.195 51.665 175.335 ;
        RECT 51.895 175.165 55.865 175.335 ;
        RECT 56.035 175.285 56.785 175.805 ;
        RECT 56.955 175.455 57.705 175.975 ;
        RECT 57.875 175.945 58.215 176.575 ;
        RECT 58.385 175.945 58.635 176.745 ;
        RECT 58.825 176.095 59.155 176.575 ;
        RECT 59.325 176.285 59.550 176.745 ;
        RECT 59.720 176.095 60.050 176.575 ;
        RECT 57.875 175.335 58.050 175.945 ;
        RECT 58.825 175.925 60.050 176.095 ;
        RECT 60.680 175.965 61.180 176.575 ;
        RECT 61.670 176.115 61.955 176.575 ;
        RECT 62.125 176.285 62.395 176.745 ;
        RECT 58.220 175.585 58.915 175.755 ;
        RECT 58.745 175.335 58.915 175.585 ;
        RECT 59.090 175.555 59.510 175.755 ;
        RECT 59.680 175.555 60.010 175.755 ;
        RECT 60.180 175.555 60.510 175.755 ;
        RECT 60.680 175.335 60.850 175.965 ;
        RECT 61.670 175.945 62.625 176.115 ;
        RECT 61.035 175.505 61.385 175.755 ;
        RECT 51.950 174.195 52.250 174.995 ;
        RECT 52.420 174.365 52.750 175.165 ;
        RECT 52.920 174.195 53.090 174.995 ;
        RECT 53.260 174.365 53.590 175.165 ;
        RECT 53.760 174.195 53.930 174.995 ;
        RECT 54.100 174.365 54.430 175.165 ;
        RECT 54.600 174.195 54.770 174.995 ;
        RECT 54.940 174.365 55.270 175.165 ;
        RECT 55.440 174.195 55.695 174.995 ;
        RECT 56.035 174.195 57.705 175.285 ;
        RECT 57.875 174.365 58.215 175.335 ;
        RECT 58.385 174.195 58.555 175.335 ;
        RECT 58.745 175.165 61.180 175.335 ;
        RECT 61.555 175.215 62.245 175.775 ;
        RECT 58.825 174.195 59.075 174.995 ;
        RECT 59.720 174.365 60.050 175.165 ;
        RECT 60.350 174.195 60.680 174.995 ;
        RECT 60.850 174.365 61.180 175.165 ;
        RECT 62.415 175.045 62.625 175.945 ;
        RECT 61.670 174.825 62.625 175.045 ;
        RECT 62.795 175.775 63.195 176.575 ;
        RECT 63.385 176.115 63.665 176.575 ;
        RECT 64.185 176.285 64.510 176.745 ;
        RECT 63.385 175.945 64.510 176.115 ;
        RECT 64.680 176.005 65.065 176.575 ;
        RECT 64.060 175.835 64.510 175.945 ;
        RECT 62.795 175.215 63.890 175.775 ;
        RECT 64.060 175.505 64.615 175.835 ;
        RECT 61.670 174.365 61.955 174.825 ;
        RECT 62.125 174.195 62.395 174.655 ;
        RECT 62.795 174.365 63.195 175.215 ;
        RECT 64.060 175.045 64.510 175.505 ;
        RECT 64.785 175.335 65.065 176.005 ;
        RECT 65.235 175.975 67.825 176.745 ;
        RECT 63.385 174.825 64.510 175.045 ;
        RECT 63.385 174.365 63.665 174.825 ;
        RECT 64.185 174.195 64.510 174.655 ;
        RECT 64.680 174.365 65.065 175.335 ;
        RECT 65.235 175.285 66.445 175.805 ;
        RECT 66.615 175.455 67.825 175.975 ;
        RECT 68.000 175.905 68.260 176.745 ;
        RECT 68.435 176.000 68.690 176.575 ;
        RECT 68.860 176.365 69.190 176.745 ;
        RECT 69.405 176.195 69.575 176.575 ;
        RECT 68.860 176.025 69.575 176.195 ;
        RECT 69.845 176.215 70.175 176.575 ;
        RECT 70.345 176.385 70.675 176.745 ;
        RECT 70.875 176.215 71.205 176.575 ;
        RECT 65.235 174.195 67.825 175.285 ;
        RECT 68.000 174.195 68.260 175.345 ;
        RECT 68.435 175.270 68.605 176.000 ;
        RECT 68.860 175.835 69.030 176.025 ;
        RECT 69.845 176.005 71.205 176.215 ;
        RECT 71.715 175.985 72.425 176.575 ;
        RECT 68.775 175.505 69.030 175.835 ;
        RECT 68.860 175.295 69.030 175.505 ;
        RECT 69.310 175.475 69.665 175.845 ;
        RECT 69.835 175.505 70.145 175.835 ;
        RECT 70.355 175.505 70.730 175.835 ;
        RECT 71.050 175.505 71.545 175.835 ;
        RECT 68.435 174.365 68.690 175.270 ;
        RECT 68.860 175.125 69.575 175.295 ;
        RECT 68.860 174.195 69.190 174.955 ;
        RECT 69.405 174.365 69.575 175.125 ;
        RECT 69.845 174.195 70.175 175.255 ;
        RECT 70.355 174.580 70.525 175.505 ;
        RECT 70.695 175.015 71.025 175.235 ;
        RECT 71.220 175.215 71.545 175.505 ;
        RECT 71.720 175.215 72.050 175.755 ;
        RECT 72.220 175.015 72.425 175.985 ;
        RECT 72.595 175.975 74.265 176.745 ;
        RECT 74.435 176.020 74.725 176.745 ;
        RECT 74.895 175.995 76.105 176.745 ;
        RECT 70.695 174.785 72.425 175.015 ;
        RECT 70.695 174.385 71.025 174.785 ;
        RECT 71.195 174.195 71.525 174.555 ;
        RECT 71.725 174.365 72.425 174.785 ;
        RECT 72.595 175.285 73.345 175.805 ;
        RECT 73.515 175.455 74.265 175.975 ;
        RECT 72.595 174.195 74.265 175.285 ;
        RECT 74.435 174.195 74.725 175.360 ;
        RECT 74.895 175.285 75.415 175.825 ;
        RECT 75.585 175.455 76.105 175.995 ;
        RECT 76.275 176.070 76.535 176.575 ;
        RECT 76.715 176.365 77.045 176.745 ;
        RECT 77.225 176.195 77.395 176.575 ;
        RECT 74.895 174.195 76.105 175.285 ;
        RECT 76.275 175.270 76.445 176.070 ;
        RECT 76.730 176.025 77.395 176.195 ;
        RECT 76.730 175.770 76.900 176.025 ;
        RECT 77.715 175.925 77.925 176.745 ;
        RECT 78.095 175.945 78.425 176.575 ;
        RECT 76.615 175.440 76.900 175.770 ;
        RECT 77.135 175.475 77.465 175.845 ;
        RECT 76.730 175.295 76.900 175.440 ;
        RECT 78.095 175.345 78.345 175.945 ;
        RECT 78.595 175.925 78.825 176.745 ;
        RECT 79.095 175.925 79.305 176.745 ;
        RECT 79.475 175.945 79.805 176.575 ;
        RECT 78.515 175.505 78.845 175.755 ;
        RECT 79.475 175.345 79.725 175.945 ;
        RECT 79.975 175.925 80.205 176.745 ;
        RECT 80.415 176.235 80.720 176.745 ;
        RECT 79.895 175.505 80.225 175.755 ;
        RECT 80.415 175.505 80.730 176.065 ;
        RECT 80.900 175.755 81.150 176.565 ;
        RECT 81.320 176.220 81.580 176.745 ;
        RECT 81.760 175.755 82.010 176.565 ;
        RECT 82.180 176.185 82.440 176.745 ;
        RECT 82.610 176.095 82.870 176.550 ;
        RECT 83.040 176.265 83.300 176.745 ;
        RECT 83.470 176.095 83.730 176.550 ;
        RECT 83.900 176.265 84.160 176.745 ;
        RECT 84.330 176.095 84.590 176.550 ;
        RECT 84.760 176.265 85.005 176.745 ;
        RECT 85.175 176.095 85.450 176.550 ;
        RECT 85.620 176.265 85.865 176.745 ;
        RECT 86.035 176.095 86.295 176.550 ;
        RECT 86.475 176.265 86.725 176.745 ;
        RECT 86.895 176.095 87.155 176.550 ;
        RECT 87.335 176.265 87.585 176.745 ;
        RECT 87.755 176.095 88.015 176.550 ;
        RECT 88.195 176.265 88.455 176.745 ;
        RECT 88.625 176.095 88.885 176.550 ;
        RECT 89.055 176.265 89.355 176.745 ;
        RECT 82.610 175.925 89.355 176.095 ;
        RECT 80.900 175.505 88.020 175.755 ;
        RECT 76.275 174.365 76.545 175.270 ;
        RECT 76.730 175.125 77.395 175.295 ;
        RECT 76.715 174.195 77.045 174.955 ;
        RECT 77.225 174.365 77.395 175.125 ;
        RECT 77.715 174.195 77.925 175.335 ;
        RECT 78.095 174.365 78.425 175.345 ;
        RECT 78.595 174.195 78.825 175.335 ;
        RECT 79.095 174.195 79.305 175.335 ;
        RECT 79.475 174.365 79.805 175.345 ;
        RECT 79.975 174.195 80.205 175.335 ;
        RECT 80.425 174.195 80.720 175.005 ;
        RECT 80.900 174.365 81.145 175.505 ;
        RECT 81.320 174.195 81.580 175.005 ;
        RECT 81.760 174.370 82.010 175.505 ;
        RECT 88.190 175.335 89.355 175.925 ;
        RECT 82.610 175.110 89.355 175.335 ;
        RECT 89.620 176.035 89.875 176.565 ;
        RECT 90.045 176.285 90.350 176.745 ;
        RECT 90.595 176.365 91.665 176.535 ;
        RECT 89.620 175.385 89.830 176.035 ;
        RECT 90.595 176.010 90.915 176.365 ;
        RECT 90.590 175.835 90.915 176.010 ;
        RECT 90.000 175.535 90.915 175.835 ;
        RECT 91.085 175.795 91.325 176.195 ;
        RECT 91.495 176.135 91.665 176.365 ;
        RECT 91.835 176.305 92.025 176.745 ;
        RECT 92.195 176.295 93.145 176.575 ;
        RECT 93.365 176.385 93.715 176.555 ;
        RECT 91.495 175.965 92.025 176.135 ;
        RECT 90.000 175.505 90.740 175.535 ;
        RECT 82.610 175.095 88.015 175.110 ;
        RECT 82.180 174.200 82.440 174.995 ;
        RECT 82.610 174.370 82.870 175.095 ;
        RECT 83.040 174.200 83.300 174.925 ;
        RECT 83.470 174.370 83.730 175.095 ;
        RECT 83.900 174.200 84.160 174.925 ;
        RECT 84.330 174.370 84.590 175.095 ;
        RECT 84.760 174.200 85.020 174.925 ;
        RECT 85.190 174.370 85.450 175.095 ;
        RECT 85.620 174.200 85.865 174.925 ;
        RECT 86.035 174.370 86.295 175.095 ;
        RECT 86.480 174.200 86.725 174.925 ;
        RECT 86.895 174.370 87.155 175.095 ;
        RECT 87.340 174.200 87.585 174.925 ;
        RECT 87.755 174.370 88.015 175.095 ;
        RECT 88.200 174.200 88.455 174.925 ;
        RECT 88.625 174.370 88.915 175.110 ;
        RECT 82.180 174.195 88.455 174.200 ;
        RECT 89.085 174.195 89.355 174.940 ;
        RECT 89.620 174.505 89.875 175.385 ;
        RECT 90.045 174.195 90.350 175.335 ;
        RECT 90.570 174.915 90.740 175.505 ;
        RECT 91.085 175.425 91.625 175.795 ;
        RECT 91.805 175.685 92.025 175.965 ;
        RECT 92.195 175.515 92.365 176.295 ;
        RECT 91.960 175.345 92.365 175.515 ;
        RECT 92.535 175.505 92.885 176.125 ;
        RECT 91.960 175.255 92.130 175.345 ;
        RECT 93.055 175.335 93.265 176.125 ;
        RECT 90.910 175.085 92.130 175.255 ;
        RECT 92.590 175.175 93.265 175.335 ;
        RECT 90.570 174.745 91.370 174.915 ;
        RECT 90.690 174.195 91.020 174.575 ;
        RECT 91.200 174.455 91.370 174.745 ;
        RECT 91.960 174.705 92.130 175.085 ;
        RECT 92.300 175.165 93.265 175.175 ;
        RECT 93.455 175.995 93.715 176.385 ;
        RECT 93.925 176.285 94.255 176.745 ;
        RECT 95.130 176.355 95.985 176.525 ;
        RECT 96.190 176.355 96.685 176.525 ;
        RECT 96.855 176.385 97.185 176.745 ;
        RECT 93.455 175.305 93.625 175.995 ;
        RECT 93.795 175.645 93.965 175.825 ;
        RECT 94.135 175.815 94.925 176.065 ;
        RECT 95.130 175.645 95.300 176.355 ;
        RECT 95.470 175.845 95.825 176.065 ;
        RECT 93.795 175.475 95.485 175.645 ;
        RECT 92.300 174.875 92.760 175.165 ;
        RECT 93.455 175.135 94.955 175.305 ;
        RECT 93.455 174.995 93.625 175.135 ;
        RECT 93.065 174.825 93.625 174.995 ;
        RECT 91.540 174.195 91.790 174.655 ;
        RECT 91.960 174.365 92.830 174.705 ;
        RECT 93.065 174.365 93.235 174.825 ;
        RECT 94.070 174.795 95.145 174.965 ;
        RECT 93.405 174.195 93.775 174.655 ;
        RECT 94.070 174.455 94.240 174.795 ;
        RECT 94.410 174.195 94.740 174.625 ;
        RECT 94.975 174.455 95.145 174.795 ;
        RECT 95.315 174.695 95.485 175.475 ;
        RECT 95.655 175.255 95.825 175.845 ;
        RECT 95.995 175.445 96.345 176.065 ;
        RECT 95.655 174.865 96.120 175.255 ;
        RECT 96.515 174.995 96.685 176.355 ;
        RECT 96.855 175.165 97.315 176.215 ;
        RECT 96.290 174.825 96.685 174.995 ;
        RECT 96.290 174.695 96.460 174.825 ;
        RECT 95.315 174.365 95.995 174.695 ;
        RECT 96.210 174.365 96.460 174.695 ;
        RECT 96.630 174.195 96.880 174.655 ;
        RECT 97.050 174.380 97.375 175.165 ;
        RECT 97.545 174.365 97.715 176.485 ;
        RECT 97.885 176.365 98.215 176.745 ;
        RECT 98.385 176.195 98.640 176.485 ;
        RECT 97.890 176.025 98.640 176.195 ;
        RECT 98.815 176.070 99.075 176.575 ;
        RECT 99.255 176.365 99.585 176.745 ;
        RECT 99.765 176.195 99.935 176.575 ;
        RECT 97.890 175.035 98.120 176.025 ;
        RECT 98.290 175.205 98.640 175.855 ;
        RECT 98.815 175.270 98.985 176.070 ;
        RECT 99.270 176.025 99.935 176.195 ;
        RECT 99.270 175.770 99.440 176.025 ;
        RECT 100.195 176.020 100.485 176.745 ;
        RECT 101.665 176.195 101.835 176.575 ;
        RECT 102.015 176.365 102.345 176.745 ;
        RECT 101.665 176.025 102.330 176.195 ;
        RECT 102.525 176.070 102.785 176.575 ;
        RECT 99.155 175.440 99.440 175.770 ;
        RECT 99.675 175.475 100.005 175.845 ;
        RECT 101.595 175.475 101.925 175.845 ;
        RECT 102.160 175.770 102.330 176.025 ;
        RECT 99.270 175.295 99.440 175.440 ;
        RECT 102.160 175.440 102.445 175.770 ;
        RECT 97.890 174.865 98.640 175.035 ;
        RECT 97.885 174.195 98.215 174.695 ;
        RECT 98.385 174.365 98.640 174.865 ;
        RECT 98.815 174.365 99.085 175.270 ;
        RECT 99.270 175.125 99.935 175.295 ;
        RECT 99.255 174.195 99.585 174.955 ;
        RECT 99.765 174.365 99.935 175.125 ;
        RECT 100.195 174.195 100.485 175.360 ;
        RECT 102.160 175.295 102.330 175.440 ;
        RECT 101.665 175.125 102.330 175.295 ;
        RECT 102.615 175.270 102.785 176.070 ;
        RECT 102.960 176.195 103.215 176.485 ;
        RECT 103.385 176.365 103.715 176.745 ;
        RECT 102.960 176.025 103.710 176.195 ;
        RECT 101.665 174.365 101.835 175.125 ;
        RECT 102.015 174.195 102.345 174.955 ;
        RECT 102.515 174.365 102.785 175.270 ;
        RECT 102.960 175.205 103.310 175.855 ;
        RECT 103.480 175.035 103.710 176.025 ;
        RECT 102.960 174.865 103.710 175.035 ;
        RECT 102.960 174.365 103.215 174.865 ;
        RECT 103.385 174.195 103.715 174.695 ;
        RECT 103.885 174.365 104.055 176.485 ;
        RECT 104.415 176.385 104.745 176.745 ;
        RECT 104.915 176.355 105.410 176.525 ;
        RECT 105.615 176.355 106.470 176.525 ;
        RECT 104.285 175.165 104.745 176.215 ;
        RECT 104.225 174.380 104.550 175.165 ;
        RECT 104.915 174.995 105.085 176.355 ;
        RECT 105.255 175.445 105.605 176.065 ;
        RECT 105.775 175.845 106.130 176.065 ;
        RECT 105.775 175.255 105.945 175.845 ;
        RECT 106.300 175.645 106.470 176.355 ;
        RECT 107.345 176.285 107.675 176.745 ;
        RECT 107.885 176.385 108.235 176.555 ;
        RECT 106.675 175.815 107.465 176.065 ;
        RECT 107.885 175.995 108.145 176.385 ;
        RECT 108.455 176.295 109.405 176.575 ;
        RECT 109.575 176.305 109.765 176.745 ;
        RECT 109.935 176.365 111.005 176.535 ;
        RECT 107.635 175.645 107.805 175.825 ;
        RECT 104.915 174.825 105.310 174.995 ;
        RECT 105.480 174.865 105.945 175.255 ;
        RECT 106.115 175.475 107.805 175.645 ;
        RECT 105.140 174.695 105.310 174.825 ;
        RECT 106.115 174.695 106.285 175.475 ;
        RECT 107.975 175.305 108.145 175.995 ;
        RECT 106.645 175.135 108.145 175.305 ;
        RECT 108.335 175.335 108.545 176.125 ;
        RECT 108.715 175.505 109.065 176.125 ;
        RECT 109.235 175.515 109.405 176.295 ;
        RECT 109.935 176.135 110.105 176.365 ;
        RECT 109.575 175.965 110.105 176.135 ;
        RECT 109.575 175.685 109.795 175.965 ;
        RECT 110.275 175.795 110.515 176.195 ;
        RECT 109.235 175.345 109.640 175.515 ;
        RECT 109.975 175.425 110.515 175.795 ;
        RECT 110.685 176.010 111.005 176.365 ;
        RECT 111.250 176.285 111.555 176.745 ;
        RECT 111.725 176.035 111.980 176.565 ;
        RECT 110.685 175.835 111.010 176.010 ;
        RECT 110.685 175.535 111.600 175.835 ;
        RECT 110.860 175.505 111.600 175.535 ;
        RECT 108.335 175.175 109.010 175.335 ;
        RECT 109.470 175.255 109.640 175.345 ;
        RECT 108.335 175.165 109.300 175.175 ;
        RECT 107.975 174.995 108.145 175.135 ;
        RECT 104.720 174.195 104.970 174.655 ;
        RECT 105.140 174.365 105.390 174.695 ;
        RECT 105.605 174.365 106.285 174.695 ;
        RECT 106.455 174.795 107.530 174.965 ;
        RECT 107.975 174.825 108.535 174.995 ;
        RECT 108.840 174.875 109.300 175.165 ;
        RECT 109.470 175.085 110.690 175.255 ;
        RECT 106.455 174.455 106.625 174.795 ;
        RECT 106.860 174.195 107.190 174.625 ;
        RECT 107.360 174.455 107.530 174.795 ;
        RECT 107.825 174.195 108.195 174.655 ;
        RECT 108.365 174.365 108.535 174.825 ;
        RECT 109.470 174.705 109.640 175.085 ;
        RECT 110.860 174.915 111.030 175.505 ;
        RECT 111.770 175.385 111.980 176.035 ;
        RECT 112.155 175.995 113.365 176.745 ;
        RECT 108.770 174.365 109.640 174.705 ;
        RECT 110.230 174.745 111.030 174.915 ;
        RECT 109.810 174.195 110.060 174.655 ;
        RECT 110.230 174.455 110.400 174.745 ;
        RECT 110.580 174.195 110.910 174.575 ;
        RECT 111.250 174.195 111.555 175.335 ;
        RECT 111.725 174.505 111.980 175.385 ;
        RECT 112.155 175.285 112.675 175.825 ;
        RECT 112.845 175.455 113.365 175.995 ;
        RECT 112.155 174.195 113.365 175.285 ;
        RECT 22.830 174.025 113.450 174.195 ;
        RECT 22.915 172.935 24.125 174.025 ;
        RECT 22.915 172.225 23.435 172.765 ;
        RECT 23.605 172.395 24.125 172.935 ;
        RECT 24.355 172.885 24.565 174.025 ;
        RECT 24.735 172.875 25.065 173.855 ;
        RECT 25.235 172.885 25.465 174.025 ;
        RECT 25.765 173.095 25.935 173.855 ;
        RECT 26.115 173.265 26.445 174.025 ;
        RECT 25.765 172.925 26.430 173.095 ;
        RECT 26.615 172.950 26.885 173.855 ;
        RECT 22.915 171.475 24.125 172.225 ;
        RECT 24.355 171.475 24.565 172.295 ;
        RECT 24.735 172.275 24.985 172.875 ;
        RECT 26.260 172.780 26.430 172.925 ;
        RECT 25.155 172.465 25.485 172.715 ;
        RECT 25.695 172.375 26.025 172.745 ;
        RECT 26.260 172.450 26.545 172.780 ;
        RECT 24.735 171.645 25.065 172.275 ;
        RECT 25.235 171.475 25.465 172.295 ;
        RECT 26.260 172.195 26.430 172.450 ;
        RECT 25.765 172.025 26.430 172.195 ;
        RECT 26.715 172.150 26.885 172.950 ;
        RECT 27.095 172.885 27.325 174.025 ;
        RECT 27.495 172.875 27.825 173.855 ;
        RECT 27.995 172.885 28.205 174.025 ;
        RECT 28.550 173.395 28.835 173.855 ;
        RECT 29.005 173.565 29.275 174.025 ;
        RECT 28.550 173.175 29.505 173.395 ;
        RECT 27.075 172.465 27.405 172.715 ;
        RECT 25.765 171.645 25.935 172.025 ;
        RECT 26.115 171.475 26.445 171.855 ;
        RECT 26.625 171.645 26.885 172.150 ;
        RECT 27.095 171.475 27.325 172.295 ;
        RECT 27.575 172.275 27.825 172.875 ;
        RECT 28.435 172.445 29.125 173.005 ;
        RECT 27.495 171.645 27.825 172.275 ;
        RECT 27.995 171.475 28.205 172.295 ;
        RECT 29.295 172.275 29.505 173.175 ;
        RECT 28.550 172.105 29.505 172.275 ;
        RECT 29.675 173.005 30.075 173.855 ;
        RECT 30.265 173.395 30.545 173.855 ;
        RECT 31.065 173.565 31.390 174.025 ;
        RECT 30.265 173.175 31.390 173.395 ;
        RECT 29.675 172.445 30.770 173.005 ;
        RECT 30.940 172.715 31.390 173.175 ;
        RECT 31.560 172.885 31.945 173.855 ;
        RECT 32.320 173.055 32.650 173.855 ;
        RECT 32.820 173.225 33.150 174.025 ;
        RECT 33.450 173.055 33.780 173.855 ;
        RECT 34.425 173.225 34.675 174.025 ;
        RECT 32.320 172.885 34.755 173.055 ;
        RECT 34.945 172.885 35.115 174.025 ;
        RECT 35.285 172.885 35.625 173.855 ;
        RECT 28.550 171.645 28.835 172.105 ;
        RECT 29.005 171.475 29.275 171.935 ;
        RECT 29.675 171.645 30.075 172.445 ;
        RECT 30.940 172.385 31.495 172.715 ;
        RECT 30.940 172.275 31.390 172.385 ;
        RECT 30.265 172.105 31.390 172.275 ;
        RECT 31.665 172.215 31.945 172.885 ;
        RECT 32.115 172.465 32.465 172.715 ;
        RECT 32.650 172.255 32.820 172.885 ;
        RECT 32.990 172.465 33.320 172.665 ;
        RECT 33.490 172.465 33.820 172.665 ;
        RECT 33.990 172.465 34.410 172.665 ;
        RECT 34.585 172.635 34.755 172.885 ;
        RECT 34.585 172.465 35.280 172.635 ;
        RECT 30.265 171.645 30.545 172.105 ;
        RECT 31.065 171.475 31.390 171.935 ;
        RECT 31.560 171.645 31.945 172.215 ;
        RECT 32.320 171.645 32.820 172.255 ;
        RECT 33.450 172.125 34.675 172.295 ;
        RECT 35.450 172.275 35.625 172.885 ;
        RECT 35.795 172.860 36.085 174.025 ;
        RECT 36.345 173.280 36.615 174.025 ;
        RECT 37.245 174.020 43.520 174.025 ;
        RECT 36.785 173.110 37.075 173.850 ;
        RECT 37.245 173.295 37.500 174.020 ;
        RECT 37.685 173.125 37.945 173.850 ;
        RECT 38.115 173.295 38.360 174.020 ;
        RECT 38.545 173.125 38.805 173.850 ;
        RECT 38.975 173.295 39.220 174.020 ;
        RECT 39.405 173.125 39.665 173.850 ;
        RECT 39.835 173.295 40.080 174.020 ;
        RECT 40.250 173.125 40.510 173.850 ;
        RECT 40.680 173.295 40.940 174.020 ;
        RECT 41.110 173.125 41.370 173.850 ;
        RECT 41.540 173.295 41.800 174.020 ;
        RECT 41.970 173.125 42.230 173.850 ;
        RECT 42.400 173.295 42.660 174.020 ;
        RECT 42.830 173.125 43.090 173.850 ;
        RECT 43.260 173.225 43.520 174.020 ;
        RECT 37.685 173.110 43.090 173.125 ;
        RECT 36.345 173.005 43.090 173.110 ;
        RECT 36.315 172.885 43.090 173.005 ;
        RECT 36.315 172.835 37.510 172.885 ;
        RECT 33.450 171.645 33.780 172.125 ;
        RECT 33.950 171.475 34.175 171.935 ;
        RECT 34.345 171.645 34.675 172.125 ;
        RECT 34.865 171.475 35.115 172.275 ;
        RECT 35.285 171.645 35.625 172.275 ;
        RECT 36.345 172.295 37.510 172.835 ;
        RECT 43.690 172.715 43.940 173.850 ;
        RECT 44.120 173.215 44.380 174.025 ;
        RECT 44.555 172.715 44.800 173.855 ;
        RECT 44.980 173.215 45.275 174.025 ;
        RECT 45.515 172.885 45.725 174.025 ;
        RECT 45.895 172.875 46.225 173.855 ;
        RECT 46.395 172.885 46.625 174.025 ;
        RECT 46.845 173.215 47.140 174.025 ;
        RECT 37.680 172.465 44.800 172.715 ;
        RECT 35.795 171.475 36.085 172.200 ;
        RECT 36.345 172.125 43.090 172.295 ;
        RECT 36.345 171.475 36.645 171.955 ;
        RECT 36.815 171.670 37.075 172.125 ;
        RECT 37.245 171.475 37.505 171.955 ;
        RECT 37.685 171.670 37.945 172.125 ;
        RECT 38.115 171.475 38.365 171.955 ;
        RECT 38.545 171.670 38.805 172.125 ;
        RECT 38.975 171.475 39.225 171.955 ;
        RECT 39.405 171.670 39.665 172.125 ;
        RECT 39.835 171.475 40.080 171.955 ;
        RECT 40.250 171.670 40.525 172.125 ;
        RECT 40.695 171.475 40.940 171.955 ;
        RECT 41.110 171.670 41.370 172.125 ;
        RECT 41.540 171.475 41.800 171.955 ;
        RECT 41.970 171.670 42.230 172.125 ;
        RECT 42.400 171.475 42.660 171.955 ;
        RECT 42.830 171.670 43.090 172.125 ;
        RECT 43.260 171.475 43.520 172.035 ;
        RECT 43.690 171.655 43.940 172.465 ;
        RECT 44.120 171.475 44.380 172.000 ;
        RECT 44.550 171.655 44.800 172.465 ;
        RECT 44.970 172.155 45.285 172.715 ;
        RECT 44.980 171.475 45.285 171.985 ;
        RECT 45.515 171.475 45.725 172.295 ;
        RECT 45.895 172.275 46.145 172.875 ;
        RECT 47.320 172.715 47.565 173.855 ;
        RECT 47.740 173.215 48.000 174.025 ;
        RECT 48.600 174.020 54.875 174.025 ;
        RECT 48.180 172.715 48.430 173.850 ;
        RECT 48.600 173.225 48.860 174.020 ;
        RECT 49.030 173.125 49.290 173.850 ;
        RECT 49.460 173.295 49.720 174.020 ;
        RECT 49.890 173.125 50.150 173.850 ;
        RECT 50.320 173.295 50.580 174.020 ;
        RECT 50.750 173.125 51.010 173.850 ;
        RECT 51.180 173.295 51.440 174.020 ;
        RECT 51.610 173.125 51.870 173.850 ;
        RECT 52.040 173.295 52.285 174.020 ;
        RECT 52.455 173.125 52.715 173.850 ;
        RECT 52.900 173.295 53.145 174.020 ;
        RECT 53.315 173.125 53.575 173.850 ;
        RECT 53.760 173.295 54.005 174.020 ;
        RECT 54.175 173.125 54.435 173.850 ;
        RECT 54.620 173.295 54.875 174.020 ;
        RECT 49.030 173.110 54.435 173.125 ;
        RECT 55.045 173.110 55.335 173.850 ;
        RECT 55.505 173.280 55.775 174.025 ;
        RECT 49.030 172.885 55.775 173.110 ;
        RECT 46.315 172.465 46.645 172.715 ;
        RECT 45.895 171.645 46.225 172.275 ;
        RECT 46.395 171.475 46.625 172.295 ;
        RECT 46.835 172.155 47.150 172.715 ;
        RECT 47.320 172.465 54.440 172.715 ;
        RECT 46.835 171.475 47.140 171.985 ;
        RECT 47.320 171.655 47.570 172.465 ;
        RECT 47.740 171.475 48.000 172.000 ;
        RECT 48.180 171.655 48.430 172.465 ;
        RECT 54.610 172.325 55.775 172.885 ;
        RECT 56.495 172.935 60.005 174.025 ;
        RECT 56.495 172.415 58.185 172.935 ;
        RECT 60.215 172.885 60.445 174.025 ;
        RECT 60.615 172.875 60.945 173.855 ;
        RECT 61.115 172.885 61.325 174.025 ;
        RECT 54.610 172.295 55.805 172.325 ;
        RECT 49.030 172.155 55.805 172.295 ;
        RECT 58.355 172.245 60.005 172.765 ;
        RECT 60.195 172.465 60.525 172.715 ;
        RECT 49.030 172.125 55.775 172.155 ;
        RECT 48.600 171.475 48.860 172.035 ;
        RECT 49.030 171.670 49.290 172.125 ;
        RECT 49.460 171.475 49.720 171.955 ;
        RECT 49.890 171.670 50.150 172.125 ;
        RECT 50.320 171.475 50.580 171.955 ;
        RECT 50.750 171.670 51.010 172.125 ;
        RECT 51.180 171.475 51.425 171.955 ;
        RECT 51.595 171.670 51.870 172.125 ;
        RECT 52.040 171.475 52.285 171.955 ;
        RECT 52.455 171.670 52.715 172.125 ;
        RECT 52.895 171.475 53.145 171.955 ;
        RECT 53.315 171.670 53.575 172.125 ;
        RECT 53.755 171.475 54.005 171.955 ;
        RECT 54.175 171.670 54.435 172.125 ;
        RECT 54.615 171.475 54.875 171.955 ;
        RECT 55.045 171.670 55.305 172.125 ;
        RECT 55.475 171.475 55.775 171.955 ;
        RECT 56.495 171.475 60.005 172.245 ;
        RECT 60.215 171.475 60.445 172.295 ;
        RECT 60.695 172.275 60.945 172.875 ;
        RECT 61.555 172.860 61.845 174.025 ;
        RECT 62.020 172.875 62.280 174.025 ;
        RECT 62.455 172.950 62.710 173.855 ;
        RECT 62.880 173.265 63.210 174.025 ;
        RECT 63.425 173.095 63.595 173.855 ;
        RECT 63.910 173.155 64.195 174.025 ;
        RECT 64.365 173.395 64.625 173.855 ;
        RECT 64.800 173.565 65.055 174.025 ;
        RECT 65.225 173.395 65.485 173.855 ;
        RECT 64.365 173.225 65.485 173.395 ;
        RECT 65.655 173.225 65.965 174.025 ;
        RECT 60.615 171.645 60.945 172.275 ;
        RECT 61.115 171.475 61.325 172.295 ;
        RECT 61.555 171.475 61.845 172.200 ;
        RECT 62.020 171.475 62.280 172.315 ;
        RECT 62.455 172.220 62.625 172.950 ;
        RECT 62.880 172.925 63.595 173.095 ;
        RECT 64.365 172.975 64.625 173.225 ;
        RECT 64.835 173.175 65.005 173.225 ;
        RECT 66.135 173.055 66.445 173.855 ;
        RECT 62.880 172.715 63.050 172.925 ;
        RECT 63.870 172.805 64.625 172.975 ;
        RECT 65.415 172.885 66.445 173.055 ;
        RECT 62.795 172.385 63.050 172.715 ;
        RECT 62.455 171.645 62.710 172.220 ;
        RECT 62.880 172.195 63.050 172.385 ;
        RECT 63.330 172.375 63.685 172.745 ;
        RECT 63.870 172.295 64.275 172.805 ;
        RECT 65.415 172.635 65.585 172.885 ;
        RECT 64.445 172.465 65.585 172.635 ;
        RECT 62.880 172.025 63.595 172.195 ;
        RECT 63.870 172.125 65.520 172.295 ;
        RECT 65.755 172.145 66.105 172.715 ;
        RECT 62.880 171.475 63.210 171.855 ;
        RECT 63.425 171.645 63.595 172.025 ;
        RECT 63.915 171.475 64.195 171.955 ;
        RECT 64.365 171.735 64.625 172.125 ;
        RECT 64.800 171.475 65.055 171.955 ;
        RECT 65.225 171.735 65.520 172.125 ;
        RECT 66.275 171.975 66.445 172.885 ;
        RECT 66.990 173.045 67.245 173.715 ;
        RECT 67.425 173.225 67.710 174.025 ;
        RECT 67.890 173.305 68.220 173.815 ;
        RECT 66.990 172.185 67.170 173.045 ;
        RECT 67.890 172.715 68.140 173.305 ;
        RECT 68.490 173.155 68.660 173.765 ;
        RECT 68.830 173.335 69.160 174.025 ;
        RECT 69.390 173.475 69.630 173.765 ;
        RECT 69.830 173.645 70.250 174.025 ;
        RECT 70.430 173.555 71.060 173.805 ;
        RECT 71.530 173.645 71.860 174.025 ;
        RECT 70.430 173.475 70.600 173.555 ;
        RECT 72.030 173.475 72.200 173.765 ;
        RECT 72.380 173.645 72.760 174.025 ;
        RECT 73.000 173.640 73.830 173.810 ;
        RECT 69.390 173.305 70.600 173.475 ;
        RECT 67.340 172.385 68.140 172.715 ;
        RECT 66.990 171.985 67.245 172.185 ;
        RECT 65.700 171.475 65.975 171.955 ;
        RECT 66.145 171.645 66.445 171.975 ;
        RECT 66.905 171.815 67.245 171.985 ;
        RECT 66.990 171.655 67.245 171.815 ;
        RECT 67.425 171.475 67.710 171.935 ;
        RECT 67.890 171.735 68.140 172.385 ;
        RECT 68.340 173.135 68.660 173.155 ;
        RECT 68.340 172.965 70.260 173.135 ;
        RECT 68.340 172.070 68.530 172.965 ;
        RECT 70.430 172.795 70.600 173.305 ;
        RECT 70.770 173.045 71.290 173.355 ;
        RECT 68.700 172.625 70.600 172.795 ;
        RECT 68.700 172.565 69.030 172.625 ;
        RECT 69.180 172.395 69.510 172.455 ;
        RECT 68.850 172.125 69.510 172.395 ;
        RECT 68.340 171.740 68.660 172.070 ;
        RECT 68.840 171.475 69.500 171.955 ;
        RECT 69.700 171.865 69.870 172.625 ;
        RECT 70.770 172.455 70.950 172.865 ;
        RECT 70.040 172.285 70.370 172.405 ;
        RECT 71.120 172.285 71.290 173.045 ;
        RECT 70.040 172.115 71.290 172.285 ;
        RECT 71.460 173.225 72.830 173.475 ;
        RECT 71.460 172.455 71.650 173.225 ;
        RECT 72.580 172.965 72.830 173.225 ;
        RECT 71.820 172.795 72.070 172.955 ;
        RECT 73.000 172.795 73.170 173.640 ;
        RECT 74.065 173.355 74.235 173.855 ;
        RECT 74.405 173.525 74.735 174.025 ;
        RECT 73.340 172.965 73.840 173.345 ;
        RECT 74.065 173.185 74.760 173.355 ;
        RECT 71.820 172.625 73.170 172.795 ;
        RECT 72.750 172.585 73.170 172.625 ;
        RECT 71.460 172.115 71.880 172.455 ;
        RECT 72.170 172.125 72.580 172.455 ;
        RECT 69.700 171.695 70.550 171.865 ;
        RECT 71.110 171.475 71.430 171.935 ;
        RECT 71.630 171.685 71.880 172.115 ;
        RECT 72.170 171.475 72.580 171.915 ;
        RECT 72.750 171.855 72.920 172.585 ;
        RECT 73.090 172.035 73.440 172.405 ;
        RECT 73.620 172.095 73.840 172.965 ;
        RECT 74.010 172.395 74.420 173.015 ;
        RECT 74.590 172.215 74.760 173.185 ;
        RECT 74.065 172.025 74.760 172.215 ;
        RECT 72.750 171.655 73.765 171.855 ;
        RECT 74.065 171.695 74.235 172.025 ;
        RECT 74.405 171.475 74.735 171.855 ;
        RECT 74.950 171.735 75.175 173.855 ;
        RECT 75.345 173.525 75.675 174.025 ;
        RECT 75.845 173.355 76.015 173.855 ;
        RECT 75.350 173.185 76.015 173.355 ;
        RECT 76.385 173.225 76.555 174.025 ;
        RECT 75.350 172.195 75.580 173.185 ;
        RECT 75.750 172.365 76.100 173.015 ;
        RECT 76.725 173.005 77.055 173.855 ;
        RECT 77.225 173.225 77.395 174.025 ;
        RECT 77.565 173.005 77.895 173.855 ;
        RECT 78.065 173.225 78.235 174.025 ;
        RECT 78.405 173.005 78.735 173.855 ;
        RECT 78.905 173.225 79.075 174.025 ;
        RECT 79.245 173.005 79.575 173.855 ;
        RECT 79.745 173.225 79.915 174.025 ;
        RECT 80.085 173.005 80.415 173.855 ;
        RECT 80.585 173.225 80.755 174.025 ;
        RECT 80.925 173.005 81.255 173.855 ;
        RECT 81.425 173.225 81.595 174.025 ;
        RECT 81.765 173.005 82.095 173.855 ;
        RECT 82.265 173.225 82.435 174.025 ;
        RECT 82.605 173.005 82.935 173.855 ;
        RECT 83.105 173.225 83.275 174.025 ;
        RECT 83.445 173.005 83.775 173.855 ;
        RECT 83.945 173.225 84.115 174.025 ;
        RECT 84.285 173.005 84.615 173.855 ;
        RECT 84.785 173.225 84.955 174.025 ;
        RECT 85.125 173.005 85.455 173.855 ;
        RECT 85.625 173.175 85.795 174.025 ;
        RECT 85.965 173.005 86.295 173.855 ;
        RECT 86.465 173.175 86.635 174.025 ;
        RECT 86.805 173.005 87.135 173.855 ;
        RECT 76.275 172.835 82.935 173.005 ;
        RECT 83.105 172.835 85.455 173.005 ;
        RECT 85.625 172.835 87.135 173.005 ;
        RECT 87.315 172.860 87.605 174.025 ;
        RECT 87.815 172.885 88.045 174.025 ;
        RECT 88.215 172.875 88.545 173.855 ;
        RECT 88.715 172.885 88.925 174.025 ;
        RECT 89.195 172.885 89.425 174.025 ;
        RECT 89.595 172.875 89.925 173.855 ;
        RECT 90.095 172.885 90.305 174.025 ;
        RECT 76.275 172.295 76.550 172.835 ;
        RECT 83.105 172.665 83.280 172.835 ;
        RECT 85.625 172.665 85.795 172.835 ;
        RECT 76.720 172.465 83.280 172.665 ;
        RECT 83.485 172.465 85.795 172.665 ;
        RECT 85.965 172.465 87.140 172.665 ;
        RECT 87.795 172.465 88.125 172.715 ;
        RECT 83.105 172.295 83.280 172.465 ;
        RECT 85.625 172.295 85.795 172.465 ;
        RECT 75.350 172.025 76.015 172.195 ;
        RECT 76.275 172.125 82.935 172.295 ;
        RECT 83.105 172.125 85.455 172.295 ;
        RECT 85.625 172.125 87.135 172.295 ;
        RECT 75.345 171.475 75.675 171.855 ;
        RECT 75.845 171.735 76.015 172.025 ;
        RECT 76.385 171.475 76.555 171.955 ;
        RECT 76.725 171.650 77.055 172.125 ;
        RECT 77.225 171.475 77.395 171.955 ;
        RECT 77.565 171.650 77.895 172.125 ;
        RECT 78.065 171.475 78.235 171.955 ;
        RECT 78.405 171.650 78.735 172.125 ;
        RECT 78.905 171.475 79.075 171.955 ;
        RECT 79.245 171.650 79.575 172.125 ;
        RECT 79.745 171.475 79.915 171.955 ;
        RECT 80.085 171.650 80.415 172.125 ;
        RECT 80.585 171.475 80.755 171.955 ;
        RECT 80.925 171.650 81.255 172.125 ;
        RECT 81.005 171.645 81.175 171.650 ;
        RECT 81.425 171.475 81.595 171.955 ;
        RECT 81.765 171.650 82.095 172.125 ;
        RECT 81.845 171.645 82.015 171.650 ;
        RECT 82.265 171.475 82.435 171.955 ;
        RECT 82.605 171.650 82.935 172.125 ;
        RECT 82.685 171.645 82.935 171.650 ;
        RECT 83.105 171.475 83.275 171.955 ;
        RECT 83.445 171.650 83.775 172.125 ;
        RECT 83.945 171.475 84.115 171.955 ;
        RECT 84.285 171.650 84.615 172.125 ;
        RECT 84.785 171.475 84.955 171.955 ;
        RECT 85.125 171.650 85.455 172.125 ;
        RECT 85.625 171.475 85.795 171.955 ;
        RECT 85.965 171.650 86.295 172.125 ;
        RECT 86.465 171.475 86.635 171.955 ;
        RECT 86.805 171.650 87.135 172.125 ;
        RECT 87.315 171.475 87.605 172.200 ;
        RECT 87.815 171.475 88.045 172.295 ;
        RECT 88.295 172.275 88.545 172.875 ;
        RECT 89.175 172.465 89.505 172.715 ;
        RECT 88.215 171.645 88.545 172.275 ;
        RECT 88.715 171.475 88.925 172.295 ;
        RECT 89.195 171.475 89.425 172.295 ;
        RECT 89.675 172.275 89.925 172.875 ;
        RECT 91.000 172.835 91.255 173.715 ;
        RECT 91.425 172.885 91.730 174.025 ;
        RECT 92.070 173.645 92.400 174.025 ;
        RECT 92.580 173.475 92.750 173.765 ;
        RECT 92.920 173.565 93.170 174.025 ;
        RECT 91.950 173.305 92.750 173.475 ;
        RECT 93.340 173.515 94.210 173.855 ;
        RECT 89.595 171.645 89.925 172.275 ;
        RECT 90.095 171.475 90.305 172.295 ;
        RECT 91.000 172.185 91.210 172.835 ;
        RECT 91.950 172.715 92.120 173.305 ;
        RECT 93.340 173.135 93.510 173.515 ;
        RECT 94.445 173.395 94.615 173.855 ;
        RECT 94.785 173.565 95.155 174.025 ;
        RECT 95.450 173.425 95.620 173.765 ;
        RECT 95.790 173.595 96.120 174.025 ;
        RECT 96.355 173.425 96.525 173.765 ;
        RECT 92.290 172.965 93.510 173.135 ;
        RECT 93.680 173.055 94.140 173.345 ;
        RECT 94.445 173.225 95.005 173.395 ;
        RECT 95.450 173.255 96.525 173.425 ;
        RECT 96.695 173.525 97.375 173.855 ;
        RECT 97.590 173.525 97.840 173.855 ;
        RECT 98.010 173.565 98.260 174.025 ;
        RECT 94.835 173.085 95.005 173.225 ;
        RECT 93.680 173.045 94.645 173.055 ;
        RECT 93.340 172.875 93.510 172.965 ;
        RECT 93.970 172.885 94.645 173.045 ;
        RECT 91.380 172.685 92.120 172.715 ;
        RECT 91.380 172.385 92.295 172.685 ;
        RECT 91.970 172.210 92.295 172.385 ;
        RECT 91.000 171.655 91.255 172.185 ;
        RECT 91.425 171.475 91.730 171.935 ;
        RECT 91.975 171.855 92.295 172.210 ;
        RECT 92.465 172.425 93.005 172.795 ;
        RECT 93.340 172.705 93.745 172.875 ;
        RECT 92.465 172.025 92.705 172.425 ;
        RECT 93.185 172.255 93.405 172.535 ;
        RECT 92.875 172.085 93.405 172.255 ;
        RECT 92.875 171.855 93.045 172.085 ;
        RECT 93.575 171.925 93.745 172.705 ;
        RECT 93.915 172.095 94.265 172.715 ;
        RECT 94.435 172.095 94.645 172.885 ;
        RECT 94.835 172.915 96.335 173.085 ;
        RECT 94.835 172.225 95.005 172.915 ;
        RECT 96.695 172.745 96.865 173.525 ;
        RECT 97.670 173.395 97.840 173.525 ;
        RECT 95.175 172.575 96.865 172.745 ;
        RECT 97.035 172.965 97.500 173.355 ;
        RECT 97.670 173.225 98.065 173.395 ;
        RECT 95.175 172.395 95.345 172.575 ;
        RECT 91.975 171.685 93.045 171.855 ;
        RECT 93.215 171.475 93.405 171.915 ;
        RECT 93.575 171.645 94.525 171.925 ;
        RECT 94.835 171.835 95.095 172.225 ;
        RECT 95.515 172.155 96.305 172.405 ;
        RECT 94.745 171.665 95.095 171.835 ;
        RECT 95.305 171.475 95.635 171.935 ;
        RECT 96.510 171.865 96.680 172.575 ;
        RECT 97.035 172.375 97.205 172.965 ;
        RECT 96.850 172.155 97.205 172.375 ;
        RECT 97.375 172.155 97.725 172.775 ;
        RECT 97.895 171.865 98.065 173.225 ;
        RECT 98.430 173.055 98.755 173.840 ;
        RECT 98.235 172.005 98.695 173.055 ;
        RECT 96.510 171.695 97.365 171.865 ;
        RECT 97.570 171.695 98.065 171.865 ;
        RECT 98.235 171.475 98.565 171.835 ;
        RECT 98.925 171.735 99.095 173.855 ;
        RECT 99.265 173.525 99.595 174.025 ;
        RECT 99.765 173.355 100.020 173.855 ;
        RECT 99.270 173.185 100.020 173.355 ;
        RECT 99.270 172.195 99.500 173.185 ;
        RECT 99.670 172.365 100.020 173.015 ;
        RECT 100.200 172.835 100.455 173.715 ;
        RECT 100.625 172.885 100.930 174.025 ;
        RECT 101.270 173.645 101.600 174.025 ;
        RECT 101.780 173.475 101.950 173.765 ;
        RECT 102.120 173.565 102.370 174.025 ;
        RECT 101.150 173.305 101.950 173.475 ;
        RECT 102.540 173.515 103.410 173.855 ;
        RECT 99.270 172.025 100.020 172.195 ;
        RECT 99.265 171.475 99.595 171.855 ;
        RECT 99.765 171.735 100.020 172.025 ;
        RECT 100.200 172.185 100.410 172.835 ;
        RECT 101.150 172.715 101.320 173.305 ;
        RECT 102.540 173.135 102.710 173.515 ;
        RECT 103.645 173.395 103.815 173.855 ;
        RECT 103.985 173.565 104.355 174.025 ;
        RECT 104.650 173.425 104.820 173.765 ;
        RECT 104.990 173.595 105.320 174.025 ;
        RECT 105.555 173.425 105.725 173.765 ;
        RECT 101.490 172.965 102.710 173.135 ;
        RECT 102.880 173.055 103.340 173.345 ;
        RECT 103.645 173.225 104.205 173.395 ;
        RECT 104.650 173.255 105.725 173.425 ;
        RECT 105.895 173.525 106.575 173.855 ;
        RECT 106.790 173.525 107.040 173.855 ;
        RECT 107.210 173.565 107.460 174.025 ;
        RECT 104.035 173.085 104.205 173.225 ;
        RECT 102.880 173.045 103.845 173.055 ;
        RECT 102.540 172.875 102.710 172.965 ;
        RECT 103.170 172.885 103.845 173.045 ;
        RECT 100.580 172.685 101.320 172.715 ;
        RECT 100.580 172.385 101.495 172.685 ;
        RECT 101.170 172.210 101.495 172.385 ;
        RECT 100.200 171.655 100.455 172.185 ;
        RECT 100.625 171.475 100.930 171.935 ;
        RECT 101.175 171.855 101.495 172.210 ;
        RECT 101.665 172.425 102.205 172.795 ;
        RECT 102.540 172.705 102.945 172.875 ;
        RECT 101.665 172.025 101.905 172.425 ;
        RECT 102.385 172.255 102.605 172.535 ;
        RECT 102.075 172.085 102.605 172.255 ;
        RECT 102.075 171.855 102.245 172.085 ;
        RECT 102.775 171.925 102.945 172.705 ;
        RECT 103.115 172.095 103.465 172.715 ;
        RECT 103.635 172.095 103.845 172.885 ;
        RECT 104.035 172.915 105.535 173.085 ;
        RECT 104.035 172.225 104.205 172.915 ;
        RECT 105.895 172.745 106.065 173.525 ;
        RECT 106.870 173.395 107.040 173.525 ;
        RECT 104.375 172.575 106.065 172.745 ;
        RECT 106.235 172.965 106.700 173.355 ;
        RECT 106.870 173.225 107.265 173.395 ;
        RECT 104.375 172.395 104.545 172.575 ;
        RECT 101.175 171.685 102.245 171.855 ;
        RECT 102.415 171.475 102.605 171.915 ;
        RECT 102.775 171.645 103.725 171.925 ;
        RECT 104.035 171.835 104.295 172.225 ;
        RECT 104.715 172.155 105.505 172.405 ;
        RECT 103.945 171.665 104.295 171.835 ;
        RECT 104.505 171.475 104.835 171.935 ;
        RECT 105.710 171.865 105.880 172.575 ;
        RECT 106.235 172.375 106.405 172.965 ;
        RECT 106.050 172.155 106.405 172.375 ;
        RECT 106.575 172.155 106.925 172.775 ;
        RECT 107.095 171.865 107.265 173.225 ;
        RECT 107.630 173.055 107.955 173.840 ;
        RECT 107.435 172.005 107.895 173.055 ;
        RECT 105.710 171.695 106.565 171.865 ;
        RECT 106.770 171.695 107.265 171.865 ;
        RECT 107.435 171.475 107.765 171.835 ;
        RECT 108.125 171.735 108.295 173.855 ;
        RECT 108.465 173.525 108.795 174.025 ;
        RECT 108.965 173.355 109.220 173.855 ;
        RECT 108.470 173.185 109.220 173.355 ;
        RECT 108.470 172.195 108.700 173.185 ;
        RECT 108.870 172.365 109.220 173.015 ;
        RECT 109.545 172.875 109.875 174.025 ;
        RECT 110.045 173.005 110.215 173.855 ;
        RECT 110.385 173.225 110.715 174.025 ;
        RECT 110.885 173.005 111.055 173.855 ;
        RECT 111.235 173.225 111.475 174.025 ;
        RECT 111.645 173.045 111.975 173.855 ;
        RECT 110.045 172.835 111.055 173.005 ;
        RECT 111.260 172.875 111.975 173.045 ;
        RECT 112.155 172.935 113.365 174.025 ;
        RECT 110.045 172.325 110.540 172.835 ;
        RECT 111.260 172.635 111.430 172.875 ;
        RECT 110.930 172.465 111.430 172.635 ;
        RECT 111.600 172.465 111.980 172.705 ;
        RECT 110.045 172.295 110.545 172.325 ;
        RECT 111.260 172.295 111.430 172.465 ;
        RECT 112.155 172.395 112.675 172.935 ;
        RECT 108.470 172.025 109.220 172.195 ;
        RECT 108.465 171.475 108.795 171.855 ;
        RECT 108.965 171.735 109.220 172.025 ;
        RECT 109.545 171.475 109.875 172.275 ;
        RECT 110.045 172.125 111.055 172.295 ;
        RECT 111.260 172.125 111.895 172.295 ;
        RECT 112.845 172.225 113.365 172.765 ;
        RECT 110.045 171.645 110.215 172.125 ;
        RECT 110.385 171.475 110.715 171.955 ;
        RECT 110.885 171.645 111.055 172.125 ;
        RECT 111.305 171.475 111.545 171.955 ;
        RECT 111.725 171.645 111.895 172.125 ;
        RECT 112.155 171.475 113.365 172.225 ;
        RECT 22.830 171.305 113.450 171.475 ;
        RECT 22.915 170.555 24.125 171.305 ;
        RECT 25.590 170.595 25.845 171.125 ;
        RECT 26.025 170.845 26.310 171.305 ;
        RECT 22.915 170.015 23.435 170.555 ;
        RECT 23.605 169.845 24.125 170.385 ;
        RECT 22.915 168.755 24.125 169.845 ;
        RECT 25.590 169.735 25.770 170.595 ;
        RECT 26.490 170.395 26.740 171.045 ;
        RECT 25.940 170.065 26.740 170.395 ;
        RECT 25.590 169.265 25.845 169.735 ;
        RECT 25.505 169.095 25.845 169.265 ;
        RECT 25.590 169.065 25.845 169.095 ;
        RECT 26.025 168.755 26.310 169.555 ;
        RECT 26.490 169.475 26.740 170.065 ;
        RECT 26.940 170.710 27.260 171.040 ;
        RECT 27.440 170.825 28.100 171.305 ;
        RECT 28.300 170.915 29.150 171.085 ;
        RECT 26.940 169.815 27.130 170.710 ;
        RECT 27.450 170.385 28.110 170.655 ;
        RECT 27.780 170.325 28.110 170.385 ;
        RECT 27.300 170.155 27.630 170.215 ;
        RECT 28.300 170.155 28.470 170.915 ;
        RECT 29.710 170.845 30.030 171.305 ;
        RECT 30.230 170.665 30.480 171.095 ;
        RECT 30.770 170.865 31.180 171.305 ;
        RECT 31.350 170.925 32.365 171.125 ;
        RECT 28.640 170.495 29.890 170.665 ;
        RECT 28.640 170.375 28.970 170.495 ;
        RECT 27.300 169.985 29.200 170.155 ;
        RECT 26.940 169.645 28.860 169.815 ;
        RECT 26.940 169.625 27.260 169.645 ;
        RECT 26.490 168.965 26.820 169.475 ;
        RECT 27.090 169.015 27.260 169.625 ;
        RECT 29.030 169.475 29.200 169.985 ;
        RECT 29.370 169.915 29.550 170.325 ;
        RECT 29.720 169.735 29.890 170.495 ;
        RECT 27.430 168.755 27.760 169.445 ;
        RECT 27.990 169.305 29.200 169.475 ;
        RECT 29.370 169.425 29.890 169.735 ;
        RECT 30.060 170.325 30.480 170.665 ;
        RECT 30.770 170.325 31.180 170.655 ;
        RECT 30.060 169.555 30.250 170.325 ;
        RECT 31.350 170.195 31.520 170.925 ;
        RECT 32.665 170.755 32.835 171.085 ;
        RECT 33.005 170.925 33.335 171.305 ;
        RECT 31.690 170.375 32.040 170.745 ;
        RECT 31.350 170.155 31.770 170.195 ;
        RECT 30.420 169.985 31.770 170.155 ;
        RECT 30.420 169.825 30.670 169.985 ;
        RECT 31.180 169.555 31.430 169.815 ;
        RECT 30.060 169.305 31.430 169.555 ;
        RECT 27.990 169.015 28.230 169.305 ;
        RECT 29.030 169.225 29.200 169.305 ;
        RECT 28.430 168.755 28.850 169.135 ;
        RECT 29.030 168.975 29.660 169.225 ;
        RECT 30.130 168.755 30.460 169.135 ;
        RECT 30.630 169.015 30.800 169.305 ;
        RECT 31.600 169.140 31.770 169.985 ;
        RECT 32.220 169.815 32.440 170.685 ;
        RECT 32.665 170.565 33.360 170.755 ;
        RECT 31.940 169.435 32.440 169.815 ;
        RECT 32.610 169.765 33.020 170.385 ;
        RECT 33.190 169.595 33.360 170.565 ;
        RECT 32.665 169.425 33.360 169.595 ;
        RECT 30.980 168.755 31.360 169.135 ;
        RECT 31.600 168.970 32.430 169.140 ;
        RECT 32.665 168.925 32.835 169.425 ;
        RECT 33.005 168.755 33.335 169.255 ;
        RECT 33.550 168.925 33.775 171.045 ;
        RECT 33.945 170.925 34.275 171.305 ;
        RECT 34.445 170.755 34.615 171.045 ;
        RECT 33.950 170.585 34.615 170.755 ;
        RECT 33.950 169.595 34.180 170.585 ;
        RECT 36.000 170.525 36.500 171.135 ;
        RECT 34.350 169.765 34.700 170.415 ;
        RECT 35.795 170.065 36.145 170.315 ;
        RECT 36.330 169.895 36.500 170.525 ;
        RECT 37.130 170.655 37.460 171.135 ;
        RECT 37.630 170.845 37.855 171.305 ;
        RECT 38.025 170.655 38.355 171.135 ;
        RECT 37.130 170.485 38.355 170.655 ;
        RECT 38.545 170.505 38.795 171.305 ;
        RECT 38.965 170.505 39.305 171.135 ;
        RECT 36.670 170.115 37.000 170.315 ;
        RECT 37.170 170.115 37.500 170.315 ;
        RECT 37.670 170.115 38.090 170.315 ;
        RECT 38.265 170.145 38.960 170.315 ;
        RECT 38.265 169.895 38.435 170.145 ;
        RECT 39.130 169.895 39.305 170.505 ;
        RECT 36.000 169.725 38.435 169.895 ;
        RECT 33.950 169.425 34.615 169.595 ;
        RECT 33.945 168.755 34.275 169.255 ;
        RECT 34.445 168.925 34.615 169.425 ;
        RECT 36.000 168.925 36.330 169.725 ;
        RECT 36.500 168.755 36.830 169.555 ;
        RECT 37.130 168.925 37.460 169.725 ;
        RECT 38.105 168.755 38.355 169.555 ;
        RECT 38.625 168.755 38.795 169.895 ;
        RECT 38.965 168.925 39.305 169.895 ;
        RECT 39.480 170.595 39.735 171.125 ;
        RECT 39.905 170.845 40.210 171.305 ;
        RECT 40.455 170.925 41.525 171.095 ;
        RECT 39.480 169.945 39.690 170.595 ;
        RECT 40.455 170.570 40.775 170.925 ;
        RECT 40.450 170.395 40.775 170.570 ;
        RECT 39.860 170.095 40.775 170.395 ;
        RECT 40.945 170.355 41.185 170.755 ;
        RECT 41.355 170.695 41.525 170.925 ;
        RECT 41.695 170.865 41.885 171.305 ;
        RECT 42.055 170.855 43.005 171.135 ;
        RECT 43.225 170.945 43.575 171.115 ;
        RECT 41.355 170.525 41.885 170.695 ;
        RECT 39.860 170.065 40.600 170.095 ;
        RECT 39.480 169.065 39.735 169.945 ;
        RECT 39.905 168.755 40.210 169.895 ;
        RECT 40.430 169.475 40.600 170.065 ;
        RECT 40.945 169.985 41.485 170.355 ;
        RECT 41.665 170.245 41.885 170.525 ;
        RECT 42.055 170.075 42.225 170.855 ;
        RECT 41.820 169.905 42.225 170.075 ;
        RECT 42.395 170.065 42.745 170.685 ;
        RECT 41.820 169.815 41.990 169.905 ;
        RECT 42.915 169.895 43.125 170.685 ;
        RECT 40.770 169.645 41.990 169.815 ;
        RECT 42.450 169.735 43.125 169.895 ;
        RECT 40.430 169.305 41.230 169.475 ;
        RECT 40.550 168.755 40.880 169.135 ;
        RECT 41.060 169.015 41.230 169.305 ;
        RECT 41.820 169.265 41.990 169.645 ;
        RECT 42.160 169.725 43.125 169.735 ;
        RECT 43.315 170.555 43.575 170.945 ;
        RECT 43.785 170.845 44.115 171.305 ;
        RECT 44.990 170.915 45.845 171.085 ;
        RECT 46.050 170.915 46.545 171.085 ;
        RECT 46.715 170.945 47.045 171.305 ;
        RECT 43.315 169.865 43.485 170.555 ;
        RECT 43.655 170.205 43.825 170.385 ;
        RECT 43.995 170.375 44.785 170.625 ;
        RECT 44.990 170.205 45.160 170.915 ;
        RECT 45.330 170.405 45.685 170.625 ;
        RECT 43.655 170.035 45.345 170.205 ;
        RECT 42.160 169.435 42.620 169.725 ;
        RECT 43.315 169.695 44.815 169.865 ;
        RECT 43.315 169.555 43.485 169.695 ;
        RECT 42.925 169.385 43.485 169.555 ;
        RECT 41.400 168.755 41.650 169.215 ;
        RECT 41.820 168.925 42.690 169.265 ;
        RECT 42.925 168.925 43.095 169.385 ;
        RECT 43.930 169.355 45.005 169.525 ;
        RECT 43.265 168.755 43.635 169.215 ;
        RECT 43.930 169.015 44.100 169.355 ;
        RECT 44.270 168.755 44.600 169.185 ;
        RECT 44.835 169.015 45.005 169.355 ;
        RECT 45.175 169.255 45.345 170.035 ;
        RECT 45.515 169.815 45.685 170.405 ;
        RECT 45.855 170.005 46.205 170.625 ;
        RECT 45.515 169.425 45.980 169.815 ;
        RECT 46.375 169.555 46.545 170.915 ;
        RECT 46.715 169.725 47.175 170.775 ;
        RECT 46.150 169.385 46.545 169.555 ;
        RECT 46.150 169.255 46.320 169.385 ;
        RECT 45.175 168.925 45.855 169.255 ;
        RECT 46.070 168.925 46.320 169.255 ;
        RECT 46.490 168.755 46.740 169.215 ;
        RECT 46.910 168.940 47.235 169.725 ;
        RECT 47.405 168.925 47.575 171.045 ;
        RECT 47.745 170.925 48.075 171.305 ;
        RECT 48.245 170.755 48.500 171.045 ;
        RECT 47.750 170.585 48.500 170.755 ;
        RECT 47.750 169.595 47.980 170.585 ;
        RECT 48.675 170.580 48.965 171.305 ;
        RECT 49.140 170.595 49.395 171.125 ;
        RECT 49.565 170.845 49.870 171.305 ;
        RECT 50.115 170.925 51.185 171.095 ;
        RECT 48.150 169.765 48.500 170.415 ;
        RECT 49.140 169.945 49.350 170.595 ;
        RECT 50.115 170.570 50.435 170.925 ;
        RECT 50.110 170.395 50.435 170.570 ;
        RECT 49.520 170.095 50.435 170.395 ;
        RECT 50.605 170.355 50.845 170.755 ;
        RECT 51.015 170.695 51.185 170.925 ;
        RECT 51.355 170.865 51.545 171.305 ;
        RECT 51.715 170.855 52.665 171.135 ;
        RECT 52.885 170.945 53.235 171.115 ;
        RECT 51.015 170.525 51.545 170.695 ;
        RECT 49.520 170.065 50.260 170.095 ;
        RECT 47.750 169.425 48.500 169.595 ;
        RECT 47.745 168.755 48.075 169.255 ;
        RECT 48.245 168.925 48.500 169.425 ;
        RECT 48.675 168.755 48.965 169.920 ;
        RECT 49.140 169.065 49.395 169.945 ;
        RECT 49.565 168.755 49.870 169.895 ;
        RECT 50.090 169.475 50.260 170.065 ;
        RECT 50.605 169.985 51.145 170.355 ;
        RECT 51.325 170.245 51.545 170.525 ;
        RECT 51.715 170.075 51.885 170.855 ;
        RECT 51.480 169.905 51.885 170.075 ;
        RECT 52.055 170.065 52.405 170.685 ;
        RECT 51.480 169.815 51.650 169.905 ;
        RECT 52.575 169.895 52.785 170.685 ;
        RECT 50.430 169.645 51.650 169.815 ;
        RECT 52.110 169.735 52.785 169.895 ;
        RECT 50.090 169.305 50.890 169.475 ;
        RECT 50.210 168.755 50.540 169.135 ;
        RECT 50.720 169.015 50.890 169.305 ;
        RECT 51.480 169.265 51.650 169.645 ;
        RECT 51.820 169.725 52.785 169.735 ;
        RECT 52.975 170.555 53.235 170.945 ;
        RECT 53.445 170.845 53.775 171.305 ;
        RECT 54.650 170.915 55.505 171.085 ;
        RECT 55.710 170.915 56.205 171.085 ;
        RECT 56.375 170.945 56.705 171.305 ;
        RECT 52.975 169.865 53.145 170.555 ;
        RECT 53.315 170.205 53.485 170.385 ;
        RECT 53.655 170.375 54.445 170.625 ;
        RECT 54.650 170.205 54.820 170.915 ;
        RECT 54.990 170.405 55.345 170.625 ;
        RECT 53.315 170.035 55.005 170.205 ;
        RECT 51.820 169.435 52.280 169.725 ;
        RECT 52.975 169.695 54.475 169.865 ;
        RECT 52.975 169.555 53.145 169.695 ;
        RECT 52.585 169.385 53.145 169.555 ;
        RECT 51.060 168.755 51.310 169.215 ;
        RECT 51.480 168.925 52.350 169.265 ;
        RECT 52.585 168.925 52.755 169.385 ;
        RECT 53.590 169.355 54.665 169.525 ;
        RECT 52.925 168.755 53.295 169.215 ;
        RECT 53.590 169.015 53.760 169.355 ;
        RECT 53.930 168.755 54.260 169.185 ;
        RECT 54.495 169.015 54.665 169.355 ;
        RECT 54.835 169.255 55.005 170.035 ;
        RECT 55.175 169.815 55.345 170.405 ;
        RECT 55.515 170.005 55.865 170.625 ;
        RECT 55.175 169.425 55.640 169.815 ;
        RECT 56.035 169.555 56.205 170.915 ;
        RECT 56.375 169.725 56.835 170.775 ;
        RECT 55.810 169.385 56.205 169.555 ;
        RECT 55.810 169.255 55.980 169.385 ;
        RECT 54.835 168.925 55.515 169.255 ;
        RECT 55.730 168.925 55.980 169.255 ;
        RECT 56.150 168.755 56.400 169.215 ;
        RECT 56.570 168.940 56.895 169.725 ;
        RECT 57.065 168.925 57.235 171.045 ;
        RECT 57.405 170.925 57.735 171.305 ;
        RECT 57.905 170.755 58.160 171.045 ;
        RECT 57.410 170.585 58.160 170.755 ;
        RECT 59.345 170.755 59.515 171.135 ;
        RECT 59.695 170.925 60.025 171.305 ;
        RECT 59.345 170.585 60.010 170.755 ;
        RECT 60.205 170.630 60.465 171.135 ;
        RECT 60.695 170.825 60.975 171.305 ;
        RECT 61.145 170.655 61.405 171.045 ;
        RECT 61.580 170.825 61.835 171.305 ;
        RECT 62.005 170.655 62.300 171.045 ;
        RECT 62.480 170.825 62.755 171.305 ;
        RECT 62.925 170.805 63.225 171.135 ;
        RECT 57.410 169.595 57.640 170.585 ;
        RECT 57.810 169.765 58.160 170.415 ;
        RECT 59.275 170.035 59.605 170.405 ;
        RECT 59.840 170.330 60.010 170.585 ;
        RECT 59.840 170.000 60.125 170.330 ;
        RECT 59.840 169.855 60.010 170.000 ;
        RECT 59.345 169.685 60.010 169.855 ;
        RECT 60.295 169.830 60.465 170.630 ;
        RECT 57.410 169.425 58.160 169.595 ;
        RECT 57.405 168.755 57.735 169.255 ;
        RECT 57.905 168.925 58.160 169.425 ;
        RECT 59.345 168.925 59.515 169.685 ;
        RECT 59.695 168.755 60.025 169.515 ;
        RECT 60.195 168.925 60.465 169.830 ;
        RECT 60.650 170.485 62.300 170.655 ;
        RECT 60.650 169.975 61.055 170.485 ;
        RECT 61.225 170.145 62.365 170.315 ;
        RECT 60.650 169.805 61.405 169.975 ;
        RECT 60.690 168.755 60.975 169.625 ;
        RECT 61.145 169.555 61.405 169.805 ;
        RECT 62.195 169.895 62.365 170.145 ;
        RECT 62.535 170.065 62.885 170.635 ;
        RECT 63.055 169.895 63.225 170.805 ;
        RECT 63.545 170.505 63.875 171.305 ;
        RECT 64.045 170.655 64.215 171.135 ;
        RECT 64.385 170.825 64.715 171.305 ;
        RECT 64.885 170.655 65.055 171.135 ;
        RECT 65.305 170.825 65.545 171.305 ;
        RECT 65.725 170.655 65.895 171.135 ;
        RECT 64.045 170.485 65.055 170.655 ;
        RECT 65.260 170.485 65.895 170.655 ;
        RECT 67.225 170.505 67.555 171.305 ;
        RECT 67.725 170.655 67.895 171.135 ;
        RECT 68.065 170.825 68.395 171.305 ;
        RECT 68.565 170.655 68.735 171.135 ;
        RECT 68.985 170.825 69.225 171.305 ;
        RECT 69.405 170.655 69.575 171.135 ;
        RECT 67.725 170.485 68.735 170.655 ;
        RECT 68.940 170.485 69.575 170.655 ;
        RECT 70.570 170.495 70.815 171.100 ;
        RECT 71.035 170.770 71.545 171.305 ;
        RECT 64.045 170.285 64.540 170.485 ;
        RECT 65.260 170.315 65.430 170.485 ;
        RECT 64.045 170.115 64.545 170.285 ;
        RECT 64.930 170.145 65.430 170.315 ;
        RECT 64.045 169.945 64.540 170.115 ;
        RECT 62.195 169.725 63.225 169.895 ;
        RECT 61.145 169.385 62.265 169.555 ;
        RECT 61.145 168.925 61.405 169.385 ;
        RECT 61.580 168.755 61.835 169.215 ;
        RECT 62.005 168.925 62.265 169.385 ;
        RECT 62.435 168.755 62.745 169.555 ;
        RECT 62.915 168.925 63.225 169.725 ;
        RECT 63.545 168.755 63.875 169.905 ;
        RECT 64.045 169.775 65.055 169.945 ;
        RECT 64.045 168.925 64.215 169.775 ;
        RECT 64.385 168.755 64.715 169.555 ;
        RECT 64.885 168.925 65.055 169.775 ;
        RECT 65.260 169.905 65.430 170.145 ;
        RECT 65.600 170.075 65.980 170.315 ;
        RECT 67.725 169.945 68.220 170.485 ;
        RECT 68.940 170.315 69.110 170.485 ;
        RECT 70.295 170.325 71.525 170.495 ;
        RECT 68.610 170.145 69.110 170.315 ;
        RECT 65.260 169.735 65.975 169.905 ;
        RECT 65.235 168.755 65.475 169.555 ;
        RECT 65.645 168.925 65.975 169.735 ;
        RECT 67.225 168.755 67.555 169.905 ;
        RECT 67.725 169.775 68.735 169.945 ;
        RECT 67.725 168.925 67.895 169.775 ;
        RECT 68.065 168.755 68.395 169.555 ;
        RECT 68.565 168.925 68.735 169.775 ;
        RECT 68.940 169.905 69.110 170.145 ;
        RECT 69.280 170.075 69.660 170.315 ;
        RECT 68.940 169.735 69.655 169.905 ;
        RECT 68.915 168.755 69.155 169.555 ;
        RECT 69.325 168.925 69.655 169.735 ;
        RECT 70.295 169.515 70.635 170.325 ;
        RECT 70.805 169.760 71.555 169.950 ;
        RECT 70.295 169.105 70.810 169.515 ;
        RECT 71.045 168.755 71.215 169.515 ;
        RECT 71.385 169.095 71.555 169.760 ;
        RECT 71.725 169.775 71.915 171.135 ;
        RECT 72.085 170.285 72.360 171.135 ;
        RECT 72.550 170.770 73.080 171.135 ;
        RECT 73.505 170.905 73.835 171.305 ;
        RECT 72.905 170.735 73.080 170.770 ;
        RECT 72.085 170.115 72.365 170.285 ;
        RECT 72.085 169.975 72.360 170.115 ;
        RECT 72.565 169.775 72.735 170.575 ;
        RECT 71.725 169.605 72.735 169.775 ;
        RECT 72.905 170.565 73.835 170.735 ;
        RECT 74.005 170.565 74.260 171.135 ;
        RECT 74.435 170.580 74.725 171.305 ;
        RECT 75.270 170.595 75.525 171.125 ;
        RECT 75.705 170.845 75.990 171.305 ;
        RECT 72.905 169.435 73.075 170.565 ;
        RECT 73.665 170.395 73.835 170.565 ;
        RECT 71.950 169.265 73.075 169.435 ;
        RECT 73.245 170.065 73.440 170.395 ;
        RECT 73.665 170.065 73.920 170.395 ;
        RECT 73.245 169.095 73.415 170.065 ;
        RECT 74.090 169.895 74.260 170.565 ;
        RECT 71.385 168.925 73.415 169.095 ;
        RECT 73.585 168.755 73.755 169.895 ;
        RECT 73.925 168.925 74.260 169.895 ;
        RECT 74.435 168.755 74.725 169.920 ;
        RECT 75.270 169.735 75.450 170.595 ;
        RECT 76.170 170.395 76.420 171.045 ;
        RECT 75.620 170.065 76.420 170.395 ;
        RECT 75.270 169.265 75.525 169.735 ;
        RECT 75.185 169.095 75.525 169.265 ;
        RECT 75.270 169.065 75.525 169.095 ;
        RECT 75.705 168.755 75.990 169.555 ;
        RECT 76.170 169.475 76.420 170.065 ;
        RECT 76.620 170.710 76.940 171.040 ;
        RECT 77.120 170.825 77.780 171.305 ;
        RECT 77.980 170.915 78.830 171.085 ;
        RECT 76.620 169.815 76.810 170.710 ;
        RECT 77.130 170.385 77.790 170.655 ;
        RECT 77.460 170.325 77.790 170.385 ;
        RECT 76.980 170.155 77.310 170.215 ;
        RECT 77.980 170.155 78.150 170.915 ;
        RECT 79.390 170.845 79.710 171.305 ;
        RECT 79.910 170.665 80.160 171.095 ;
        RECT 80.450 170.865 80.860 171.305 ;
        RECT 81.030 170.925 82.045 171.125 ;
        RECT 78.320 170.495 79.570 170.665 ;
        RECT 78.320 170.375 78.650 170.495 ;
        RECT 76.980 169.985 78.880 170.155 ;
        RECT 76.620 169.645 78.540 169.815 ;
        RECT 76.620 169.625 76.940 169.645 ;
        RECT 76.170 168.965 76.500 169.475 ;
        RECT 76.770 169.015 76.940 169.625 ;
        RECT 78.710 169.475 78.880 169.985 ;
        RECT 79.050 169.915 79.230 170.325 ;
        RECT 79.400 169.735 79.570 170.495 ;
        RECT 77.110 168.755 77.440 169.445 ;
        RECT 77.670 169.305 78.880 169.475 ;
        RECT 79.050 169.425 79.570 169.735 ;
        RECT 79.740 170.325 80.160 170.665 ;
        RECT 80.450 170.325 80.860 170.655 ;
        RECT 79.740 169.555 79.930 170.325 ;
        RECT 81.030 170.195 81.200 170.925 ;
        RECT 82.345 170.755 82.515 171.085 ;
        RECT 82.685 170.925 83.015 171.305 ;
        RECT 81.370 170.375 81.720 170.745 ;
        RECT 81.030 170.155 81.450 170.195 ;
        RECT 80.100 169.985 81.450 170.155 ;
        RECT 80.100 169.825 80.350 169.985 ;
        RECT 80.860 169.555 81.110 169.815 ;
        RECT 79.740 169.305 81.110 169.555 ;
        RECT 77.670 169.015 77.910 169.305 ;
        RECT 78.710 169.225 78.880 169.305 ;
        RECT 78.110 168.755 78.530 169.135 ;
        RECT 78.710 168.975 79.340 169.225 ;
        RECT 79.810 168.755 80.140 169.135 ;
        RECT 80.310 169.015 80.480 169.305 ;
        RECT 81.280 169.140 81.450 169.985 ;
        RECT 81.900 169.815 82.120 170.685 ;
        RECT 82.345 170.565 83.040 170.755 ;
        RECT 81.620 169.435 82.120 169.815 ;
        RECT 82.290 169.765 82.700 170.385 ;
        RECT 82.870 169.595 83.040 170.565 ;
        RECT 82.345 169.425 83.040 169.595 ;
        RECT 80.660 168.755 81.040 169.135 ;
        RECT 81.280 168.970 82.110 169.140 ;
        RECT 82.345 168.925 82.515 169.425 ;
        RECT 82.685 168.755 83.015 169.255 ;
        RECT 83.230 168.925 83.455 171.045 ;
        RECT 83.625 170.925 83.955 171.305 ;
        RECT 84.125 170.755 84.295 171.045 ;
        RECT 85.105 170.825 85.405 171.305 ;
        RECT 83.630 170.585 84.295 170.755 ;
        RECT 85.575 170.655 85.835 171.110 ;
        RECT 86.005 170.825 86.265 171.305 ;
        RECT 86.445 170.655 86.705 171.110 ;
        RECT 86.875 170.825 87.125 171.305 ;
        RECT 87.305 170.655 87.565 171.110 ;
        RECT 87.735 170.825 87.985 171.305 ;
        RECT 88.165 170.655 88.425 171.110 ;
        RECT 88.595 170.825 88.840 171.305 ;
        RECT 89.010 170.655 89.285 171.110 ;
        RECT 89.455 170.825 89.700 171.305 ;
        RECT 89.870 170.655 90.130 171.110 ;
        RECT 90.300 170.825 90.560 171.305 ;
        RECT 90.730 170.655 90.990 171.110 ;
        RECT 91.160 170.825 91.420 171.305 ;
        RECT 91.590 170.655 91.850 171.110 ;
        RECT 92.020 170.745 92.280 171.305 ;
        RECT 83.630 169.595 83.860 170.585 ;
        RECT 85.105 170.485 91.850 170.655 ;
        RECT 84.030 169.765 84.380 170.415 ;
        RECT 85.105 169.895 86.270 170.485 ;
        RECT 92.450 170.315 92.700 171.125 ;
        RECT 92.880 170.780 93.140 171.305 ;
        RECT 93.310 170.315 93.560 171.125 ;
        RECT 93.740 170.795 94.045 171.305 ;
        RECT 86.440 170.065 93.560 170.315 ;
        RECT 93.730 170.065 94.045 170.625 ;
        RECT 94.490 170.495 94.735 171.100 ;
        RECT 94.955 170.770 95.465 171.305 ;
        RECT 94.215 170.325 95.445 170.495 ;
        RECT 85.105 169.670 91.850 169.895 ;
        RECT 83.630 169.425 84.295 169.595 ;
        RECT 83.625 168.755 83.955 169.255 ;
        RECT 84.125 168.925 84.295 169.425 ;
        RECT 85.105 168.755 85.375 169.500 ;
        RECT 85.545 168.930 85.835 169.670 ;
        RECT 86.445 169.655 91.850 169.670 ;
        RECT 86.005 168.760 86.260 169.485 ;
        RECT 86.445 168.930 86.705 169.655 ;
        RECT 86.875 168.760 87.120 169.485 ;
        RECT 87.305 168.930 87.565 169.655 ;
        RECT 87.735 168.760 87.980 169.485 ;
        RECT 88.165 168.930 88.425 169.655 ;
        RECT 88.595 168.760 88.840 169.485 ;
        RECT 89.010 168.930 89.270 169.655 ;
        RECT 89.440 168.760 89.700 169.485 ;
        RECT 89.870 168.930 90.130 169.655 ;
        RECT 90.300 168.760 90.560 169.485 ;
        RECT 90.730 168.930 90.990 169.655 ;
        RECT 91.160 168.760 91.420 169.485 ;
        RECT 91.590 168.930 91.850 169.655 ;
        RECT 92.020 168.760 92.280 169.555 ;
        RECT 92.450 168.930 92.700 170.065 ;
        RECT 86.005 168.755 92.280 168.760 ;
        RECT 92.880 168.755 93.140 169.565 ;
        RECT 93.315 168.925 93.560 170.065 ;
        RECT 93.740 168.755 94.035 169.565 ;
        RECT 94.215 169.515 94.555 170.325 ;
        RECT 94.725 169.760 95.475 169.950 ;
        RECT 94.215 169.105 94.730 169.515 ;
        RECT 94.965 168.755 95.135 169.515 ;
        RECT 95.305 169.095 95.475 169.760 ;
        RECT 95.645 169.775 95.835 171.135 ;
        RECT 96.005 170.965 96.280 171.135 ;
        RECT 96.005 170.795 96.285 170.965 ;
        RECT 96.005 169.975 96.280 170.795 ;
        RECT 96.470 170.770 97.000 171.135 ;
        RECT 97.425 170.905 97.755 171.305 ;
        RECT 96.825 170.735 97.000 170.770 ;
        RECT 96.485 169.775 96.655 170.575 ;
        RECT 95.645 169.605 96.655 169.775 ;
        RECT 96.825 170.565 97.755 170.735 ;
        RECT 97.925 170.565 98.180 171.135 ;
        RECT 98.360 170.905 98.695 171.305 ;
        RECT 98.865 170.735 99.070 171.135 ;
        RECT 99.280 170.825 99.555 171.305 ;
        RECT 99.765 170.805 100.025 171.135 ;
        RECT 96.825 169.435 96.995 170.565 ;
        RECT 97.585 170.395 97.755 170.565 ;
        RECT 95.870 169.265 96.995 169.435 ;
        RECT 97.165 170.065 97.360 170.395 ;
        RECT 97.585 170.065 97.840 170.395 ;
        RECT 97.165 169.095 97.335 170.065 ;
        RECT 98.010 169.895 98.180 170.565 ;
        RECT 95.305 168.925 97.335 169.095 ;
        RECT 97.505 168.755 97.675 169.895 ;
        RECT 97.845 168.925 98.180 169.895 ;
        RECT 98.385 170.565 99.070 170.735 ;
        RECT 98.385 169.535 98.725 170.565 ;
        RECT 98.895 169.895 99.145 170.395 ;
        RECT 99.325 170.065 99.685 170.645 ;
        RECT 99.855 169.895 100.025 170.805 ;
        RECT 100.195 170.580 100.485 171.305 ;
        RECT 100.660 170.565 100.915 171.135 ;
        RECT 101.085 170.905 101.415 171.305 ;
        RECT 101.840 170.770 102.370 171.135 ;
        RECT 101.840 170.735 102.015 170.770 ;
        RECT 101.085 170.565 102.015 170.735 ;
        RECT 98.895 169.725 100.025 169.895 ;
        RECT 98.385 169.360 99.050 169.535 ;
        RECT 98.360 168.755 98.695 169.180 ;
        RECT 98.865 168.955 99.050 169.360 ;
        RECT 99.255 168.755 99.585 169.535 ;
        RECT 99.755 168.955 100.025 169.725 ;
        RECT 100.195 168.755 100.485 169.920 ;
        RECT 100.660 169.895 100.830 170.565 ;
        RECT 101.085 170.395 101.255 170.565 ;
        RECT 101.000 170.065 101.255 170.395 ;
        RECT 101.480 170.065 101.675 170.395 ;
        RECT 100.660 168.925 100.995 169.895 ;
        RECT 101.165 168.755 101.335 169.895 ;
        RECT 101.505 169.095 101.675 170.065 ;
        RECT 101.845 169.435 102.015 170.565 ;
        RECT 102.185 169.775 102.355 170.575 ;
        RECT 102.560 170.285 102.835 171.135 ;
        RECT 102.555 170.115 102.835 170.285 ;
        RECT 102.560 169.975 102.835 170.115 ;
        RECT 103.005 169.775 103.195 171.135 ;
        RECT 103.375 170.770 103.885 171.305 ;
        RECT 104.105 170.495 104.350 171.100 ;
        RECT 104.795 170.565 105.180 171.135 ;
        RECT 105.350 170.845 105.675 171.305 ;
        RECT 106.195 170.675 106.475 171.135 ;
        RECT 103.395 170.325 104.625 170.495 ;
        RECT 102.185 169.605 103.195 169.775 ;
        RECT 103.365 169.760 104.115 169.950 ;
        RECT 101.845 169.265 102.970 169.435 ;
        RECT 103.365 169.095 103.535 169.760 ;
        RECT 104.285 169.515 104.625 170.325 ;
        RECT 101.505 168.925 103.535 169.095 ;
        RECT 103.705 168.755 103.875 169.515 ;
        RECT 104.110 169.105 104.625 169.515 ;
        RECT 104.795 169.895 105.075 170.565 ;
        RECT 105.350 170.505 106.475 170.675 ;
        RECT 105.350 170.395 105.800 170.505 ;
        RECT 105.245 170.065 105.800 170.395 ;
        RECT 106.665 170.335 107.065 171.135 ;
        RECT 107.465 170.845 107.735 171.305 ;
        RECT 107.905 170.675 108.190 171.135 ;
        RECT 108.575 170.840 108.825 171.305 ;
        RECT 104.795 168.925 105.180 169.895 ;
        RECT 105.350 169.605 105.800 170.065 ;
        RECT 105.970 169.775 107.065 170.335 ;
        RECT 105.350 169.385 106.475 169.605 ;
        RECT 105.350 168.755 105.675 169.215 ;
        RECT 106.195 168.925 106.475 169.385 ;
        RECT 106.665 168.925 107.065 169.775 ;
        RECT 107.235 170.505 108.190 170.675 ;
        RECT 108.995 170.665 109.165 171.135 ;
        RECT 109.415 170.845 109.585 171.305 ;
        RECT 109.835 170.665 110.005 171.135 ;
        RECT 110.255 170.845 110.425 171.305 ;
        RECT 110.675 170.665 110.845 171.135 ;
        RECT 111.215 170.845 111.480 171.305 ;
        RECT 107.235 169.605 107.445 170.505 ;
        RECT 108.475 170.485 110.845 170.665 ;
        RECT 112.155 170.555 113.365 171.305 ;
        RECT 107.615 169.775 108.305 170.335 ;
        RECT 108.475 169.895 108.825 170.485 ;
        RECT 108.995 170.065 111.505 170.315 ;
        RECT 108.475 169.725 110.925 169.895 ;
        RECT 108.475 169.705 109.245 169.725 ;
        RECT 107.235 169.385 108.190 169.605 ;
        RECT 107.465 168.755 107.735 169.215 ;
        RECT 107.905 168.925 108.190 169.385 ;
        RECT 108.575 168.755 108.745 169.215 ;
        RECT 108.915 168.925 109.245 169.705 ;
        RECT 109.415 168.755 109.585 169.555 ;
        RECT 109.755 168.925 110.085 169.725 ;
        RECT 110.255 168.755 110.425 169.555 ;
        RECT 110.595 168.925 110.925 169.725 ;
        RECT 111.185 168.755 111.480 169.895 ;
        RECT 112.155 169.845 112.675 170.385 ;
        RECT 112.845 170.015 113.365 170.555 ;
        RECT 112.155 168.755 113.365 169.845 ;
        RECT 22.830 168.585 113.450 168.755 ;
        RECT 22.915 167.495 24.125 168.585 ;
        RECT 22.915 166.785 23.435 167.325 ;
        RECT 23.605 166.955 24.125 167.495 ;
        RECT 24.300 167.445 24.635 168.415 ;
        RECT 24.805 167.445 24.975 168.585 ;
        RECT 25.145 168.245 27.175 168.415 ;
        RECT 22.915 166.035 24.125 166.785 ;
        RECT 24.300 166.775 24.470 167.445 ;
        RECT 25.145 167.275 25.315 168.245 ;
        RECT 24.640 166.945 24.895 167.275 ;
        RECT 25.120 166.945 25.315 167.275 ;
        RECT 25.485 167.905 26.610 168.075 ;
        RECT 24.725 166.775 24.895 166.945 ;
        RECT 25.485 166.775 25.655 167.905 ;
        RECT 24.300 166.205 24.555 166.775 ;
        RECT 24.725 166.605 25.655 166.775 ;
        RECT 25.825 167.565 26.835 167.735 ;
        RECT 25.825 166.765 25.995 167.565 ;
        RECT 26.200 167.225 26.475 167.365 ;
        RECT 26.195 167.055 26.475 167.225 ;
        RECT 25.480 166.570 25.655 166.605 ;
        RECT 24.725 166.035 25.055 166.435 ;
        RECT 25.480 166.205 26.010 166.570 ;
        RECT 26.200 166.205 26.475 167.055 ;
        RECT 26.645 166.205 26.835 167.565 ;
        RECT 27.005 167.580 27.175 168.245 ;
        RECT 27.345 167.825 27.515 168.585 ;
        RECT 27.750 167.825 28.265 168.235 ;
        RECT 27.005 167.390 27.755 167.580 ;
        RECT 27.925 167.015 28.265 167.825 ;
        RECT 27.035 166.845 28.265 167.015 ;
        RECT 28.435 167.825 28.950 168.235 ;
        RECT 29.185 167.825 29.355 168.585 ;
        RECT 29.525 168.245 31.555 168.415 ;
        RECT 28.435 167.015 28.775 167.825 ;
        RECT 29.525 167.580 29.695 168.245 ;
        RECT 30.090 167.905 31.215 168.075 ;
        RECT 28.945 167.390 29.695 167.580 ;
        RECT 29.865 167.565 30.875 167.735 ;
        RECT 28.435 166.845 29.665 167.015 ;
        RECT 27.015 166.035 27.525 166.570 ;
        RECT 27.745 166.240 27.990 166.845 ;
        RECT 28.710 166.240 28.955 166.845 ;
        RECT 29.175 166.035 29.685 166.570 ;
        RECT 29.865 166.205 30.055 167.565 ;
        RECT 30.225 166.545 30.500 167.365 ;
        RECT 30.705 166.765 30.875 167.565 ;
        RECT 31.045 166.775 31.215 167.905 ;
        RECT 31.385 167.275 31.555 168.245 ;
        RECT 31.725 167.445 31.895 168.585 ;
        RECT 32.065 167.445 32.400 168.415 ;
        RECT 32.575 167.750 32.960 168.585 ;
        RECT 33.130 167.580 33.390 168.385 ;
        RECT 33.560 167.750 33.820 168.585 ;
        RECT 33.990 167.580 34.245 168.385 ;
        RECT 34.420 167.750 34.680 168.585 ;
        RECT 34.850 167.580 35.105 168.385 ;
        RECT 35.280 167.750 35.625 168.585 ;
        RECT 31.385 166.945 31.580 167.275 ;
        RECT 31.805 166.945 32.060 167.275 ;
        RECT 31.805 166.775 31.975 166.945 ;
        RECT 32.230 166.775 32.400 167.445 ;
        RECT 31.045 166.605 31.975 166.775 ;
        RECT 31.045 166.570 31.220 166.605 ;
        RECT 30.225 166.375 30.505 166.545 ;
        RECT 30.225 166.205 30.500 166.375 ;
        RECT 30.690 166.205 31.220 166.570 ;
        RECT 31.645 166.035 31.975 166.435 ;
        RECT 32.145 166.205 32.400 166.775 ;
        RECT 32.575 167.410 35.605 167.580 ;
        RECT 35.795 167.420 36.085 168.585 ;
        RECT 36.255 167.825 36.770 168.235 ;
        RECT 37.005 167.825 37.175 168.585 ;
        RECT 37.345 168.245 39.375 168.415 ;
        RECT 32.575 166.845 32.875 167.410 ;
        RECT 33.050 167.015 35.265 167.240 ;
        RECT 35.435 166.845 35.605 167.410 ;
        RECT 36.255 167.015 36.595 167.825 ;
        RECT 37.345 167.580 37.515 168.245 ;
        RECT 37.910 167.905 39.035 168.075 ;
        RECT 36.765 167.390 37.515 167.580 ;
        RECT 37.685 167.565 38.695 167.735 ;
        RECT 36.255 166.845 37.485 167.015 ;
        RECT 32.575 166.675 35.605 166.845 ;
        RECT 33.095 166.035 33.395 166.505 ;
        RECT 33.565 166.230 33.820 166.675 ;
        RECT 33.990 166.035 34.250 166.505 ;
        RECT 34.420 166.230 34.680 166.675 ;
        RECT 34.850 166.035 35.145 166.505 ;
        RECT 35.795 166.035 36.085 166.760 ;
        RECT 36.530 166.240 36.775 166.845 ;
        RECT 36.995 166.035 37.505 166.570 ;
        RECT 37.685 166.205 37.875 167.565 ;
        RECT 38.045 166.885 38.320 167.365 ;
        RECT 38.045 166.715 38.325 166.885 ;
        RECT 38.525 166.765 38.695 167.565 ;
        RECT 38.865 166.775 39.035 167.905 ;
        RECT 39.205 167.275 39.375 168.245 ;
        RECT 39.545 167.445 39.715 168.585 ;
        RECT 39.885 167.445 40.220 168.415 ;
        RECT 40.435 167.445 40.665 168.585 ;
        RECT 39.205 166.945 39.400 167.275 ;
        RECT 39.625 166.945 39.880 167.275 ;
        RECT 39.625 166.775 39.795 166.945 ;
        RECT 40.050 166.775 40.220 167.445 ;
        RECT 40.835 167.435 41.165 168.415 ;
        RECT 41.335 167.445 41.545 168.585 ;
        RECT 41.890 167.955 42.175 168.415 ;
        RECT 42.345 168.125 42.615 168.585 ;
        RECT 41.890 167.735 42.845 167.955 ;
        RECT 40.415 167.025 40.745 167.275 ;
        RECT 38.045 166.205 38.320 166.715 ;
        RECT 38.865 166.605 39.795 166.775 ;
        RECT 38.865 166.570 39.040 166.605 ;
        RECT 38.510 166.205 39.040 166.570 ;
        RECT 39.465 166.035 39.795 166.435 ;
        RECT 39.965 166.205 40.220 166.775 ;
        RECT 40.435 166.035 40.665 166.855 ;
        RECT 40.915 166.835 41.165 167.435 ;
        RECT 41.775 167.005 42.465 167.565 ;
        RECT 40.835 166.205 41.165 166.835 ;
        RECT 41.335 166.035 41.545 166.855 ;
        RECT 42.635 166.835 42.845 167.735 ;
        RECT 41.890 166.665 42.845 166.835 ;
        RECT 43.015 167.565 43.415 168.415 ;
        RECT 43.605 167.955 43.885 168.415 ;
        RECT 44.405 168.125 44.730 168.585 ;
        RECT 43.605 167.735 44.730 167.955 ;
        RECT 43.015 167.005 44.110 167.565 ;
        RECT 44.280 167.275 44.730 167.735 ;
        RECT 44.900 167.445 45.285 168.415 ;
        RECT 41.890 166.205 42.175 166.665 ;
        RECT 42.345 166.035 42.615 166.495 ;
        RECT 43.015 166.205 43.415 167.005 ;
        RECT 44.280 166.945 44.835 167.275 ;
        RECT 44.280 166.835 44.730 166.945 ;
        RECT 43.605 166.665 44.730 166.835 ;
        RECT 45.005 166.775 45.285 167.445 ;
        RECT 45.455 167.825 45.970 168.235 ;
        RECT 46.205 167.825 46.375 168.585 ;
        RECT 46.545 168.245 48.575 168.415 ;
        RECT 45.455 167.015 45.795 167.825 ;
        RECT 46.545 167.580 46.715 168.245 ;
        RECT 47.110 167.905 48.235 168.075 ;
        RECT 45.965 167.390 46.715 167.580 ;
        RECT 46.885 167.565 47.895 167.735 ;
        RECT 45.455 166.845 46.685 167.015 ;
        RECT 43.605 166.205 43.885 166.665 ;
        RECT 44.405 166.035 44.730 166.495 ;
        RECT 44.900 166.205 45.285 166.775 ;
        RECT 45.730 166.240 45.975 166.845 ;
        RECT 46.195 166.035 46.705 166.570 ;
        RECT 46.885 166.205 47.075 167.565 ;
        RECT 47.245 167.225 47.520 167.365 ;
        RECT 47.245 167.055 47.525 167.225 ;
        RECT 47.245 166.205 47.520 167.055 ;
        RECT 47.725 166.765 47.895 167.565 ;
        RECT 48.065 166.775 48.235 167.905 ;
        RECT 48.405 167.275 48.575 168.245 ;
        RECT 48.745 167.445 48.915 168.585 ;
        RECT 49.085 167.445 49.420 168.415 ;
        RECT 49.685 167.655 49.855 168.415 ;
        RECT 50.035 167.825 50.365 168.585 ;
        RECT 49.685 167.485 50.350 167.655 ;
        RECT 50.535 167.510 50.805 168.415 ;
        RECT 48.405 166.945 48.600 167.275 ;
        RECT 48.825 166.945 49.080 167.275 ;
        RECT 48.825 166.775 48.995 166.945 ;
        RECT 49.250 166.775 49.420 167.445 ;
        RECT 50.180 167.340 50.350 167.485 ;
        RECT 49.615 166.935 49.945 167.305 ;
        RECT 50.180 167.010 50.465 167.340 ;
        RECT 48.065 166.605 48.995 166.775 ;
        RECT 48.065 166.570 48.240 166.605 ;
        RECT 47.710 166.205 48.240 166.570 ;
        RECT 48.665 166.035 48.995 166.435 ;
        RECT 49.165 166.205 49.420 166.775 ;
        RECT 50.180 166.755 50.350 167.010 ;
        RECT 49.685 166.585 50.350 166.755 ;
        RECT 50.635 166.710 50.805 167.510 ;
        RECT 51.015 167.445 51.245 168.585 ;
        RECT 51.415 167.435 51.745 168.415 ;
        RECT 51.915 167.445 52.125 168.585 ;
        RECT 50.995 167.025 51.325 167.275 ;
        RECT 49.685 166.205 49.855 166.585 ;
        RECT 50.035 166.035 50.365 166.415 ;
        RECT 50.545 166.205 50.805 166.710 ;
        RECT 51.015 166.035 51.245 166.855 ;
        RECT 51.495 166.835 51.745 167.435 ;
        RECT 52.360 167.395 52.615 168.275 ;
        RECT 52.785 167.445 53.090 168.585 ;
        RECT 53.430 168.205 53.760 168.585 ;
        RECT 53.940 168.035 54.110 168.325 ;
        RECT 54.280 168.125 54.530 168.585 ;
        RECT 53.310 167.865 54.110 168.035 ;
        RECT 54.700 168.075 55.570 168.415 ;
        RECT 51.415 166.205 51.745 166.835 ;
        RECT 51.915 166.035 52.125 166.855 ;
        RECT 52.360 166.745 52.570 167.395 ;
        RECT 53.310 167.275 53.480 167.865 ;
        RECT 54.700 167.695 54.870 168.075 ;
        RECT 55.805 167.955 55.975 168.415 ;
        RECT 56.145 168.125 56.515 168.585 ;
        RECT 56.810 167.985 56.980 168.325 ;
        RECT 57.150 168.155 57.480 168.585 ;
        RECT 57.715 167.985 57.885 168.325 ;
        RECT 53.650 167.525 54.870 167.695 ;
        RECT 55.040 167.615 55.500 167.905 ;
        RECT 55.805 167.785 56.365 167.955 ;
        RECT 56.810 167.815 57.885 167.985 ;
        RECT 58.055 168.085 58.735 168.415 ;
        RECT 58.950 168.085 59.200 168.415 ;
        RECT 59.370 168.125 59.620 168.585 ;
        RECT 56.195 167.645 56.365 167.785 ;
        RECT 55.040 167.605 56.005 167.615 ;
        RECT 54.700 167.435 54.870 167.525 ;
        RECT 55.330 167.445 56.005 167.605 ;
        RECT 52.740 167.245 53.480 167.275 ;
        RECT 52.740 166.945 53.655 167.245 ;
        RECT 53.330 166.770 53.655 166.945 ;
        RECT 52.360 166.215 52.615 166.745 ;
        RECT 52.785 166.035 53.090 166.495 ;
        RECT 53.335 166.415 53.655 166.770 ;
        RECT 53.825 166.985 54.365 167.355 ;
        RECT 54.700 167.265 55.105 167.435 ;
        RECT 53.825 166.585 54.065 166.985 ;
        RECT 54.545 166.815 54.765 167.095 ;
        RECT 54.235 166.645 54.765 166.815 ;
        RECT 54.235 166.415 54.405 166.645 ;
        RECT 54.935 166.485 55.105 167.265 ;
        RECT 55.275 166.655 55.625 167.275 ;
        RECT 55.795 166.655 56.005 167.445 ;
        RECT 56.195 167.475 57.695 167.645 ;
        RECT 56.195 166.785 56.365 167.475 ;
        RECT 58.055 167.305 58.225 168.085 ;
        RECT 59.030 167.955 59.200 168.085 ;
        RECT 56.535 167.135 58.225 167.305 ;
        RECT 58.395 167.525 58.860 167.915 ;
        RECT 59.030 167.785 59.425 167.955 ;
        RECT 56.535 166.955 56.705 167.135 ;
        RECT 53.335 166.245 54.405 166.415 ;
        RECT 54.575 166.035 54.765 166.475 ;
        RECT 54.935 166.205 55.885 166.485 ;
        RECT 56.195 166.395 56.455 166.785 ;
        RECT 56.875 166.715 57.665 166.965 ;
        RECT 56.105 166.225 56.455 166.395 ;
        RECT 56.665 166.035 56.995 166.495 ;
        RECT 57.870 166.425 58.040 167.135 ;
        RECT 58.395 166.935 58.565 167.525 ;
        RECT 58.210 166.715 58.565 166.935 ;
        RECT 58.735 166.715 59.085 167.335 ;
        RECT 59.255 166.425 59.425 167.785 ;
        RECT 59.790 167.615 60.115 168.400 ;
        RECT 59.595 166.565 60.055 167.615 ;
        RECT 57.870 166.255 58.725 166.425 ;
        RECT 58.930 166.255 59.425 166.425 ;
        RECT 59.595 166.035 59.925 166.395 ;
        RECT 60.285 166.295 60.455 168.415 ;
        RECT 60.625 168.085 60.955 168.585 ;
        RECT 61.125 167.915 61.380 168.415 ;
        RECT 60.630 167.745 61.380 167.915 ;
        RECT 60.630 166.755 60.860 167.745 ;
        RECT 61.030 166.925 61.380 167.575 ;
        RECT 61.555 167.420 61.845 168.585 ;
        RECT 62.940 167.435 63.200 168.585 ;
        RECT 63.375 167.510 63.630 168.415 ;
        RECT 63.800 167.825 64.130 168.585 ;
        RECT 64.345 167.655 64.515 168.415 ;
        RECT 60.630 166.585 61.380 166.755 ;
        RECT 60.625 166.035 60.955 166.415 ;
        RECT 61.125 166.295 61.380 166.585 ;
        RECT 61.555 166.035 61.845 166.760 ;
        RECT 62.940 166.035 63.200 166.875 ;
        RECT 63.375 166.780 63.545 167.510 ;
        RECT 63.800 167.485 64.515 167.655 ;
        RECT 63.800 167.275 63.970 167.485 ;
        RECT 64.925 167.435 65.255 168.585 ;
        RECT 65.425 167.565 65.595 168.415 ;
        RECT 65.765 167.785 66.095 168.585 ;
        RECT 66.265 167.565 66.435 168.415 ;
        RECT 66.615 167.785 66.855 168.585 ;
        RECT 67.025 167.605 67.355 168.415 ;
        RECT 65.425 167.395 66.435 167.565 ;
        RECT 66.640 167.435 67.355 167.605 ;
        RECT 67.540 167.435 67.800 168.585 ;
        RECT 67.975 167.510 68.230 168.415 ;
        RECT 68.400 167.825 68.730 168.585 ;
        RECT 68.945 167.655 69.115 168.415 ;
        RECT 63.715 166.945 63.970 167.275 ;
        RECT 63.375 166.205 63.630 166.780 ;
        RECT 63.800 166.755 63.970 166.945 ;
        RECT 64.250 166.935 64.605 167.305 ;
        RECT 65.425 166.855 65.920 167.395 ;
        RECT 66.640 167.195 66.810 167.435 ;
        RECT 66.310 167.025 66.810 167.195 ;
        RECT 66.980 167.025 67.360 167.265 ;
        RECT 66.640 166.855 66.810 167.025 ;
        RECT 63.800 166.585 64.515 166.755 ;
        RECT 63.800 166.035 64.130 166.415 ;
        RECT 64.345 166.205 64.515 166.585 ;
        RECT 64.925 166.035 65.255 166.835 ;
        RECT 65.425 166.685 66.435 166.855 ;
        RECT 66.640 166.685 67.275 166.855 ;
        RECT 65.425 166.205 65.595 166.685 ;
        RECT 65.765 166.035 66.095 166.515 ;
        RECT 66.265 166.205 66.435 166.685 ;
        RECT 66.685 166.035 66.925 166.515 ;
        RECT 67.105 166.205 67.275 166.685 ;
        RECT 67.540 166.035 67.800 166.875 ;
        RECT 67.975 166.780 68.145 167.510 ;
        RECT 68.400 167.485 69.115 167.655 ;
        RECT 69.375 167.615 69.685 168.415 ;
        RECT 69.855 167.785 70.165 168.585 ;
        RECT 70.335 167.955 70.595 168.415 ;
        RECT 70.765 168.125 71.020 168.585 ;
        RECT 71.195 167.955 71.455 168.415 ;
        RECT 70.335 167.785 71.455 167.955 ;
        RECT 68.400 167.275 68.570 167.485 ;
        RECT 69.375 167.445 70.405 167.615 ;
        RECT 68.315 166.945 68.570 167.275 ;
        RECT 67.975 166.205 68.230 166.780 ;
        RECT 68.400 166.755 68.570 166.945 ;
        RECT 68.850 166.935 69.205 167.305 ;
        RECT 68.400 166.585 69.115 166.755 ;
        RECT 68.400 166.035 68.730 166.415 ;
        RECT 68.945 166.205 69.115 166.585 ;
        RECT 69.375 166.535 69.545 167.445 ;
        RECT 69.715 166.705 70.065 167.275 ;
        RECT 70.235 167.195 70.405 167.445 ;
        RECT 71.195 167.535 71.455 167.785 ;
        RECT 71.625 167.715 71.910 168.585 ;
        RECT 72.225 167.655 72.395 168.415 ;
        RECT 72.610 167.825 72.940 168.585 ;
        RECT 71.195 167.365 71.950 167.535 ;
        RECT 72.225 167.485 72.940 167.655 ;
        RECT 73.110 167.510 73.365 168.415 ;
        RECT 70.235 167.025 71.375 167.195 ;
        RECT 71.545 166.855 71.950 167.365 ;
        RECT 72.135 166.935 72.490 167.305 ;
        RECT 72.770 167.275 72.940 167.485 ;
        RECT 72.770 166.945 73.025 167.275 ;
        RECT 70.300 166.685 71.950 166.855 ;
        RECT 72.770 166.755 72.940 166.945 ;
        RECT 73.195 166.780 73.365 167.510 ;
        RECT 73.540 167.435 73.800 168.585 ;
        RECT 74.440 167.445 74.775 168.415 ;
        RECT 74.945 167.445 75.115 168.585 ;
        RECT 75.285 168.245 77.315 168.415 ;
        RECT 69.375 166.205 69.675 166.535 ;
        RECT 69.845 166.035 70.120 166.515 ;
        RECT 70.300 166.295 70.595 166.685 ;
        RECT 70.765 166.035 71.020 166.515 ;
        RECT 71.195 166.295 71.455 166.685 ;
        RECT 72.225 166.585 72.940 166.755 ;
        RECT 71.625 166.035 71.905 166.515 ;
        RECT 72.225 166.205 72.395 166.585 ;
        RECT 72.610 166.035 72.940 166.415 ;
        RECT 73.110 166.205 73.365 166.780 ;
        RECT 73.540 166.035 73.800 166.875 ;
        RECT 74.440 166.775 74.610 167.445 ;
        RECT 75.285 167.275 75.455 168.245 ;
        RECT 74.780 166.945 75.035 167.275 ;
        RECT 75.260 166.945 75.455 167.275 ;
        RECT 75.625 167.905 76.750 168.075 ;
        RECT 74.865 166.775 75.035 166.945 ;
        RECT 75.625 166.775 75.795 167.905 ;
        RECT 74.440 166.205 74.695 166.775 ;
        RECT 74.865 166.605 75.795 166.775 ;
        RECT 75.965 167.565 76.975 167.735 ;
        RECT 75.965 166.765 76.135 167.565 ;
        RECT 75.620 166.570 75.795 166.605 ;
        RECT 74.865 166.035 75.195 166.435 ;
        RECT 75.620 166.205 76.150 166.570 ;
        RECT 76.340 166.545 76.615 167.365 ;
        RECT 76.335 166.375 76.615 166.545 ;
        RECT 76.340 166.205 76.615 166.375 ;
        RECT 76.785 166.205 76.975 167.565 ;
        RECT 77.145 167.580 77.315 168.245 ;
        RECT 77.485 167.825 77.655 168.585 ;
        RECT 77.890 167.825 78.405 168.235 ;
        RECT 77.145 167.390 77.895 167.580 ;
        RECT 78.065 167.015 78.405 167.825 ;
        RECT 77.175 166.845 78.405 167.015 ;
        RECT 79.035 167.825 79.550 168.235 ;
        RECT 79.785 167.825 79.955 168.585 ;
        RECT 80.125 168.245 82.155 168.415 ;
        RECT 79.035 167.015 79.375 167.825 ;
        RECT 80.125 167.580 80.295 168.245 ;
        RECT 80.690 167.905 81.815 168.075 ;
        RECT 79.545 167.390 80.295 167.580 ;
        RECT 80.465 167.565 81.475 167.735 ;
        RECT 79.035 166.845 80.265 167.015 ;
        RECT 77.155 166.035 77.665 166.570 ;
        RECT 77.885 166.240 78.130 166.845 ;
        RECT 79.310 166.240 79.555 166.845 ;
        RECT 79.775 166.035 80.285 166.570 ;
        RECT 80.465 166.205 80.655 167.565 ;
        RECT 80.825 167.225 81.100 167.365 ;
        RECT 80.825 167.055 81.105 167.225 ;
        RECT 80.825 166.205 81.100 167.055 ;
        RECT 81.305 166.765 81.475 167.565 ;
        RECT 81.645 166.775 81.815 167.905 ;
        RECT 81.985 167.275 82.155 168.245 ;
        RECT 82.325 167.445 82.495 168.585 ;
        RECT 82.665 167.445 83.000 168.415 ;
        RECT 81.985 166.945 82.180 167.275 ;
        RECT 82.405 166.945 82.660 167.275 ;
        RECT 82.405 166.775 82.575 166.945 ;
        RECT 82.830 166.775 83.000 167.445 ;
        RECT 83.175 167.825 83.690 168.235 ;
        RECT 83.925 167.825 84.095 168.585 ;
        RECT 84.265 168.245 86.295 168.415 ;
        RECT 83.175 167.015 83.515 167.825 ;
        RECT 84.265 167.580 84.435 168.245 ;
        RECT 84.830 167.905 85.955 168.075 ;
        RECT 83.685 167.390 84.435 167.580 ;
        RECT 84.605 167.565 85.615 167.735 ;
        RECT 83.175 166.845 84.405 167.015 ;
        RECT 81.645 166.605 82.575 166.775 ;
        RECT 81.645 166.570 81.820 166.605 ;
        RECT 81.290 166.205 81.820 166.570 ;
        RECT 82.245 166.035 82.575 166.435 ;
        RECT 82.745 166.205 83.000 166.775 ;
        RECT 83.450 166.240 83.695 166.845 ;
        RECT 83.915 166.035 84.425 166.570 ;
        RECT 84.605 166.205 84.795 167.565 ;
        RECT 84.965 167.225 85.240 167.365 ;
        RECT 84.965 167.055 85.245 167.225 ;
        RECT 84.965 166.205 85.240 167.055 ;
        RECT 85.445 166.765 85.615 167.565 ;
        RECT 85.785 166.775 85.955 167.905 ;
        RECT 86.125 167.275 86.295 168.245 ;
        RECT 86.465 167.445 86.635 168.585 ;
        RECT 86.805 167.445 87.140 168.415 ;
        RECT 86.125 166.945 86.320 167.275 ;
        RECT 86.545 166.945 86.800 167.275 ;
        RECT 86.545 166.775 86.715 166.945 ;
        RECT 86.970 166.775 87.140 167.445 ;
        RECT 87.315 167.420 87.605 168.585 ;
        RECT 88.150 168.245 88.405 168.275 ;
        RECT 88.065 168.075 88.405 168.245 ;
        RECT 88.150 167.605 88.405 168.075 ;
        RECT 88.585 167.785 88.870 168.585 ;
        RECT 89.050 167.865 89.380 168.375 ;
        RECT 85.785 166.605 86.715 166.775 ;
        RECT 85.785 166.570 85.960 166.605 ;
        RECT 85.430 166.205 85.960 166.570 ;
        RECT 86.385 166.035 86.715 166.435 ;
        RECT 86.885 166.205 87.140 166.775 ;
        RECT 87.315 166.035 87.605 166.760 ;
        RECT 88.150 166.745 88.330 167.605 ;
        RECT 89.050 167.275 89.300 167.865 ;
        RECT 89.650 167.715 89.820 168.325 ;
        RECT 89.990 167.895 90.320 168.585 ;
        RECT 90.550 168.035 90.790 168.325 ;
        RECT 90.990 168.205 91.410 168.585 ;
        RECT 91.590 168.115 92.220 168.365 ;
        RECT 92.690 168.205 93.020 168.585 ;
        RECT 91.590 168.035 91.760 168.115 ;
        RECT 93.190 168.035 93.360 168.325 ;
        RECT 93.540 168.205 93.920 168.585 ;
        RECT 94.160 168.200 94.990 168.370 ;
        RECT 90.550 167.865 91.760 168.035 ;
        RECT 88.500 166.945 89.300 167.275 ;
        RECT 88.150 166.215 88.405 166.745 ;
        RECT 88.585 166.035 88.870 166.495 ;
        RECT 89.050 166.295 89.300 166.945 ;
        RECT 89.500 167.695 89.820 167.715 ;
        RECT 89.500 167.525 91.420 167.695 ;
        RECT 89.500 166.630 89.690 167.525 ;
        RECT 91.590 167.355 91.760 167.865 ;
        RECT 91.930 167.605 92.450 167.915 ;
        RECT 89.860 167.185 91.760 167.355 ;
        RECT 89.860 167.125 90.190 167.185 ;
        RECT 90.340 166.955 90.670 167.015 ;
        RECT 90.010 166.685 90.670 166.955 ;
        RECT 89.500 166.300 89.820 166.630 ;
        RECT 90.000 166.035 90.660 166.515 ;
        RECT 90.860 166.425 91.030 167.185 ;
        RECT 91.930 167.015 92.110 167.425 ;
        RECT 91.200 166.845 91.530 166.965 ;
        RECT 92.280 166.845 92.450 167.605 ;
        RECT 91.200 166.675 92.450 166.845 ;
        RECT 92.620 167.785 93.990 168.035 ;
        RECT 92.620 167.015 92.810 167.785 ;
        RECT 93.740 167.525 93.990 167.785 ;
        RECT 92.980 167.355 93.230 167.515 ;
        RECT 94.160 167.355 94.330 168.200 ;
        RECT 95.225 167.915 95.395 168.415 ;
        RECT 95.565 168.085 95.895 168.585 ;
        RECT 94.500 167.525 95.000 167.905 ;
        RECT 95.225 167.745 95.920 167.915 ;
        RECT 92.980 167.185 94.330 167.355 ;
        RECT 93.910 167.145 94.330 167.185 ;
        RECT 92.620 166.675 93.040 167.015 ;
        RECT 93.330 166.685 93.740 167.015 ;
        RECT 90.860 166.255 91.710 166.425 ;
        RECT 92.270 166.035 92.590 166.495 ;
        RECT 92.790 166.245 93.040 166.675 ;
        RECT 93.330 166.035 93.740 166.475 ;
        RECT 93.910 166.415 94.080 167.145 ;
        RECT 94.250 166.595 94.600 166.965 ;
        RECT 94.780 166.655 95.000 167.525 ;
        RECT 95.170 166.955 95.580 167.575 ;
        RECT 95.750 166.775 95.920 167.745 ;
        RECT 95.225 166.585 95.920 166.775 ;
        RECT 93.910 166.215 94.925 166.415 ;
        RECT 95.225 166.255 95.395 166.585 ;
        RECT 95.565 166.035 95.895 166.415 ;
        RECT 96.110 166.295 96.335 168.415 ;
        RECT 96.505 168.085 96.835 168.585 ;
        RECT 97.005 167.915 97.175 168.415 ;
        RECT 96.510 167.745 97.175 167.915 ;
        RECT 98.010 167.955 98.295 168.415 ;
        RECT 98.465 168.125 98.735 168.585 ;
        RECT 96.510 166.755 96.740 167.745 ;
        RECT 98.010 167.735 98.965 167.955 ;
        RECT 96.910 166.925 97.260 167.575 ;
        RECT 97.895 167.005 98.585 167.565 ;
        RECT 98.755 166.835 98.965 167.735 ;
        RECT 96.510 166.585 97.175 166.755 ;
        RECT 96.505 166.035 96.835 166.415 ;
        RECT 97.005 166.295 97.175 166.585 ;
        RECT 98.010 166.665 98.965 166.835 ;
        RECT 99.135 167.565 99.535 168.415 ;
        RECT 99.725 167.955 100.005 168.415 ;
        RECT 100.525 168.125 100.850 168.585 ;
        RECT 99.725 167.735 100.850 167.955 ;
        RECT 99.135 167.005 100.230 167.565 ;
        RECT 100.400 167.275 100.850 167.735 ;
        RECT 101.020 167.445 101.405 168.415 ;
        RECT 98.010 166.205 98.295 166.665 ;
        RECT 98.465 166.035 98.735 166.495 ;
        RECT 99.135 166.205 99.535 167.005 ;
        RECT 100.400 166.945 100.955 167.275 ;
        RECT 100.400 166.835 100.850 166.945 ;
        RECT 99.725 166.665 100.850 166.835 ;
        RECT 101.125 166.775 101.405 167.445 ;
        RECT 101.575 167.825 102.090 168.235 ;
        RECT 102.325 167.825 102.495 168.585 ;
        RECT 102.665 168.245 104.695 168.415 ;
        RECT 101.575 167.015 101.915 167.825 ;
        RECT 102.665 167.580 102.835 168.245 ;
        RECT 103.230 167.905 104.355 168.075 ;
        RECT 102.085 167.390 102.835 167.580 ;
        RECT 103.005 167.565 104.015 167.735 ;
        RECT 101.575 166.845 102.805 167.015 ;
        RECT 99.725 166.205 100.005 166.665 ;
        RECT 100.525 166.035 100.850 166.495 ;
        RECT 101.020 166.205 101.405 166.775 ;
        RECT 101.850 166.240 102.095 166.845 ;
        RECT 102.315 166.035 102.825 166.570 ;
        RECT 103.005 166.205 103.195 167.565 ;
        RECT 103.365 166.545 103.640 167.365 ;
        RECT 103.845 166.765 104.015 167.565 ;
        RECT 104.185 166.775 104.355 167.905 ;
        RECT 104.525 167.275 104.695 168.245 ;
        RECT 104.865 167.445 105.035 168.585 ;
        RECT 105.205 167.445 105.540 168.415 ;
        RECT 104.525 166.945 104.720 167.275 ;
        RECT 104.945 166.945 105.200 167.275 ;
        RECT 104.945 166.775 105.115 166.945 ;
        RECT 105.370 166.775 105.540 167.445 ;
        RECT 104.185 166.605 105.115 166.775 ;
        RECT 104.185 166.570 104.360 166.605 ;
        RECT 103.365 166.375 103.645 166.545 ;
        RECT 103.365 166.205 103.640 166.375 ;
        RECT 103.830 166.205 104.360 166.570 ;
        RECT 104.785 166.035 105.115 166.435 ;
        RECT 105.285 166.205 105.540 166.775 ;
        RECT 105.715 167.445 106.100 168.415 ;
        RECT 106.270 168.125 106.595 168.585 ;
        RECT 107.115 167.955 107.395 168.415 ;
        RECT 106.270 167.735 107.395 167.955 ;
        RECT 105.715 166.775 105.995 167.445 ;
        RECT 106.270 167.275 106.720 167.735 ;
        RECT 107.585 167.565 107.985 168.415 ;
        RECT 108.385 168.125 108.655 168.585 ;
        RECT 108.825 167.955 109.110 168.415 ;
        RECT 106.165 166.945 106.720 167.275 ;
        RECT 106.890 167.005 107.985 167.565 ;
        RECT 106.270 166.835 106.720 166.945 ;
        RECT 105.715 166.205 106.100 166.775 ;
        RECT 106.270 166.665 107.395 166.835 ;
        RECT 106.270 166.035 106.595 166.495 ;
        RECT 107.115 166.205 107.395 166.665 ;
        RECT 107.585 166.205 107.985 167.005 ;
        RECT 108.155 167.735 109.110 167.955 ;
        RECT 108.155 166.835 108.365 167.735 ;
        RECT 108.535 167.005 109.225 167.565 ;
        RECT 109.545 167.435 109.875 168.585 ;
        RECT 110.045 167.565 110.215 168.415 ;
        RECT 110.385 167.785 110.715 168.585 ;
        RECT 110.885 167.565 111.055 168.415 ;
        RECT 111.235 167.785 111.475 168.585 ;
        RECT 111.645 167.605 111.975 168.415 ;
        RECT 110.045 167.395 111.055 167.565 ;
        RECT 111.260 167.435 111.975 167.605 ;
        RECT 112.155 167.495 113.365 168.585 ;
        RECT 110.045 166.885 110.540 167.395 ;
        RECT 111.260 167.195 111.430 167.435 ;
        RECT 110.930 167.025 111.430 167.195 ;
        RECT 111.600 167.025 111.980 167.265 ;
        RECT 110.045 166.855 110.545 166.885 ;
        RECT 111.260 166.855 111.430 167.025 ;
        RECT 112.155 166.955 112.675 167.495 ;
        RECT 108.155 166.665 109.110 166.835 ;
        RECT 108.385 166.035 108.655 166.495 ;
        RECT 108.825 166.205 109.110 166.665 ;
        RECT 109.545 166.035 109.875 166.835 ;
        RECT 110.045 166.685 111.055 166.855 ;
        RECT 111.260 166.685 111.895 166.855 ;
        RECT 112.845 166.785 113.365 167.325 ;
        RECT 110.045 166.205 110.215 166.685 ;
        RECT 110.385 166.035 110.715 166.515 ;
        RECT 110.885 166.205 111.055 166.685 ;
        RECT 111.305 166.035 111.545 166.515 ;
        RECT 111.725 166.205 111.895 166.685 ;
        RECT 112.155 166.035 113.365 166.785 ;
        RECT 22.830 165.865 113.450 166.035 ;
        RECT 22.915 165.115 24.125 165.865 ;
        RECT 24.670 165.155 24.925 165.685 ;
        RECT 25.105 165.405 25.390 165.865 ;
        RECT 22.915 164.575 23.435 165.115 ;
        RECT 23.605 164.405 24.125 164.945 ;
        RECT 24.670 164.505 24.850 165.155 ;
        RECT 25.570 164.955 25.820 165.605 ;
        RECT 25.020 164.625 25.820 164.955 ;
        RECT 22.915 163.315 24.125 164.405 ;
        RECT 24.585 164.335 24.850 164.505 ;
        RECT 24.670 164.295 24.850 164.335 ;
        RECT 24.670 163.625 24.925 164.295 ;
        RECT 25.105 163.315 25.390 164.115 ;
        RECT 25.570 164.035 25.820 164.625 ;
        RECT 26.020 165.270 26.340 165.600 ;
        RECT 26.520 165.385 27.180 165.865 ;
        RECT 27.380 165.475 28.230 165.645 ;
        RECT 26.020 164.375 26.210 165.270 ;
        RECT 26.530 164.945 27.190 165.215 ;
        RECT 26.860 164.885 27.190 164.945 ;
        RECT 26.380 164.715 26.710 164.775 ;
        RECT 27.380 164.715 27.550 165.475 ;
        RECT 28.790 165.405 29.110 165.865 ;
        RECT 29.310 165.225 29.560 165.655 ;
        RECT 29.850 165.425 30.260 165.865 ;
        RECT 30.430 165.485 31.445 165.685 ;
        RECT 27.720 165.055 28.970 165.225 ;
        RECT 27.720 164.935 28.050 165.055 ;
        RECT 26.380 164.545 28.280 164.715 ;
        RECT 26.020 164.205 27.940 164.375 ;
        RECT 26.020 164.185 26.340 164.205 ;
        RECT 25.570 163.525 25.900 164.035 ;
        RECT 26.170 163.575 26.340 164.185 ;
        RECT 28.110 164.035 28.280 164.545 ;
        RECT 28.450 164.475 28.630 164.885 ;
        RECT 28.800 164.295 28.970 165.055 ;
        RECT 26.510 163.315 26.840 164.005 ;
        RECT 27.070 163.865 28.280 164.035 ;
        RECT 28.450 163.985 28.970 164.295 ;
        RECT 29.140 164.885 29.560 165.225 ;
        RECT 29.850 164.885 30.260 165.215 ;
        RECT 29.140 164.115 29.330 164.885 ;
        RECT 30.430 164.755 30.600 165.485 ;
        RECT 31.745 165.315 31.915 165.645 ;
        RECT 32.085 165.485 32.415 165.865 ;
        RECT 30.770 164.935 31.120 165.305 ;
        RECT 30.430 164.715 30.850 164.755 ;
        RECT 29.500 164.545 30.850 164.715 ;
        RECT 29.500 164.385 29.750 164.545 ;
        RECT 30.260 164.115 30.510 164.375 ;
        RECT 29.140 163.865 30.510 164.115 ;
        RECT 27.070 163.575 27.310 163.865 ;
        RECT 28.110 163.785 28.280 163.865 ;
        RECT 27.510 163.315 27.930 163.695 ;
        RECT 28.110 163.535 28.740 163.785 ;
        RECT 29.210 163.315 29.540 163.695 ;
        RECT 29.710 163.575 29.880 163.865 ;
        RECT 30.680 163.700 30.850 164.545 ;
        RECT 31.300 164.375 31.520 165.245 ;
        RECT 31.745 165.125 32.440 165.315 ;
        RECT 31.020 163.995 31.520 164.375 ;
        RECT 31.690 164.325 32.100 164.945 ;
        RECT 32.270 164.155 32.440 165.125 ;
        RECT 31.745 163.985 32.440 164.155 ;
        RECT 30.060 163.315 30.440 163.695 ;
        RECT 30.680 163.530 31.510 163.700 ;
        RECT 31.745 163.485 31.915 163.985 ;
        RECT 32.085 163.315 32.415 163.815 ;
        RECT 32.630 163.485 32.855 165.605 ;
        RECT 33.025 165.485 33.355 165.865 ;
        RECT 33.525 165.315 33.695 165.605 ;
        RECT 33.030 165.145 33.695 165.315 ;
        RECT 34.070 165.235 34.355 165.695 ;
        RECT 34.525 165.405 34.795 165.865 ;
        RECT 33.030 164.155 33.260 165.145 ;
        RECT 34.070 165.065 35.025 165.235 ;
        RECT 33.430 164.325 33.780 164.975 ;
        RECT 33.955 164.335 34.645 164.895 ;
        RECT 34.815 164.165 35.025 165.065 ;
        RECT 33.030 163.985 33.695 164.155 ;
        RECT 33.025 163.315 33.355 163.815 ;
        RECT 33.525 163.485 33.695 163.985 ;
        RECT 34.070 163.945 35.025 164.165 ;
        RECT 35.195 164.895 35.595 165.695 ;
        RECT 35.785 165.235 36.065 165.695 ;
        RECT 36.585 165.405 36.910 165.865 ;
        RECT 35.785 165.065 36.910 165.235 ;
        RECT 37.080 165.125 37.465 165.695 ;
        RECT 36.460 164.955 36.910 165.065 ;
        RECT 35.195 164.335 36.290 164.895 ;
        RECT 36.460 164.625 37.015 164.955 ;
        RECT 34.070 163.485 34.355 163.945 ;
        RECT 34.525 163.315 34.795 163.775 ;
        RECT 35.195 163.485 35.595 164.335 ;
        RECT 36.460 164.165 36.910 164.625 ;
        RECT 37.185 164.455 37.465 165.125 ;
        RECT 37.750 165.235 38.035 165.695 ;
        RECT 38.205 165.405 38.475 165.865 ;
        RECT 37.750 165.065 38.705 165.235 ;
        RECT 35.785 163.945 36.910 164.165 ;
        RECT 35.785 163.485 36.065 163.945 ;
        RECT 36.585 163.315 36.910 163.775 ;
        RECT 37.080 163.485 37.465 164.455 ;
        RECT 37.635 164.335 38.325 164.895 ;
        RECT 38.495 164.165 38.705 165.065 ;
        RECT 37.750 163.945 38.705 164.165 ;
        RECT 38.875 164.895 39.275 165.695 ;
        RECT 39.465 165.235 39.745 165.695 ;
        RECT 40.265 165.405 40.590 165.865 ;
        RECT 39.465 165.065 40.590 165.235 ;
        RECT 40.760 165.125 41.145 165.695 ;
        RECT 40.140 164.955 40.590 165.065 ;
        RECT 38.875 164.335 39.970 164.895 ;
        RECT 40.140 164.625 40.695 164.955 ;
        RECT 37.750 163.485 38.035 163.945 ;
        RECT 38.205 163.315 38.475 163.775 ;
        RECT 38.875 163.485 39.275 164.335 ;
        RECT 40.140 164.165 40.590 164.625 ;
        RECT 40.865 164.455 41.145 165.125 ;
        RECT 41.430 165.235 41.715 165.695 ;
        RECT 41.885 165.405 42.155 165.865 ;
        RECT 41.430 165.065 42.385 165.235 ;
        RECT 39.465 163.945 40.590 164.165 ;
        RECT 39.465 163.485 39.745 163.945 ;
        RECT 40.265 163.315 40.590 163.775 ;
        RECT 40.760 163.485 41.145 164.455 ;
        RECT 41.315 164.335 42.005 164.895 ;
        RECT 42.175 164.165 42.385 165.065 ;
        RECT 41.430 163.945 42.385 164.165 ;
        RECT 42.555 164.895 42.955 165.695 ;
        RECT 43.145 165.235 43.425 165.695 ;
        RECT 43.945 165.405 44.270 165.865 ;
        RECT 43.145 165.065 44.270 165.235 ;
        RECT 44.440 165.125 44.825 165.695 ;
        RECT 43.820 164.955 44.270 165.065 ;
        RECT 42.555 164.335 43.650 164.895 ;
        RECT 43.820 164.625 44.375 164.955 ;
        RECT 41.430 163.485 41.715 163.945 ;
        RECT 41.885 163.315 42.155 163.775 ;
        RECT 42.555 163.485 42.955 164.335 ;
        RECT 43.820 164.165 44.270 164.625 ;
        RECT 44.545 164.455 44.825 165.125 ;
        RECT 45.110 165.235 45.395 165.695 ;
        RECT 45.565 165.405 45.835 165.865 ;
        RECT 45.110 165.065 46.065 165.235 ;
        RECT 43.145 163.945 44.270 164.165 ;
        RECT 43.145 163.485 43.425 163.945 ;
        RECT 43.945 163.315 44.270 163.775 ;
        RECT 44.440 163.485 44.825 164.455 ;
        RECT 44.995 164.335 45.685 164.895 ;
        RECT 45.855 164.165 46.065 165.065 ;
        RECT 45.110 163.945 46.065 164.165 ;
        RECT 46.235 164.895 46.635 165.695 ;
        RECT 46.825 165.235 47.105 165.695 ;
        RECT 47.625 165.405 47.950 165.865 ;
        RECT 46.825 165.065 47.950 165.235 ;
        RECT 48.120 165.125 48.505 165.695 ;
        RECT 48.675 165.140 48.965 165.865 ;
        RECT 47.500 164.955 47.950 165.065 ;
        RECT 46.235 164.335 47.330 164.895 ;
        RECT 47.500 164.625 48.055 164.955 ;
        RECT 45.110 163.485 45.395 163.945 ;
        RECT 45.565 163.315 45.835 163.775 ;
        RECT 46.235 163.485 46.635 164.335 ;
        RECT 47.500 164.165 47.950 164.625 ;
        RECT 48.225 164.455 48.505 165.125 ;
        RECT 49.595 165.095 51.265 165.865 ;
        RECT 46.825 163.945 47.950 164.165 ;
        RECT 46.825 163.485 47.105 163.945 ;
        RECT 47.625 163.315 47.950 163.775 ;
        RECT 48.120 163.485 48.505 164.455 ;
        RECT 48.675 163.315 48.965 164.480 ;
        RECT 49.595 164.405 50.345 164.925 ;
        RECT 50.515 164.575 51.265 165.095 ;
        RECT 51.440 165.125 51.695 165.695 ;
        RECT 51.865 165.465 52.195 165.865 ;
        RECT 52.620 165.330 53.150 165.695 ;
        RECT 52.620 165.295 52.795 165.330 ;
        RECT 51.865 165.125 52.795 165.295 ;
        RECT 53.340 165.185 53.615 165.695 ;
        RECT 51.440 164.455 51.610 165.125 ;
        RECT 51.865 164.955 52.035 165.125 ;
        RECT 51.780 164.625 52.035 164.955 ;
        RECT 52.260 164.625 52.455 164.955 ;
        RECT 49.595 163.315 51.265 164.405 ;
        RECT 51.440 163.485 51.775 164.455 ;
        RECT 51.945 163.315 52.115 164.455 ;
        RECT 52.285 163.655 52.455 164.625 ;
        RECT 52.625 163.995 52.795 165.125 ;
        RECT 52.965 164.335 53.135 165.135 ;
        RECT 53.335 165.015 53.615 165.185 ;
        RECT 53.340 164.535 53.615 165.015 ;
        RECT 53.785 164.335 53.975 165.695 ;
        RECT 54.155 165.330 54.665 165.865 ;
        RECT 54.885 165.055 55.130 165.660 ;
        RECT 55.850 165.055 56.095 165.660 ;
        RECT 56.315 165.330 56.825 165.865 ;
        RECT 54.175 164.885 55.405 165.055 ;
        RECT 52.965 164.165 53.975 164.335 ;
        RECT 54.145 164.320 54.895 164.510 ;
        RECT 52.625 163.825 53.750 163.995 ;
        RECT 54.145 163.655 54.315 164.320 ;
        RECT 55.065 164.075 55.405 164.885 ;
        RECT 52.285 163.485 54.315 163.655 ;
        RECT 54.485 163.315 54.655 164.075 ;
        RECT 54.890 163.665 55.405 164.075 ;
        RECT 55.575 164.885 56.805 165.055 ;
        RECT 55.575 164.075 55.915 164.885 ;
        RECT 56.085 164.320 56.835 164.510 ;
        RECT 55.575 163.665 56.090 164.075 ;
        RECT 56.325 163.315 56.495 164.075 ;
        RECT 56.665 163.655 56.835 164.320 ;
        RECT 57.005 164.335 57.195 165.695 ;
        RECT 57.365 164.845 57.640 165.695 ;
        RECT 57.830 165.330 58.360 165.695 ;
        RECT 58.785 165.465 59.115 165.865 ;
        RECT 58.185 165.295 58.360 165.330 ;
        RECT 57.365 164.675 57.645 164.845 ;
        RECT 57.365 164.535 57.640 164.675 ;
        RECT 57.845 164.335 58.015 165.135 ;
        RECT 57.005 164.165 58.015 164.335 ;
        RECT 58.185 165.125 59.115 165.295 ;
        RECT 59.285 165.125 59.540 165.695 ;
        RECT 58.185 163.995 58.355 165.125 ;
        RECT 58.945 164.955 59.115 165.125 ;
        RECT 57.230 163.825 58.355 163.995 ;
        RECT 58.525 164.625 58.720 164.955 ;
        RECT 58.945 164.625 59.200 164.955 ;
        RECT 58.525 163.655 58.695 164.625 ;
        RECT 59.370 164.455 59.540 165.125 ;
        RECT 56.665 163.485 58.695 163.655 ;
        RECT 58.865 163.315 59.035 164.455 ;
        RECT 59.205 163.485 59.540 164.455 ;
        RECT 59.720 165.155 59.975 165.685 ;
        RECT 60.145 165.405 60.450 165.865 ;
        RECT 60.695 165.485 61.765 165.655 ;
        RECT 59.720 164.505 59.930 165.155 ;
        RECT 60.695 165.130 61.015 165.485 ;
        RECT 60.690 164.955 61.015 165.130 ;
        RECT 60.100 164.655 61.015 164.955 ;
        RECT 61.185 164.915 61.425 165.315 ;
        RECT 61.595 165.255 61.765 165.485 ;
        RECT 61.935 165.425 62.125 165.865 ;
        RECT 62.295 165.415 63.245 165.695 ;
        RECT 63.465 165.505 63.815 165.675 ;
        RECT 61.595 165.085 62.125 165.255 ;
        RECT 60.100 164.625 60.840 164.655 ;
        RECT 59.720 163.625 59.975 164.505 ;
        RECT 60.145 163.315 60.450 164.455 ;
        RECT 60.670 164.035 60.840 164.625 ;
        RECT 61.185 164.545 61.725 164.915 ;
        RECT 61.905 164.805 62.125 165.085 ;
        RECT 62.295 164.635 62.465 165.415 ;
        RECT 62.060 164.465 62.465 164.635 ;
        RECT 62.635 164.625 62.985 165.245 ;
        RECT 62.060 164.375 62.230 164.465 ;
        RECT 63.155 164.455 63.365 165.245 ;
        RECT 61.010 164.205 62.230 164.375 ;
        RECT 62.690 164.295 63.365 164.455 ;
        RECT 60.670 163.865 61.470 164.035 ;
        RECT 60.790 163.315 61.120 163.695 ;
        RECT 61.300 163.575 61.470 163.865 ;
        RECT 62.060 163.825 62.230 164.205 ;
        RECT 62.400 164.285 63.365 164.295 ;
        RECT 63.555 165.115 63.815 165.505 ;
        RECT 64.025 165.405 64.355 165.865 ;
        RECT 65.230 165.475 66.085 165.645 ;
        RECT 66.290 165.475 66.785 165.645 ;
        RECT 66.955 165.505 67.285 165.865 ;
        RECT 63.555 164.425 63.725 165.115 ;
        RECT 63.895 164.765 64.065 164.945 ;
        RECT 64.235 164.935 65.025 165.185 ;
        RECT 65.230 164.765 65.400 165.475 ;
        RECT 65.570 164.965 65.925 165.185 ;
        RECT 63.895 164.595 65.585 164.765 ;
        RECT 62.400 163.995 62.860 164.285 ;
        RECT 63.555 164.255 65.055 164.425 ;
        RECT 63.555 164.115 63.725 164.255 ;
        RECT 63.165 163.945 63.725 164.115 ;
        RECT 61.640 163.315 61.890 163.775 ;
        RECT 62.060 163.485 62.930 163.825 ;
        RECT 63.165 163.485 63.335 163.945 ;
        RECT 64.170 163.915 65.245 164.085 ;
        RECT 63.505 163.315 63.875 163.775 ;
        RECT 64.170 163.575 64.340 163.915 ;
        RECT 64.510 163.315 64.840 163.745 ;
        RECT 65.075 163.575 65.245 163.915 ;
        RECT 65.415 163.815 65.585 164.595 ;
        RECT 65.755 164.375 65.925 164.965 ;
        RECT 66.095 164.565 66.445 165.185 ;
        RECT 65.755 163.985 66.220 164.375 ;
        RECT 66.615 164.115 66.785 165.475 ;
        RECT 66.955 164.285 67.415 165.335 ;
        RECT 66.390 163.945 66.785 164.115 ;
        RECT 66.390 163.815 66.560 163.945 ;
        RECT 65.415 163.485 66.095 163.815 ;
        RECT 66.310 163.485 66.560 163.815 ;
        RECT 66.730 163.315 66.980 163.775 ;
        RECT 67.150 163.500 67.475 164.285 ;
        RECT 67.645 163.485 67.815 165.605 ;
        RECT 67.985 165.485 68.315 165.865 ;
        RECT 68.485 165.315 68.740 165.605 ;
        RECT 67.990 165.145 68.740 165.315 ;
        RECT 69.005 165.315 69.175 165.695 ;
        RECT 69.390 165.485 69.720 165.865 ;
        RECT 69.005 165.145 69.720 165.315 ;
        RECT 67.990 164.155 68.220 165.145 ;
        RECT 68.390 164.325 68.740 164.975 ;
        RECT 68.915 164.595 69.270 164.965 ;
        RECT 69.550 164.955 69.720 165.145 ;
        RECT 69.890 165.120 70.145 165.695 ;
        RECT 69.550 164.625 69.805 164.955 ;
        RECT 69.550 164.415 69.720 164.625 ;
        RECT 69.005 164.245 69.720 164.415 ;
        RECT 69.975 164.390 70.145 165.120 ;
        RECT 70.320 165.025 70.580 165.865 ;
        RECT 70.960 165.085 71.460 165.695 ;
        RECT 70.755 164.625 71.105 164.875 ;
        RECT 67.990 163.985 68.740 164.155 ;
        RECT 67.985 163.315 68.315 163.815 ;
        RECT 68.485 163.485 68.740 163.985 ;
        RECT 69.005 163.485 69.175 164.245 ;
        RECT 69.390 163.315 69.720 164.075 ;
        RECT 69.890 163.485 70.145 164.390 ;
        RECT 70.320 163.315 70.580 164.465 ;
        RECT 71.290 164.455 71.460 165.085 ;
        RECT 72.090 165.215 72.420 165.695 ;
        RECT 72.590 165.405 72.815 165.865 ;
        RECT 72.985 165.215 73.315 165.695 ;
        RECT 72.090 165.045 73.315 165.215 ;
        RECT 73.505 165.065 73.755 165.865 ;
        RECT 73.925 165.065 74.265 165.695 ;
        RECT 74.435 165.140 74.725 165.865 ;
        RECT 74.985 165.315 75.155 165.695 ;
        RECT 75.335 165.485 75.665 165.865 ;
        RECT 74.985 165.145 75.650 165.315 ;
        RECT 75.845 165.190 76.105 165.695 ;
        RECT 71.630 164.675 71.960 164.875 ;
        RECT 72.130 164.675 72.460 164.875 ;
        RECT 72.630 164.675 73.050 164.875 ;
        RECT 73.225 164.705 73.920 164.875 ;
        RECT 73.225 164.455 73.395 164.705 ;
        RECT 74.090 164.455 74.265 165.065 ;
        RECT 74.915 164.595 75.245 164.965 ;
        RECT 75.480 164.890 75.650 165.145 ;
        RECT 75.480 164.560 75.765 164.890 ;
        RECT 70.960 164.285 73.395 164.455 ;
        RECT 70.960 163.485 71.290 164.285 ;
        RECT 71.460 163.315 71.790 164.115 ;
        RECT 72.090 163.485 72.420 164.285 ;
        RECT 73.065 163.315 73.315 164.115 ;
        RECT 73.585 163.315 73.755 164.455 ;
        RECT 73.925 163.485 74.265 164.455 ;
        RECT 74.435 163.315 74.725 164.480 ;
        RECT 75.480 164.415 75.650 164.560 ;
        RECT 74.985 164.245 75.650 164.415 ;
        RECT 75.935 164.390 76.105 165.190 ;
        RECT 76.550 165.055 76.795 165.660 ;
        RECT 77.015 165.330 77.525 165.865 ;
        RECT 74.985 163.485 75.155 164.245 ;
        RECT 75.335 163.315 75.665 164.075 ;
        RECT 75.835 163.485 76.105 164.390 ;
        RECT 76.275 164.885 77.505 165.055 ;
        RECT 76.275 164.075 76.615 164.885 ;
        RECT 76.785 164.320 77.535 164.510 ;
        RECT 76.275 163.665 76.790 164.075 ;
        RECT 77.025 163.315 77.195 164.075 ;
        RECT 77.365 163.655 77.535 164.320 ;
        RECT 77.705 164.335 77.895 165.695 ;
        RECT 78.065 164.845 78.340 165.695 ;
        RECT 78.530 165.330 79.060 165.695 ;
        RECT 79.485 165.465 79.815 165.865 ;
        RECT 78.885 165.295 79.060 165.330 ;
        RECT 78.065 164.675 78.345 164.845 ;
        RECT 78.065 164.535 78.340 164.675 ;
        RECT 78.545 164.335 78.715 165.135 ;
        RECT 77.705 164.165 78.715 164.335 ;
        RECT 78.885 165.125 79.815 165.295 ;
        RECT 79.985 165.125 80.240 165.695 ;
        RECT 78.885 163.995 79.055 165.125 ;
        RECT 79.645 164.955 79.815 165.125 ;
        RECT 77.930 163.825 79.055 163.995 ;
        RECT 79.225 164.625 79.420 164.955 ;
        RECT 79.645 164.625 79.900 164.955 ;
        RECT 79.225 163.655 79.395 164.625 ;
        RECT 80.070 164.455 80.240 165.125 ;
        RECT 80.790 165.155 81.045 165.685 ;
        RECT 81.225 165.405 81.510 165.865 ;
        RECT 80.790 164.845 80.970 165.155 ;
        RECT 81.690 164.955 81.940 165.605 ;
        RECT 80.705 164.675 80.970 164.845 ;
        RECT 77.365 163.485 79.395 163.655 ;
        RECT 79.565 163.315 79.735 164.455 ;
        RECT 79.905 163.485 80.240 164.455 ;
        RECT 80.790 164.295 80.970 164.675 ;
        RECT 81.140 164.625 81.940 164.955 ;
        RECT 80.790 163.625 81.045 164.295 ;
        RECT 81.225 163.315 81.510 164.115 ;
        RECT 81.690 164.035 81.940 164.625 ;
        RECT 82.140 165.270 82.460 165.600 ;
        RECT 82.640 165.385 83.300 165.865 ;
        RECT 83.500 165.475 84.350 165.645 ;
        RECT 82.140 164.375 82.330 165.270 ;
        RECT 82.650 164.945 83.310 165.215 ;
        RECT 82.980 164.885 83.310 164.945 ;
        RECT 82.500 164.715 82.830 164.775 ;
        RECT 83.500 164.715 83.670 165.475 ;
        RECT 84.910 165.405 85.230 165.865 ;
        RECT 85.430 165.225 85.680 165.655 ;
        RECT 85.970 165.425 86.380 165.865 ;
        RECT 86.550 165.485 87.565 165.685 ;
        RECT 83.840 165.055 85.090 165.225 ;
        RECT 83.840 164.935 84.170 165.055 ;
        RECT 82.500 164.545 84.400 164.715 ;
        RECT 82.140 164.205 84.060 164.375 ;
        RECT 82.140 164.185 82.460 164.205 ;
        RECT 81.690 163.525 82.020 164.035 ;
        RECT 82.290 163.575 82.460 164.185 ;
        RECT 84.230 164.035 84.400 164.545 ;
        RECT 84.570 164.475 84.750 164.885 ;
        RECT 84.920 164.295 85.090 165.055 ;
        RECT 82.630 163.315 82.960 164.005 ;
        RECT 83.190 163.865 84.400 164.035 ;
        RECT 84.570 163.985 85.090 164.295 ;
        RECT 85.260 164.885 85.680 165.225 ;
        RECT 85.970 164.885 86.380 165.215 ;
        RECT 85.260 164.115 85.450 164.885 ;
        RECT 86.550 164.755 86.720 165.485 ;
        RECT 87.865 165.315 88.035 165.645 ;
        RECT 88.205 165.485 88.535 165.865 ;
        RECT 86.890 164.935 87.240 165.305 ;
        RECT 86.550 164.715 86.970 164.755 ;
        RECT 85.620 164.545 86.970 164.715 ;
        RECT 85.620 164.385 85.870 164.545 ;
        RECT 86.380 164.115 86.630 164.375 ;
        RECT 85.260 163.865 86.630 164.115 ;
        RECT 83.190 163.575 83.430 163.865 ;
        RECT 84.230 163.785 84.400 163.865 ;
        RECT 83.630 163.315 84.050 163.695 ;
        RECT 84.230 163.535 84.860 163.785 ;
        RECT 85.330 163.315 85.660 163.695 ;
        RECT 85.830 163.575 86.000 163.865 ;
        RECT 86.800 163.700 86.970 164.545 ;
        RECT 87.420 164.375 87.640 165.245 ;
        RECT 87.865 165.125 88.560 165.315 ;
        RECT 87.140 163.995 87.640 164.375 ;
        RECT 87.810 164.325 88.220 164.945 ;
        RECT 88.390 164.155 88.560 165.125 ;
        RECT 87.865 163.985 88.560 164.155 ;
        RECT 86.180 163.315 86.560 163.695 ;
        RECT 86.800 163.530 87.630 163.700 ;
        RECT 87.865 163.485 88.035 163.985 ;
        RECT 88.205 163.315 88.535 163.815 ;
        RECT 88.750 163.485 88.975 165.605 ;
        RECT 89.145 165.485 89.475 165.865 ;
        RECT 89.645 165.315 89.815 165.605 ;
        RECT 89.150 165.145 89.815 165.315 ;
        RECT 89.150 164.155 89.380 165.145 ;
        RECT 90.280 165.085 90.780 165.695 ;
        RECT 89.550 164.325 89.900 164.975 ;
        RECT 90.075 164.625 90.425 164.875 ;
        RECT 90.610 164.455 90.780 165.085 ;
        RECT 91.410 165.215 91.740 165.695 ;
        RECT 91.910 165.405 92.135 165.865 ;
        RECT 92.305 165.215 92.635 165.695 ;
        RECT 91.410 165.045 92.635 165.215 ;
        RECT 92.825 165.065 93.075 165.865 ;
        RECT 93.245 165.065 93.585 165.695 ;
        RECT 93.960 165.085 94.460 165.695 ;
        RECT 90.950 164.675 91.280 164.875 ;
        RECT 91.450 164.675 91.780 164.875 ;
        RECT 91.950 164.675 92.370 164.875 ;
        RECT 92.545 164.705 93.240 164.875 ;
        RECT 92.545 164.455 92.715 164.705 ;
        RECT 93.410 164.455 93.585 165.065 ;
        RECT 93.755 164.625 94.105 164.875 ;
        RECT 94.290 164.455 94.460 165.085 ;
        RECT 95.090 165.215 95.420 165.695 ;
        RECT 95.590 165.405 95.815 165.865 ;
        RECT 95.985 165.215 96.315 165.695 ;
        RECT 95.090 165.045 96.315 165.215 ;
        RECT 96.505 165.065 96.755 165.865 ;
        RECT 96.925 165.065 97.265 165.695 ;
        RECT 94.630 164.675 94.960 164.875 ;
        RECT 95.130 164.675 95.460 164.875 ;
        RECT 95.630 164.675 96.050 164.875 ;
        RECT 96.225 164.705 96.920 164.875 ;
        RECT 96.225 164.455 96.395 164.705 ;
        RECT 97.090 164.455 97.265 165.065 ;
        RECT 90.280 164.285 92.715 164.455 ;
        RECT 89.150 163.985 89.815 164.155 ;
        RECT 89.145 163.315 89.475 163.815 ;
        RECT 89.645 163.485 89.815 163.985 ;
        RECT 90.280 163.485 90.610 164.285 ;
        RECT 90.780 163.315 91.110 164.115 ;
        RECT 91.410 163.485 91.740 164.285 ;
        RECT 92.385 163.315 92.635 164.115 ;
        RECT 92.905 163.315 93.075 164.455 ;
        RECT 93.245 163.485 93.585 164.455 ;
        RECT 93.960 164.285 96.395 164.455 ;
        RECT 93.960 163.485 94.290 164.285 ;
        RECT 94.460 163.315 94.790 164.115 ;
        RECT 95.090 163.485 95.420 164.285 ;
        RECT 96.065 163.315 96.315 164.115 ;
        RECT 96.585 163.315 96.755 164.455 ;
        RECT 96.925 163.485 97.265 164.455 ;
        RECT 97.435 165.190 97.695 165.695 ;
        RECT 97.875 165.485 98.205 165.865 ;
        RECT 98.385 165.315 98.555 165.695 ;
        RECT 97.435 164.390 97.605 165.190 ;
        RECT 97.890 165.145 98.555 165.315 ;
        RECT 98.905 165.315 99.075 165.695 ;
        RECT 99.255 165.485 99.585 165.865 ;
        RECT 98.905 165.145 99.570 165.315 ;
        RECT 99.765 165.190 100.025 165.695 ;
        RECT 97.890 164.890 98.060 165.145 ;
        RECT 97.775 164.560 98.060 164.890 ;
        RECT 98.295 164.595 98.625 164.965 ;
        RECT 98.835 164.595 99.165 164.965 ;
        RECT 99.400 164.890 99.570 165.145 ;
        RECT 97.890 164.415 98.060 164.560 ;
        RECT 99.400 164.560 99.685 164.890 ;
        RECT 99.400 164.415 99.570 164.560 ;
        RECT 97.435 163.485 97.705 164.390 ;
        RECT 97.890 164.245 98.555 164.415 ;
        RECT 97.875 163.315 98.205 164.075 ;
        RECT 98.385 163.485 98.555 164.245 ;
        RECT 98.905 164.245 99.570 164.415 ;
        RECT 99.855 164.390 100.025 165.190 ;
        RECT 100.195 165.140 100.485 165.865 ;
        RECT 101.155 165.045 101.385 165.865 ;
        RECT 101.555 165.065 101.885 165.695 ;
        RECT 101.135 164.625 101.465 164.875 ;
        RECT 98.905 163.485 99.075 164.245 ;
        RECT 99.255 163.315 99.585 164.075 ;
        RECT 99.755 163.485 100.025 164.390 ;
        RECT 100.195 163.315 100.485 164.480 ;
        RECT 101.635 164.465 101.885 165.065 ;
        RECT 102.055 165.045 102.265 165.865 ;
        RECT 102.500 165.155 102.755 165.685 ;
        RECT 102.925 165.405 103.230 165.865 ;
        RECT 103.475 165.485 104.545 165.655 ;
        RECT 101.155 163.315 101.385 164.455 ;
        RECT 101.555 163.485 101.885 164.465 ;
        RECT 102.500 164.505 102.710 165.155 ;
        RECT 103.475 165.130 103.795 165.485 ;
        RECT 103.470 164.955 103.795 165.130 ;
        RECT 102.880 164.655 103.795 164.955 ;
        RECT 103.965 164.915 104.205 165.315 ;
        RECT 104.375 165.255 104.545 165.485 ;
        RECT 104.715 165.425 104.905 165.865 ;
        RECT 105.075 165.415 106.025 165.695 ;
        RECT 106.245 165.505 106.595 165.675 ;
        RECT 104.375 165.085 104.905 165.255 ;
        RECT 102.880 164.625 103.620 164.655 ;
        RECT 102.055 163.315 102.265 164.455 ;
        RECT 102.500 163.625 102.755 164.505 ;
        RECT 102.925 163.315 103.230 164.455 ;
        RECT 103.450 164.035 103.620 164.625 ;
        RECT 103.965 164.545 104.505 164.915 ;
        RECT 104.685 164.805 104.905 165.085 ;
        RECT 105.075 164.635 105.245 165.415 ;
        RECT 104.840 164.465 105.245 164.635 ;
        RECT 105.415 164.625 105.765 165.245 ;
        RECT 104.840 164.375 105.010 164.465 ;
        RECT 105.935 164.455 106.145 165.245 ;
        RECT 103.790 164.205 105.010 164.375 ;
        RECT 105.470 164.295 106.145 164.455 ;
        RECT 103.450 163.865 104.250 164.035 ;
        RECT 103.570 163.315 103.900 163.695 ;
        RECT 104.080 163.575 104.250 163.865 ;
        RECT 104.840 163.825 105.010 164.205 ;
        RECT 105.180 164.285 106.145 164.295 ;
        RECT 106.335 165.115 106.595 165.505 ;
        RECT 106.805 165.405 107.135 165.865 ;
        RECT 108.010 165.475 108.865 165.645 ;
        RECT 109.070 165.475 109.565 165.645 ;
        RECT 109.735 165.505 110.065 165.865 ;
        RECT 106.335 164.425 106.505 165.115 ;
        RECT 106.675 164.765 106.845 164.945 ;
        RECT 107.015 164.935 107.805 165.185 ;
        RECT 108.010 164.765 108.180 165.475 ;
        RECT 108.350 164.965 108.705 165.185 ;
        RECT 106.675 164.595 108.365 164.765 ;
        RECT 105.180 163.995 105.640 164.285 ;
        RECT 106.335 164.255 107.835 164.425 ;
        RECT 106.335 164.115 106.505 164.255 ;
        RECT 105.945 163.945 106.505 164.115 ;
        RECT 104.420 163.315 104.670 163.775 ;
        RECT 104.840 163.485 105.710 163.825 ;
        RECT 105.945 163.485 106.115 163.945 ;
        RECT 106.950 163.915 108.025 164.085 ;
        RECT 106.285 163.315 106.655 163.775 ;
        RECT 106.950 163.575 107.120 163.915 ;
        RECT 107.290 163.315 107.620 163.745 ;
        RECT 107.855 163.575 108.025 163.915 ;
        RECT 108.195 163.815 108.365 164.595 ;
        RECT 108.535 164.375 108.705 164.965 ;
        RECT 108.875 164.565 109.225 165.185 ;
        RECT 108.535 163.985 109.000 164.375 ;
        RECT 109.395 164.115 109.565 165.475 ;
        RECT 109.735 164.285 110.195 165.335 ;
        RECT 109.170 163.945 109.565 164.115 ;
        RECT 109.170 163.815 109.340 163.945 ;
        RECT 108.195 163.485 108.875 163.815 ;
        RECT 109.090 163.485 109.340 163.815 ;
        RECT 109.510 163.315 109.760 163.775 ;
        RECT 109.930 163.500 110.255 164.285 ;
        RECT 110.425 163.485 110.595 165.605 ;
        RECT 110.765 165.485 111.095 165.865 ;
        RECT 111.265 165.315 111.520 165.605 ;
        RECT 110.770 165.145 111.520 165.315 ;
        RECT 110.770 164.155 111.000 165.145 ;
        RECT 112.155 165.115 113.365 165.865 ;
        RECT 111.170 164.325 111.520 164.975 ;
        RECT 112.155 164.405 112.675 164.945 ;
        RECT 112.845 164.575 113.365 165.115 ;
        RECT 110.770 163.985 111.520 164.155 ;
        RECT 110.765 163.315 111.095 163.815 ;
        RECT 111.265 163.485 111.520 163.985 ;
        RECT 112.155 163.315 113.365 164.405 ;
        RECT 22.830 163.145 113.450 163.315 ;
        RECT 22.915 162.055 24.125 163.145 ;
        RECT 22.915 161.345 23.435 161.885 ;
        RECT 23.605 161.515 24.125 162.055 ;
        RECT 24.670 162.165 24.925 162.835 ;
        RECT 25.105 162.345 25.390 163.145 ;
        RECT 25.570 162.425 25.900 162.935 ;
        RECT 22.915 160.595 24.125 161.345 ;
        RECT 24.670 161.305 24.850 162.165 ;
        RECT 25.570 161.835 25.820 162.425 ;
        RECT 26.170 162.275 26.340 162.885 ;
        RECT 26.510 162.455 26.840 163.145 ;
        RECT 27.070 162.595 27.310 162.885 ;
        RECT 27.510 162.765 27.930 163.145 ;
        RECT 28.110 162.675 28.740 162.925 ;
        RECT 29.210 162.765 29.540 163.145 ;
        RECT 28.110 162.595 28.280 162.675 ;
        RECT 29.710 162.595 29.880 162.885 ;
        RECT 30.060 162.765 30.440 163.145 ;
        RECT 30.680 162.760 31.510 162.930 ;
        RECT 27.070 162.425 28.280 162.595 ;
        RECT 25.020 161.505 25.820 161.835 ;
        RECT 24.670 161.105 24.925 161.305 ;
        RECT 24.585 160.935 24.925 161.105 ;
        RECT 24.670 160.775 24.925 160.935 ;
        RECT 25.105 160.595 25.390 161.055 ;
        RECT 25.570 160.855 25.820 161.505 ;
        RECT 26.020 162.255 26.340 162.275 ;
        RECT 26.020 162.085 27.940 162.255 ;
        RECT 26.020 161.190 26.210 162.085 ;
        RECT 28.110 161.915 28.280 162.425 ;
        RECT 28.450 162.165 28.970 162.475 ;
        RECT 26.380 161.745 28.280 161.915 ;
        RECT 26.380 161.685 26.710 161.745 ;
        RECT 26.860 161.515 27.190 161.575 ;
        RECT 26.530 161.245 27.190 161.515 ;
        RECT 26.020 160.860 26.340 161.190 ;
        RECT 26.520 160.595 27.180 161.075 ;
        RECT 27.380 160.985 27.550 161.745 ;
        RECT 28.450 161.575 28.630 161.985 ;
        RECT 27.720 161.405 28.050 161.525 ;
        RECT 28.800 161.405 28.970 162.165 ;
        RECT 27.720 161.235 28.970 161.405 ;
        RECT 29.140 162.345 30.510 162.595 ;
        RECT 29.140 161.575 29.330 162.345 ;
        RECT 30.260 162.085 30.510 162.345 ;
        RECT 29.500 161.915 29.750 162.075 ;
        RECT 30.680 161.915 30.850 162.760 ;
        RECT 31.745 162.475 31.915 162.975 ;
        RECT 32.085 162.645 32.415 163.145 ;
        RECT 31.020 162.085 31.520 162.465 ;
        RECT 31.745 162.305 32.440 162.475 ;
        RECT 29.500 161.745 30.850 161.915 ;
        RECT 30.430 161.705 30.850 161.745 ;
        RECT 29.140 161.235 29.560 161.575 ;
        RECT 29.850 161.245 30.260 161.575 ;
        RECT 27.380 160.815 28.230 160.985 ;
        RECT 28.790 160.595 29.110 161.055 ;
        RECT 29.310 160.805 29.560 161.235 ;
        RECT 29.850 160.595 30.260 161.035 ;
        RECT 30.430 160.975 30.600 161.705 ;
        RECT 30.770 161.155 31.120 161.525 ;
        RECT 31.300 161.215 31.520 162.085 ;
        RECT 31.690 161.515 32.100 162.135 ;
        RECT 32.270 161.335 32.440 162.305 ;
        RECT 31.745 161.145 32.440 161.335 ;
        RECT 30.430 160.775 31.445 160.975 ;
        RECT 31.745 160.815 31.915 161.145 ;
        RECT 32.085 160.595 32.415 160.975 ;
        RECT 32.630 160.855 32.855 162.975 ;
        RECT 33.025 162.645 33.355 163.145 ;
        RECT 33.525 162.475 33.695 162.975 ;
        RECT 33.030 162.305 33.695 162.475 ;
        RECT 33.030 161.315 33.260 162.305 ;
        RECT 33.430 161.485 33.780 162.135 ;
        RECT 33.955 162.070 34.225 162.975 ;
        RECT 34.395 162.385 34.725 163.145 ;
        RECT 34.905 162.215 35.075 162.975 ;
        RECT 33.030 161.145 33.695 161.315 ;
        RECT 33.025 160.595 33.355 160.975 ;
        RECT 33.525 160.855 33.695 161.145 ;
        RECT 33.955 161.270 34.125 162.070 ;
        RECT 34.410 162.045 35.075 162.215 ;
        RECT 34.410 161.900 34.580 162.045 ;
        RECT 35.795 161.980 36.085 163.145 ;
        RECT 36.315 162.005 36.525 163.145 ;
        RECT 36.695 161.995 37.025 162.975 ;
        RECT 37.195 162.005 37.425 163.145 ;
        RECT 37.635 162.070 37.905 162.975 ;
        RECT 38.075 162.385 38.405 163.145 ;
        RECT 38.585 162.215 38.755 162.975 ;
        RECT 39.390 162.805 39.645 162.835 ;
        RECT 39.305 162.635 39.645 162.805 ;
        RECT 34.295 161.570 34.580 161.900 ;
        RECT 34.410 161.315 34.580 161.570 ;
        RECT 34.815 161.495 35.145 161.865 ;
        RECT 33.955 160.765 34.215 161.270 ;
        RECT 34.410 161.145 35.075 161.315 ;
        RECT 34.395 160.595 34.725 160.975 ;
        RECT 34.905 160.765 35.075 161.145 ;
        RECT 35.795 160.595 36.085 161.320 ;
        RECT 36.315 160.595 36.525 161.415 ;
        RECT 36.695 161.395 36.945 161.995 ;
        RECT 37.115 161.585 37.445 161.835 ;
        RECT 36.695 160.765 37.025 161.395 ;
        RECT 37.195 160.595 37.425 161.415 ;
        RECT 37.635 161.270 37.805 162.070 ;
        RECT 38.090 162.045 38.755 162.215 ;
        RECT 39.390 162.165 39.645 162.635 ;
        RECT 39.825 162.345 40.110 163.145 ;
        RECT 40.290 162.425 40.620 162.935 ;
        RECT 38.090 161.900 38.260 162.045 ;
        RECT 37.975 161.570 38.260 161.900 ;
        RECT 38.090 161.315 38.260 161.570 ;
        RECT 38.495 161.495 38.825 161.865 ;
        RECT 37.635 160.765 37.895 161.270 ;
        RECT 38.090 161.145 38.755 161.315 ;
        RECT 38.075 160.595 38.405 160.975 ;
        RECT 38.585 160.765 38.755 161.145 ;
        RECT 39.390 161.305 39.570 162.165 ;
        RECT 40.290 161.835 40.540 162.425 ;
        RECT 40.890 162.275 41.060 162.885 ;
        RECT 41.230 162.455 41.560 163.145 ;
        RECT 41.790 162.595 42.030 162.885 ;
        RECT 42.230 162.765 42.650 163.145 ;
        RECT 42.830 162.675 43.460 162.925 ;
        RECT 43.930 162.765 44.260 163.145 ;
        RECT 42.830 162.595 43.000 162.675 ;
        RECT 44.430 162.595 44.600 162.885 ;
        RECT 44.780 162.765 45.160 163.145 ;
        RECT 45.400 162.760 46.230 162.930 ;
        RECT 41.790 162.425 43.000 162.595 ;
        RECT 39.740 161.505 40.540 161.835 ;
        RECT 39.390 160.775 39.645 161.305 ;
        RECT 39.825 160.595 40.110 161.055 ;
        RECT 40.290 160.855 40.540 161.505 ;
        RECT 40.740 162.255 41.060 162.275 ;
        RECT 40.740 162.085 42.660 162.255 ;
        RECT 40.740 161.190 40.930 162.085 ;
        RECT 42.830 161.915 43.000 162.425 ;
        RECT 43.170 162.165 43.690 162.475 ;
        RECT 41.100 161.745 43.000 161.915 ;
        RECT 41.100 161.685 41.430 161.745 ;
        RECT 41.580 161.515 41.910 161.575 ;
        RECT 41.250 161.245 41.910 161.515 ;
        RECT 40.740 160.860 41.060 161.190 ;
        RECT 41.240 160.595 41.900 161.075 ;
        RECT 42.100 160.985 42.270 161.745 ;
        RECT 43.170 161.575 43.350 161.985 ;
        RECT 42.440 161.405 42.770 161.525 ;
        RECT 43.520 161.405 43.690 162.165 ;
        RECT 42.440 161.235 43.690 161.405 ;
        RECT 43.860 162.345 45.230 162.595 ;
        RECT 43.860 161.575 44.050 162.345 ;
        RECT 44.980 162.085 45.230 162.345 ;
        RECT 44.220 161.915 44.470 162.075 ;
        RECT 45.400 161.915 45.570 162.760 ;
        RECT 46.465 162.475 46.635 162.975 ;
        RECT 46.805 162.645 47.135 163.145 ;
        RECT 45.740 162.085 46.240 162.465 ;
        RECT 46.465 162.305 47.160 162.475 ;
        RECT 44.220 161.745 45.570 161.915 ;
        RECT 45.150 161.705 45.570 161.745 ;
        RECT 43.860 161.235 44.280 161.575 ;
        RECT 44.570 161.245 44.980 161.575 ;
        RECT 42.100 160.815 42.950 160.985 ;
        RECT 43.510 160.595 43.830 161.055 ;
        RECT 44.030 160.805 44.280 161.235 ;
        RECT 44.570 160.595 44.980 161.035 ;
        RECT 45.150 160.975 45.320 161.705 ;
        RECT 45.490 161.155 45.840 161.525 ;
        RECT 46.020 161.215 46.240 162.085 ;
        RECT 46.410 161.515 46.820 162.135 ;
        RECT 46.990 161.335 47.160 162.305 ;
        RECT 46.465 161.145 47.160 161.335 ;
        RECT 45.150 160.775 46.165 160.975 ;
        RECT 46.465 160.815 46.635 161.145 ;
        RECT 46.805 160.595 47.135 160.975 ;
        RECT 47.350 160.855 47.575 162.975 ;
        RECT 47.745 162.645 48.075 163.145 ;
        RECT 48.245 162.475 48.415 162.975 ;
        RECT 47.750 162.305 48.415 162.475 ;
        RECT 47.750 161.315 47.980 162.305 ;
        RECT 48.150 161.485 48.500 162.135 ;
        RECT 48.680 162.005 49.015 162.975 ;
        RECT 49.185 162.005 49.355 163.145 ;
        RECT 49.525 162.805 51.555 162.975 ;
        RECT 48.680 161.335 48.850 162.005 ;
        RECT 49.525 161.835 49.695 162.805 ;
        RECT 49.020 161.505 49.275 161.835 ;
        RECT 49.500 161.505 49.695 161.835 ;
        RECT 49.865 162.465 50.990 162.635 ;
        RECT 49.105 161.335 49.275 161.505 ;
        RECT 49.865 161.335 50.035 162.465 ;
        RECT 47.750 161.145 48.415 161.315 ;
        RECT 47.745 160.595 48.075 160.975 ;
        RECT 48.245 160.855 48.415 161.145 ;
        RECT 48.680 160.765 48.935 161.335 ;
        RECT 49.105 161.165 50.035 161.335 ;
        RECT 50.205 162.125 51.215 162.295 ;
        RECT 50.205 161.325 50.375 162.125 ;
        RECT 50.580 161.785 50.855 161.925 ;
        RECT 50.575 161.615 50.855 161.785 ;
        RECT 49.860 161.130 50.035 161.165 ;
        RECT 49.105 160.595 49.435 160.995 ;
        RECT 49.860 160.765 50.390 161.130 ;
        RECT 50.580 160.765 50.855 161.615 ;
        RECT 51.025 160.765 51.215 162.125 ;
        RECT 51.385 162.140 51.555 162.805 ;
        RECT 51.725 162.385 51.895 163.145 ;
        RECT 52.130 162.385 52.645 162.795 ;
        RECT 51.385 161.950 52.135 162.140 ;
        RECT 52.305 161.575 52.645 162.385 ;
        RECT 53.850 162.515 54.135 162.975 ;
        RECT 54.305 162.685 54.575 163.145 ;
        RECT 53.850 162.295 54.805 162.515 ;
        RECT 51.415 161.405 52.645 161.575 ;
        RECT 53.735 161.565 54.425 162.125 ;
        RECT 51.395 160.595 51.905 161.130 ;
        RECT 52.125 160.800 52.370 161.405 ;
        RECT 54.595 161.395 54.805 162.295 ;
        RECT 53.850 161.225 54.805 161.395 ;
        RECT 54.975 162.125 55.375 162.975 ;
        RECT 55.565 162.515 55.845 162.975 ;
        RECT 56.365 162.685 56.690 163.145 ;
        RECT 55.565 162.295 56.690 162.515 ;
        RECT 54.975 161.565 56.070 162.125 ;
        RECT 56.240 161.835 56.690 162.295 ;
        RECT 56.860 162.005 57.245 162.975 ;
        RECT 53.850 160.765 54.135 161.225 ;
        RECT 54.305 160.595 54.575 161.055 ;
        RECT 54.975 160.765 55.375 161.565 ;
        RECT 56.240 161.505 56.795 161.835 ;
        RECT 56.240 161.395 56.690 161.505 ;
        RECT 55.565 161.225 56.690 161.395 ;
        RECT 56.965 161.335 57.245 162.005 ;
        RECT 55.565 160.765 55.845 161.225 ;
        RECT 56.365 160.595 56.690 161.055 ;
        RECT 56.860 160.765 57.245 161.335 ;
        RECT 57.420 162.005 57.755 162.975 ;
        RECT 57.925 162.005 58.095 163.145 ;
        RECT 58.265 162.805 60.295 162.975 ;
        RECT 57.420 161.335 57.590 162.005 ;
        RECT 58.265 161.835 58.435 162.805 ;
        RECT 57.760 161.505 58.015 161.835 ;
        RECT 58.240 161.505 58.435 161.835 ;
        RECT 58.605 162.465 59.730 162.635 ;
        RECT 57.845 161.335 58.015 161.505 ;
        RECT 58.605 161.335 58.775 162.465 ;
        RECT 57.420 160.765 57.675 161.335 ;
        RECT 57.845 161.165 58.775 161.335 ;
        RECT 58.945 162.125 59.955 162.295 ;
        RECT 58.945 161.325 59.115 162.125 ;
        RECT 59.320 161.785 59.595 161.925 ;
        RECT 59.315 161.615 59.595 161.785 ;
        RECT 58.600 161.130 58.775 161.165 ;
        RECT 57.845 160.595 58.175 160.995 ;
        RECT 58.600 160.765 59.130 161.130 ;
        RECT 59.320 160.765 59.595 161.615 ;
        RECT 59.765 160.765 59.955 162.125 ;
        RECT 60.125 162.140 60.295 162.805 ;
        RECT 60.465 162.385 60.635 163.145 ;
        RECT 60.870 162.385 61.385 162.795 ;
        RECT 60.125 161.950 60.875 162.140 ;
        RECT 61.045 161.575 61.385 162.385 ;
        RECT 61.555 161.980 61.845 163.145 ;
        RECT 62.015 162.005 62.355 162.975 ;
        RECT 62.525 162.005 62.695 163.145 ;
        RECT 62.965 162.345 63.215 163.145 ;
        RECT 63.860 162.175 64.190 162.975 ;
        RECT 64.490 162.345 64.820 163.145 ;
        RECT 64.990 162.175 65.320 162.975 ;
        RECT 62.885 162.005 65.320 162.175 ;
        RECT 65.785 162.215 65.955 162.975 ;
        RECT 66.135 162.385 66.465 163.145 ;
        RECT 65.785 162.045 66.450 162.215 ;
        RECT 66.635 162.070 66.905 162.975 ;
        RECT 60.155 161.405 61.385 161.575 ;
        RECT 60.135 160.595 60.645 161.130 ;
        RECT 60.865 160.800 61.110 161.405 ;
        RECT 62.015 161.395 62.190 162.005 ;
        RECT 62.885 161.755 63.055 162.005 ;
        RECT 62.360 161.585 63.055 161.755 ;
        RECT 63.230 161.585 63.650 161.785 ;
        RECT 63.820 161.585 64.150 161.785 ;
        RECT 64.320 161.585 64.650 161.785 ;
        RECT 61.555 160.595 61.845 161.320 ;
        RECT 62.015 160.765 62.355 161.395 ;
        RECT 62.525 160.595 62.775 161.395 ;
        RECT 62.965 161.245 64.190 161.415 ;
        RECT 62.965 160.765 63.295 161.245 ;
        RECT 63.465 160.595 63.690 161.055 ;
        RECT 63.860 160.765 64.190 161.245 ;
        RECT 64.820 161.375 64.990 162.005 ;
        RECT 66.280 161.900 66.450 162.045 ;
        RECT 65.175 161.585 65.525 161.835 ;
        RECT 65.715 161.495 66.045 161.865 ;
        RECT 66.280 161.570 66.565 161.900 ;
        RECT 64.820 160.765 65.320 161.375 ;
        RECT 66.280 161.315 66.450 161.570 ;
        RECT 65.785 161.145 66.450 161.315 ;
        RECT 66.735 161.270 66.905 162.070 ;
        RECT 67.280 162.175 67.610 162.975 ;
        RECT 67.780 162.345 68.110 163.145 ;
        RECT 68.410 162.175 68.740 162.975 ;
        RECT 69.385 162.345 69.635 163.145 ;
        RECT 67.280 162.005 69.715 162.175 ;
        RECT 69.905 162.005 70.075 163.145 ;
        RECT 70.245 162.005 70.585 162.975 ;
        RECT 67.075 161.585 67.425 161.835 ;
        RECT 67.610 161.375 67.780 162.005 ;
        RECT 67.950 161.585 68.280 161.785 ;
        RECT 68.450 161.585 68.780 161.785 ;
        RECT 68.950 161.585 69.370 161.785 ;
        RECT 69.545 161.755 69.715 162.005 ;
        RECT 69.545 161.585 70.240 161.755 ;
        RECT 65.785 160.765 65.955 161.145 ;
        RECT 66.135 160.595 66.465 160.975 ;
        RECT 66.645 160.765 66.905 161.270 ;
        RECT 67.280 160.765 67.780 161.375 ;
        RECT 68.410 161.245 69.635 161.415 ;
        RECT 70.410 161.395 70.585 162.005 ;
        RECT 68.410 160.765 68.740 161.245 ;
        RECT 68.910 160.595 69.135 161.055 ;
        RECT 69.305 160.765 69.635 161.245 ;
        RECT 69.825 160.595 70.075 161.395 ;
        RECT 70.245 160.765 70.585 161.395 ;
        RECT 70.755 162.005 71.095 162.975 ;
        RECT 71.265 162.005 71.435 163.145 ;
        RECT 71.705 162.345 71.955 163.145 ;
        RECT 72.600 162.175 72.930 162.975 ;
        RECT 73.230 162.345 73.560 163.145 ;
        RECT 73.730 162.175 74.060 162.975 ;
        RECT 71.625 162.005 74.060 162.175 ;
        RECT 74.810 162.165 75.065 162.835 ;
        RECT 75.245 162.345 75.530 163.145 ;
        RECT 75.710 162.425 76.040 162.935 ;
        RECT 74.810 162.125 74.990 162.165 ;
        RECT 70.755 161.395 70.930 162.005 ;
        RECT 71.625 161.755 71.795 162.005 ;
        RECT 71.100 161.585 71.795 161.755 ;
        RECT 71.970 161.585 72.390 161.785 ;
        RECT 72.560 161.585 72.890 161.785 ;
        RECT 73.060 161.585 73.390 161.785 ;
        RECT 70.755 160.765 71.095 161.395 ;
        RECT 71.265 160.595 71.515 161.395 ;
        RECT 71.705 161.245 72.930 161.415 ;
        RECT 71.705 160.765 72.035 161.245 ;
        RECT 72.205 160.595 72.430 161.055 ;
        RECT 72.600 160.765 72.930 161.245 ;
        RECT 73.560 161.375 73.730 162.005 ;
        RECT 74.725 161.955 74.990 162.125 ;
        RECT 73.915 161.585 74.265 161.835 ;
        RECT 73.560 160.765 74.060 161.375 ;
        RECT 74.810 161.305 74.990 161.955 ;
        RECT 75.710 161.835 75.960 162.425 ;
        RECT 76.310 162.275 76.480 162.885 ;
        RECT 76.650 162.455 76.980 163.145 ;
        RECT 77.210 162.595 77.450 162.885 ;
        RECT 77.650 162.765 78.070 163.145 ;
        RECT 78.250 162.675 78.880 162.925 ;
        RECT 79.350 162.765 79.680 163.145 ;
        RECT 78.250 162.595 78.420 162.675 ;
        RECT 79.850 162.595 80.020 162.885 ;
        RECT 80.200 162.765 80.580 163.145 ;
        RECT 80.820 162.760 81.650 162.930 ;
        RECT 77.210 162.425 78.420 162.595 ;
        RECT 75.160 161.505 75.960 161.835 ;
        RECT 74.810 160.775 75.065 161.305 ;
        RECT 75.245 160.595 75.530 161.055 ;
        RECT 75.710 160.855 75.960 161.505 ;
        RECT 76.160 162.255 76.480 162.275 ;
        RECT 76.160 162.085 78.080 162.255 ;
        RECT 76.160 161.190 76.350 162.085 ;
        RECT 78.250 161.915 78.420 162.425 ;
        RECT 78.590 162.165 79.110 162.475 ;
        RECT 76.520 161.745 78.420 161.915 ;
        RECT 76.520 161.685 76.850 161.745 ;
        RECT 77.000 161.515 77.330 161.575 ;
        RECT 76.670 161.245 77.330 161.515 ;
        RECT 76.160 160.860 76.480 161.190 ;
        RECT 76.660 160.595 77.320 161.075 ;
        RECT 77.520 160.985 77.690 161.745 ;
        RECT 78.590 161.575 78.770 161.985 ;
        RECT 77.860 161.405 78.190 161.525 ;
        RECT 78.940 161.405 79.110 162.165 ;
        RECT 77.860 161.235 79.110 161.405 ;
        RECT 79.280 162.345 80.650 162.595 ;
        RECT 79.280 161.575 79.470 162.345 ;
        RECT 80.400 162.085 80.650 162.345 ;
        RECT 79.640 161.915 79.890 162.075 ;
        RECT 80.820 161.915 80.990 162.760 ;
        RECT 81.885 162.475 82.055 162.975 ;
        RECT 82.225 162.645 82.555 163.145 ;
        RECT 81.160 162.085 81.660 162.465 ;
        RECT 81.885 162.305 82.580 162.475 ;
        RECT 79.640 161.745 80.990 161.915 ;
        RECT 80.570 161.705 80.990 161.745 ;
        RECT 79.280 161.235 79.700 161.575 ;
        RECT 79.990 161.245 80.400 161.575 ;
        RECT 77.520 160.815 78.370 160.985 ;
        RECT 78.930 160.595 79.250 161.055 ;
        RECT 79.450 160.805 79.700 161.235 ;
        RECT 79.990 160.595 80.400 161.035 ;
        RECT 80.570 160.975 80.740 161.705 ;
        RECT 80.910 161.155 81.260 161.525 ;
        RECT 81.440 161.215 81.660 162.085 ;
        RECT 81.830 161.515 82.240 162.135 ;
        RECT 82.410 161.335 82.580 162.305 ;
        RECT 81.885 161.145 82.580 161.335 ;
        RECT 80.570 160.775 81.585 160.975 ;
        RECT 81.885 160.815 82.055 161.145 ;
        RECT 82.225 160.595 82.555 160.975 ;
        RECT 82.770 160.855 82.995 162.975 ;
        RECT 83.165 162.645 83.495 163.145 ;
        RECT 83.665 162.475 83.835 162.975 ;
        RECT 83.170 162.305 83.835 162.475 ;
        RECT 83.170 161.315 83.400 162.305 ;
        RECT 83.570 161.485 83.920 162.135 ;
        RECT 84.155 162.005 84.365 163.145 ;
        RECT 84.535 161.995 84.865 162.975 ;
        RECT 85.035 162.005 85.265 163.145 ;
        RECT 86.025 162.215 86.195 162.975 ;
        RECT 86.375 162.385 86.705 163.145 ;
        RECT 86.025 162.045 86.690 162.215 ;
        RECT 86.875 162.070 87.145 162.975 ;
        RECT 83.170 161.145 83.835 161.315 ;
        RECT 83.165 160.595 83.495 160.975 ;
        RECT 83.665 160.855 83.835 161.145 ;
        RECT 84.155 160.595 84.365 161.415 ;
        RECT 84.535 161.395 84.785 161.995 ;
        RECT 86.520 161.900 86.690 162.045 ;
        RECT 84.955 161.585 85.285 161.835 ;
        RECT 85.955 161.495 86.285 161.865 ;
        RECT 86.520 161.570 86.805 161.900 ;
        RECT 84.535 160.765 84.865 161.395 ;
        RECT 85.035 160.595 85.265 161.415 ;
        RECT 86.520 161.315 86.690 161.570 ;
        RECT 86.025 161.145 86.690 161.315 ;
        RECT 86.975 161.270 87.145 162.070 ;
        RECT 87.315 161.980 87.605 163.145 ;
        RECT 87.775 162.055 88.985 163.145 ;
        RECT 87.775 161.515 88.295 162.055 ;
        RECT 89.155 162.005 89.495 162.975 ;
        RECT 89.665 162.005 89.835 163.145 ;
        RECT 90.105 162.345 90.355 163.145 ;
        RECT 91.000 162.175 91.330 162.975 ;
        RECT 91.630 162.345 91.960 163.145 ;
        RECT 92.130 162.175 92.460 162.975 ;
        RECT 90.025 162.005 92.460 162.175 ;
        RECT 92.835 162.005 93.175 162.975 ;
        RECT 93.345 162.005 93.515 163.145 ;
        RECT 93.785 162.345 94.035 163.145 ;
        RECT 94.680 162.175 95.010 162.975 ;
        RECT 95.310 162.345 95.640 163.145 ;
        RECT 95.810 162.175 96.140 162.975 ;
        RECT 93.705 162.005 96.140 162.175 ;
        RECT 96.515 162.005 96.855 162.975 ;
        RECT 97.025 162.005 97.195 163.145 ;
        RECT 97.465 162.345 97.715 163.145 ;
        RECT 98.360 162.175 98.690 162.975 ;
        RECT 98.990 162.345 99.320 163.145 ;
        RECT 99.490 162.175 99.820 162.975 ;
        RECT 97.385 162.005 99.820 162.175 ;
        RECT 101.155 162.005 101.385 163.145 ;
        RECT 88.465 161.345 88.985 161.885 ;
        RECT 86.025 160.765 86.195 161.145 ;
        RECT 86.375 160.595 86.705 160.975 ;
        RECT 86.885 160.765 87.145 161.270 ;
        RECT 87.315 160.595 87.605 161.320 ;
        RECT 87.775 160.595 88.985 161.345 ;
        RECT 89.155 161.395 89.330 162.005 ;
        RECT 90.025 161.755 90.195 162.005 ;
        RECT 89.500 161.585 90.195 161.755 ;
        RECT 90.370 161.585 90.790 161.785 ;
        RECT 90.960 161.585 91.290 161.785 ;
        RECT 91.460 161.585 91.790 161.785 ;
        RECT 89.155 160.765 89.495 161.395 ;
        RECT 89.665 160.595 89.915 161.395 ;
        RECT 90.105 161.245 91.330 161.415 ;
        RECT 90.105 160.765 90.435 161.245 ;
        RECT 90.605 160.595 90.830 161.055 ;
        RECT 91.000 160.765 91.330 161.245 ;
        RECT 91.960 161.375 92.130 162.005 ;
        RECT 92.315 161.585 92.665 161.835 ;
        RECT 92.835 161.395 93.010 162.005 ;
        RECT 93.705 161.755 93.875 162.005 ;
        RECT 93.180 161.585 93.875 161.755 ;
        RECT 94.050 161.585 94.470 161.785 ;
        RECT 94.640 161.585 94.970 161.785 ;
        RECT 95.140 161.585 95.470 161.785 ;
        RECT 91.960 160.765 92.460 161.375 ;
        RECT 92.835 160.765 93.175 161.395 ;
        RECT 93.345 160.595 93.595 161.395 ;
        RECT 93.785 161.245 95.010 161.415 ;
        RECT 93.785 160.765 94.115 161.245 ;
        RECT 94.285 160.595 94.510 161.055 ;
        RECT 94.680 160.765 95.010 161.245 ;
        RECT 95.640 161.375 95.810 162.005 ;
        RECT 95.995 161.585 96.345 161.835 ;
        RECT 96.515 161.395 96.690 162.005 ;
        RECT 97.385 161.755 97.555 162.005 ;
        RECT 96.860 161.585 97.555 161.755 ;
        RECT 97.730 161.585 98.150 161.785 ;
        RECT 98.320 161.585 98.650 161.785 ;
        RECT 98.820 161.585 99.150 161.785 ;
        RECT 95.640 160.765 96.140 161.375 ;
        RECT 96.515 160.765 96.855 161.395 ;
        RECT 97.025 160.595 97.275 161.395 ;
        RECT 97.465 161.245 98.690 161.415 ;
        RECT 97.465 160.765 97.795 161.245 ;
        RECT 97.965 160.595 98.190 161.055 ;
        RECT 98.360 160.765 98.690 161.245 ;
        RECT 99.320 161.375 99.490 162.005 ;
        RECT 101.555 161.995 101.885 162.975 ;
        RECT 102.055 162.005 102.265 163.145 ;
        RECT 102.585 162.475 102.755 162.975 ;
        RECT 102.925 162.645 103.255 163.145 ;
        RECT 102.585 162.305 103.250 162.475 ;
        RECT 99.675 161.585 100.025 161.835 ;
        RECT 101.135 161.585 101.465 161.835 ;
        RECT 99.320 160.765 99.820 161.375 ;
        RECT 101.155 160.595 101.385 161.415 ;
        RECT 101.635 161.395 101.885 161.995 ;
        RECT 102.500 161.485 102.850 162.135 ;
        RECT 101.555 160.765 101.885 161.395 ;
        RECT 102.055 160.595 102.265 161.415 ;
        RECT 103.020 161.315 103.250 162.305 ;
        RECT 102.585 161.145 103.250 161.315 ;
        RECT 102.585 160.855 102.755 161.145 ;
        RECT 102.925 160.595 103.255 160.975 ;
        RECT 103.425 160.855 103.650 162.975 ;
        RECT 103.865 162.645 104.195 163.145 ;
        RECT 104.365 162.475 104.535 162.975 ;
        RECT 104.770 162.760 105.600 162.930 ;
        RECT 105.840 162.765 106.220 163.145 ;
        RECT 103.840 162.305 104.535 162.475 ;
        RECT 103.840 161.335 104.010 162.305 ;
        RECT 104.180 161.515 104.590 162.135 ;
        RECT 104.760 162.085 105.260 162.465 ;
        RECT 103.840 161.145 104.535 161.335 ;
        RECT 104.760 161.215 104.980 162.085 ;
        RECT 105.430 161.915 105.600 162.760 ;
        RECT 106.400 162.595 106.570 162.885 ;
        RECT 106.740 162.765 107.070 163.145 ;
        RECT 107.540 162.675 108.170 162.925 ;
        RECT 108.350 162.765 108.770 163.145 ;
        RECT 108.000 162.595 108.170 162.675 ;
        RECT 108.970 162.595 109.210 162.885 ;
        RECT 105.770 162.345 107.140 162.595 ;
        RECT 105.770 162.085 106.020 162.345 ;
        RECT 106.530 161.915 106.780 162.075 ;
        RECT 105.430 161.745 106.780 161.915 ;
        RECT 105.430 161.705 105.850 161.745 ;
        RECT 105.160 161.155 105.510 161.525 ;
        RECT 103.865 160.595 104.195 160.975 ;
        RECT 104.365 160.815 104.535 161.145 ;
        RECT 105.680 160.975 105.850 161.705 ;
        RECT 106.950 161.575 107.140 162.345 ;
        RECT 106.020 161.245 106.430 161.575 ;
        RECT 106.720 161.235 107.140 161.575 ;
        RECT 107.310 162.165 107.830 162.475 ;
        RECT 108.000 162.425 109.210 162.595 ;
        RECT 109.440 162.455 109.770 163.145 ;
        RECT 107.310 161.405 107.480 162.165 ;
        RECT 107.650 161.575 107.830 161.985 ;
        RECT 108.000 161.915 108.170 162.425 ;
        RECT 109.940 162.275 110.110 162.885 ;
        RECT 110.380 162.425 110.710 162.935 ;
        RECT 109.940 162.255 110.260 162.275 ;
        RECT 108.340 162.085 110.260 162.255 ;
        RECT 108.000 161.745 109.900 161.915 ;
        RECT 108.230 161.405 108.560 161.525 ;
        RECT 107.310 161.235 108.560 161.405 ;
        RECT 104.835 160.775 105.850 160.975 ;
        RECT 106.020 160.595 106.430 161.035 ;
        RECT 106.720 160.805 106.970 161.235 ;
        RECT 107.170 160.595 107.490 161.055 ;
        RECT 108.730 160.985 108.900 161.745 ;
        RECT 109.570 161.685 109.900 161.745 ;
        RECT 109.090 161.515 109.420 161.575 ;
        RECT 109.090 161.245 109.750 161.515 ;
        RECT 110.070 161.190 110.260 162.085 ;
        RECT 108.050 160.815 108.900 160.985 ;
        RECT 109.100 160.595 109.760 161.075 ;
        RECT 109.940 160.860 110.260 161.190 ;
        RECT 110.460 161.835 110.710 162.425 ;
        RECT 110.890 162.345 111.175 163.145 ;
        RECT 111.355 162.165 111.610 162.835 ;
        RECT 110.460 161.505 111.260 161.835 ;
        RECT 110.460 160.855 110.710 161.505 ;
        RECT 111.430 161.305 111.610 162.165 ;
        RECT 112.155 162.055 113.365 163.145 ;
        RECT 112.155 161.515 112.675 162.055 ;
        RECT 112.845 161.345 113.365 161.885 ;
        RECT 111.355 161.105 111.610 161.305 ;
        RECT 110.890 160.595 111.175 161.055 ;
        RECT 111.355 160.935 111.695 161.105 ;
        RECT 111.355 160.775 111.610 160.935 ;
        RECT 112.155 160.595 113.365 161.345 ;
        RECT 22.830 160.425 113.450 160.595 ;
        RECT 22.915 159.675 24.125 160.425 ;
        RECT 22.915 159.135 23.435 159.675 ;
        RECT 25.490 159.615 25.735 160.220 ;
        RECT 25.955 159.890 26.465 160.425 ;
        RECT 23.605 158.965 24.125 159.505 ;
        RECT 22.915 157.875 24.125 158.965 ;
        RECT 25.215 159.445 26.445 159.615 ;
        RECT 25.215 158.635 25.555 159.445 ;
        RECT 25.725 158.880 26.475 159.070 ;
        RECT 25.215 158.225 25.730 158.635 ;
        RECT 25.965 157.875 26.135 158.635 ;
        RECT 26.305 158.215 26.475 158.880 ;
        RECT 26.645 158.895 26.835 160.255 ;
        RECT 27.005 159.405 27.280 160.255 ;
        RECT 27.470 159.890 28.000 160.255 ;
        RECT 28.425 160.025 28.755 160.425 ;
        RECT 27.825 159.855 28.000 159.890 ;
        RECT 27.005 159.235 27.285 159.405 ;
        RECT 27.005 159.095 27.280 159.235 ;
        RECT 27.485 158.895 27.655 159.695 ;
        RECT 26.645 158.725 27.655 158.895 ;
        RECT 27.825 159.685 28.755 159.855 ;
        RECT 28.925 159.685 29.180 160.255 ;
        RECT 27.825 158.555 27.995 159.685 ;
        RECT 28.585 159.515 28.755 159.685 ;
        RECT 26.870 158.385 27.995 158.555 ;
        RECT 28.165 159.185 28.360 159.515 ;
        RECT 28.585 159.185 28.840 159.515 ;
        RECT 28.165 158.215 28.335 159.185 ;
        RECT 29.010 159.015 29.180 159.685 ;
        RECT 29.730 159.715 29.985 160.245 ;
        RECT 30.165 159.965 30.450 160.425 ;
        RECT 29.730 159.065 29.910 159.715 ;
        RECT 30.630 159.515 30.880 160.165 ;
        RECT 30.080 159.185 30.880 159.515 ;
        RECT 26.305 158.045 28.335 158.215 ;
        RECT 28.505 157.875 28.675 159.015 ;
        RECT 28.845 158.045 29.180 159.015 ;
        RECT 29.645 158.895 29.910 159.065 ;
        RECT 29.730 158.855 29.910 158.895 ;
        RECT 29.730 158.185 29.985 158.855 ;
        RECT 30.165 157.875 30.450 158.675 ;
        RECT 30.630 158.595 30.880 159.185 ;
        RECT 31.080 159.830 31.400 160.160 ;
        RECT 31.580 159.945 32.240 160.425 ;
        RECT 32.440 160.035 33.290 160.205 ;
        RECT 31.080 158.935 31.270 159.830 ;
        RECT 31.590 159.505 32.250 159.775 ;
        RECT 31.920 159.445 32.250 159.505 ;
        RECT 31.440 159.275 31.770 159.335 ;
        RECT 32.440 159.275 32.610 160.035 ;
        RECT 33.850 159.965 34.170 160.425 ;
        RECT 34.370 159.785 34.620 160.215 ;
        RECT 34.910 159.985 35.320 160.425 ;
        RECT 35.490 160.045 36.505 160.245 ;
        RECT 32.780 159.615 34.030 159.785 ;
        RECT 32.780 159.495 33.110 159.615 ;
        RECT 31.440 159.105 33.340 159.275 ;
        RECT 31.080 158.765 33.000 158.935 ;
        RECT 31.080 158.745 31.400 158.765 ;
        RECT 30.630 158.085 30.960 158.595 ;
        RECT 31.230 158.135 31.400 158.745 ;
        RECT 33.170 158.595 33.340 159.105 ;
        RECT 33.510 159.035 33.690 159.445 ;
        RECT 33.860 158.855 34.030 159.615 ;
        RECT 31.570 157.875 31.900 158.565 ;
        RECT 32.130 158.425 33.340 158.595 ;
        RECT 33.510 158.545 34.030 158.855 ;
        RECT 34.200 159.445 34.620 159.785 ;
        RECT 34.910 159.445 35.320 159.775 ;
        RECT 34.200 158.675 34.390 159.445 ;
        RECT 35.490 159.315 35.660 160.045 ;
        RECT 36.805 159.875 36.975 160.205 ;
        RECT 37.145 160.045 37.475 160.425 ;
        RECT 35.830 159.495 36.180 159.865 ;
        RECT 35.490 159.275 35.910 159.315 ;
        RECT 34.560 159.105 35.910 159.275 ;
        RECT 34.560 158.945 34.810 159.105 ;
        RECT 35.320 158.675 35.570 158.935 ;
        RECT 34.200 158.425 35.570 158.675 ;
        RECT 32.130 158.135 32.370 158.425 ;
        RECT 33.170 158.345 33.340 158.425 ;
        RECT 32.570 157.875 32.990 158.255 ;
        RECT 33.170 158.095 33.800 158.345 ;
        RECT 34.270 157.875 34.600 158.255 ;
        RECT 34.770 158.135 34.940 158.425 ;
        RECT 35.740 158.260 35.910 159.105 ;
        RECT 36.360 158.935 36.580 159.805 ;
        RECT 36.805 159.685 37.500 159.875 ;
        RECT 36.080 158.555 36.580 158.935 ;
        RECT 36.750 158.885 37.160 159.505 ;
        RECT 37.330 158.715 37.500 159.685 ;
        RECT 36.805 158.545 37.500 158.715 ;
        RECT 35.120 157.875 35.500 158.255 ;
        RECT 35.740 158.090 36.570 158.260 ;
        RECT 36.805 158.045 36.975 158.545 ;
        RECT 37.145 157.875 37.475 158.375 ;
        RECT 37.690 158.045 37.915 160.165 ;
        RECT 38.085 160.045 38.415 160.425 ;
        RECT 38.585 159.875 38.755 160.165 ;
        RECT 38.090 159.705 38.755 159.875 ;
        RECT 38.090 158.715 38.320 159.705 ;
        RECT 39.020 159.685 39.275 160.255 ;
        RECT 39.445 160.025 39.775 160.425 ;
        RECT 40.200 159.890 40.730 160.255 ;
        RECT 40.920 160.085 41.195 160.255 ;
        RECT 40.915 159.915 41.195 160.085 ;
        RECT 40.200 159.855 40.375 159.890 ;
        RECT 39.445 159.685 40.375 159.855 ;
        RECT 38.490 158.885 38.840 159.535 ;
        RECT 39.020 159.015 39.190 159.685 ;
        RECT 39.445 159.515 39.615 159.685 ;
        RECT 39.360 159.185 39.615 159.515 ;
        RECT 39.840 159.185 40.035 159.515 ;
        RECT 38.090 158.545 38.755 158.715 ;
        RECT 38.085 157.875 38.415 158.375 ;
        RECT 38.585 158.045 38.755 158.545 ;
        RECT 39.020 158.045 39.355 159.015 ;
        RECT 39.525 157.875 39.695 159.015 ;
        RECT 39.865 158.215 40.035 159.185 ;
        RECT 40.205 158.555 40.375 159.685 ;
        RECT 40.545 158.895 40.715 159.695 ;
        RECT 40.920 159.095 41.195 159.915 ;
        RECT 41.365 158.895 41.555 160.255 ;
        RECT 41.735 159.890 42.245 160.425 ;
        RECT 42.465 159.615 42.710 160.220 ;
        RECT 43.705 159.875 43.875 160.255 ;
        RECT 44.055 160.045 44.385 160.425 ;
        RECT 43.705 159.705 44.370 159.875 ;
        RECT 44.565 159.750 44.825 160.255 ;
        RECT 41.755 159.445 42.985 159.615 ;
        RECT 40.545 158.725 41.555 158.895 ;
        RECT 41.725 158.880 42.475 159.070 ;
        RECT 40.205 158.385 41.330 158.555 ;
        RECT 41.725 158.215 41.895 158.880 ;
        RECT 42.645 158.635 42.985 159.445 ;
        RECT 43.635 159.155 43.965 159.525 ;
        RECT 44.200 159.450 44.370 159.705 ;
        RECT 44.200 159.120 44.485 159.450 ;
        RECT 44.200 158.975 44.370 159.120 ;
        RECT 39.865 158.045 41.895 158.215 ;
        RECT 42.065 157.875 42.235 158.635 ;
        RECT 42.470 158.225 42.985 158.635 ;
        RECT 43.705 158.805 44.370 158.975 ;
        RECT 44.655 158.950 44.825 159.750 ;
        RECT 45.200 159.645 45.700 160.255 ;
        RECT 44.995 159.185 45.345 159.435 ;
        RECT 45.530 159.015 45.700 159.645 ;
        RECT 46.330 159.775 46.660 160.255 ;
        RECT 46.830 159.965 47.055 160.425 ;
        RECT 47.225 159.775 47.555 160.255 ;
        RECT 46.330 159.605 47.555 159.775 ;
        RECT 47.745 159.625 47.995 160.425 ;
        RECT 48.165 159.625 48.505 160.255 ;
        RECT 48.675 159.700 48.965 160.425 ;
        RECT 49.135 159.675 50.345 160.425 ;
        RECT 50.605 159.875 50.775 160.255 ;
        RECT 50.955 160.045 51.285 160.425 ;
        RECT 50.605 159.705 51.270 159.875 ;
        RECT 51.465 159.750 51.725 160.255 ;
        RECT 45.870 159.235 46.200 159.435 ;
        RECT 46.370 159.235 46.700 159.435 ;
        RECT 46.870 159.235 47.290 159.435 ;
        RECT 47.465 159.265 48.160 159.435 ;
        RECT 47.465 159.015 47.635 159.265 ;
        RECT 48.330 159.015 48.505 159.625 ;
        RECT 43.705 158.045 43.875 158.805 ;
        RECT 44.055 157.875 44.385 158.635 ;
        RECT 44.555 158.045 44.825 158.950 ;
        RECT 45.200 158.845 47.635 159.015 ;
        RECT 45.200 158.045 45.530 158.845 ;
        RECT 45.700 157.875 46.030 158.675 ;
        RECT 46.330 158.045 46.660 158.845 ;
        RECT 47.305 157.875 47.555 158.675 ;
        RECT 47.825 157.875 47.995 159.015 ;
        RECT 48.165 158.045 48.505 159.015 ;
        RECT 48.675 157.875 48.965 159.040 ;
        RECT 49.135 158.965 49.655 159.505 ;
        RECT 49.825 159.135 50.345 159.675 ;
        RECT 50.535 159.155 50.865 159.525 ;
        RECT 51.100 159.450 51.270 159.705 ;
        RECT 51.100 159.120 51.385 159.450 ;
        RECT 51.100 158.975 51.270 159.120 ;
        RECT 49.135 157.875 50.345 158.965 ;
        RECT 50.605 158.805 51.270 158.975 ;
        RECT 51.555 158.950 51.725 159.750 ;
        RECT 50.605 158.045 50.775 158.805 ;
        RECT 50.955 157.875 51.285 158.635 ;
        RECT 51.455 158.045 51.725 158.950 ;
        RECT 51.895 159.625 52.235 160.255 ;
        RECT 52.405 159.625 52.655 160.425 ;
        RECT 52.845 159.775 53.175 160.255 ;
        RECT 53.345 159.965 53.570 160.425 ;
        RECT 53.740 159.775 54.070 160.255 ;
        RECT 51.895 159.015 52.070 159.625 ;
        RECT 52.845 159.605 54.070 159.775 ;
        RECT 54.700 159.645 55.200 160.255 ;
        RECT 55.780 159.645 56.280 160.255 ;
        RECT 52.240 159.265 52.935 159.435 ;
        RECT 52.765 159.015 52.935 159.265 ;
        RECT 53.110 159.235 53.530 159.435 ;
        RECT 53.700 159.235 54.030 159.435 ;
        RECT 54.200 159.235 54.530 159.435 ;
        RECT 54.700 159.015 54.870 159.645 ;
        RECT 55.055 159.185 55.405 159.435 ;
        RECT 55.575 159.185 55.925 159.435 ;
        RECT 56.110 159.015 56.280 159.645 ;
        RECT 56.910 159.775 57.240 160.255 ;
        RECT 57.410 159.965 57.635 160.425 ;
        RECT 57.805 159.775 58.135 160.255 ;
        RECT 56.910 159.605 58.135 159.775 ;
        RECT 58.325 159.625 58.575 160.425 ;
        RECT 58.745 159.625 59.085 160.255 ;
        RECT 59.345 159.945 59.645 160.425 ;
        RECT 59.815 159.775 60.075 160.230 ;
        RECT 60.245 159.945 60.505 160.425 ;
        RECT 60.685 159.775 60.945 160.230 ;
        RECT 61.115 159.945 61.365 160.425 ;
        RECT 61.545 159.775 61.805 160.230 ;
        RECT 61.975 159.945 62.225 160.425 ;
        RECT 62.405 159.775 62.665 160.230 ;
        RECT 62.835 159.945 63.080 160.425 ;
        RECT 63.250 159.775 63.525 160.230 ;
        RECT 63.695 159.945 63.940 160.425 ;
        RECT 64.110 159.775 64.370 160.230 ;
        RECT 64.540 159.945 64.800 160.425 ;
        RECT 64.970 159.775 65.230 160.230 ;
        RECT 65.400 159.945 65.660 160.425 ;
        RECT 65.830 159.775 66.090 160.230 ;
        RECT 66.260 159.865 66.520 160.425 ;
        RECT 56.450 159.235 56.780 159.435 ;
        RECT 56.950 159.235 57.280 159.435 ;
        RECT 57.450 159.235 57.870 159.435 ;
        RECT 58.045 159.265 58.740 159.435 ;
        RECT 58.045 159.015 58.215 159.265 ;
        RECT 58.910 159.015 59.085 159.625 ;
        RECT 51.895 158.045 52.235 159.015 ;
        RECT 52.405 157.875 52.575 159.015 ;
        RECT 52.765 158.845 55.200 159.015 ;
        RECT 52.845 157.875 53.095 158.675 ;
        RECT 53.740 158.045 54.070 158.845 ;
        RECT 54.370 157.875 54.700 158.675 ;
        RECT 54.870 158.045 55.200 158.845 ;
        RECT 55.780 158.845 58.215 159.015 ;
        RECT 55.780 158.045 56.110 158.845 ;
        RECT 56.280 157.875 56.610 158.675 ;
        RECT 56.910 158.045 57.240 158.845 ;
        RECT 57.885 157.875 58.135 158.675 ;
        RECT 58.405 157.875 58.575 159.015 ;
        RECT 58.745 158.045 59.085 159.015 ;
        RECT 59.345 159.605 66.090 159.775 ;
        RECT 59.345 159.015 60.510 159.605 ;
        RECT 66.690 159.435 66.940 160.245 ;
        RECT 67.120 159.900 67.380 160.425 ;
        RECT 67.550 159.435 67.800 160.245 ;
        RECT 67.980 159.915 68.285 160.425 ;
        RECT 68.545 159.875 68.715 160.255 ;
        RECT 68.930 160.045 69.260 160.425 ;
        RECT 60.680 159.185 67.800 159.435 ;
        RECT 67.970 159.185 68.285 159.745 ;
        RECT 68.545 159.705 69.260 159.875 ;
        RECT 59.345 158.790 66.090 159.015 ;
        RECT 59.345 157.875 59.615 158.620 ;
        RECT 59.785 158.050 60.075 158.790 ;
        RECT 60.685 158.775 66.090 158.790 ;
        RECT 60.245 157.880 60.500 158.605 ;
        RECT 60.685 158.050 60.945 158.775 ;
        RECT 61.115 157.880 61.360 158.605 ;
        RECT 61.545 158.050 61.805 158.775 ;
        RECT 61.975 157.880 62.220 158.605 ;
        RECT 62.405 158.050 62.665 158.775 ;
        RECT 62.835 157.880 63.080 158.605 ;
        RECT 63.250 158.050 63.510 158.775 ;
        RECT 63.680 157.880 63.940 158.605 ;
        RECT 64.110 158.050 64.370 158.775 ;
        RECT 64.540 157.880 64.800 158.605 ;
        RECT 64.970 158.050 65.230 158.775 ;
        RECT 65.400 157.880 65.660 158.605 ;
        RECT 65.830 158.050 66.090 158.775 ;
        RECT 66.260 157.880 66.520 158.675 ;
        RECT 66.690 158.050 66.940 159.185 ;
        RECT 60.245 157.875 66.520 157.880 ;
        RECT 67.120 157.875 67.380 158.685 ;
        RECT 67.555 158.045 67.800 159.185 ;
        RECT 68.455 159.155 68.810 159.525 ;
        RECT 69.090 159.515 69.260 159.705 ;
        RECT 69.430 159.680 69.685 160.255 ;
        RECT 69.090 159.185 69.345 159.515 ;
        RECT 69.090 158.975 69.260 159.185 ;
        RECT 68.545 158.805 69.260 158.975 ;
        RECT 69.515 158.950 69.685 159.680 ;
        RECT 69.860 159.585 70.120 160.425 ;
        RECT 70.755 159.625 71.095 160.255 ;
        RECT 71.265 159.625 71.515 160.425 ;
        RECT 71.705 159.775 72.035 160.255 ;
        RECT 72.205 159.965 72.430 160.425 ;
        RECT 72.600 159.775 72.930 160.255 ;
        RECT 67.980 157.875 68.275 158.685 ;
        RECT 68.545 158.045 68.715 158.805 ;
        RECT 68.930 157.875 69.260 158.635 ;
        RECT 69.430 158.045 69.685 158.950 ;
        RECT 69.860 157.875 70.120 159.025 ;
        RECT 70.755 159.015 70.930 159.625 ;
        RECT 71.705 159.605 72.930 159.775 ;
        RECT 73.560 159.645 74.060 160.255 ;
        RECT 74.435 159.700 74.725 160.425 ;
        RECT 74.985 159.875 75.155 160.255 ;
        RECT 75.370 160.045 75.700 160.425 ;
        RECT 74.985 159.705 75.700 159.875 ;
        RECT 71.100 159.265 71.795 159.435 ;
        RECT 71.625 159.015 71.795 159.265 ;
        RECT 71.970 159.235 72.390 159.435 ;
        RECT 72.560 159.235 72.890 159.435 ;
        RECT 73.060 159.235 73.390 159.435 ;
        RECT 73.560 159.015 73.730 159.645 ;
        RECT 73.915 159.185 74.265 159.435 ;
        RECT 74.895 159.155 75.250 159.525 ;
        RECT 75.530 159.515 75.700 159.705 ;
        RECT 75.870 159.680 76.125 160.255 ;
        RECT 75.530 159.185 75.785 159.515 ;
        RECT 70.755 158.045 71.095 159.015 ;
        RECT 71.265 157.875 71.435 159.015 ;
        RECT 71.625 158.845 74.060 159.015 ;
        RECT 71.705 157.875 71.955 158.675 ;
        RECT 72.600 158.045 72.930 158.845 ;
        RECT 73.230 157.875 73.560 158.675 ;
        RECT 73.730 158.045 74.060 158.845 ;
        RECT 74.435 157.875 74.725 159.040 ;
        RECT 75.530 158.975 75.700 159.185 ;
        RECT 74.985 158.805 75.700 158.975 ;
        RECT 75.955 158.950 76.125 159.680 ;
        RECT 76.300 159.585 76.560 160.425 ;
        RECT 77.255 159.605 77.465 160.425 ;
        RECT 77.635 159.625 77.965 160.255 ;
        RECT 77.635 159.025 77.885 159.625 ;
        RECT 78.135 159.605 78.365 160.425 ;
        RECT 78.635 159.605 78.845 160.425 ;
        RECT 79.015 159.625 79.345 160.255 ;
        RECT 78.055 159.185 78.385 159.435 ;
        RECT 79.015 159.025 79.265 159.625 ;
        RECT 79.515 159.605 79.745 160.425 ;
        RECT 80.045 159.875 80.215 160.255 ;
        RECT 80.395 160.045 80.725 160.425 ;
        RECT 80.045 159.705 80.710 159.875 ;
        RECT 80.905 159.750 81.165 160.255 ;
        RECT 79.435 159.185 79.765 159.435 ;
        RECT 79.975 159.155 80.305 159.525 ;
        RECT 80.540 159.450 80.710 159.705 ;
        RECT 80.540 159.120 80.825 159.450 ;
        RECT 74.985 158.045 75.155 158.805 ;
        RECT 75.370 157.875 75.700 158.635 ;
        RECT 75.870 158.045 76.125 158.950 ;
        RECT 76.300 157.875 76.560 159.025 ;
        RECT 77.255 157.875 77.465 159.015 ;
        RECT 77.635 158.045 77.965 159.025 ;
        RECT 78.135 157.875 78.365 159.015 ;
        RECT 78.635 157.875 78.845 159.015 ;
        RECT 79.015 158.045 79.345 159.025 ;
        RECT 79.515 157.875 79.745 159.015 ;
        RECT 80.540 158.975 80.710 159.120 ;
        RECT 80.045 158.805 80.710 158.975 ;
        RECT 80.995 158.950 81.165 159.750 ;
        RECT 81.425 159.875 81.595 160.255 ;
        RECT 81.775 160.045 82.105 160.425 ;
        RECT 81.425 159.705 82.090 159.875 ;
        RECT 82.285 159.750 82.545 160.255 ;
        RECT 81.355 159.155 81.685 159.525 ;
        RECT 81.920 159.450 82.090 159.705 ;
        RECT 81.920 159.120 82.205 159.450 ;
        RECT 81.920 158.975 82.090 159.120 ;
        RECT 80.045 158.045 80.215 158.805 ;
        RECT 80.395 157.875 80.725 158.635 ;
        RECT 80.895 158.045 81.165 158.950 ;
        RECT 81.425 158.805 82.090 158.975 ;
        RECT 82.375 158.950 82.545 159.750 ;
        RECT 81.425 158.045 81.595 158.805 ;
        RECT 81.775 157.875 82.105 158.635 ;
        RECT 82.275 158.045 82.545 158.950 ;
        RECT 82.720 159.715 82.975 160.245 ;
        RECT 83.145 159.965 83.450 160.425 ;
        RECT 83.695 160.045 84.765 160.215 ;
        RECT 82.720 159.065 82.930 159.715 ;
        RECT 83.695 159.690 84.015 160.045 ;
        RECT 83.690 159.515 84.015 159.690 ;
        RECT 83.100 159.215 84.015 159.515 ;
        RECT 84.185 159.475 84.425 159.875 ;
        RECT 84.595 159.815 84.765 160.045 ;
        RECT 84.935 159.985 85.125 160.425 ;
        RECT 85.295 159.975 86.245 160.255 ;
        RECT 86.465 160.065 86.815 160.235 ;
        RECT 84.595 159.645 85.125 159.815 ;
        RECT 83.100 159.185 83.840 159.215 ;
        RECT 82.720 158.185 82.975 159.065 ;
        RECT 83.145 157.875 83.450 159.015 ;
        RECT 83.670 158.595 83.840 159.185 ;
        RECT 84.185 159.105 84.725 159.475 ;
        RECT 84.905 159.365 85.125 159.645 ;
        RECT 85.295 159.195 85.465 159.975 ;
        RECT 85.060 159.025 85.465 159.195 ;
        RECT 85.635 159.185 85.985 159.805 ;
        RECT 85.060 158.935 85.230 159.025 ;
        RECT 86.155 159.015 86.365 159.805 ;
        RECT 84.010 158.765 85.230 158.935 ;
        RECT 85.690 158.855 86.365 159.015 ;
        RECT 83.670 158.425 84.470 158.595 ;
        RECT 83.790 157.875 84.120 158.255 ;
        RECT 84.300 158.135 84.470 158.425 ;
        RECT 85.060 158.385 85.230 158.765 ;
        RECT 85.400 158.845 86.365 158.855 ;
        RECT 86.555 159.675 86.815 160.065 ;
        RECT 87.025 159.965 87.355 160.425 ;
        RECT 88.230 160.035 89.085 160.205 ;
        RECT 89.290 160.035 89.785 160.205 ;
        RECT 89.955 160.065 90.285 160.425 ;
        RECT 86.555 158.985 86.725 159.675 ;
        RECT 86.895 159.325 87.065 159.505 ;
        RECT 87.235 159.495 88.025 159.745 ;
        RECT 88.230 159.325 88.400 160.035 ;
        RECT 88.570 159.525 88.925 159.745 ;
        RECT 86.895 159.155 88.585 159.325 ;
        RECT 85.400 158.555 85.860 158.845 ;
        RECT 86.555 158.815 88.055 158.985 ;
        RECT 86.555 158.675 86.725 158.815 ;
        RECT 86.165 158.505 86.725 158.675 ;
        RECT 84.640 157.875 84.890 158.335 ;
        RECT 85.060 158.045 85.930 158.385 ;
        RECT 86.165 158.045 86.335 158.505 ;
        RECT 87.170 158.475 88.245 158.645 ;
        RECT 86.505 157.875 86.875 158.335 ;
        RECT 87.170 158.135 87.340 158.475 ;
        RECT 87.510 157.875 87.840 158.305 ;
        RECT 88.075 158.135 88.245 158.475 ;
        RECT 88.415 158.375 88.585 159.155 ;
        RECT 88.755 158.935 88.925 159.525 ;
        RECT 89.095 159.125 89.445 159.745 ;
        RECT 88.755 158.545 89.220 158.935 ;
        RECT 89.615 158.675 89.785 160.035 ;
        RECT 89.955 158.845 90.415 159.895 ;
        RECT 89.390 158.505 89.785 158.675 ;
        RECT 89.390 158.375 89.560 158.505 ;
        RECT 88.415 158.045 89.095 158.375 ;
        RECT 89.310 158.045 89.560 158.375 ;
        RECT 89.730 157.875 89.980 158.335 ;
        RECT 90.150 158.060 90.475 158.845 ;
        RECT 90.645 158.045 90.815 160.165 ;
        RECT 90.985 160.045 91.315 160.425 ;
        RECT 91.485 159.875 91.740 160.165 ;
        RECT 90.990 159.705 91.740 159.875 ;
        RECT 90.990 158.715 91.220 159.705 ;
        RECT 92.835 159.625 93.175 160.255 ;
        RECT 93.345 159.625 93.595 160.425 ;
        RECT 93.785 159.775 94.115 160.255 ;
        RECT 94.285 159.965 94.510 160.425 ;
        RECT 94.680 159.775 95.010 160.255 ;
        RECT 91.390 158.885 91.740 159.535 ;
        RECT 92.835 159.015 93.010 159.625 ;
        RECT 93.785 159.605 95.010 159.775 ;
        RECT 95.640 159.645 96.140 160.255 ;
        RECT 93.180 159.265 93.875 159.435 ;
        RECT 93.705 159.015 93.875 159.265 ;
        RECT 94.050 159.235 94.470 159.435 ;
        RECT 94.640 159.235 94.970 159.435 ;
        RECT 95.140 159.235 95.470 159.435 ;
        RECT 95.640 159.015 95.810 159.645 ;
        RECT 96.515 159.625 96.855 160.255 ;
        RECT 97.025 159.625 97.275 160.425 ;
        RECT 97.465 159.775 97.795 160.255 ;
        RECT 97.965 159.965 98.190 160.425 ;
        RECT 98.360 159.775 98.690 160.255 ;
        RECT 95.995 159.185 96.345 159.435 ;
        RECT 96.515 159.015 96.690 159.625 ;
        RECT 97.465 159.605 98.690 159.775 ;
        RECT 99.320 159.645 99.820 160.255 ;
        RECT 100.195 159.700 100.485 160.425 ;
        RECT 96.860 159.265 97.555 159.435 ;
        RECT 97.385 159.015 97.555 159.265 ;
        RECT 97.730 159.235 98.150 159.435 ;
        RECT 98.320 159.235 98.650 159.435 ;
        RECT 98.820 159.235 99.150 159.435 ;
        RECT 99.320 159.015 99.490 159.645 ;
        RECT 101.850 159.615 102.095 160.220 ;
        RECT 102.315 159.890 102.825 160.425 ;
        RECT 101.575 159.445 102.805 159.615 ;
        RECT 99.675 159.185 100.025 159.435 ;
        RECT 90.990 158.545 91.740 158.715 ;
        RECT 90.985 157.875 91.315 158.375 ;
        RECT 91.485 158.045 91.740 158.545 ;
        RECT 92.835 158.045 93.175 159.015 ;
        RECT 93.345 157.875 93.515 159.015 ;
        RECT 93.705 158.845 96.140 159.015 ;
        RECT 93.785 157.875 94.035 158.675 ;
        RECT 94.680 158.045 95.010 158.845 ;
        RECT 95.310 157.875 95.640 158.675 ;
        RECT 95.810 158.045 96.140 158.845 ;
        RECT 96.515 158.045 96.855 159.015 ;
        RECT 97.025 157.875 97.195 159.015 ;
        RECT 97.385 158.845 99.820 159.015 ;
        RECT 97.465 157.875 97.715 158.675 ;
        RECT 98.360 158.045 98.690 158.845 ;
        RECT 98.990 157.875 99.320 158.675 ;
        RECT 99.490 158.045 99.820 158.845 ;
        RECT 100.195 157.875 100.485 159.040 ;
        RECT 101.575 158.635 101.915 159.445 ;
        RECT 102.085 158.880 102.835 159.070 ;
        RECT 101.575 158.225 102.090 158.635 ;
        RECT 102.325 157.875 102.495 158.635 ;
        RECT 102.665 158.215 102.835 158.880 ;
        RECT 103.005 158.895 103.195 160.255 ;
        RECT 103.365 160.085 103.640 160.255 ;
        RECT 103.365 159.915 103.645 160.085 ;
        RECT 103.365 159.095 103.640 159.915 ;
        RECT 103.830 159.890 104.360 160.255 ;
        RECT 104.785 160.025 105.115 160.425 ;
        RECT 104.185 159.855 104.360 159.890 ;
        RECT 103.845 158.895 104.015 159.695 ;
        RECT 103.005 158.725 104.015 158.895 ;
        RECT 104.185 159.685 105.115 159.855 ;
        RECT 105.285 159.685 105.540 160.255 ;
        RECT 104.185 158.555 104.355 159.685 ;
        RECT 104.945 159.515 105.115 159.685 ;
        RECT 103.230 158.385 104.355 158.555 ;
        RECT 104.525 159.185 104.720 159.515 ;
        RECT 104.945 159.185 105.200 159.515 ;
        RECT 104.525 158.215 104.695 159.185 ;
        RECT 105.370 159.015 105.540 159.685 ;
        RECT 102.665 158.045 104.695 158.215 ;
        RECT 104.865 157.875 105.035 159.015 ;
        RECT 105.205 158.045 105.540 159.015 ;
        RECT 105.720 159.685 105.975 160.255 ;
        RECT 106.145 160.025 106.475 160.425 ;
        RECT 106.900 159.890 107.430 160.255 ;
        RECT 106.900 159.855 107.075 159.890 ;
        RECT 106.145 159.685 107.075 159.855 ;
        RECT 107.620 159.745 107.895 160.255 ;
        RECT 105.720 159.015 105.890 159.685 ;
        RECT 106.145 159.515 106.315 159.685 ;
        RECT 106.060 159.185 106.315 159.515 ;
        RECT 106.540 159.185 106.735 159.515 ;
        RECT 105.720 158.045 106.055 159.015 ;
        RECT 106.225 157.875 106.395 159.015 ;
        RECT 106.565 158.215 106.735 159.185 ;
        RECT 106.905 158.555 107.075 159.685 ;
        RECT 107.245 158.895 107.415 159.695 ;
        RECT 107.615 159.575 107.895 159.745 ;
        RECT 107.620 159.095 107.895 159.575 ;
        RECT 108.065 158.895 108.255 160.255 ;
        RECT 108.435 159.890 108.945 160.425 ;
        RECT 109.165 159.615 109.410 160.220 ;
        RECT 109.855 159.750 110.115 160.255 ;
        RECT 110.295 160.045 110.625 160.425 ;
        RECT 110.805 159.875 110.975 160.255 ;
        RECT 108.455 159.445 109.685 159.615 ;
        RECT 107.245 158.725 108.255 158.895 ;
        RECT 108.425 158.880 109.175 159.070 ;
        RECT 106.905 158.385 108.030 158.555 ;
        RECT 108.425 158.215 108.595 158.880 ;
        RECT 109.345 158.635 109.685 159.445 ;
        RECT 106.565 158.045 108.595 158.215 ;
        RECT 108.765 157.875 108.935 158.635 ;
        RECT 109.170 158.225 109.685 158.635 ;
        RECT 109.855 158.950 110.025 159.750 ;
        RECT 110.310 159.705 110.975 159.875 ;
        RECT 110.310 159.450 110.480 159.705 ;
        RECT 112.155 159.675 113.365 160.425 ;
        RECT 110.195 159.120 110.480 159.450 ;
        RECT 110.715 159.155 111.045 159.525 ;
        RECT 110.310 158.975 110.480 159.120 ;
        RECT 109.855 158.045 110.125 158.950 ;
        RECT 110.310 158.805 110.975 158.975 ;
        RECT 110.295 157.875 110.625 158.635 ;
        RECT 110.805 158.045 110.975 158.805 ;
        RECT 112.155 158.965 112.675 159.505 ;
        RECT 112.845 159.135 113.365 159.675 ;
        RECT 112.155 157.875 113.365 158.965 ;
        RECT 22.830 157.705 113.450 157.875 ;
        RECT 22.915 156.615 24.125 157.705 ;
        RECT 22.915 155.905 23.435 156.445 ;
        RECT 23.605 156.075 24.125 156.615 ;
        RECT 24.295 156.615 27.805 157.705 ;
        RECT 24.295 156.095 25.985 156.615 ;
        RECT 28.035 156.565 28.245 157.705 ;
        RECT 28.415 156.555 28.745 157.535 ;
        RECT 28.915 156.565 29.145 157.705 ;
        RECT 29.445 156.775 29.615 157.535 ;
        RECT 29.795 156.945 30.125 157.705 ;
        RECT 29.445 156.605 30.110 156.775 ;
        RECT 30.295 156.630 30.565 157.535 ;
        RECT 26.155 155.925 27.805 156.445 ;
        RECT 22.915 155.155 24.125 155.905 ;
        RECT 24.295 155.155 27.805 155.925 ;
        RECT 28.035 155.155 28.245 155.975 ;
        RECT 28.415 155.955 28.665 156.555 ;
        RECT 29.940 156.460 30.110 156.605 ;
        RECT 28.835 156.145 29.165 156.395 ;
        RECT 29.375 156.055 29.705 156.425 ;
        RECT 29.940 156.130 30.225 156.460 ;
        RECT 28.415 155.325 28.745 155.955 ;
        RECT 28.915 155.155 29.145 155.975 ;
        RECT 29.940 155.875 30.110 156.130 ;
        RECT 29.445 155.705 30.110 155.875 ;
        RECT 30.395 155.830 30.565 156.630 ;
        RECT 30.775 156.565 31.005 157.705 ;
        RECT 31.175 156.555 31.505 157.535 ;
        RECT 31.675 156.565 31.885 157.705 ;
        RECT 32.320 156.735 32.650 157.535 ;
        RECT 32.820 156.905 33.150 157.705 ;
        RECT 33.450 156.735 33.780 157.535 ;
        RECT 34.425 156.905 34.675 157.705 ;
        RECT 32.320 156.565 34.755 156.735 ;
        RECT 34.945 156.565 35.115 157.705 ;
        RECT 35.285 156.565 35.625 157.535 ;
        RECT 30.755 156.145 31.085 156.395 ;
        RECT 29.445 155.325 29.615 155.705 ;
        RECT 29.795 155.155 30.125 155.535 ;
        RECT 30.305 155.325 30.565 155.830 ;
        RECT 30.775 155.155 31.005 155.975 ;
        RECT 31.255 155.955 31.505 156.555 ;
        RECT 32.115 156.145 32.465 156.395 ;
        RECT 31.175 155.325 31.505 155.955 ;
        RECT 31.675 155.155 31.885 155.975 ;
        RECT 32.650 155.935 32.820 156.565 ;
        RECT 32.990 156.145 33.320 156.345 ;
        RECT 33.490 156.145 33.820 156.345 ;
        RECT 33.990 156.145 34.410 156.345 ;
        RECT 34.585 156.315 34.755 156.565 ;
        RECT 34.585 156.145 35.280 156.315 ;
        RECT 32.320 155.325 32.820 155.935 ;
        RECT 33.450 155.805 34.675 155.975 ;
        RECT 35.450 155.955 35.625 156.565 ;
        RECT 35.795 156.540 36.085 157.705 ;
        RECT 36.715 156.615 38.385 157.705 ;
        RECT 36.715 156.095 37.465 156.615 ;
        RECT 38.555 156.565 38.895 157.535 ;
        RECT 39.065 156.565 39.235 157.705 ;
        RECT 39.505 156.905 39.755 157.705 ;
        RECT 40.400 156.735 40.730 157.535 ;
        RECT 41.030 156.905 41.360 157.705 ;
        RECT 41.530 156.735 41.860 157.535 ;
        RECT 39.425 156.565 41.860 156.735 ;
        RECT 42.695 156.565 43.035 157.535 ;
        RECT 43.205 156.565 43.375 157.705 ;
        RECT 43.645 156.905 43.895 157.705 ;
        RECT 44.540 156.735 44.870 157.535 ;
        RECT 45.170 156.905 45.500 157.705 ;
        RECT 45.670 156.735 46.000 157.535 ;
        RECT 43.565 156.565 46.000 156.735 ;
        RECT 46.750 156.725 47.005 157.395 ;
        RECT 47.185 156.905 47.470 157.705 ;
        RECT 47.650 156.985 47.980 157.495 ;
        RECT 33.450 155.325 33.780 155.805 ;
        RECT 33.950 155.155 34.175 155.615 ;
        RECT 34.345 155.325 34.675 155.805 ;
        RECT 34.865 155.155 35.115 155.955 ;
        RECT 35.285 155.325 35.625 155.955 ;
        RECT 37.635 155.925 38.385 156.445 ;
        RECT 35.795 155.155 36.085 155.880 ;
        RECT 36.715 155.155 38.385 155.925 ;
        RECT 38.555 155.955 38.730 156.565 ;
        RECT 39.425 156.315 39.595 156.565 ;
        RECT 38.900 156.145 39.595 156.315 ;
        RECT 39.770 156.145 40.190 156.345 ;
        RECT 40.360 156.145 40.690 156.345 ;
        RECT 40.860 156.145 41.190 156.345 ;
        RECT 38.555 155.325 38.895 155.955 ;
        RECT 39.065 155.155 39.315 155.955 ;
        RECT 39.505 155.805 40.730 155.975 ;
        RECT 39.505 155.325 39.835 155.805 ;
        RECT 40.005 155.155 40.230 155.615 ;
        RECT 40.400 155.325 40.730 155.805 ;
        RECT 41.360 155.935 41.530 156.565 ;
        RECT 41.715 156.145 42.065 156.395 ;
        RECT 42.695 155.955 42.870 156.565 ;
        RECT 43.565 156.315 43.735 156.565 ;
        RECT 43.040 156.145 43.735 156.315 ;
        RECT 43.910 156.145 44.330 156.345 ;
        RECT 44.500 156.145 44.830 156.345 ;
        RECT 45.000 156.145 45.330 156.345 ;
        RECT 41.360 155.325 41.860 155.935 ;
        RECT 42.695 155.325 43.035 155.955 ;
        RECT 43.205 155.155 43.455 155.955 ;
        RECT 43.645 155.805 44.870 155.975 ;
        RECT 43.645 155.325 43.975 155.805 ;
        RECT 44.145 155.155 44.370 155.615 ;
        RECT 44.540 155.325 44.870 155.805 ;
        RECT 45.500 155.935 45.670 156.565 ;
        RECT 45.855 156.145 46.205 156.395 ;
        RECT 45.500 155.325 46.000 155.935 ;
        RECT 46.750 155.865 46.930 156.725 ;
        RECT 47.650 156.395 47.900 156.985 ;
        RECT 48.250 156.835 48.420 157.445 ;
        RECT 48.590 157.015 48.920 157.705 ;
        RECT 49.150 157.155 49.390 157.445 ;
        RECT 49.590 157.325 50.010 157.705 ;
        RECT 50.190 157.235 50.820 157.485 ;
        RECT 51.290 157.325 51.620 157.705 ;
        RECT 50.190 157.155 50.360 157.235 ;
        RECT 51.790 157.155 51.960 157.445 ;
        RECT 52.140 157.325 52.520 157.705 ;
        RECT 52.760 157.320 53.590 157.490 ;
        RECT 49.150 156.985 50.360 157.155 ;
        RECT 47.100 156.065 47.900 156.395 ;
        RECT 46.750 155.665 47.005 155.865 ;
        RECT 46.665 155.495 47.005 155.665 ;
        RECT 46.750 155.335 47.005 155.495 ;
        RECT 47.185 155.155 47.470 155.615 ;
        RECT 47.650 155.415 47.900 156.065 ;
        RECT 48.100 156.815 48.420 156.835 ;
        RECT 48.100 156.645 50.020 156.815 ;
        RECT 48.100 155.750 48.290 156.645 ;
        RECT 50.190 156.475 50.360 156.985 ;
        RECT 50.530 156.725 51.050 157.035 ;
        RECT 48.460 156.305 50.360 156.475 ;
        RECT 48.460 156.245 48.790 156.305 ;
        RECT 48.940 156.075 49.270 156.135 ;
        RECT 48.610 155.805 49.270 156.075 ;
        RECT 48.100 155.420 48.420 155.750 ;
        RECT 48.600 155.155 49.260 155.635 ;
        RECT 49.460 155.545 49.630 156.305 ;
        RECT 50.530 156.135 50.710 156.545 ;
        RECT 49.800 155.965 50.130 156.085 ;
        RECT 50.880 155.965 51.050 156.725 ;
        RECT 49.800 155.795 51.050 155.965 ;
        RECT 51.220 156.905 52.590 157.155 ;
        RECT 51.220 156.135 51.410 156.905 ;
        RECT 52.340 156.645 52.590 156.905 ;
        RECT 51.580 156.475 51.830 156.635 ;
        RECT 52.760 156.475 52.930 157.320 ;
        RECT 53.825 157.035 53.995 157.535 ;
        RECT 54.165 157.205 54.495 157.705 ;
        RECT 53.100 156.645 53.600 157.025 ;
        RECT 53.825 156.865 54.520 157.035 ;
        RECT 51.580 156.305 52.930 156.475 ;
        RECT 52.510 156.265 52.930 156.305 ;
        RECT 51.220 155.795 51.640 156.135 ;
        RECT 51.930 155.805 52.340 156.135 ;
        RECT 49.460 155.375 50.310 155.545 ;
        RECT 50.870 155.155 51.190 155.615 ;
        RECT 51.390 155.365 51.640 155.795 ;
        RECT 51.930 155.155 52.340 155.595 ;
        RECT 52.510 155.535 52.680 156.265 ;
        RECT 52.850 155.715 53.200 156.085 ;
        RECT 53.380 155.775 53.600 156.645 ;
        RECT 53.770 156.075 54.180 156.695 ;
        RECT 54.350 155.895 54.520 156.865 ;
        RECT 53.825 155.705 54.520 155.895 ;
        RECT 52.510 155.335 53.525 155.535 ;
        RECT 53.825 155.375 53.995 155.705 ;
        RECT 54.165 155.155 54.495 155.535 ;
        RECT 54.710 155.415 54.935 157.535 ;
        RECT 55.105 157.205 55.435 157.705 ;
        RECT 55.605 157.035 55.775 157.535 ;
        RECT 55.110 156.865 55.775 157.035 ;
        RECT 55.110 155.875 55.340 156.865 ;
        RECT 55.510 156.045 55.860 156.695 ;
        RECT 56.075 156.565 56.305 157.705 ;
        RECT 56.475 156.555 56.805 157.535 ;
        RECT 56.975 156.565 57.185 157.705 ;
        RECT 57.530 157.075 57.815 157.535 ;
        RECT 57.985 157.245 58.255 157.705 ;
        RECT 57.530 156.855 58.485 157.075 ;
        RECT 56.055 156.145 56.385 156.395 ;
        RECT 55.110 155.705 55.775 155.875 ;
        RECT 55.105 155.155 55.435 155.535 ;
        RECT 55.605 155.415 55.775 155.705 ;
        RECT 56.075 155.155 56.305 155.975 ;
        RECT 56.555 155.955 56.805 156.555 ;
        RECT 57.415 156.125 58.105 156.685 ;
        RECT 56.475 155.325 56.805 155.955 ;
        RECT 56.975 155.155 57.185 155.975 ;
        RECT 58.275 155.955 58.485 156.855 ;
        RECT 57.530 155.785 58.485 155.955 ;
        RECT 58.655 156.685 59.055 157.535 ;
        RECT 59.245 157.075 59.525 157.535 ;
        RECT 60.045 157.245 60.370 157.705 ;
        RECT 59.245 156.855 60.370 157.075 ;
        RECT 58.655 156.125 59.750 156.685 ;
        RECT 59.920 156.395 60.370 156.855 ;
        RECT 60.540 156.565 60.925 157.535 ;
        RECT 57.530 155.325 57.815 155.785 ;
        RECT 57.985 155.155 58.255 155.615 ;
        RECT 58.655 155.325 59.055 156.125 ;
        RECT 59.920 156.065 60.475 156.395 ;
        RECT 59.920 155.955 60.370 156.065 ;
        RECT 59.245 155.785 60.370 155.955 ;
        RECT 60.645 155.895 60.925 156.565 ;
        RECT 61.555 156.540 61.845 157.705 ;
        RECT 62.075 156.565 62.285 157.705 ;
        RECT 62.455 156.555 62.785 157.535 ;
        RECT 62.955 156.565 63.185 157.705 ;
        RECT 63.400 156.555 63.660 157.705 ;
        RECT 63.835 156.630 64.090 157.535 ;
        RECT 64.260 156.945 64.590 157.705 ;
        RECT 64.805 156.775 64.975 157.535 ;
        RECT 59.245 155.325 59.525 155.785 ;
        RECT 60.045 155.155 60.370 155.615 ;
        RECT 60.540 155.325 60.925 155.895 ;
        RECT 61.555 155.155 61.845 155.880 ;
        RECT 62.075 155.155 62.285 155.975 ;
        RECT 62.455 155.955 62.705 156.555 ;
        RECT 62.875 156.145 63.205 156.395 ;
        RECT 62.455 155.325 62.785 155.955 ;
        RECT 62.955 155.155 63.185 155.975 ;
        RECT 63.400 155.155 63.660 155.995 ;
        RECT 63.835 155.900 64.005 156.630 ;
        RECT 64.260 156.605 64.975 156.775 ;
        RECT 65.325 156.775 65.495 157.535 ;
        RECT 65.710 156.945 66.040 157.705 ;
        RECT 65.325 156.605 66.040 156.775 ;
        RECT 66.210 156.630 66.465 157.535 ;
        RECT 64.260 156.395 64.430 156.605 ;
        RECT 64.175 156.065 64.430 156.395 ;
        RECT 63.835 155.325 64.090 155.900 ;
        RECT 64.260 155.875 64.430 156.065 ;
        RECT 64.710 156.055 65.065 156.425 ;
        RECT 65.235 156.055 65.590 156.425 ;
        RECT 65.870 156.395 66.040 156.605 ;
        RECT 65.870 156.065 66.125 156.395 ;
        RECT 65.870 155.875 66.040 156.065 ;
        RECT 66.295 155.900 66.465 156.630 ;
        RECT 66.640 156.555 66.900 157.705 ;
        RECT 67.165 156.775 67.335 157.535 ;
        RECT 67.550 156.945 67.880 157.705 ;
        RECT 67.165 156.605 67.880 156.775 ;
        RECT 68.050 156.630 68.305 157.535 ;
        RECT 67.075 156.055 67.430 156.425 ;
        RECT 67.710 156.395 67.880 156.605 ;
        RECT 67.710 156.065 67.965 156.395 ;
        RECT 64.260 155.705 64.975 155.875 ;
        RECT 64.260 155.155 64.590 155.535 ;
        RECT 64.805 155.325 64.975 155.705 ;
        RECT 65.325 155.705 66.040 155.875 ;
        RECT 65.325 155.325 65.495 155.705 ;
        RECT 65.710 155.155 66.040 155.535 ;
        RECT 66.210 155.325 66.465 155.900 ;
        RECT 66.640 155.155 66.900 155.995 ;
        RECT 67.710 155.875 67.880 156.065 ;
        RECT 68.135 155.900 68.305 156.630 ;
        RECT 68.480 156.555 68.740 157.705 ;
        RECT 69.005 156.775 69.175 157.535 ;
        RECT 69.390 156.945 69.720 157.705 ;
        RECT 69.005 156.605 69.720 156.775 ;
        RECT 69.890 156.630 70.145 157.535 ;
        RECT 68.915 156.055 69.270 156.425 ;
        RECT 69.550 156.395 69.720 156.605 ;
        RECT 69.550 156.065 69.805 156.395 ;
        RECT 67.165 155.705 67.880 155.875 ;
        RECT 67.165 155.325 67.335 155.705 ;
        RECT 67.550 155.155 67.880 155.535 ;
        RECT 68.050 155.325 68.305 155.900 ;
        RECT 68.480 155.155 68.740 155.995 ;
        RECT 69.550 155.875 69.720 156.065 ;
        RECT 69.975 155.900 70.145 156.630 ;
        RECT 70.320 156.555 70.580 157.705 ;
        RECT 70.765 156.645 71.095 157.705 ;
        RECT 71.275 156.395 71.445 157.365 ;
        RECT 71.615 157.115 71.945 157.515 ;
        RECT 72.115 157.345 72.445 157.705 ;
        RECT 72.645 157.115 73.345 157.535 ;
        RECT 71.615 156.885 73.345 157.115 ;
        RECT 71.615 156.665 71.945 156.885 ;
        RECT 72.140 156.395 72.465 156.685 ;
        RECT 70.755 156.065 71.065 156.395 ;
        RECT 71.275 156.065 71.650 156.395 ;
        RECT 71.970 156.065 72.465 156.395 ;
        RECT 72.640 156.145 72.970 156.685 ;
        RECT 69.005 155.705 69.720 155.875 ;
        RECT 69.005 155.325 69.175 155.705 ;
        RECT 69.390 155.155 69.720 155.535 ;
        RECT 69.890 155.325 70.145 155.900 ;
        RECT 70.320 155.155 70.580 155.995 ;
        RECT 73.140 155.915 73.345 156.885 ;
        RECT 73.605 156.775 73.775 157.535 ;
        RECT 73.990 156.945 74.320 157.705 ;
        RECT 73.605 156.605 74.320 156.775 ;
        RECT 74.490 156.630 74.745 157.535 ;
        RECT 73.515 156.055 73.870 156.425 ;
        RECT 74.150 156.395 74.320 156.605 ;
        RECT 74.150 156.065 74.405 156.395 ;
        RECT 70.765 155.685 72.125 155.895 ;
        RECT 70.765 155.325 71.095 155.685 ;
        RECT 71.265 155.155 71.595 155.515 ;
        RECT 71.795 155.325 72.125 155.685 ;
        RECT 72.635 155.325 73.345 155.915 ;
        RECT 74.150 155.875 74.320 156.065 ;
        RECT 74.575 155.900 74.745 156.630 ;
        RECT 74.920 156.555 75.180 157.705 ;
        RECT 75.815 156.615 77.485 157.705 ;
        RECT 75.815 156.095 76.565 156.615 ;
        RECT 77.695 156.565 77.925 157.705 ;
        RECT 78.095 156.555 78.425 157.535 ;
        RECT 78.595 156.565 78.805 157.705 ;
        RECT 79.150 157.075 79.435 157.535 ;
        RECT 79.605 157.245 79.875 157.705 ;
        RECT 79.150 156.855 80.105 157.075 ;
        RECT 73.605 155.705 74.320 155.875 ;
        RECT 73.605 155.325 73.775 155.705 ;
        RECT 73.990 155.155 74.320 155.535 ;
        RECT 74.490 155.325 74.745 155.900 ;
        RECT 74.920 155.155 75.180 155.995 ;
        RECT 76.735 155.925 77.485 156.445 ;
        RECT 77.675 156.145 78.005 156.395 ;
        RECT 75.815 155.155 77.485 155.925 ;
        RECT 77.695 155.155 77.925 155.975 ;
        RECT 78.175 155.955 78.425 156.555 ;
        RECT 79.035 156.125 79.725 156.685 ;
        RECT 78.095 155.325 78.425 155.955 ;
        RECT 78.595 155.155 78.805 155.975 ;
        RECT 79.895 155.955 80.105 156.855 ;
        RECT 79.150 155.785 80.105 155.955 ;
        RECT 80.275 156.685 80.675 157.535 ;
        RECT 80.865 157.075 81.145 157.535 ;
        RECT 81.665 157.245 81.990 157.705 ;
        RECT 80.865 156.855 81.990 157.075 ;
        RECT 80.275 156.125 81.370 156.685 ;
        RECT 81.540 156.395 81.990 156.855 ;
        RECT 82.160 156.565 82.545 157.535 ;
        RECT 79.150 155.325 79.435 155.785 ;
        RECT 79.605 155.155 79.875 155.615 ;
        RECT 80.275 155.325 80.675 156.125 ;
        RECT 81.540 156.065 82.095 156.395 ;
        RECT 81.540 155.955 81.990 156.065 ;
        RECT 80.865 155.785 81.990 155.955 ;
        RECT 82.265 155.895 82.545 156.565 ;
        RECT 82.715 156.945 83.230 157.355 ;
        RECT 83.465 156.945 83.635 157.705 ;
        RECT 83.805 157.365 85.835 157.535 ;
        RECT 82.715 156.135 83.055 156.945 ;
        RECT 83.805 156.700 83.975 157.365 ;
        RECT 84.370 157.025 85.495 157.195 ;
        RECT 83.225 156.510 83.975 156.700 ;
        RECT 84.145 156.685 85.155 156.855 ;
        RECT 82.715 155.965 83.945 156.135 ;
        RECT 80.865 155.325 81.145 155.785 ;
        RECT 81.665 155.155 81.990 155.615 ;
        RECT 82.160 155.325 82.545 155.895 ;
        RECT 82.990 155.360 83.235 155.965 ;
        RECT 83.455 155.155 83.965 155.690 ;
        RECT 84.145 155.325 84.335 156.685 ;
        RECT 84.505 155.665 84.780 156.485 ;
        RECT 84.985 155.885 85.155 156.685 ;
        RECT 85.325 155.895 85.495 157.025 ;
        RECT 85.665 156.395 85.835 157.365 ;
        RECT 86.005 156.565 86.175 157.705 ;
        RECT 86.345 156.565 86.680 157.535 ;
        RECT 85.665 156.065 85.860 156.395 ;
        RECT 86.085 156.065 86.340 156.395 ;
        RECT 86.085 155.895 86.255 156.065 ;
        RECT 86.510 155.895 86.680 156.565 ;
        RECT 87.315 156.540 87.605 157.705 ;
        RECT 88.240 157.195 89.895 157.485 ;
        RECT 88.240 156.855 89.830 157.025 ;
        RECT 90.065 156.905 90.345 157.705 ;
        RECT 88.240 156.565 88.560 156.855 ;
        RECT 89.660 156.735 89.830 156.855 ;
        RECT 88.755 156.515 89.470 156.685 ;
        RECT 89.660 156.565 90.385 156.735 ;
        RECT 90.555 156.565 90.825 157.535 ;
        RECT 91.000 157.195 92.655 157.485 ;
        RECT 91.000 156.855 92.590 157.025 ;
        RECT 92.825 156.905 93.105 157.705 ;
        RECT 91.000 156.565 91.320 156.855 ;
        RECT 92.420 156.735 92.590 156.855 ;
        RECT 85.325 155.725 86.255 155.895 ;
        RECT 85.325 155.690 85.500 155.725 ;
        RECT 84.505 155.495 84.785 155.665 ;
        RECT 84.505 155.325 84.780 155.495 ;
        RECT 84.970 155.325 85.500 155.690 ;
        RECT 85.925 155.155 86.255 155.555 ;
        RECT 86.425 155.325 86.680 155.895 ;
        RECT 87.315 155.155 87.605 155.880 ;
        RECT 88.240 155.825 88.590 156.395 ;
        RECT 88.760 156.065 89.470 156.515 ;
        RECT 90.215 156.395 90.385 156.565 ;
        RECT 89.640 156.065 90.045 156.395 ;
        RECT 90.215 156.065 90.485 156.395 ;
        RECT 90.215 155.895 90.385 156.065 ;
        RECT 88.775 155.725 90.385 155.895 ;
        RECT 90.655 155.830 90.825 156.565 ;
        RECT 91.515 156.515 92.230 156.685 ;
        RECT 92.420 156.565 93.145 156.735 ;
        RECT 93.315 156.565 93.585 157.535 ;
        RECT 88.245 155.155 88.575 155.655 ;
        RECT 88.775 155.375 88.945 155.725 ;
        RECT 89.145 155.155 89.475 155.555 ;
        RECT 89.645 155.375 89.815 155.725 ;
        RECT 89.985 155.155 90.365 155.555 ;
        RECT 90.555 155.485 90.825 155.830 ;
        RECT 91.000 155.825 91.350 156.395 ;
        RECT 91.520 156.065 92.230 156.515 ;
        RECT 92.975 156.395 93.145 156.565 ;
        RECT 92.400 156.065 92.805 156.395 ;
        RECT 92.975 156.065 93.245 156.395 ;
        RECT 92.975 155.895 93.145 156.065 ;
        RECT 91.535 155.725 93.145 155.895 ;
        RECT 93.415 155.830 93.585 156.565 ;
        RECT 91.005 155.155 91.335 155.655 ;
        RECT 91.535 155.375 91.705 155.725 ;
        RECT 91.905 155.155 92.235 155.555 ;
        RECT 92.405 155.375 92.575 155.725 ;
        RECT 92.745 155.155 93.125 155.555 ;
        RECT 93.315 155.485 93.585 155.830 ;
        RECT 93.755 156.565 94.095 157.535 ;
        RECT 94.265 156.565 94.435 157.705 ;
        RECT 94.705 156.905 94.955 157.705 ;
        RECT 95.600 156.735 95.930 157.535 ;
        RECT 96.230 156.905 96.560 157.705 ;
        RECT 96.730 156.735 97.060 157.535 ;
        RECT 94.625 156.565 97.060 156.735 ;
        RECT 97.895 156.565 98.235 157.535 ;
        RECT 98.405 156.565 98.575 157.705 ;
        RECT 98.845 156.905 99.095 157.705 ;
        RECT 99.740 156.735 100.070 157.535 ;
        RECT 100.370 156.905 100.700 157.705 ;
        RECT 100.870 156.735 101.200 157.535 ;
        RECT 98.765 156.565 101.200 156.735 ;
        RECT 101.575 156.615 102.785 157.705 ;
        RECT 102.955 156.945 103.470 157.355 ;
        RECT 103.705 156.945 103.875 157.705 ;
        RECT 104.045 157.365 106.075 157.535 ;
        RECT 93.755 156.005 93.930 156.565 ;
        RECT 94.625 156.315 94.795 156.565 ;
        RECT 94.100 156.145 94.795 156.315 ;
        RECT 94.965 156.175 95.390 156.345 ;
        RECT 94.970 156.145 95.390 156.175 ;
        RECT 95.560 156.145 95.890 156.345 ;
        RECT 96.060 156.145 96.390 156.345 ;
        RECT 93.755 155.955 93.985 156.005 ;
        RECT 93.755 155.325 94.095 155.955 ;
        RECT 94.265 155.155 94.515 155.955 ;
        RECT 94.705 155.805 95.930 155.975 ;
        RECT 94.705 155.325 95.035 155.805 ;
        RECT 95.205 155.155 95.430 155.615 ;
        RECT 95.600 155.325 95.930 155.805 ;
        RECT 96.560 155.935 96.730 156.565 ;
        RECT 96.915 156.145 97.265 156.395 ;
        RECT 97.895 155.955 98.070 156.565 ;
        RECT 98.765 156.315 98.935 156.565 ;
        RECT 98.240 156.145 98.935 156.315 ;
        RECT 99.110 156.145 99.530 156.345 ;
        RECT 99.700 156.145 100.030 156.345 ;
        RECT 100.200 156.145 100.530 156.345 ;
        RECT 96.560 155.325 97.060 155.935 ;
        RECT 97.895 155.325 98.235 155.955 ;
        RECT 98.405 155.155 98.655 155.955 ;
        RECT 98.845 155.805 100.070 155.975 ;
        RECT 98.845 155.325 99.175 155.805 ;
        RECT 99.345 155.155 99.570 155.615 ;
        RECT 99.740 155.325 100.070 155.805 ;
        RECT 100.700 155.935 100.870 156.565 ;
        RECT 101.055 156.145 101.405 156.395 ;
        RECT 101.575 156.075 102.095 156.615 ;
        RECT 100.700 155.325 101.200 155.935 ;
        RECT 102.265 155.905 102.785 156.445 ;
        RECT 102.955 156.135 103.295 156.945 ;
        RECT 104.045 156.700 104.215 157.365 ;
        RECT 104.610 157.025 105.735 157.195 ;
        RECT 103.465 156.510 104.215 156.700 ;
        RECT 104.385 156.685 105.395 156.855 ;
        RECT 102.955 155.965 104.185 156.135 ;
        RECT 101.575 155.155 102.785 155.905 ;
        RECT 103.230 155.360 103.475 155.965 ;
        RECT 103.695 155.155 104.205 155.690 ;
        RECT 104.385 155.325 104.575 156.685 ;
        RECT 104.745 156.345 105.020 156.485 ;
        RECT 104.745 156.175 105.025 156.345 ;
        RECT 104.745 155.325 105.020 156.175 ;
        RECT 105.225 155.885 105.395 156.685 ;
        RECT 105.565 155.895 105.735 157.025 ;
        RECT 105.905 156.395 106.075 157.365 ;
        RECT 106.245 156.565 106.415 157.705 ;
        RECT 106.585 156.565 106.920 157.535 ;
        RECT 107.210 157.075 107.495 157.535 ;
        RECT 107.665 157.245 107.935 157.705 ;
        RECT 107.210 156.855 108.165 157.075 ;
        RECT 105.905 156.065 106.100 156.395 ;
        RECT 106.325 156.065 106.580 156.395 ;
        RECT 106.325 155.895 106.495 156.065 ;
        RECT 106.750 155.895 106.920 156.565 ;
        RECT 107.095 156.125 107.785 156.685 ;
        RECT 107.955 155.955 108.165 156.855 ;
        RECT 105.565 155.725 106.495 155.895 ;
        RECT 105.565 155.690 105.740 155.725 ;
        RECT 105.210 155.325 105.740 155.690 ;
        RECT 106.165 155.155 106.495 155.555 ;
        RECT 106.665 155.325 106.920 155.895 ;
        RECT 107.210 155.785 108.165 155.955 ;
        RECT 108.335 156.685 108.735 157.535 ;
        RECT 108.925 157.075 109.205 157.535 ;
        RECT 109.725 157.245 110.050 157.705 ;
        RECT 108.925 156.855 110.050 157.075 ;
        RECT 108.335 156.125 109.430 156.685 ;
        RECT 109.600 156.395 110.050 156.855 ;
        RECT 110.220 156.565 110.605 157.535 ;
        RECT 107.210 155.325 107.495 155.785 ;
        RECT 107.665 155.155 107.935 155.615 ;
        RECT 108.335 155.325 108.735 156.125 ;
        RECT 109.600 156.065 110.155 156.395 ;
        RECT 109.600 155.955 110.050 156.065 ;
        RECT 108.925 155.785 110.050 155.955 ;
        RECT 110.325 155.895 110.605 156.565 ;
        RECT 108.925 155.325 109.205 155.785 ;
        RECT 109.725 155.155 110.050 155.615 ;
        RECT 110.220 155.325 110.605 155.895 ;
        RECT 110.775 156.630 111.045 157.535 ;
        RECT 111.215 156.945 111.545 157.705 ;
        RECT 111.725 156.775 111.895 157.535 ;
        RECT 110.775 155.830 110.945 156.630 ;
        RECT 111.230 156.605 111.895 156.775 ;
        RECT 112.155 156.615 113.365 157.705 ;
        RECT 111.230 156.460 111.400 156.605 ;
        RECT 111.115 156.130 111.400 156.460 ;
        RECT 111.230 155.875 111.400 156.130 ;
        RECT 111.635 156.055 111.965 156.425 ;
        RECT 112.155 156.075 112.675 156.615 ;
        RECT 112.845 155.905 113.365 156.445 ;
        RECT 110.775 155.325 111.035 155.830 ;
        RECT 111.230 155.705 111.895 155.875 ;
        RECT 111.215 155.155 111.545 155.535 ;
        RECT 111.725 155.325 111.895 155.705 ;
        RECT 112.155 155.155 113.365 155.905 ;
        RECT 22.830 154.985 113.450 155.155 ;
        RECT 22.915 154.235 24.125 154.985 ;
        RECT 22.915 153.695 23.435 154.235 ;
        RECT 24.755 154.215 26.425 154.985 ;
        RECT 23.605 153.525 24.125 154.065 ;
        RECT 22.915 152.435 24.125 153.525 ;
        RECT 24.755 153.525 25.505 154.045 ;
        RECT 25.675 153.695 26.425 154.215 ;
        RECT 26.635 154.165 26.865 154.985 ;
        RECT 27.035 154.185 27.365 154.815 ;
        RECT 26.615 153.745 26.945 153.995 ;
        RECT 27.115 153.585 27.365 154.185 ;
        RECT 27.535 154.165 27.745 154.985 ;
        RECT 28.250 154.175 28.495 154.780 ;
        RECT 28.715 154.450 29.225 154.985 ;
        RECT 24.755 152.435 26.425 153.525 ;
        RECT 26.635 152.435 26.865 153.575 ;
        RECT 27.035 152.605 27.365 153.585 ;
        RECT 27.975 154.005 29.205 154.175 ;
        RECT 27.535 152.435 27.745 153.575 ;
        RECT 27.975 153.195 28.315 154.005 ;
        RECT 28.485 153.440 29.235 153.630 ;
        RECT 27.975 152.785 28.490 153.195 ;
        RECT 28.725 152.435 28.895 153.195 ;
        RECT 29.065 152.775 29.235 153.440 ;
        RECT 29.405 153.455 29.595 154.815 ;
        RECT 29.765 153.965 30.040 154.815 ;
        RECT 30.230 154.450 30.760 154.815 ;
        RECT 31.185 154.585 31.515 154.985 ;
        RECT 30.585 154.415 30.760 154.450 ;
        RECT 29.765 153.795 30.045 153.965 ;
        RECT 29.765 153.655 30.040 153.795 ;
        RECT 30.245 153.455 30.415 154.255 ;
        RECT 29.405 153.285 30.415 153.455 ;
        RECT 30.585 154.245 31.515 154.415 ;
        RECT 31.685 154.245 31.940 154.815 ;
        RECT 30.585 153.115 30.755 154.245 ;
        RECT 31.345 154.075 31.515 154.245 ;
        RECT 29.630 152.945 30.755 153.115 ;
        RECT 30.925 153.745 31.120 154.075 ;
        RECT 31.345 153.745 31.600 154.075 ;
        RECT 30.925 152.775 31.095 153.745 ;
        RECT 31.770 153.575 31.940 154.245 ;
        RECT 32.575 154.215 35.165 154.985 ;
        RECT 29.065 152.605 31.095 152.775 ;
        RECT 31.265 152.435 31.435 153.575 ;
        RECT 31.605 152.605 31.940 153.575 ;
        RECT 32.575 153.525 33.785 154.045 ;
        RECT 33.955 153.695 35.165 154.215 ;
        RECT 35.335 154.310 35.605 154.655 ;
        RECT 35.795 154.585 36.175 154.985 ;
        RECT 36.345 154.415 36.515 154.765 ;
        RECT 36.685 154.585 37.015 154.985 ;
        RECT 37.215 154.415 37.385 154.765 ;
        RECT 37.585 154.485 37.915 154.985 ;
        RECT 35.335 153.575 35.505 154.310 ;
        RECT 35.775 154.245 37.385 154.415 ;
        RECT 35.775 154.075 35.945 154.245 ;
        RECT 35.675 153.745 35.945 154.075 ;
        RECT 36.115 153.745 36.520 154.075 ;
        RECT 35.775 153.575 35.945 153.745 ;
        RECT 32.575 152.435 35.165 153.525 ;
        RECT 35.335 152.605 35.605 153.575 ;
        RECT 35.775 153.405 36.500 153.575 ;
        RECT 36.690 153.455 37.400 154.075 ;
        RECT 37.570 153.745 37.920 154.315 ;
        RECT 38.095 154.185 38.435 154.815 ;
        RECT 38.605 154.185 38.855 154.985 ;
        RECT 39.045 154.335 39.375 154.815 ;
        RECT 39.545 154.525 39.770 154.985 ;
        RECT 39.940 154.335 40.270 154.815 ;
        RECT 38.095 154.135 38.325 154.185 ;
        RECT 39.045 154.165 40.270 154.335 ;
        RECT 40.900 154.205 41.400 154.815 ;
        RECT 41.785 154.485 42.115 154.985 ;
        RECT 42.315 154.415 42.485 154.765 ;
        RECT 42.685 154.585 43.015 154.985 ;
        RECT 43.185 154.415 43.355 154.765 ;
        RECT 43.525 154.585 43.905 154.985 ;
        RECT 38.095 153.575 38.270 154.135 ;
        RECT 38.440 153.825 39.135 153.995 ;
        RECT 38.965 153.575 39.135 153.825 ;
        RECT 39.310 153.795 39.730 153.995 ;
        RECT 39.900 153.795 40.230 153.995 ;
        RECT 40.400 153.795 40.730 153.995 ;
        RECT 40.900 153.575 41.070 154.205 ;
        RECT 41.255 153.745 41.605 153.995 ;
        RECT 41.780 153.745 42.130 154.315 ;
        RECT 42.315 154.245 43.925 154.415 ;
        RECT 44.095 154.310 44.365 154.655 ;
        RECT 43.755 154.075 43.925 154.245 ;
        RECT 42.300 153.625 43.010 154.075 ;
        RECT 43.180 153.745 43.585 154.075 ;
        RECT 43.755 153.745 44.025 154.075 ;
        RECT 36.330 153.285 36.500 153.405 ;
        RECT 37.600 153.285 37.920 153.575 ;
        RECT 35.815 152.435 36.095 153.235 ;
        RECT 36.330 153.115 37.920 153.285 ;
        RECT 36.265 152.655 37.920 152.945 ;
        RECT 38.095 152.605 38.435 153.575 ;
        RECT 38.605 152.435 38.775 153.575 ;
        RECT 38.965 153.405 41.400 153.575 ;
        RECT 39.045 152.435 39.295 153.235 ;
        RECT 39.940 152.605 40.270 153.405 ;
        RECT 40.570 152.435 40.900 153.235 ;
        RECT 41.070 152.605 41.400 153.405 ;
        RECT 41.780 153.285 42.100 153.575 ;
        RECT 42.295 153.455 43.010 153.625 ;
        RECT 43.755 153.575 43.925 153.745 ;
        RECT 44.195 153.575 44.365 154.310 ;
        RECT 44.810 154.175 45.055 154.780 ;
        RECT 45.275 154.450 45.785 154.985 ;
        RECT 43.200 153.405 43.925 153.575 ;
        RECT 43.200 153.285 43.370 153.405 ;
        RECT 41.780 153.115 43.370 153.285 ;
        RECT 41.780 152.655 43.435 152.945 ;
        RECT 43.605 152.435 43.885 153.235 ;
        RECT 44.095 152.605 44.365 153.575 ;
        RECT 44.535 154.005 45.765 154.175 ;
        RECT 44.535 153.195 44.875 154.005 ;
        RECT 45.045 153.440 45.795 153.630 ;
        RECT 44.535 152.785 45.050 153.195 ;
        RECT 45.285 152.435 45.455 153.195 ;
        RECT 45.625 152.775 45.795 153.440 ;
        RECT 45.965 153.455 46.155 154.815 ;
        RECT 46.325 153.965 46.600 154.815 ;
        RECT 46.790 154.450 47.320 154.815 ;
        RECT 47.745 154.585 48.075 154.985 ;
        RECT 47.145 154.415 47.320 154.450 ;
        RECT 46.325 153.795 46.605 153.965 ;
        RECT 46.325 153.655 46.600 153.795 ;
        RECT 46.805 153.455 46.975 154.255 ;
        RECT 45.965 153.285 46.975 153.455 ;
        RECT 47.145 154.245 48.075 154.415 ;
        RECT 48.245 154.245 48.500 154.815 ;
        RECT 48.675 154.260 48.965 154.985 ;
        RECT 47.145 153.115 47.315 154.245 ;
        RECT 47.905 154.075 48.075 154.245 ;
        RECT 46.190 152.945 47.315 153.115 ;
        RECT 47.485 153.745 47.680 154.075 ;
        RECT 47.905 153.745 48.160 154.075 ;
        RECT 47.485 152.775 47.655 153.745 ;
        RECT 48.330 153.575 48.500 154.245 ;
        RECT 49.135 154.185 49.475 154.815 ;
        RECT 49.645 154.185 49.895 154.985 ;
        RECT 50.085 154.335 50.415 154.815 ;
        RECT 50.585 154.525 50.810 154.985 ;
        RECT 50.980 154.335 51.310 154.815 ;
        RECT 45.625 152.605 47.655 152.775 ;
        RECT 47.825 152.435 47.995 153.575 ;
        RECT 48.165 152.605 48.500 153.575 ;
        RECT 48.675 152.435 48.965 153.600 ;
        RECT 49.135 153.575 49.310 154.185 ;
        RECT 50.085 154.165 51.310 154.335 ;
        RECT 51.940 154.205 52.440 154.815 ;
        RECT 53.365 154.435 53.535 154.815 ;
        RECT 53.715 154.605 54.045 154.985 ;
        RECT 53.365 154.265 54.030 154.435 ;
        RECT 54.225 154.310 54.485 154.815 ;
        RECT 49.480 153.825 50.175 153.995 ;
        RECT 50.005 153.575 50.175 153.825 ;
        RECT 50.350 153.795 50.770 153.995 ;
        RECT 50.940 153.795 51.270 153.995 ;
        RECT 51.440 153.795 51.770 153.995 ;
        RECT 51.940 153.575 52.110 154.205 ;
        RECT 52.295 153.745 52.645 153.995 ;
        RECT 53.295 153.715 53.625 154.085 ;
        RECT 53.860 154.010 54.030 154.265 ;
        RECT 53.860 153.680 54.145 154.010 ;
        RECT 49.135 152.605 49.475 153.575 ;
        RECT 49.645 152.435 49.815 153.575 ;
        RECT 50.005 153.405 52.440 153.575 ;
        RECT 53.860 153.535 54.030 153.680 ;
        RECT 50.085 152.435 50.335 153.235 ;
        RECT 50.980 152.605 51.310 153.405 ;
        RECT 51.610 152.435 51.940 153.235 ;
        RECT 52.110 152.605 52.440 153.405 ;
        RECT 53.365 153.365 54.030 153.535 ;
        RECT 54.315 153.510 54.485 154.310 ;
        RECT 53.365 152.605 53.535 153.365 ;
        RECT 53.715 152.435 54.045 153.195 ;
        RECT 54.215 152.605 54.485 153.510 ;
        RECT 55.030 154.275 55.285 154.805 ;
        RECT 55.465 154.525 55.750 154.985 ;
        RECT 55.030 153.415 55.210 154.275 ;
        RECT 55.930 154.075 56.180 154.725 ;
        RECT 55.380 153.745 56.180 154.075 ;
        RECT 55.030 153.285 55.285 153.415 ;
        RECT 54.945 153.115 55.285 153.285 ;
        RECT 55.030 152.745 55.285 153.115 ;
        RECT 55.465 152.435 55.750 153.235 ;
        RECT 55.930 153.155 56.180 153.745 ;
        RECT 56.380 154.390 56.700 154.720 ;
        RECT 56.880 154.505 57.540 154.985 ;
        RECT 57.740 154.595 58.590 154.765 ;
        RECT 56.380 153.495 56.570 154.390 ;
        RECT 56.890 154.065 57.550 154.335 ;
        RECT 57.220 154.005 57.550 154.065 ;
        RECT 56.740 153.835 57.070 153.895 ;
        RECT 57.740 153.835 57.910 154.595 ;
        RECT 59.150 154.525 59.470 154.985 ;
        RECT 59.670 154.345 59.920 154.775 ;
        RECT 60.210 154.545 60.620 154.985 ;
        RECT 60.790 154.605 61.805 154.805 ;
        RECT 58.080 154.175 59.330 154.345 ;
        RECT 58.080 154.055 58.410 154.175 ;
        RECT 56.740 153.665 58.640 153.835 ;
        RECT 56.380 153.325 58.300 153.495 ;
        RECT 56.380 153.305 56.700 153.325 ;
        RECT 55.930 152.645 56.260 153.155 ;
        RECT 56.530 152.695 56.700 153.305 ;
        RECT 58.470 153.155 58.640 153.665 ;
        RECT 58.810 153.595 58.990 154.005 ;
        RECT 59.160 153.415 59.330 154.175 ;
        RECT 56.870 152.435 57.200 153.125 ;
        RECT 57.430 152.985 58.640 153.155 ;
        RECT 58.810 153.105 59.330 153.415 ;
        RECT 59.500 154.005 59.920 154.345 ;
        RECT 60.210 154.005 60.620 154.335 ;
        RECT 59.500 153.235 59.690 154.005 ;
        RECT 60.790 153.875 60.960 154.605 ;
        RECT 62.105 154.435 62.275 154.765 ;
        RECT 62.445 154.605 62.775 154.985 ;
        RECT 61.130 154.055 61.480 154.425 ;
        RECT 60.790 153.835 61.210 153.875 ;
        RECT 59.860 153.665 61.210 153.835 ;
        RECT 59.860 153.505 60.110 153.665 ;
        RECT 60.620 153.235 60.870 153.495 ;
        RECT 59.500 152.985 60.870 153.235 ;
        RECT 57.430 152.695 57.670 152.985 ;
        RECT 58.470 152.905 58.640 152.985 ;
        RECT 57.870 152.435 58.290 152.815 ;
        RECT 58.470 152.655 59.100 152.905 ;
        RECT 59.570 152.435 59.900 152.815 ;
        RECT 60.070 152.695 60.240 152.985 ;
        RECT 61.040 152.820 61.210 153.665 ;
        RECT 61.660 153.495 61.880 154.365 ;
        RECT 62.105 154.245 62.800 154.435 ;
        RECT 61.380 153.115 61.880 153.495 ;
        RECT 62.050 153.445 62.460 154.065 ;
        RECT 62.630 153.275 62.800 154.245 ;
        RECT 62.105 153.105 62.800 153.275 ;
        RECT 60.420 152.435 60.800 152.815 ;
        RECT 61.040 152.650 61.870 152.820 ;
        RECT 62.105 152.605 62.275 153.105 ;
        RECT 62.445 152.435 62.775 152.935 ;
        RECT 62.990 152.605 63.215 154.725 ;
        RECT 63.385 154.605 63.715 154.985 ;
        RECT 63.885 154.435 64.055 154.725 ;
        RECT 63.390 154.265 64.055 154.435 ;
        RECT 64.315 154.485 64.575 154.815 ;
        RECT 64.745 154.625 65.075 154.985 ;
        RECT 65.330 154.605 66.630 154.815 ;
        RECT 63.390 153.275 63.620 154.265 ;
        RECT 63.790 153.445 64.140 154.095 ;
        RECT 64.315 153.285 64.485 154.485 ;
        RECT 65.330 154.455 65.500 154.605 ;
        RECT 64.745 154.330 65.500 154.455 ;
        RECT 64.655 154.285 65.500 154.330 ;
        RECT 64.655 154.165 64.925 154.285 ;
        RECT 64.655 153.590 64.825 154.165 ;
        RECT 65.055 153.725 65.465 154.030 ;
        RECT 65.755 153.995 65.965 154.395 ;
        RECT 65.635 153.785 65.965 153.995 ;
        RECT 66.210 153.995 66.430 154.395 ;
        RECT 66.905 154.220 67.360 154.985 ;
        RECT 67.595 154.505 67.875 154.985 ;
        RECT 68.045 154.335 68.305 154.725 ;
        RECT 68.480 154.505 68.735 154.985 ;
        RECT 68.905 154.335 69.200 154.725 ;
        RECT 69.380 154.505 69.655 154.985 ;
        RECT 69.825 154.485 70.125 154.815 ;
        RECT 67.550 154.165 69.200 154.335 ;
        RECT 66.210 153.785 66.685 153.995 ;
        RECT 66.875 153.795 67.365 153.995 ;
        RECT 67.550 153.655 67.955 154.165 ;
        RECT 68.125 153.825 69.265 153.995 ;
        RECT 64.655 153.555 64.855 153.590 ;
        RECT 66.185 153.555 67.360 153.615 ;
        RECT 64.655 153.445 67.360 153.555 ;
        RECT 67.550 153.485 68.305 153.655 ;
        RECT 64.715 153.385 66.515 153.445 ;
        RECT 66.185 153.355 66.515 153.385 ;
        RECT 63.390 153.105 64.055 153.275 ;
        RECT 63.385 152.435 63.715 152.935 ;
        RECT 63.885 152.605 64.055 153.105 ;
        RECT 64.315 152.605 64.575 153.285 ;
        RECT 64.745 152.435 64.995 153.215 ;
        RECT 65.245 153.185 66.080 153.195 ;
        RECT 66.670 153.185 66.855 153.275 ;
        RECT 65.245 152.985 66.855 153.185 ;
        RECT 65.245 152.605 65.495 152.985 ;
        RECT 66.625 152.945 66.855 152.985 ;
        RECT 67.105 152.825 67.360 153.445 ;
        RECT 65.665 152.435 66.020 152.815 ;
        RECT 67.025 152.605 67.360 152.825 ;
        RECT 67.590 152.435 67.875 153.305 ;
        RECT 68.045 153.235 68.305 153.485 ;
        RECT 69.095 153.575 69.265 153.825 ;
        RECT 69.435 153.745 69.785 154.315 ;
        RECT 69.955 153.575 70.125 154.485 ;
        RECT 70.295 154.235 71.505 154.985 ;
        RECT 69.095 153.405 70.125 153.575 ;
        RECT 68.045 153.065 69.165 153.235 ;
        RECT 68.045 152.605 68.305 153.065 ;
        RECT 68.480 152.435 68.735 152.895 ;
        RECT 68.905 152.605 69.165 153.065 ;
        RECT 69.335 152.435 69.645 153.235 ;
        RECT 69.815 152.605 70.125 153.405 ;
        RECT 70.295 153.525 70.815 154.065 ;
        RECT 70.985 153.695 71.505 154.235 ;
        RECT 71.675 154.485 71.975 154.815 ;
        RECT 72.145 154.505 72.420 154.985 ;
        RECT 71.675 153.575 71.845 154.485 ;
        RECT 72.600 154.335 72.895 154.725 ;
        RECT 73.065 154.505 73.320 154.985 ;
        RECT 73.495 154.335 73.755 154.725 ;
        RECT 73.925 154.505 74.205 154.985 ;
        RECT 72.015 153.745 72.365 154.315 ;
        RECT 72.600 154.165 74.250 154.335 ;
        RECT 74.435 154.260 74.725 154.985 ;
        RECT 75.355 154.215 77.025 154.985 ;
        RECT 72.535 153.825 73.675 153.995 ;
        RECT 72.535 153.575 72.705 153.825 ;
        RECT 73.845 153.655 74.250 154.165 ;
        RECT 70.295 152.435 71.505 153.525 ;
        RECT 71.675 153.405 72.705 153.575 ;
        RECT 73.495 153.485 74.250 153.655 ;
        RECT 71.675 152.605 71.985 153.405 ;
        RECT 73.495 153.235 73.755 153.485 ;
        RECT 72.155 152.435 72.465 153.235 ;
        RECT 72.635 153.065 73.755 153.235 ;
        RECT 72.635 152.605 72.895 153.065 ;
        RECT 73.065 152.435 73.320 152.895 ;
        RECT 73.495 152.605 73.755 153.065 ;
        RECT 73.925 152.435 74.210 153.305 ;
        RECT 74.435 152.435 74.725 153.600 ;
        RECT 75.355 153.525 76.105 154.045 ;
        RECT 76.275 153.695 77.025 154.215 ;
        RECT 77.570 154.275 77.825 154.805 ;
        RECT 78.005 154.525 78.290 154.985 ;
        RECT 75.355 152.435 77.025 153.525 ;
        RECT 77.570 153.415 77.750 154.275 ;
        RECT 78.470 154.075 78.720 154.725 ;
        RECT 77.920 153.745 78.720 154.075 ;
        RECT 77.570 152.945 77.825 153.415 ;
        RECT 77.485 152.775 77.825 152.945 ;
        RECT 77.570 152.745 77.825 152.775 ;
        RECT 78.005 152.435 78.290 153.235 ;
        RECT 78.470 153.155 78.720 153.745 ;
        RECT 78.920 154.390 79.240 154.720 ;
        RECT 79.420 154.505 80.080 154.985 ;
        RECT 80.280 154.595 81.130 154.765 ;
        RECT 78.920 153.495 79.110 154.390 ;
        RECT 79.430 154.065 80.090 154.335 ;
        RECT 79.760 154.005 80.090 154.065 ;
        RECT 79.280 153.835 79.610 153.895 ;
        RECT 80.280 153.835 80.450 154.595 ;
        RECT 81.690 154.525 82.010 154.985 ;
        RECT 82.210 154.345 82.460 154.775 ;
        RECT 82.750 154.545 83.160 154.985 ;
        RECT 83.330 154.605 84.345 154.805 ;
        RECT 80.620 154.175 81.870 154.345 ;
        RECT 80.620 154.055 80.950 154.175 ;
        RECT 79.280 153.665 81.180 153.835 ;
        RECT 78.920 153.325 80.840 153.495 ;
        RECT 78.920 153.305 79.240 153.325 ;
        RECT 78.470 152.645 78.800 153.155 ;
        RECT 79.070 152.695 79.240 153.305 ;
        RECT 81.010 153.155 81.180 153.665 ;
        RECT 81.350 153.595 81.530 154.005 ;
        RECT 81.700 153.415 81.870 154.175 ;
        RECT 79.410 152.435 79.740 153.125 ;
        RECT 79.970 152.985 81.180 153.155 ;
        RECT 81.350 153.105 81.870 153.415 ;
        RECT 82.040 154.005 82.460 154.345 ;
        RECT 82.750 154.005 83.160 154.335 ;
        RECT 82.040 153.235 82.230 154.005 ;
        RECT 83.330 153.875 83.500 154.605 ;
        RECT 84.645 154.435 84.815 154.765 ;
        RECT 84.985 154.605 85.315 154.985 ;
        RECT 83.670 154.055 84.020 154.425 ;
        RECT 83.330 153.835 83.750 153.875 ;
        RECT 82.400 153.665 83.750 153.835 ;
        RECT 82.400 153.505 82.650 153.665 ;
        RECT 83.160 153.235 83.410 153.495 ;
        RECT 82.040 152.985 83.410 153.235 ;
        RECT 79.970 152.695 80.210 152.985 ;
        RECT 81.010 152.905 81.180 152.985 ;
        RECT 80.410 152.435 80.830 152.815 ;
        RECT 81.010 152.655 81.640 152.905 ;
        RECT 82.110 152.435 82.440 152.815 ;
        RECT 82.610 152.695 82.780 152.985 ;
        RECT 83.580 152.820 83.750 153.665 ;
        RECT 84.200 153.495 84.420 154.365 ;
        RECT 84.645 154.245 85.340 154.435 ;
        RECT 83.920 153.115 84.420 153.495 ;
        RECT 84.590 153.445 85.000 154.065 ;
        RECT 85.170 153.275 85.340 154.245 ;
        RECT 84.645 153.105 85.340 153.275 ;
        RECT 82.960 152.435 83.340 152.815 ;
        RECT 83.580 152.650 84.410 152.820 ;
        RECT 84.645 152.605 84.815 153.105 ;
        RECT 84.985 152.435 85.315 152.935 ;
        RECT 85.530 152.605 85.755 154.725 ;
        RECT 85.925 154.605 86.255 154.985 ;
        RECT 86.425 154.435 86.595 154.725 ;
        RECT 85.930 154.265 86.595 154.435 ;
        RECT 87.865 154.435 88.035 154.815 ;
        RECT 88.215 154.605 88.545 154.985 ;
        RECT 87.865 154.265 88.530 154.435 ;
        RECT 88.725 154.310 88.985 154.815 ;
        RECT 85.930 153.275 86.160 154.265 ;
        RECT 86.330 153.445 86.680 154.095 ;
        RECT 87.795 153.715 88.125 154.085 ;
        RECT 88.360 154.010 88.530 154.265 ;
        RECT 88.360 153.680 88.645 154.010 ;
        RECT 88.360 153.535 88.530 153.680 ;
        RECT 87.865 153.365 88.530 153.535 ;
        RECT 88.815 153.510 88.985 154.310 ;
        RECT 89.155 154.215 92.665 154.985 ;
        RECT 85.930 153.105 86.595 153.275 ;
        RECT 85.925 152.435 86.255 152.935 ;
        RECT 86.425 152.605 86.595 153.105 ;
        RECT 87.865 152.605 88.035 153.365 ;
        RECT 88.215 152.435 88.545 153.195 ;
        RECT 88.715 152.605 88.985 153.510 ;
        RECT 89.155 153.525 90.845 154.045 ;
        RECT 91.015 153.695 92.665 154.215 ;
        RECT 92.835 154.310 93.105 154.655 ;
        RECT 93.295 154.585 93.675 154.985 ;
        RECT 93.845 154.415 94.015 154.765 ;
        RECT 94.185 154.585 94.515 154.985 ;
        RECT 94.715 154.415 94.885 154.765 ;
        RECT 95.085 154.485 95.415 154.985 ;
        RECT 92.835 153.575 93.005 154.310 ;
        RECT 93.275 154.245 94.885 154.415 ;
        RECT 93.275 154.075 93.445 154.245 ;
        RECT 93.175 153.745 93.445 154.075 ;
        RECT 93.615 153.745 94.020 154.075 ;
        RECT 93.275 153.575 93.445 153.745 ;
        RECT 89.155 152.435 92.665 153.525 ;
        RECT 92.835 152.605 93.105 153.575 ;
        RECT 93.275 153.405 94.000 153.575 ;
        RECT 94.190 153.455 94.900 154.075 ;
        RECT 95.070 153.745 95.420 154.315 ;
        RECT 95.595 154.310 95.865 154.655 ;
        RECT 96.055 154.585 96.435 154.985 ;
        RECT 96.605 154.415 96.775 154.765 ;
        RECT 96.945 154.585 97.275 154.985 ;
        RECT 97.475 154.415 97.645 154.765 ;
        RECT 97.845 154.485 98.175 154.985 ;
        RECT 95.595 153.575 95.765 154.310 ;
        RECT 96.035 154.245 97.645 154.415 ;
        RECT 96.035 154.075 96.205 154.245 ;
        RECT 95.935 153.745 96.205 154.075 ;
        RECT 96.375 153.745 96.780 154.075 ;
        RECT 96.035 153.575 96.205 153.745 ;
        RECT 96.950 153.625 97.660 154.075 ;
        RECT 97.830 153.745 98.180 154.315 ;
        RECT 98.355 154.215 100.025 154.985 ;
        RECT 100.195 154.260 100.485 154.985 ;
        RECT 93.830 153.285 94.000 153.405 ;
        RECT 95.100 153.285 95.420 153.575 ;
        RECT 93.315 152.435 93.595 153.235 ;
        RECT 93.830 153.115 95.420 153.285 ;
        RECT 93.765 152.655 95.420 152.945 ;
        RECT 95.595 152.605 95.865 153.575 ;
        RECT 96.035 153.405 96.760 153.575 ;
        RECT 96.950 153.455 97.665 153.625 ;
        RECT 96.590 153.285 96.760 153.405 ;
        RECT 97.860 153.285 98.180 153.575 ;
        RECT 96.075 152.435 96.355 153.235 ;
        RECT 96.590 153.115 98.180 153.285 ;
        RECT 98.355 153.525 99.105 154.045 ;
        RECT 99.275 153.695 100.025 154.215 ;
        RECT 101.155 154.165 101.385 154.985 ;
        RECT 101.555 154.185 101.885 154.815 ;
        RECT 101.135 153.745 101.465 153.995 ;
        RECT 96.525 152.655 98.180 152.945 ;
        RECT 98.355 152.435 100.025 153.525 ;
        RECT 100.195 152.435 100.485 153.600 ;
        RECT 101.635 153.585 101.885 154.185 ;
        RECT 102.055 154.165 102.265 154.985 ;
        RECT 102.870 154.275 103.125 154.805 ;
        RECT 103.305 154.525 103.590 154.985 ;
        RECT 101.155 152.435 101.385 153.575 ;
        RECT 101.555 152.605 101.885 153.585 ;
        RECT 102.055 152.435 102.265 153.575 ;
        RECT 102.870 153.415 103.050 154.275 ;
        RECT 103.770 154.075 104.020 154.725 ;
        RECT 103.220 153.745 104.020 154.075 ;
        RECT 102.870 152.945 103.125 153.415 ;
        RECT 102.785 152.775 103.125 152.945 ;
        RECT 102.870 152.745 103.125 152.775 ;
        RECT 103.305 152.435 103.590 153.235 ;
        RECT 103.770 153.155 104.020 153.745 ;
        RECT 104.220 154.390 104.540 154.720 ;
        RECT 104.720 154.505 105.380 154.985 ;
        RECT 105.580 154.595 106.430 154.765 ;
        RECT 104.220 153.495 104.410 154.390 ;
        RECT 104.730 154.065 105.390 154.335 ;
        RECT 105.060 154.005 105.390 154.065 ;
        RECT 104.580 153.835 104.910 153.895 ;
        RECT 105.580 153.835 105.750 154.595 ;
        RECT 106.990 154.525 107.310 154.985 ;
        RECT 107.510 154.345 107.760 154.775 ;
        RECT 108.050 154.545 108.460 154.985 ;
        RECT 108.630 154.605 109.645 154.805 ;
        RECT 105.920 154.175 107.170 154.345 ;
        RECT 105.920 154.055 106.250 154.175 ;
        RECT 104.580 153.665 106.480 153.835 ;
        RECT 104.220 153.325 106.140 153.495 ;
        RECT 104.220 153.305 104.540 153.325 ;
        RECT 103.770 152.645 104.100 153.155 ;
        RECT 104.370 152.695 104.540 153.305 ;
        RECT 106.310 153.155 106.480 153.665 ;
        RECT 106.650 153.595 106.830 154.005 ;
        RECT 107.000 153.415 107.170 154.175 ;
        RECT 104.710 152.435 105.040 153.125 ;
        RECT 105.270 152.985 106.480 153.155 ;
        RECT 106.650 153.105 107.170 153.415 ;
        RECT 107.340 154.005 107.760 154.345 ;
        RECT 108.050 154.005 108.460 154.335 ;
        RECT 107.340 153.235 107.530 154.005 ;
        RECT 108.630 153.875 108.800 154.605 ;
        RECT 109.945 154.435 110.115 154.765 ;
        RECT 110.285 154.605 110.615 154.985 ;
        RECT 108.970 154.055 109.320 154.425 ;
        RECT 108.630 153.835 109.050 153.875 ;
        RECT 107.700 153.665 109.050 153.835 ;
        RECT 107.700 153.505 107.950 153.665 ;
        RECT 108.460 153.235 108.710 153.495 ;
        RECT 107.340 152.985 108.710 153.235 ;
        RECT 105.270 152.695 105.510 152.985 ;
        RECT 106.310 152.905 106.480 152.985 ;
        RECT 105.710 152.435 106.130 152.815 ;
        RECT 106.310 152.655 106.940 152.905 ;
        RECT 107.410 152.435 107.740 152.815 ;
        RECT 107.910 152.695 108.080 152.985 ;
        RECT 108.880 152.820 109.050 153.665 ;
        RECT 109.500 153.495 109.720 154.365 ;
        RECT 109.945 154.245 110.640 154.435 ;
        RECT 109.220 153.115 109.720 153.495 ;
        RECT 109.890 153.445 110.300 154.065 ;
        RECT 110.470 153.275 110.640 154.245 ;
        RECT 109.945 153.105 110.640 153.275 ;
        RECT 108.260 152.435 108.640 152.815 ;
        RECT 108.880 152.650 109.710 152.820 ;
        RECT 109.945 152.605 110.115 153.105 ;
        RECT 110.285 152.435 110.615 152.935 ;
        RECT 110.830 152.605 111.055 154.725 ;
        RECT 111.225 154.605 111.555 154.985 ;
        RECT 111.725 154.435 111.895 154.725 ;
        RECT 111.230 154.265 111.895 154.435 ;
        RECT 111.230 153.275 111.460 154.265 ;
        RECT 112.155 154.235 113.365 154.985 ;
        RECT 111.630 153.445 111.980 154.095 ;
        RECT 112.155 153.525 112.675 154.065 ;
        RECT 112.845 153.695 113.365 154.235 ;
        RECT 111.230 153.105 111.895 153.275 ;
        RECT 111.225 152.435 111.555 152.935 ;
        RECT 111.725 152.605 111.895 153.105 ;
        RECT 112.155 152.435 113.365 153.525 ;
        RECT 22.830 152.265 113.450 152.435 ;
        RECT 22.915 151.175 24.125 152.265 ;
        RECT 25.130 151.285 25.385 151.955 ;
        RECT 25.565 151.465 25.850 152.265 ;
        RECT 26.030 151.545 26.360 152.055 ;
        RECT 25.130 151.245 25.310 151.285 ;
        RECT 22.915 150.465 23.435 151.005 ;
        RECT 23.605 150.635 24.125 151.175 ;
        RECT 25.045 151.075 25.310 151.245 ;
        RECT 22.915 149.715 24.125 150.465 ;
        RECT 25.130 150.425 25.310 151.075 ;
        RECT 26.030 150.955 26.280 151.545 ;
        RECT 26.630 151.395 26.800 152.005 ;
        RECT 26.970 151.575 27.300 152.265 ;
        RECT 27.530 151.715 27.770 152.005 ;
        RECT 27.970 151.885 28.390 152.265 ;
        RECT 28.570 151.795 29.200 152.045 ;
        RECT 29.670 151.885 30.000 152.265 ;
        RECT 28.570 151.715 28.740 151.795 ;
        RECT 30.170 151.715 30.340 152.005 ;
        RECT 30.520 151.885 30.900 152.265 ;
        RECT 31.140 151.880 31.970 152.050 ;
        RECT 27.530 151.545 28.740 151.715 ;
        RECT 25.480 150.625 26.280 150.955 ;
        RECT 25.130 149.895 25.385 150.425 ;
        RECT 25.565 149.715 25.850 150.175 ;
        RECT 26.030 149.975 26.280 150.625 ;
        RECT 26.480 151.375 26.800 151.395 ;
        RECT 26.480 151.205 28.400 151.375 ;
        RECT 26.480 150.310 26.670 151.205 ;
        RECT 28.570 151.035 28.740 151.545 ;
        RECT 28.910 151.285 29.430 151.595 ;
        RECT 26.840 150.865 28.740 151.035 ;
        RECT 26.840 150.805 27.170 150.865 ;
        RECT 27.320 150.635 27.650 150.695 ;
        RECT 26.990 150.365 27.650 150.635 ;
        RECT 26.480 149.980 26.800 150.310 ;
        RECT 26.980 149.715 27.640 150.195 ;
        RECT 27.840 150.105 28.010 150.865 ;
        RECT 28.910 150.695 29.090 151.105 ;
        RECT 28.180 150.525 28.510 150.645 ;
        RECT 29.260 150.525 29.430 151.285 ;
        RECT 28.180 150.355 29.430 150.525 ;
        RECT 29.600 151.465 30.970 151.715 ;
        RECT 29.600 150.695 29.790 151.465 ;
        RECT 30.720 151.205 30.970 151.465 ;
        RECT 29.960 151.035 30.210 151.195 ;
        RECT 31.140 151.035 31.310 151.880 ;
        RECT 32.205 151.595 32.375 152.095 ;
        RECT 32.545 151.765 32.875 152.265 ;
        RECT 31.480 151.205 31.980 151.585 ;
        RECT 32.205 151.425 32.900 151.595 ;
        RECT 29.960 150.865 31.310 151.035 ;
        RECT 30.890 150.825 31.310 150.865 ;
        RECT 29.600 150.355 30.020 150.695 ;
        RECT 30.310 150.365 30.720 150.695 ;
        RECT 27.840 149.935 28.690 150.105 ;
        RECT 29.250 149.715 29.570 150.175 ;
        RECT 29.770 149.925 30.020 150.355 ;
        RECT 30.310 149.715 30.720 150.155 ;
        RECT 30.890 150.095 31.060 150.825 ;
        RECT 31.230 150.275 31.580 150.645 ;
        RECT 31.760 150.335 31.980 151.205 ;
        RECT 32.150 150.635 32.560 151.255 ;
        RECT 32.730 150.455 32.900 151.425 ;
        RECT 32.205 150.265 32.900 150.455 ;
        RECT 30.890 149.895 31.905 150.095 ;
        RECT 32.205 149.935 32.375 150.265 ;
        RECT 32.545 149.715 32.875 150.095 ;
        RECT 33.090 149.975 33.315 152.095 ;
        RECT 33.485 151.765 33.815 152.265 ;
        RECT 33.985 151.595 34.155 152.095 ;
        RECT 33.490 151.425 34.155 151.595 ;
        RECT 33.490 150.435 33.720 151.425 ;
        RECT 33.890 150.605 34.240 151.255 ;
        RECT 34.415 151.190 34.685 152.095 ;
        RECT 34.855 151.505 35.185 152.265 ;
        RECT 35.365 151.335 35.535 152.095 ;
        RECT 33.490 150.265 34.155 150.435 ;
        RECT 33.485 149.715 33.815 150.095 ;
        RECT 33.985 149.975 34.155 150.265 ;
        RECT 34.415 150.390 34.585 151.190 ;
        RECT 34.870 151.165 35.535 151.335 ;
        RECT 34.870 151.020 35.040 151.165 ;
        RECT 35.795 151.100 36.085 152.265 ;
        RECT 36.255 151.125 36.525 152.095 ;
        RECT 36.735 151.465 37.015 152.265 ;
        RECT 37.185 151.755 38.840 152.045 ;
        RECT 37.250 151.415 38.840 151.585 ;
        RECT 37.250 151.295 37.420 151.415 ;
        RECT 36.695 151.125 37.420 151.295 ;
        RECT 34.755 150.690 35.040 151.020 ;
        RECT 34.870 150.435 35.040 150.690 ;
        RECT 35.275 150.615 35.605 150.985 ;
        RECT 34.415 149.885 34.675 150.390 ;
        RECT 34.870 150.265 35.535 150.435 ;
        RECT 34.855 149.715 35.185 150.095 ;
        RECT 35.365 149.885 35.535 150.265 ;
        RECT 35.795 149.715 36.085 150.440 ;
        RECT 36.255 150.390 36.425 151.125 ;
        RECT 36.695 150.955 36.865 151.125 ;
        RECT 36.595 150.625 36.865 150.955 ;
        RECT 37.035 150.625 37.440 150.955 ;
        RECT 37.610 150.625 38.320 151.245 ;
        RECT 38.520 151.125 38.840 151.415 ;
        RECT 39.015 151.125 39.285 152.095 ;
        RECT 39.495 151.465 39.775 152.265 ;
        RECT 39.945 151.755 41.600 152.045 ;
        RECT 40.010 151.415 41.600 151.585 ;
        RECT 40.010 151.295 40.180 151.415 ;
        RECT 39.455 151.125 40.180 151.295 ;
        RECT 36.695 150.455 36.865 150.625 ;
        RECT 36.255 150.045 36.525 150.390 ;
        RECT 36.695 150.285 38.305 150.455 ;
        RECT 38.490 150.385 38.840 150.955 ;
        RECT 39.015 150.390 39.185 151.125 ;
        RECT 39.455 150.955 39.625 151.125 ;
        RECT 39.355 150.625 39.625 150.955 ;
        RECT 39.795 150.625 40.200 150.955 ;
        RECT 40.370 150.625 41.080 151.245 ;
        RECT 41.280 151.125 41.600 151.415 ;
        RECT 41.775 151.125 42.115 152.095 ;
        RECT 42.285 151.125 42.455 152.265 ;
        RECT 42.725 151.465 42.975 152.265 ;
        RECT 43.620 151.295 43.950 152.095 ;
        RECT 44.250 151.465 44.580 152.265 ;
        RECT 44.750 151.295 45.080 152.095 ;
        RECT 42.645 151.125 45.080 151.295 ;
        RECT 45.455 151.125 45.795 152.095 ;
        RECT 45.965 151.125 46.135 152.265 ;
        RECT 46.405 151.465 46.655 152.265 ;
        RECT 47.300 151.295 47.630 152.095 ;
        RECT 47.930 151.465 48.260 152.265 ;
        RECT 48.430 151.295 48.760 152.095 ;
        RECT 46.325 151.125 48.760 151.295 ;
        RECT 49.595 151.505 50.110 151.915 ;
        RECT 50.345 151.505 50.515 152.265 ;
        RECT 50.685 151.925 52.715 152.095 ;
        RECT 39.455 150.455 39.625 150.625 ;
        RECT 36.715 149.715 37.095 150.115 ;
        RECT 37.265 149.935 37.435 150.285 ;
        RECT 37.605 149.715 37.935 150.115 ;
        RECT 38.135 149.935 38.305 150.285 ;
        RECT 38.505 149.715 38.835 150.215 ;
        RECT 39.015 150.045 39.285 150.390 ;
        RECT 39.455 150.285 41.065 150.455 ;
        RECT 41.250 150.385 41.600 150.955 ;
        RECT 41.775 150.515 41.950 151.125 ;
        RECT 42.645 150.875 42.815 151.125 ;
        RECT 42.120 150.705 42.815 150.875 ;
        RECT 42.990 150.705 43.410 150.905 ;
        RECT 43.580 150.705 43.910 150.905 ;
        RECT 44.080 150.705 44.410 150.905 ;
        RECT 39.475 149.715 39.855 150.115 ;
        RECT 40.025 149.935 40.195 150.285 ;
        RECT 40.365 149.715 40.695 150.115 ;
        RECT 40.895 149.935 41.065 150.285 ;
        RECT 41.265 149.715 41.595 150.215 ;
        RECT 41.775 149.885 42.115 150.515 ;
        RECT 42.285 149.715 42.535 150.515 ;
        RECT 42.725 150.365 43.950 150.535 ;
        RECT 42.725 149.885 43.055 150.365 ;
        RECT 43.225 149.715 43.450 150.175 ;
        RECT 43.620 149.885 43.950 150.365 ;
        RECT 44.580 150.495 44.750 151.125 ;
        RECT 44.935 150.705 45.285 150.955 ;
        RECT 45.455 150.565 45.630 151.125 ;
        RECT 46.325 150.875 46.495 151.125 ;
        RECT 45.800 150.705 46.495 150.875 ;
        RECT 46.670 150.705 47.090 150.905 ;
        RECT 47.260 150.705 47.590 150.905 ;
        RECT 47.760 150.705 48.090 150.905 ;
        RECT 45.455 150.515 45.685 150.565 ;
        RECT 44.580 149.885 45.080 150.495 ;
        RECT 45.455 149.885 45.795 150.515 ;
        RECT 45.965 149.715 46.215 150.515 ;
        RECT 46.405 150.365 47.630 150.535 ;
        RECT 46.405 149.885 46.735 150.365 ;
        RECT 46.905 149.715 47.130 150.175 ;
        RECT 47.300 149.885 47.630 150.365 ;
        RECT 48.260 150.495 48.430 151.125 ;
        RECT 48.615 150.705 48.965 150.955 ;
        RECT 49.595 150.695 49.935 151.505 ;
        RECT 50.685 151.260 50.855 151.925 ;
        RECT 51.250 151.585 52.375 151.755 ;
        RECT 50.105 151.070 50.855 151.260 ;
        RECT 51.025 151.245 52.035 151.415 ;
        RECT 49.595 150.525 50.825 150.695 ;
        RECT 48.260 149.885 48.760 150.495 ;
        RECT 49.870 149.920 50.115 150.525 ;
        RECT 50.335 149.715 50.845 150.250 ;
        RECT 51.025 149.885 51.215 151.245 ;
        RECT 51.385 150.565 51.660 151.045 ;
        RECT 51.385 150.395 51.665 150.565 ;
        RECT 51.865 150.445 52.035 151.245 ;
        RECT 52.205 150.455 52.375 151.585 ;
        RECT 52.545 150.955 52.715 151.925 ;
        RECT 52.885 151.125 53.055 152.265 ;
        RECT 53.225 151.125 53.560 152.095 ;
        RECT 52.545 150.625 52.740 150.955 ;
        RECT 52.965 150.625 53.220 150.955 ;
        RECT 52.965 150.455 53.135 150.625 ;
        RECT 53.390 150.455 53.560 151.125 ;
        RECT 51.385 149.885 51.660 150.395 ;
        RECT 52.205 150.285 53.135 150.455 ;
        RECT 52.205 150.250 52.380 150.285 ;
        RECT 51.850 149.885 52.380 150.250 ;
        RECT 52.805 149.715 53.135 150.115 ;
        RECT 53.305 149.885 53.560 150.455 ;
        RECT 54.195 151.125 54.535 152.095 ;
        RECT 54.705 151.125 54.875 152.265 ;
        RECT 55.145 151.465 55.395 152.265 ;
        RECT 56.040 151.295 56.370 152.095 ;
        RECT 56.670 151.465 57.000 152.265 ;
        RECT 57.170 151.295 57.500 152.095 ;
        RECT 57.990 151.635 58.275 152.095 ;
        RECT 58.445 151.805 58.715 152.265 ;
        RECT 57.990 151.415 58.945 151.635 ;
        RECT 55.065 151.125 57.500 151.295 ;
        RECT 54.195 150.515 54.370 151.125 ;
        RECT 55.065 150.875 55.235 151.125 ;
        RECT 54.540 150.705 55.235 150.875 ;
        RECT 55.410 150.705 55.830 150.905 ;
        RECT 56.000 150.705 56.330 150.905 ;
        RECT 56.500 150.705 56.830 150.905 ;
        RECT 54.195 149.885 54.535 150.515 ;
        RECT 54.705 149.715 54.955 150.515 ;
        RECT 55.145 150.365 56.370 150.535 ;
        RECT 55.145 149.885 55.475 150.365 ;
        RECT 55.645 149.715 55.870 150.175 ;
        RECT 56.040 149.885 56.370 150.365 ;
        RECT 57.000 150.495 57.170 151.125 ;
        RECT 57.355 150.705 57.705 150.955 ;
        RECT 57.875 150.685 58.565 151.245 ;
        RECT 58.735 150.515 58.945 151.415 ;
        RECT 57.000 149.885 57.500 150.495 ;
        RECT 57.990 150.345 58.945 150.515 ;
        RECT 59.115 151.245 59.515 152.095 ;
        RECT 59.705 151.635 59.985 152.095 ;
        RECT 60.505 151.805 60.830 152.265 ;
        RECT 59.705 151.415 60.830 151.635 ;
        RECT 59.115 150.685 60.210 151.245 ;
        RECT 60.380 150.955 60.830 151.415 ;
        RECT 61.000 151.125 61.385 152.095 ;
        RECT 57.990 149.885 58.275 150.345 ;
        RECT 58.445 149.715 58.715 150.175 ;
        RECT 59.115 149.885 59.515 150.685 ;
        RECT 60.380 150.625 60.935 150.955 ;
        RECT 60.380 150.515 60.830 150.625 ;
        RECT 59.705 150.345 60.830 150.515 ;
        RECT 61.105 150.455 61.385 151.125 ;
        RECT 61.555 151.100 61.845 152.265 ;
        RECT 59.705 149.885 59.985 150.345 ;
        RECT 60.505 149.715 60.830 150.175 ;
        RECT 61.000 149.885 61.385 150.455 ;
        RECT 62.020 151.075 62.275 151.955 ;
        RECT 62.445 151.125 62.750 152.265 ;
        RECT 63.090 151.885 63.420 152.265 ;
        RECT 63.600 151.715 63.770 152.005 ;
        RECT 63.940 151.805 64.190 152.265 ;
        RECT 62.970 151.545 63.770 151.715 ;
        RECT 64.360 151.755 65.230 152.095 ;
        RECT 61.555 149.715 61.845 150.440 ;
        RECT 62.020 150.425 62.230 151.075 ;
        RECT 62.970 150.955 63.140 151.545 ;
        RECT 64.360 151.375 64.530 151.755 ;
        RECT 65.465 151.635 65.635 152.095 ;
        RECT 65.805 151.805 66.175 152.265 ;
        RECT 66.470 151.665 66.640 152.005 ;
        RECT 66.810 151.835 67.140 152.265 ;
        RECT 67.375 151.665 67.545 152.005 ;
        RECT 63.310 151.205 64.530 151.375 ;
        RECT 64.700 151.295 65.160 151.585 ;
        RECT 65.465 151.465 66.025 151.635 ;
        RECT 66.470 151.495 67.545 151.665 ;
        RECT 67.715 151.765 68.395 152.095 ;
        RECT 68.610 151.765 68.860 152.095 ;
        RECT 69.030 151.805 69.280 152.265 ;
        RECT 65.855 151.325 66.025 151.465 ;
        RECT 64.700 151.285 65.665 151.295 ;
        RECT 64.360 151.115 64.530 151.205 ;
        RECT 64.990 151.125 65.665 151.285 ;
        RECT 62.400 150.925 63.140 150.955 ;
        RECT 62.400 150.625 63.315 150.925 ;
        RECT 62.990 150.450 63.315 150.625 ;
        RECT 62.020 149.895 62.275 150.425 ;
        RECT 62.445 149.715 62.750 150.175 ;
        RECT 62.995 150.095 63.315 150.450 ;
        RECT 63.485 150.665 64.025 151.035 ;
        RECT 64.360 150.945 64.765 151.115 ;
        RECT 63.485 150.265 63.725 150.665 ;
        RECT 64.205 150.495 64.425 150.775 ;
        RECT 63.895 150.325 64.425 150.495 ;
        RECT 63.895 150.095 64.065 150.325 ;
        RECT 64.595 150.165 64.765 150.945 ;
        RECT 64.935 150.335 65.285 150.955 ;
        RECT 65.455 150.335 65.665 151.125 ;
        RECT 65.855 151.155 67.355 151.325 ;
        RECT 65.855 150.465 66.025 151.155 ;
        RECT 67.715 150.985 67.885 151.765 ;
        RECT 68.690 151.635 68.860 151.765 ;
        RECT 66.195 150.815 67.885 150.985 ;
        RECT 68.055 151.205 68.520 151.595 ;
        RECT 68.690 151.465 69.085 151.635 ;
        RECT 66.195 150.635 66.365 150.815 ;
        RECT 62.995 149.925 64.065 150.095 ;
        RECT 64.235 149.715 64.425 150.155 ;
        RECT 64.595 149.885 65.545 150.165 ;
        RECT 65.855 150.075 66.115 150.465 ;
        RECT 66.535 150.395 67.325 150.645 ;
        RECT 65.765 149.905 66.115 150.075 ;
        RECT 66.325 149.715 66.655 150.175 ;
        RECT 67.530 150.105 67.700 150.815 ;
        RECT 68.055 150.615 68.225 151.205 ;
        RECT 67.870 150.395 68.225 150.615 ;
        RECT 68.395 150.395 68.745 151.015 ;
        RECT 68.915 150.105 69.085 151.465 ;
        RECT 69.450 151.295 69.775 152.080 ;
        RECT 69.255 150.245 69.715 151.295 ;
        RECT 67.530 149.935 68.385 150.105 ;
        RECT 68.590 149.935 69.085 150.105 ;
        RECT 69.255 149.715 69.585 150.075 ;
        RECT 69.945 149.975 70.115 152.095 ;
        RECT 70.285 151.765 70.615 152.265 ;
        RECT 70.785 151.595 71.040 152.095 ;
        RECT 70.290 151.425 71.040 151.595 ;
        RECT 70.290 150.435 70.520 151.425 ;
        RECT 70.690 150.605 71.040 151.255 ;
        RECT 71.215 151.125 71.485 152.095 ;
        RECT 71.695 151.465 71.975 152.265 ;
        RECT 72.145 151.755 73.800 152.045 ;
        RECT 72.210 151.415 73.800 151.585 ;
        RECT 72.210 151.295 72.380 151.415 ;
        RECT 71.655 151.125 72.380 151.295 ;
        RECT 70.290 150.265 71.040 150.435 ;
        RECT 70.285 149.715 70.615 150.095 ;
        RECT 70.785 149.975 71.040 150.265 ;
        RECT 71.215 150.390 71.385 151.125 ;
        RECT 71.655 150.955 71.825 151.125 ;
        RECT 72.570 151.075 73.285 151.245 ;
        RECT 73.480 151.125 73.800 151.415 ;
        RECT 73.975 151.125 74.315 152.095 ;
        RECT 74.485 151.125 74.655 152.265 ;
        RECT 74.925 151.465 75.175 152.265 ;
        RECT 75.820 151.295 76.150 152.095 ;
        RECT 76.450 151.465 76.780 152.265 ;
        RECT 76.950 151.295 77.280 152.095 ;
        RECT 74.845 151.125 77.280 151.295 ;
        RECT 78.115 151.505 78.630 151.915 ;
        RECT 78.865 151.505 79.035 152.265 ;
        RECT 79.205 151.925 81.235 152.095 ;
        RECT 71.555 150.625 71.825 150.955 ;
        RECT 71.995 150.625 72.400 150.955 ;
        RECT 72.570 150.625 73.280 151.075 ;
        RECT 71.655 150.455 71.825 150.625 ;
        RECT 71.215 150.045 71.485 150.390 ;
        RECT 71.655 150.285 73.265 150.455 ;
        RECT 73.450 150.385 73.800 150.955 ;
        RECT 73.975 150.565 74.150 151.125 ;
        RECT 74.845 150.875 75.015 151.125 ;
        RECT 74.320 150.705 75.015 150.875 ;
        RECT 75.190 150.705 75.610 150.905 ;
        RECT 75.780 150.705 76.110 150.905 ;
        RECT 76.280 150.705 76.610 150.905 ;
        RECT 73.975 150.515 74.205 150.565 ;
        RECT 71.675 149.715 72.055 150.115 ;
        RECT 72.225 149.935 72.395 150.285 ;
        RECT 72.565 149.715 72.895 150.115 ;
        RECT 73.095 149.935 73.265 150.285 ;
        RECT 73.465 149.715 73.795 150.215 ;
        RECT 73.975 149.885 74.315 150.515 ;
        RECT 74.485 149.715 74.735 150.515 ;
        RECT 74.925 150.365 76.150 150.535 ;
        RECT 74.925 149.885 75.255 150.365 ;
        RECT 75.425 149.715 75.650 150.175 ;
        RECT 75.820 149.885 76.150 150.365 ;
        RECT 76.780 150.495 76.950 151.125 ;
        RECT 77.135 150.705 77.485 150.955 ;
        RECT 78.115 150.695 78.455 151.505 ;
        RECT 79.205 151.260 79.375 151.925 ;
        RECT 79.770 151.585 80.895 151.755 ;
        RECT 78.625 151.070 79.375 151.260 ;
        RECT 79.545 151.245 80.555 151.415 ;
        RECT 78.115 150.525 79.345 150.695 ;
        RECT 76.780 149.885 77.280 150.495 ;
        RECT 78.390 149.920 78.635 150.525 ;
        RECT 78.855 149.715 79.365 150.250 ;
        RECT 79.545 149.885 79.735 151.245 ;
        RECT 79.905 150.225 80.180 151.045 ;
        RECT 80.385 150.445 80.555 151.245 ;
        RECT 80.725 150.455 80.895 151.585 ;
        RECT 81.065 150.955 81.235 151.925 ;
        RECT 81.405 151.125 81.575 152.265 ;
        RECT 81.745 151.125 82.080 152.095 ;
        RECT 81.065 150.625 81.260 150.955 ;
        RECT 81.485 150.625 81.740 150.955 ;
        RECT 81.485 150.455 81.655 150.625 ;
        RECT 81.910 150.455 82.080 151.125 ;
        RECT 80.725 150.285 81.655 150.455 ;
        RECT 80.725 150.250 80.900 150.285 ;
        RECT 79.905 150.055 80.185 150.225 ;
        RECT 79.905 149.885 80.180 150.055 ;
        RECT 80.370 149.885 80.900 150.250 ;
        RECT 81.325 149.715 81.655 150.115 ;
        RECT 81.825 149.885 82.080 150.455 ;
        RECT 82.260 151.125 82.595 152.095 ;
        RECT 82.765 151.125 82.935 152.265 ;
        RECT 83.105 151.925 85.135 152.095 ;
        RECT 82.260 150.455 82.430 151.125 ;
        RECT 83.105 150.955 83.275 151.925 ;
        RECT 82.600 150.625 82.855 150.955 ;
        RECT 83.080 150.625 83.275 150.955 ;
        RECT 83.445 151.585 84.570 151.755 ;
        RECT 82.685 150.455 82.855 150.625 ;
        RECT 83.445 150.455 83.615 151.585 ;
        RECT 82.260 149.885 82.515 150.455 ;
        RECT 82.685 150.285 83.615 150.455 ;
        RECT 83.785 151.245 84.795 151.415 ;
        RECT 83.785 150.445 83.955 151.245 ;
        RECT 84.160 150.905 84.435 151.045 ;
        RECT 84.155 150.735 84.435 150.905 ;
        RECT 83.440 150.250 83.615 150.285 ;
        RECT 82.685 149.715 83.015 150.115 ;
        RECT 83.440 149.885 83.970 150.250 ;
        RECT 84.160 149.885 84.435 150.735 ;
        RECT 84.605 149.885 84.795 151.245 ;
        RECT 84.965 151.260 85.135 151.925 ;
        RECT 85.305 151.505 85.475 152.265 ;
        RECT 85.710 151.505 86.225 151.915 ;
        RECT 84.965 151.070 85.715 151.260 ;
        RECT 85.885 150.695 86.225 151.505 ;
        RECT 87.315 151.100 87.605 152.265 ;
        RECT 88.240 151.830 93.585 152.265 ;
        RECT 84.995 150.525 86.225 150.695 ;
        RECT 89.830 150.580 90.180 151.830 ;
        RECT 93.960 151.295 94.290 152.095 ;
        RECT 94.460 151.465 94.790 152.265 ;
        RECT 95.090 151.295 95.420 152.095 ;
        RECT 96.065 151.465 96.315 152.265 ;
        RECT 93.960 151.125 96.395 151.295 ;
        RECT 96.585 151.125 96.755 152.265 ;
        RECT 96.925 151.125 97.265 152.095 ;
        RECT 84.975 149.715 85.485 150.250 ;
        RECT 85.705 149.920 85.950 150.525 ;
        RECT 87.315 149.715 87.605 150.440 ;
        RECT 91.660 150.260 92.000 151.090 ;
        RECT 93.755 150.705 94.105 150.955 ;
        RECT 94.290 150.495 94.460 151.125 ;
        RECT 94.630 150.705 94.960 150.905 ;
        RECT 95.130 150.705 95.460 150.905 ;
        RECT 95.630 150.705 96.050 150.905 ;
        RECT 96.225 150.875 96.395 151.125 ;
        RECT 96.225 150.705 96.920 150.875 ;
        RECT 88.240 149.715 93.585 150.260 ;
        RECT 93.960 149.885 94.460 150.495 ;
        RECT 95.090 150.365 96.315 150.535 ;
        RECT 97.090 150.515 97.265 151.125 ;
        RECT 95.090 149.885 95.420 150.365 ;
        RECT 95.590 149.715 95.815 150.175 ;
        RECT 95.985 149.885 96.315 150.365 ;
        RECT 96.505 149.715 96.755 150.515 ;
        RECT 96.925 149.885 97.265 150.515 ;
        RECT 97.435 151.125 97.775 152.095 ;
        RECT 97.945 151.125 98.115 152.265 ;
        RECT 98.385 151.465 98.635 152.265 ;
        RECT 99.280 151.295 99.610 152.095 ;
        RECT 99.910 151.465 100.240 152.265 ;
        RECT 100.410 151.295 100.740 152.095 ;
        RECT 98.305 151.125 100.740 151.295 ;
        RECT 101.615 151.125 101.845 152.265 ;
        RECT 97.435 151.075 97.665 151.125 ;
        RECT 97.435 150.515 97.610 151.075 ;
        RECT 98.305 150.875 98.475 151.125 ;
        RECT 97.780 150.705 98.475 150.875 ;
        RECT 98.650 150.705 99.070 150.905 ;
        RECT 99.240 150.705 99.570 150.905 ;
        RECT 99.740 150.705 100.070 150.905 ;
        RECT 97.435 149.885 97.775 150.515 ;
        RECT 97.945 149.715 98.195 150.515 ;
        RECT 98.385 150.365 99.610 150.535 ;
        RECT 98.385 149.885 98.715 150.365 ;
        RECT 98.885 149.715 99.110 150.175 ;
        RECT 99.280 149.885 99.610 150.365 ;
        RECT 100.240 150.495 100.410 151.125 ;
        RECT 102.015 151.115 102.345 152.095 ;
        RECT 102.515 151.125 102.725 152.265 ;
        RECT 102.955 151.505 103.470 151.915 ;
        RECT 103.705 151.505 103.875 152.265 ;
        RECT 104.045 151.925 106.075 152.095 ;
        RECT 100.595 150.705 100.945 150.955 ;
        RECT 101.595 150.705 101.925 150.955 ;
        RECT 100.240 149.885 100.740 150.495 ;
        RECT 101.615 149.715 101.845 150.535 ;
        RECT 102.095 150.515 102.345 151.115 ;
        RECT 102.955 150.695 103.295 151.505 ;
        RECT 104.045 151.260 104.215 151.925 ;
        RECT 104.610 151.585 105.735 151.755 ;
        RECT 103.465 151.070 104.215 151.260 ;
        RECT 104.385 151.245 105.395 151.415 ;
        RECT 102.015 149.885 102.345 150.515 ;
        RECT 102.515 149.715 102.725 150.535 ;
        RECT 102.955 150.525 104.185 150.695 ;
        RECT 103.230 149.920 103.475 150.525 ;
        RECT 103.695 149.715 104.205 150.250 ;
        RECT 104.385 149.885 104.575 151.245 ;
        RECT 104.745 150.905 105.020 151.045 ;
        RECT 104.745 150.735 105.025 150.905 ;
        RECT 104.745 149.885 105.020 150.735 ;
        RECT 105.225 150.445 105.395 151.245 ;
        RECT 105.565 150.455 105.735 151.585 ;
        RECT 105.905 150.955 106.075 151.925 ;
        RECT 106.245 151.125 106.415 152.265 ;
        RECT 106.585 151.125 106.920 152.095 ;
        RECT 108.105 151.335 108.275 152.095 ;
        RECT 108.455 151.505 108.785 152.265 ;
        RECT 108.105 151.165 108.770 151.335 ;
        RECT 108.955 151.190 109.225 152.095 ;
        RECT 105.905 150.625 106.100 150.955 ;
        RECT 106.325 150.625 106.580 150.955 ;
        RECT 106.325 150.455 106.495 150.625 ;
        RECT 106.750 150.455 106.920 151.125 ;
        RECT 108.600 151.020 108.770 151.165 ;
        RECT 108.035 150.615 108.365 150.985 ;
        RECT 108.600 150.690 108.885 151.020 ;
        RECT 105.565 150.285 106.495 150.455 ;
        RECT 105.565 150.250 105.740 150.285 ;
        RECT 105.210 149.885 105.740 150.250 ;
        RECT 106.165 149.715 106.495 150.115 ;
        RECT 106.665 149.885 106.920 150.455 ;
        RECT 108.600 150.435 108.770 150.690 ;
        RECT 108.105 150.265 108.770 150.435 ;
        RECT 109.055 150.390 109.225 151.190 ;
        RECT 109.395 151.175 111.985 152.265 ;
        RECT 112.155 151.175 113.365 152.265 ;
        RECT 109.395 150.655 110.605 151.175 ;
        RECT 110.775 150.485 111.985 151.005 ;
        RECT 112.155 150.635 112.675 151.175 ;
        RECT 108.105 149.885 108.275 150.265 ;
        RECT 108.455 149.715 108.785 150.095 ;
        RECT 108.965 149.885 109.225 150.390 ;
        RECT 109.395 149.715 111.985 150.485 ;
        RECT 112.845 150.465 113.365 151.005 ;
        RECT 112.155 149.715 113.365 150.465 ;
        RECT 22.830 149.545 113.450 149.715 ;
        RECT 22.915 148.795 24.125 149.545 ;
        RECT 24.670 148.835 24.925 149.365 ;
        RECT 25.105 149.085 25.390 149.545 ;
        RECT 22.915 148.255 23.435 148.795 ;
        RECT 23.605 148.085 24.125 148.625 ;
        RECT 22.915 146.995 24.125 148.085 ;
        RECT 24.670 147.975 24.850 148.835 ;
        RECT 25.570 148.635 25.820 149.285 ;
        RECT 25.020 148.305 25.820 148.635 ;
        RECT 24.670 147.505 24.925 147.975 ;
        RECT 24.585 147.335 24.925 147.505 ;
        RECT 24.670 147.305 24.925 147.335 ;
        RECT 25.105 146.995 25.390 147.795 ;
        RECT 25.570 147.715 25.820 148.305 ;
        RECT 26.020 148.950 26.340 149.280 ;
        RECT 26.520 149.065 27.180 149.545 ;
        RECT 27.380 149.155 28.230 149.325 ;
        RECT 26.020 148.055 26.210 148.950 ;
        RECT 26.530 148.625 27.190 148.895 ;
        RECT 26.860 148.565 27.190 148.625 ;
        RECT 26.380 148.395 26.710 148.455 ;
        RECT 27.380 148.395 27.550 149.155 ;
        RECT 28.790 149.085 29.110 149.545 ;
        RECT 29.310 148.905 29.560 149.335 ;
        RECT 29.850 149.105 30.260 149.545 ;
        RECT 30.430 149.165 31.445 149.365 ;
        RECT 27.720 148.735 28.970 148.905 ;
        RECT 27.720 148.615 28.050 148.735 ;
        RECT 26.380 148.225 28.280 148.395 ;
        RECT 26.020 147.885 27.940 148.055 ;
        RECT 26.020 147.865 26.340 147.885 ;
        RECT 25.570 147.205 25.900 147.715 ;
        RECT 26.170 147.255 26.340 147.865 ;
        RECT 28.110 147.715 28.280 148.225 ;
        RECT 28.450 148.155 28.630 148.565 ;
        RECT 28.800 147.975 28.970 148.735 ;
        RECT 26.510 146.995 26.840 147.685 ;
        RECT 27.070 147.545 28.280 147.715 ;
        RECT 28.450 147.665 28.970 147.975 ;
        RECT 29.140 148.565 29.560 148.905 ;
        RECT 29.850 148.565 30.260 148.895 ;
        RECT 29.140 147.795 29.330 148.565 ;
        RECT 30.430 148.435 30.600 149.165 ;
        RECT 31.745 148.995 31.915 149.325 ;
        RECT 32.085 149.165 32.415 149.545 ;
        RECT 30.770 148.615 31.120 148.985 ;
        RECT 30.430 148.395 30.850 148.435 ;
        RECT 29.500 148.225 30.850 148.395 ;
        RECT 29.500 148.065 29.750 148.225 ;
        RECT 30.260 147.795 30.510 148.055 ;
        RECT 29.140 147.545 30.510 147.795 ;
        RECT 27.070 147.255 27.310 147.545 ;
        RECT 28.110 147.465 28.280 147.545 ;
        RECT 27.510 146.995 27.930 147.375 ;
        RECT 28.110 147.215 28.740 147.465 ;
        RECT 29.210 146.995 29.540 147.375 ;
        RECT 29.710 147.255 29.880 147.545 ;
        RECT 30.680 147.380 30.850 148.225 ;
        RECT 31.300 148.055 31.520 148.925 ;
        RECT 31.745 148.805 32.440 148.995 ;
        RECT 31.020 147.675 31.520 148.055 ;
        RECT 31.690 148.005 32.100 148.625 ;
        RECT 32.270 147.835 32.440 148.805 ;
        RECT 31.745 147.665 32.440 147.835 ;
        RECT 30.060 146.995 30.440 147.375 ;
        RECT 30.680 147.210 31.510 147.380 ;
        RECT 31.745 147.165 31.915 147.665 ;
        RECT 32.085 146.995 32.415 147.495 ;
        RECT 32.630 147.165 32.855 149.285 ;
        RECT 33.025 149.165 33.355 149.545 ;
        RECT 33.525 148.995 33.695 149.285 ;
        RECT 33.030 148.825 33.695 148.995 ;
        RECT 33.030 147.835 33.260 148.825 ;
        RECT 33.960 148.805 34.215 149.375 ;
        RECT 34.385 149.145 34.715 149.545 ;
        RECT 35.140 149.010 35.670 149.375 ;
        RECT 35.860 149.205 36.135 149.375 ;
        RECT 35.855 149.035 36.135 149.205 ;
        RECT 35.140 148.975 35.315 149.010 ;
        RECT 34.385 148.805 35.315 148.975 ;
        RECT 33.430 148.005 33.780 148.655 ;
        RECT 33.960 148.135 34.130 148.805 ;
        RECT 34.385 148.635 34.555 148.805 ;
        RECT 34.300 148.305 34.555 148.635 ;
        RECT 34.780 148.305 34.975 148.635 ;
        RECT 33.030 147.665 33.695 147.835 ;
        RECT 33.025 146.995 33.355 147.495 ;
        RECT 33.525 147.165 33.695 147.665 ;
        RECT 33.960 147.165 34.295 148.135 ;
        RECT 34.465 146.995 34.635 148.135 ;
        RECT 34.805 147.335 34.975 148.305 ;
        RECT 35.145 147.675 35.315 148.805 ;
        RECT 35.485 148.015 35.655 148.815 ;
        RECT 35.860 148.215 36.135 149.035 ;
        RECT 36.305 148.015 36.495 149.375 ;
        RECT 36.675 149.010 37.185 149.545 ;
        RECT 37.405 148.735 37.650 149.340 ;
        RECT 38.755 148.915 39.085 149.275 ;
        RECT 39.705 149.085 39.955 149.545 ;
        RECT 40.125 149.085 40.685 149.375 ;
        RECT 36.695 148.565 37.925 148.735 ;
        RECT 38.755 148.725 40.145 148.915 ;
        RECT 35.485 147.845 36.495 148.015 ;
        RECT 36.665 148.000 37.415 148.190 ;
        RECT 35.145 147.505 36.270 147.675 ;
        RECT 36.665 147.335 36.835 148.000 ;
        RECT 37.585 147.755 37.925 148.565 ;
        RECT 39.975 148.635 40.145 148.725 ;
        RECT 38.570 148.305 39.245 148.555 ;
        RECT 39.465 148.305 39.805 148.555 ;
        RECT 39.975 148.305 40.265 148.635 ;
        RECT 38.570 147.945 38.835 148.305 ;
        RECT 39.975 148.055 40.145 148.305 ;
        RECT 34.805 147.165 36.835 147.335 ;
        RECT 37.005 146.995 37.175 147.755 ;
        RECT 37.410 147.345 37.925 147.755 ;
        RECT 39.205 147.885 40.145 148.055 ;
        RECT 38.755 146.995 39.035 147.665 ;
        RECT 39.205 147.335 39.505 147.885 ;
        RECT 40.435 147.715 40.685 149.085 ;
        RECT 41.055 148.915 41.385 149.275 ;
        RECT 42.005 149.085 42.255 149.545 ;
        RECT 42.425 149.085 42.985 149.375 ;
        RECT 41.055 148.725 42.445 148.915 ;
        RECT 42.275 148.635 42.445 148.725 ;
        RECT 40.870 148.305 41.545 148.555 ;
        RECT 41.765 148.305 42.105 148.555 ;
        RECT 42.275 148.305 42.565 148.635 ;
        RECT 40.870 147.945 41.135 148.305 ;
        RECT 42.275 148.055 42.445 148.305 ;
        RECT 39.705 146.995 40.035 147.715 ;
        RECT 40.225 147.165 40.685 147.715 ;
        RECT 41.505 147.885 42.445 148.055 ;
        RECT 41.055 146.995 41.335 147.665 ;
        RECT 41.505 147.335 41.805 147.885 ;
        RECT 42.735 147.715 42.985 149.085 ;
        RECT 42.005 146.995 42.335 147.715 ;
        RECT 42.525 147.165 42.985 147.715 ;
        RECT 43.155 149.085 43.715 149.375 ;
        RECT 43.885 149.085 44.135 149.545 ;
        RECT 43.155 147.715 43.405 149.085 ;
        RECT 44.755 148.915 45.085 149.275 ;
        RECT 43.695 148.725 45.085 148.915 ;
        RECT 45.455 148.775 47.125 149.545 ;
        RECT 43.695 148.635 43.865 148.725 ;
        RECT 43.575 148.305 43.865 148.635 ;
        RECT 44.035 148.305 44.375 148.555 ;
        RECT 44.595 148.305 45.270 148.555 ;
        RECT 43.695 148.055 43.865 148.305 ;
        RECT 43.695 147.885 44.635 148.055 ;
        RECT 45.005 147.945 45.270 148.305 ;
        RECT 45.455 148.085 46.205 148.605 ;
        RECT 46.375 148.255 47.125 148.775 ;
        RECT 47.335 148.725 47.565 149.545 ;
        RECT 47.735 148.745 48.065 149.375 ;
        RECT 47.315 148.305 47.645 148.555 ;
        RECT 47.815 148.145 48.065 148.745 ;
        RECT 48.235 148.725 48.445 149.545 ;
        RECT 48.675 148.820 48.965 149.545 ;
        RECT 49.510 149.205 49.765 149.365 ;
        RECT 49.425 149.035 49.765 149.205 ;
        RECT 49.945 149.085 50.230 149.545 ;
        RECT 49.510 148.835 49.765 149.035 ;
        RECT 43.155 147.165 43.615 147.715 ;
        RECT 43.805 146.995 44.135 147.715 ;
        RECT 44.335 147.335 44.635 147.885 ;
        RECT 44.805 146.995 45.085 147.665 ;
        RECT 45.455 146.995 47.125 148.085 ;
        RECT 47.335 146.995 47.565 148.135 ;
        RECT 47.735 147.165 48.065 148.145 ;
        RECT 48.235 146.995 48.445 148.135 ;
        RECT 48.675 146.995 48.965 148.160 ;
        RECT 49.510 147.975 49.690 148.835 ;
        RECT 50.410 148.635 50.660 149.285 ;
        RECT 49.860 148.305 50.660 148.635 ;
        RECT 49.510 147.305 49.765 147.975 ;
        RECT 49.945 146.995 50.230 147.795 ;
        RECT 50.410 147.715 50.660 148.305 ;
        RECT 50.860 148.950 51.180 149.280 ;
        RECT 51.360 149.065 52.020 149.545 ;
        RECT 52.220 149.155 53.070 149.325 ;
        RECT 50.860 148.055 51.050 148.950 ;
        RECT 51.370 148.625 52.030 148.895 ;
        RECT 51.700 148.565 52.030 148.625 ;
        RECT 51.220 148.395 51.550 148.455 ;
        RECT 52.220 148.395 52.390 149.155 ;
        RECT 53.630 149.085 53.950 149.545 ;
        RECT 54.150 148.905 54.400 149.335 ;
        RECT 54.690 149.105 55.100 149.545 ;
        RECT 55.270 149.165 56.285 149.365 ;
        RECT 52.560 148.735 53.810 148.905 ;
        RECT 52.560 148.615 52.890 148.735 ;
        RECT 51.220 148.225 53.120 148.395 ;
        RECT 50.860 147.885 52.780 148.055 ;
        RECT 50.860 147.865 51.180 147.885 ;
        RECT 50.410 147.205 50.740 147.715 ;
        RECT 51.010 147.255 51.180 147.865 ;
        RECT 52.950 147.715 53.120 148.225 ;
        RECT 53.290 148.155 53.470 148.565 ;
        RECT 53.640 147.975 53.810 148.735 ;
        RECT 51.350 146.995 51.680 147.685 ;
        RECT 51.910 147.545 53.120 147.715 ;
        RECT 53.290 147.665 53.810 147.975 ;
        RECT 53.980 148.565 54.400 148.905 ;
        RECT 54.690 148.565 55.100 148.895 ;
        RECT 53.980 147.795 54.170 148.565 ;
        RECT 55.270 148.435 55.440 149.165 ;
        RECT 56.585 148.995 56.755 149.325 ;
        RECT 56.925 149.165 57.255 149.545 ;
        RECT 55.610 148.615 55.960 148.985 ;
        RECT 55.270 148.395 55.690 148.435 ;
        RECT 54.340 148.225 55.690 148.395 ;
        RECT 54.340 148.065 54.590 148.225 ;
        RECT 55.100 147.795 55.350 148.055 ;
        RECT 53.980 147.545 55.350 147.795 ;
        RECT 51.910 147.255 52.150 147.545 ;
        RECT 52.950 147.465 53.120 147.545 ;
        RECT 52.350 146.995 52.770 147.375 ;
        RECT 52.950 147.215 53.580 147.465 ;
        RECT 54.050 146.995 54.380 147.375 ;
        RECT 54.550 147.255 54.720 147.545 ;
        RECT 55.520 147.380 55.690 148.225 ;
        RECT 56.140 148.055 56.360 148.925 ;
        RECT 56.585 148.805 57.280 148.995 ;
        RECT 55.860 147.675 56.360 148.055 ;
        RECT 56.530 148.005 56.940 148.625 ;
        RECT 57.110 147.835 57.280 148.805 ;
        RECT 56.585 147.665 57.280 147.835 ;
        RECT 54.900 146.995 55.280 147.375 ;
        RECT 55.520 147.210 56.350 147.380 ;
        RECT 56.585 147.165 56.755 147.665 ;
        RECT 56.925 146.995 57.255 147.495 ;
        RECT 57.470 147.165 57.695 149.285 ;
        RECT 57.865 149.165 58.195 149.545 ;
        RECT 58.365 148.995 58.535 149.285 ;
        RECT 57.870 148.825 58.535 148.995 ;
        RECT 57.870 147.835 58.100 148.825 ;
        RECT 58.795 148.775 60.465 149.545 ;
        RECT 58.270 148.005 58.620 148.655 ;
        RECT 58.795 148.085 59.545 148.605 ;
        RECT 59.715 148.255 60.465 148.775 ;
        RECT 60.675 148.725 60.905 149.545 ;
        RECT 61.075 148.745 61.405 149.375 ;
        RECT 60.655 148.305 60.985 148.555 ;
        RECT 61.155 148.145 61.405 148.745 ;
        RECT 61.575 148.725 61.785 149.545 ;
        RECT 62.290 148.735 62.535 149.340 ;
        RECT 62.755 149.010 63.265 149.545 ;
        RECT 57.870 147.665 58.535 147.835 ;
        RECT 57.865 146.995 58.195 147.495 ;
        RECT 58.365 147.165 58.535 147.665 ;
        RECT 58.795 146.995 60.465 148.085 ;
        RECT 60.675 146.995 60.905 148.135 ;
        RECT 61.075 147.165 61.405 148.145 ;
        RECT 62.015 148.565 63.245 148.735 ;
        RECT 61.575 146.995 61.785 148.135 ;
        RECT 62.015 147.755 62.355 148.565 ;
        RECT 62.525 148.000 63.275 148.190 ;
        RECT 62.015 147.345 62.530 147.755 ;
        RECT 62.765 146.995 62.935 147.755 ;
        RECT 63.105 147.335 63.275 148.000 ;
        RECT 63.445 148.015 63.635 149.375 ;
        RECT 63.805 148.865 64.080 149.375 ;
        RECT 64.270 149.010 64.800 149.375 ;
        RECT 65.225 149.145 65.555 149.545 ;
        RECT 64.625 148.975 64.800 149.010 ;
        RECT 63.805 148.695 64.085 148.865 ;
        RECT 63.805 148.215 64.080 148.695 ;
        RECT 64.285 148.015 64.455 148.815 ;
        RECT 63.445 147.845 64.455 148.015 ;
        RECT 64.625 148.805 65.555 148.975 ;
        RECT 65.725 148.805 65.980 149.375 ;
        RECT 66.245 148.995 66.415 149.375 ;
        RECT 66.595 149.165 66.925 149.545 ;
        RECT 66.245 148.825 66.910 148.995 ;
        RECT 67.105 148.870 67.365 149.375 ;
        RECT 68.005 149.045 68.335 149.545 ;
        RECT 68.535 148.975 68.705 149.325 ;
        RECT 68.905 149.145 69.235 149.545 ;
        RECT 69.405 148.975 69.575 149.325 ;
        RECT 69.745 149.145 70.125 149.545 ;
        RECT 64.625 147.675 64.795 148.805 ;
        RECT 65.385 148.635 65.555 148.805 ;
        RECT 63.670 147.505 64.795 147.675 ;
        RECT 64.965 148.305 65.160 148.635 ;
        RECT 65.385 148.305 65.640 148.635 ;
        RECT 64.965 147.335 65.135 148.305 ;
        RECT 65.810 148.135 65.980 148.805 ;
        RECT 66.175 148.275 66.505 148.645 ;
        RECT 66.740 148.570 66.910 148.825 ;
        RECT 63.105 147.165 65.135 147.335 ;
        RECT 65.305 146.995 65.475 148.135 ;
        RECT 65.645 147.165 65.980 148.135 ;
        RECT 66.740 148.240 67.025 148.570 ;
        RECT 66.740 148.095 66.910 148.240 ;
        RECT 66.245 147.925 66.910 148.095 ;
        RECT 67.195 148.070 67.365 148.870 ;
        RECT 68.000 148.305 68.350 148.875 ;
        RECT 68.535 148.805 70.145 148.975 ;
        RECT 70.315 148.870 70.585 149.215 ;
        RECT 69.975 148.635 70.145 148.805 ;
        RECT 66.245 147.165 66.415 147.925 ;
        RECT 66.595 146.995 66.925 147.755 ;
        RECT 67.095 147.165 67.365 148.070 ;
        RECT 68.000 147.845 68.320 148.135 ;
        RECT 68.520 148.015 69.230 148.635 ;
        RECT 69.400 148.305 69.805 148.635 ;
        RECT 69.975 148.305 70.245 148.635 ;
        RECT 69.975 148.135 70.145 148.305 ;
        RECT 70.415 148.135 70.585 148.870 ;
        RECT 69.420 147.965 70.145 148.135 ;
        RECT 69.420 147.845 69.590 147.965 ;
        RECT 68.000 147.675 69.590 147.845 ;
        RECT 68.000 147.215 69.655 147.505 ;
        RECT 69.825 146.995 70.105 147.795 ;
        RECT 70.315 147.165 70.585 148.135 ;
        RECT 70.755 148.745 71.095 149.375 ;
        RECT 71.265 148.745 71.515 149.545 ;
        RECT 71.705 148.895 72.035 149.375 ;
        RECT 72.205 149.085 72.430 149.545 ;
        RECT 72.600 148.895 72.930 149.375 ;
        RECT 70.755 148.695 70.985 148.745 ;
        RECT 71.705 148.725 72.930 148.895 ;
        RECT 73.560 148.765 74.060 149.375 ;
        RECT 74.435 148.820 74.725 149.545 ;
        RECT 70.755 148.135 70.930 148.695 ;
        RECT 71.100 148.385 71.795 148.555 ;
        RECT 71.625 148.135 71.795 148.385 ;
        RECT 71.970 148.355 72.390 148.555 ;
        RECT 72.560 148.355 72.890 148.555 ;
        RECT 73.060 148.355 73.390 148.555 ;
        RECT 73.560 148.135 73.730 148.765 ;
        RECT 75.875 148.725 76.085 149.545 ;
        RECT 76.255 148.745 76.585 149.375 ;
        RECT 73.915 148.305 74.265 148.555 ;
        RECT 70.755 147.165 71.095 148.135 ;
        RECT 71.265 146.995 71.435 148.135 ;
        RECT 71.625 147.965 74.060 148.135 ;
        RECT 71.705 146.995 71.955 147.795 ;
        RECT 72.600 147.165 72.930 147.965 ;
        RECT 73.230 146.995 73.560 147.795 ;
        RECT 73.730 147.165 74.060 147.965 ;
        RECT 74.435 146.995 74.725 148.160 ;
        RECT 76.255 148.145 76.505 148.745 ;
        RECT 76.755 148.725 76.985 149.545 ;
        RECT 77.570 148.835 77.825 149.365 ;
        RECT 78.005 149.085 78.290 149.545 ;
        RECT 76.675 148.305 77.005 148.555 ;
        RECT 77.570 148.185 77.750 148.835 ;
        RECT 78.470 148.635 78.720 149.285 ;
        RECT 77.920 148.305 78.720 148.635 ;
        RECT 75.875 146.995 76.085 148.135 ;
        RECT 76.255 147.165 76.585 148.145 ;
        RECT 76.755 146.995 76.985 148.135 ;
        RECT 77.485 148.015 77.750 148.185 ;
        RECT 77.570 147.975 77.750 148.015 ;
        RECT 77.570 147.305 77.825 147.975 ;
        RECT 78.005 146.995 78.290 147.795 ;
        RECT 78.470 147.715 78.720 148.305 ;
        RECT 78.920 148.950 79.240 149.280 ;
        RECT 79.420 149.065 80.080 149.545 ;
        RECT 80.280 149.155 81.130 149.325 ;
        RECT 78.920 148.055 79.110 148.950 ;
        RECT 79.430 148.625 80.090 148.895 ;
        RECT 79.760 148.565 80.090 148.625 ;
        RECT 79.280 148.395 79.610 148.455 ;
        RECT 80.280 148.395 80.450 149.155 ;
        RECT 81.690 149.085 82.010 149.545 ;
        RECT 82.210 148.905 82.460 149.335 ;
        RECT 82.750 149.105 83.160 149.545 ;
        RECT 83.330 149.165 84.345 149.365 ;
        RECT 80.620 148.735 81.870 148.905 ;
        RECT 80.620 148.615 80.950 148.735 ;
        RECT 79.280 148.225 81.180 148.395 ;
        RECT 78.920 147.885 80.840 148.055 ;
        RECT 78.920 147.865 79.240 147.885 ;
        RECT 78.470 147.205 78.800 147.715 ;
        RECT 79.070 147.255 79.240 147.865 ;
        RECT 81.010 147.715 81.180 148.225 ;
        RECT 81.350 148.155 81.530 148.565 ;
        RECT 81.700 147.975 81.870 148.735 ;
        RECT 79.410 146.995 79.740 147.685 ;
        RECT 79.970 147.545 81.180 147.715 ;
        RECT 81.350 147.665 81.870 147.975 ;
        RECT 82.040 148.565 82.460 148.905 ;
        RECT 82.750 148.565 83.160 148.895 ;
        RECT 82.040 147.795 82.230 148.565 ;
        RECT 83.330 148.435 83.500 149.165 ;
        RECT 84.645 148.995 84.815 149.325 ;
        RECT 84.985 149.165 85.315 149.545 ;
        RECT 83.670 148.615 84.020 148.985 ;
        RECT 83.330 148.395 83.750 148.435 ;
        RECT 82.400 148.225 83.750 148.395 ;
        RECT 82.400 148.065 82.650 148.225 ;
        RECT 83.160 147.795 83.410 148.055 ;
        RECT 82.040 147.545 83.410 147.795 ;
        RECT 79.970 147.255 80.210 147.545 ;
        RECT 81.010 147.465 81.180 147.545 ;
        RECT 80.410 146.995 80.830 147.375 ;
        RECT 81.010 147.215 81.640 147.465 ;
        RECT 82.110 146.995 82.440 147.375 ;
        RECT 82.610 147.255 82.780 147.545 ;
        RECT 83.580 147.380 83.750 148.225 ;
        RECT 84.200 148.055 84.420 148.925 ;
        RECT 84.645 148.805 85.340 148.995 ;
        RECT 83.920 147.675 84.420 148.055 ;
        RECT 84.590 148.005 85.000 148.625 ;
        RECT 85.170 147.835 85.340 148.805 ;
        RECT 84.645 147.665 85.340 147.835 ;
        RECT 82.960 146.995 83.340 147.375 ;
        RECT 83.580 147.210 84.410 147.380 ;
        RECT 84.645 147.165 84.815 147.665 ;
        RECT 84.985 146.995 85.315 147.495 ;
        RECT 85.530 147.165 85.755 149.285 ;
        RECT 85.925 149.165 86.255 149.545 ;
        RECT 86.425 148.995 86.595 149.285 ;
        RECT 85.930 148.825 86.595 148.995 ;
        RECT 86.855 148.870 87.115 149.375 ;
        RECT 87.295 149.165 87.625 149.545 ;
        RECT 87.805 148.995 87.975 149.375 ;
        RECT 89.165 149.045 89.495 149.545 ;
        RECT 85.930 147.835 86.160 148.825 ;
        RECT 86.330 148.005 86.680 148.655 ;
        RECT 86.855 148.070 87.025 148.870 ;
        RECT 87.310 148.825 87.975 148.995 ;
        RECT 89.695 148.975 89.865 149.325 ;
        RECT 90.065 149.145 90.395 149.545 ;
        RECT 90.565 148.975 90.735 149.325 ;
        RECT 90.905 149.145 91.285 149.545 ;
        RECT 87.310 148.570 87.480 148.825 ;
        RECT 87.195 148.240 87.480 148.570 ;
        RECT 87.715 148.275 88.045 148.645 ;
        RECT 89.160 148.305 89.510 148.875 ;
        RECT 89.695 148.805 91.305 148.975 ;
        RECT 91.475 148.870 91.745 149.215 ;
        RECT 91.135 148.635 91.305 148.805 ;
        RECT 87.310 148.095 87.480 148.240 ;
        RECT 85.930 147.665 86.595 147.835 ;
        RECT 85.925 146.995 86.255 147.495 ;
        RECT 86.425 147.165 86.595 147.665 ;
        RECT 86.855 147.165 87.125 148.070 ;
        RECT 87.310 147.925 87.975 148.095 ;
        RECT 87.295 146.995 87.625 147.755 ;
        RECT 87.805 147.165 87.975 147.925 ;
        RECT 89.160 147.845 89.480 148.135 ;
        RECT 89.680 148.015 90.390 148.635 ;
        RECT 90.560 148.305 90.965 148.635 ;
        RECT 91.135 148.305 91.405 148.635 ;
        RECT 91.135 148.135 91.305 148.305 ;
        RECT 91.575 148.135 91.745 148.870 ;
        RECT 90.580 147.965 91.305 148.135 ;
        RECT 90.580 147.845 90.750 147.965 ;
        RECT 89.160 147.675 90.750 147.845 ;
        RECT 89.160 147.215 90.815 147.505 ;
        RECT 90.985 146.995 91.265 147.795 ;
        RECT 91.475 147.165 91.745 148.135 ;
        RECT 91.915 148.745 92.255 149.375 ;
        RECT 92.425 148.745 92.675 149.545 ;
        RECT 92.865 148.895 93.195 149.375 ;
        RECT 93.365 149.085 93.590 149.545 ;
        RECT 93.760 148.895 94.090 149.375 ;
        RECT 91.915 148.695 92.145 148.745 ;
        RECT 92.865 148.725 94.090 148.895 ;
        RECT 94.720 148.765 95.220 149.375 ;
        RECT 95.605 149.045 95.935 149.545 ;
        RECT 96.135 148.975 96.305 149.325 ;
        RECT 96.505 149.145 96.835 149.545 ;
        RECT 97.005 148.975 97.175 149.325 ;
        RECT 97.345 149.145 97.725 149.545 ;
        RECT 91.915 148.135 92.090 148.695 ;
        RECT 92.260 148.385 92.955 148.555 ;
        RECT 92.785 148.135 92.955 148.385 ;
        RECT 93.130 148.355 93.550 148.555 ;
        RECT 93.720 148.355 94.050 148.555 ;
        RECT 94.220 148.355 94.550 148.555 ;
        RECT 94.720 148.135 94.890 148.765 ;
        RECT 95.075 148.305 95.425 148.555 ;
        RECT 95.600 148.305 95.950 148.875 ;
        RECT 96.135 148.805 97.745 148.975 ;
        RECT 97.915 148.870 98.185 149.215 ;
        RECT 97.575 148.635 97.745 148.805 ;
        RECT 91.915 147.165 92.255 148.135 ;
        RECT 92.425 146.995 92.595 148.135 ;
        RECT 92.785 147.965 95.220 148.135 ;
        RECT 92.865 146.995 93.115 147.795 ;
        RECT 93.760 147.165 94.090 147.965 ;
        RECT 94.390 146.995 94.720 147.795 ;
        RECT 94.890 147.165 95.220 147.965 ;
        RECT 95.600 147.845 95.920 148.135 ;
        RECT 96.120 148.015 96.830 148.635 ;
        RECT 97.000 148.305 97.405 148.635 ;
        RECT 97.575 148.305 97.845 148.635 ;
        RECT 97.575 148.135 97.745 148.305 ;
        RECT 98.015 148.135 98.185 148.870 ;
        RECT 98.355 148.775 100.025 149.545 ;
        RECT 100.195 148.820 100.485 149.545 ;
        RECT 100.655 148.775 102.325 149.545 ;
        RECT 97.020 147.965 97.745 148.135 ;
        RECT 97.020 147.845 97.190 147.965 ;
        RECT 95.600 147.675 97.190 147.845 ;
        RECT 95.600 147.215 97.255 147.505 ;
        RECT 97.425 146.995 97.705 147.795 ;
        RECT 97.915 147.165 98.185 148.135 ;
        RECT 98.355 148.085 99.105 148.605 ;
        RECT 99.275 148.255 100.025 148.775 ;
        RECT 98.355 146.995 100.025 148.085 ;
        RECT 100.195 146.995 100.485 148.160 ;
        RECT 100.655 148.085 101.405 148.605 ;
        RECT 101.575 148.255 102.325 148.775 ;
        RECT 102.870 148.835 103.125 149.365 ;
        RECT 103.305 149.085 103.590 149.545 ;
        RECT 100.655 146.995 102.325 148.085 ;
        RECT 102.870 147.975 103.050 148.835 ;
        RECT 103.770 148.635 104.020 149.285 ;
        RECT 103.220 148.305 104.020 148.635 ;
        RECT 102.870 147.505 103.125 147.975 ;
        RECT 102.785 147.335 103.125 147.505 ;
        RECT 102.870 147.305 103.125 147.335 ;
        RECT 103.305 146.995 103.590 147.795 ;
        RECT 103.770 147.715 104.020 148.305 ;
        RECT 104.220 148.950 104.540 149.280 ;
        RECT 104.720 149.065 105.380 149.545 ;
        RECT 105.580 149.155 106.430 149.325 ;
        RECT 104.220 148.055 104.410 148.950 ;
        RECT 104.730 148.625 105.390 148.895 ;
        RECT 105.060 148.565 105.390 148.625 ;
        RECT 104.580 148.395 104.910 148.455 ;
        RECT 105.580 148.395 105.750 149.155 ;
        RECT 106.990 149.085 107.310 149.545 ;
        RECT 107.510 148.905 107.760 149.335 ;
        RECT 108.050 149.105 108.460 149.545 ;
        RECT 108.630 149.165 109.645 149.365 ;
        RECT 105.920 148.735 107.170 148.905 ;
        RECT 105.920 148.615 106.250 148.735 ;
        RECT 104.580 148.225 106.480 148.395 ;
        RECT 104.220 147.885 106.140 148.055 ;
        RECT 104.220 147.865 104.540 147.885 ;
        RECT 103.770 147.205 104.100 147.715 ;
        RECT 104.370 147.255 104.540 147.865 ;
        RECT 106.310 147.715 106.480 148.225 ;
        RECT 106.650 148.155 106.830 148.565 ;
        RECT 107.000 147.975 107.170 148.735 ;
        RECT 104.710 146.995 105.040 147.685 ;
        RECT 105.270 147.545 106.480 147.715 ;
        RECT 106.650 147.665 107.170 147.975 ;
        RECT 107.340 148.565 107.760 148.905 ;
        RECT 108.050 148.565 108.460 148.895 ;
        RECT 107.340 147.795 107.530 148.565 ;
        RECT 108.630 148.435 108.800 149.165 ;
        RECT 109.945 148.995 110.115 149.325 ;
        RECT 110.285 149.165 110.615 149.545 ;
        RECT 108.970 148.615 109.320 148.985 ;
        RECT 108.630 148.395 109.050 148.435 ;
        RECT 107.700 148.225 109.050 148.395 ;
        RECT 107.700 148.065 107.950 148.225 ;
        RECT 108.460 147.795 108.710 148.055 ;
        RECT 107.340 147.545 108.710 147.795 ;
        RECT 105.270 147.255 105.510 147.545 ;
        RECT 106.310 147.465 106.480 147.545 ;
        RECT 105.710 146.995 106.130 147.375 ;
        RECT 106.310 147.215 106.940 147.465 ;
        RECT 107.410 146.995 107.740 147.375 ;
        RECT 107.910 147.255 108.080 147.545 ;
        RECT 108.880 147.380 109.050 148.225 ;
        RECT 109.500 148.055 109.720 148.925 ;
        RECT 109.945 148.805 110.640 148.995 ;
        RECT 109.220 147.675 109.720 148.055 ;
        RECT 109.890 148.005 110.300 148.625 ;
        RECT 110.470 147.835 110.640 148.805 ;
        RECT 109.945 147.665 110.640 147.835 ;
        RECT 108.260 146.995 108.640 147.375 ;
        RECT 108.880 147.210 109.710 147.380 ;
        RECT 109.945 147.165 110.115 147.665 ;
        RECT 110.285 146.995 110.615 147.495 ;
        RECT 110.830 147.165 111.055 149.285 ;
        RECT 111.225 149.165 111.555 149.545 ;
        RECT 111.725 148.995 111.895 149.285 ;
        RECT 111.230 148.825 111.895 148.995 ;
        RECT 111.230 147.835 111.460 148.825 ;
        RECT 112.155 148.795 113.365 149.545 ;
        RECT 111.630 148.005 111.980 148.655 ;
        RECT 112.155 148.085 112.675 148.625 ;
        RECT 112.845 148.255 113.365 148.795 ;
        RECT 111.230 147.665 111.895 147.835 ;
        RECT 111.225 146.995 111.555 147.495 ;
        RECT 111.725 147.165 111.895 147.665 ;
        RECT 112.155 146.995 113.365 148.085 ;
        RECT 22.830 146.825 113.450 146.995 ;
        RECT 22.915 145.735 24.125 146.825 ;
        RECT 22.915 145.025 23.435 145.565 ;
        RECT 23.605 145.195 24.125 145.735 ;
        RECT 24.815 145.685 25.025 146.825 ;
        RECT 25.195 145.675 25.525 146.655 ;
        RECT 25.695 145.685 25.925 146.825 ;
        RECT 26.225 146.155 26.395 146.655 ;
        RECT 26.565 146.325 26.895 146.825 ;
        RECT 26.225 145.985 26.890 146.155 ;
        RECT 22.915 144.275 24.125 145.025 ;
        RECT 24.815 144.275 25.025 145.095 ;
        RECT 25.195 145.075 25.445 145.675 ;
        RECT 25.615 145.265 25.945 145.515 ;
        RECT 26.140 145.165 26.490 145.815 ;
        RECT 25.195 144.445 25.525 145.075 ;
        RECT 25.695 144.275 25.925 145.095 ;
        RECT 26.660 144.995 26.890 145.985 ;
        RECT 26.225 144.825 26.890 144.995 ;
        RECT 26.225 144.535 26.395 144.825 ;
        RECT 26.565 144.275 26.895 144.655 ;
        RECT 27.065 144.535 27.290 146.655 ;
        RECT 27.505 146.325 27.835 146.825 ;
        RECT 28.005 146.155 28.175 146.655 ;
        RECT 28.410 146.440 29.240 146.610 ;
        RECT 29.480 146.445 29.860 146.825 ;
        RECT 27.480 145.985 28.175 146.155 ;
        RECT 27.480 145.015 27.650 145.985 ;
        RECT 27.820 145.195 28.230 145.815 ;
        RECT 28.400 145.765 28.900 146.145 ;
        RECT 27.480 144.825 28.175 145.015 ;
        RECT 28.400 144.895 28.620 145.765 ;
        RECT 29.070 145.595 29.240 146.440 ;
        RECT 30.040 146.275 30.210 146.565 ;
        RECT 30.380 146.445 30.710 146.825 ;
        RECT 31.180 146.355 31.810 146.605 ;
        RECT 31.990 146.445 32.410 146.825 ;
        RECT 31.640 146.275 31.810 146.355 ;
        RECT 32.610 146.275 32.850 146.565 ;
        RECT 29.410 146.025 30.780 146.275 ;
        RECT 29.410 145.765 29.660 146.025 ;
        RECT 30.170 145.595 30.420 145.755 ;
        RECT 29.070 145.425 30.420 145.595 ;
        RECT 29.070 145.385 29.490 145.425 ;
        RECT 28.800 144.835 29.150 145.205 ;
        RECT 27.505 144.275 27.835 144.655 ;
        RECT 28.005 144.495 28.175 144.825 ;
        RECT 29.320 144.655 29.490 145.385 ;
        RECT 30.590 145.255 30.780 146.025 ;
        RECT 29.660 144.925 30.070 145.255 ;
        RECT 30.360 144.915 30.780 145.255 ;
        RECT 30.950 145.845 31.470 146.155 ;
        RECT 31.640 146.105 32.850 146.275 ;
        RECT 33.080 146.135 33.410 146.825 ;
        RECT 30.950 145.085 31.120 145.845 ;
        RECT 31.290 145.255 31.470 145.665 ;
        RECT 31.640 145.595 31.810 146.105 ;
        RECT 33.580 145.955 33.750 146.565 ;
        RECT 34.020 146.105 34.350 146.615 ;
        RECT 33.580 145.935 33.900 145.955 ;
        RECT 31.980 145.765 33.900 145.935 ;
        RECT 31.640 145.425 33.540 145.595 ;
        RECT 31.870 145.085 32.200 145.205 ;
        RECT 30.950 144.915 32.200 145.085 ;
        RECT 28.475 144.455 29.490 144.655 ;
        RECT 29.660 144.275 30.070 144.715 ;
        RECT 30.360 144.485 30.610 144.915 ;
        RECT 30.810 144.275 31.130 144.735 ;
        RECT 32.370 144.665 32.540 145.425 ;
        RECT 33.210 145.365 33.540 145.425 ;
        RECT 32.730 145.195 33.060 145.255 ;
        RECT 32.730 144.925 33.390 145.195 ;
        RECT 33.710 144.870 33.900 145.765 ;
        RECT 31.690 144.495 32.540 144.665 ;
        RECT 32.740 144.275 33.400 144.755 ;
        RECT 33.580 144.540 33.900 144.870 ;
        RECT 34.100 145.515 34.350 146.105 ;
        RECT 34.530 146.025 34.815 146.825 ;
        RECT 34.995 146.485 35.250 146.515 ;
        RECT 34.995 146.315 35.335 146.485 ;
        RECT 34.995 145.845 35.250 146.315 ;
        RECT 34.100 145.185 34.900 145.515 ;
        RECT 34.100 144.535 34.350 145.185 ;
        RECT 35.070 144.985 35.250 145.845 ;
        RECT 35.795 145.660 36.085 146.825 ;
        RECT 36.915 146.155 37.195 146.825 ;
        RECT 37.365 145.935 37.665 146.485 ;
        RECT 37.865 146.105 38.195 146.825 ;
        RECT 38.385 146.105 38.845 146.655 ;
        RECT 36.730 145.515 36.995 145.875 ;
        RECT 37.365 145.765 38.305 145.935 ;
        RECT 38.135 145.515 38.305 145.765 ;
        RECT 36.730 145.265 37.405 145.515 ;
        RECT 37.625 145.265 37.965 145.515 ;
        RECT 38.135 145.185 38.425 145.515 ;
        RECT 38.135 145.095 38.305 145.185 ;
        RECT 34.530 144.275 34.815 144.735 ;
        RECT 34.995 144.455 35.250 144.985 ;
        RECT 35.795 144.275 36.085 145.000 ;
        RECT 36.915 144.905 38.305 145.095 ;
        RECT 36.915 144.545 37.245 144.905 ;
        RECT 38.595 144.735 38.845 146.105 ;
        RECT 37.865 144.275 38.115 144.735 ;
        RECT 38.285 144.445 38.845 144.735 ;
        RECT 39.020 145.685 39.355 146.655 ;
        RECT 39.525 145.685 39.695 146.825 ;
        RECT 39.865 146.485 41.895 146.655 ;
        RECT 39.020 145.015 39.190 145.685 ;
        RECT 39.865 145.515 40.035 146.485 ;
        RECT 39.360 145.185 39.615 145.515 ;
        RECT 39.840 145.185 40.035 145.515 ;
        RECT 40.205 146.145 41.330 146.315 ;
        RECT 39.445 145.015 39.615 145.185 ;
        RECT 40.205 145.015 40.375 146.145 ;
        RECT 39.020 144.445 39.275 145.015 ;
        RECT 39.445 144.845 40.375 145.015 ;
        RECT 40.545 145.805 41.555 145.975 ;
        RECT 40.545 145.005 40.715 145.805 ;
        RECT 40.200 144.810 40.375 144.845 ;
        RECT 39.445 144.275 39.775 144.675 ;
        RECT 40.200 144.445 40.730 144.810 ;
        RECT 40.920 144.785 41.195 145.605 ;
        RECT 40.915 144.615 41.195 144.785 ;
        RECT 40.920 144.445 41.195 144.615 ;
        RECT 41.365 144.445 41.555 145.805 ;
        RECT 41.725 145.820 41.895 146.485 ;
        RECT 42.065 146.065 42.235 146.825 ;
        RECT 42.470 146.065 42.985 146.475 ;
        RECT 44.275 146.155 44.555 146.825 ;
        RECT 41.725 145.630 42.475 145.820 ;
        RECT 42.645 145.255 42.985 146.065 ;
        RECT 44.725 145.935 45.025 146.485 ;
        RECT 45.225 146.105 45.555 146.825 ;
        RECT 45.745 146.105 46.205 146.655 ;
        RECT 46.575 146.155 46.855 146.825 ;
        RECT 44.090 145.515 44.355 145.875 ;
        RECT 44.725 145.765 45.665 145.935 ;
        RECT 45.495 145.515 45.665 145.765 ;
        RECT 44.090 145.265 44.765 145.515 ;
        RECT 44.985 145.265 45.325 145.515 ;
        RECT 41.755 145.085 42.985 145.255 ;
        RECT 45.495 145.185 45.785 145.515 ;
        RECT 45.495 145.095 45.665 145.185 ;
        RECT 41.735 144.275 42.245 144.810 ;
        RECT 42.465 144.480 42.710 145.085 ;
        RECT 44.275 144.905 45.665 145.095 ;
        RECT 44.275 144.545 44.605 144.905 ;
        RECT 45.955 144.735 46.205 146.105 ;
        RECT 47.025 145.935 47.325 146.485 ;
        RECT 47.525 146.105 47.855 146.825 ;
        RECT 48.045 146.105 48.505 146.655 ;
        RECT 46.390 145.515 46.655 145.875 ;
        RECT 47.025 145.765 47.965 145.935 ;
        RECT 47.795 145.515 47.965 145.765 ;
        RECT 46.390 145.265 47.065 145.515 ;
        RECT 47.285 145.265 47.625 145.515 ;
        RECT 47.795 145.185 48.085 145.515 ;
        RECT 47.795 145.095 47.965 145.185 ;
        RECT 45.225 144.275 45.475 144.735 ;
        RECT 45.645 144.445 46.205 144.735 ;
        RECT 46.575 144.905 47.965 145.095 ;
        RECT 46.575 144.545 46.905 144.905 ;
        RECT 48.255 144.735 48.505 146.105 ;
        RECT 49.135 145.735 51.725 146.825 ;
        RECT 51.900 146.315 53.555 146.605 ;
        RECT 51.900 145.975 53.490 146.145 ;
        RECT 53.725 146.025 54.005 146.825 ;
        RECT 49.135 145.215 50.345 145.735 ;
        RECT 51.900 145.685 52.220 145.975 ;
        RECT 53.320 145.855 53.490 145.975 ;
        RECT 50.515 145.045 51.725 145.565 ;
        RECT 47.525 144.275 47.775 144.735 ;
        RECT 47.945 144.445 48.505 144.735 ;
        RECT 49.135 144.275 51.725 145.045 ;
        RECT 51.900 144.945 52.250 145.515 ;
        RECT 52.420 145.185 53.130 145.805 ;
        RECT 53.320 145.685 54.045 145.855 ;
        RECT 54.215 145.685 54.485 146.655 ;
        RECT 53.875 145.515 54.045 145.685 ;
        RECT 53.300 145.185 53.705 145.515 ;
        RECT 53.875 145.185 54.145 145.515 ;
        RECT 53.875 145.015 54.045 145.185 ;
        RECT 52.435 144.845 54.045 145.015 ;
        RECT 54.315 144.950 54.485 145.685 ;
        RECT 54.655 145.735 57.245 146.825 ;
        RECT 57.420 146.315 59.075 146.605 ;
        RECT 57.420 145.975 59.010 146.145 ;
        RECT 59.245 146.025 59.525 146.825 ;
        RECT 54.655 145.215 55.865 145.735 ;
        RECT 57.420 145.685 57.740 145.975 ;
        RECT 58.840 145.855 59.010 145.975 ;
        RECT 56.035 145.045 57.245 145.565 ;
        RECT 51.905 144.275 52.235 144.775 ;
        RECT 52.435 144.495 52.605 144.845 ;
        RECT 52.805 144.275 53.135 144.675 ;
        RECT 53.305 144.495 53.475 144.845 ;
        RECT 53.645 144.275 54.025 144.675 ;
        RECT 54.215 144.605 54.485 144.950 ;
        RECT 54.655 144.275 57.245 145.045 ;
        RECT 57.420 144.945 57.770 145.515 ;
        RECT 57.940 145.185 58.650 145.805 ;
        RECT 58.840 145.685 59.565 145.855 ;
        RECT 59.735 145.685 60.005 146.655 ;
        RECT 59.395 145.515 59.565 145.685 ;
        RECT 58.820 145.185 59.225 145.515 ;
        RECT 59.395 145.185 59.665 145.515 ;
        RECT 59.395 145.015 59.565 145.185 ;
        RECT 57.955 144.845 59.565 145.015 ;
        RECT 59.835 144.950 60.005 145.685 ;
        RECT 60.175 145.735 61.385 146.825 ;
        RECT 60.175 145.195 60.695 145.735 ;
        RECT 61.555 145.660 61.845 146.825 ;
        RECT 62.015 146.065 62.530 146.475 ;
        RECT 62.765 146.065 62.935 146.825 ;
        RECT 63.105 146.485 65.135 146.655 ;
        RECT 60.865 145.025 61.385 145.565 ;
        RECT 62.015 145.255 62.355 146.065 ;
        RECT 63.105 145.820 63.275 146.485 ;
        RECT 63.670 146.145 64.795 146.315 ;
        RECT 62.525 145.630 63.275 145.820 ;
        RECT 63.445 145.805 64.455 145.975 ;
        RECT 62.015 145.085 63.245 145.255 ;
        RECT 57.425 144.275 57.755 144.775 ;
        RECT 57.955 144.495 58.125 144.845 ;
        RECT 58.325 144.275 58.655 144.675 ;
        RECT 58.825 144.495 58.995 144.845 ;
        RECT 59.165 144.275 59.545 144.675 ;
        RECT 59.735 144.605 60.005 144.950 ;
        RECT 60.175 144.275 61.385 145.025 ;
        RECT 61.555 144.275 61.845 145.000 ;
        RECT 62.290 144.480 62.535 145.085 ;
        RECT 62.755 144.275 63.265 144.810 ;
        RECT 63.445 144.445 63.635 145.805 ;
        RECT 63.805 145.465 64.080 145.605 ;
        RECT 63.805 145.295 64.085 145.465 ;
        RECT 63.805 144.445 64.080 145.295 ;
        RECT 64.285 145.005 64.455 145.805 ;
        RECT 64.625 145.015 64.795 146.145 ;
        RECT 64.965 145.515 65.135 146.485 ;
        RECT 65.305 145.685 65.475 146.825 ;
        RECT 65.645 145.685 65.980 146.655 ;
        RECT 64.965 145.185 65.160 145.515 ;
        RECT 65.385 145.185 65.640 145.515 ;
        RECT 65.385 145.015 65.555 145.185 ;
        RECT 65.810 145.015 65.980 145.685 ;
        RECT 64.625 144.845 65.555 145.015 ;
        RECT 64.625 144.810 64.800 144.845 ;
        RECT 64.270 144.445 64.800 144.810 ;
        RECT 65.225 144.275 65.555 144.675 ;
        RECT 65.725 144.445 65.980 145.015 ;
        RECT 66.155 145.855 66.425 146.625 ;
        RECT 66.595 146.045 66.925 146.825 ;
        RECT 67.130 146.220 67.315 146.625 ;
        RECT 67.485 146.400 67.820 146.825 ;
        RECT 67.130 146.045 67.795 146.220 ;
        RECT 66.155 145.685 67.285 145.855 ;
        RECT 66.155 144.775 66.325 145.685 ;
        RECT 66.495 144.935 66.855 145.515 ;
        RECT 67.035 145.185 67.285 145.685 ;
        RECT 67.455 145.015 67.795 146.045 ;
        RECT 68.085 145.895 68.255 146.655 ;
        RECT 68.435 146.065 68.765 146.825 ;
        RECT 68.085 145.725 68.750 145.895 ;
        RECT 68.935 145.750 69.205 146.655 ;
        RECT 68.580 145.580 68.750 145.725 ;
        RECT 68.015 145.175 68.345 145.545 ;
        RECT 68.580 145.250 68.865 145.580 ;
        RECT 67.110 144.845 67.795 145.015 ;
        RECT 68.580 144.995 68.750 145.250 ;
        RECT 66.155 144.445 66.415 144.775 ;
        RECT 66.625 144.275 66.900 144.755 ;
        RECT 67.110 144.445 67.315 144.845 ;
        RECT 68.085 144.825 68.750 144.995 ;
        RECT 69.035 144.950 69.205 145.750 ;
        RECT 69.375 145.735 70.585 146.825 ;
        RECT 70.755 145.735 74.265 146.825 ;
        RECT 74.640 145.855 74.970 146.655 ;
        RECT 75.140 146.025 75.470 146.825 ;
        RECT 75.770 145.855 76.100 146.655 ;
        RECT 76.745 146.025 76.995 146.825 ;
        RECT 69.375 145.195 69.895 145.735 ;
        RECT 70.065 145.025 70.585 145.565 ;
        RECT 70.755 145.215 72.445 145.735 ;
        RECT 74.640 145.685 77.075 145.855 ;
        RECT 77.265 145.685 77.435 146.825 ;
        RECT 77.605 145.685 77.945 146.655 ;
        RECT 72.615 145.045 74.265 145.565 ;
        RECT 74.435 145.265 74.785 145.515 ;
        RECT 74.970 145.055 75.140 145.685 ;
        RECT 75.310 145.265 75.640 145.465 ;
        RECT 75.810 145.265 76.140 145.465 ;
        RECT 76.310 145.265 76.730 145.465 ;
        RECT 76.905 145.435 77.075 145.685 ;
        RECT 76.905 145.265 77.600 145.435 ;
        RECT 67.485 144.275 67.820 144.675 ;
        RECT 68.085 144.445 68.255 144.825 ;
        RECT 68.435 144.275 68.765 144.655 ;
        RECT 68.945 144.445 69.205 144.950 ;
        RECT 69.375 144.275 70.585 145.025 ;
        RECT 70.755 144.275 74.265 145.045 ;
        RECT 74.640 144.445 75.140 145.055 ;
        RECT 75.770 144.925 76.995 145.095 ;
        RECT 77.770 145.075 77.945 145.685 ;
        RECT 78.115 145.735 79.325 146.825 ;
        RECT 79.495 146.065 80.010 146.475 ;
        RECT 80.245 146.065 80.415 146.825 ;
        RECT 80.585 146.485 82.615 146.655 ;
        RECT 78.115 145.195 78.635 145.735 ;
        RECT 75.770 144.445 76.100 144.925 ;
        RECT 76.270 144.275 76.495 144.735 ;
        RECT 76.665 144.445 76.995 144.925 ;
        RECT 77.185 144.275 77.435 145.075 ;
        RECT 77.605 144.445 77.945 145.075 ;
        RECT 78.805 145.025 79.325 145.565 ;
        RECT 79.495 145.255 79.835 146.065 ;
        RECT 80.585 145.820 80.755 146.485 ;
        RECT 81.150 146.145 82.275 146.315 ;
        RECT 80.005 145.630 80.755 145.820 ;
        RECT 80.925 145.805 81.935 145.975 ;
        RECT 79.495 145.085 80.725 145.255 ;
        RECT 78.115 144.275 79.325 145.025 ;
        RECT 79.770 144.480 80.015 145.085 ;
        RECT 80.235 144.275 80.745 144.810 ;
        RECT 80.925 144.445 81.115 145.805 ;
        RECT 81.285 145.125 81.560 145.605 ;
        RECT 81.285 144.955 81.565 145.125 ;
        RECT 81.765 145.005 81.935 145.805 ;
        RECT 82.105 145.015 82.275 146.145 ;
        RECT 82.445 145.515 82.615 146.485 ;
        RECT 82.785 145.685 82.955 146.825 ;
        RECT 83.125 145.685 83.460 146.655 ;
        RECT 83.725 145.895 83.895 146.655 ;
        RECT 84.075 146.065 84.405 146.825 ;
        RECT 83.725 145.725 84.390 145.895 ;
        RECT 84.575 145.750 84.845 146.655 ;
        RECT 82.445 145.185 82.640 145.515 ;
        RECT 82.865 145.185 83.120 145.515 ;
        RECT 82.865 145.015 83.035 145.185 ;
        RECT 83.290 145.015 83.460 145.685 ;
        RECT 84.220 145.580 84.390 145.725 ;
        RECT 83.655 145.175 83.985 145.545 ;
        RECT 84.220 145.250 84.505 145.580 ;
        RECT 81.285 144.445 81.560 144.955 ;
        RECT 82.105 144.845 83.035 145.015 ;
        RECT 82.105 144.810 82.280 144.845 ;
        RECT 81.750 144.445 82.280 144.810 ;
        RECT 82.705 144.275 83.035 144.675 ;
        RECT 83.205 144.445 83.460 145.015 ;
        RECT 84.220 144.995 84.390 145.250 ;
        RECT 83.725 144.825 84.390 144.995 ;
        RECT 84.675 144.950 84.845 145.750 ;
        RECT 85.475 145.735 87.145 146.825 ;
        RECT 85.475 145.215 86.225 145.735 ;
        RECT 87.315 145.660 87.605 146.825 ;
        RECT 87.975 146.155 88.255 146.825 ;
        RECT 88.425 145.935 88.725 146.485 ;
        RECT 88.925 146.105 89.255 146.825 ;
        RECT 89.445 146.105 89.905 146.655 ;
        RECT 86.395 145.045 87.145 145.565 ;
        RECT 87.790 145.515 88.055 145.875 ;
        RECT 88.425 145.765 89.365 145.935 ;
        RECT 89.195 145.515 89.365 145.765 ;
        RECT 87.790 145.265 88.465 145.515 ;
        RECT 88.685 145.265 89.025 145.515 ;
        RECT 89.195 145.185 89.485 145.515 ;
        RECT 89.195 145.095 89.365 145.185 ;
        RECT 83.725 144.445 83.895 144.825 ;
        RECT 84.075 144.275 84.405 144.655 ;
        RECT 84.585 144.445 84.845 144.950 ;
        RECT 85.475 144.275 87.145 145.045 ;
        RECT 87.315 144.275 87.605 145.000 ;
        RECT 87.975 144.905 89.365 145.095 ;
        RECT 87.975 144.545 88.305 144.905 ;
        RECT 89.655 144.735 89.905 146.105 ;
        RECT 90.075 146.065 90.590 146.475 ;
        RECT 90.825 146.065 90.995 146.825 ;
        RECT 91.165 146.485 93.195 146.655 ;
        RECT 90.075 145.255 90.415 146.065 ;
        RECT 91.165 145.820 91.335 146.485 ;
        RECT 91.730 146.145 92.855 146.315 ;
        RECT 90.585 145.630 91.335 145.820 ;
        RECT 91.505 145.805 92.515 145.975 ;
        RECT 90.075 145.085 91.305 145.255 ;
        RECT 88.925 144.275 89.175 144.735 ;
        RECT 89.345 144.445 89.905 144.735 ;
        RECT 90.350 144.480 90.595 145.085 ;
        RECT 90.815 144.275 91.325 144.810 ;
        RECT 91.505 144.445 91.695 145.805 ;
        RECT 91.865 145.125 92.140 145.605 ;
        RECT 91.865 144.955 92.145 145.125 ;
        RECT 92.345 145.005 92.515 145.805 ;
        RECT 92.685 145.015 92.855 146.145 ;
        RECT 93.025 145.515 93.195 146.485 ;
        RECT 93.365 145.685 93.535 146.825 ;
        RECT 93.705 145.685 94.040 146.655 ;
        RECT 93.025 145.185 93.220 145.515 ;
        RECT 93.445 145.185 93.700 145.515 ;
        RECT 93.445 145.015 93.615 145.185 ;
        RECT 93.870 145.015 94.040 145.685 ;
        RECT 91.865 144.445 92.140 144.955 ;
        RECT 92.685 144.845 93.615 145.015 ;
        RECT 92.685 144.810 92.860 144.845 ;
        RECT 92.330 144.445 92.860 144.810 ;
        RECT 93.285 144.275 93.615 144.675 ;
        RECT 93.785 144.445 94.040 145.015 ;
        RECT 94.215 146.105 94.675 146.655 ;
        RECT 94.865 146.105 95.195 146.825 ;
        RECT 94.215 144.735 94.465 146.105 ;
        RECT 95.395 145.935 95.695 146.485 ;
        RECT 95.865 146.155 96.145 146.825 ;
        RECT 94.755 145.765 95.695 145.935 ;
        RECT 96.975 146.105 97.435 146.655 ;
        RECT 97.625 146.105 97.955 146.825 ;
        RECT 94.755 145.515 94.925 145.765 ;
        RECT 96.065 145.515 96.330 145.875 ;
        RECT 94.635 145.185 94.925 145.515 ;
        RECT 95.095 145.265 95.435 145.515 ;
        RECT 95.655 145.265 96.330 145.515 ;
        RECT 94.755 145.095 94.925 145.185 ;
        RECT 94.755 144.905 96.145 145.095 ;
        RECT 94.215 144.445 94.775 144.735 ;
        RECT 94.945 144.275 95.195 144.735 ;
        RECT 95.815 144.545 96.145 144.905 ;
        RECT 96.975 144.735 97.225 146.105 ;
        RECT 98.155 145.935 98.455 146.485 ;
        RECT 98.625 146.155 98.905 146.825 ;
        RECT 97.515 145.765 98.455 145.935 ;
        RECT 97.515 145.515 97.685 145.765 ;
        RECT 98.825 145.515 99.090 145.875 ;
        RECT 97.395 145.185 97.685 145.515 ;
        RECT 97.855 145.265 98.195 145.515 ;
        RECT 98.415 145.265 99.090 145.515 ;
        RECT 99.275 145.735 101.865 146.825 ;
        RECT 102.035 146.065 102.550 146.475 ;
        RECT 102.785 146.065 102.955 146.825 ;
        RECT 103.125 146.485 105.155 146.655 ;
        RECT 99.275 145.215 100.485 145.735 ;
        RECT 97.515 145.095 97.685 145.185 ;
        RECT 97.515 144.905 98.905 145.095 ;
        RECT 100.655 145.045 101.865 145.565 ;
        RECT 102.035 145.255 102.375 146.065 ;
        RECT 103.125 145.820 103.295 146.485 ;
        RECT 103.690 146.145 104.815 146.315 ;
        RECT 102.545 145.630 103.295 145.820 ;
        RECT 103.465 145.805 104.475 145.975 ;
        RECT 102.035 145.085 103.265 145.255 ;
        RECT 96.975 144.445 97.535 144.735 ;
        RECT 97.705 144.275 97.955 144.735 ;
        RECT 98.575 144.545 98.905 144.905 ;
        RECT 99.275 144.275 101.865 145.045 ;
        RECT 102.310 144.480 102.555 145.085 ;
        RECT 102.775 144.275 103.285 144.810 ;
        RECT 103.465 144.445 103.655 145.805 ;
        RECT 103.825 145.465 104.100 145.605 ;
        RECT 103.825 145.295 104.105 145.465 ;
        RECT 103.825 144.445 104.100 145.295 ;
        RECT 104.305 145.005 104.475 145.805 ;
        RECT 104.645 145.015 104.815 146.145 ;
        RECT 104.985 145.515 105.155 146.485 ;
        RECT 105.325 145.685 105.495 146.825 ;
        RECT 105.665 145.685 106.000 146.655 ;
        RECT 104.985 145.185 105.180 145.515 ;
        RECT 105.405 145.185 105.660 145.515 ;
        RECT 105.405 145.015 105.575 145.185 ;
        RECT 105.830 145.015 106.000 145.685 ;
        RECT 106.175 145.735 107.385 146.825 ;
        RECT 107.645 145.895 107.815 146.655 ;
        RECT 107.995 146.065 108.325 146.825 ;
        RECT 106.175 145.195 106.695 145.735 ;
        RECT 107.645 145.725 108.310 145.895 ;
        RECT 108.495 145.750 108.765 146.655 ;
        RECT 108.140 145.580 108.310 145.725 ;
        RECT 106.865 145.025 107.385 145.565 ;
        RECT 107.575 145.175 107.905 145.545 ;
        RECT 108.140 145.250 108.425 145.580 ;
        RECT 104.645 144.845 105.575 145.015 ;
        RECT 104.645 144.810 104.820 144.845 ;
        RECT 104.290 144.445 104.820 144.810 ;
        RECT 105.245 144.275 105.575 144.675 ;
        RECT 105.745 144.445 106.000 145.015 ;
        RECT 106.175 144.275 107.385 145.025 ;
        RECT 108.140 144.995 108.310 145.250 ;
        RECT 107.645 144.825 108.310 144.995 ;
        RECT 108.595 144.950 108.765 145.750 ;
        RECT 109.395 145.735 111.985 146.825 ;
        RECT 112.155 145.735 113.365 146.825 ;
        RECT 109.395 145.215 110.605 145.735 ;
        RECT 110.775 145.045 111.985 145.565 ;
        RECT 112.155 145.195 112.675 145.735 ;
        RECT 107.645 144.445 107.815 144.825 ;
        RECT 107.995 144.275 108.325 144.655 ;
        RECT 108.505 144.445 108.765 144.950 ;
        RECT 109.395 144.275 111.985 145.045 ;
        RECT 112.845 145.025 113.365 145.565 ;
        RECT 112.155 144.275 113.365 145.025 ;
        RECT 22.830 144.105 113.450 144.275 ;
        RECT 22.915 143.355 24.125 144.105 ;
        RECT 22.915 142.815 23.435 143.355 ;
        RECT 24.755 143.335 26.425 144.105 ;
        RECT 23.605 142.645 24.125 143.185 ;
        RECT 22.915 141.555 24.125 142.645 ;
        RECT 24.755 142.645 25.505 143.165 ;
        RECT 25.675 142.815 26.425 143.335 ;
        RECT 26.635 143.285 26.865 144.105 ;
        RECT 27.035 143.305 27.365 143.935 ;
        RECT 26.615 142.865 26.945 143.115 ;
        RECT 27.115 142.705 27.365 143.305 ;
        RECT 27.535 143.285 27.745 144.105 ;
        RECT 28.065 143.555 28.235 143.935 ;
        RECT 28.415 143.725 28.745 144.105 ;
        RECT 28.065 143.385 28.730 143.555 ;
        RECT 28.925 143.430 29.185 143.935 ;
        RECT 27.995 142.835 28.325 143.205 ;
        RECT 28.560 143.130 28.730 143.385 ;
        RECT 24.755 141.555 26.425 142.645 ;
        RECT 26.635 141.555 26.865 142.695 ;
        RECT 27.035 141.725 27.365 142.705 ;
        RECT 28.560 142.800 28.845 143.130 ;
        RECT 27.535 141.555 27.745 142.695 ;
        RECT 28.560 142.655 28.730 142.800 ;
        RECT 28.065 142.485 28.730 142.655 ;
        RECT 29.015 142.630 29.185 143.430 ;
        RECT 28.065 141.725 28.235 142.485 ;
        RECT 28.415 141.555 28.745 142.315 ;
        RECT 28.915 141.725 29.185 142.630 ;
        RECT 29.355 143.430 29.615 143.935 ;
        RECT 29.795 143.725 30.125 144.105 ;
        RECT 30.305 143.555 30.475 143.935 ;
        RECT 29.355 142.630 29.525 143.430 ;
        RECT 29.810 143.385 30.475 143.555 ;
        RECT 29.810 143.130 29.980 143.385 ;
        RECT 30.775 143.285 31.005 144.105 ;
        RECT 31.175 143.305 31.505 143.935 ;
        RECT 29.695 142.800 29.980 143.130 ;
        RECT 30.215 142.835 30.545 143.205 ;
        RECT 30.755 142.865 31.085 143.115 ;
        RECT 29.810 142.655 29.980 142.800 ;
        RECT 31.255 142.705 31.505 143.305 ;
        RECT 31.675 143.285 31.885 144.105 ;
        RECT 32.120 143.365 32.375 143.935 ;
        RECT 32.545 143.705 32.875 144.105 ;
        RECT 33.300 143.570 33.830 143.935 ;
        RECT 34.020 143.765 34.295 143.935 ;
        RECT 34.015 143.595 34.295 143.765 ;
        RECT 33.300 143.535 33.475 143.570 ;
        RECT 32.545 143.365 33.475 143.535 ;
        RECT 29.355 141.725 29.625 142.630 ;
        RECT 29.810 142.485 30.475 142.655 ;
        RECT 29.795 141.555 30.125 142.315 ;
        RECT 30.305 141.725 30.475 142.485 ;
        RECT 30.775 141.555 31.005 142.695 ;
        RECT 31.175 141.725 31.505 142.705 ;
        RECT 32.120 142.695 32.290 143.365 ;
        RECT 32.545 143.195 32.715 143.365 ;
        RECT 32.460 142.865 32.715 143.195 ;
        RECT 32.940 142.865 33.135 143.195 ;
        RECT 31.675 141.555 31.885 142.695 ;
        RECT 32.120 141.725 32.455 142.695 ;
        RECT 32.625 141.555 32.795 142.695 ;
        RECT 32.965 141.895 33.135 142.865 ;
        RECT 33.305 142.235 33.475 143.365 ;
        RECT 33.645 142.575 33.815 143.375 ;
        RECT 34.020 142.775 34.295 143.595 ;
        RECT 34.465 142.575 34.655 143.935 ;
        RECT 34.835 143.570 35.345 144.105 ;
        RECT 35.565 143.295 35.810 143.900 ;
        RECT 36.345 143.555 36.515 143.845 ;
        RECT 36.685 143.725 37.015 144.105 ;
        RECT 36.345 143.385 37.010 143.555 ;
        RECT 34.855 143.125 36.085 143.295 ;
        RECT 33.645 142.405 34.655 142.575 ;
        RECT 34.825 142.560 35.575 142.750 ;
        RECT 33.305 142.065 34.430 142.235 ;
        RECT 34.825 141.895 34.995 142.560 ;
        RECT 35.745 142.315 36.085 143.125 ;
        RECT 36.260 142.565 36.610 143.215 ;
        RECT 36.780 142.395 37.010 143.385 ;
        RECT 32.965 141.725 34.995 141.895 ;
        RECT 35.165 141.555 35.335 142.315 ;
        RECT 35.570 141.905 36.085 142.315 ;
        RECT 36.345 142.225 37.010 142.395 ;
        RECT 36.345 141.725 36.515 142.225 ;
        RECT 36.685 141.555 37.015 142.055 ;
        RECT 37.185 141.725 37.410 143.845 ;
        RECT 37.625 143.725 37.955 144.105 ;
        RECT 38.125 143.555 38.295 143.885 ;
        RECT 38.595 143.725 39.610 143.925 ;
        RECT 37.600 143.365 38.295 143.555 ;
        RECT 37.600 142.395 37.770 143.365 ;
        RECT 37.940 142.565 38.350 143.185 ;
        RECT 38.520 142.615 38.740 143.485 ;
        RECT 38.920 143.175 39.270 143.545 ;
        RECT 39.440 142.995 39.610 143.725 ;
        RECT 39.780 143.665 40.190 144.105 ;
        RECT 40.480 143.465 40.730 143.895 ;
        RECT 40.930 143.645 41.250 144.105 ;
        RECT 41.810 143.715 42.660 143.885 ;
        RECT 39.780 143.125 40.190 143.455 ;
        RECT 40.480 143.125 40.900 143.465 ;
        RECT 39.190 142.955 39.610 142.995 ;
        RECT 39.190 142.785 40.540 142.955 ;
        RECT 37.600 142.225 38.295 142.395 ;
        RECT 38.520 142.235 39.020 142.615 ;
        RECT 37.625 141.555 37.955 142.055 ;
        RECT 38.125 141.725 38.295 142.225 ;
        RECT 39.190 141.940 39.360 142.785 ;
        RECT 40.290 142.625 40.540 142.785 ;
        RECT 39.530 142.355 39.780 142.615 ;
        RECT 40.710 142.355 40.900 143.125 ;
        RECT 39.530 142.105 40.900 142.355 ;
        RECT 41.070 143.295 42.320 143.465 ;
        RECT 41.070 142.535 41.240 143.295 ;
        RECT 41.990 143.175 42.320 143.295 ;
        RECT 41.410 142.715 41.590 143.125 ;
        RECT 42.490 142.955 42.660 143.715 ;
        RECT 42.860 143.625 43.520 144.105 ;
        RECT 43.700 143.510 44.020 143.840 ;
        RECT 42.850 143.185 43.510 143.455 ;
        RECT 42.850 143.125 43.180 143.185 ;
        RECT 43.330 142.955 43.660 143.015 ;
        RECT 41.760 142.785 43.660 142.955 ;
        RECT 41.070 142.225 41.590 142.535 ;
        RECT 41.760 142.275 41.930 142.785 ;
        RECT 43.830 142.615 44.020 143.510 ;
        RECT 42.100 142.445 44.020 142.615 ;
        RECT 43.700 142.425 44.020 142.445 ;
        RECT 44.220 143.195 44.470 143.845 ;
        RECT 44.650 143.645 44.935 144.105 ;
        RECT 45.115 143.765 45.370 143.925 ;
        RECT 45.115 143.595 45.455 143.765 ;
        RECT 45.115 143.395 45.370 143.595 ;
        RECT 44.220 142.865 45.020 143.195 ;
        RECT 41.760 142.105 42.970 142.275 ;
        RECT 38.530 141.770 39.360 141.940 ;
        RECT 39.600 141.555 39.980 141.935 ;
        RECT 40.160 141.815 40.330 142.105 ;
        RECT 41.760 142.025 41.930 142.105 ;
        RECT 40.500 141.555 40.830 141.935 ;
        RECT 41.300 141.775 41.930 142.025 ;
        RECT 42.110 141.555 42.530 141.935 ;
        RECT 42.730 141.815 42.970 142.105 ;
        RECT 43.200 141.555 43.530 142.245 ;
        RECT 43.700 141.815 43.870 142.425 ;
        RECT 44.220 142.275 44.470 142.865 ;
        RECT 45.190 142.535 45.370 143.395 ;
        RECT 44.140 141.765 44.470 142.275 ;
        RECT 44.650 141.555 44.935 142.355 ;
        RECT 45.115 141.865 45.370 142.535 ;
        RECT 45.915 143.430 46.185 143.775 ;
        RECT 46.375 143.705 46.755 144.105 ;
        RECT 46.925 143.535 47.095 143.885 ;
        RECT 47.265 143.705 47.595 144.105 ;
        RECT 47.795 143.535 47.965 143.885 ;
        RECT 48.165 143.605 48.495 144.105 ;
        RECT 45.915 142.695 46.085 143.430 ;
        RECT 46.355 143.365 47.965 143.535 ;
        RECT 46.355 143.195 46.525 143.365 ;
        RECT 46.255 142.865 46.525 143.195 ;
        RECT 46.695 142.865 47.100 143.195 ;
        RECT 46.355 142.695 46.525 142.865 ;
        RECT 45.915 141.725 46.185 142.695 ;
        RECT 46.355 142.525 47.080 142.695 ;
        RECT 47.270 142.575 47.980 143.195 ;
        RECT 48.150 142.865 48.500 143.435 ;
        RECT 48.675 143.380 48.965 144.105 ;
        RECT 49.175 143.285 49.405 144.105 ;
        RECT 49.575 143.305 49.905 143.935 ;
        RECT 49.155 142.865 49.485 143.115 ;
        RECT 46.910 142.405 47.080 142.525 ;
        RECT 48.180 142.405 48.500 142.695 ;
        RECT 46.395 141.555 46.675 142.355 ;
        RECT 46.910 142.235 48.500 142.405 ;
        RECT 46.845 141.775 48.500 142.065 ;
        RECT 48.675 141.555 48.965 142.720 ;
        RECT 49.655 142.705 49.905 143.305 ;
        RECT 50.075 143.285 50.285 144.105 ;
        RECT 50.520 143.365 50.775 143.935 ;
        RECT 50.945 143.705 51.275 144.105 ;
        RECT 51.700 143.570 52.230 143.935 ;
        RECT 52.420 143.765 52.695 143.935 ;
        RECT 52.415 143.595 52.695 143.765 ;
        RECT 51.700 143.535 51.875 143.570 ;
        RECT 50.945 143.365 51.875 143.535 ;
        RECT 49.175 141.555 49.405 142.695 ;
        RECT 49.575 141.725 49.905 142.705 ;
        RECT 50.520 142.695 50.690 143.365 ;
        RECT 50.945 143.195 51.115 143.365 ;
        RECT 50.860 142.865 51.115 143.195 ;
        RECT 51.340 142.865 51.535 143.195 ;
        RECT 50.075 141.555 50.285 142.695 ;
        RECT 50.520 141.725 50.855 142.695 ;
        RECT 51.025 141.555 51.195 142.695 ;
        RECT 51.365 141.895 51.535 142.865 ;
        RECT 51.705 142.235 51.875 143.365 ;
        RECT 52.045 142.575 52.215 143.375 ;
        RECT 52.420 142.775 52.695 143.595 ;
        RECT 52.865 142.575 53.055 143.935 ;
        RECT 53.235 143.570 53.745 144.105 ;
        RECT 53.965 143.295 54.210 143.900 ;
        RECT 55.115 143.335 56.785 144.105 ;
        RECT 53.255 143.125 54.485 143.295 ;
        RECT 52.045 142.405 53.055 142.575 ;
        RECT 53.225 142.560 53.975 142.750 ;
        RECT 51.705 142.065 52.830 142.235 ;
        RECT 53.225 141.895 53.395 142.560 ;
        RECT 54.145 142.315 54.485 143.125 ;
        RECT 51.365 141.725 53.395 141.895 ;
        RECT 53.565 141.555 53.735 142.315 ;
        RECT 53.970 141.905 54.485 142.315 ;
        RECT 55.115 142.645 55.865 143.165 ;
        RECT 56.035 142.815 56.785 143.335 ;
        RECT 56.955 143.305 57.295 143.935 ;
        RECT 57.465 143.305 57.715 144.105 ;
        RECT 57.905 143.455 58.235 143.935 ;
        RECT 58.405 143.645 58.630 144.105 ;
        RECT 58.800 143.455 59.130 143.935 ;
        RECT 56.955 142.695 57.130 143.305 ;
        RECT 57.905 143.285 59.130 143.455 ;
        RECT 59.760 143.325 60.260 143.935 ;
        RECT 61.010 143.395 61.265 143.925 ;
        RECT 61.445 143.645 61.730 144.105 ;
        RECT 57.300 142.945 57.995 143.115 ;
        RECT 57.825 142.695 57.995 142.945 ;
        RECT 58.170 142.915 58.590 143.115 ;
        RECT 58.760 142.915 59.090 143.115 ;
        RECT 59.260 142.915 59.590 143.115 ;
        RECT 59.760 142.695 59.930 143.325 ;
        RECT 60.115 142.865 60.465 143.115 ;
        RECT 55.115 141.555 56.785 142.645 ;
        RECT 56.955 141.725 57.295 142.695 ;
        RECT 57.465 141.555 57.635 142.695 ;
        RECT 57.825 142.525 60.260 142.695 ;
        RECT 57.905 141.555 58.155 142.355 ;
        RECT 58.800 141.725 59.130 142.525 ;
        RECT 59.430 141.555 59.760 142.355 ;
        RECT 59.930 141.725 60.260 142.525 ;
        RECT 61.010 142.535 61.190 143.395 ;
        RECT 61.910 143.195 62.160 143.845 ;
        RECT 61.360 142.865 62.160 143.195 ;
        RECT 61.010 142.065 61.265 142.535 ;
        RECT 60.925 141.895 61.265 142.065 ;
        RECT 61.010 141.865 61.265 141.895 ;
        RECT 61.445 141.555 61.730 142.355 ;
        RECT 61.910 142.275 62.160 142.865 ;
        RECT 62.360 143.510 62.680 143.840 ;
        RECT 62.860 143.625 63.520 144.105 ;
        RECT 63.720 143.715 64.570 143.885 ;
        RECT 62.360 142.615 62.550 143.510 ;
        RECT 62.870 143.185 63.530 143.455 ;
        RECT 63.200 143.125 63.530 143.185 ;
        RECT 62.720 142.955 63.050 143.015 ;
        RECT 63.720 142.955 63.890 143.715 ;
        RECT 65.130 143.645 65.450 144.105 ;
        RECT 65.650 143.465 65.900 143.895 ;
        RECT 66.190 143.665 66.600 144.105 ;
        RECT 66.770 143.725 67.785 143.925 ;
        RECT 64.060 143.295 65.310 143.465 ;
        RECT 64.060 143.175 64.390 143.295 ;
        RECT 62.720 142.785 64.620 142.955 ;
        RECT 62.360 142.445 64.280 142.615 ;
        RECT 62.360 142.425 62.680 142.445 ;
        RECT 61.910 141.765 62.240 142.275 ;
        RECT 62.510 141.815 62.680 142.425 ;
        RECT 64.450 142.275 64.620 142.785 ;
        RECT 64.790 142.715 64.970 143.125 ;
        RECT 65.140 142.535 65.310 143.295 ;
        RECT 62.850 141.555 63.180 142.245 ;
        RECT 63.410 142.105 64.620 142.275 ;
        RECT 64.790 142.225 65.310 142.535 ;
        RECT 65.480 143.125 65.900 143.465 ;
        RECT 66.190 143.125 66.600 143.455 ;
        RECT 65.480 142.355 65.670 143.125 ;
        RECT 66.770 142.995 66.940 143.725 ;
        RECT 68.085 143.555 68.255 143.885 ;
        RECT 68.425 143.725 68.755 144.105 ;
        RECT 67.110 143.175 67.460 143.545 ;
        RECT 66.770 142.955 67.190 142.995 ;
        RECT 65.840 142.785 67.190 142.955 ;
        RECT 65.840 142.625 66.090 142.785 ;
        RECT 66.600 142.355 66.850 142.615 ;
        RECT 65.480 142.105 66.850 142.355 ;
        RECT 63.410 141.815 63.650 142.105 ;
        RECT 64.450 142.025 64.620 142.105 ;
        RECT 63.850 141.555 64.270 141.935 ;
        RECT 64.450 141.775 65.080 142.025 ;
        RECT 65.550 141.555 65.880 141.935 ;
        RECT 66.050 141.815 66.220 142.105 ;
        RECT 67.020 141.940 67.190 142.785 ;
        RECT 67.640 142.615 67.860 143.485 ;
        RECT 68.085 143.365 68.780 143.555 ;
        RECT 67.360 142.235 67.860 142.615 ;
        RECT 68.030 142.565 68.440 143.185 ;
        RECT 68.610 142.395 68.780 143.365 ;
        RECT 68.085 142.225 68.780 142.395 ;
        RECT 66.400 141.555 66.780 141.935 ;
        RECT 67.020 141.770 67.850 141.940 ;
        RECT 68.085 141.725 68.255 142.225 ;
        RECT 68.425 141.555 68.755 142.055 ;
        RECT 68.970 141.725 69.195 143.845 ;
        RECT 69.365 143.725 69.695 144.105 ;
        RECT 69.865 143.555 70.035 143.845 ;
        RECT 69.370 143.385 70.035 143.555 ;
        RECT 69.370 142.395 69.600 143.385 ;
        RECT 70.960 143.325 71.460 143.935 ;
        RECT 69.770 142.565 70.120 143.215 ;
        RECT 70.755 142.865 71.105 143.115 ;
        RECT 71.290 142.695 71.460 143.325 ;
        RECT 72.090 143.455 72.420 143.935 ;
        RECT 72.590 143.645 72.815 144.105 ;
        RECT 72.985 143.455 73.315 143.935 ;
        RECT 72.090 143.285 73.315 143.455 ;
        RECT 73.505 143.305 73.755 144.105 ;
        RECT 73.925 143.305 74.265 143.935 ;
        RECT 74.435 143.380 74.725 144.105 ;
        RECT 74.905 143.605 75.235 144.105 ;
        RECT 75.435 143.535 75.605 143.885 ;
        RECT 75.805 143.705 76.135 144.105 ;
        RECT 76.305 143.535 76.475 143.885 ;
        RECT 76.645 143.705 77.025 144.105 ;
        RECT 71.630 142.915 71.960 143.115 ;
        RECT 72.130 142.915 72.460 143.115 ;
        RECT 72.630 142.915 73.050 143.115 ;
        RECT 73.225 142.945 73.920 143.115 ;
        RECT 73.225 142.695 73.395 142.945 ;
        RECT 74.090 142.695 74.265 143.305 ;
        RECT 74.900 142.865 75.250 143.435 ;
        RECT 75.435 143.365 77.045 143.535 ;
        RECT 77.215 143.430 77.485 143.775 ;
        RECT 78.030 143.765 78.285 143.925 ;
        RECT 77.945 143.595 78.285 143.765 ;
        RECT 78.465 143.645 78.750 144.105 ;
        RECT 76.875 143.195 77.045 143.365 ;
        RECT 75.420 142.745 76.130 143.195 ;
        RECT 76.300 142.865 76.705 143.195 ;
        RECT 76.875 142.865 77.145 143.195 ;
        RECT 70.960 142.525 73.395 142.695 ;
        RECT 69.370 142.225 70.035 142.395 ;
        RECT 69.365 141.555 69.695 142.055 ;
        RECT 69.865 141.725 70.035 142.225 ;
        RECT 70.960 141.725 71.290 142.525 ;
        RECT 71.460 141.555 71.790 142.355 ;
        RECT 72.090 141.725 72.420 142.525 ;
        RECT 73.065 141.555 73.315 142.355 ;
        RECT 73.585 141.555 73.755 142.695 ;
        RECT 73.925 141.725 74.265 142.695 ;
        RECT 74.435 141.555 74.725 142.720 ;
        RECT 74.900 142.405 75.220 142.695 ;
        RECT 75.415 142.575 76.130 142.745 ;
        RECT 76.875 142.695 77.045 142.865 ;
        RECT 77.315 142.695 77.485 143.430 ;
        RECT 76.320 142.525 77.045 142.695 ;
        RECT 76.320 142.405 76.490 142.525 ;
        RECT 74.900 142.235 76.490 142.405 ;
        RECT 74.900 141.775 76.555 142.065 ;
        RECT 76.725 141.555 77.005 142.355 ;
        RECT 77.215 141.725 77.485 142.695 ;
        RECT 78.030 143.395 78.285 143.595 ;
        RECT 78.030 142.535 78.210 143.395 ;
        RECT 78.930 143.195 79.180 143.845 ;
        RECT 78.380 142.865 79.180 143.195 ;
        RECT 78.030 141.865 78.285 142.535 ;
        RECT 78.465 141.555 78.750 142.355 ;
        RECT 78.930 142.275 79.180 142.865 ;
        RECT 79.380 143.510 79.700 143.840 ;
        RECT 79.880 143.625 80.540 144.105 ;
        RECT 80.740 143.715 81.590 143.885 ;
        RECT 79.380 142.615 79.570 143.510 ;
        RECT 79.890 143.185 80.550 143.455 ;
        RECT 80.220 143.125 80.550 143.185 ;
        RECT 79.740 142.955 80.070 143.015 ;
        RECT 80.740 142.955 80.910 143.715 ;
        RECT 82.150 143.645 82.470 144.105 ;
        RECT 82.670 143.465 82.920 143.895 ;
        RECT 83.210 143.665 83.620 144.105 ;
        RECT 83.790 143.725 84.805 143.925 ;
        RECT 81.080 143.295 82.330 143.465 ;
        RECT 81.080 143.175 81.410 143.295 ;
        RECT 79.740 142.785 81.640 142.955 ;
        RECT 79.380 142.445 81.300 142.615 ;
        RECT 79.380 142.425 79.700 142.445 ;
        RECT 78.930 141.765 79.260 142.275 ;
        RECT 79.530 141.815 79.700 142.425 ;
        RECT 81.470 142.275 81.640 142.785 ;
        RECT 81.810 142.715 81.990 143.125 ;
        RECT 82.160 142.535 82.330 143.295 ;
        RECT 79.870 141.555 80.200 142.245 ;
        RECT 80.430 142.105 81.640 142.275 ;
        RECT 81.810 142.225 82.330 142.535 ;
        RECT 82.500 143.125 82.920 143.465 ;
        RECT 83.210 143.125 83.620 143.455 ;
        RECT 82.500 142.355 82.690 143.125 ;
        RECT 83.790 142.995 83.960 143.725 ;
        RECT 85.105 143.555 85.275 143.885 ;
        RECT 85.445 143.725 85.775 144.105 ;
        RECT 84.130 143.175 84.480 143.545 ;
        RECT 83.790 142.955 84.210 142.995 ;
        RECT 82.860 142.785 84.210 142.955 ;
        RECT 82.860 142.625 83.110 142.785 ;
        RECT 83.620 142.355 83.870 142.615 ;
        RECT 82.500 142.105 83.870 142.355 ;
        RECT 80.430 141.815 80.670 142.105 ;
        RECT 81.470 142.025 81.640 142.105 ;
        RECT 80.870 141.555 81.290 141.935 ;
        RECT 81.470 141.775 82.100 142.025 ;
        RECT 82.570 141.555 82.900 141.935 ;
        RECT 83.070 141.815 83.240 142.105 ;
        RECT 84.040 141.940 84.210 142.785 ;
        RECT 84.660 142.615 84.880 143.485 ;
        RECT 85.105 143.365 85.800 143.555 ;
        RECT 84.380 142.235 84.880 142.615 ;
        RECT 85.050 142.565 85.460 143.185 ;
        RECT 85.630 142.395 85.800 143.365 ;
        RECT 85.105 142.225 85.800 142.395 ;
        RECT 83.420 141.555 83.800 141.935 ;
        RECT 84.040 141.770 84.870 141.940 ;
        RECT 85.105 141.725 85.275 142.225 ;
        RECT 85.445 141.555 85.775 142.055 ;
        RECT 85.990 141.725 86.215 143.845 ;
        RECT 86.385 143.725 86.715 144.105 ;
        RECT 86.885 143.555 87.055 143.845 ;
        RECT 87.690 143.765 87.945 143.925 ;
        RECT 87.605 143.595 87.945 143.765 ;
        RECT 88.125 143.645 88.410 144.105 ;
        RECT 86.390 143.385 87.055 143.555 ;
        RECT 87.690 143.395 87.945 143.595 ;
        RECT 86.390 142.395 86.620 143.385 ;
        RECT 86.790 142.565 87.140 143.215 ;
        RECT 87.690 142.535 87.870 143.395 ;
        RECT 88.590 143.195 88.840 143.845 ;
        RECT 88.040 142.865 88.840 143.195 ;
        RECT 86.390 142.225 87.055 142.395 ;
        RECT 86.385 141.555 86.715 142.055 ;
        RECT 86.885 141.725 87.055 142.225 ;
        RECT 87.690 141.865 87.945 142.535 ;
        RECT 88.125 141.555 88.410 142.355 ;
        RECT 88.590 142.275 88.840 142.865 ;
        RECT 89.040 143.510 89.360 143.840 ;
        RECT 89.540 143.625 90.200 144.105 ;
        RECT 90.400 143.715 91.250 143.885 ;
        RECT 89.040 142.615 89.230 143.510 ;
        RECT 89.550 143.185 90.210 143.455 ;
        RECT 89.880 143.125 90.210 143.185 ;
        RECT 89.400 142.955 89.730 143.015 ;
        RECT 90.400 142.955 90.570 143.715 ;
        RECT 91.810 143.645 92.130 144.105 ;
        RECT 92.330 143.465 92.580 143.895 ;
        RECT 92.870 143.665 93.280 144.105 ;
        RECT 93.450 143.725 94.465 143.925 ;
        RECT 90.740 143.295 91.990 143.465 ;
        RECT 90.740 143.175 91.070 143.295 ;
        RECT 89.400 142.785 91.300 142.955 ;
        RECT 89.040 142.445 90.960 142.615 ;
        RECT 89.040 142.425 89.360 142.445 ;
        RECT 88.590 141.765 88.920 142.275 ;
        RECT 89.190 141.815 89.360 142.425 ;
        RECT 91.130 142.275 91.300 142.785 ;
        RECT 91.470 142.715 91.650 143.125 ;
        RECT 91.820 142.535 91.990 143.295 ;
        RECT 89.530 141.555 89.860 142.245 ;
        RECT 90.090 142.105 91.300 142.275 ;
        RECT 91.470 142.225 91.990 142.535 ;
        RECT 92.160 143.125 92.580 143.465 ;
        RECT 92.870 143.125 93.280 143.455 ;
        RECT 92.160 142.355 92.350 143.125 ;
        RECT 93.450 142.995 93.620 143.725 ;
        RECT 94.765 143.555 94.935 143.885 ;
        RECT 95.105 143.725 95.435 144.105 ;
        RECT 93.790 143.175 94.140 143.545 ;
        RECT 93.450 142.955 93.870 142.995 ;
        RECT 92.520 142.785 93.870 142.955 ;
        RECT 92.520 142.625 92.770 142.785 ;
        RECT 93.280 142.355 93.530 142.615 ;
        RECT 92.160 142.105 93.530 142.355 ;
        RECT 90.090 141.815 90.330 142.105 ;
        RECT 91.130 142.025 91.300 142.105 ;
        RECT 90.530 141.555 90.950 141.935 ;
        RECT 91.130 141.775 91.760 142.025 ;
        RECT 92.230 141.555 92.560 141.935 ;
        RECT 92.730 141.815 92.900 142.105 ;
        RECT 93.700 141.940 93.870 142.785 ;
        RECT 94.320 142.615 94.540 143.485 ;
        RECT 94.765 143.365 95.460 143.555 ;
        RECT 94.040 142.235 94.540 142.615 ;
        RECT 94.710 142.565 95.120 143.185 ;
        RECT 95.290 142.395 95.460 143.365 ;
        RECT 94.765 142.225 95.460 142.395 ;
        RECT 93.080 141.555 93.460 141.935 ;
        RECT 93.700 141.770 94.530 141.940 ;
        RECT 94.765 141.725 94.935 142.225 ;
        RECT 95.105 141.555 95.435 142.055 ;
        RECT 95.650 141.725 95.875 143.845 ;
        RECT 96.045 143.725 96.375 144.105 ;
        RECT 96.545 143.555 96.715 143.845 ;
        RECT 96.050 143.385 96.715 143.555 ;
        RECT 96.975 143.645 97.535 143.935 ;
        RECT 97.705 143.645 97.955 144.105 ;
        RECT 96.050 142.395 96.280 143.385 ;
        RECT 96.450 142.565 96.800 143.215 ;
        RECT 96.050 142.225 96.715 142.395 ;
        RECT 96.045 141.555 96.375 142.055 ;
        RECT 96.545 141.725 96.715 142.225 ;
        RECT 96.975 142.275 97.225 143.645 ;
        RECT 98.575 143.475 98.905 143.835 ;
        RECT 97.515 143.285 98.905 143.475 ;
        RECT 100.195 143.380 100.485 144.105 ;
        RECT 100.695 143.285 100.925 144.105 ;
        RECT 101.095 143.305 101.425 143.935 ;
        RECT 97.515 143.195 97.685 143.285 ;
        RECT 97.395 142.865 97.685 143.195 ;
        RECT 97.855 142.865 98.195 143.115 ;
        RECT 98.415 142.865 99.090 143.115 ;
        RECT 100.675 142.865 101.005 143.115 ;
        RECT 97.515 142.615 97.685 142.865 ;
        RECT 97.515 142.445 98.455 142.615 ;
        RECT 98.825 142.505 99.090 142.865 ;
        RECT 96.975 141.725 97.435 142.275 ;
        RECT 97.625 141.555 97.955 142.275 ;
        RECT 98.155 141.895 98.455 142.445 ;
        RECT 98.625 141.555 98.905 142.225 ;
        RECT 100.195 141.555 100.485 142.720 ;
        RECT 101.175 142.705 101.425 143.305 ;
        RECT 101.595 143.285 101.805 144.105 ;
        RECT 102.410 143.765 102.665 143.925 ;
        RECT 102.325 143.595 102.665 143.765 ;
        RECT 102.845 143.645 103.130 144.105 ;
        RECT 102.410 143.395 102.665 143.595 ;
        RECT 100.695 141.555 100.925 142.695 ;
        RECT 101.095 141.725 101.425 142.705 ;
        RECT 101.595 141.555 101.805 142.695 ;
        RECT 102.410 142.535 102.590 143.395 ;
        RECT 103.310 143.195 103.560 143.845 ;
        RECT 102.760 142.865 103.560 143.195 ;
        RECT 102.410 141.865 102.665 142.535 ;
        RECT 102.845 141.555 103.130 142.355 ;
        RECT 103.310 142.275 103.560 142.865 ;
        RECT 103.760 143.510 104.080 143.840 ;
        RECT 104.260 143.625 104.920 144.105 ;
        RECT 105.120 143.715 105.970 143.885 ;
        RECT 103.760 142.615 103.950 143.510 ;
        RECT 104.270 143.185 104.930 143.455 ;
        RECT 104.600 143.125 104.930 143.185 ;
        RECT 104.120 142.955 104.450 143.015 ;
        RECT 105.120 142.955 105.290 143.715 ;
        RECT 106.530 143.645 106.850 144.105 ;
        RECT 107.050 143.465 107.300 143.895 ;
        RECT 107.590 143.665 108.000 144.105 ;
        RECT 108.170 143.725 109.185 143.925 ;
        RECT 105.460 143.295 106.710 143.465 ;
        RECT 105.460 143.175 105.790 143.295 ;
        RECT 104.120 142.785 106.020 142.955 ;
        RECT 103.760 142.445 105.680 142.615 ;
        RECT 103.760 142.425 104.080 142.445 ;
        RECT 103.310 141.765 103.640 142.275 ;
        RECT 103.910 141.815 104.080 142.425 ;
        RECT 105.850 142.275 106.020 142.785 ;
        RECT 106.190 142.715 106.370 143.125 ;
        RECT 106.540 142.535 106.710 143.295 ;
        RECT 104.250 141.555 104.580 142.245 ;
        RECT 104.810 142.105 106.020 142.275 ;
        RECT 106.190 142.225 106.710 142.535 ;
        RECT 106.880 143.125 107.300 143.465 ;
        RECT 107.590 143.125 108.000 143.455 ;
        RECT 106.880 142.355 107.070 143.125 ;
        RECT 108.170 142.995 108.340 143.725 ;
        RECT 109.485 143.555 109.655 143.885 ;
        RECT 109.825 143.725 110.155 144.105 ;
        RECT 108.510 143.175 108.860 143.545 ;
        RECT 108.170 142.955 108.590 142.995 ;
        RECT 107.240 142.785 108.590 142.955 ;
        RECT 107.240 142.625 107.490 142.785 ;
        RECT 108.000 142.355 108.250 142.615 ;
        RECT 106.880 142.105 108.250 142.355 ;
        RECT 104.810 141.815 105.050 142.105 ;
        RECT 105.850 142.025 106.020 142.105 ;
        RECT 105.250 141.555 105.670 141.935 ;
        RECT 105.850 141.775 106.480 142.025 ;
        RECT 106.950 141.555 107.280 141.935 ;
        RECT 107.450 141.815 107.620 142.105 ;
        RECT 108.420 141.940 108.590 142.785 ;
        RECT 109.040 142.615 109.260 143.485 ;
        RECT 109.485 143.365 110.180 143.555 ;
        RECT 108.760 142.235 109.260 142.615 ;
        RECT 109.430 142.565 109.840 143.185 ;
        RECT 110.010 142.395 110.180 143.365 ;
        RECT 109.485 142.225 110.180 142.395 ;
        RECT 107.800 141.555 108.180 141.935 ;
        RECT 108.420 141.770 109.250 141.940 ;
        RECT 109.485 141.725 109.655 142.225 ;
        RECT 109.825 141.555 110.155 142.055 ;
        RECT 110.370 141.725 110.595 143.845 ;
        RECT 110.765 143.725 111.095 144.105 ;
        RECT 111.265 143.555 111.435 143.845 ;
        RECT 110.770 143.385 111.435 143.555 ;
        RECT 110.770 142.395 111.000 143.385 ;
        RECT 112.155 143.355 113.365 144.105 ;
        RECT 111.170 142.565 111.520 143.215 ;
        RECT 112.155 142.645 112.675 143.185 ;
        RECT 112.845 142.815 113.365 143.355 ;
        RECT 110.770 142.225 111.435 142.395 ;
        RECT 110.765 141.555 111.095 142.055 ;
        RECT 111.265 141.725 111.435 142.225 ;
        RECT 112.155 141.555 113.365 142.645 ;
        RECT 22.830 141.385 113.450 141.555 ;
        RECT 22.915 140.295 24.125 141.385 ;
        RECT 22.915 139.585 23.435 140.125 ;
        RECT 23.605 139.755 24.125 140.295 ;
        RECT 24.295 140.295 25.965 141.385 ;
        RECT 24.295 139.775 25.045 140.295 ;
        RECT 26.175 140.245 26.405 141.385 ;
        RECT 26.575 140.235 26.905 141.215 ;
        RECT 27.075 140.245 27.285 141.385 ;
        RECT 27.515 140.310 27.785 141.215 ;
        RECT 27.955 140.625 28.285 141.385 ;
        RECT 28.465 140.455 28.635 141.215 ;
        RECT 25.215 139.605 25.965 140.125 ;
        RECT 26.155 139.825 26.485 140.075 ;
        RECT 22.915 138.835 24.125 139.585 ;
        RECT 24.295 138.835 25.965 139.605 ;
        RECT 26.175 138.835 26.405 139.655 ;
        RECT 26.655 139.635 26.905 140.235 ;
        RECT 26.575 139.005 26.905 139.635 ;
        RECT 27.075 138.835 27.285 139.655 ;
        RECT 27.515 139.510 27.685 140.310 ;
        RECT 27.970 140.285 28.635 140.455 ;
        RECT 27.970 140.140 28.140 140.285 ;
        RECT 27.855 139.810 28.140 140.140 ;
        RECT 28.900 140.245 29.235 141.215 ;
        RECT 29.405 140.245 29.575 141.385 ;
        RECT 29.745 141.045 31.775 141.215 ;
        RECT 27.970 139.555 28.140 139.810 ;
        RECT 28.375 139.735 28.705 140.105 ;
        RECT 28.900 139.575 29.070 140.245 ;
        RECT 29.745 140.075 29.915 141.045 ;
        RECT 29.240 139.745 29.495 140.075 ;
        RECT 29.720 139.745 29.915 140.075 ;
        RECT 30.085 140.705 31.210 140.875 ;
        RECT 29.325 139.575 29.495 139.745 ;
        RECT 30.085 139.575 30.255 140.705 ;
        RECT 27.515 139.005 27.775 139.510 ;
        RECT 27.970 139.385 28.635 139.555 ;
        RECT 27.955 138.835 28.285 139.215 ;
        RECT 28.465 139.005 28.635 139.385 ;
        RECT 28.900 139.005 29.155 139.575 ;
        RECT 29.325 139.405 30.255 139.575 ;
        RECT 30.425 140.365 31.435 140.535 ;
        RECT 30.425 139.565 30.595 140.365 ;
        RECT 30.800 139.685 31.075 140.165 ;
        RECT 30.795 139.515 31.075 139.685 ;
        RECT 30.080 139.370 30.255 139.405 ;
        RECT 29.325 138.835 29.655 139.235 ;
        RECT 30.080 139.005 30.610 139.370 ;
        RECT 30.800 139.005 31.075 139.515 ;
        RECT 31.245 139.005 31.435 140.365 ;
        RECT 31.605 140.380 31.775 141.045 ;
        RECT 31.945 140.625 32.115 141.385 ;
        RECT 32.350 140.625 32.865 141.035 ;
        RECT 31.605 140.190 32.355 140.380 ;
        RECT 32.525 139.815 32.865 140.625 ;
        RECT 33.090 140.515 33.375 141.385 ;
        RECT 33.545 140.755 33.805 141.215 ;
        RECT 33.980 140.925 34.235 141.385 ;
        RECT 34.405 140.755 34.665 141.215 ;
        RECT 33.545 140.585 34.665 140.755 ;
        RECT 34.835 140.585 35.145 141.385 ;
        RECT 33.545 140.335 33.805 140.585 ;
        RECT 35.315 140.415 35.625 141.215 ;
        RECT 31.635 139.645 32.865 139.815 ;
        RECT 33.050 140.165 33.805 140.335 ;
        RECT 34.595 140.245 35.625 140.415 ;
        RECT 33.050 139.655 33.455 140.165 ;
        RECT 34.595 139.995 34.765 140.245 ;
        RECT 33.625 139.825 34.765 139.995 ;
        RECT 31.615 138.835 32.125 139.370 ;
        RECT 32.345 139.040 32.590 139.645 ;
        RECT 33.050 139.485 34.700 139.655 ;
        RECT 34.935 139.505 35.285 140.075 ;
        RECT 33.095 138.835 33.375 139.315 ;
        RECT 33.545 139.095 33.805 139.485 ;
        RECT 33.980 138.835 34.235 139.315 ;
        RECT 34.405 139.095 34.700 139.485 ;
        RECT 35.455 139.335 35.625 140.245 ;
        RECT 35.795 140.220 36.085 141.385 ;
        RECT 36.365 140.585 36.535 141.385 ;
        RECT 36.705 140.365 37.035 141.215 ;
        RECT 37.205 140.585 37.375 141.385 ;
        RECT 37.545 140.365 37.875 141.215 ;
        RECT 38.045 140.585 38.215 141.385 ;
        RECT 38.385 140.365 38.715 141.215 ;
        RECT 38.885 140.585 39.055 141.385 ;
        RECT 39.225 140.365 39.555 141.215 ;
        RECT 39.725 140.585 39.895 141.385 ;
        RECT 40.065 140.365 40.395 141.215 ;
        RECT 40.565 140.585 40.735 141.385 ;
        RECT 40.905 140.365 41.235 141.215 ;
        RECT 41.405 140.585 41.575 141.385 ;
        RECT 41.745 140.365 42.075 141.215 ;
        RECT 42.245 140.585 42.415 141.385 ;
        RECT 42.585 140.365 42.915 141.215 ;
        RECT 43.085 140.585 43.255 141.385 ;
        RECT 43.425 140.365 43.755 141.215 ;
        RECT 43.925 140.585 44.095 141.385 ;
        RECT 44.265 140.365 44.595 141.215 ;
        RECT 44.765 140.585 44.935 141.385 ;
        RECT 45.105 140.365 45.435 141.215 ;
        RECT 45.605 140.535 45.775 141.385 ;
        RECT 45.945 140.365 46.275 141.215 ;
        RECT 46.445 140.535 46.615 141.385 ;
        RECT 46.785 140.365 47.115 141.215 ;
        RECT 47.670 141.045 47.925 141.075 ;
        RECT 47.585 140.875 47.925 141.045 ;
        RECT 36.255 140.195 42.915 140.365 ;
        RECT 43.085 140.195 45.435 140.365 ;
        RECT 45.605 140.195 47.115 140.365 ;
        RECT 47.670 140.405 47.925 140.875 ;
        RECT 48.105 140.585 48.390 141.385 ;
        RECT 48.570 140.665 48.900 141.175 ;
        RECT 36.255 139.655 36.530 140.195 ;
        RECT 43.085 140.025 43.260 140.195 ;
        RECT 45.605 140.025 45.775 140.195 ;
        RECT 36.700 139.825 43.260 140.025 ;
        RECT 43.465 139.825 45.775 140.025 ;
        RECT 45.945 139.825 47.120 140.025 ;
        RECT 43.085 139.655 43.260 139.825 ;
        RECT 45.605 139.655 45.775 139.825 ;
        RECT 34.880 138.835 35.155 139.315 ;
        RECT 35.325 139.005 35.625 139.335 ;
        RECT 35.795 138.835 36.085 139.560 ;
        RECT 36.255 139.485 42.915 139.655 ;
        RECT 43.085 139.485 45.435 139.655 ;
        RECT 45.605 139.485 47.115 139.655 ;
        RECT 36.365 138.835 36.535 139.315 ;
        RECT 36.705 139.010 37.035 139.485 ;
        RECT 37.205 138.835 37.375 139.315 ;
        RECT 37.545 139.010 37.875 139.485 ;
        RECT 38.045 138.835 38.215 139.315 ;
        RECT 38.385 139.010 38.715 139.485 ;
        RECT 38.885 138.835 39.055 139.315 ;
        RECT 39.225 139.010 39.555 139.485 ;
        RECT 39.725 138.835 39.895 139.315 ;
        RECT 40.065 139.010 40.395 139.485 ;
        RECT 40.565 138.835 40.735 139.315 ;
        RECT 40.905 139.010 41.235 139.485 ;
        RECT 40.985 139.005 41.155 139.010 ;
        RECT 41.405 138.835 41.575 139.315 ;
        RECT 41.745 139.010 42.075 139.485 ;
        RECT 41.825 139.005 41.995 139.010 ;
        RECT 42.245 138.835 42.415 139.315 ;
        RECT 42.585 139.010 42.915 139.485 ;
        RECT 42.665 139.005 42.915 139.010 ;
        RECT 43.085 138.835 43.255 139.315 ;
        RECT 43.425 139.010 43.755 139.485 ;
        RECT 43.925 138.835 44.095 139.315 ;
        RECT 44.265 139.010 44.595 139.485 ;
        RECT 44.765 138.835 44.935 139.315 ;
        RECT 45.105 139.010 45.435 139.485 ;
        RECT 45.605 138.835 45.775 139.315 ;
        RECT 45.945 139.010 46.275 139.485 ;
        RECT 46.445 138.835 46.615 139.315 ;
        RECT 46.785 139.010 47.115 139.485 ;
        RECT 47.670 139.545 47.850 140.405 ;
        RECT 48.570 140.075 48.820 140.665 ;
        RECT 49.170 140.515 49.340 141.125 ;
        RECT 49.510 140.695 49.840 141.385 ;
        RECT 50.070 140.835 50.310 141.125 ;
        RECT 50.510 141.005 50.930 141.385 ;
        RECT 51.110 140.915 51.740 141.165 ;
        RECT 52.210 141.005 52.540 141.385 ;
        RECT 51.110 140.835 51.280 140.915 ;
        RECT 52.710 140.835 52.880 141.125 ;
        RECT 53.060 141.005 53.440 141.385 ;
        RECT 53.680 141.000 54.510 141.170 ;
        RECT 50.070 140.665 51.280 140.835 ;
        RECT 48.020 139.745 48.820 140.075 ;
        RECT 47.670 139.015 47.925 139.545 ;
        RECT 48.105 138.835 48.390 139.295 ;
        RECT 48.570 139.095 48.820 139.745 ;
        RECT 49.020 140.495 49.340 140.515 ;
        RECT 49.020 140.325 50.940 140.495 ;
        RECT 49.020 139.430 49.210 140.325 ;
        RECT 51.110 140.155 51.280 140.665 ;
        RECT 51.450 140.405 51.970 140.715 ;
        RECT 49.380 139.985 51.280 140.155 ;
        RECT 49.380 139.925 49.710 139.985 ;
        RECT 49.860 139.755 50.190 139.815 ;
        RECT 49.530 139.485 50.190 139.755 ;
        RECT 49.020 139.100 49.340 139.430 ;
        RECT 49.520 138.835 50.180 139.315 ;
        RECT 50.380 139.225 50.550 139.985 ;
        RECT 51.450 139.815 51.630 140.225 ;
        RECT 50.720 139.645 51.050 139.765 ;
        RECT 51.800 139.645 51.970 140.405 ;
        RECT 50.720 139.475 51.970 139.645 ;
        RECT 52.140 140.585 53.510 140.835 ;
        RECT 52.140 139.815 52.330 140.585 ;
        RECT 53.260 140.325 53.510 140.585 ;
        RECT 52.500 140.155 52.750 140.315 ;
        RECT 53.680 140.155 53.850 141.000 ;
        RECT 54.745 140.715 54.915 141.215 ;
        RECT 55.085 140.885 55.415 141.385 ;
        RECT 54.020 140.325 54.520 140.705 ;
        RECT 54.745 140.545 55.440 140.715 ;
        RECT 52.500 139.985 53.850 140.155 ;
        RECT 53.430 139.945 53.850 139.985 ;
        RECT 52.140 139.475 52.560 139.815 ;
        RECT 52.850 139.485 53.260 139.815 ;
        RECT 50.380 139.055 51.230 139.225 ;
        RECT 51.790 138.835 52.110 139.295 ;
        RECT 52.310 139.045 52.560 139.475 ;
        RECT 52.850 138.835 53.260 139.275 ;
        RECT 53.430 139.215 53.600 139.945 ;
        RECT 53.770 139.395 54.120 139.765 ;
        RECT 54.300 139.455 54.520 140.325 ;
        RECT 54.690 139.755 55.100 140.375 ;
        RECT 55.270 139.575 55.440 140.545 ;
        RECT 54.745 139.385 55.440 139.575 ;
        RECT 53.430 139.015 54.445 139.215 ;
        RECT 54.745 139.055 54.915 139.385 ;
        RECT 55.085 138.835 55.415 139.215 ;
        RECT 55.630 139.095 55.855 141.215 ;
        RECT 56.025 140.885 56.355 141.385 ;
        RECT 56.525 140.715 56.695 141.215 ;
        RECT 56.960 140.875 58.615 141.165 ;
        RECT 56.030 140.545 56.695 140.715 ;
        RECT 56.030 139.555 56.260 140.545 ;
        RECT 56.960 140.535 58.550 140.705 ;
        RECT 58.785 140.585 59.065 141.385 ;
        RECT 56.430 139.725 56.780 140.375 ;
        RECT 56.960 140.245 57.280 140.535 ;
        RECT 58.380 140.415 58.550 140.535 ;
        RECT 57.475 140.195 58.190 140.365 ;
        RECT 58.380 140.245 59.105 140.415 ;
        RECT 59.275 140.245 59.545 141.215 ;
        RECT 56.030 139.385 56.695 139.555 ;
        RECT 56.960 139.505 57.310 140.075 ;
        RECT 57.480 139.745 58.190 140.195 ;
        RECT 58.935 140.075 59.105 140.245 ;
        RECT 58.360 139.745 58.765 140.075 ;
        RECT 58.935 139.745 59.205 140.075 ;
        RECT 58.935 139.575 59.105 139.745 ;
        RECT 56.025 138.835 56.355 139.215 ;
        RECT 56.525 139.095 56.695 139.385 ;
        RECT 57.495 139.405 59.105 139.575 ;
        RECT 59.375 139.510 59.545 140.245 ;
        RECT 59.715 140.295 61.385 141.385 ;
        RECT 59.715 139.775 60.465 140.295 ;
        RECT 61.555 140.220 61.845 141.385 ;
        RECT 62.975 140.245 63.205 141.385 ;
        RECT 63.375 140.235 63.705 141.215 ;
        RECT 63.875 140.245 64.085 141.385 ;
        RECT 64.320 140.960 64.655 141.385 ;
        RECT 64.825 140.780 65.010 141.185 ;
        RECT 64.345 140.605 65.010 140.780 ;
        RECT 65.215 140.605 65.545 141.385 ;
        RECT 60.635 139.605 61.385 140.125 ;
        RECT 62.955 139.825 63.285 140.075 ;
        RECT 56.965 138.835 57.295 139.335 ;
        RECT 57.495 139.055 57.665 139.405 ;
        RECT 57.865 138.835 58.195 139.235 ;
        RECT 58.365 139.055 58.535 139.405 ;
        RECT 58.705 138.835 59.085 139.235 ;
        RECT 59.275 139.165 59.545 139.510 ;
        RECT 59.715 138.835 61.385 139.605 ;
        RECT 61.555 138.835 61.845 139.560 ;
        RECT 62.975 138.835 63.205 139.655 ;
        RECT 63.455 139.635 63.705 140.235 ;
        RECT 63.375 139.005 63.705 139.635 ;
        RECT 63.875 138.835 64.085 139.655 ;
        RECT 64.345 139.575 64.685 140.605 ;
        RECT 65.715 140.415 65.985 141.185 ;
        RECT 64.855 140.245 65.985 140.415 ;
        RECT 64.855 139.745 65.105 140.245 ;
        RECT 64.345 139.405 65.030 139.575 ;
        RECT 65.285 139.495 65.645 140.075 ;
        RECT 64.320 138.835 64.655 139.235 ;
        RECT 64.825 139.005 65.030 139.405 ;
        RECT 65.815 139.335 65.985 140.245 ;
        RECT 65.240 138.835 65.515 139.315 ;
        RECT 65.725 139.005 65.985 139.335 ;
        RECT 66.155 140.665 66.615 141.215 ;
        RECT 66.805 140.665 67.135 141.385 ;
        RECT 66.155 139.295 66.405 140.665 ;
        RECT 67.335 140.495 67.635 141.045 ;
        RECT 67.805 140.715 68.085 141.385 ;
        RECT 66.695 140.325 67.635 140.495 ;
        RECT 66.695 140.075 66.865 140.325 ;
        RECT 68.005 140.075 68.270 140.435 ;
        RECT 66.575 139.745 66.865 140.075 ;
        RECT 67.035 139.825 67.375 140.075 ;
        RECT 67.595 139.825 68.270 140.075 ;
        RECT 68.455 140.415 68.765 141.215 ;
        RECT 68.935 140.585 69.245 141.385 ;
        RECT 69.415 140.755 69.675 141.215 ;
        RECT 69.845 140.925 70.100 141.385 ;
        RECT 70.275 140.755 70.535 141.215 ;
        RECT 69.415 140.585 70.535 140.755 ;
        RECT 68.455 140.245 69.485 140.415 ;
        RECT 66.695 139.655 66.865 139.745 ;
        RECT 66.695 139.465 68.085 139.655 ;
        RECT 66.155 139.005 66.715 139.295 ;
        RECT 66.885 138.835 67.135 139.295 ;
        RECT 67.755 139.105 68.085 139.465 ;
        RECT 68.455 139.335 68.625 140.245 ;
        RECT 68.795 139.505 69.145 140.075 ;
        RECT 69.315 139.995 69.485 140.245 ;
        RECT 70.275 140.335 70.535 140.585 ;
        RECT 70.705 140.515 70.990 141.385 ;
        RECT 72.225 140.640 72.495 141.385 ;
        RECT 73.125 141.380 79.400 141.385 ;
        RECT 72.665 140.470 72.955 141.210 ;
        RECT 73.125 140.655 73.380 141.380 ;
        RECT 73.565 140.485 73.825 141.210 ;
        RECT 73.995 140.655 74.240 141.380 ;
        RECT 74.425 140.485 74.685 141.210 ;
        RECT 74.855 140.655 75.100 141.380 ;
        RECT 75.285 140.485 75.545 141.210 ;
        RECT 75.715 140.655 75.960 141.380 ;
        RECT 76.130 140.485 76.390 141.210 ;
        RECT 76.560 140.655 76.820 141.380 ;
        RECT 76.990 140.485 77.250 141.210 ;
        RECT 77.420 140.655 77.680 141.380 ;
        RECT 77.850 140.485 78.110 141.210 ;
        RECT 78.280 140.655 78.540 141.380 ;
        RECT 78.710 140.485 78.970 141.210 ;
        RECT 79.140 140.585 79.400 141.380 ;
        RECT 73.565 140.470 78.970 140.485 ;
        RECT 72.225 140.365 78.970 140.470 ;
        RECT 70.275 140.165 71.030 140.335 ;
        RECT 72.195 140.245 78.970 140.365 ;
        RECT 72.195 140.195 73.390 140.245 ;
        RECT 69.315 139.825 70.455 139.995 ;
        RECT 70.625 139.655 71.030 140.165 ;
        RECT 69.380 139.485 71.030 139.655 ;
        RECT 72.225 139.655 73.390 140.195 ;
        RECT 79.570 140.075 79.820 141.210 ;
        RECT 80.000 140.575 80.260 141.385 ;
        RECT 80.435 140.075 80.680 141.215 ;
        RECT 80.860 140.575 81.155 141.385 ;
        RECT 81.335 140.665 81.795 141.215 ;
        RECT 81.985 140.665 82.315 141.385 ;
        RECT 73.560 139.825 80.680 140.075 ;
        RECT 72.225 139.485 78.970 139.655 ;
        RECT 68.455 139.005 68.755 139.335 ;
        RECT 68.925 138.835 69.200 139.315 ;
        RECT 69.380 139.095 69.675 139.485 ;
        RECT 69.845 138.835 70.100 139.315 ;
        RECT 70.275 139.095 70.535 139.485 ;
        RECT 70.705 138.835 70.985 139.315 ;
        RECT 72.225 138.835 72.525 139.315 ;
        RECT 72.695 139.030 72.955 139.485 ;
        RECT 73.125 138.835 73.385 139.315 ;
        RECT 73.565 139.030 73.825 139.485 ;
        RECT 73.995 138.835 74.245 139.315 ;
        RECT 74.425 139.030 74.685 139.485 ;
        RECT 74.855 138.835 75.105 139.315 ;
        RECT 75.285 139.030 75.545 139.485 ;
        RECT 75.715 138.835 75.960 139.315 ;
        RECT 76.130 139.030 76.405 139.485 ;
        RECT 76.575 138.835 76.820 139.315 ;
        RECT 76.990 139.030 77.250 139.485 ;
        RECT 77.420 138.835 77.680 139.315 ;
        RECT 77.850 139.030 78.110 139.485 ;
        RECT 78.280 138.835 78.540 139.315 ;
        RECT 78.710 139.030 78.970 139.485 ;
        RECT 79.140 138.835 79.400 139.395 ;
        RECT 79.570 139.015 79.820 139.825 ;
        RECT 80.000 138.835 80.260 139.360 ;
        RECT 80.430 139.015 80.680 139.825 ;
        RECT 80.850 139.515 81.165 140.075 ;
        RECT 80.860 138.835 81.165 139.345 ;
        RECT 81.335 139.295 81.585 140.665 ;
        RECT 82.515 140.495 82.815 141.045 ;
        RECT 82.985 140.715 83.265 141.385 ;
        RECT 81.875 140.325 82.815 140.495 ;
        RECT 81.875 140.075 82.045 140.325 ;
        RECT 83.185 140.075 83.450 140.435 ;
        RECT 83.695 140.245 83.905 141.385 ;
        RECT 81.755 139.745 82.045 140.075 ;
        RECT 82.215 139.825 82.555 140.075 ;
        RECT 82.775 139.825 83.450 140.075 ;
        RECT 84.075 140.235 84.405 141.215 ;
        RECT 84.575 140.245 84.805 141.385 ;
        RECT 85.215 140.715 85.495 141.385 ;
        RECT 85.665 140.495 85.965 141.045 ;
        RECT 86.165 140.665 86.495 141.385 ;
        RECT 86.685 140.665 87.145 141.215 ;
        RECT 81.875 139.655 82.045 139.745 ;
        RECT 81.875 139.465 83.265 139.655 ;
        RECT 81.335 139.005 81.895 139.295 ;
        RECT 82.065 138.835 82.315 139.295 ;
        RECT 82.935 139.105 83.265 139.465 ;
        RECT 83.695 138.835 83.905 139.655 ;
        RECT 84.075 139.635 84.325 140.235 ;
        RECT 85.030 140.075 85.295 140.435 ;
        RECT 85.665 140.325 86.605 140.495 ;
        RECT 86.435 140.075 86.605 140.325 ;
        RECT 84.495 139.825 84.825 140.075 ;
        RECT 85.030 139.825 85.705 140.075 ;
        RECT 85.925 139.825 86.265 140.075 ;
        RECT 86.435 139.745 86.725 140.075 ;
        RECT 86.435 139.655 86.605 139.745 ;
        RECT 84.075 139.005 84.405 139.635 ;
        RECT 84.575 138.835 84.805 139.655 ;
        RECT 85.215 139.465 86.605 139.655 ;
        RECT 85.215 139.105 85.545 139.465 ;
        RECT 86.895 139.295 87.145 140.665 ;
        RECT 87.315 140.220 87.605 141.385 ;
        RECT 87.785 140.575 88.080 141.385 ;
        RECT 88.260 140.075 88.505 141.215 ;
        RECT 88.680 140.575 88.940 141.385 ;
        RECT 89.540 141.380 95.815 141.385 ;
        RECT 89.120 140.075 89.370 141.210 ;
        RECT 89.540 140.585 89.800 141.380 ;
        RECT 89.970 140.485 90.230 141.210 ;
        RECT 90.400 140.655 90.660 141.380 ;
        RECT 90.830 140.485 91.090 141.210 ;
        RECT 91.260 140.655 91.520 141.380 ;
        RECT 91.690 140.485 91.950 141.210 ;
        RECT 92.120 140.655 92.380 141.380 ;
        RECT 92.550 140.485 92.810 141.210 ;
        RECT 92.980 140.655 93.225 141.380 ;
        RECT 93.395 140.485 93.655 141.210 ;
        RECT 93.840 140.655 94.085 141.380 ;
        RECT 94.255 140.485 94.515 141.210 ;
        RECT 94.700 140.655 94.945 141.380 ;
        RECT 95.115 140.485 95.375 141.210 ;
        RECT 95.560 140.655 95.815 141.380 ;
        RECT 89.970 140.470 95.375 140.485 ;
        RECT 95.985 140.470 96.275 141.210 ;
        RECT 96.445 140.640 96.715 141.385 ;
        RECT 96.975 140.665 97.435 141.215 ;
        RECT 97.625 140.665 97.955 141.385 ;
        RECT 89.970 140.245 96.715 140.470 ;
        RECT 86.165 138.835 86.415 139.295 ;
        RECT 86.585 139.005 87.145 139.295 ;
        RECT 87.315 138.835 87.605 139.560 ;
        RECT 87.775 139.515 88.090 140.075 ;
        RECT 88.260 139.825 95.380 140.075 ;
        RECT 87.775 138.835 88.080 139.345 ;
        RECT 88.260 139.015 88.510 139.825 ;
        RECT 88.680 138.835 88.940 139.360 ;
        RECT 89.120 139.015 89.370 139.825 ;
        RECT 95.550 139.655 96.715 140.245 ;
        RECT 89.970 139.485 96.715 139.655 ;
        RECT 89.540 138.835 89.800 139.395 ;
        RECT 89.970 139.030 90.230 139.485 ;
        RECT 90.400 138.835 90.660 139.315 ;
        RECT 90.830 139.030 91.090 139.485 ;
        RECT 91.260 138.835 91.520 139.315 ;
        RECT 91.690 139.030 91.950 139.485 ;
        RECT 92.120 138.835 92.365 139.315 ;
        RECT 92.535 139.030 92.810 139.485 ;
        RECT 92.980 138.835 93.225 139.315 ;
        RECT 93.395 139.030 93.655 139.485 ;
        RECT 93.835 138.835 94.085 139.315 ;
        RECT 94.255 139.030 94.515 139.485 ;
        RECT 94.695 138.835 94.945 139.315 ;
        RECT 95.115 139.030 95.375 139.485 ;
        RECT 95.555 138.835 95.815 139.315 ;
        RECT 95.985 139.030 96.245 139.485 ;
        RECT 96.415 138.835 96.715 139.315 ;
        RECT 96.975 139.295 97.225 140.665 ;
        RECT 98.155 140.495 98.455 141.045 ;
        RECT 98.625 140.715 98.905 141.385 ;
        RECT 97.515 140.325 98.455 140.495 ;
        RECT 97.515 140.075 97.685 140.325 ;
        RECT 98.825 140.075 99.090 140.435 ;
        RECT 97.395 139.745 97.685 140.075 ;
        RECT 97.855 139.825 98.195 140.075 ;
        RECT 98.415 139.825 99.090 140.075 ;
        RECT 99.275 140.295 100.485 141.385 ;
        RECT 101.030 140.405 101.285 141.075 ;
        RECT 101.465 140.585 101.750 141.385 ;
        RECT 101.930 140.665 102.260 141.175 ;
        RECT 99.275 139.755 99.795 140.295 ;
        RECT 97.515 139.655 97.685 139.745 ;
        RECT 97.515 139.465 98.905 139.655 ;
        RECT 99.965 139.585 100.485 140.125 ;
        RECT 101.030 139.685 101.210 140.405 ;
        RECT 101.930 140.075 102.180 140.665 ;
        RECT 102.530 140.515 102.700 141.125 ;
        RECT 102.870 140.695 103.200 141.385 ;
        RECT 103.430 140.835 103.670 141.125 ;
        RECT 103.870 141.005 104.290 141.385 ;
        RECT 104.470 140.915 105.100 141.165 ;
        RECT 105.570 141.005 105.900 141.385 ;
        RECT 104.470 140.835 104.640 140.915 ;
        RECT 106.070 140.835 106.240 141.125 ;
        RECT 106.420 141.005 106.800 141.385 ;
        RECT 107.040 141.000 107.870 141.170 ;
        RECT 103.430 140.665 104.640 140.835 ;
        RECT 101.380 139.745 102.180 140.075 ;
        RECT 96.975 139.005 97.535 139.295 ;
        RECT 97.705 138.835 97.955 139.295 ;
        RECT 98.575 139.105 98.905 139.465 ;
        RECT 99.275 138.835 100.485 139.585 ;
        RECT 100.945 139.545 101.210 139.685 ;
        RECT 100.945 139.515 101.285 139.545 ;
        RECT 101.030 139.015 101.285 139.515 ;
        RECT 101.465 138.835 101.750 139.295 ;
        RECT 101.930 139.095 102.180 139.745 ;
        RECT 102.380 140.495 102.700 140.515 ;
        RECT 102.380 140.325 104.300 140.495 ;
        RECT 102.380 139.430 102.570 140.325 ;
        RECT 104.470 140.155 104.640 140.665 ;
        RECT 104.810 140.405 105.330 140.715 ;
        RECT 102.740 139.985 104.640 140.155 ;
        RECT 102.740 139.925 103.070 139.985 ;
        RECT 103.220 139.755 103.550 139.815 ;
        RECT 102.890 139.485 103.550 139.755 ;
        RECT 102.380 139.100 102.700 139.430 ;
        RECT 102.880 138.835 103.540 139.315 ;
        RECT 103.740 139.225 103.910 139.985 ;
        RECT 104.810 139.815 104.990 140.225 ;
        RECT 104.080 139.645 104.410 139.765 ;
        RECT 105.160 139.645 105.330 140.405 ;
        RECT 104.080 139.475 105.330 139.645 ;
        RECT 105.500 140.585 106.870 140.835 ;
        RECT 105.500 139.815 105.690 140.585 ;
        RECT 106.620 140.325 106.870 140.585 ;
        RECT 105.860 140.155 106.110 140.315 ;
        RECT 107.040 140.155 107.210 141.000 ;
        RECT 108.105 140.715 108.275 141.215 ;
        RECT 108.445 140.885 108.775 141.385 ;
        RECT 107.380 140.325 107.880 140.705 ;
        RECT 108.105 140.545 108.800 140.715 ;
        RECT 105.860 139.985 107.210 140.155 ;
        RECT 106.790 139.945 107.210 139.985 ;
        RECT 105.500 139.475 105.920 139.815 ;
        RECT 106.210 139.485 106.620 139.815 ;
        RECT 103.740 139.055 104.590 139.225 ;
        RECT 105.150 138.835 105.470 139.295 ;
        RECT 105.670 139.045 105.920 139.475 ;
        RECT 106.210 138.835 106.620 139.275 ;
        RECT 106.790 139.215 106.960 139.945 ;
        RECT 107.130 139.395 107.480 139.765 ;
        RECT 107.660 139.455 107.880 140.325 ;
        RECT 108.050 139.755 108.460 140.375 ;
        RECT 108.630 139.575 108.800 140.545 ;
        RECT 108.105 139.385 108.800 139.575 ;
        RECT 106.790 139.015 107.805 139.215 ;
        RECT 108.105 139.055 108.275 139.385 ;
        RECT 108.445 138.835 108.775 139.215 ;
        RECT 108.990 139.095 109.215 141.215 ;
        RECT 109.385 140.885 109.715 141.385 ;
        RECT 109.885 140.715 110.055 141.215 ;
        RECT 109.390 140.545 110.055 140.715 ;
        RECT 109.390 139.555 109.620 140.545 ;
        RECT 109.790 139.725 110.140 140.375 ;
        RECT 110.315 140.295 111.985 141.385 ;
        RECT 112.155 140.295 113.365 141.385 ;
        RECT 110.315 139.775 111.065 140.295 ;
        RECT 111.235 139.605 111.985 140.125 ;
        RECT 112.155 139.755 112.675 140.295 ;
        RECT 109.390 139.385 110.055 139.555 ;
        RECT 109.385 138.835 109.715 139.215 ;
        RECT 109.885 139.095 110.055 139.385 ;
        RECT 110.315 138.835 111.985 139.605 ;
        RECT 112.845 139.585 113.365 140.125 ;
        RECT 112.155 138.835 113.365 139.585 ;
        RECT 22.830 138.665 113.450 138.835 ;
        RECT 22.915 137.915 24.125 138.665 ;
        RECT 24.845 138.115 25.015 138.405 ;
        RECT 25.185 138.285 25.515 138.665 ;
        RECT 24.845 137.945 25.510 138.115 ;
        RECT 22.915 137.375 23.435 137.915 ;
        RECT 23.605 137.205 24.125 137.745 ;
        RECT 22.915 136.115 24.125 137.205 ;
        RECT 24.760 137.125 25.110 137.775 ;
        RECT 25.280 136.955 25.510 137.945 ;
        RECT 24.845 136.785 25.510 136.955 ;
        RECT 24.845 136.285 25.015 136.785 ;
        RECT 25.185 136.115 25.515 136.615 ;
        RECT 25.685 136.285 25.910 138.405 ;
        RECT 26.125 138.285 26.455 138.665 ;
        RECT 26.625 138.115 26.795 138.445 ;
        RECT 27.095 138.285 28.110 138.485 ;
        RECT 26.100 137.925 26.795 138.115 ;
        RECT 26.100 136.955 26.270 137.925 ;
        RECT 26.440 137.125 26.850 137.745 ;
        RECT 27.020 137.175 27.240 138.045 ;
        RECT 27.420 137.735 27.770 138.105 ;
        RECT 27.940 137.555 28.110 138.285 ;
        RECT 28.280 138.225 28.690 138.665 ;
        RECT 28.980 138.025 29.230 138.455 ;
        RECT 29.430 138.205 29.750 138.665 ;
        RECT 30.310 138.275 31.160 138.445 ;
        RECT 28.280 137.685 28.690 138.015 ;
        RECT 28.980 137.685 29.400 138.025 ;
        RECT 27.690 137.515 28.110 137.555 ;
        RECT 27.690 137.345 29.040 137.515 ;
        RECT 26.100 136.785 26.795 136.955 ;
        RECT 27.020 136.795 27.520 137.175 ;
        RECT 26.125 136.115 26.455 136.615 ;
        RECT 26.625 136.285 26.795 136.785 ;
        RECT 27.690 136.500 27.860 137.345 ;
        RECT 28.790 137.185 29.040 137.345 ;
        RECT 28.030 136.915 28.280 137.175 ;
        RECT 29.210 136.915 29.400 137.685 ;
        RECT 28.030 136.665 29.400 136.915 ;
        RECT 29.570 137.855 30.820 138.025 ;
        RECT 29.570 137.095 29.740 137.855 ;
        RECT 30.490 137.735 30.820 137.855 ;
        RECT 29.910 137.275 30.090 137.685 ;
        RECT 30.990 137.515 31.160 138.275 ;
        RECT 31.360 138.185 32.020 138.665 ;
        RECT 32.200 138.070 32.520 138.400 ;
        RECT 31.350 137.745 32.010 138.015 ;
        RECT 31.350 137.685 31.680 137.745 ;
        RECT 31.830 137.515 32.160 137.575 ;
        RECT 30.260 137.345 32.160 137.515 ;
        RECT 29.570 136.785 30.090 137.095 ;
        RECT 30.260 136.835 30.430 137.345 ;
        RECT 32.330 137.175 32.520 138.070 ;
        RECT 30.600 137.005 32.520 137.175 ;
        RECT 32.200 136.985 32.520 137.005 ;
        RECT 32.720 137.755 32.970 138.405 ;
        RECT 33.150 138.205 33.435 138.665 ;
        RECT 33.615 138.325 33.870 138.485 ;
        RECT 33.615 138.155 33.955 138.325 ;
        RECT 33.615 137.955 33.870 138.155 ;
        RECT 32.720 137.425 33.520 137.755 ;
        RECT 30.260 136.665 31.470 136.835 ;
        RECT 27.030 136.330 27.860 136.500 ;
        RECT 28.100 136.115 28.480 136.495 ;
        RECT 28.660 136.375 28.830 136.665 ;
        RECT 30.260 136.585 30.430 136.665 ;
        RECT 29.000 136.115 29.330 136.495 ;
        RECT 29.800 136.335 30.430 136.585 ;
        RECT 30.610 136.115 31.030 136.495 ;
        RECT 31.230 136.375 31.470 136.665 ;
        RECT 31.700 136.115 32.030 136.805 ;
        RECT 32.200 136.375 32.370 136.985 ;
        RECT 32.720 136.835 32.970 137.425 ;
        RECT 33.690 137.095 33.870 137.955 ;
        RECT 34.505 138.115 34.675 138.495 ;
        RECT 34.855 138.285 35.185 138.665 ;
        RECT 34.505 137.945 35.170 138.115 ;
        RECT 35.365 137.990 35.625 138.495 ;
        RECT 35.885 138.185 36.185 138.665 ;
        RECT 36.355 138.015 36.615 138.470 ;
        RECT 36.785 138.185 37.045 138.665 ;
        RECT 37.225 138.015 37.485 138.470 ;
        RECT 37.655 138.185 37.905 138.665 ;
        RECT 38.085 138.015 38.345 138.470 ;
        RECT 38.515 138.185 38.765 138.665 ;
        RECT 38.945 138.015 39.205 138.470 ;
        RECT 39.375 138.185 39.620 138.665 ;
        RECT 39.790 138.015 40.065 138.470 ;
        RECT 40.235 138.185 40.480 138.665 ;
        RECT 40.650 138.015 40.910 138.470 ;
        RECT 41.080 138.185 41.340 138.665 ;
        RECT 41.510 138.015 41.770 138.470 ;
        RECT 41.940 138.185 42.200 138.665 ;
        RECT 42.370 138.015 42.630 138.470 ;
        RECT 42.800 138.105 43.060 138.665 ;
        RECT 34.435 137.395 34.765 137.765 ;
        RECT 35.000 137.690 35.170 137.945 ;
        RECT 35.000 137.360 35.285 137.690 ;
        RECT 35.000 137.215 35.170 137.360 ;
        RECT 32.640 136.325 32.970 136.835 ;
        RECT 33.150 136.115 33.435 136.915 ;
        RECT 33.615 136.425 33.870 137.095 ;
        RECT 34.505 137.045 35.170 137.215 ;
        RECT 35.455 137.190 35.625 137.990 ;
        RECT 34.505 136.285 34.675 137.045 ;
        RECT 34.855 136.115 35.185 136.875 ;
        RECT 35.355 136.285 35.625 137.190 ;
        RECT 35.885 137.845 42.630 138.015 ;
        RECT 35.885 137.255 37.050 137.845 ;
        RECT 43.230 137.675 43.480 138.485 ;
        RECT 43.660 138.140 43.920 138.665 ;
        RECT 44.090 137.675 44.340 138.485 ;
        RECT 44.520 138.155 44.825 138.665 ;
        RECT 37.220 137.425 44.340 137.675 ;
        RECT 44.510 137.425 44.825 137.985 ;
        RECT 44.995 137.865 45.335 138.495 ;
        RECT 45.505 137.865 45.755 138.665 ;
        RECT 45.945 138.015 46.275 138.495 ;
        RECT 46.445 138.205 46.670 138.665 ;
        RECT 46.840 138.015 47.170 138.495 ;
        RECT 35.885 137.030 42.630 137.255 ;
        RECT 35.885 136.115 36.155 136.860 ;
        RECT 36.325 136.290 36.615 137.030 ;
        RECT 37.225 137.015 42.630 137.030 ;
        RECT 36.785 136.120 37.040 136.845 ;
        RECT 37.225 136.290 37.485 137.015 ;
        RECT 37.655 136.120 37.900 136.845 ;
        RECT 38.085 136.290 38.345 137.015 ;
        RECT 38.515 136.120 38.760 136.845 ;
        RECT 38.945 136.290 39.205 137.015 ;
        RECT 39.375 136.120 39.620 136.845 ;
        RECT 39.790 136.290 40.050 137.015 ;
        RECT 40.220 136.120 40.480 136.845 ;
        RECT 40.650 136.290 40.910 137.015 ;
        RECT 41.080 136.120 41.340 136.845 ;
        RECT 41.510 136.290 41.770 137.015 ;
        RECT 41.940 136.120 42.200 136.845 ;
        RECT 42.370 136.290 42.630 137.015 ;
        RECT 42.800 136.120 43.060 136.915 ;
        RECT 43.230 136.290 43.480 137.425 ;
        RECT 36.785 136.115 43.060 136.120 ;
        RECT 43.660 136.115 43.920 136.925 ;
        RECT 44.095 136.285 44.340 137.425 ;
        RECT 44.995 137.255 45.170 137.865 ;
        RECT 45.945 137.845 47.170 138.015 ;
        RECT 47.800 137.885 48.300 138.495 ;
        RECT 48.675 137.940 48.965 138.665 ;
        RECT 49.135 138.155 49.440 138.665 ;
        RECT 45.340 137.505 46.035 137.675 ;
        RECT 45.865 137.255 46.035 137.505 ;
        RECT 46.210 137.475 46.630 137.675 ;
        RECT 46.800 137.475 47.130 137.675 ;
        RECT 47.300 137.475 47.630 137.675 ;
        RECT 47.800 137.255 47.970 137.885 ;
        RECT 48.155 137.425 48.505 137.675 ;
        RECT 49.135 137.425 49.450 137.985 ;
        RECT 49.620 137.675 49.870 138.485 ;
        RECT 50.040 138.140 50.300 138.665 ;
        RECT 50.480 137.675 50.730 138.485 ;
        RECT 50.900 138.105 51.160 138.665 ;
        RECT 51.330 138.015 51.590 138.470 ;
        RECT 51.760 138.185 52.020 138.665 ;
        RECT 52.190 138.015 52.450 138.470 ;
        RECT 52.620 138.185 52.880 138.665 ;
        RECT 53.050 138.015 53.310 138.470 ;
        RECT 53.480 138.185 53.725 138.665 ;
        RECT 53.895 138.015 54.170 138.470 ;
        RECT 54.340 138.185 54.585 138.665 ;
        RECT 54.755 138.015 55.015 138.470 ;
        RECT 55.195 138.185 55.445 138.665 ;
        RECT 55.615 138.015 55.875 138.470 ;
        RECT 56.055 138.185 56.305 138.665 ;
        RECT 56.475 138.015 56.735 138.470 ;
        RECT 56.915 138.185 57.175 138.665 ;
        RECT 57.345 138.015 57.605 138.470 ;
        RECT 57.775 138.185 58.075 138.665 ;
        RECT 51.330 137.845 58.075 138.015 ;
        RECT 49.620 137.425 56.740 137.675 ;
        RECT 44.520 136.115 44.815 136.925 ;
        RECT 44.995 136.285 45.335 137.255 ;
        RECT 45.505 136.115 45.675 137.255 ;
        RECT 45.865 137.085 48.300 137.255 ;
        RECT 45.945 136.115 46.195 136.915 ;
        RECT 46.840 136.285 47.170 137.085 ;
        RECT 47.470 136.115 47.800 136.915 ;
        RECT 47.970 136.285 48.300 137.085 ;
        RECT 48.675 136.115 48.965 137.280 ;
        RECT 49.145 136.115 49.440 136.925 ;
        RECT 49.620 136.285 49.865 137.425 ;
        RECT 50.040 136.115 50.300 136.925 ;
        RECT 50.480 136.290 50.730 137.425 ;
        RECT 56.910 137.255 58.075 137.845 ;
        RECT 51.330 137.030 58.075 137.255 ;
        RECT 58.795 137.865 59.135 138.495 ;
        RECT 59.305 137.865 59.555 138.665 ;
        RECT 59.745 138.015 60.075 138.495 ;
        RECT 60.245 138.205 60.470 138.665 ;
        RECT 60.640 138.015 60.970 138.495 ;
        RECT 58.795 137.255 58.970 137.865 ;
        RECT 59.745 137.845 60.970 138.015 ;
        RECT 61.600 137.885 62.100 138.495 ;
        RECT 59.140 137.505 59.835 137.675 ;
        RECT 59.665 137.255 59.835 137.505 ;
        RECT 60.010 137.475 60.430 137.675 ;
        RECT 60.600 137.475 60.930 137.675 ;
        RECT 61.100 137.475 61.430 137.675 ;
        RECT 61.600 137.255 61.770 137.885 ;
        RECT 62.750 137.855 62.995 138.460 ;
        RECT 63.215 138.130 63.725 138.665 ;
        RECT 62.475 137.685 63.705 137.855 ;
        RECT 61.955 137.425 62.305 137.675 ;
        RECT 51.330 137.015 56.735 137.030 ;
        RECT 50.900 136.120 51.160 136.915 ;
        RECT 51.330 136.290 51.590 137.015 ;
        RECT 51.760 136.120 52.020 136.845 ;
        RECT 52.190 136.290 52.450 137.015 ;
        RECT 52.620 136.120 52.880 136.845 ;
        RECT 53.050 136.290 53.310 137.015 ;
        RECT 53.480 136.120 53.740 136.845 ;
        RECT 53.910 136.290 54.170 137.015 ;
        RECT 54.340 136.120 54.585 136.845 ;
        RECT 54.755 136.290 55.015 137.015 ;
        RECT 55.200 136.120 55.445 136.845 ;
        RECT 55.615 136.290 55.875 137.015 ;
        RECT 56.060 136.120 56.305 136.845 ;
        RECT 56.475 136.290 56.735 137.015 ;
        RECT 56.920 136.120 57.175 136.845 ;
        RECT 57.345 136.290 57.635 137.030 ;
        RECT 50.900 136.115 57.175 136.120 ;
        RECT 57.805 136.115 58.075 136.860 ;
        RECT 58.795 136.285 59.135 137.255 ;
        RECT 59.305 136.115 59.475 137.255 ;
        RECT 59.665 137.085 62.100 137.255 ;
        RECT 59.745 136.115 59.995 136.915 ;
        RECT 60.640 136.285 60.970 137.085 ;
        RECT 61.270 136.115 61.600 136.915 ;
        RECT 61.770 136.285 62.100 137.085 ;
        RECT 62.475 136.875 62.815 137.685 ;
        RECT 62.985 137.120 63.735 137.310 ;
        RECT 62.475 136.465 62.990 136.875 ;
        RECT 63.225 136.115 63.395 136.875 ;
        RECT 63.565 136.455 63.735 137.120 ;
        RECT 63.905 137.135 64.095 138.495 ;
        RECT 64.265 138.325 64.540 138.495 ;
        RECT 64.265 138.155 64.545 138.325 ;
        RECT 64.265 137.335 64.540 138.155 ;
        RECT 64.730 138.130 65.260 138.495 ;
        RECT 65.685 138.265 66.015 138.665 ;
        RECT 65.085 138.095 65.260 138.130 ;
        RECT 64.745 137.135 64.915 137.935 ;
        RECT 63.905 136.965 64.915 137.135 ;
        RECT 65.085 137.925 66.015 138.095 ;
        RECT 66.185 137.925 66.440 138.495 ;
        RECT 65.085 136.795 65.255 137.925 ;
        RECT 65.845 137.755 66.015 137.925 ;
        RECT 64.130 136.625 65.255 136.795 ;
        RECT 65.425 137.425 65.620 137.755 ;
        RECT 65.845 137.425 66.100 137.755 ;
        RECT 65.425 136.455 65.595 137.425 ;
        RECT 66.270 137.255 66.440 137.925 ;
        RECT 63.565 136.285 65.595 136.455 ;
        RECT 65.765 136.115 65.935 137.255 ;
        RECT 66.105 136.285 66.440 137.255 ;
        RECT 67.075 138.205 67.635 138.495 ;
        RECT 67.805 138.205 68.055 138.665 ;
        RECT 67.075 136.835 67.325 138.205 ;
        RECT 68.675 138.035 69.005 138.395 ;
        RECT 67.615 137.845 69.005 138.035 ;
        RECT 69.575 138.035 69.905 138.395 ;
        RECT 70.525 138.205 70.775 138.665 ;
        RECT 70.945 138.205 71.505 138.495 ;
        RECT 69.575 137.845 70.965 138.035 ;
        RECT 67.615 137.755 67.785 137.845 ;
        RECT 67.495 137.425 67.785 137.755 ;
        RECT 70.795 137.755 70.965 137.845 ;
        RECT 67.955 137.425 68.295 137.675 ;
        RECT 68.515 137.425 69.190 137.675 ;
        RECT 67.615 137.175 67.785 137.425 ;
        RECT 67.615 137.005 68.555 137.175 ;
        RECT 68.925 137.065 69.190 137.425 ;
        RECT 69.390 137.425 70.065 137.675 ;
        RECT 70.285 137.425 70.625 137.675 ;
        RECT 70.795 137.425 71.085 137.755 ;
        RECT 69.390 137.065 69.655 137.425 ;
        RECT 70.795 137.175 70.965 137.425 ;
        RECT 67.075 136.285 67.535 136.835 ;
        RECT 67.725 136.115 68.055 136.835 ;
        RECT 68.255 136.455 68.555 137.005 ;
        RECT 70.025 137.005 70.965 137.175 ;
        RECT 68.725 136.115 69.005 136.785 ;
        RECT 69.575 136.115 69.855 136.785 ;
        RECT 70.025 136.455 70.325 137.005 ;
        RECT 71.255 136.835 71.505 138.205 ;
        RECT 70.525 136.115 70.855 136.835 ;
        RECT 71.045 136.285 71.505 136.835 ;
        RECT 71.675 137.990 71.945 138.335 ;
        RECT 72.135 138.265 72.515 138.665 ;
        RECT 72.685 138.095 72.855 138.445 ;
        RECT 73.025 138.265 73.355 138.665 ;
        RECT 73.555 138.095 73.725 138.445 ;
        RECT 73.925 138.165 74.255 138.665 ;
        RECT 71.675 137.255 71.845 137.990 ;
        RECT 72.115 137.925 73.725 138.095 ;
        RECT 72.115 137.755 72.285 137.925 ;
        RECT 72.015 137.425 72.285 137.755 ;
        RECT 72.455 137.425 72.860 137.755 ;
        RECT 72.115 137.255 72.285 137.425 ;
        RECT 71.675 136.285 71.945 137.255 ;
        RECT 72.115 137.085 72.840 137.255 ;
        RECT 73.030 137.135 73.740 137.755 ;
        RECT 73.910 137.425 74.260 137.995 ;
        RECT 74.435 137.940 74.725 138.665 ;
        RECT 76.090 137.855 76.335 138.460 ;
        RECT 76.555 138.130 77.065 138.665 ;
        RECT 75.815 137.685 77.045 137.855 ;
        RECT 72.670 136.965 72.840 137.085 ;
        RECT 73.940 136.965 74.260 137.255 ;
        RECT 72.155 136.115 72.435 136.915 ;
        RECT 72.670 136.795 74.260 136.965 ;
        RECT 72.605 136.335 74.260 136.625 ;
        RECT 74.435 136.115 74.725 137.280 ;
        RECT 75.815 136.875 76.155 137.685 ;
        RECT 76.325 137.120 77.075 137.310 ;
        RECT 75.815 136.465 76.330 136.875 ;
        RECT 76.565 136.115 76.735 136.875 ;
        RECT 76.905 136.455 77.075 137.120 ;
        RECT 77.245 137.135 77.435 138.495 ;
        RECT 77.605 137.645 77.880 138.495 ;
        RECT 78.070 138.130 78.600 138.495 ;
        RECT 79.025 138.265 79.355 138.665 ;
        RECT 78.425 138.095 78.600 138.130 ;
        RECT 77.605 137.475 77.885 137.645 ;
        RECT 77.605 137.335 77.880 137.475 ;
        RECT 78.085 137.135 78.255 137.935 ;
        RECT 77.245 136.965 78.255 137.135 ;
        RECT 78.425 137.925 79.355 138.095 ;
        RECT 79.525 137.925 79.780 138.495 ;
        RECT 78.425 136.795 78.595 137.925 ;
        RECT 79.185 137.755 79.355 137.925 ;
        RECT 77.470 136.625 78.595 136.795 ;
        RECT 78.765 137.425 78.960 137.755 ;
        RECT 79.185 137.425 79.440 137.755 ;
        RECT 78.765 136.455 78.935 137.425 ;
        RECT 79.610 137.255 79.780 137.925 ;
        RECT 81.150 137.855 81.395 138.460 ;
        RECT 81.615 138.130 82.125 138.665 ;
        RECT 76.905 136.285 78.935 136.455 ;
        RECT 79.105 136.115 79.275 137.255 ;
        RECT 79.445 136.285 79.780 137.255 ;
        RECT 80.875 137.685 82.105 137.855 ;
        RECT 80.875 136.875 81.215 137.685 ;
        RECT 81.385 137.120 82.135 137.310 ;
        RECT 80.875 136.465 81.390 136.875 ;
        RECT 81.625 136.115 81.795 136.875 ;
        RECT 81.965 136.455 82.135 137.120 ;
        RECT 82.305 137.135 82.495 138.495 ;
        RECT 82.665 138.325 82.940 138.495 ;
        RECT 82.665 138.155 82.945 138.325 ;
        RECT 82.665 137.335 82.940 138.155 ;
        RECT 83.130 138.130 83.660 138.495 ;
        RECT 84.085 138.265 84.415 138.665 ;
        RECT 83.485 138.095 83.660 138.130 ;
        RECT 83.145 137.135 83.315 137.935 ;
        RECT 82.305 136.965 83.315 137.135 ;
        RECT 83.485 137.925 84.415 138.095 ;
        RECT 84.585 137.925 84.840 138.495 ;
        RECT 85.105 138.115 85.275 138.405 ;
        RECT 85.445 138.285 85.775 138.665 ;
        RECT 85.105 137.945 85.770 138.115 ;
        RECT 83.485 136.795 83.655 137.925 ;
        RECT 84.245 137.755 84.415 137.925 ;
        RECT 82.530 136.625 83.655 136.795 ;
        RECT 83.825 137.425 84.020 137.755 ;
        RECT 84.245 137.425 84.500 137.755 ;
        RECT 83.825 136.455 83.995 137.425 ;
        RECT 84.670 137.255 84.840 137.925 ;
        RECT 81.965 136.285 83.995 136.455 ;
        RECT 84.165 136.115 84.335 137.255 ;
        RECT 84.505 136.285 84.840 137.255 ;
        RECT 85.020 137.125 85.370 137.775 ;
        RECT 85.540 136.955 85.770 137.945 ;
        RECT 85.105 136.785 85.770 136.955 ;
        RECT 85.105 136.285 85.275 136.785 ;
        RECT 85.445 136.115 85.775 136.615 ;
        RECT 85.945 136.285 86.170 138.405 ;
        RECT 86.385 138.285 86.715 138.665 ;
        RECT 86.885 138.115 87.055 138.445 ;
        RECT 87.355 138.285 88.370 138.485 ;
        RECT 86.360 137.925 87.055 138.115 ;
        RECT 86.360 136.955 86.530 137.925 ;
        RECT 86.700 137.125 87.110 137.745 ;
        RECT 87.280 137.175 87.500 138.045 ;
        RECT 87.680 137.735 88.030 138.105 ;
        RECT 88.200 137.555 88.370 138.285 ;
        RECT 88.540 138.225 88.950 138.665 ;
        RECT 89.240 138.025 89.490 138.455 ;
        RECT 89.690 138.205 90.010 138.665 ;
        RECT 90.570 138.275 91.420 138.445 ;
        RECT 88.540 137.685 88.950 138.015 ;
        RECT 89.240 137.685 89.660 138.025 ;
        RECT 87.950 137.515 88.370 137.555 ;
        RECT 87.950 137.345 89.300 137.515 ;
        RECT 86.360 136.785 87.055 136.955 ;
        RECT 87.280 136.795 87.780 137.175 ;
        RECT 86.385 136.115 86.715 136.615 ;
        RECT 86.885 136.285 87.055 136.785 ;
        RECT 87.950 136.500 88.120 137.345 ;
        RECT 89.050 137.185 89.300 137.345 ;
        RECT 88.290 136.915 88.540 137.175 ;
        RECT 89.470 136.915 89.660 137.685 ;
        RECT 88.290 136.665 89.660 136.915 ;
        RECT 89.830 137.855 91.080 138.025 ;
        RECT 89.830 137.095 90.000 137.855 ;
        RECT 90.750 137.735 91.080 137.855 ;
        RECT 90.170 137.275 90.350 137.685 ;
        RECT 91.250 137.515 91.420 138.275 ;
        RECT 91.620 138.185 92.280 138.665 ;
        RECT 92.460 138.070 92.780 138.400 ;
        RECT 91.610 137.745 92.270 138.015 ;
        RECT 91.610 137.685 91.940 137.745 ;
        RECT 92.090 137.515 92.420 137.575 ;
        RECT 90.520 137.345 92.420 137.515 ;
        RECT 89.830 136.785 90.350 137.095 ;
        RECT 90.520 136.835 90.690 137.345 ;
        RECT 92.590 137.175 92.780 138.070 ;
        RECT 90.860 137.005 92.780 137.175 ;
        RECT 92.460 136.985 92.780 137.005 ;
        RECT 92.980 137.755 93.230 138.405 ;
        RECT 93.410 138.205 93.695 138.665 ;
        RECT 93.875 138.325 94.130 138.485 ;
        RECT 93.875 138.155 94.215 138.325 ;
        RECT 93.875 137.955 94.130 138.155 ;
        RECT 92.980 137.425 93.780 137.755 ;
        RECT 90.520 136.665 91.730 136.835 ;
        RECT 87.290 136.330 88.120 136.500 ;
        RECT 88.360 136.115 88.740 136.495 ;
        RECT 88.920 136.375 89.090 136.665 ;
        RECT 90.520 136.585 90.690 136.665 ;
        RECT 89.260 136.115 89.590 136.495 ;
        RECT 90.060 136.335 90.690 136.585 ;
        RECT 90.870 136.115 91.290 136.495 ;
        RECT 91.490 136.375 91.730 136.665 ;
        RECT 91.960 136.115 92.290 136.805 ;
        RECT 92.460 136.375 92.630 136.985 ;
        RECT 92.980 136.835 93.230 137.425 ;
        RECT 93.950 137.095 94.130 137.955 ;
        RECT 94.765 138.115 94.935 138.495 ;
        RECT 95.115 138.285 95.445 138.665 ;
        RECT 94.765 137.945 95.430 138.115 ;
        RECT 95.625 137.990 95.885 138.495 ;
        RECT 94.695 137.395 95.025 137.765 ;
        RECT 95.260 137.690 95.430 137.945 ;
        RECT 95.260 137.360 95.545 137.690 ;
        RECT 95.260 137.215 95.430 137.360 ;
        RECT 92.900 136.325 93.230 136.835 ;
        RECT 93.410 136.115 93.695 136.915 ;
        RECT 93.875 136.425 94.130 137.095 ;
        RECT 94.765 137.045 95.430 137.215 ;
        RECT 95.715 137.190 95.885 137.990 ;
        RECT 96.330 137.855 96.575 138.460 ;
        RECT 96.795 138.130 97.305 138.665 ;
        RECT 94.765 136.285 94.935 137.045 ;
        RECT 95.115 136.115 95.445 136.875 ;
        RECT 95.615 136.285 95.885 137.190 ;
        RECT 96.055 137.685 97.285 137.855 ;
        RECT 96.055 136.875 96.395 137.685 ;
        RECT 96.565 137.120 97.315 137.310 ;
        RECT 96.055 136.465 96.570 136.875 ;
        RECT 96.805 136.115 96.975 136.875 ;
        RECT 97.145 136.455 97.315 137.120 ;
        RECT 97.485 137.135 97.675 138.495 ;
        RECT 97.845 138.325 98.120 138.495 ;
        RECT 97.845 138.155 98.125 138.325 ;
        RECT 97.845 137.335 98.120 138.155 ;
        RECT 98.310 138.130 98.840 138.495 ;
        RECT 99.265 138.265 99.595 138.665 ;
        RECT 98.665 138.095 98.840 138.130 ;
        RECT 98.325 137.135 98.495 137.935 ;
        RECT 97.485 136.965 98.495 137.135 ;
        RECT 98.665 137.925 99.595 138.095 ;
        RECT 99.765 137.925 100.020 138.495 ;
        RECT 100.195 137.940 100.485 138.665 ;
        RECT 98.665 136.795 98.835 137.925 ;
        RECT 99.425 137.755 99.595 137.925 ;
        RECT 97.710 136.625 98.835 136.795 ;
        RECT 99.005 137.425 99.200 137.755 ;
        RECT 99.425 137.425 99.680 137.755 ;
        RECT 99.005 136.455 99.175 137.425 ;
        RECT 99.850 137.255 100.020 137.925 ;
        RECT 100.930 137.855 101.175 138.460 ;
        RECT 101.395 138.130 101.905 138.665 ;
        RECT 100.655 137.685 101.885 137.855 ;
        RECT 97.145 136.285 99.175 136.455 ;
        RECT 99.345 136.115 99.515 137.255 ;
        RECT 99.685 136.285 100.020 137.255 ;
        RECT 100.195 136.115 100.485 137.280 ;
        RECT 100.655 136.875 100.995 137.685 ;
        RECT 101.165 137.120 101.915 137.310 ;
        RECT 100.655 136.465 101.170 136.875 ;
        RECT 101.405 136.115 101.575 136.875 ;
        RECT 101.745 136.455 101.915 137.120 ;
        RECT 102.085 137.135 102.275 138.495 ;
        RECT 102.445 137.645 102.720 138.495 ;
        RECT 102.910 138.130 103.440 138.495 ;
        RECT 103.865 138.265 104.195 138.665 ;
        RECT 103.265 138.095 103.440 138.130 ;
        RECT 102.445 137.475 102.725 137.645 ;
        RECT 102.445 137.335 102.720 137.475 ;
        RECT 102.925 137.135 103.095 137.935 ;
        RECT 102.085 136.965 103.095 137.135 ;
        RECT 103.265 137.925 104.195 138.095 ;
        RECT 104.365 137.925 104.620 138.495 ;
        RECT 103.265 136.795 103.435 137.925 ;
        RECT 104.025 137.755 104.195 137.925 ;
        RECT 102.310 136.625 103.435 136.795 ;
        RECT 103.605 137.425 103.800 137.755 ;
        RECT 104.025 137.425 104.280 137.755 ;
        RECT 103.605 136.455 103.775 137.425 ;
        RECT 104.450 137.255 104.620 137.925 ;
        RECT 104.855 137.845 105.065 138.665 ;
        RECT 105.235 137.865 105.565 138.495 ;
        RECT 105.235 137.265 105.485 137.865 ;
        RECT 105.735 137.845 105.965 138.665 ;
        RECT 106.265 138.115 106.435 138.495 ;
        RECT 106.615 138.285 106.945 138.665 ;
        RECT 106.265 137.945 106.930 138.115 ;
        RECT 107.125 137.990 107.385 138.495 ;
        RECT 105.655 137.425 105.985 137.675 ;
        RECT 106.195 137.395 106.525 137.765 ;
        RECT 106.760 137.690 106.930 137.945 ;
        RECT 106.760 137.360 107.045 137.690 ;
        RECT 101.745 136.285 103.775 136.455 ;
        RECT 103.945 136.115 104.115 137.255 ;
        RECT 104.285 136.285 104.620 137.255 ;
        RECT 104.855 136.115 105.065 137.255 ;
        RECT 105.235 136.285 105.565 137.265 ;
        RECT 105.735 136.115 105.965 137.255 ;
        RECT 106.760 137.215 106.930 137.360 ;
        RECT 106.265 137.045 106.930 137.215 ;
        RECT 107.215 137.190 107.385 137.990 ;
        RECT 107.645 138.115 107.815 138.495 ;
        RECT 107.995 138.285 108.325 138.665 ;
        RECT 107.645 137.945 108.310 138.115 ;
        RECT 108.505 137.990 108.765 138.495 ;
        RECT 107.575 137.395 107.905 137.765 ;
        RECT 108.140 137.690 108.310 137.945 ;
        RECT 108.140 137.360 108.425 137.690 ;
        RECT 108.140 137.215 108.310 137.360 ;
        RECT 106.265 136.285 106.435 137.045 ;
        RECT 106.615 136.115 106.945 136.875 ;
        RECT 107.115 136.285 107.385 137.190 ;
        RECT 107.645 137.045 108.310 137.215 ;
        RECT 108.595 137.190 108.765 137.990 ;
        RECT 109.395 137.895 111.985 138.665 ;
        RECT 112.155 137.915 113.365 138.665 ;
        RECT 107.645 136.285 107.815 137.045 ;
        RECT 107.995 136.115 108.325 136.875 ;
        RECT 108.495 136.285 108.765 137.190 ;
        RECT 109.395 137.205 110.605 137.725 ;
        RECT 110.775 137.375 111.985 137.895 ;
        RECT 112.155 137.205 112.675 137.745 ;
        RECT 112.845 137.375 113.365 137.915 ;
        RECT 109.395 136.115 111.985 137.205 ;
        RECT 112.155 136.115 113.365 137.205 ;
        RECT 22.830 135.945 113.450 136.115 ;
        RECT 22.915 134.855 24.125 135.945 ;
        RECT 22.915 134.145 23.435 134.685 ;
        RECT 23.605 134.315 24.125 134.855 ;
        RECT 24.355 134.805 24.565 135.945 ;
        RECT 24.735 134.795 25.065 135.775 ;
        RECT 25.235 134.805 25.465 135.945 ;
        RECT 25.765 135.015 25.935 135.775 ;
        RECT 26.115 135.185 26.445 135.945 ;
        RECT 25.765 134.845 26.430 135.015 ;
        RECT 26.615 134.870 26.885 135.775 ;
        RECT 22.915 133.395 24.125 134.145 ;
        RECT 24.355 133.395 24.565 134.215 ;
        RECT 24.735 134.195 24.985 134.795 ;
        RECT 26.260 134.700 26.430 134.845 ;
        RECT 25.155 134.385 25.485 134.635 ;
        RECT 25.695 134.295 26.025 134.665 ;
        RECT 26.260 134.370 26.545 134.700 ;
        RECT 24.735 133.565 25.065 134.195 ;
        RECT 25.235 133.395 25.465 134.215 ;
        RECT 26.260 134.115 26.430 134.370 ;
        RECT 25.765 133.945 26.430 134.115 ;
        RECT 26.715 134.070 26.885 134.870 ;
        RECT 27.095 134.805 27.325 135.945 ;
        RECT 27.495 134.795 27.825 135.775 ;
        RECT 27.995 134.805 28.205 135.945 ;
        RECT 28.440 134.805 28.775 135.775 ;
        RECT 28.945 134.805 29.115 135.945 ;
        RECT 29.285 135.605 31.315 135.775 ;
        RECT 27.075 134.385 27.405 134.635 ;
        RECT 25.765 133.565 25.935 133.945 ;
        RECT 26.115 133.395 26.445 133.775 ;
        RECT 26.625 133.565 26.885 134.070 ;
        RECT 27.095 133.395 27.325 134.215 ;
        RECT 27.575 134.195 27.825 134.795 ;
        RECT 27.495 133.565 27.825 134.195 ;
        RECT 27.995 133.395 28.205 134.215 ;
        RECT 28.440 134.135 28.610 134.805 ;
        RECT 29.285 134.635 29.455 135.605 ;
        RECT 28.780 134.305 29.035 134.635 ;
        RECT 29.260 134.305 29.455 134.635 ;
        RECT 29.625 135.265 30.750 135.435 ;
        RECT 28.865 134.135 29.035 134.305 ;
        RECT 29.625 134.135 29.795 135.265 ;
        RECT 28.440 133.565 28.695 134.135 ;
        RECT 28.865 133.965 29.795 134.135 ;
        RECT 29.965 134.925 30.975 135.095 ;
        RECT 29.965 134.125 30.135 134.925 ;
        RECT 30.340 134.245 30.615 134.725 ;
        RECT 30.335 134.075 30.615 134.245 ;
        RECT 29.620 133.930 29.795 133.965 ;
        RECT 28.865 133.395 29.195 133.795 ;
        RECT 29.620 133.565 30.150 133.930 ;
        RECT 30.340 133.565 30.615 134.075 ;
        RECT 30.785 133.565 30.975 134.925 ;
        RECT 31.145 134.940 31.315 135.605 ;
        RECT 31.485 135.185 31.655 135.945 ;
        RECT 31.890 135.185 32.405 135.595 ;
        RECT 33.695 135.275 33.975 135.945 ;
        RECT 31.145 134.750 31.895 134.940 ;
        RECT 32.065 134.375 32.405 135.185 ;
        RECT 34.145 135.055 34.445 135.605 ;
        RECT 34.645 135.225 34.975 135.945 ;
        RECT 35.165 135.225 35.625 135.775 ;
        RECT 33.510 134.635 33.775 134.995 ;
        RECT 34.145 134.885 35.085 135.055 ;
        RECT 34.915 134.635 35.085 134.885 ;
        RECT 33.510 134.385 34.185 134.635 ;
        RECT 34.405 134.385 34.745 134.635 ;
        RECT 31.175 134.205 32.405 134.375 ;
        RECT 34.915 134.305 35.205 134.635 ;
        RECT 34.915 134.215 35.085 134.305 ;
        RECT 31.155 133.395 31.665 133.930 ;
        RECT 31.885 133.600 32.130 134.205 ;
        RECT 33.695 134.025 35.085 134.215 ;
        RECT 33.695 133.665 34.025 134.025 ;
        RECT 35.375 133.855 35.625 135.225 ;
        RECT 35.795 134.780 36.085 135.945 ;
        RECT 36.345 135.275 36.515 135.775 ;
        RECT 36.685 135.445 37.015 135.945 ;
        RECT 36.345 135.105 37.010 135.275 ;
        RECT 36.260 134.285 36.610 134.935 ;
        RECT 34.645 133.395 34.895 133.855 ;
        RECT 35.065 133.565 35.625 133.855 ;
        RECT 35.795 133.395 36.085 134.120 ;
        RECT 36.780 134.115 37.010 135.105 ;
        RECT 36.345 133.945 37.010 134.115 ;
        RECT 36.345 133.655 36.515 133.945 ;
        RECT 36.685 133.395 37.015 133.775 ;
        RECT 37.185 133.655 37.410 135.775 ;
        RECT 37.625 135.445 37.955 135.945 ;
        RECT 38.125 135.275 38.295 135.775 ;
        RECT 38.530 135.560 39.360 135.730 ;
        RECT 39.600 135.565 39.980 135.945 ;
        RECT 37.600 135.105 38.295 135.275 ;
        RECT 37.600 134.135 37.770 135.105 ;
        RECT 37.940 134.315 38.350 134.935 ;
        RECT 38.520 134.885 39.020 135.265 ;
        RECT 37.600 133.945 38.295 134.135 ;
        RECT 38.520 134.015 38.740 134.885 ;
        RECT 39.190 134.715 39.360 135.560 ;
        RECT 40.160 135.395 40.330 135.685 ;
        RECT 40.500 135.565 40.830 135.945 ;
        RECT 41.300 135.475 41.930 135.725 ;
        RECT 42.110 135.565 42.530 135.945 ;
        RECT 41.760 135.395 41.930 135.475 ;
        RECT 42.730 135.395 42.970 135.685 ;
        RECT 39.530 135.145 40.900 135.395 ;
        RECT 39.530 134.885 39.780 135.145 ;
        RECT 40.290 134.715 40.540 134.875 ;
        RECT 39.190 134.545 40.540 134.715 ;
        RECT 39.190 134.505 39.610 134.545 ;
        RECT 38.920 133.955 39.270 134.325 ;
        RECT 37.625 133.395 37.955 133.775 ;
        RECT 38.125 133.615 38.295 133.945 ;
        RECT 39.440 133.775 39.610 134.505 ;
        RECT 40.710 134.375 40.900 135.145 ;
        RECT 39.780 134.045 40.190 134.375 ;
        RECT 40.480 134.035 40.900 134.375 ;
        RECT 41.070 134.965 41.590 135.275 ;
        RECT 41.760 135.225 42.970 135.395 ;
        RECT 43.200 135.255 43.530 135.945 ;
        RECT 41.070 134.205 41.240 134.965 ;
        RECT 41.410 134.375 41.590 134.785 ;
        RECT 41.760 134.715 41.930 135.225 ;
        RECT 43.700 135.075 43.870 135.685 ;
        RECT 44.140 135.225 44.470 135.735 ;
        RECT 43.700 135.055 44.020 135.075 ;
        RECT 42.100 134.885 44.020 135.055 ;
        RECT 41.760 134.545 43.660 134.715 ;
        RECT 41.990 134.205 42.320 134.325 ;
        RECT 41.070 134.035 42.320 134.205 ;
        RECT 38.595 133.575 39.610 133.775 ;
        RECT 39.780 133.395 40.190 133.835 ;
        RECT 40.480 133.605 40.730 134.035 ;
        RECT 40.930 133.395 41.250 133.855 ;
        RECT 42.490 133.785 42.660 134.545 ;
        RECT 43.330 134.485 43.660 134.545 ;
        RECT 42.850 134.315 43.180 134.375 ;
        RECT 42.850 134.045 43.510 134.315 ;
        RECT 43.830 133.990 44.020 134.885 ;
        RECT 41.810 133.615 42.660 133.785 ;
        RECT 42.860 133.395 43.520 133.875 ;
        RECT 43.700 133.660 44.020 133.990 ;
        RECT 44.220 134.635 44.470 135.225 ;
        RECT 44.650 135.145 44.935 135.945 ;
        RECT 45.115 135.605 45.370 135.635 ;
        RECT 45.115 135.435 45.455 135.605 ;
        RECT 45.920 135.435 47.575 135.725 ;
        RECT 45.115 134.965 45.370 135.435 ;
        RECT 44.220 134.305 45.020 134.635 ;
        RECT 44.220 133.655 44.470 134.305 ;
        RECT 45.190 134.105 45.370 134.965 ;
        RECT 45.920 135.095 47.510 135.265 ;
        RECT 47.745 135.145 48.025 135.945 ;
        RECT 45.920 134.805 46.240 135.095 ;
        RECT 47.340 134.975 47.510 135.095 ;
        RECT 46.435 134.755 47.150 134.925 ;
        RECT 47.340 134.805 48.065 134.975 ;
        RECT 48.235 134.805 48.505 135.775 ;
        RECT 48.880 134.975 49.210 135.775 ;
        RECT 49.380 135.145 49.710 135.945 ;
        RECT 50.010 134.975 50.340 135.775 ;
        RECT 50.985 135.145 51.235 135.945 ;
        RECT 48.880 134.805 51.315 134.975 ;
        RECT 51.505 134.805 51.675 135.945 ;
        RECT 51.845 134.805 52.185 135.775 ;
        RECT 52.410 135.145 52.710 135.945 ;
        RECT 52.880 134.975 53.210 135.775 ;
        RECT 53.380 135.145 53.550 135.945 ;
        RECT 53.720 134.975 54.050 135.775 ;
        RECT 54.220 135.145 54.390 135.945 ;
        RECT 54.560 134.975 54.890 135.775 ;
        RECT 55.060 135.145 55.230 135.945 ;
        RECT 55.400 134.975 55.730 135.775 ;
        RECT 55.900 135.145 56.155 135.945 ;
        RECT 44.650 133.395 44.935 133.855 ;
        RECT 45.115 133.575 45.370 134.105 ;
        RECT 45.920 134.065 46.270 134.635 ;
        RECT 46.440 134.305 47.150 134.755 ;
        RECT 47.895 134.635 48.065 134.805 ;
        RECT 47.320 134.305 47.725 134.635 ;
        RECT 47.895 134.305 48.165 134.635 ;
        RECT 47.895 134.135 48.065 134.305 ;
        RECT 46.455 133.965 48.065 134.135 ;
        RECT 48.335 134.070 48.505 134.805 ;
        RECT 48.675 134.385 49.025 134.635 ;
        RECT 49.210 134.175 49.380 134.805 ;
        RECT 49.550 134.385 49.880 134.585 ;
        RECT 50.050 134.385 50.380 134.585 ;
        RECT 50.550 134.385 50.970 134.585 ;
        RECT 51.145 134.555 51.315 134.805 ;
        RECT 51.145 134.385 51.840 134.555 ;
        RECT 45.925 133.395 46.255 133.895 ;
        RECT 46.455 133.615 46.625 133.965 ;
        RECT 46.825 133.395 47.155 133.795 ;
        RECT 47.325 133.615 47.495 133.965 ;
        RECT 47.665 133.395 48.045 133.795 ;
        RECT 48.235 133.725 48.505 134.070 ;
        RECT 48.880 133.565 49.380 134.175 ;
        RECT 50.010 134.045 51.235 134.215 ;
        RECT 52.010 134.195 52.185 134.805 ;
        RECT 50.010 133.565 50.340 134.045 ;
        RECT 50.510 133.395 50.735 133.855 ;
        RECT 50.905 133.565 51.235 134.045 ;
        RECT 51.425 133.395 51.675 134.195 ;
        RECT 51.845 133.565 52.185 134.195 ;
        RECT 52.355 134.805 56.325 134.975 ;
        RECT 52.355 134.215 52.675 134.805 ;
        RECT 52.875 134.585 55.730 134.635 ;
        RECT 52.875 134.415 55.805 134.585 ;
        RECT 52.875 134.385 55.730 134.415 ;
        RECT 55.980 134.215 56.325 134.805 ;
        RECT 52.355 134.025 56.325 134.215 ;
        RECT 56.495 134.805 56.835 135.775 ;
        RECT 57.005 134.805 57.175 135.945 ;
        RECT 57.445 135.145 57.695 135.945 ;
        RECT 58.340 134.975 58.670 135.775 ;
        RECT 58.970 135.145 59.300 135.945 ;
        RECT 59.470 134.975 59.800 135.775 ;
        RECT 57.365 134.805 59.800 134.975 ;
        RECT 60.215 134.805 60.445 135.945 ;
        RECT 56.495 134.195 56.670 134.805 ;
        RECT 57.365 134.555 57.535 134.805 ;
        RECT 56.840 134.385 57.535 134.555 ;
        RECT 57.710 134.385 58.130 134.585 ;
        RECT 58.300 134.385 58.630 134.585 ;
        RECT 58.800 134.385 59.130 134.585 ;
        RECT 52.405 133.395 52.710 133.855 ;
        RECT 52.880 133.565 53.210 134.025 ;
        RECT 53.380 133.395 53.550 133.855 ;
        RECT 53.720 133.565 54.050 134.025 ;
        RECT 54.220 133.395 54.390 133.855 ;
        RECT 54.560 133.565 54.890 134.025 ;
        RECT 55.060 133.395 55.230 133.855 ;
        RECT 55.400 133.565 55.730 134.025 ;
        RECT 55.900 133.395 56.155 133.855 ;
        RECT 56.495 133.565 56.835 134.195 ;
        RECT 57.005 133.395 57.255 134.195 ;
        RECT 57.445 134.045 58.670 134.215 ;
        RECT 57.445 133.565 57.775 134.045 ;
        RECT 57.945 133.395 58.170 133.855 ;
        RECT 58.340 133.565 58.670 134.045 ;
        RECT 59.300 134.175 59.470 134.805 ;
        RECT 60.615 134.795 60.945 135.775 ;
        RECT 61.115 134.805 61.325 135.945 ;
        RECT 59.655 134.385 60.005 134.635 ;
        RECT 60.195 134.385 60.525 134.635 ;
        RECT 59.300 133.565 59.800 134.175 ;
        RECT 60.215 133.395 60.445 134.215 ;
        RECT 60.695 134.195 60.945 134.795 ;
        RECT 61.555 134.780 61.845 135.945 ;
        RECT 62.390 135.605 62.645 135.635 ;
        RECT 62.305 135.435 62.645 135.605 ;
        RECT 62.390 134.965 62.645 135.435 ;
        RECT 62.825 135.145 63.110 135.945 ;
        RECT 63.290 135.225 63.620 135.735 ;
        RECT 60.615 133.565 60.945 134.195 ;
        RECT 61.115 133.395 61.325 134.215 ;
        RECT 61.555 133.395 61.845 134.120 ;
        RECT 62.390 134.105 62.570 134.965 ;
        RECT 63.290 134.635 63.540 135.225 ;
        RECT 63.890 135.075 64.060 135.685 ;
        RECT 64.230 135.255 64.560 135.945 ;
        RECT 64.790 135.395 65.030 135.685 ;
        RECT 65.230 135.565 65.650 135.945 ;
        RECT 65.830 135.475 66.460 135.725 ;
        RECT 66.930 135.565 67.260 135.945 ;
        RECT 65.830 135.395 66.000 135.475 ;
        RECT 67.430 135.395 67.600 135.685 ;
        RECT 67.780 135.565 68.160 135.945 ;
        RECT 68.400 135.560 69.230 135.730 ;
        RECT 64.790 135.225 66.000 135.395 ;
        RECT 62.740 134.305 63.540 134.635 ;
        RECT 62.390 133.575 62.645 134.105 ;
        RECT 62.825 133.395 63.110 133.855 ;
        RECT 63.290 133.655 63.540 134.305 ;
        RECT 63.740 135.055 64.060 135.075 ;
        RECT 63.740 134.885 65.660 135.055 ;
        RECT 63.740 133.990 63.930 134.885 ;
        RECT 65.830 134.715 66.000 135.225 ;
        RECT 66.170 134.965 66.690 135.275 ;
        RECT 64.100 134.545 66.000 134.715 ;
        RECT 64.100 134.485 64.430 134.545 ;
        RECT 64.580 134.315 64.910 134.375 ;
        RECT 64.250 134.045 64.910 134.315 ;
        RECT 63.740 133.660 64.060 133.990 ;
        RECT 64.240 133.395 64.900 133.875 ;
        RECT 65.100 133.785 65.270 134.545 ;
        RECT 66.170 134.375 66.350 134.785 ;
        RECT 65.440 134.205 65.770 134.325 ;
        RECT 66.520 134.205 66.690 134.965 ;
        RECT 65.440 134.035 66.690 134.205 ;
        RECT 66.860 135.145 68.230 135.395 ;
        RECT 66.860 134.375 67.050 135.145 ;
        RECT 67.980 134.885 68.230 135.145 ;
        RECT 67.220 134.715 67.470 134.875 ;
        RECT 68.400 134.715 68.570 135.560 ;
        RECT 69.465 135.275 69.635 135.775 ;
        RECT 69.805 135.445 70.135 135.945 ;
        RECT 68.740 134.885 69.240 135.265 ;
        RECT 69.465 135.105 70.160 135.275 ;
        RECT 67.220 134.545 68.570 134.715 ;
        RECT 68.150 134.505 68.570 134.545 ;
        RECT 66.860 134.035 67.280 134.375 ;
        RECT 67.570 134.045 67.980 134.375 ;
        RECT 65.100 133.615 65.950 133.785 ;
        RECT 66.510 133.395 66.830 133.855 ;
        RECT 67.030 133.605 67.280 134.035 ;
        RECT 67.570 133.395 67.980 133.835 ;
        RECT 68.150 133.775 68.320 134.505 ;
        RECT 68.490 133.955 68.840 134.325 ;
        RECT 69.020 134.015 69.240 134.885 ;
        RECT 69.410 134.315 69.820 134.935 ;
        RECT 69.990 134.135 70.160 135.105 ;
        RECT 69.465 133.945 70.160 134.135 ;
        RECT 68.150 133.575 69.165 133.775 ;
        RECT 69.465 133.615 69.635 133.945 ;
        RECT 69.805 133.395 70.135 133.775 ;
        RECT 70.350 133.655 70.575 135.775 ;
        RECT 70.745 135.445 71.075 135.945 ;
        RECT 71.245 135.275 71.415 135.775 ;
        RECT 70.750 135.105 71.415 135.275 ;
        RECT 72.135 135.110 72.520 135.945 ;
        RECT 70.750 134.115 70.980 135.105 ;
        RECT 72.690 134.940 72.950 135.745 ;
        RECT 73.120 135.110 73.380 135.945 ;
        RECT 73.550 134.940 73.805 135.745 ;
        RECT 73.980 135.110 74.240 135.945 ;
        RECT 74.410 134.940 74.665 135.745 ;
        RECT 74.840 135.110 75.185 135.945 ;
        RECT 75.730 135.605 75.985 135.635 ;
        RECT 75.645 135.435 75.985 135.605 ;
        RECT 75.730 134.965 75.985 135.435 ;
        RECT 76.165 135.145 76.450 135.945 ;
        RECT 76.630 135.225 76.960 135.735 ;
        RECT 71.150 134.285 71.500 134.935 ;
        RECT 72.135 134.770 75.165 134.940 ;
        RECT 72.135 134.205 72.435 134.770 ;
        RECT 72.610 134.375 74.825 134.600 ;
        RECT 74.995 134.205 75.165 134.770 ;
        RECT 70.750 133.945 71.415 134.115 ;
        RECT 72.135 134.035 75.165 134.205 ;
        RECT 75.730 134.105 75.910 134.965 ;
        RECT 76.630 134.635 76.880 135.225 ;
        RECT 77.230 135.075 77.400 135.685 ;
        RECT 77.570 135.255 77.900 135.945 ;
        RECT 78.130 135.395 78.370 135.685 ;
        RECT 78.570 135.565 78.990 135.945 ;
        RECT 79.170 135.475 79.800 135.725 ;
        RECT 80.270 135.565 80.600 135.945 ;
        RECT 79.170 135.395 79.340 135.475 ;
        RECT 80.770 135.395 80.940 135.685 ;
        RECT 81.120 135.565 81.500 135.945 ;
        RECT 81.740 135.560 82.570 135.730 ;
        RECT 78.130 135.225 79.340 135.395 ;
        RECT 76.080 134.305 76.880 134.635 ;
        RECT 70.745 133.395 71.075 133.775 ;
        RECT 71.245 133.655 71.415 133.945 ;
        RECT 72.655 133.395 72.955 133.865 ;
        RECT 73.125 133.590 73.380 134.035 ;
        RECT 73.550 133.395 73.810 133.865 ;
        RECT 73.980 133.590 74.240 134.035 ;
        RECT 74.410 133.395 74.705 133.865 ;
        RECT 75.730 133.575 75.985 134.105 ;
        RECT 76.165 133.395 76.450 133.855 ;
        RECT 76.630 133.655 76.880 134.305 ;
        RECT 77.080 135.055 77.400 135.075 ;
        RECT 77.080 134.885 79.000 135.055 ;
        RECT 77.080 133.990 77.270 134.885 ;
        RECT 79.170 134.715 79.340 135.225 ;
        RECT 79.510 134.965 80.030 135.275 ;
        RECT 77.440 134.545 79.340 134.715 ;
        RECT 77.440 134.485 77.770 134.545 ;
        RECT 77.920 134.315 78.250 134.375 ;
        RECT 77.590 134.045 78.250 134.315 ;
        RECT 77.080 133.660 77.400 133.990 ;
        RECT 77.580 133.395 78.240 133.875 ;
        RECT 78.440 133.785 78.610 134.545 ;
        RECT 79.510 134.375 79.690 134.785 ;
        RECT 78.780 134.205 79.110 134.325 ;
        RECT 79.860 134.205 80.030 134.965 ;
        RECT 78.780 134.035 80.030 134.205 ;
        RECT 80.200 135.145 81.570 135.395 ;
        RECT 80.200 134.375 80.390 135.145 ;
        RECT 81.320 134.885 81.570 135.145 ;
        RECT 80.560 134.715 80.810 134.875 ;
        RECT 81.740 134.715 81.910 135.560 ;
        RECT 82.805 135.275 82.975 135.775 ;
        RECT 83.145 135.445 83.475 135.945 ;
        RECT 82.080 134.885 82.580 135.265 ;
        RECT 82.805 135.105 83.500 135.275 ;
        RECT 80.560 134.545 81.910 134.715 ;
        RECT 81.490 134.505 81.910 134.545 ;
        RECT 80.200 134.035 80.620 134.375 ;
        RECT 80.910 134.045 81.320 134.375 ;
        RECT 78.440 133.615 79.290 133.785 ;
        RECT 79.850 133.395 80.170 133.855 ;
        RECT 80.370 133.605 80.620 134.035 ;
        RECT 80.910 133.395 81.320 133.835 ;
        RECT 81.490 133.775 81.660 134.505 ;
        RECT 81.830 133.955 82.180 134.325 ;
        RECT 82.360 134.015 82.580 134.885 ;
        RECT 82.750 134.315 83.160 134.935 ;
        RECT 83.330 134.135 83.500 135.105 ;
        RECT 82.805 133.945 83.500 134.135 ;
        RECT 81.490 133.575 82.505 133.775 ;
        RECT 82.805 133.615 82.975 133.945 ;
        RECT 83.145 133.395 83.475 133.775 ;
        RECT 83.690 133.655 83.915 135.775 ;
        RECT 84.085 135.445 84.415 135.945 ;
        RECT 84.585 135.275 84.755 135.775 ;
        RECT 84.090 135.105 84.755 135.275 ;
        RECT 84.090 134.115 84.320 135.105 ;
        RECT 84.490 134.285 84.840 134.935 ;
        RECT 85.975 134.805 86.205 135.945 ;
        RECT 86.375 134.795 86.705 135.775 ;
        RECT 86.875 134.805 87.085 135.945 ;
        RECT 85.955 134.385 86.285 134.635 ;
        RECT 84.090 133.945 84.755 134.115 ;
        RECT 84.085 133.395 84.415 133.775 ;
        RECT 84.585 133.655 84.755 133.945 ;
        RECT 85.975 133.395 86.205 134.215 ;
        RECT 86.455 134.195 86.705 134.795 ;
        RECT 87.315 134.780 87.605 135.945 ;
        RECT 88.735 134.805 88.965 135.945 ;
        RECT 89.135 134.795 89.465 135.775 ;
        RECT 89.635 134.805 89.845 135.945 ;
        RECT 90.075 134.870 90.345 135.775 ;
        RECT 90.515 135.185 90.845 135.945 ;
        RECT 91.025 135.015 91.195 135.775 ;
        RECT 88.715 134.385 89.045 134.635 ;
        RECT 86.375 133.565 86.705 134.195 ;
        RECT 86.875 133.395 87.085 134.215 ;
        RECT 87.315 133.395 87.605 134.120 ;
        RECT 88.735 133.395 88.965 134.215 ;
        RECT 89.215 134.195 89.465 134.795 ;
        RECT 89.135 133.565 89.465 134.195 ;
        RECT 89.635 133.395 89.845 134.215 ;
        RECT 90.075 134.070 90.245 134.870 ;
        RECT 90.530 134.845 91.195 135.015 ;
        RECT 92.290 134.965 92.545 135.635 ;
        RECT 92.725 135.145 93.010 135.945 ;
        RECT 93.190 135.225 93.520 135.735 ;
        RECT 92.290 134.925 92.470 134.965 ;
        RECT 90.530 134.700 90.700 134.845 ;
        RECT 92.205 134.755 92.470 134.925 ;
        RECT 90.415 134.370 90.700 134.700 ;
        RECT 90.530 134.115 90.700 134.370 ;
        RECT 90.935 134.295 91.265 134.665 ;
        RECT 90.075 133.565 90.335 134.070 ;
        RECT 90.530 133.945 91.195 134.115 ;
        RECT 90.515 133.395 90.845 133.775 ;
        RECT 91.025 133.565 91.195 133.945 ;
        RECT 92.290 134.105 92.470 134.755 ;
        RECT 93.190 134.635 93.440 135.225 ;
        RECT 93.790 135.075 93.960 135.685 ;
        RECT 94.130 135.255 94.460 135.945 ;
        RECT 94.690 135.395 94.930 135.685 ;
        RECT 95.130 135.565 95.550 135.945 ;
        RECT 95.730 135.475 96.360 135.725 ;
        RECT 96.830 135.565 97.160 135.945 ;
        RECT 95.730 135.395 95.900 135.475 ;
        RECT 97.330 135.395 97.500 135.685 ;
        RECT 97.680 135.565 98.060 135.945 ;
        RECT 98.300 135.560 99.130 135.730 ;
        RECT 94.690 135.225 95.900 135.395 ;
        RECT 92.640 134.305 93.440 134.635 ;
        RECT 92.290 133.575 92.545 134.105 ;
        RECT 92.725 133.395 93.010 133.855 ;
        RECT 93.190 133.655 93.440 134.305 ;
        RECT 93.640 135.055 93.960 135.075 ;
        RECT 93.640 134.885 95.560 135.055 ;
        RECT 93.640 133.990 93.830 134.885 ;
        RECT 95.730 134.715 95.900 135.225 ;
        RECT 96.070 134.965 96.590 135.275 ;
        RECT 94.000 134.545 95.900 134.715 ;
        RECT 94.000 134.485 94.330 134.545 ;
        RECT 94.480 134.315 94.810 134.375 ;
        RECT 94.150 134.045 94.810 134.315 ;
        RECT 93.640 133.660 93.960 133.990 ;
        RECT 94.140 133.395 94.800 133.875 ;
        RECT 95.000 133.785 95.170 134.545 ;
        RECT 96.070 134.375 96.250 134.785 ;
        RECT 95.340 134.205 95.670 134.325 ;
        RECT 96.420 134.205 96.590 134.965 ;
        RECT 95.340 134.035 96.590 134.205 ;
        RECT 96.760 135.145 98.130 135.395 ;
        RECT 96.760 134.375 96.950 135.145 ;
        RECT 97.880 134.885 98.130 135.145 ;
        RECT 97.120 134.715 97.370 134.875 ;
        RECT 98.300 134.715 98.470 135.560 ;
        RECT 99.365 135.275 99.535 135.775 ;
        RECT 99.705 135.445 100.035 135.945 ;
        RECT 98.640 134.885 99.140 135.265 ;
        RECT 99.365 135.105 100.060 135.275 ;
        RECT 97.120 134.545 98.470 134.715 ;
        RECT 98.050 134.505 98.470 134.545 ;
        RECT 96.760 134.035 97.180 134.375 ;
        RECT 97.470 134.045 97.880 134.375 ;
        RECT 95.000 133.615 95.850 133.785 ;
        RECT 96.410 133.395 96.730 133.855 ;
        RECT 96.930 133.605 97.180 134.035 ;
        RECT 97.470 133.395 97.880 133.835 ;
        RECT 98.050 133.775 98.220 134.505 ;
        RECT 98.390 133.955 98.740 134.325 ;
        RECT 98.920 134.015 99.140 134.885 ;
        RECT 99.310 134.315 99.720 134.935 ;
        RECT 99.890 134.135 100.060 135.105 ;
        RECT 99.365 133.945 100.060 134.135 ;
        RECT 98.050 133.575 99.065 133.775 ;
        RECT 99.365 133.615 99.535 133.945 ;
        RECT 99.705 133.395 100.035 133.775 ;
        RECT 100.250 133.655 100.475 135.775 ;
        RECT 100.645 135.445 100.975 135.945 ;
        RECT 101.145 135.275 101.315 135.775 ;
        RECT 102.410 135.605 102.665 135.635 ;
        RECT 102.325 135.435 102.665 135.605 ;
        RECT 100.650 135.105 101.315 135.275 ;
        RECT 100.650 134.115 100.880 135.105 ;
        RECT 102.410 134.965 102.665 135.435 ;
        RECT 102.845 135.145 103.130 135.945 ;
        RECT 103.310 135.225 103.640 135.735 ;
        RECT 101.050 134.285 101.400 134.935 ;
        RECT 100.650 133.945 101.315 134.115 ;
        RECT 100.645 133.395 100.975 133.775 ;
        RECT 101.145 133.655 101.315 133.945 ;
        RECT 102.410 134.105 102.590 134.965 ;
        RECT 103.310 134.635 103.560 135.225 ;
        RECT 103.910 135.075 104.080 135.685 ;
        RECT 104.250 135.255 104.580 135.945 ;
        RECT 104.810 135.395 105.050 135.685 ;
        RECT 105.250 135.565 105.670 135.945 ;
        RECT 105.850 135.475 106.480 135.725 ;
        RECT 106.950 135.565 107.280 135.945 ;
        RECT 105.850 135.395 106.020 135.475 ;
        RECT 107.450 135.395 107.620 135.685 ;
        RECT 107.800 135.565 108.180 135.945 ;
        RECT 108.420 135.560 109.250 135.730 ;
        RECT 104.810 135.225 106.020 135.395 ;
        RECT 102.760 134.305 103.560 134.635 ;
        RECT 102.410 133.575 102.665 134.105 ;
        RECT 102.845 133.395 103.130 133.855 ;
        RECT 103.310 133.655 103.560 134.305 ;
        RECT 103.760 135.055 104.080 135.075 ;
        RECT 103.760 134.885 105.680 135.055 ;
        RECT 103.760 133.990 103.950 134.885 ;
        RECT 105.850 134.715 106.020 135.225 ;
        RECT 106.190 134.965 106.710 135.275 ;
        RECT 104.120 134.545 106.020 134.715 ;
        RECT 104.120 134.485 104.450 134.545 ;
        RECT 104.600 134.315 104.930 134.375 ;
        RECT 104.270 134.045 104.930 134.315 ;
        RECT 103.760 133.660 104.080 133.990 ;
        RECT 104.260 133.395 104.920 133.875 ;
        RECT 105.120 133.785 105.290 134.545 ;
        RECT 106.190 134.375 106.370 134.785 ;
        RECT 105.460 134.205 105.790 134.325 ;
        RECT 106.540 134.205 106.710 134.965 ;
        RECT 105.460 134.035 106.710 134.205 ;
        RECT 106.880 135.145 108.250 135.395 ;
        RECT 106.880 134.375 107.070 135.145 ;
        RECT 108.000 134.885 108.250 135.145 ;
        RECT 107.240 134.715 107.490 134.875 ;
        RECT 108.420 134.715 108.590 135.560 ;
        RECT 109.485 135.275 109.655 135.775 ;
        RECT 109.825 135.445 110.155 135.945 ;
        RECT 108.760 134.885 109.260 135.265 ;
        RECT 109.485 135.105 110.180 135.275 ;
        RECT 107.240 134.545 108.590 134.715 ;
        RECT 108.170 134.505 108.590 134.545 ;
        RECT 106.880 134.035 107.300 134.375 ;
        RECT 107.590 134.045 108.000 134.375 ;
        RECT 105.120 133.615 105.970 133.785 ;
        RECT 106.530 133.395 106.850 133.855 ;
        RECT 107.050 133.605 107.300 134.035 ;
        RECT 107.590 133.395 108.000 133.835 ;
        RECT 108.170 133.775 108.340 134.505 ;
        RECT 108.510 133.955 108.860 134.325 ;
        RECT 109.040 134.015 109.260 134.885 ;
        RECT 109.430 134.315 109.840 134.935 ;
        RECT 110.010 134.135 110.180 135.105 ;
        RECT 109.485 133.945 110.180 134.135 ;
        RECT 108.170 133.575 109.185 133.775 ;
        RECT 109.485 133.615 109.655 133.945 ;
        RECT 109.825 133.395 110.155 133.775 ;
        RECT 110.370 133.655 110.595 135.775 ;
        RECT 110.765 135.445 111.095 135.945 ;
        RECT 111.265 135.275 111.435 135.775 ;
        RECT 110.770 135.105 111.435 135.275 ;
        RECT 110.770 134.115 111.000 135.105 ;
        RECT 111.170 134.285 111.520 134.935 ;
        RECT 112.155 134.855 113.365 135.945 ;
        RECT 112.155 134.315 112.675 134.855 ;
        RECT 112.845 134.145 113.365 134.685 ;
        RECT 110.770 133.945 111.435 134.115 ;
        RECT 110.765 133.395 111.095 133.775 ;
        RECT 111.265 133.655 111.435 133.945 ;
        RECT 112.155 133.395 113.365 134.145 ;
        RECT 22.830 133.225 113.450 133.395 ;
        RECT 22.915 132.475 24.125 133.225 ;
        RECT 24.670 132.515 24.925 133.045 ;
        RECT 25.105 132.765 25.390 133.225 ;
        RECT 22.915 131.935 23.435 132.475 ;
        RECT 23.605 131.765 24.125 132.305 ;
        RECT 22.915 130.675 24.125 131.765 ;
        RECT 24.670 131.655 24.850 132.515 ;
        RECT 25.570 132.315 25.820 132.965 ;
        RECT 25.020 131.985 25.820 132.315 ;
        RECT 24.670 131.185 24.925 131.655 ;
        RECT 24.585 131.015 24.925 131.185 ;
        RECT 24.670 130.985 24.925 131.015 ;
        RECT 25.105 130.675 25.390 131.475 ;
        RECT 25.570 131.395 25.820 131.985 ;
        RECT 26.020 132.630 26.340 132.960 ;
        RECT 26.520 132.745 27.180 133.225 ;
        RECT 27.380 132.835 28.230 133.005 ;
        RECT 26.020 131.735 26.210 132.630 ;
        RECT 26.530 132.305 27.190 132.575 ;
        RECT 26.860 132.245 27.190 132.305 ;
        RECT 26.380 132.075 26.710 132.135 ;
        RECT 27.380 132.075 27.550 132.835 ;
        RECT 28.790 132.765 29.110 133.225 ;
        RECT 29.310 132.585 29.560 133.015 ;
        RECT 29.850 132.785 30.260 133.225 ;
        RECT 30.430 132.845 31.445 133.045 ;
        RECT 27.720 132.415 28.970 132.585 ;
        RECT 27.720 132.295 28.050 132.415 ;
        RECT 26.380 131.905 28.280 132.075 ;
        RECT 26.020 131.565 27.940 131.735 ;
        RECT 26.020 131.545 26.340 131.565 ;
        RECT 25.570 130.885 25.900 131.395 ;
        RECT 26.170 130.935 26.340 131.545 ;
        RECT 28.110 131.395 28.280 131.905 ;
        RECT 28.450 131.835 28.630 132.245 ;
        RECT 28.800 131.655 28.970 132.415 ;
        RECT 26.510 130.675 26.840 131.365 ;
        RECT 27.070 131.225 28.280 131.395 ;
        RECT 28.450 131.345 28.970 131.655 ;
        RECT 29.140 132.245 29.560 132.585 ;
        RECT 29.850 132.245 30.260 132.575 ;
        RECT 29.140 131.475 29.330 132.245 ;
        RECT 30.430 132.115 30.600 132.845 ;
        RECT 31.745 132.675 31.915 133.005 ;
        RECT 32.085 132.845 32.415 133.225 ;
        RECT 30.770 132.295 31.120 132.665 ;
        RECT 30.430 132.075 30.850 132.115 ;
        RECT 29.500 131.905 30.850 132.075 ;
        RECT 29.500 131.745 29.750 131.905 ;
        RECT 30.260 131.475 30.510 131.735 ;
        RECT 29.140 131.225 30.510 131.475 ;
        RECT 27.070 130.935 27.310 131.225 ;
        RECT 28.110 131.145 28.280 131.225 ;
        RECT 27.510 130.675 27.930 131.055 ;
        RECT 28.110 130.895 28.740 131.145 ;
        RECT 29.210 130.675 29.540 131.055 ;
        RECT 29.710 130.935 29.880 131.225 ;
        RECT 30.680 131.060 30.850 131.905 ;
        RECT 31.300 131.735 31.520 132.605 ;
        RECT 31.745 132.485 32.440 132.675 ;
        RECT 31.020 131.355 31.520 131.735 ;
        RECT 31.690 131.685 32.100 132.305 ;
        RECT 32.270 131.515 32.440 132.485 ;
        RECT 31.745 131.345 32.440 131.515 ;
        RECT 30.060 130.675 30.440 131.055 ;
        RECT 30.680 130.890 31.510 131.060 ;
        RECT 31.745 130.845 31.915 131.345 ;
        RECT 32.085 130.675 32.415 131.175 ;
        RECT 32.630 130.845 32.855 132.965 ;
        RECT 33.025 132.845 33.355 133.225 ;
        RECT 33.525 132.675 33.695 132.965 ;
        RECT 33.030 132.505 33.695 132.675 ;
        RECT 33.030 131.515 33.260 132.505 ;
        RECT 34.690 132.415 34.935 133.020 ;
        RECT 35.155 132.690 35.665 133.225 ;
        RECT 33.430 131.685 33.780 132.335 ;
        RECT 34.415 132.245 35.645 132.415 ;
        RECT 33.030 131.345 33.695 131.515 ;
        RECT 33.025 130.675 33.355 131.175 ;
        RECT 33.525 130.845 33.695 131.345 ;
        RECT 34.415 131.435 34.755 132.245 ;
        RECT 34.925 131.680 35.675 131.870 ;
        RECT 34.415 131.025 34.930 131.435 ;
        RECT 35.165 130.675 35.335 131.435 ;
        RECT 35.505 131.015 35.675 131.680 ;
        RECT 35.845 131.695 36.035 133.055 ;
        RECT 36.205 132.205 36.480 133.055 ;
        RECT 36.670 132.690 37.200 133.055 ;
        RECT 37.625 132.825 37.955 133.225 ;
        RECT 37.025 132.655 37.200 132.690 ;
        RECT 36.205 132.035 36.485 132.205 ;
        RECT 36.205 131.895 36.480 132.035 ;
        RECT 36.685 131.695 36.855 132.495 ;
        RECT 35.845 131.525 36.855 131.695 ;
        RECT 37.025 132.485 37.955 132.655 ;
        RECT 38.125 132.485 38.380 133.055 ;
        RECT 37.025 131.355 37.195 132.485 ;
        RECT 37.785 132.315 37.955 132.485 ;
        RECT 36.070 131.185 37.195 131.355 ;
        RECT 37.365 131.985 37.560 132.315 ;
        RECT 37.785 131.985 38.040 132.315 ;
        RECT 37.365 131.015 37.535 131.985 ;
        RECT 38.210 131.815 38.380 132.485 ;
        RECT 35.505 130.845 37.535 131.015 ;
        RECT 37.705 130.675 37.875 131.815 ;
        RECT 38.045 130.845 38.380 131.815 ;
        RECT 38.560 132.485 38.815 133.055 ;
        RECT 38.985 132.825 39.315 133.225 ;
        RECT 39.740 132.690 40.270 133.055 ;
        RECT 39.740 132.655 39.915 132.690 ;
        RECT 38.985 132.485 39.915 132.655 ;
        RECT 38.560 131.815 38.730 132.485 ;
        RECT 38.985 132.315 39.155 132.485 ;
        RECT 38.900 131.985 39.155 132.315 ;
        RECT 39.380 131.985 39.575 132.315 ;
        RECT 38.560 130.845 38.895 131.815 ;
        RECT 39.065 130.675 39.235 131.815 ;
        RECT 39.405 131.015 39.575 131.985 ;
        RECT 39.745 131.355 39.915 132.485 ;
        RECT 40.085 131.695 40.255 132.495 ;
        RECT 40.460 132.205 40.735 133.055 ;
        RECT 40.455 132.035 40.735 132.205 ;
        RECT 40.460 131.895 40.735 132.035 ;
        RECT 40.905 131.695 41.095 133.055 ;
        RECT 41.275 132.690 41.785 133.225 ;
        RECT 42.005 132.415 42.250 133.020 ;
        RECT 42.700 132.485 42.955 133.055 ;
        RECT 43.125 132.825 43.455 133.225 ;
        RECT 43.880 132.690 44.410 133.055 ;
        RECT 44.600 132.885 44.875 133.055 ;
        RECT 44.595 132.715 44.875 132.885 ;
        RECT 43.880 132.655 44.055 132.690 ;
        RECT 43.125 132.485 44.055 132.655 ;
        RECT 41.295 132.245 42.525 132.415 ;
        RECT 40.085 131.525 41.095 131.695 ;
        RECT 41.265 131.680 42.015 131.870 ;
        RECT 39.745 131.185 40.870 131.355 ;
        RECT 41.265 131.015 41.435 131.680 ;
        RECT 42.185 131.435 42.525 132.245 ;
        RECT 39.405 130.845 41.435 131.015 ;
        RECT 41.605 130.675 41.775 131.435 ;
        RECT 42.010 131.025 42.525 131.435 ;
        RECT 42.700 131.815 42.870 132.485 ;
        RECT 43.125 132.315 43.295 132.485 ;
        RECT 43.040 131.985 43.295 132.315 ;
        RECT 43.520 131.985 43.715 132.315 ;
        RECT 42.700 130.845 43.035 131.815 ;
        RECT 43.205 130.675 43.375 131.815 ;
        RECT 43.545 131.015 43.715 131.985 ;
        RECT 43.885 131.355 44.055 132.485 ;
        RECT 44.225 131.695 44.395 132.495 ;
        RECT 44.600 131.895 44.875 132.715 ;
        RECT 45.045 131.695 45.235 133.055 ;
        RECT 45.415 132.690 45.925 133.225 ;
        RECT 46.145 132.415 46.390 133.020 ;
        RECT 45.435 132.245 46.665 132.415 ;
        RECT 46.875 132.405 47.105 133.225 ;
        RECT 47.275 132.425 47.605 133.055 ;
        RECT 44.225 131.525 45.235 131.695 ;
        RECT 45.405 131.680 46.155 131.870 ;
        RECT 43.885 131.185 45.010 131.355 ;
        RECT 45.405 131.015 45.575 131.680 ;
        RECT 46.325 131.435 46.665 132.245 ;
        RECT 46.855 131.985 47.185 132.235 ;
        RECT 47.355 131.825 47.605 132.425 ;
        RECT 47.775 132.405 47.985 133.225 ;
        RECT 48.675 132.500 48.965 133.225 ;
        RECT 49.135 132.550 49.405 132.895 ;
        RECT 49.595 132.825 49.975 133.225 ;
        RECT 50.145 132.655 50.315 133.005 ;
        RECT 50.485 132.825 50.815 133.225 ;
        RECT 51.015 132.655 51.185 133.005 ;
        RECT 51.385 132.725 51.715 133.225 ;
        RECT 43.545 130.845 45.575 131.015 ;
        RECT 45.745 130.675 45.915 131.435 ;
        RECT 46.150 131.025 46.665 131.435 ;
        RECT 46.875 130.675 47.105 131.815 ;
        RECT 47.275 130.845 47.605 131.825 ;
        RECT 47.775 130.675 47.985 131.815 ;
        RECT 48.675 130.675 48.965 131.840 ;
        RECT 49.135 131.815 49.305 132.550 ;
        RECT 49.575 132.485 51.185 132.655 ;
        RECT 51.985 132.675 52.155 133.055 ;
        RECT 52.335 132.845 52.665 133.225 ;
        RECT 49.575 132.315 49.745 132.485 ;
        RECT 49.475 131.985 49.745 132.315 ;
        RECT 49.915 131.985 50.320 132.315 ;
        RECT 49.575 131.815 49.745 131.985 ;
        RECT 50.490 131.865 51.200 132.315 ;
        RECT 51.370 131.985 51.720 132.555 ;
        RECT 51.985 132.505 52.650 132.675 ;
        RECT 52.845 132.550 53.105 133.055 ;
        RECT 51.915 131.955 52.245 132.325 ;
        RECT 52.480 132.250 52.650 132.505 ;
        RECT 52.480 131.920 52.765 132.250 ;
        RECT 49.135 130.845 49.405 131.815 ;
        RECT 49.575 131.645 50.300 131.815 ;
        RECT 50.490 131.695 51.205 131.865 ;
        RECT 50.130 131.525 50.300 131.645 ;
        RECT 51.400 131.525 51.720 131.815 ;
        RECT 52.480 131.775 52.650 131.920 ;
        RECT 49.615 130.675 49.895 131.475 ;
        RECT 50.130 131.355 51.720 131.525 ;
        RECT 51.985 131.605 52.650 131.775 ;
        RECT 52.935 131.750 53.105 132.550 ;
        RECT 53.550 132.415 53.795 133.020 ;
        RECT 54.015 132.690 54.525 133.225 ;
        RECT 50.065 130.895 51.720 131.185 ;
        RECT 51.985 130.845 52.155 131.605 ;
        RECT 52.335 130.675 52.665 131.435 ;
        RECT 52.835 130.845 53.105 131.750 ;
        RECT 53.275 132.245 54.505 132.415 ;
        RECT 53.275 131.435 53.615 132.245 ;
        RECT 53.785 131.680 54.535 131.870 ;
        RECT 53.275 131.025 53.790 131.435 ;
        RECT 54.025 130.675 54.195 131.435 ;
        RECT 54.365 131.015 54.535 131.680 ;
        RECT 54.705 131.695 54.895 133.055 ;
        RECT 55.065 132.545 55.340 133.055 ;
        RECT 55.530 132.690 56.060 133.055 ;
        RECT 56.485 132.825 56.815 133.225 ;
        RECT 55.885 132.655 56.060 132.690 ;
        RECT 55.065 132.375 55.345 132.545 ;
        RECT 55.065 131.895 55.340 132.375 ;
        RECT 55.545 131.695 55.715 132.495 ;
        RECT 54.705 131.525 55.715 131.695 ;
        RECT 55.885 132.485 56.815 132.655 ;
        RECT 56.985 132.485 57.240 133.055 ;
        RECT 55.885 131.355 56.055 132.485 ;
        RECT 56.645 132.315 56.815 132.485 ;
        RECT 54.930 131.185 56.055 131.355 ;
        RECT 56.225 131.985 56.420 132.315 ;
        RECT 56.645 131.985 56.900 132.315 ;
        RECT 56.225 131.015 56.395 131.985 ;
        RECT 57.070 131.815 57.240 132.485 ;
        RECT 57.690 132.415 57.935 133.020 ;
        RECT 58.155 132.690 58.665 133.225 ;
        RECT 54.365 130.845 56.395 131.015 ;
        RECT 56.565 130.675 56.735 131.815 ;
        RECT 56.905 130.845 57.240 131.815 ;
        RECT 57.415 132.245 58.645 132.415 ;
        RECT 57.415 131.435 57.755 132.245 ;
        RECT 57.925 131.680 58.675 131.870 ;
        RECT 57.415 131.025 57.930 131.435 ;
        RECT 58.165 130.675 58.335 131.435 ;
        RECT 58.505 131.015 58.675 131.680 ;
        RECT 58.845 131.695 59.035 133.055 ;
        RECT 59.205 132.205 59.480 133.055 ;
        RECT 59.670 132.690 60.200 133.055 ;
        RECT 60.625 132.825 60.955 133.225 ;
        RECT 60.025 132.655 60.200 132.690 ;
        RECT 59.205 132.035 59.485 132.205 ;
        RECT 59.205 131.895 59.480 132.035 ;
        RECT 59.685 131.695 59.855 132.495 ;
        RECT 58.845 131.525 59.855 131.695 ;
        RECT 60.025 132.485 60.955 132.655 ;
        RECT 61.125 132.485 61.380 133.055 ;
        RECT 60.025 131.355 60.195 132.485 ;
        RECT 60.785 132.315 60.955 132.485 ;
        RECT 59.070 131.185 60.195 131.355 ;
        RECT 60.365 131.985 60.560 132.315 ;
        RECT 60.785 131.985 61.040 132.315 ;
        RECT 60.365 131.015 60.535 131.985 ;
        RECT 61.210 131.815 61.380 132.485 ;
        RECT 62.290 132.415 62.535 133.020 ;
        RECT 62.755 132.690 63.265 133.225 ;
        RECT 58.505 130.845 60.535 131.015 ;
        RECT 60.705 130.675 60.875 131.815 ;
        RECT 61.045 130.845 61.380 131.815 ;
        RECT 62.015 132.245 63.245 132.415 ;
        RECT 62.015 131.435 62.355 132.245 ;
        RECT 62.525 131.680 63.275 131.870 ;
        RECT 62.015 131.025 62.530 131.435 ;
        RECT 62.765 130.675 62.935 131.435 ;
        RECT 63.105 131.015 63.275 131.680 ;
        RECT 63.445 131.695 63.635 133.055 ;
        RECT 63.805 132.885 64.080 133.055 ;
        RECT 63.805 132.715 64.085 132.885 ;
        RECT 63.805 131.895 64.080 132.715 ;
        RECT 64.270 132.690 64.800 133.055 ;
        RECT 65.225 132.825 65.555 133.225 ;
        RECT 64.625 132.655 64.800 132.690 ;
        RECT 64.285 131.695 64.455 132.495 ;
        RECT 63.445 131.525 64.455 131.695 ;
        RECT 64.625 132.485 65.555 132.655 ;
        RECT 65.725 132.485 65.980 133.055 ;
        RECT 66.705 132.675 66.875 133.055 ;
        RECT 67.055 132.845 67.385 133.225 ;
        RECT 66.705 132.505 67.370 132.675 ;
        RECT 67.565 132.550 67.825 133.055 ;
        RECT 64.625 131.355 64.795 132.485 ;
        RECT 65.385 132.315 65.555 132.485 ;
        RECT 63.670 131.185 64.795 131.355 ;
        RECT 64.965 131.985 65.160 132.315 ;
        RECT 65.385 131.985 65.640 132.315 ;
        RECT 64.965 131.015 65.135 131.985 ;
        RECT 65.810 131.815 65.980 132.485 ;
        RECT 66.635 131.955 66.965 132.325 ;
        RECT 67.200 132.250 67.370 132.505 ;
        RECT 63.105 130.845 65.135 131.015 ;
        RECT 65.305 130.675 65.475 131.815 ;
        RECT 65.645 130.845 65.980 131.815 ;
        RECT 67.200 131.920 67.485 132.250 ;
        RECT 67.200 131.775 67.370 131.920 ;
        RECT 66.705 131.605 67.370 131.775 ;
        RECT 67.655 131.750 67.825 132.550 ;
        RECT 68.195 132.595 68.525 132.955 ;
        RECT 69.145 132.765 69.395 133.225 ;
        RECT 69.565 132.765 70.125 133.055 ;
        RECT 68.195 132.405 69.585 132.595 ;
        RECT 69.415 132.315 69.585 132.405 ;
        RECT 66.705 130.845 66.875 131.605 ;
        RECT 67.055 130.675 67.385 131.435 ;
        RECT 67.555 130.845 67.825 131.750 ;
        RECT 68.010 131.985 68.685 132.235 ;
        RECT 68.905 131.985 69.245 132.235 ;
        RECT 69.415 131.985 69.705 132.315 ;
        RECT 68.010 131.625 68.275 131.985 ;
        RECT 69.415 131.735 69.585 131.985 ;
        RECT 68.645 131.565 69.585 131.735 ;
        RECT 68.195 130.675 68.475 131.345 ;
        RECT 68.645 131.015 68.945 131.565 ;
        RECT 69.875 131.395 70.125 132.765 ;
        RECT 70.570 132.415 70.815 133.020 ;
        RECT 71.035 132.690 71.545 133.225 ;
        RECT 69.145 130.675 69.475 131.395 ;
        RECT 69.665 130.845 70.125 131.395 ;
        RECT 70.295 132.245 71.525 132.415 ;
        RECT 70.295 131.435 70.635 132.245 ;
        RECT 70.805 131.680 71.555 131.870 ;
        RECT 70.295 131.025 70.810 131.435 ;
        RECT 71.045 130.675 71.215 131.435 ;
        RECT 71.385 131.015 71.555 131.680 ;
        RECT 71.725 131.695 71.915 133.055 ;
        RECT 72.085 132.885 72.360 133.055 ;
        RECT 72.085 132.715 72.365 132.885 ;
        RECT 72.085 131.895 72.360 132.715 ;
        RECT 72.550 132.690 73.080 133.055 ;
        RECT 73.505 132.825 73.835 133.225 ;
        RECT 72.905 132.655 73.080 132.690 ;
        RECT 72.565 131.695 72.735 132.495 ;
        RECT 71.725 131.525 72.735 131.695 ;
        RECT 72.905 132.485 73.835 132.655 ;
        RECT 74.005 132.485 74.260 133.055 ;
        RECT 74.435 132.500 74.725 133.225 ;
        RECT 72.905 131.355 73.075 132.485 ;
        RECT 73.665 132.315 73.835 132.485 ;
        RECT 71.950 131.185 73.075 131.355 ;
        RECT 73.245 131.985 73.440 132.315 ;
        RECT 73.665 131.985 73.920 132.315 ;
        RECT 73.245 131.015 73.415 131.985 ;
        RECT 74.090 131.815 74.260 132.485 ;
        RECT 75.630 132.415 75.875 133.020 ;
        RECT 76.095 132.690 76.605 133.225 ;
        RECT 75.355 132.245 76.585 132.415 ;
        RECT 71.385 130.845 73.415 131.015 ;
        RECT 73.585 130.675 73.755 131.815 ;
        RECT 73.925 130.845 74.260 131.815 ;
        RECT 74.435 130.675 74.725 131.840 ;
        RECT 75.355 131.435 75.695 132.245 ;
        RECT 75.865 131.680 76.615 131.870 ;
        RECT 75.355 131.025 75.870 131.435 ;
        RECT 76.105 130.675 76.275 131.435 ;
        RECT 76.445 131.015 76.615 131.680 ;
        RECT 76.785 131.695 76.975 133.055 ;
        RECT 77.145 132.545 77.420 133.055 ;
        RECT 77.610 132.690 78.140 133.055 ;
        RECT 78.565 132.825 78.895 133.225 ;
        RECT 77.965 132.655 78.140 132.690 ;
        RECT 77.145 132.375 77.425 132.545 ;
        RECT 77.145 131.895 77.420 132.375 ;
        RECT 77.625 131.695 77.795 132.495 ;
        RECT 76.785 131.525 77.795 131.695 ;
        RECT 77.965 132.485 78.895 132.655 ;
        RECT 79.065 132.485 79.320 133.055 ;
        RECT 77.965 131.355 78.135 132.485 ;
        RECT 78.725 132.315 78.895 132.485 ;
        RECT 77.010 131.185 78.135 131.355 ;
        RECT 78.305 131.985 78.500 132.315 ;
        RECT 78.725 131.985 78.980 132.315 ;
        RECT 78.305 131.015 78.475 131.985 ;
        RECT 79.150 131.815 79.320 132.485 ;
        RECT 76.445 130.845 78.475 131.015 ;
        RECT 78.645 130.675 78.815 131.815 ;
        RECT 78.985 130.845 79.320 131.815 ;
        RECT 79.495 132.550 79.755 133.055 ;
        RECT 79.935 132.845 80.265 133.225 ;
        RECT 80.445 132.675 80.615 133.055 ;
        RECT 79.495 131.750 79.665 132.550 ;
        RECT 79.950 132.505 80.615 132.675 ;
        RECT 80.965 132.675 81.135 133.055 ;
        RECT 81.315 132.845 81.645 133.225 ;
        RECT 80.965 132.505 81.630 132.675 ;
        RECT 81.825 132.550 82.085 133.055 ;
        RECT 79.950 132.250 80.120 132.505 ;
        RECT 79.835 131.920 80.120 132.250 ;
        RECT 80.355 131.955 80.685 132.325 ;
        RECT 80.895 131.955 81.225 132.325 ;
        RECT 81.460 132.250 81.630 132.505 ;
        RECT 79.950 131.775 80.120 131.920 ;
        RECT 81.460 131.920 81.745 132.250 ;
        RECT 81.460 131.775 81.630 131.920 ;
        RECT 79.495 130.845 79.765 131.750 ;
        RECT 79.950 131.605 80.615 131.775 ;
        RECT 79.935 130.675 80.265 131.435 ;
        RECT 80.445 130.845 80.615 131.605 ;
        RECT 80.965 131.605 81.630 131.775 ;
        RECT 81.915 131.750 82.085 132.550 ;
        RECT 82.255 132.475 83.465 133.225 ;
        RECT 80.965 130.845 81.135 131.605 ;
        RECT 81.315 130.675 81.645 131.435 ;
        RECT 81.815 130.845 82.085 131.750 ;
        RECT 82.255 131.765 82.775 132.305 ;
        RECT 82.945 131.935 83.465 132.475 ;
        RECT 83.675 132.405 83.905 133.225 ;
        RECT 84.075 132.425 84.405 133.055 ;
        RECT 83.655 131.985 83.985 132.235 ;
        RECT 84.155 131.825 84.405 132.425 ;
        RECT 84.575 132.405 84.785 133.225 ;
        RECT 85.390 132.515 85.645 133.045 ;
        RECT 85.825 132.765 86.110 133.225 ;
        RECT 82.255 130.675 83.465 131.765 ;
        RECT 83.675 130.675 83.905 131.815 ;
        RECT 84.075 130.845 84.405 131.825 ;
        RECT 84.575 130.675 84.785 131.815 ;
        RECT 85.390 131.655 85.570 132.515 ;
        RECT 86.290 132.315 86.540 132.965 ;
        RECT 85.740 131.985 86.540 132.315 ;
        RECT 85.390 131.525 85.645 131.655 ;
        RECT 85.305 131.355 85.645 131.525 ;
        RECT 85.390 130.985 85.645 131.355 ;
        RECT 85.825 130.675 86.110 131.475 ;
        RECT 86.290 131.395 86.540 131.985 ;
        RECT 86.740 132.630 87.060 132.960 ;
        RECT 87.240 132.745 87.900 133.225 ;
        RECT 88.100 132.835 88.950 133.005 ;
        RECT 86.740 131.735 86.930 132.630 ;
        RECT 87.250 132.305 87.910 132.575 ;
        RECT 87.580 132.245 87.910 132.305 ;
        RECT 87.100 132.075 87.430 132.135 ;
        RECT 88.100 132.075 88.270 132.835 ;
        RECT 89.510 132.765 89.830 133.225 ;
        RECT 90.030 132.585 90.280 133.015 ;
        RECT 90.570 132.785 90.980 133.225 ;
        RECT 91.150 132.845 92.165 133.045 ;
        RECT 88.440 132.415 89.690 132.585 ;
        RECT 88.440 132.295 88.770 132.415 ;
        RECT 87.100 131.905 89.000 132.075 ;
        RECT 86.740 131.565 88.660 131.735 ;
        RECT 86.740 131.545 87.060 131.565 ;
        RECT 86.290 130.885 86.620 131.395 ;
        RECT 86.890 130.935 87.060 131.545 ;
        RECT 88.830 131.395 89.000 131.905 ;
        RECT 89.170 131.835 89.350 132.245 ;
        RECT 89.520 131.655 89.690 132.415 ;
        RECT 87.230 130.675 87.560 131.365 ;
        RECT 87.790 131.225 89.000 131.395 ;
        RECT 89.170 131.345 89.690 131.655 ;
        RECT 89.860 132.245 90.280 132.585 ;
        RECT 90.570 132.245 90.980 132.575 ;
        RECT 89.860 131.475 90.050 132.245 ;
        RECT 91.150 132.115 91.320 132.845 ;
        RECT 92.465 132.675 92.635 133.005 ;
        RECT 92.805 132.845 93.135 133.225 ;
        RECT 91.490 132.295 91.840 132.665 ;
        RECT 91.150 132.075 91.570 132.115 ;
        RECT 90.220 131.905 91.570 132.075 ;
        RECT 90.220 131.745 90.470 131.905 ;
        RECT 90.980 131.475 91.230 131.735 ;
        RECT 89.860 131.225 91.230 131.475 ;
        RECT 87.790 130.935 88.030 131.225 ;
        RECT 88.830 131.145 89.000 131.225 ;
        RECT 88.230 130.675 88.650 131.055 ;
        RECT 88.830 130.895 89.460 131.145 ;
        RECT 89.930 130.675 90.260 131.055 ;
        RECT 90.430 130.935 90.600 131.225 ;
        RECT 91.400 131.060 91.570 131.905 ;
        RECT 92.020 131.735 92.240 132.605 ;
        RECT 92.465 132.485 93.160 132.675 ;
        RECT 91.740 131.355 92.240 131.735 ;
        RECT 92.410 131.685 92.820 132.305 ;
        RECT 92.990 131.515 93.160 132.485 ;
        RECT 92.465 131.345 93.160 131.515 ;
        RECT 90.780 130.675 91.160 131.055 ;
        RECT 91.400 130.890 92.230 131.060 ;
        RECT 92.465 130.845 92.635 131.345 ;
        RECT 92.805 130.675 93.135 131.175 ;
        RECT 93.350 130.845 93.575 132.965 ;
        RECT 93.745 132.845 94.075 133.225 ;
        RECT 94.245 132.675 94.415 132.965 ;
        RECT 93.750 132.505 94.415 132.675 ;
        RECT 93.750 131.515 93.980 132.505 ;
        RECT 94.715 132.405 94.945 133.225 ;
        RECT 95.115 132.425 95.445 133.055 ;
        RECT 94.150 131.685 94.500 132.335 ;
        RECT 94.695 131.985 95.025 132.235 ;
        RECT 95.195 131.825 95.445 132.425 ;
        RECT 95.615 132.405 95.825 133.225 ;
        RECT 96.330 132.415 96.575 133.020 ;
        RECT 96.795 132.690 97.305 133.225 ;
        RECT 93.750 131.345 94.415 131.515 ;
        RECT 93.745 130.675 94.075 131.175 ;
        RECT 94.245 130.845 94.415 131.345 ;
        RECT 94.715 130.675 94.945 131.815 ;
        RECT 95.115 130.845 95.445 131.825 ;
        RECT 96.055 132.245 97.285 132.415 ;
        RECT 95.615 130.675 95.825 131.815 ;
        RECT 96.055 131.435 96.395 132.245 ;
        RECT 96.565 131.680 97.315 131.870 ;
        RECT 96.055 131.025 96.570 131.435 ;
        RECT 96.805 130.675 96.975 131.435 ;
        RECT 97.145 131.015 97.315 131.680 ;
        RECT 97.485 131.695 97.675 133.055 ;
        RECT 97.845 132.885 98.120 133.055 ;
        RECT 97.845 132.715 98.125 132.885 ;
        RECT 97.845 131.895 98.120 132.715 ;
        RECT 98.310 132.690 98.840 133.055 ;
        RECT 99.265 132.825 99.595 133.225 ;
        RECT 98.665 132.655 98.840 132.690 ;
        RECT 98.325 131.695 98.495 132.495 ;
        RECT 97.485 131.525 98.495 131.695 ;
        RECT 98.665 132.485 99.595 132.655 ;
        RECT 99.765 132.485 100.020 133.055 ;
        RECT 100.195 132.500 100.485 133.225 ;
        RECT 101.030 132.515 101.285 133.045 ;
        RECT 101.465 132.765 101.750 133.225 ;
        RECT 98.665 131.355 98.835 132.485 ;
        RECT 99.425 132.315 99.595 132.485 ;
        RECT 97.710 131.185 98.835 131.355 ;
        RECT 99.005 131.985 99.200 132.315 ;
        RECT 99.425 131.985 99.680 132.315 ;
        RECT 99.005 131.015 99.175 131.985 ;
        RECT 99.850 131.815 100.020 132.485 ;
        RECT 101.030 131.865 101.210 132.515 ;
        RECT 101.930 132.315 102.180 132.965 ;
        RECT 101.380 131.985 102.180 132.315 ;
        RECT 97.145 130.845 99.175 131.015 ;
        RECT 99.345 130.675 99.515 131.815 ;
        RECT 99.685 130.845 100.020 131.815 ;
        RECT 100.195 130.675 100.485 131.840 ;
        RECT 100.945 131.695 101.210 131.865 ;
        RECT 101.030 131.655 101.210 131.695 ;
        RECT 101.030 130.985 101.285 131.655 ;
        RECT 101.465 130.675 101.750 131.475 ;
        RECT 101.930 131.395 102.180 131.985 ;
        RECT 102.380 132.630 102.700 132.960 ;
        RECT 102.880 132.745 103.540 133.225 ;
        RECT 103.740 132.835 104.590 133.005 ;
        RECT 102.380 131.735 102.570 132.630 ;
        RECT 102.890 132.305 103.550 132.575 ;
        RECT 103.220 132.245 103.550 132.305 ;
        RECT 102.740 132.075 103.070 132.135 ;
        RECT 103.740 132.075 103.910 132.835 ;
        RECT 105.150 132.765 105.470 133.225 ;
        RECT 105.670 132.585 105.920 133.015 ;
        RECT 106.210 132.785 106.620 133.225 ;
        RECT 106.790 132.845 107.805 133.045 ;
        RECT 104.080 132.415 105.330 132.585 ;
        RECT 104.080 132.295 104.410 132.415 ;
        RECT 102.740 131.905 104.640 132.075 ;
        RECT 102.380 131.565 104.300 131.735 ;
        RECT 102.380 131.545 102.700 131.565 ;
        RECT 101.930 130.885 102.260 131.395 ;
        RECT 102.530 130.935 102.700 131.545 ;
        RECT 104.470 131.395 104.640 131.905 ;
        RECT 104.810 131.835 104.990 132.245 ;
        RECT 105.160 131.655 105.330 132.415 ;
        RECT 102.870 130.675 103.200 131.365 ;
        RECT 103.430 131.225 104.640 131.395 ;
        RECT 104.810 131.345 105.330 131.655 ;
        RECT 105.500 132.245 105.920 132.585 ;
        RECT 106.210 132.245 106.620 132.575 ;
        RECT 105.500 131.475 105.690 132.245 ;
        RECT 106.790 132.115 106.960 132.845 ;
        RECT 108.105 132.675 108.275 133.005 ;
        RECT 108.445 132.845 108.775 133.225 ;
        RECT 107.130 132.295 107.480 132.665 ;
        RECT 106.790 132.075 107.210 132.115 ;
        RECT 105.860 131.905 107.210 132.075 ;
        RECT 105.860 131.745 106.110 131.905 ;
        RECT 106.620 131.475 106.870 131.735 ;
        RECT 105.500 131.225 106.870 131.475 ;
        RECT 103.430 130.935 103.670 131.225 ;
        RECT 104.470 131.145 104.640 131.225 ;
        RECT 103.870 130.675 104.290 131.055 ;
        RECT 104.470 130.895 105.100 131.145 ;
        RECT 105.570 130.675 105.900 131.055 ;
        RECT 106.070 130.935 106.240 131.225 ;
        RECT 107.040 131.060 107.210 131.905 ;
        RECT 107.660 131.735 107.880 132.605 ;
        RECT 108.105 132.485 108.800 132.675 ;
        RECT 107.380 131.355 107.880 131.735 ;
        RECT 108.050 131.685 108.460 132.305 ;
        RECT 108.630 131.515 108.800 132.485 ;
        RECT 108.105 131.345 108.800 131.515 ;
        RECT 106.420 130.675 106.800 131.055 ;
        RECT 107.040 130.890 107.870 131.060 ;
        RECT 108.105 130.845 108.275 131.345 ;
        RECT 108.445 130.675 108.775 131.175 ;
        RECT 108.990 130.845 109.215 132.965 ;
        RECT 109.385 132.845 109.715 133.225 ;
        RECT 109.885 132.675 110.055 132.965 ;
        RECT 109.390 132.505 110.055 132.675 ;
        RECT 109.390 131.515 109.620 132.505 ;
        RECT 110.315 132.455 111.985 133.225 ;
        RECT 112.155 132.475 113.365 133.225 ;
        RECT 109.790 131.685 110.140 132.335 ;
        RECT 110.315 131.765 111.065 132.285 ;
        RECT 111.235 131.935 111.985 132.455 ;
        RECT 112.155 131.765 112.675 132.305 ;
        RECT 112.845 131.935 113.365 132.475 ;
        RECT 109.390 131.345 110.055 131.515 ;
        RECT 109.385 130.675 109.715 131.175 ;
        RECT 109.885 130.845 110.055 131.345 ;
        RECT 110.315 130.675 111.985 131.765 ;
        RECT 112.155 130.675 113.365 131.765 ;
        RECT 22.830 130.505 113.450 130.675 ;
        RECT 22.915 129.415 24.125 130.505 ;
        RECT 25.305 129.835 25.475 130.335 ;
        RECT 25.645 130.005 25.975 130.505 ;
        RECT 25.305 129.665 25.970 129.835 ;
        RECT 22.915 128.705 23.435 129.245 ;
        RECT 23.605 128.875 24.125 129.415 ;
        RECT 25.220 128.845 25.570 129.495 ;
        RECT 22.915 127.955 24.125 128.705 ;
        RECT 25.740 128.675 25.970 129.665 ;
        RECT 25.305 128.505 25.970 128.675 ;
        RECT 25.305 128.215 25.475 128.505 ;
        RECT 25.645 127.955 25.975 128.335 ;
        RECT 26.145 128.215 26.370 130.335 ;
        RECT 26.585 130.005 26.915 130.505 ;
        RECT 27.085 129.835 27.255 130.335 ;
        RECT 27.490 130.120 28.320 130.290 ;
        RECT 28.560 130.125 28.940 130.505 ;
        RECT 26.560 129.665 27.255 129.835 ;
        RECT 26.560 128.695 26.730 129.665 ;
        RECT 26.900 128.875 27.310 129.495 ;
        RECT 27.480 129.445 27.980 129.825 ;
        RECT 26.560 128.505 27.255 128.695 ;
        RECT 27.480 128.575 27.700 129.445 ;
        RECT 28.150 129.275 28.320 130.120 ;
        RECT 29.120 129.955 29.290 130.245 ;
        RECT 29.460 130.125 29.790 130.505 ;
        RECT 30.260 130.035 30.890 130.285 ;
        RECT 31.070 130.125 31.490 130.505 ;
        RECT 30.720 129.955 30.890 130.035 ;
        RECT 31.690 129.955 31.930 130.245 ;
        RECT 28.490 129.705 29.860 129.955 ;
        RECT 28.490 129.445 28.740 129.705 ;
        RECT 29.250 129.275 29.500 129.435 ;
        RECT 28.150 129.105 29.500 129.275 ;
        RECT 28.150 129.065 28.570 129.105 ;
        RECT 27.880 128.515 28.230 128.885 ;
        RECT 26.585 127.955 26.915 128.335 ;
        RECT 27.085 128.175 27.255 128.505 ;
        RECT 28.400 128.335 28.570 129.065 ;
        RECT 29.670 128.935 29.860 129.705 ;
        RECT 28.740 128.605 29.150 128.935 ;
        RECT 29.440 128.595 29.860 128.935 ;
        RECT 30.030 129.525 30.550 129.835 ;
        RECT 30.720 129.785 31.930 129.955 ;
        RECT 32.160 129.815 32.490 130.505 ;
        RECT 30.030 128.765 30.200 129.525 ;
        RECT 30.370 128.935 30.550 129.345 ;
        RECT 30.720 129.275 30.890 129.785 ;
        RECT 32.660 129.635 32.830 130.245 ;
        RECT 33.100 129.785 33.430 130.295 ;
        RECT 32.660 129.615 32.980 129.635 ;
        RECT 31.060 129.445 32.980 129.615 ;
        RECT 30.720 129.105 32.620 129.275 ;
        RECT 30.950 128.765 31.280 128.885 ;
        RECT 30.030 128.595 31.280 128.765 ;
        RECT 27.555 128.135 28.570 128.335 ;
        RECT 28.740 127.955 29.150 128.395 ;
        RECT 29.440 128.165 29.690 128.595 ;
        RECT 29.890 127.955 30.210 128.415 ;
        RECT 31.450 128.345 31.620 129.105 ;
        RECT 32.290 129.045 32.620 129.105 ;
        RECT 31.810 128.875 32.140 128.935 ;
        RECT 31.810 128.605 32.470 128.875 ;
        RECT 32.790 128.550 32.980 129.445 ;
        RECT 30.770 128.175 31.620 128.345 ;
        RECT 31.820 127.955 32.480 128.435 ;
        RECT 32.660 128.220 32.980 128.550 ;
        RECT 33.180 129.195 33.430 129.785 ;
        RECT 33.610 129.705 33.895 130.505 ;
        RECT 34.075 129.525 34.330 130.195 ;
        RECT 33.180 128.865 33.980 129.195 ;
        RECT 33.180 128.215 33.430 128.865 ;
        RECT 34.150 128.805 34.330 129.525 ;
        RECT 35.795 129.340 36.085 130.505 ;
        RECT 37.175 129.430 37.445 130.335 ;
        RECT 37.615 129.745 37.945 130.505 ;
        RECT 38.125 129.575 38.295 130.335 ;
        RECT 39.105 129.835 39.275 130.335 ;
        RECT 39.445 130.005 39.775 130.505 ;
        RECT 39.105 129.665 39.770 129.835 ;
        RECT 34.150 128.665 34.415 128.805 ;
        RECT 34.075 128.635 34.415 128.665 ;
        RECT 33.610 127.955 33.895 128.415 ;
        RECT 34.075 128.135 34.330 128.635 ;
        RECT 35.795 127.955 36.085 128.680 ;
        RECT 37.175 128.630 37.345 129.430 ;
        RECT 37.630 129.405 38.295 129.575 ;
        RECT 37.630 129.260 37.800 129.405 ;
        RECT 37.515 128.930 37.800 129.260 ;
        RECT 37.630 128.675 37.800 128.930 ;
        RECT 38.035 128.855 38.365 129.225 ;
        RECT 39.020 128.845 39.370 129.495 ;
        RECT 39.540 128.675 39.770 129.665 ;
        RECT 37.175 128.125 37.435 128.630 ;
        RECT 37.630 128.505 38.295 128.675 ;
        RECT 37.615 127.955 37.945 128.335 ;
        RECT 38.125 128.125 38.295 128.505 ;
        RECT 39.105 128.505 39.770 128.675 ;
        RECT 39.105 128.215 39.275 128.505 ;
        RECT 39.445 127.955 39.775 128.335 ;
        RECT 39.945 128.215 40.170 130.335 ;
        RECT 40.385 130.005 40.715 130.505 ;
        RECT 40.885 129.835 41.055 130.335 ;
        RECT 41.290 130.120 42.120 130.290 ;
        RECT 42.360 130.125 42.740 130.505 ;
        RECT 40.360 129.665 41.055 129.835 ;
        RECT 40.360 128.695 40.530 129.665 ;
        RECT 40.700 128.875 41.110 129.495 ;
        RECT 41.280 129.445 41.780 129.825 ;
        RECT 40.360 128.505 41.055 128.695 ;
        RECT 41.280 128.575 41.500 129.445 ;
        RECT 41.950 129.275 42.120 130.120 ;
        RECT 42.920 129.955 43.090 130.245 ;
        RECT 43.260 130.125 43.590 130.505 ;
        RECT 44.060 130.035 44.690 130.285 ;
        RECT 44.870 130.125 45.290 130.505 ;
        RECT 44.520 129.955 44.690 130.035 ;
        RECT 45.490 129.955 45.730 130.245 ;
        RECT 42.290 129.705 43.660 129.955 ;
        RECT 42.290 129.445 42.540 129.705 ;
        RECT 43.050 129.275 43.300 129.435 ;
        RECT 41.950 129.105 43.300 129.275 ;
        RECT 41.950 129.065 42.370 129.105 ;
        RECT 41.680 128.515 42.030 128.885 ;
        RECT 40.385 127.955 40.715 128.335 ;
        RECT 40.885 128.175 41.055 128.505 ;
        RECT 42.200 128.335 42.370 129.065 ;
        RECT 43.470 128.935 43.660 129.705 ;
        RECT 42.540 128.605 42.950 128.935 ;
        RECT 43.240 128.595 43.660 128.935 ;
        RECT 43.830 129.525 44.350 129.835 ;
        RECT 44.520 129.785 45.730 129.955 ;
        RECT 45.960 129.815 46.290 130.505 ;
        RECT 43.830 128.765 44.000 129.525 ;
        RECT 44.170 128.935 44.350 129.345 ;
        RECT 44.520 129.275 44.690 129.785 ;
        RECT 46.460 129.635 46.630 130.245 ;
        RECT 46.900 129.785 47.230 130.295 ;
        RECT 46.460 129.615 46.780 129.635 ;
        RECT 44.860 129.445 46.780 129.615 ;
        RECT 44.520 129.105 46.420 129.275 ;
        RECT 44.750 128.765 45.080 128.885 ;
        RECT 43.830 128.595 45.080 128.765 ;
        RECT 41.355 128.135 42.370 128.335 ;
        RECT 42.540 127.955 42.950 128.395 ;
        RECT 43.240 128.165 43.490 128.595 ;
        RECT 43.690 127.955 44.010 128.415 ;
        RECT 45.250 128.345 45.420 129.105 ;
        RECT 46.090 129.045 46.420 129.105 ;
        RECT 45.610 128.875 45.940 128.935 ;
        RECT 45.610 128.605 46.270 128.875 ;
        RECT 46.590 128.550 46.780 129.445 ;
        RECT 44.570 128.175 45.420 128.345 ;
        RECT 45.620 127.955 46.280 128.435 ;
        RECT 46.460 128.220 46.780 128.550 ;
        RECT 46.980 129.195 47.230 129.785 ;
        RECT 47.410 129.705 47.695 130.505 ;
        RECT 47.875 130.165 48.130 130.195 ;
        RECT 47.875 129.995 48.215 130.165 ;
        RECT 47.875 129.525 48.130 129.995 ;
        RECT 46.980 128.865 47.780 129.195 ;
        RECT 46.980 128.215 47.230 128.865 ;
        RECT 47.950 128.665 48.130 129.525 ;
        RECT 47.410 127.955 47.695 128.415 ;
        RECT 47.875 128.135 48.130 128.665 ;
        RECT 49.135 129.785 49.595 130.335 ;
        RECT 49.785 129.785 50.115 130.505 ;
        RECT 49.135 128.415 49.385 129.785 ;
        RECT 50.315 129.615 50.615 130.165 ;
        RECT 50.785 129.835 51.065 130.505 ;
        RECT 52.270 130.165 52.525 130.195 ;
        RECT 52.185 129.995 52.525 130.165 ;
        RECT 49.675 129.445 50.615 129.615 ;
        RECT 49.675 129.195 49.845 129.445 ;
        RECT 50.985 129.195 51.250 129.555 ;
        RECT 49.555 128.865 49.845 129.195 ;
        RECT 50.015 128.945 50.355 129.195 ;
        RECT 50.575 128.945 51.250 129.195 ;
        RECT 52.270 129.525 52.525 129.995 ;
        RECT 52.705 129.705 52.990 130.505 ;
        RECT 53.170 129.785 53.500 130.295 ;
        RECT 49.675 128.775 49.845 128.865 ;
        RECT 49.675 128.585 51.065 128.775 ;
        RECT 49.135 128.125 49.695 128.415 ;
        RECT 49.865 127.955 50.115 128.415 ;
        RECT 50.735 128.225 51.065 128.585 ;
        RECT 52.270 128.665 52.450 129.525 ;
        RECT 53.170 129.195 53.420 129.785 ;
        RECT 53.770 129.635 53.940 130.245 ;
        RECT 54.110 129.815 54.440 130.505 ;
        RECT 54.670 129.955 54.910 130.245 ;
        RECT 55.110 130.125 55.530 130.505 ;
        RECT 55.710 130.035 56.340 130.285 ;
        RECT 56.810 130.125 57.140 130.505 ;
        RECT 55.710 129.955 55.880 130.035 ;
        RECT 57.310 129.955 57.480 130.245 ;
        RECT 57.660 130.125 58.040 130.505 ;
        RECT 58.280 130.120 59.110 130.290 ;
        RECT 54.670 129.785 55.880 129.955 ;
        RECT 52.620 128.865 53.420 129.195 ;
        RECT 52.270 128.135 52.525 128.665 ;
        RECT 52.705 127.955 52.990 128.415 ;
        RECT 53.170 128.215 53.420 128.865 ;
        RECT 53.620 129.615 53.940 129.635 ;
        RECT 53.620 129.445 55.540 129.615 ;
        RECT 53.620 128.550 53.810 129.445 ;
        RECT 55.710 129.275 55.880 129.785 ;
        RECT 56.050 129.525 56.570 129.835 ;
        RECT 53.980 129.105 55.880 129.275 ;
        RECT 53.980 129.045 54.310 129.105 ;
        RECT 54.460 128.875 54.790 128.935 ;
        RECT 54.130 128.605 54.790 128.875 ;
        RECT 53.620 128.220 53.940 128.550 ;
        RECT 54.120 127.955 54.780 128.435 ;
        RECT 54.980 128.345 55.150 129.105 ;
        RECT 56.050 128.935 56.230 129.345 ;
        RECT 55.320 128.765 55.650 128.885 ;
        RECT 56.400 128.765 56.570 129.525 ;
        RECT 55.320 128.595 56.570 128.765 ;
        RECT 56.740 129.705 58.110 129.955 ;
        RECT 56.740 128.935 56.930 129.705 ;
        RECT 57.860 129.445 58.110 129.705 ;
        RECT 57.100 129.275 57.350 129.435 ;
        RECT 58.280 129.275 58.450 130.120 ;
        RECT 59.345 129.835 59.515 130.335 ;
        RECT 59.685 130.005 60.015 130.505 ;
        RECT 58.620 129.445 59.120 129.825 ;
        RECT 59.345 129.665 60.040 129.835 ;
        RECT 57.100 129.105 58.450 129.275 ;
        RECT 58.030 129.065 58.450 129.105 ;
        RECT 56.740 128.595 57.160 128.935 ;
        RECT 57.450 128.605 57.860 128.935 ;
        RECT 54.980 128.175 55.830 128.345 ;
        RECT 56.390 127.955 56.710 128.415 ;
        RECT 56.910 128.165 57.160 128.595 ;
        RECT 57.450 127.955 57.860 128.395 ;
        RECT 58.030 128.335 58.200 129.065 ;
        RECT 58.370 128.515 58.720 128.885 ;
        RECT 58.900 128.575 59.120 129.445 ;
        RECT 59.290 128.875 59.700 129.495 ;
        RECT 59.870 128.695 60.040 129.665 ;
        RECT 59.345 128.505 60.040 128.695 ;
        RECT 58.030 128.135 59.045 128.335 ;
        RECT 59.345 128.175 59.515 128.505 ;
        RECT 59.685 127.955 60.015 128.335 ;
        RECT 60.230 128.215 60.455 130.335 ;
        RECT 60.625 130.005 60.955 130.505 ;
        RECT 61.125 129.835 61.295 130.335 ;
        RECT 60.630 129.665 61.295 129.835 ;
        RECT 60.630 128.675 60.860 129.665 ;
        RECT 61.030 128.845 61.380 129.495 ;
        RECT 61.555 129.340 61.845 130.505 ;
        RECT 62.390 130.165 62.645 130.195 ;
        RECT 62.305 129.995 62.645 130.165 ;
        RECT 62.390 129.525 62.645 129.995 ;
        RECT 62.825 129.705 63.110 130.505 ;
        RECT 63.290 129.785 63.620 130.295 ;
        RECT 60.630 128.505 61.295 128.675 ;
        RECT 60.625 127.955 60.955 128.335 ;
        RECT 61.125 128.215 61.295 128.505 ;
        RECT 61.555 127.955 61.845 128.680 ;
        RECT 62.390 128.665 62.570 129.525 ;
        RECT 63.290 129.195 63.540 129.785 ;
        RECT 63.890 129.635 64.060 130.245 ;
        RECT 64.230 129.815 64.560 130.505 ;
        RECT 64.790 129.955 65.030 130.245 ;
        RECT 65.230 130.125 65.650 130.505 ;
        RECT 65.830 130.035 66.460 130.285 ;
        RECT 66.930 130.125 67.260 130.505 ;
        RECT 65.830 129.955 66.000 130.035 ;
        RECT 67.430 129.955 67.600 130.245 ;
        RECT 67.780 130.125 68.160 130.505 ;
        RECT 68.400 130.120 69.230 130.290 ;
        RECT 64.790 129.785 66.000 129.955 ;
        RECT 62.740 128.865 63.540 129.195 ;
        RECT 62.390 128.135 62.645 128.665 ;
        RECT 62.825 127.955 63.110 128.415 ;
        RECT 63.290 128.215 63.540 128.865 ;
        RECT 63.740 129.615 64.060 129.635 ;
        RECT 63.740 129.445 65.660 129.615 ;
        RECT 63.740 128.550 63.930 129.445 ;
        RECT 65.830 129.275 66.000 129.785 ;
        RECT 66.170 129.525 66.690 129.835 ;
        RECT 64.100 129.105 66.000 129.275 ;
        RECT 64.100 129.045 64.430 129.105 ;
        RECT 64.580 128.875 64.910 128.935 ;
        RECT 64.250 128.605 64.910 128.875 ;
        RECT 63.740 128.220 64.060 128.550 ;
        RECT 64.240 127.955 64.900 128.435 ;
        RECT 65.100 128.345 65.270 129.105 ;
        RECT 66.170 128.935 66.350 129.345 ;
        RECT 65.440 128.765 65.770 128.885 ;
        RECT 66.520 128.765 66.690 129.525 ;
        RECT 65.440 128.595 66.690 128.765 ;
        RECT 66.860 129.705 68.230 129.955 ;
        RECT 66.860 128.935 67.050 129.705 ;
        RECT 67.980 129.445 68.230 129.705 ;
        RECT 67.220 129.275 67.470 129.435 ;
        RECT 68.400 129.275 68.570 130.120 ;
        RECT 69.465 129.835 69.635 130.335 ;
        RECT 69.805 130.005 70.135 130.505 ;
        RECT 68.740 129.445 69.240 129.825 ;
        RECT 69.465 129.665 70.160 129.835 ;
        RECT 67.220 129.105 68.570 129.275 ;
        RECT 68.150 129.065 68.570 129.105 ;
        RECT 66.860 128.595 67.280 128.935 ;
        RECT 67.570 128.605 67.980 128.935 ;
        RECT 65.100 128.175 65.950 128.345 ;
        RECT 66.510 127.955 66.830 128.415 ;
        RECT 67.030 128.165 67.280 128.595 ;
        RECT 67.570 127.955 67.980 128.395 ;
        RECT 68.150 128.335 68.320 129.065 ;
        RECT 68.490 128.515 68.840 128.885 ;
        RECT 69.020 128.575 69.240 129.445 ;
        RECT 69.410 128.875 69.820 129.495 ;
        RECT 69.990 128.695 70.160 129.665 ;
        RECT 69.465 128.505 70.160 128.695 ;
        RECT 68.150 128.135 69.165 128.335 ;
        RECT 69.465 128.175 69.635 128.505 ;
        RECT 69.805 127.955 70.135 128.335 ;
        RECT 70.350 128.215 70.575 130.335 ;
        RECT 70.745 130.005 71.075 130.505 ;
        RECT 71.245 129.835 71.415 130.335 ;
        RECT 70.750 129.665 71.415 129.835 ;
        RECT 72.050 129.825 72.305 130.195 ;
        RECT 70.750 128.675 70.980 129.665 ;
        RECT 71.965 129.655 72.305 129.825 ;
        RECT 72.485 129.705 72.770 130.505 ;
        RECT 72.950 129.785 73.280 130.295 ;
        RECT 72.050 129.525 72.305 129.655 ;
        RECT 71.150 128.845 71.500 129.495 ;
        RECT 70.750 128.505 71.415 128.675 ;
        RECT 70.745 127.955 71.075 128.335 ;
        RECT 71.245 128.215 71.415 128.505 ;
        RECT 72.050 128.665 72.230 129.525 ;
        RECT 72.950 129.195 73.200 129.785 ;
        RECT 73.550 129.635 73.720 130.245 ;
        RECT 73.890 129.815 74.220 130.505 ;
        RECT 74.450 129.955 74.690 130.245 ;
        RECT 74.890 130.125 75.310 130.505 ;
        RECT 75.490 130.035 76.120 130.285 ;
        RECT 76.590 130.125 76.920 130.505 ;
        RECT 75.490 129.955 75.660 130.035 ;
        RECT 77.090 129.955 77.260 130.245 ;
        RECT 77.440 130.125 77.820 130.505 ;
        RECT 78.060 130.120 78.890 130.290 ;
        RECT 74.450 129.785 75.660 129.955 ;
        RECT 72.400 128.865 73.200 129.195 ;
        RECT 72.050 128.135 72.305 128.665 ;
        RECT 72.485 127.955 72.770 128.415 ;
        RECT 72.950 128.215 73.200 128.865 ;
        RECT 73.400 129.615 73.720 129.635 ;
        RECT 73.400 129.445 75.320 129.615 ;
        RECT 73.400 128.550 73.590 129.445 ;
        RECT 75.490 129.275 75.660 129.785 ;
        RECT 75.830 129.525 76.350 129.835 ;
        RECT 73.760 129.105 75.660 129.275 ;
        RECT 73.760 129.045 74.090 129.105 ;
        RECT 74.240 128.875 74.570 128.935 ;
        RECT 73.910 128.605 74.570 128.875 ;
        RECT 73.400 128.220 73.720 128.550 ;
        RECT 73.900 127.955 74.560 128.435 ;
        RECT 74.760 128.345 74.930 129.105 ;
        RECT 75.830 128.935 76.010 129.345 ;
        RECT 75.100 128.765 75.430 128.885 ;
        RECT 76.180 128.765 76.350 129.525 ;
        RECT 75.100 128.595 76.350 128.765 ;
        RECT 76.520 129.705 77.890 129.955 ;
        RECT 76.520 128.935 76.710 129.705 ;
        RECT 77.640 129.445 77.890 129.705 ;
        RECT 76.880 129.275 77.130 129.435 ;
        RECT 78.060 129.275 78.230 130.120 ;
        RECT 79.125 129.835 79.295 130.335 ;
        RECT 79.465 130.005 79.795 130.505 ;
        RECT 78.400 129.445 78.900 129.825 ;
        RECT 79.125 129.665 79.820 129.835 ;
        RECT 76.880 129.105 78.230 129.275 ;
        RECT 77.810 129.065 78.230 129.105 ;
        RECT 76.520 128.595 76.940 128.935 ;
        RECT 77.230 128.605 77.640 128.935 ;
        RECT 74.760 128.175 75.610 128.345 ;
        RECT 76.170 127.955 76.490 128.415 ;
        RECT 76.690 128.165 76.940 128.595 ;
        RECT 77.230 127.955 77.640 128.395 ;
        RECT 77.810 128.335 77.980 129.065 ;
        RECT 78.150 128.515 78.500 128.885 ;
        RECT 78.680 128.575 78.900 129.445 ;
        RECT 79.070 128.875 79.480 129.495 ;
        RECT 79.650 128.695 79.820 129.665 ;
        RECT 79.125 128.505 79.820 128.695 ;
        RECT 77.810 128.135 78.825 128.335 ;
        RECT 79.125 128.175 79.295 128.505 ;
        RECT 79.465 127.955 79.795 128.335 ;
        RECT 80.010 128.215 80.235 130.335 ;
        RECT 80.405 130.005 80.735 130.505 ;
        RECT 80.905 129.835 81.075 130.335 ;
        RECT 80.410 129.665 81.075 129.835 ;
        RECT 80.410 128.675 80.640 129.665 ;
        RECT 80.810 128.845 81.160 129.495 ;
        RECT 81.395 129.365 81.605 130.505 ;
        RECT 81.775 129.355 82.105 130.335 ;
        RECT 82.275 129.365 82.505 130.505 ;
        RECT 83.175 129.745 83.690 130.155 ;
        RECT 83.925 129.745 84.095 130.505 ;
        RECT 84.265 130.165 86.295 130.335 ;
        RECT 80.410 128.505 81.075 128.675 ;
        RECT 80.405 127.955 80.735 128.335 ;
        RECT 80.905 128.215 81.075 128.505 ;
        RECT 81.395 127.955 81.605 128.775 ;
        RECT 81.775 128.755 82.025 129.355 ;
        RECT 82.195 128.945 82.525 129.195 ;
        RECT 83.175 128.935 83.515 129.745 ;
        RECT 84.265 129.500 84.435 130.165 ;
        RECT 84.830 129.825 85.955 129.995 ;
        RECT 83.685 129.310 84.435 129.500 ;
        RECT 84.605 129.485 85.615 129.655 ;
        RECT 81.775 128.125 82.105 128.755 ;
        RECT 82.275 127.955 82.505 128.775 ;
        RECT 83.175 128.765 84.405 128.935 ;
        RECT 83.450 128.160 83.695 128.765 ;
        RECT 83.915 127.955 84.425 128.490 ;
        RECT 84.605 128.125 84.795 129.485 ;
        RECT 84.965 128.465 85.240 129.285 ;
        RECT 85.445 128.685 85.615 129.485 ;
        RECT 85.785 128.695 85.955 129.825 ;
        RECT 86.125 129.195 86.295 130.165 ;
        RECT 86.465 129.365 86.635 130.505 ;
        RECT 86.805 129.365 87.140 130.335 ;
        RECT 86.125 128.865 86.320 129.195 ;
        RECT 86.545 128.865 86.800 129.195 ;
        RECT 86.545 128.695 86.715 128.865 ;
        RECT 86.970 128.695 87.140 129.365 ;
        RECT 87.315 129.340 87.605 130.505 ;
        RECT 87.815 129.365 88.045 130.505 ;
        RECT 88.215 129.355 88.545 130.335 ;
        RECT 88.715 129.365 88.925 130.505 ;
        RECT 89.245 129.575 89.415 130.335 ;
        RECT 89.595 129.745 89.925 130.505 ;
        RECT 89.245 129.405 89.910 129.575 ;
        RECT 90.095 129.430 90.365 130.335 ;
        RECT 87.795 128.945 88.125 129.195 ;
        RECT 85.785 128.525 86.715 128.695 ;
        RECT 85.785 128.490 85.960 128.525 ;
        RECT 84.965 128.295 85.245 128.465 ;
        RECT 84.965 128.125 85.240 128.295 ;
        RECT 85.430 128.125 85.960 128.490 ;
        RECT 86.385 127.955 86.715 128.355 ;
        RECT 86.885 128.125 87.140 128.695 ;
        RECT 87.315 127.955 87.605 128.680 ;
        RECT 87.815 127.955 88.045 128.775 ;
        RECT 88.295 128.755 88.545 129.355 ;
        RECT 89.740 129.260 89.910 129.405 ;
        RECT 89.175 128.855 89.505 129.225 ;
        RECT 89.740 128.930 90.025 129.260 ;
        RECT 88.215 128.125 88.545 128.755 ;
        RECT 88.715 127.955 88.925 128.775 ;
        RECT 89.740 128.675 89.910 128.930 ;
        RECT 89.245 128.505 89.910 128.675 ;
        RECT 90.195 128.630 90.365 129.430 ;
        RECT 90.995 129.745 91.510 130.155 ;
        RECT 91.745 129.745 91.915 130.505 ;
        RECT 92.085 130.165 94.115 130.335 ;
        RECT 90.995 128.935 91.335 129.745 ;
        RECT 92.085 129.500 92.255 130.165 ;
        RECT 92.650 129.825 93.775 129.995 ;
        RECT 91.505 129.310 92.255 129.500 ;
        RECT 92.425 129.485 93.435 129.655 ;
        RECT 90.995 128.765 92.225 128.935 ;
        RECT 89.245 128.125 89.415 128.505 ;
        RECT 89.595 127.955 89.925 128.335 ;
        RECT 90.105 128.125 90.365 128.630 ;
        RECT 91.270 128.160 91.515 128.765 ;
        RECT 91.735 127.955 92.245 128.490 ;
        RECT 92.425 128.125 92.615 129.485 ;
        RECT 92.785 128.805 93.060 129.285 ;
        RECT 92.785 128.635 93.065 128.805 ;
        RECT 93.265 128.685 93.435 129.485 ;
        RECT 93.605 128.695 93.775 129.825 ;
        RECT 93.945 129.195 94.115 130.165 ;
        RECT 94.285 129.365 94.455 130.505 ;
        RECT 94.625 129.365 94.960 130.335 ;
        RECT 93.945 128.865 94.140 129.195 ;
        RECT 94.365 128.865 94.620 129.195 ;
        RECT 94.365 128.695 94.535 128.865 ;
        RECT 94.790 128.695 94.960 129.365 ;
        RECT 92.785 128.125 93.060 128.635 ;
        RECT 93.605 128.525 94.535 128.695 ;
        RECT 93.605 128.490 93.780 128.525 ;
        RECT 93.250 128.125 93.780 128.490 ;
        RECT 94.205 127.955 94.535 128.355 ;
        RECT 94.705 128.125 94.960 128.695 ;
        RECT 95.135 129.430 95.405 130.335 ;
        RECT 95.575 129.745 95.905 130.505 ;
        RECT 96.085 129.575 96.255 130.335 ;
        RECT 95.135 128.630 95.305 129.430 ;
        RECT 95.590 129.405 96.255 129.575 ;
        RECT 96.515 129.415 98.185 130.505 ;
        RECT 98.445 129.575 98.615 130.335 ;
        RECT 98.795 129.745 99.125 130.505 ;
        RECT 95.590 129.260 95.760 129.405 ;
        RECT 95.475 128.930 95.760 129.260 ;
        RECT 95.590 128.675 95.760 128.930 ;
        RECT 95.995 128.855 96.325 129.225 ;
        RECT 96.515 128.895 97.265 129.415 ;
        RECT 98.445 129.405 99.110 129.575 ;
        RECT 99.295 129.430 99.565 130.335 ;
        RECT 98.940 129.260 99.110 129.405 ;
        RECT 97.435 128.725 98.185 129.245 ;
        RECT 98.375 128.855 98.705 129.225 ;
        RECT 98.940 128.930 99.225 129.260 ;
        RECT 95.135 128.125 95.395 128.630 ;
        RECT 95.590 128.505 96.255 128.675 ;
        RECT 95.575 127.955 95.905 128.335 ;
        RECT 96.085 128.125 96.255 128.505 ;
        RECT 96.515 127.955 98.185 128.725 ;
        RECT 98.940 128.675 99.110 128.930 ;
        RECT 98.445 128.505 99.110 128.675 ;
        RECT 99.395 128.630 99.565 129.430 ;
        RECT 99.735 129.745 100.250 130.155 ;
        RECT 100.485 129.745 100.655 130.505 ;
        RECT 100.825 130.165 102.855 130.335 ;
        RECT 99.735 128.935 100.075 129.745 ;
        RECT 100.825 129.500 100.995 130.165 ;
        RECT 101.390 129.825 102.515 129.995 ;
        RECT 100.245 129.310 100.995 129.500 ;
        RECT 101.165 129.485 102.175 129.655 ;
        RECT 99.735 128.765 100.965 128.935 ;
        RECT 98.445 128.125 98.615 128.505 ;
        RECT 98.795 127.955 99.125 128.335 ;
        RECT 99.305 128.125 99.565 128.630 ;
        RECT 100.010 128.160 100.255 128.765 ;
        RECT 100.475 127.955 100.985 128.490 ;
        RECT 101.165 128.125 101.355 129.485 ;
        RECT 101.525 129.145 101.800 129.285 ;
        RECT 101.525 128.975 101.805 129.145 ;
        RECT 101.525 128.125 101.800 128.975 ;
        RECT 102.005 128.685 102.175 129.485 ;
        RECT 102.345 128.695 102.515 129.825 ;
        RECT 102.685 129.195 102.855 130.165 ;
        RECT 103.025 129.365 103.195 130.505 ;
        RECT 103.365 129.365 103.700 130.335 ;
        RECT 103.915 129.365 104.145 130.505 ;
        RECT 102.685 128.865 102.880 129.195 ;
        RECT 103.105 128.865 103.360 129.195 ;
        RECT 103.105 128.695 103.275 128.865 ;
        RECT 103.530 128.695 103.700 129.365 ;
        RECT 104.315 129.355 104.645 130.335 ;
        RECT 104.815 129.365 105.025 130.505 ;
        RECT 105.295 129.365 105.525 130.505 ;
        RECT 105.695 129.355 106.025 130.335 ;
        RECT 106.195 129.365 106.405 130.505 ;
        RECT 106.725 129.575 106.895 130.335 ;
        RECT 107.075 129.745 107.405 130.505 ;
        RECT 106.725 129.405 107.390 129.575 ;
        RECT 107.575 129.430 107.845 130.335 ;
        RECT 103.895 128.945 104.225 129.195 ;
        RECT 102.345 128.525 103.275 128.695 ;
        RECT 102.345 128.490 102.520 128.525 ;
        RECT 101.990 128.125 102.520 128.490 ;
        RECT 102.945 127.955 103.275 128.355 ;
        RECT 103.445 128.125 103.700 128.695 ;
        RECT 103.915 127.955 104.145 128.775 ;
        RECT 104.395 128.755 104.645 129.355 ;
        RECT 105.275 128.945 105.605 129.195 ;
        RECT 104.315 128.125 104.645 128.755 ;
        RECT 104.815 127.955 105.025 128.775 ;
        RECT 105.295 127.955 105.525 128.775 ;
        RECT 105.775 128.755 106.025 129.355 ;
        RECT 107.220 129.260 107.390 129.405 ;
        RECT 106.655 128.855 106.985 129.225 ;
        RECT 107.220 128.930 107.505 129.260 ;
        RECT 105.695 128.125 106.025 128.755 ;
        RECT 106.195 127.955 106.405 128.775 ;
        RECT 107.220 128.675 107.390 128.930 ;
        RECT 106.725 128.505 107.390 128.675 ;
        RECT 107.675 128.630 107.845 129.430 ;
        RECT 108.475 129.415 111.985 130.505 ;
        RECT 112.155 129.415 113.365 130.505 ;
        RECT 108.475 128.895 110.165 129.415 ;
        RECT 110.335 128.725 111.985 129.245 ;
        RECT 112.155 128.875 112.675 129.415 ;
        RECT 106.725 128.125 106.895 128.505 ;
        RECT 107.075 127.955 107.405 128.335 ;
        RECT 107.585 128.125 107.845 128.630 ;
        RECT 108.475 127.955 111.985 128.725 ;
        RECT 112.845 128.705 113.365 129.245 ;
        RECT 112.155 127.955 113.365 128.705 ;
        RECT 22.830 127.785 113.450 127.955 ;
        RECT 22.915 127.035 24.125 127.785 ;
        RECT 22.915 126.495 23.435 127.035 ;
        RECT 24.355 126.965 24.565 127.785 ;
        RECT 24.735 126.985 25.065 127.615 ;
        RECT 23.605 126.325 24.125 126.865 ;
        RECT 24.735 126.385 24.985 126.985 ;
        RECT 25.235 126.965 25.465 127.785 ;
        RECT 25.715 126.965 25.945 127.785 ;
        RECT 26.115 126.985 26.445 127.615 ;
        RECT 25.155 126.545 25.485 126.795 ;
        RECT 25.695 126.545 26.025 126.795 ;
        RECT 26.195 126.385 26.445 126.985 ;
        RECT 26.615 126.965 26.825 127.785 ;
        RECT 27.145 127.235 27.315 127.615 ;
        RECT 27.495 127.405 27.825 127.785 ;
        RECT 27.145 127.065 27.810 127.235 ;
        RECT 28.005 127.110 28.265 127.615 ;
        RECT 27.075 126.515 27.405 126.885 ;
        RECT 27.640 126.810 27.810 127.065 ;
        RECT 22.915 125.235 24.125 126.325 ;
        RECT 24.355 125.235 24.565 126.375 ;
        RECT 24.735 125.405 25.065 126.385 ;
        RECT 25.235 125.235 25.465 126.375 ;
        RECT 25.715 125.235 25.945 126.375 ;
        RECT 26.115 125.405 26.445 126.385 ;
        RECT 27.640 126.480 27.925 126.810 ;
        RECT 26.615 125.235 26.825 126.375 ;
        RECT 27.640 126.335 27.810 126.480 ;
        RECT 27.145 126.165 27.810 126.335 ;
        RECT 28.095 126.310 28.265 127.110 ;
        RECT 27.145 125.405 27.315 126.165 ;
        RECT 27.495 125.235 27.825 125.995 ;
        RECT 27.995 125.405 28.265 126.310 ;
        RECT 28.440 127.045 28.695 127.615 ;
        RECT 28.865 127.385 29.195 127.785 ;
        RECT 29.620 127.250 30.150 127.615 ;
        RECT 29.620 127.215 29.795 127.250 ;
        RECT 28.865 127.045 29.795 127.215 ;
        RECT 28.440 126.375 28.610 127.045 ;
        RECT 28.865 126.875 29.035 127.045 ;
        RECT 28.780 126.545 29.035 126.875 ;
        RECT 29.260 126.545 29.455 126.875 ;
        RECT 28.440 125.405 28.775 126.375 ;
        RECT 28.945 125.235 29.115 126.375 ;
        RECT 29.285 125.575 29.455 126.545 ;
        RECT 29.625 125.915 29.795 127.045 ;
        RECT 29.965 126.255 30.135 127.055 ;
        RECT 30.340 126.765 30.615 127.615 ;
        RECT 30.335 126.595 30.615 126.765 ;
        RECT 30.340 126.455 30.615 126.595 ;
        RECT 30.785 126.255 30.975 127.615 ;
        RECT 31.155 127.250 31.665 127.785 ;
        RECT 31.885 126.975 32.130 127.580 ;
        RECT 32.950 127.445 33.205 127.605 ;
        RECT 32.865 127.275 33.205 127.445 ;
        RECT 33.385 127.325 33.670 127.785 ;
        RECT 32.950 127.075 33.205 127.275 ;
        RECT 31.175 126.805 32.405 126.975 ;
        RECT 29.965 126.085 30.975 126.255 ;
        RECT 31.145 126.240 31.895 126.430 ;
        RECT 29.625 125.745 30.750 125.915 ;
        RECT 31.145 125.575 31.315 126.240 ;
        RECT 32.065 125.995 32.405 126.805 ;
        RECT 29.285 125.405 31.315 125.575 ;
        RECT 31.485 125.235 31.655 125.995 ;
        RECT 31.890 125.585 32.405 125.995 ;
        RECT 32.950 126.215 33.130 127.075 ;
        RECT 33.850 126.875 34.100 127.525 ;
        RECT 33.300 126.545 34.100 126.875 ;
        RECT 32.950 125.545 33.205 126.215 ;
        RECT 33.385 125.235 33.670 126.035 ;
        RECT 33.850 125.955 34.100 126.545 ;
        RECT 34.300 127.190 34.620 127.520 ;
        RECT 34.800 127.305 35.460 127.785 ;
        RECT 35.660 127.395 36.510 127.565 ;
        RECT 34.300 126.295 34.490 127.190 ;
        RECT 34.810 126.865 35.470 127.135 ;
        RECT 35.140 126.805 35.470 126.865 ;
        RECT 34.660 126.635 34.990 126.695 ;
        RECT 35.660 126.635 35.830 127.395 ;
        RECT 37.070 127.325 37.390 127.785 ;
        RECT 37.590 127.145 37.840 127.575 ;
        RECT 38.130 127.345 38.540 127.785 ;
        RECT 38.710 127.405 39.725 127.605 ;
        RECT 36.000 126.975 37.250 127.145 ;
        RECT 36.000 126.855 36.330 126.975 ;
        RECT 34.660 126.465 36.560 126.635 ;
        RECT 34.300 126.125 36.220 126.295 ;
        RECT 34.300 126.105 34.620 126.125 ;
        RECT 33.850 125.445 34.180 125.955 ;
        RECT 34.450 125.495 34.620 126.105 ;
        RECT 36.390 125.955 36.560 126.465 ;
        RECT 36.730 126.395 36.910 126.805 ;
        RECT 37.080 126.215 37.250 126.975 ;
        RECT 34.790 125.235 35.120 125.925 ;
        RECT 35.350 125.785 36.560 125.955 ;
        RECT 36.730 125.905 37.250 126.215 ;
        RECT 37.420 126.805 37.840 127.145 ;
        RECT 38.130 126.805 38.540 127.135 ;
        RECT 37.420 126.035 37.610 126.805 ;
        RECT 38.710 126.675 38.880 127.405 ;
        RECT 40.025 127.235 40.195 127.565 ;
        RECT 40.365 127.405 40.695 127.785 ;
        RECT 39.050 126.855 39.400 127.225 ;
        RECT 38.710 126.635 39.130 126.675 ;
        RECT 37.780 126.465 39.130 126.635 ;
        RECT 37.780 126.305 38.030 126.465 ;
        RECT 38.540 126.035 38.790 126.295 ;
        RECT 37.420 125.785 38.790 126.035 ;
        RECT 35.350 125.495 35.590 125.785 ;
        RECT 36.390 125.705 36.560 125.785 ;
        RECT 35.790 125.235 36.210 125.615 ;
        RECT 36.390 125.455 37.020 125.705 ;
        RECT 37.490 125.235 37.820 125.615 ;
        RECT 37.990 125.495 38.160 125.785 ;
        RECT 38.960 125.620 39.130 126.465 ;
        RECT 39.580 126.295 39.800 127.165 ;
        RECT 40.025 127.045 40.720 127.235 ;
        RECT 39.300 125.915 39.800 126.295 ;
        RECT 39.970 126.245 40.380 126.865 ;
        RECT 40.550 126.075 40.720 127.045 ;
        RECT 40.025 125.905 40.720 126.075 ;
        RECT 38.340 125.235 38.720 125.615 ;
        RECT 38.960 125.450 39.790 125.620 ;
        RECT 40.025 125.405 40.195 125.905 ;
        RECT 40.365 125.235 40.695 125.735 ;
        RECT 40.910 125.405 41.135 127.525 ;
        RECT 41.305 127.405 41.635 127.785 ;
        RECT 41.805 127.235 41.975 127.525 ;
        RECT 41.310 127.065 41.975 127.235 ;
        RECT 42.435 127.155 42.765 127.515 ;
        RECT 43.385 127.325 43.635 127.785 ;
        RECT 43.805 127.325 44.365 127.615 ;
        RECT 41.310 126.075 41.540 127.065 ;
        RECT 42.435 126.965 43.825 127.155 ;
        RECT 41.710 126.245 42.060 126.895 ;
        RECT 43.655 126.875 43.825 126.965 ;
        RECT 42.250 126.545 42.925 126.795 ;
        RECT 43.145 126.545 43.485 126.795 ;
        RECT 43.655 126.545 43.945 126.875 ;
        RECT 42.250 126.185 42.515 126.545 ;
        RECT 43.655 126.295 43.825 126.545 ;
        RECT 42.885 126.125 43.825 126.295 ;
        RECT 41.310 125.905 41.975 126.075 ;
        RECT 41.305 125.235 41.635 125.735 ;
        RECT 41.805 125.405 41.975 125.905 ;
        RECT 42.435 125.235 42.715 125.905 ;
        RECT 42.885 125.575 43.185 126.125 ;
        RECT 44.115 125.955 44.365 127.325 ;
        RECT 44.685 126.985 45.015 127.785 ;
        RECT 45.185 127.135 45.355 127.615 ;
        RECT 45.525 127.305 45.855 127.785 ;
        RECT 46.025 127.135 46.195 127.615 ;
        RECT 46.445 127.305 46.685 127.785 ;
        RECT 46.865 127.135 47.035 127.615 ;
        RECT 45.185 126.965 46.195 127.135 ;
        RECT 46.400 126.965 47.035 127.135 ;
        RECT 47.335 126.965 47.565 127.785 ;
        RECT 47.735 126.985 48.065 127.615 ;
        RECT 45.185 126.935 45.685 126.965 ;
        RECT 45.185 126.425 45.680 126.935 ;
        RECT 46.400 126.795 46.570 126.965 ;
        RECT 46.070 126.625 46.570 126.795 ;
        RECT 43.385 125.235 43.715 125.955 ;
        RECT 43.905 125.405 44.365 125.955 ;
        RECT 44.685 125.235 45.015 126.385 ;
        RECT 45.185 126.255 46.195 126.425 ;
        RECT 45.185 125.405 45.355 126.255 ;
        RECT 45.525 125.235 45.855 126.035 ;
        RECT 46.025 125.405 46.195 126.255 ;
        RECT 46.400 126.385 46.570 126.625 ;
        RECT 46.740 126.555 47.120 126.795 ;
        RECT 47.315 126.545 47.645 126.795 ;
        RECT 47.815 126.385 48.065 126.985 ;
        RECT 48.235 126.965 48.445 127.785 ;
        RECT 48.675 127.060 48.965 127.785 ;
        RECT 49.510 127.445 49.765 127.605 ;
        RECT 49.425 127.275 49.765 127.445 ;
        RECT 49.945 127.325 50.230 127.785 ;
        RECT 49.510 127.075 49.765 127.275 ;
        RECT 46.400 126.215 47.115 126.385 ;
        RECT 46.375 125.235 46.615 126.035 ;
        RECT 46.785 125.405 47.115 126.215 ;
        RECT 47.335 125.235 47.565 126.375 ;
        RECT 47.735 125.405 48.065 126.385 ;
        RECT 48.235 125.235 48.445 126.375 ;
        RECT 48.675 125.235 48.965 126.400 ;
        RECT 49.510 126.215 49.690 127.075 ;
        RECT 50.410 126.875 50.660 127.525 ;
        RECT 49.860 126.545 50.660 126.875 ;
        RECT 49.510 125.545 49.765 126.215 ;
        RECT 49.945 125.235 50.230 126.035 ;
        RECT 50.410 125.955 50.660 126.545 ;
        RECT 50.860 127.190 51.180 127.520 ;
        RECT 51.360 127.305 52.020 127.785 ;
        RECT 52.220 127.395 53.070 127.565 ;
        RECT 50.860 126.295 51.050 127.190 ;
        RECT 51.370 126.865 52.030 127.135 ;
        RECT 51.700 126.805 52.030 126.865 ;
        RECT 51.220 126.635 51.550 126.695 ;
        RECT 52.220 126.635 52.390 127.395 ;
        RECT 53.630 127.325 53.950 127.785 ;
        RECT 54.150 127.145 54.400 127.575 ;
        RECT 54.690 127.345 55.100 127.785 ;
        RECT 55.270 127.405 56.285 127.605 ;
        RECT 52.560 126.975 53.810 127.145 ;
        RECT 52.560 126.855 52.890 126.975 ;
        RECT 51.220 126.465 53.120 126.635 ;
        RECT 50.860 126.125 52.780 126.295 ;
        RECT 50.860 126.105 51.180 126.125 ;
        RECT 50.410 125.445 50.740 125.955 ;
        RECT 51.010 125.495 51.180 126.105 ;
        RECT 52.950 125.955 53.120 126.465 ;
        RECT 53.290 126.395 53.470 126.805 ;
        RECT 53.640 126.215 53.810 126.975 ;
        RECT 51.350 125.235 51.680 125.925 ;
        RECT 51.910 125.785 53.120 125.955 ;
        RECT 53.290 125.905 53.810 126.215 ;
        RECT 53.980 126.805 54.400 127.145 ;
        RECT 54.690 126.805 55.100 127.135 ;
        RECT 53.980 126.035 54.170 126.805 ;
        RECT 55.270 126.675 55.440 127.405 ;
        RECT 56.585 127.235 56.755 127.565 ;
        RECT 56.925 127.405 57.255 127.785 ;
        RECT 55.610 126.855 55.960 127.225 ;
        RECT 55.270 126.635 55.690 126.675 ;
        RECT 54.340 126.465 55.690 126.635 ;
        RECT 54.340 126.305 54.590 126.465 ;
        RECT 55.100 126.035 55.350 126.295 ;
        RECT 53.980 125.785 55.350 126.035 ;
        RECT 51.910 125.495 52.150 125.785 ;
        RECT 52.950 125.705 53.120 125.785 ;
        RECT 52.350 125.235 52.770 125.615 ;
        RECT 52.950 125.455 53.580 125.705 ;
        RECT 54.050 125.235 54.380 125.615 ;
        RECT 54.550 125.495 54.720 125.785 ;
        RECT 55.520 125.620 55.690 126.465 ;
        RECT 56.140 126.295 56.360 127.165 ;
        RECT 56.585 127.045 57.280 127.235 ;
        RECT 55.860 125.915 56.360 126.295 ;
        RECT 56.530 126.245 56.940 126.865 ;
        RECT 57.110 126.075 57.280 127.045 ;
        RECT 56.585 125.905 57.280 126.075 ;
        RECT 54.900 125.235 55.280 125.615 ;
        RECT 55.520 125.450 56.350 125.620 ;
        RECT 56.585 125.405 56.755 125.905 ;
        RECT 56.925 125.235 57.255 125.735 ;
        RECT 57.470 125.405 57.695 127.525 ;
        RECT 57.865 127.405 58.195 127.785 ;
        RECT 58.365 127.235 58.535 127.525 ;
        RECT 57.870 127.065 58.535 127.235 ;
        RECT 57.870 126.075 58.100 127.065 ;
        RECT 58.855 126.965 59.065 127.785 ;
        RECT 59.235 126.985 59.565 127.615 ;
        RECT 58.270 126.245 58.620 126.895 ;
        RECT 59.235 126.385 59.485 126.985 ;
        RECT 59.735 126.965 59.965 127.785 ;
        RECT 60.635 127.110 60.895 127.615 ;
        RECT 61.075 127.405 61.405 127.785 ;
        RECT 61.585 127.235 61.755 127.615 ;
        RECT 59.655 126.545 59.985 126.795 ;
        RECT 57.870 125.905 58.535 126.075 ;
        RECT 57.865 125.235 58.195 125.735 ;
        RECT 58.365 125.405 58.535 125.905 ;
        RECT 58.855 125.235 59.065 126.375 ;
        RECT 59.235 125.405 59.565 126.385 ;
        RECT 59.735 125.235 59.965 126.375 ;
        RECT 60.635 126.310 60.805 127.110 ;
        RECT 61.090 127.065 61.755 127.235 ;
        RECT 61.090 126.810 61.260 127.065 ;
        RECT 62.015 127.015 63.685 127.785 ;
        RECT 60.975 126.480 61.260 126.810 ;
        RECT 61.495 126.515 61.825 126.885 ;
        RECT 61.090 126.335 61.260 126.480 ;
        RECT 60.635 125.405 60.905 126.310 ;
        RECT 61.090 126.165 61.755 126.335 ;
        RECT 61.075 125.235 61.405 125.995 ;
        RECT 61.585 125.405 61.755 126.165 ;
        RECT 62.015 126.325 62.765 126.845 ;
        RECT 62.935 126.495 63.685 127.015 ;
        RECT 63.895 126.965 64.125 127.785 ;
        RECT 64.295 126.985 64.625 127.615 ;
        RECT 63.875 126.545 64.205 126.795 ;
        RECT 64.375 126.385 64.625 126.985 ;
        RECT 64.795 126.965 65.005 127.785 ;
        RECT 66.245 127.235 66.415 127.615 ;
        RECT 66.595 127.405 66.925 127.785 ;
        RECT 66.245 127.065 66.910 127.235 ;
        RECT 67.105 127.110 67.365 127.615 ;
        RECT 66.175 126.515 66.505 126.885 ;
        RECT 66.740 126.810 66.910 127.065 ;
        RECT 62.015 125.235 63.685 126.325 ;
        RECT 63.895 125.235 64.125 126.375 ;
        RECT 64.295 125.405 64.625 126.385 ;
        RECT 66.740 126.480 67.025 126.810 ;
        RECT 64.795 125.235 65.005 126.375 ;
        RECT 66.740 126.335 66.910 126.480 ;
        RECT 66.245 126.165 66.910 126.335 ;
        RECT 67.195 126.310 67.365 127.110 ;
        RECT 67.535 127.015 70.125 127.785 ;
        RECT 66.245 125.405 66.415 126.165 ;
        RECT 66.595 125.235 66.925 125.995 ;
        RECT 67.095 125.405 67.365 126.310 ;
        RECT 67.535 126.325 68.745 126.845 ;
        RECT 68.915 126.495 70.125 127.015 ;
        RECT 70.335 126.965 70.565 127.785 ;
        RECT 70.735 126.985 71.065 127.615 ;
        RECT 70.315 126.545 70.645 126.795 ;
        RECT 70.815 126.385 71.065 126.985 ;
        RECT 71.235 126.965 71.445 127.785 ;
        RECT 71.715 126.965 71.945 127.785 ;
        RECT 72.115 126.985 72.445 127.615 ;
        RECT 71.695 126.545 72.025 126.795 ;
        RECT 72.195 126.385 72.445 126.985 ;
        RECT 72.615 126.965 72.825 127.785 ;
        RECT 73.055 127.035 74.265 127.785 ;
        RECT 74.435 127.060 74.725 127.785 ;
        RECT 75.270 127.445 75.525 127.605 ;
        RECT 75.185 127.275 75.525 127.445 ;
        RECT 75.705 127.325 75.990 127.785 ;
        RECT 75.270 127.075 75.525 127.275 ;
        RECT 67.535 125.235 70.125 126.325 ;
        RECT 70.335 125.235 70.565 126.375 ;
        RECT 70.735 125.405 71.065 126.385 ;
        RECT 71.235 125.235 71.445 126.375 ;
        RECT 71.715 125.235 71.945 126.375 ;
        RECT 72.115 125.405 72.445 126.385 ;
        RECT 72.615 125.235 72.825 126.375 ;
        RECT 73.055 126.325 73.575 126.865 ;
        RECT 73.745 126.495 74.265 127.035 ;
        RECT 73.055 125.235 74.265 126.325 ;
        RECT 74.435 125.235 74.725 126.400 ;
        RECT 75.270 126.215 75.450 127.075 ;
        RECT 76.170 126.875 76.420 127.525 ;
        RECT 75.620 126.545 76.420 126.875 ;
        RECT 75.270 125.545 75.525 126.215 ;
        RECT 75.705 125.235 75.990 126.035 ;
        RECT 76.170 125.955 76.420 126.545 ;
        RECT 76.620 127.190 76.940 127.520 ;
        RECT 77.120 127.305 77.780 127.785 ;
        RECT 77.980 127.395 78.830 127.565 ;
        RECT 76.620 126.295 76.810 127.190 ;
        RECT 77.130 126.865 77.790 127.135 ;
        RECT 77.460 126.805 77.790 126.865 ;
        RECT 76.980 126.635 77.310 126.695 ;
        RECT 77.980 126.635 78.150 127.395 ;
        RECT 79.390 127.325 79.710 127.785 ;
        RECT 79.910 127.145 80.160 127.575 ;
        RECT 80.450 127.345 80.860 127.785 ;
        RECT 81.030 127.405 82.045 127.605 ;
        RECT 78.320 126.975 79.570 127.145 ;
        RECT 78.320 126.855 78.650 126.975 ;
        RECT 76.980 126.465 78.880 126.635 ;
        RECT 76.620 126.125 78.540 126.295 ;
        RECT 76.620 126.105 76.940 126.125 ;
        RECT 76.170 125.445 76.500 125.955 ;
        RECT 76.770 125.495 76.940 126.105 ;
        RECT 78.710 125.955 78.880 126.465 ;
        RECT 79.050 126.395 79.230 126.805 ;
        RECT 79.400 126.215 79.570 126.975 ;
        RECT 77.110 125.235 77.440 125.925 ;
        RECT 77.670 125.785 78.880 125.955 ;
        RECT 79.050 125.905 79.570 126.215 ;
        RECT 79.740 126.805 80.160 127.145 ;
        RECT 80.450 126.805 80.860 127.135 ;
        RECT 79.740 126.035 79.930 126.805 ;
        RECT 81.030 126.675 81.200 127.405 ;
        RECT 82.345 127.235 82.515 127.565 ;
        RECT 82.685 127.405 83.015 127.785 ;
        RECT 81.370 126.855 81.720 127.225 ;
        RECT 81.030 126.635 81.450 126.675 ;
        RECT 80.100 126.465 81.450 126.635 ;
        RECT 80.100 126.305 80.350 126.465 ;
        RECT 80.860 126.035 81.110 126.295 ;
        RECT 79.740 125.785 81.110 126.035 ;
        RECT 77.670 125.495 77.910 125.785 ;
        RECT 78.710 125.705 78.880 125.785 ;
        RECT 78.110 125.235 78.530 125.615 ;
        RECT 78.710 125.455 79.340 125.705 ;
        RECT 79.810 125.235 80.140 125.615 ;
        RECT 80.310 125.495 80.480 125.785 ;
        RECT 81.280 125.620 81.450 126.465 ;
        RECT 81.900 126.295 82.120 127.165 ;
        RECT 82.345 127.045 83.040 127.235 ;
        RECT 81.620 125.915 82.120 126.295 ;
        RECT 82.290 126.245 82.700 126.865 ;
        RECT 82.870 126.075 83.040 127.045 ;
        RECT 82.345 125.905 83.040 126.075 ;
        RECT 80.660 125.235 81.040 125.615 ;
        RECT 81.280 125.450 82.110 125.620 ;
        RECT 82.345 125.405 82.515 125.905 ;
        RECT 82.685 125.235 83.015 125.735 ;
        RECT 83.230 125.405 83.455 127.525 ;
        RECT 83.625 127.405 83.955 127.785 ;
        RECT 84.125 127.235 84.295 127.525 ;
        RECT 84.930 127.445 85.185 127.605 ;
        RECT 84.845 127.275 85.185 127.445 ;
        RECT 85.365 127.325 85.650 127.785 ;
        RECT 83.630 127.065 84.295 127.235 ;
        RECT 84.930 127.075 85.185 127.275 ;
        RECT 83.630 126.075 83.860 127.065 ;
        RECT 84.030 126.245 84.380 126.895 ;
        RECT 84.930 126.215 85.110 127.075 ;
        RECT 85.830 126.875 86.080 127.525 ;
        RECT 85.280 126.545 86.080 126.875 ;
        RECT 83.630 125.905 84.295 126.075 ;
        RECT 83.625 125.235 83.955 125.735 ;
        RECT 84.125 125.405 84.295 125.905 ;
        RECT 84.930 125.545 85.185 126.215 ;
        RECT 85.365 125.235 85.650 126.035 ;
        RECT 85.830 125.955 86.080 126.545 ;
        RECT 86.280 127.190 86.600 127.520 ;
        RECT 86.780 127.305 87.440 127.785 ;
        RECT 87.640 127.395 88.490 127.565 ;
        RECT 86.280 126.295 86.470 127.190 ;
        RECT 86.790 126.865 87.450 127.135 ;
        RECT 87.120 126.805 87.450 126.865 ;
        RECT 86.640 126.635 86.970 126.695 ;
        RECT 87.640 126.635 87.810 127.395 ;
        RECT 89.050 127.325 89.370 127.785 ;
        RECT 89.570 127.145 89.820 127.575 ;
        RECT 90.110 127.345 90.520 127.785 ;
        RECT 90.690 127.405 91.705 127.605 ;
        RECT 87.980 126.975 89.230 127.145 ;
        RECT 87.980 126.855 88.310 126.975 ;
        RECT 86.640 126.465 88.540 126.635 ;
        RECT 86.280 126.125 88.200 126.295 ;
        RECT 86.280 126.105 86.600 126.125 ;
        RECT 85.830 125.445 86.160 125.955 ;
        RECT 86.430 125.495 86.600 126.105 ;
        RECT 88.370 125.955 88.540 126.465 ;
        RECT 88.710 126.395 88.890 126.805 ;
        RECT 89.060 126.215 89.230 126.975 ;
        RECT 86.770 125.235 87.100 125.925 ;
        RECT 87.330 125.785 88.540 125.955 ;
        RECT 88.710 125.905 89.230 126.215 ;
        RECT 89.400 126.805 89.820 127.145 ;
        RECT 90.110 126.805 90.520 127.135 ;
        RECT 89.400 126.035 89.590 126.805 ;
        RECT 90.690 126.675 90.860 127.405 ;
        RECT 92.005 127.235 92.175 127.565 ;
        RECT 92.345 127.405 92.675 127.785 ;
        RECT 91.030 126.855 91.380 127.225 ;
        RECT 90.690 126.635 91.110 126.675 ;
        RECT 89.760 126.465 91.110 126.635 ;
        RECT 89.760 126.305 90.010 126.465 ;
        RECT 90.520 126.035 90.770 126.295 ;
        RECT 89.400 125.785 90.770 126.035 ;
        RECT 87.330 125.495 87.570 125.785 ;
        RECT 88.370 125.705 88.540 125.785 ;
        RECT 87.770 125.235 88.190 125.615 ;
        RECT 88.370 125.455 89.000 125.705 ;
        RECT 89.470 125.235 89.800 125.615 ;
        RECT 89.970 125.495 90.140 125.785 ;
        RECT 90.940 125.620 91.110 126.465 ;
        RECT 91.560 126.295 91.780 127.165 ;
        RECT 92.005 127.045 92.700 127.235 ;
        RECT 91.280 125.915 91.780 126.295 ;
        RECT 91.950 126.245 92.360 126.865 ;
        RECT 92.530 126.075 92.700 127.045 ;
        RECT 92.005 125.905 92.700 126.075 ;
        RECT 90.320 125.235 90.700 125.615 ;
        RECT 90.940 125.450 91.770 125.620 ;
        RECT 92.005 125.405 92.175 125.905 ;
        RECT 92.345 125.235 92.675 125.735 ;
        RECT 92.890 125.405 93.115 127.525 ;
        RECT 93.285 127.405 93.615 127.785 ;
        RECT 93.785 127.235 93.955 127.525 ;
        RECT 94.680 127.240 100.025 127.785 ;
        RECT 93.290 127.065 93.955 127.235 ;
        RECT 93.290 126.075 93.520 127.065 ;
        RECT 93.690 126.245 94.040 126.895 ;
        RECT 93.290 125.905 93.955 126.075 ;
        RECT 93.285 125.235 93.615 125.735 ;
        RECT 93.785 125.405 93.955 125.905 ;
        RECT 96.270 125.670 96.620 126.920 ;
        RECT 98.100 126.410 98.440 127.240 ;
        RECT 100.195 127.060 100.485 127.785 ;
        RECT 100.660 127.240 106.005 127.785 ;
        RECT 94.680 125.235 100.025 125.670 ;
        RECT 100.195 125.235 100.485 126.400 ;
        RECT 102.250 125.670 102.600 126.920 ;
        RECT 104.080 126.410 104.420 127.240 ;
        RECT 106.215 126.965 106.445 127.785 ;
        RECT 106.615 126.985 106.945 127.615 ;
        RECT 106.195 126.545 106.525 126.795 ;
        RECT 106.695 126.385 106.945 126.985 ;
        RECT 107.115 126.965 107.325 127.785 ;
        RECT 107.555 127.035 108.765 127.785 ;
        RECT 100.660 125.235 106.005 125.670 ;
        RECT 106.215 125.235 106.445 126.375 ;
        RECT 106.615 125.405 106.945 126.385 ;
        RECT 107.115 125.235 107.325 126.375 ;
        RECT 107.555 126.325 108.075 126.865 ;
        RECT 108.245 126.495 108.765 127.035 ;
        RECT 108.935 127.110 109.195 127.615 ;
        RECT 109.375 127.405 109.705 127.785 ;
        RECT 109.885 127.235 110.055 127.615 ;
        RECT 107.555 125.235 108.765 126.325 ;
        RECT 108.935 126.310 109.105 127.110 ;
        RECT 109.390 127.065 110.055 127.235 ;
        RECT 110.775 127.110 111.035 127.615 ;
        RECT 111.215 127.405 111.545 127.785 ;
        RECT 111.725 127.235 111.895 127.615 ;
        RECT 109.390 126.810 109.560 127.065 ;
        RECT 109.275 126.480 109.560 126.810 ;
        RECT 109.795 126.515 110.125 126.885 ;
        RECT 109.390 126.335 109.560 126.480 ;
        RECT 108.935 125.405 109.205 126.310 ;
        RECT 109.390 126.165 110.055 126.335 ;
        RECT 109.375 125.235 109.705 125.995 ;
        RECT 109.885 125.405 110.055 126.165 ;
        RECT 110.775 126.310 110.955 127.110 ;
        RECT 111.230 127.065 111.895 127.235 ;
        RECT 111.230 126.810 111.400 127.065 ;
        RECT 112.155 127.035 113.365 127.785 ;
        RECT 111.125 126.480 111.400 126.810 ;
        RECT 111.625 126.515 111.965 126.885 ;
        RECT 111.230 126.335 111.400 126.480 ;
        RECT 110.775 125.405 111.045 126.310 ;
        RECT 111.230 126.165 111.905 126.335 ;
        RECT 111.215 125.235 111.545 125.995 ;
        RECT 111.725 125.405 111.905 126.165 ;
        RECT 112.155 126.325 112.675 126.865 ;
        RECT 112.845 126.495 113.365 127.035 ;
        RECT 112.155 125.235 113.365 126.325 ;
        RECT 22.830 125.065 113.450 125.235 ;
        RECT 22.915 123.975 24.125 125.065 ;
        RECT 24.605 124.225 24.775 125.065 ;
        RECT 24.985 124.055 25.235 124.895 ;
        RECT 25.445 124.225 25.615 125.065 ;
        RECT 25.785 124.055 26.075 124.895 ;
        RECT 22.915 123.265 23.435 123.805 ;
        RECT 23.605 123.435 24.125 123.975 ;
        RECT 24.350 123.885 26.075 124.055 ;
        RECT 26.285 124.005 26.455 125.065 ;
        RECT 26.750 124.685 27.080 125.065 ;
        RECT 27.260 124.515 27.430 124.805 ;
        RECT 27.600 124.605 27.850 125.065 ;
        RECT 26.630 124.345 27.430 124.515 ;
        RECT 28.020 124.555 28.890 124.895 ;
        RECT 24.350 123.335 24.760 123.885 ;
        RECT 26.630 123.725 26.800 124.345 ;
        RECT 28.020 124.175 28.190 124.555 ;
        RECT 29.125 124.435 29.295 124.895 ;
        RECT 29.465 124.605 29.835 125.065 ;
        RECT 30.130 124.465 30.300 124.805 ;
        RECT 30.470 124.635 30.800 125.065 ;
        RECT 31.035 124.465 31.205 124.805 ;
        RECT 26.970 124.005 28.190 124.175 ;
        RECT 28.360 124.095 28.820 124.385 ;
        RECT 29.125 124.265 29.685 124.435 ;
        RECT 30.130 124.295 31.205 124.465 ;
        RECT 31.375 124.565 32.055 124.895 ;
        RECT 32.270 124.565 32.520 124.895 ;
        RECT 32.690 124.605 32.940 125.065 ;
        RECT 29.515 124.125 29.685 124.265 ;
        RECT 28.360 124.085 29.325 124.095 ;
        RECT 28.020 123.915 28.190 124.005 ;
        RECT 28.650 123.925 29.325 124.085 ;
        RECT 26.630 123.715 26.975 123.725 ;
        RECT 24.945 123.505 26.975 123.715 ;
        RECT 22.915 122.515 24.125 123.265 ;
        RECT 24.350 123.165 26.115 123.335 ;
        RECT 24.605 122.515 24.775 122.985 ;
        RECT 24.945 122.685 25.275 123.165 ;
        RECT 25.445 122.515 25.615 122.985 ;
        RECT 25.785 122.685 26.115 123.165 ;
        RECT 26.285 122.515 26.455 123.325 ;
        RECT 26.650 123.250 26.975 123.505 ;
        RECT 26.655 122.895 26.975 123.250 ;
        RECT 27.145 123.465 27.685 123.835 ;
        RECT 28.020 123.745 28.425 123.915 ;
        RECT 27.145 123.065 27.385 123.465 ;
        RECT 27.865 123.295 28.085 123.575 ;
        RECT 27.555 123.125 28.085 123.295 ;
        RECT 27.555 122.895 27.725 123.125 ;
        RECT 28.255 122.965 28.425 123.745 ;
        RECT 28.595 123.135 28.945 123.755 ;
        RECT 29.115 123.135 29.325 123.925 ;
        RECT 29.515 123.955 31.015 124.125 ;
        RECT 29.515 123.265 29.685 123.955 ;
        RECT 31.375 123.785 31.545 124.565 ;
        RECT 32.350 124.435 32.520 124.565 ;
        RECT 29.855 123.615 31.545 123.785 ;
        RECT 31.715 124.005 32.180 124.395 ;
        RECT 32.350 124.265 32.745 124.435 ;
        RECT 29.855 123.435 30.025 123.615 ;
        RECT 26.655 122.725 27.725 122.895 ;
        RECT 27.895 122.515 28.085 122.955 ;
        RECT 28.255 122.685 29.205 122.965 ;
        RECT 29.515 122.875 29.775 123.265 ;
        RECT 30.195 123.195 30.985 123.445 ;
        RECT 29.425 122.705 29.775 122.875 ;
        RECT 29.985 122.515 30.315 122.975 ;
        RECT 31.190 122.905 31.360 123.615 ;
        RECT 31.715 123.415 31.885 124.005 ;
        RECT 31.530 123.195 31.885 123.415 ;
        RECT 32.055 123.195 32.405 123.815 ;
        RECT 32.575 122.905 32.745 124.265 ;
        RECT 33.110 124.095 33.435 124.880 ;
        RECT 32.915 123.045 33.375 124.095 ;
        RECT 31.190 122.735 32.045 122.905 ;
        RECT 32.250 122.735 32.745 122.905 ;
        RECT 32.915 122.515 33.245 122.875 ;
        RECT 33.605 122.775 33.775 124.895 ;
        RECT 33.945 124.565 34.275 125.065 ;
        RECT 34.445 124.395 34.700 124.895 ;
        RECT 33.950 124.225 34.700 124.395 ;
        RECT 33.950 123.235 34.180 124.225 ;
        RECT 34.350 123.405 34.700 124.055 ;
        RECT 35.795 123.900 36.085 125.065 ;
        RECT 37.265 124.135 37.435 124.895 ;
        RECT 37.615 124.305 37.945 125.065 ;
        RECT 37.265 123.965 37.930 124.135 ;
        RECT 38.115 123.990 38.385 124.895 ;
        RECT 37.760 123.820 37.930 123.965 ;
        RECT 37.195 123.415 37.525 123.785 ;
        RECT 37.760 123.490 38.045 123.820 ;
        RECT 33.950 123.065 34.700 123.235 ;
        RECT 33.945 122.515 34.275 122.895 ;
        RECT 34.445 122.775 34.700 123.065 ;
        RECT 35.795 122.515 36.085 123.240 ;
        RECT 37.760 123.235 37.930 123.490 ;
        RECT 37.265 123.065 37.930 123.235 ;
        RECT 38.215 123.190 38.385 123.990 ;
        RECT 38.645 124.135 38.815 124.895 ;
        RECT 38.995 124.305 39.325 125.065 ;
        RECT 38.645 123.965 39.310 124.135 ;
        RECT 39.495 123.990 39.765 124.895 ;
        RECT 40.595 124.395 40.875 125.065 ;
        RECT 41.045 124.175 41.345 124.725 ;
        RECT 41.545 124.345 41.875 125.065 ;
        RECT 42.065 124.345 42.525 124.895 ;
        RECT 39.140 123.820 39.310 123.965 ;
        RECT 38.575 123.415 38.905 123.785 ;
        RECT 39.140 123.490 39.425 123.820 ;
        RECT 39.140 123.235 39.310 123.490 ;
        RECT 37.265 122.685 37.435 123.065 ;
        RECT 37.615 122.515 37.945 122.895 ;
        RECT 38.125 122.685 38.385 123.190 ;
        RECT 38.645 123.065 39.310 123.235 ;
        RECT 39.595 123.190 39.765 123.990 ;
        RECT 40.410 123.755 40.675 124.115 ;
        RECT 41.045 124.005 41.985 124.175 ;
        RECT 41.815 123.755 41.985 124.005 ;
        RECT 40.410 123.505 41.085 123.755 ;
        RECT 41.305 123.505 41.645 123.755 ;
        RECT 41.815 123.425 42.105 123.755 ;
        RECT 41.815 123.335 41.985 123.425 ;
        RECT 38.645 122.685 38.815 123.065 ;
        RECT 38.995 122.515 39.325 122.895 ;
        RECT 39.505 122.685 39.765 123.190 ;
        RECT 40.595 123.145 41.985 123.335 ;
        RECT 40.595 122.785 40.925 123.145 ;
        RECT 42.275 122.975 42.525 124.345 ;
        RECT 43.005 124.225 43.175 125.065 ;
        RECT 43.385 124.055 43.635 124.895 ;
        RECT 43.845 124.225 44.015 125.065 ;
        RECT 44.185 124.055 44.475 124.895 ;
        RECT 42.750 123.885 44.475 124.055 ;
        RECT 44.685 124.005 44.855 125.065 ;
        RECT 45.150 124.685 45.480 125.065 ;
        RECT 45.660 124.515 45.830 124.805 ;
        RECT 46.000 124.605 46.250 125.065 ;
        RECT 45.030 124.345 45.830 124.515 ;
        RECT 46.420 124.555 47.290 124.895 ;
        RECT 42.750 123.335 43.160 123.885 ;
        RECT 45.030 123.725 45.200 124.345 ;
        RECT 46.420 124.175 46.590 124.555 ;
        RECT 47.525 124.435 47.695 124.895 ;
        RECT 47.865 124.605 48.235 125.065 ;
        RECT 48.530 124.465 48.700 124.805 ;
        RECT 48.870 124.635 49.200 125.065 ;
        RECT 49.435 124.465 49.605 124.805 ;
        RECT 45.370 124.005 46.590 124.175 ;
        RECT 46.760 124.095 47.220 124.385 ;
        RECT 47.525 124.265 48.085 124.435 ;
        RECT 48.530 124.295 49.605 124.465 ;
        RECT 49.775 124.565 50.455 124.895 ;
        RECT 50.670 124.565 50.920 124.895 ;
        RECT 51.090 124.605 51.340 125.065 ;
        RECT 47.915 124.125 48.085 124.265 ;
        RECT 46.760 124.085 47.725 124.095 ;
        RECT 46.420 123.915 46.590 124.005 ;
        RECT 47.050 123.925 47.725 124.085 ;
        RECT 45.030 123.715 45.375 123.725 ;
        RECT 43.345 123.505 45.375 123.715 ;
        RECT 42.750 123.165 44.515 123.335 ;
        RECT 41.545 122.515 41.795 122.975 ;
        RECT 41.965 122.685 42.525 122.975 ;
        RECT 43.005 122.515 43.175 122.985 ;
        RECT 43.345 122.685 43.675 123.165 ;
        RECT 43.845 122.515 44.015 122.985 ;
        RECT 44.185 122.685 44.515 123.165 ;
        RECT 44.685 122.515 44.855 123.325 ;
        RECT 45.050 123.250 45.375 123.505 ;
        RECT 45.055 122.895 45.375 123.250 ;
        RECT 45.545 123.465 46.085 123.835 ;
        RECT 46.420 123.745 46.825 123.915 ;
        RECT 45.545 123.065 45.785 123.465 ;
        RECT 46.265 123.295 46.485 123.575 ;
        RECT 45.955 123.125 46.485 123.295 ;
        RECT 45.955 122.895 46.125 123.125 ;
        RECT 46.655 122.965 46.825 123.745 ;
        RECT 46.995 123.135 47.345 123.755 ;
        RECT 47.515 123.135 47.725 123.925 ;
        RECT 47.915 123.955 49.415 124.125 ;
        RECT 47.915 123.265 48.085 123.955 ;
        RECT 49.775 123.785 49.945 124.565 ;
        RECT 50.750 124.435 50.920 124.565 ;
        RECT 48.255 123.615 49.945 123.785 ;
        RECT 50.115 124.005 50.580 124.395 ;
        RECT 50.750 124.265 51.145 124.435 ;
        RECT 48.255 123.435 48.425 123.615 ;
        RECT 45.055 122.725 46.125 122.895 ;
        RECT 46.295 122.515 46.485 122.955 ;
        RECT 46.655 122.685 47.605 122.965 ;
        RECT 47.915 122.875 48.175 123.265 ;
        RECT 48.595 123.195 49.385 123.445 ;
        RECT 47.825 122.705 48.175 122.875 ;
        RECT 48.385 122.515 48.715 122.975 ;
        RECT 49.590 122.905 49.760 123.615 ;
        RECT 50.115 123.415 50.285 124.005 ;
        RECT 49.930 123.195 50.285 123.415 ;
        RECT 50.455 123.195 50.805 123.815 ;
        RECT 50.975 122.905 51.145 124.265 ;
        RECT 51.510 124.095 51.835 124.880 ;
        RECT 51.315 123.045 51.775 124.095 ;
        RECT 49.590 122.735 50.445 122.905 ;
        RECT 50.650 122.735 51.145 122.905 ;
        RECT 51.315 122.515 51.645 122.875 ;
        RECT 52.005 122.775 52.175 124.895 ;
        RECT 52.345 124.565 52.675 125.065 ;
        RECT 52.845 124.395 53.100 124.895 ;
        RECT 52.350 124.225 53.100 124.395 ;
        RECT 52.350 123.235 52.580 124.225 ;
        RECT 52.750 123.405 53.100 124.055 ;
        RECT 53.275 123.975 55.865 125.065 ;
        RECT 56.035 123.990 56.305 124.895 ;
        RECT 56.475 124.305 56.805 125.065 ;
        RECT 56.985 124.135 57.155 124.895 ;
        RECT 53.275 123.455 54.485 123.975 ;
        RECT 54.655 123.285 55.865 123.805 ;
        RECT 52.350 123.065 53.100 123.235 ;
        RECT 52.345 122.515 52.675 122.895 ;
        RECT 52.845 122.775 53.100 123.065 ;
        RECT 53.275 122.515 55.865 123.285 ;
        RECT 56.035 123.190 56.205 123.990 ;
        RECT 56.490 123.965 57.155 124.135 ;
        RECT 57.415 123.975 58.625 125.065 ;
        RECT 58.885 124.135 59.055 124.895 ;
        RECT 59.235 124.305 59.565 125.065 ;
        RECT 56.490 123.820 56.660 123.965 ;
        RECT 56.375 123.490 56.660 123.820 ;
        RECT 56.490 123.235 56.660 123.490 ;
        RECT 56.895 123.415 57.225 123.785 ;
        RECT 57.415 123.435 57.935 123.975 ;
        RECT 58.885 123.965 59.550 124.135 ;
        RECT 59.735 123.990 60.005 124.895 ;
        RECT 59.380 123.820 59.550 123.965 ;
        RECT 58.105 123.265 58.625 123.805 ;
        RECT 58.815 123.415 59.145 123.785 ;
        RECT 59.380 123.490 59.665 123.820 ;
        RECT 56.035 122.685 56.295 123.190 ;
        RECT 56.490 123.065 57.155 123.235 ;
        RECT 56.475 122.515 56.805 122.895 ;
        RECT 56.985 122.685 57.155 123.065 ;
        RECT 57.415 122.515 58.625 123.265 ;
        RECT 59.380 123.235 59.550 123.490 ;
        RECT 58.885 123.065 59.550 123.235 ;
        RECT 59.835 123.190 60.005 123.990 ;
        RECT 60.175 123.975 61.385 125.065 ;
        RECT 60.175 123.435 60.695 123.975 ;
        RECT 61.555 123.900 61.845 125.065 ;
        RECT 62.015 123.975 63.685 125.065 ;
        RECT 63.945 124.135 64.115 124.895 ;
        RECT 64.295 124.305 64.625 125.065 ;
        RECT 60.865 123.265 61.385 123.805 ;
        RECT 62.015 123.455 62.765 123.975 ;
        RECT 63.945 123.965 64.610 124.135 ;
        RECT 64.795 123.990 65.065 124.895 ;
        RECT 64.440 123.820 64.610 123.965 ;
        RECT 62.935 123.285 63.685 123.805 ;
        RECT 63.875 123.415 64.205 123.785 ;
        RECT 64.440 123.490 64.725 123.820 ;
        RECT 58.885 122.685 59.055 123.065 ;
        RECT 59.235 122.515 59.565 122.895 ;
        RECT 59.745 122.685 60.005 123.190 ;
        RECT 60.175 122.515 61.385 123.265 ;
        RECT 61.555 122.515 61.845 123.240 ;
        RECT 62.015 122.515 63.685 123.285 ;
        RECT 64.440 123.235 64.610 123.490 ;
        RECT 63.945 123.065 64.610 123.235 ;
        RECT 64.895 123.190 65.065 123.990 ;
        RECT 65.695 123.975 69.205 125.065 ;
        RECT 69.380 124.630 74.725 125.065 ;
        RECT 65.695 123.455 67.385 123.975 ;
        RECT 67.555 123.285 69.205 123.805 ;
        RECT 70.970 123.380 71.320 124.630 ;
        RECT 74.985 124.135 75.155 124.895 ;
        RECT 75.335 124.305 75.665 125.065 ;
        RECT 74.985 123.965 75.650 124.135 ;
        RECT 75.835 123.990 76.105 124.895 ;
        RECT 63.945 122.685 64.115 123.065 ;
        RECT 64.295 122.515 64.625 122.895 ;
        RECT 64.805 122.685 65.065 123.190 ;
        RECT 65.695 122.515 69.205 123.285 ;
        RECT 72.800 123.060 73.140 123.890 ;
        RECT 75.480 123.820 75.650 123.965 ;
        RECT 74.915 123.415 75.245 123.785 ;
        RECT 75.480 123.490 75.765 123.820 ;
        RECT 75.480 123.235 75.650 123.490 ;
        RECT 74.985 123.065 75.650 123.235 ;
        RECT 75.935 123.190 76.105 123.990 ;
        RECT 76.285 124.085 76.615 124.895 ;
        RECT 76.785 124.265 77.025 125.065 ;
        RECT 76.285 123.915 77.000 124.085 ;
        RECT 76.280 123.505 76.660 123.745 ;
        RECT 76.830 123.675 77.000 123.915 ;
        RECT 77.205 124.045 77.375 124.895 ;
        RECT 77.545 124.265 77.875 125.065 ;
        RECT 78.045 124.045 78.215 124.895 ;
        RECT 77.205 123.875 78.215 124.045 ;
        RECT 78.385 123.915 78.715 125.065 ;
        RECT 79.125 124.135 79.295 124.895 ;
        RECT 79.475 124.305 79.805 125.065 ;
        RECT 79.125 123.965 79.790 124.135 ;
        RECT 79.975 123.990 80.245 124.895 ;
        RECT 76.830 123.505 77.330 123.675 ;
        RECT 76.830 123.335 77.000 123.505 ;
        RECT 77.720 123.365 78.215 123.875 ;
        RECT 79.620 123.820 79.790 123.965 ;
        RECT 79.055 123.415 79.385 123.785 ;
        RECT 79.620 123.490 79.905 123.820 ;
        RECT 77.715 123.335 78.215 123.365 ;
        RECT 69.380 122.515 74.725 123.060 ;
        RECT 74.985 122.685 75.155 123.065 ;
        RECT 75.335 122.515 75.665 122.895 ;
        RECT 75.845 122.685 76.105 123.190 ;
        RECT 76.365 123.165 77.000 123.335 ;
        RECT 77.205 123.165 78.215 123.335 ;
        RECT 76.365 122.685 76.535 123.165 ;
        RECT 76.715 122.515 76.955 122.995 ;
        RECT 77.205 122.685 77.375 123.165 ;
        RECT 77.545 122.515 77.875 122.995 ;
        RECT 78.045 122.685 78.215 123.165 ;
        RECT 78.385 122.515 78.715 123.315 ;
        RECT 79.620 123.235 79.790 123.490 ;
        RECT 79.125 123.065 79.790 123.235 ;
        RECT 80.075 123.190 80.245 123.990 ;
        RECT 80.415 123.975 81.625 125.065 ;
        RECT 81.800 124.630 87.145 125.065 ;
        RECT 80.415 123.435 80.935 123.975 ;
        RECT 81.105 123.265 81.625 123.805 ;
        RECT 83.390 123.380 83.740 124.630 ;
        RECT 87.315 123.900 87.605 125.065 ;
        RECT 87.775 123.975 88.985 125.065 ;
        RECT 89.155 123.975 92.665 125.065 ;
        RECT 92.925 124.135 93.095 124.895 ;
        RECT 93.275 124.305 93.605 125.065 ;
        RECT 79.125 122.685 79.295 123.065 ;
        RECT 79.475 122.515 79.805 122.895 ;
        RECT 79.985 122.685 80.245 123.190 ;
        RECT 80.415 122.515 81.625 123.265 ;
        RECT 85.220 123.060 85.560 123.890 ;
        RECT 87.775 123.435 88.295 123.975 ;
        RECT 88.465 123.265 88.985 123.805 ;
        RECT 89.155 123.455 90.845 123.975 ;
        RECT 92.925 123.965 93.590 124.135 ;
        RECT 93.775 123.990 94.045 124.895 ;
        RECT 93.420 123.820 93.590 123.965 ;
        RECT 91.015 123.285 92.665 123.805 ;
        RECT 92.855 123.415 93.185 123.785 ;
        RECT 93.420 123.490 93.705 123.820 ;
        RECT 81.800 122.515 87.145 123.060 ;
        RECT 87.315 122.515 87.605 123.240 ;
        RECT 87.775 122.515 88.985 123.265 ;
        RECT 89.155 122.515 92.665 123.285 ;
        RECT 93.420 123.235 93.590 123.490 ;
        RECT 92.925 123.065 93.590 123.235 ;
        RECT 93.875 123.190 94.045 123.990 ;
        RECT 95.225 124.135 95.395 124.895 ;
        RECT 95.575 124.305 95.905 125.065 ;
        RECT 95.225 123.965 95.890 124.135 ;
        RECT 96.075 123.990 96.345 124.895 ;
        RECT 95.720 123.820 95.890 123.965 ;
        RECT 95.155 123.415 95.485 123.785 ;
        RECT 95.720 123.490 96.005 123.820 ;
        RECT 95.720 123.235 95.890 123.490 ;
        RECT 92.925 122.685 93.095 123.065 ;
        RECT 93.275 122.515 93.605 122.895 ;
        RECT 93.785 122.685 94.045 123.190 ;
        RECT 95.225 123.065 95.890 123.235 ;
        RECT 96.175 123.190 96.345 123.990 ;
        RECT 96.605 124.135 96.775 124.895 ;
        RECT 96.955 124.305 97.285 125.065 ;
        RECT 96.605 123.965 97.270 124.135 ;
        RECT 97.455 123.990 97.725 124.895 ;
        RECT 97.100 123.820 97.270 123.965 ;
        RECT 96.535 123.415 96.865 123.785 ;
        RECT 97.100 123.490 97.385 123.820 ;
        RECT 97.100 123.235 97.270 123.490 ;
        RECT 95.225 122.685 95.395 123.065 ;
        RECT 95.575 122.515 95.905 122.895 ;
        RECT 96.085 122.685 96.345 123.190 ;
        RECT 96.605 123.065 97.270 123.235 ;
        RECT 97.555 123.190 97.725 123.990 ;
        RECT 97.985 124.135 98.155 124.895 ;
        RECT 98.335 124.305 98.665 125.065 ;
        RECT 97.985 123.965 98.650 124.135 ;
        RECT 98.835 123.990 99.105 124.895 ;
        RECT 98.480 123.820 98.650 123.965 ;
        RECT 97.915 123.415 98.245 123.785 ;
        RECT 98.480 123.490 98.765 123.820 ;
        RECT 98.480 123.235 98.650 123.490 ;
        RECT 96.605 122.685 96.775 123.065 ;
        RECT 96.955 122.515 97.285 122.895 ;
        RECT 97.465 122.685 97.725 123.190 ;
        RECT 97.985 123.065 98.650 123.235 ;
        RECT 98.935 123.190 99.105 123.990 ;
        RECT 100.235 123.925 100.465 125.065 ;
        RECT 100.635 123.915 100.965 124.895 ;
        RECT 101.135 123.925 101.345 125.065 ;
        RECT 101.580 124.395 101.835 124.895 ;
        RECT 102.005 124.565 102.335 125.065 ;
        RECT 101.580 124.225 102.330 124.395 ;
        RECT 100.215 123.505 100.545 123.755 ;
        RECT 97.985 122.685 98.155 123.065 ;
        RECT 98.335 122.515 98.665 122.895 ;
        RECT 98.845 122.685 99.105 123.190 ;
        RECT 100.235 122.515 100.465 123.335 ;
        RECT 100.715 123.315 100.965 123.915 ;
        RECT 101.580 123.405 101.930 124.055 ;
        RECT 100.635 122.685 100.965 123.315 ;
        RECT 101.135 122.515 101.345 123.335 ;
        RECT 102.100 123.235 102.330 124.225 ;
        RECT 101.580 123.065 102.330 123.235 ;
        RECT 101.580 122.775 101.835 123.065 ;
        RECT 102.005 122.515 102.335 122.895 ;
        RECT 102.505 122.775 102.675 124.895 ;
        RECT 102.845 124.095 103.170 124.880 ;
        RECT 103.340 124.605 103.590 125.065 ;
        RECT 103.760 124.565 104.010 124.895 ;
        RECT 104.225 124.565 104.905 124.895 ;
        RECT 103.760 124.435 103.930 124.565 ;
        RECT 103.535 124.265 103.930 124.435 ;
        RECT 102.905 123.045 103.365 124.095 ;
        RECT 103.535 122.905 103.705 124.265 ;
        RECT 104.100 124.005 104.565 124.395 ;
        RECT 103.875 123.195 104.225 123.815 ;
        RECT 104.395 123.415 104.565 124.005 ;
        RECT 104.735 123.785 104.905 124.565 ;
        RECT 105.075 124.465 105.245 124.805 ;
        RECT 105.480 124.635 105.810 125.065 ;
        RECT 105.980 124.465 106.150 124.805 ;
        RECT 106.445 124.605 106.815 125.065 ;
        RECT 105.075 124.295 106.150 124.465 ;
        RECT 106.985 124.435 107.155 124.895 ;
        RECT 107.390 124.555 108.260 124.895 ;
        RECT 108.430 124.605 108.680 125.065 ;
        RECT 106.595 124.265 107.155 124.435 ;
        RECT 106.595 124.125 106.765 124.265 ;
        RECT 105.265 123.955 106.765 124.125 ;
        RECT 107.460 124.095 107.920 124.385 ;
        RECT 104.735 123.615 106.425 123.785 ;
        RECT 104.395 123.195 104.750 123.415 ;
        RECT 104.920 122.905 105.090 123.615 ;
        RECT 105.295 123.195 106.085 123.445 ;
        RECT 106.255 123.435 106.425 123.615 ;
        RECT 106.595 123.265 106.765 123.955 ;
        RECT 103.035 122.515 103.365 122.875 ;
        RECT 103.535 122.735 104.030 122.905 ;
        RECT 104.235 122.735 105.090 122.905 ;
        RECT 105.965 122.515 106.295 122.975 ;
        RECT 106.505 122.875 106.765 123.265 ;
        RECT 106.955 124.085 107.920 124.095 ;
        RECT 108.090 124.175 108.260 124.555 ;
        RECT 108.850 124.515 109.020 124.805 ;
        RECT 109.200 124.685 109.530 125.065 ;
        RECT 108.850 124.345 109.650 124.515 ;
        RECT 106.955 123.925 107.630 124.085 ;
        RECT 108.090 124.005 109.310 124.175 ;
        RECT 106.955 123.135 107.165 123.925 ;
        RECT 108.090 123.915 108.260 124.005 ;
        RECT 107.335 123.135 107.685 123.755 ;
        RECT 107.855 123.745 108.260 123.915 ;
        RECT 107.855 122.965 108.025 123.745 ;
        RECT 108.195 123.295 108.415 123.575 ;
        RECT 108.595 123.465 109.135 123.835 ;
        RECT 109.480 123.725 109.650 124.345 ;
        RECT 109.825 124.005 109.995 125.065 ;
        RECT 110.205 124.055 110.495 124.895 ;
        RECT 110.665 124.225 110.835 125.065 ;
        RECT 111.045 124.055 111.295 124.895 ;
        RECT 111.505 124.225 111.675 125.065 ;
        RECT 110.205 123.885 111.930 124.055 ;
        RECT 108.195 123.125 108.725 123.295 ;
        RECT 106.505 122.705 106.855 122.875 ;
        RECT 107.075 122.685 108.025 122.965 ;
        RECT 108.195 122.515 108.385 122.955 ;
        RECT 108.555 122.895 108.725 123.125 ;
        RECT 108.895 123.065 109.135 123.465 ;
        RECT 109.305 123.715 109.650 123.725 ;
        RECT 109.305 123.505 111.335 123.715 ;
        RECT 109.305 123.250 109.630 123.505 ;
        RECT 111.520 123.335 111.930 123.885 ;
        RECT 112.155 123.975 113.365 125.065 ;
        RECT 112.155 123.435 112.675 123.975 ;
        RECT 109.305 122.895 109.625 123.250 ;
        RECT 108.555 122.725 109.625 122.895 ;
        RECT 109.825 122.515 109.995 123.325 ;
        RECT 110.165 123.165 111.930 123.335 ;
        RECT 112.845 123.265 113.365 123.805 ;
        RECT 110.165 122.685 110.495 123.165 ;
        RECT 110.665 122.515 110.835 122.985 ;
        RECT 111.005 122.685 111.335 123.165 ;
        RECT 111.505 122.515 111.675 122.985 ;
        RECT 112.155 122.515 113.365 123.265 ;
        RECT 22.830 122.345 113.450 122.515 ;
        RECT 22.915 121.595 24.125 122.345 ;
        RECT 24.385 121.795 24.555 122.175 ;
        RECT 24.735 121.965 25.065 122.345 ;
        RECT 24.385 121.625 25.050 121.795 ;
        RECT 25.245 121.670 25.505 122.175 ;
        RECT 22.915 121.055 23.435 121.595 ;
        RECT 23.605 120.885 24.125 121.425 ;
        RECT 24.315 121.075 24.645 121.445 ;
        RECT 24.880 121.370 25.050 121.625 ;
        RECT 24.880 121.040 25.165 121.370 ;
        RECT 24.880 120.895 25.050 121.040 ;
        RECT 22.915 119.795 24.125 120.885 ;
        RECT 24.385 120.725 25.050 120.895 ;
        RECT 25.335 120.870 25.505 121.670 ;
        RECT 25.735 121.525 25.945 122.345 ;
        RECT 26.115 121.545 26.445 122.175 ;
        RECT 26.115 120.945 26.365 121.545 ;
        RECT 26.615 121.525 26.845 122.345 ;
        RECT 27.825 121.875 27.995 122.345 ;
        RECT 28.165 121.695 28.495 122.175 ;
        RECT 28.665 121.875 28.835 122.345 ;
        RECT 29.005 121.695 29.335 122.175 ;
        RECT 27.570 121.525 29.335 121.695 ;
        RECT 29.505 121.535 29.675 122.345 ;
        RECT 29.875 121.965 30.945 122.135 ;
        RECT 29.875 121.610 30.195 121.965 ;
        RECT 26.535 121.105 26.865 121.355 ;
        RECT 27.570 120.975 27.980 121.525 ;
        RECT 29.870 121.355 30.195 121.610 ;
        RECT 28.165 121.145 30.195 121.355 ;
        RECT 29.850 121.135 30.195 121.145 ;
        RECT 30.365 121.395 30.605 121.795 ;
        RECT 30.775 121.735 30.945 121.965 ;
        RECT 31.115 121.905 31.305 122.345 ;
        RECT 31.475 121.895 32.425 122.175 ;
        RECT 32.645 121.985 32.995 122.155 ;
        RECT 30.775 121.565 31.305 121.735 ;
        RECT 24.385 119.965 24.555 120.725 ;
        RECT 24.735 119.795 25.065 120.555 ;
        RECT 25.235 119.965 25.505 120.870 ;
        RECT 25.735 119.795 25.945 120.935 ;
        RECT 26.115 119.965 26.445 120.945 ;
        RECT 26.615 119.795 26.845 120.935 ;
        RECT 27.570 120.805 29.295 120.975 ;
        RECT 27.825 119.795 27.995 120.635 ;
        RECT 28.205 119.965 28.455 120.805 ;
        RECT 28.665 119.795 28.835 120.635 ;
        RECT 29.005 119.965 29.295 120.805 ;
        RECT 29.505 119.795 29.675 120.855 ;
        RECT 29.850 120.515 30.020 121.135 ;
        RECT 30.365 121.025 30.905 121.395 ;
        RECT 31.085 121.285 31.305 121.565 ;
        RECT 31.475 121.115 31.645 121.895 ;
        RECT 31.240 120.945 31.645 121.115 ;
        RECT 31.815 121.105 32.165 121.725 ;
        RECT 31.240 120.855 31.410 120.945 ;
        RECT 32.335 120.935 32.545 121.725 ;
        RECT 30.190 120.685 31.410 120.855 ;
        RECT 31.870 120.775 32.545 120.935 ;
        RECT 29.850 120.345 30.650 120.515 ;
        RECT 29.970 119.795 30.300 120.175 ;
        RECT 30.480 120.055 30.650 120.345 ;
        RECT 31.240 120.305 31.410 120.685 ;
        RECT 31.580 120.765 32.545 120.775 ;
        RECT 32.735 121.595 32.995 121.985 ;
        RECT 33.205 121.885 33.535 122.345 ;
        RECT 34.410 121.955 35.265 122.125 ;
        RECT 35.470 121.955 35.965 122.125 ;
        RECT 36.135 121.985 36.465 122.345 ;
        RECT 32.735 120.905 32.905 121.595 ;
        RECT 33.075 121.245 33.245 121.425 ;
        RECT 33.415 121.415 34.205 121.665 ;
        RECT 34.410 121.245 34.580 121.955 ;
        RECT 34.750 121.445 35.105 121.665 ;
        RECT 33.075 121.075 34.765 121.245 ;
        RECT 31.580 120.475 32.040 120.765 ;
        RECT 32.735 120.735 34.235 120.905 ;
        RECT 32.735 120.595 32.905 120.735 ;
        RECT 32.345 120.425 32.905 120.595 ;
        RECT 30.820 119.795 31.070 120.255 ;
        RECT 31.240 119.965 32.110 120.305 ;
        RECT 32.345 119.965 32.515 120.425 ;
        RECT 33.350 120.395 34.425 120.565 ;
        RECT 32.685 119.795 33.055 120.255 ;
        RECT 33.350 120.055 33.520 120.395 ;
        RECT 33.690 119.795 34.020 120.225 ;
        RECT 34.255 120.055 34.425 120.395 ;
        RECT 34.595 120.295 34.765 121.075 ;
        RECT 34.935 120.855 35.105 121.445 ;
        RECT 35.275 121.045 35.625 121.665 ;
        RECT 34.935 120.465 35.400 120.855 ;
        RECT 35.795 120.595 35.965 121.955 ;
        RECT 36.135 120.765 36.595 121.815 ;
        RECT 35.570 120.425 35.965 120.595 ;
        RECT 35.570 120.295 35.740 120.425 ;
        RECT 34.595 119.965 35.275 120.295 ;
        RECT 35.490 119.965 35.740 120.295 ;
        RECT 35.910 119.795 36.160 120.255 ;
        RECT 36.330 119.980 36.655 120.765 ;
        RECT 36.825 119.965 36.995 122.085 ;
        RECT 37.165 121.965 37.495 122.345 ;
        RECT 37.665 121.795 37.920 122.085 ;
        RECT 38.405 121.875 38.575 122.345 ;
        RECT 37.170 121.625 37.920 121.795 ;
        RECT 38.745 121.695 39.075 122.175 ;
        RECT 39.245 121.875 39.415 122.345 ;
        RECT 39.585 121.695 39.915 122.175 ;
        RECT 37.170 120.635 37.400 121.625 ;
        RECT 38.150 121.525 39.915 121.695 ;
        RECT 40.085 121.535 40.255 122.345 ;
        RECT 40.455 121.965 41.525 122.135 ;
        RECT 40.455 121.610 40.775 121.965 ;
        RECT 37.570 120.805 37.920 121.455 ;
        RECT 38.150 120.975 38.560 121.525 ;
        RECT 40.450 121.355 40.775 121.610 ;
        RECT 38.745 121.145 40.775 121.355 ;
        RECT 40.430 121.135 40.775 121.145 ;
        RECT 40.945 121.395 41.185 121.795 ;
        RECT 41.355 121.735 41.525 121.965 ;
        RECT 41.695 121.905 41.885 122.345 ;
        RECT 42.055 121.895 43.005 122.175 ;
        RECT 43.225 121.985 43.575 122.155 ;
        RECT 41.355 121.565 41.885 121.735 ;
        RECT 38.150 120.805 39.875 120.975 ;
        RECT 37.170 120.465 37.920 120.635 ;
        RECT 37.165 119.795 37.495 120.295 ;
        RECT 37.665 119.965 37.920 120.465 ;
        RECT 38.405 119.795 38.575 120.635 ;
        RECT 38.785 119.965 39.035 120.805 ;
        RECT 39.245 119.795 39.415 120.635 ;
        RECT 39.585 119.965 39.875 120.805 ;
        RECT 40.085 119.795 40.255 120.855 ;
        RECT 40.430 120.515 40.600 121.135 ;
        RECT 40.945 121.025 41.485 121.395 ;
        RECT 41.665 121.285 41.885 121.565 ;
        RECT 42.055 121.115 42.225 121.895 ;
        RECT 41.820 120.945 42.225 121.115 ;
        RECT 42.395 121.105 42.745 121.725 ;
        RECT 41.820 120.855 41.990 120.945 ;
        RECT 42.915 120.935 43.125 121.725 ;
        RECT 40.770 120.685 41.990 120.855 ;
        RECT 42.450 120.775 43.125 120.935 ;
        RECT 40.430 120.345 41.230 120.515 ;
        RECT 40.550 119.795 40.880 120.175 ;
        RECT 41.060 120.055 41.230 120.345 ;
        RECT 41.820 120.305 41.990 120.685 ;
        RECT 42.160 120.765 43.125 120.775 ;
        RECT 43.315 121.595 43.575 121.985 ;
        RECT 43.785 121.885 44.115 122.345 ;
        RECT 44.990 121.955 45.845 122.125 ;
        RECT 46.050 121.955 46.545 122.125 ;
        RECT 46.715 121.985 47.045 122.345 ;
        RECT 43.315 120.905 43.485 121.595 ;
        RECT 43.655 121.245 43.825 121.425 ;
        RECT 43.995 121.415 44.785 121.665 ;
        RECT 44.990 121.245 45.160 121.955 ;
        RECT 45.330 121.445 45.685 121.665 ;
        RECT 43.655 121.075 45.345 121.245 ;
        RECT 42.160 120.475 42.620 120.765 ;
        RECT 43.315 120.735 44.815 120.905 ;
        RECT 43.315 120.595 43.485 120.735 ;
        RECT 42.925 120.425 43.485 120.595 ;
        RECT 41.400 119.795 41.650 120.255 ;
        RECT 41.820 119.965 42.690 120.305 ;
        RECT 42.925 119.965 43.095 120.425 ;
        RECT 43.930 120.395 45.005 120.565 ;
        RECT 43.265 119.795 43.635 120.255 ;
        RECT 43.930 120.055 44.100 120.395 ;
        RECT 44.270 119.795 44.600 120.225 ;
        RECT 44.835 120.055 45.005 120.395 ;
        RECT 45.175 120.295 45.345 121.075 ;
        RECT 45.515 120.855 45.685 121.445 ;
        RECT 45.855 121.045 46.205 121.665 ;
        RECT 45.515 120.465 45.980 120.855 ;
        RECT 46.375 120.595 46.545 121.955 ;
        RECT 46.715 120.765 47.175 121.815 ;
        RECT 46.150 120.425 46.545 120.595 ;
        RECT 46.150 120.295 46.320 120.425 ;
        RECT 45.175 119.965 45.855 120.295 ;
        RECT 46.070 119.965 46.320 120.295 ;
        RECT 46.490 119.795 46.740 120.255 ;
        RECT 46.910 119.980 47.235 120.765 ;
        RECT 47.405 119.965 47.575 122.085 ;
        RECT 47.745 121.965 48.075 122.345 ;
        RECT 48.245 121.795 48.500 122.085 ;
        RECT 47.750 121.625 48.500 121.795 ;
        RECT 47.750 120.635 47.980 121.625 ;
        RECT 48.675 121.620 48.965 122.345 ;
        RECT 50.145 121.795 50.315 122.175 ;
        RECT 50.495 121.965 50.825 122.345 ;
        RECT 50.145 121.625 50.810 121.795 ;
        RECT 51.005 121.670 51.265 122.175 ;
        RECT 48.150 120.805 48.500 121.455 ;
        RECT 50.075 121.075 50.405 121.445 ;
        RECT 50.640 121.370 50.810 121.625 ;
        RECT 50.640 121.040 50.925 121.370 ;
        RECT 47.750 120.465 48.500 120.635 ;
        RECT 47.745 119.795 48.075 120.295 ;
        RECT 48.245 119.965 48.500 120.465 ;
        RECT 48.675 119.795 48.965 120.960 ;
        RECT 50.640 120.895 50.810 121.040 ;
        RECT 50.145 120.725 50.810 120.895 ;
        RECT 51.095 120.870 51.265 121.670 ;
        RECT 51.955 121.525 52.165 122.345 ;
        RECT 52.335 121.545 52.665 122.175 ;
        RECT 52.335 120.945 52.585 121.545 ;
        RECT 52.835 121.525 53.065 122.345 ;
        RECT 54.195 121.670 54.455 122.175 ;
        RECT 54.635 121.965 54.965 122.345 ;
        RECT 55.145 121.795 55.315 122.175 ;
        RECT 52.755 121.105 53.085 121.355 ;
        RECT 50.145 119.965 50.315 120.725 ;
        RECT 50.495 119.795 50.825 120.555 ;
        RECT 50.995 119.965 51.265 120.870 ;
        RECT 51.955 119.795 52.165 120.935 ;
        RECT 52.335 119.965 52.665 120.945 ;
        RECT 52.835 119.795 53.065 120.935 ;
        RECT 54.195 120.870 54.365 121.670 ;
        RECT 54.650 121.625 55.315 121.795 ;
        RECT 55.665 121.695 55.835 122.175 ;
        RECT 56.015 121.865 56.255 122.345 ;
        RECT 56.505 121.695 56.675 122.175 ;
        RECT 56.845 121.865 57.175 122.345 ;
        RECT 57.345 121.695 57.515 122.175 ;
        RECT 54.650 121.370 54.820 121.625 ;
        RECT 55.665 121.525 56.300 121.695 ;
        RECT 56.505 121.525 57.515 121.695 ;
        RECT 57.685 121.545 58.015 122.345 ;
        RECT 58.645 121.875 58.815 122.345 ;
        RECT 58.985 121.695 59.315 122.175 ;
        RECT 59.485 121.875 59.655 122.345 ;
        RECT 59.825 121.695 60.155 122.175 ;
        RECT 54.535 121.040 54.820 121.370 ;
        RECT 55.055 121.075 55.385 121.445 ;
        RECT 56.130 121.355 56.300 121.525 ;
        RECT 55.580 121.115 55.960 121.355 ;
        RECT 56.130 121.185 56.630 121.355 ;
        RECT 54.650 120.895 54.820 121.040 ;
        RECT 56.130 120.945 56.300 121.185 ;
        RECT 57.020 120.985 57.515 121.525 ;
        RECT 54.195 119.965 54.465 120.870 ;
        RECT 54.650 120.725 55.315 120.895 ;
        RECT 54.635 119.795 54.965 120.555 ;
        RECT 55.145 119.965 55.315 120.725 ;
        RECT 55.585 120.775 56.300 120.945 ;
        RECT 56.505 120.815 57.515 120.985 ;
        RECT 58.390 121.525 60.155 121.695 ;
        RECT 60.325 121.535 60.495 122.345 ;
        RECT 60.695 121.965 61.765 122.135 ;
        RECT 60.695 121.610 61.015 121.965 ;
        RECT 58.390 120.975 58.800 121.525 ;
        RECT 60.690 121.355 61.015 121.610 ;
        RECT 58.985 121.145 61.015 121.355 ;
        RECT 60.670 121.135 61.015 121.145 ;
        RECT 61.185 121.395 61.425 121.795 ;
        RECT 61.595 121.735 61.765 121.965 ;
        RECT 61.935 121.905 62.125 122.345 ;
        RECT 62.295 121.895 63.245 122.175 ;
        RECT 63.465 121.985 63.815 122.155 ;
        RECT 61.595 121.565 62.125 121.735 ;
        RECT 55.585 119.965 55.915 120.775 ;
        RECT 56.085 119.795 56.325 120.595 ;
        RECT 56.505 119.965 56.675 120.815 ;
        RECT 56.845 119.795 57.175 120.595 ;
        RECT 57.345 119.965 57.515 120.815 ;
        RECT 57.685 119.795 58.015 120.945 ;
        RECT 58.390 120.805 60.115 120.975 ;
        RECT 58.645 119.795 58.815 120.635 ;
        RECT 59.025 119.965 59.275 120.805 ;
        RECT 59.485 119.795 59.655 120.635 ;
        RECT 59.825 119.965 60.115 120.805 ;
        RECT 60.325 119.795 60.495 120.855 ;
        RECT 60.670 120.515 60.840 121.135 ;
        RECT 61.185 121.025 61.725 121.395 ;
        RECT 61.905 121.285 62.125 121.565 ;
        RECT 62.295 121.115 62.465 121.895 ;
        RECT 62.060 120.945 62.465 121.115 ;
        RECT 62.635 121.105 62.985 121.725 ;
        RECT 62.060 120.855 62.230 120.945 ;
        RECT 63.155 120.935 63.365 121.725 ;
        RECT 61.010 120.685 62.230 120.855 ;
        RECT 62.690 120.775 63.365 120.935 ;
        RECT 60.670 120.345 61.470 120.515 ;
        RECT 60.790 119.795 61.120 120.175 ;
        RECT 61.300 120.055 61.470 120.345 ;
        RECT 62.060 120.305 62.230 120.685 ;
        RECT 62.400 120.765 63.365 120.775 ;
        RECT 63.555 121.595 63.815 121.985 ;
        RECT 64.025 121.885 64.355 122.345 ;
        RECT 65.230 121.955 66.085 122.125 ;
        RECT 66.290 121.955 66.785 122.125 ;
        RECT 66.955 121.985 67.285 122.345 ;
        RECT 63.555 120.905 63.725 121.595 ;
        RECT 63.895 121.245 64.065 121.425 ;
        RECT 64.235 121.415 65.025 121.665 ;
        RECT 65.230 121.245 65.400 121.955 ;
        RECT 65.570 121.445 65.925 121.665 ;
        RECT 63.895 121.075 65.585 121.245 ;
        RECT 62.400 120.475 62.860 120.765 ;
        RECT 63.555 120.735 65.055 120.905 ;
        RECT 63.555 120.595 63.725 120.735 ;
        RECT 63.165 120.425 63.725 120.595 ;
        RECT 61.640 119.795 61.890 120.255 ;
        RECT 62.060 119.965 62.930 120.305 ;
        RECT 63.165 119.965 63.335 120.425 ;
        RECT 64.170 120.395 65.245 120.565 ;
        RECT 63.505 119.795 63.875 120.255 ;
        RECT 64.170 120.055 64.340 120.395 ;
        RECT 64.510 119.795 64.840 120.225 ;
        RECT 65.075 120.055 65.245 120.395 ;
        RECT 65.415 120.295 65.585 121.075 ;
        RECT 65.755 120.855 65.925 121.445 ;
        RECT 66.095 121.045 66.445 121.665 ;
        RECT 65.755 120.465 66.220 120.855 ;
        RECT 66.615 120.595 66.785 121.955 ;
        RECT 66.955 120.765 67.415 121.815 ;
        RECT 66.390 120.425 66.785 120.595 ;
        RECT 66.390 120.295 66.560 120.425 ;
        RECT 65.415 119.965 66.095 120.295 ;
        RECT 66.310 119.965 66.560 120.295 ;
        RECT 66.730 119.795 66.980 120.255 ;
        RECT 67.150 119.980 67.475 120.765 ;
        RECT 67.645 119.965 67.815 122.085 ;
        RECT 67.985 121.965 68.315 122.345 ;
        RECT 68.485 121.795 68.740 122.085 ;
        RECT 67.990 121.625 68.740 121.795 ;
        RECT 69.005 121.795 69.175 122.175 ;
        RECT 69.355 121.965 69.685 122.345 ;
        RECT 69.005 121.625 69.670 121.795 ;
        RECT 69.865 121.670 70.125 122.175 ;
        RECT 67.990 120.635 68.220 121.625 ;
        RECT 68.390 120.805 68.740 121.455 ;
        RECT 68.935 121.075 69.265 121.445 ;
        RECT 69.500 121.370 69.670 121.625 ;
        RECT 69.500 121.040 69.785 121.370 ;
        RECT 69.500 120.895 69.670 121.040 ;
        RECT 69.005 120.725 69.670 120.895 ;
        RECT 69.955 120.870 70.125 121.670 ;
        RECT 70.385 121.795 70.555 122.175 ;
        RECT 70.735 121.965 71.065 122.345 ;
        RECT 70.385 121.625 71.050 121.795 ;
        RECT 71.245 121.670 71.505 122.175 ;
        RECT 70.315 121.075 70.645 121.445 ;
        RECT 70.880 121.370 71.050 121.625 ;
        RECT 70.880 121.040 71.165 121.370 ;
        RECT 70.880 120.895 71.050 121.040 ;
        RECT 67.990 120.465 68.740 120.635 ;
        RECT 67.985 119.795 68.315 120.295 ;
        RECT 68.485 119.965 68.740 120.465 ;
        RECT 69.005 119.965 69.175 120.725 ;
        RECT 69.355 119.795 69.685 120.555 ;
        RECT 69.855 119.965 70.125 120.870 ;
        RECT 70.385 120.725 71.050 120.895 ;
        RECT 71.335 120.870 71.505 121.670 ;
        RECT 71.765 121.795 71.935 122.175 ;
        RECT 72.115 121.965 72.445 122.345 ;
        RECT 71.765 121.625 72.430 121.795 ;
        RECT 72.625 121.670 72.885 122.175 ;
        RECT 71.695 121.075 72.025 121.445 ;
        RECT 72.260 121.370 72.430 121.625 ;
        RECT 72.260 121.040 72.545 121.370 ;
        RECT 72.260 120.895 72.430 121.040 ;
        RECT 70.385 119.965 70.555 120.725 ;
        RECT 70.735 119.795 71.065 120.555 ;
        RECT 71.235 119.965 71.505 120.870 ;
        RECT 71.765 120.725 72.430 120.895 ;
        RECT 72.715 120.870 72.885 121.670 ;
        RECT 73.115 121.525 73.325 122.345 ;
        RECT 73.495 121.545 73.825 122.175 ;
        RECT 73.495 120.945 73.745 121.545 ;
        RECT 73.995 121.525 74.225 122.345 ;
        RECT 74.435 121.620 74.725 122.345 ;
        RECT 75.205 121.875 75.375 122.345 ;
        RECT 75.545 121.695 75.875 122.175 ;
        RECT 76.045 121.875 76.215 122.345 ;
        RECT 76.385 121.695 76.715 122.175 ;
        RECT 74.950 121.525 76.715 121.695 ;
        RECT 76.885 121.535 77.055 122.345 ;
        RECT 77.255 121.965 78.325 122.135 ;
        RECT 77.255 121.610 77.575 121.965 ;
        RECT 73.915 121.105 74.245 121.355 ;
        RECT 74.950 120.975 75.360 121.525 ;
        RECT 77.250 121.355 77.575 121.610 ;
        RECT 75.545 121.145 77.575 121.355 ;
        RECT 77.230 121.135 77.575 121.145 ;
        RECT 77.745 121.395 77.985 121.795 ;
        RECT 78.155 121.735 78.325 121.965 ;
        RECT 78.495 121.905 78.685 122.345 ;
        RECT 78.855 121.895 79.805 122.175 ;
        RECT 80.025 121.985 80.375 122.155 ;
        RECT 78.155 121.565 78.685 121.735 ;
        RECT 71.765 119.965 71.935 120.725 ;
        RECT 72.115 119.795 72.445 120.555 ;
        RECT 72.615 119.965 72.885 120.870 ;
        RECT 73.115 119.795 73.325 120.935 ;
        RECT 73.495 119.965 73.825 120.945 ;
        RECT 73.995 119.795 74.225 120.935 ;
        RECT 74.435 119.795 74.725 120.960 ;
        RECT 74.950 120.805 76.675 120.975 ;
        RECT 75.205 119.795 75.375 120.635 ;
        RECT 75.585 119.965 75.835 120.805 ;
        RECT 76.045 119.795 76.215 120.635 ;
        RECT 76.385 119.965 76.675 120.805 ;
        RECT 76.885 119.795 77.055 120.855 ;
        RECT 77.230 120.515 77.400 121.135 ;
        RECT 77.745 121.025 78.285 121.395 ;
        RECT 78.465 121.285 78.685 121.565 ;
        RECT 78.855 121.115 79.025 121.895 ;
        RECT 78.620 120.945 79.025 121.115 ;
        RECT 79.195 121.105 79.545 121.725 ;
        RECT 78.620 120.855 78.790 120.945 ;
        RECT 79.715 120.935 79.925 121.725 ;
        RECT 77.570 120.685 78.790 120.855 ;
        RECT 79.250 120.775 79.925 120.935 ;
        RECT 77.230 120.345 78.030 120.515 ;
        RECT 77.350 119.795 77.680 120.175 ;
        RECT 77.860 120.055 78.030 120.345 ;
        RECT 78.620 120.305 78.790 120.685 ;
        RECT 78.960 120.765 79.925 120.775 ;
        RECT 80.115 121.595 80.375 121.985 ;
        RECT 80.585 121.885 80.915 122.345 ;
        RECT 81.790 121.955 82.645 122.125 ;
        RECT 82.850 121.955 83.345 122.125 ;
        RECT 83.515 121.985 83.845 122.345 ;
        RECT 80.115 120.905 80.285 121.595 ;
        RECT 80.455 121.245 80.625 121.425 ;
        RECT 80.795 121.415 81.585 121.665 ;
        RECT 81.790 121.245 81.960 121.955 ;
        RECT 82.130 121.445 82.485 121.665 ;
        RECT 80.455 121.075 82.145 121.245 ;
        RECT 78.960 120.475 79.420 120.765 ;
        RECT 80.115 120.735 81.615 120.905 ;
        RECT 80.115 120.595 80.285 120.735 ;
        RECT 79.725 120.425 80.285 120.595 ;
        RECT 78.200 119.795 78.450 120.255 ;
        RECT 78.620 119.965 79.490 120.305 ;
        RECT 79.725 119.965 79.895 120.425 ;
        RECT 80.730 120.395 81.805 120.565 ;
        RECT 80.065 119.795 80.435 120.255 ;
        RECT 80.730 120.055 80.900 120.395 ;
        RECT 81.070 119.795 81.400 120.225 ;
        RECT 81.635 120.055 81.805 120.395 ;
        RECT 81.975 120.295 82.145 121.075 ;
        RECT 82.315 120.855 82.485 121.445 ;
        RECT 82.655 121.045 83.005 121.665 ;
        RECT 82.315 120.465 82.780 120.855 ;
        RECT 83.175 120.595 83.345 121.955 ;
        RECT 83.515 120.765 83.975 121.815 ;
        RECT 82.950 120.425 83.345 120.595 ;
        RECT 82.950 120.295 83.120 120.425 ;
        RECT 81.975 119.965 82.655 120.295 ;
        RECT 82.870 119.965 83.120 120.295 ;
        RECT 83.290 119.795 83.540 120.255 ;
        RECT 83.710 119.980 84.035 120.765 ;
        RECT 84.205 119.965 84.375 122.085 ;
        RECT 84.545 121.965 84.875 122.345 ;
        RECT 85.045 121.795 85.300 122.085 ;
        RECT 84.550 121.625 85.300 121.795 ;
        RECT 86.485 121.795 86.655 122.175 ;
        RECT 86.835 121.965 87.165 122.345 ;
        RECT 86.485 121.625 87.150 121.795 ;
        RECT 87.345 121.670 87.605 122.175 ;
        RECT 88.085 121.875 88.255 122.345 ;
        RECT 88.425 121.695 88.755 122.175 ;
        RECT 88.925 121.875 89.095 122.345 ;
        RECT 89.265 121.695 89.595 122.175 ;
        RECT 84.550 120.635 84.780 121.625 ;
        RECT 84.950 120.805 85.300 121.455 ;
        RECT 86.415 121.075 86.745 121.445 ;
        RECT 86.980 121.370 87.150 121.625 ;
        RECT 86.980 121.040 87.265 121.370 ;
        RECT 86.980 120.895 87.150 121.040 ;
        RECT 86.485 120.725 87.150 120.895 ;
        RECT 87.435 120.870 87.605 121.670 ;
        RECT 84.550 120.465 85.300 120.635 ;
        RECT 84.545 119.795 84.875 120.295 ;
        RECT 85.045 119.965 85.300 120.465 ;
        RECT 86.485 119.965 86.655 120.725 ;
        RECT 86.835 119.795 87.165 120.555 ;
        RECT 87.335 119.965 87.605 120.870 ;
        RECT 87.830 121.525 89.595 121.695 ;
        RECT 89.765 121.535 89.935 122.345 ;
        RECT 90.135 121.965 91.205 122.135 ;
        RECT 90.135 121.610 90.455 121.965 ;
        RECT 87.830 120.975 88.240 121.525 ;
        RECT 90.130 121.355 90.455 121.610 ;
        RECT 88.425 121.145 90.455 121.355 ;
        RECT 90.110 121.135 90.455 121.145 ;
        RECT 90.625 121.395 90.865 121.795 ;
        RECT 91.035 121.735 91.205 121.965 ;
        RECT 91.375 121.905 91.565 122.345 ;
        RECT 91.735 121.895 92.685 122.175 ;
        RECT 92.905 121.985 93.255 122.155 ;
        RECT 91.035 121.565 91.565 121.735 ;
        RECT 87.830 120.805 89.555 120.975 ;
        RECT 88.085 119.795 88.255 120.635 ;
        RECT 88.465 119.965 88.715 120.805 ;
        RECT 88.925 119.795 89.095 120.635 ;
        RECT 89.265 119.965 89.555 120.805 ;
        RECT 89.765 119.795 89.935 120.855 ;
        RECT 90.110 120.515 90.280 121.135 ;
        RECT 90.625 121.025 91.165 121.395 ;
        RECT 91.345 121.285 91.565 121.565 ;
        RECT 91.735 121.115 91.905 121.895 ;
        RECT 91.500 120.945 91.905 121.115 ;
        RECT 92.075 121.105 92.425 121.725 ;
        RECT 91.500 120.855 91.670 120.945 ;
        RECT 92.595 120.935 92.805 121.725 ;
        RECT 90.450 120.685 91.670 120.855 ;
        RECT 92.130 120.775 92.805 120.935 ;
        RECT 90.110 120.345 90.910 120.515 ;
        RECT 90.230 119.795 90.560 120.175 ;
        RECT 90.740 120.055 90.910 120.345 ;
        RECT 91.500 120.305 91.670 120.685 ;
        RECT 91.840 120.765 92.805 120.775 ;
        RECT 92.995 121.595 93.255 121.985 ;
        RECT 93.465 121.885 93.795 122.345 ;
        RECT 94.670 121.955 95.525 122.125 ;
        RECT 95.730 121.955 96.225 122.125 ;
        RECT 96.395 121.985 96.725 122.345 ;
        RECT 92.995 120.905 93.165 121.595 ;
        RECT 93.335 121.245 93.505 121.425 ;
        RECT 93.675 121.415 94.465 121.665 ;
        RECT 94.670 121.245 94.840 121.955 ;
        RECT 95.010 121.445 95.365 121.665 ;
        RECT 93.335 121.075 95.025 121.245 ;
        RECT 91.840 120.475 92.300 120.765 ;
        RECT 92.995 120.735 94.495 120.905 ;
        RECT 92.995 120.595 93.165 120.735 ;
        RECT 92.605 120.425 93.165 120.595 ;
        RECT 91.080 119.795 91.330 120.255 ;
        RECT 91.500 119.965 92.370 120.305 ;
        RECT 92.605 119.965 92.775 120.425 ;
        RECT 93.610 120.395 94.685 120.565 ;
        RECT 92.945 119.795 93.315 120.255 ;
        RECT 93.610 120.055 93.780 120.395 ;
        RECT 93.950 119.795 94.280 120.225 ;
        RECT 94.515 120.055 94.685 120.395 ;
        RECT 94.855 120.295 95.025 121.075 ;
        RECT 95.195 120.855 95.365 121.445 ;
        RECT 95.535 121.045 95.885 121.665 ;
        RECT 95.195 120.465 95.660 120.855 ;
        RECT 96.055 120.595 96.225 121.955 ;
        RECT 96.395 120.765 96.855 121.815 ;
        RECT 95.830 120.425 96.225 120.595 ;
        RECT 95.830 120.295 96.000 120.425 ;
        RECT 94.855 119.965 95.535 120.295 ;
        RECT 95.750 119.965 96.000 120.295 ;
        RECT 96.170 119.795 96.420 120.255 ;
        RECT 96.590 119.980 96.915 120.765 ;
        RECT 97.085 119.965 97.255 122.085 ;
        RECT 97.425 121.965 97.755 122.345 ;
        RECT 97.925 121.795 98.180 122.085 ;
        RECT 97.430 121.625 98.180 121.795 ;
        RECT 98.355 121.670 98.615 122.175 ;
        RECT 98.795 121.965 99.125 122.345 ;
        RECT 99.305 121.795 99.475 122.175 ;
        RECT 97.430 120.635 97.660 121.625 ;
        RECT 97.830 120.805 98.180 121.455 ;
        RECT 98.355 120.870 98.525 121.670 ;
        RECT 98.810 121.625 99.475 121.795 ;
        RECT 98.810 121.370 98.980 121.625 ;
        RECT 100.195 121.620 100.485 122.345 ;
        RECT 101.580 121.795 101.835 122.085 ;
        RECT 102.005 121.965 102.335 122.345 ;
        RECT 101.580 121.625 102.330 121.795 ;
        RECT 98.695 121.040 98.980 121.370 ;
        RECT 99.215 121.075 99.545 121.445 ;
        RECT 98.810 120.895 98.980 121.040 ;
        RECT 97.430 120.465 98.180 120.635 ;
        RECT 97.425 119.795 97.755 120.295 ;
        RECT 97.925 119.965 98.180 120.465 ;
        RECT 98.355 119.965 98.625 120.870 ;
        RECT 98.810 120.725 99.475 120.895 ;
        RECT 98.795 119.795 99.125 120.555 ;
        RECT 99.305 119.965 99.475 120.725 ;
        RECT 100.195 119.795 100.485 120.960 ;
        RECT 101.580 120.805 101.930 121.455 ;
        RECT 102.100 120.635 102.330 121.625 ;
        RECT 101.580 120.465 102.330 120.635 ;
        RECT 101.580 119.965 101.835 120.465 ;
        RECT 102.005 119.795 102.335 120.295 ;
        RECT 102.505 119.965 102.675 122.085 ;
        RECT 103.035 121.985 103.365 122.345 ;
        RECT 103.535 121.955 104.030 122.125 ;
        RECT 104.235 121.955 105.090 122.125 ;
        RECT 102.905 120.765 103.365 121.815 ;
        RECT 102.845 119.980 103.170 120.765 ;
        RECT 103.535 120.595 103.705 121.955 ;
        RECT 103.875 121.045 104.225 121.665 ;
        RECT 104.395 121.445 104.750 121.665 ;
        RECT 104.395 120.855 104.565 121.445 ;
        RECT 104.920 121.245 105.090 121.955 ;
        RECT 105.965 121.885 106.295 122.345 ;
        RECT 106.505 121.985 106.855 122.155 ;
        RECT 105.295 121.415 106.085 121.665 ;
        RECT 106.505 121.595 106.765 121.985 ;
        RECT 107.075 121.895 108.025 122.175 ;
        RECT 108.195 121.905 108.385 122.345 ;
        RECT 108.555 121.965 109.625 122.135 ;
        RECT 106.255 121.245 106.425 121.425 ;
        RECT 103.535 120.425 103.930 120.595 ;
        RECT 104.100 120.465 104.565 120.855 ;
        RECT 104.735 121.075 106.425 121.245 ;
        RECT 103.760 120.295 103.930 120.425 ;
        RECT 104.735 120.295 104.905 121.075 ;
        RECT 106.595 120.905 106.765 121.595 ;
        RECT 105.265 120.735 106.765 120.905 ;
        RECT 106.955 120.935 107.165 121.725 ;
        RECT 107.335 121.105 107.685 121.725 ;
        RECT 107.855 121.115 108.025 121.895 ;
        RECT 108.555 121.735 108.725 121.965 ;
        RECT 108.195 121.565 108.725 121.735 ;
        RECT 108.195 121.285 108.415 121.565 ;
        RECT 108.895 121.395 109.135 121.795 ;
        RECT 107.855 120.945 108.260 121.115 ;
        RECT 108.595 121.025 109.135 121.395 ;
        RECT 109.305 121.610 109.625 121.965 ;
        RECT 109.305 121.355 109.630 121.610 ;
        RECT 109.825 121.535 109.995 122.345 ;
        RECT 110.165 121.695 110.495 122.175 ;
        RECT 110.665 121.875 110.835 122.345 ;
        RECT 111.005 121.695 111.335 122.175 ;
        RECT 111.505 121.875 111.675 122.345 ;
        RECT 110.165 121.525 111.930 121.695 ;
        RECT 112.155 121.595 113.365 122.345 ;
        RECT 109.305 121.145 111.335 121.355 ;
        RECT 109.305 121.135 109.650 121.145 ;
        RECT 106.955 120.775 107.630 120.935 ;
        RECT 108.090 120.855 108.260 120.945 ;
        RECT 106.955 120.765 107.920 120.775 ;
        RECT 106.595 120.595 106.765 120.735 ;
        RECT 103.340 119.795 103.590 120.255 ;
        RECT 103.760 119.965 104.010 120.295 ;
        RECT 104.225 119.965 104.905 120.295 ;
        RECT 105.075 120.395 106.150 120.565 ;
        RECT 106.595 120.425 107.155 120.595 ;
        RECT 107.460 120.475 107.920 120.765 ;
        RECT 108.090 120.685 109.310 120.855 ;
        RECT 105.075 120.055 105.245 120.395 ;
        RECT 105.480 119.795 105.810 120.225 ;
        RECT 105.980 120.055 106.150 120.395 ;
        RECT 106.445 119.795 106.815 120.255 ;
        RECT 106.985 119.965 107.155 120.425 ;
        RECT 108.090 120.305 108.260 120.685 ;
        RECT 109.480 120.515 109.650 121.135 ;
        RECT 111.520 120.975 111.930 121.525 ;
        RECT 107.390 119.965 108.260 120.305 ;
        RECT 108.850 120.345 109.650 120.515 ;
        RECT 108.430 119.795 108.680 120.255 ;
        RECT 108.850 120.055 109.020 120.345 ;
        RECT 109.200 119.795 109.530 120.175 ;
        RECT 109.825 119.795 109.995 120.855 ;
        RECT 110.205 120.805 111.930 120.975 ;
        RECT 112.155 120.885 112.675 121.425 ;
        RECT 112.845 121.055 113.365 121.595 ;
        RECT 110.205 119.965 110.495 120.805 ;
        RECT 110.665 119.795 110.835 120.635 ;
        RECT 111.045 119.965 111.295 120.805 ;
        RECT 111.505 119.795 111.675 120.635 ;
        RECT 112.155 119.795 113.365 120.885 ;
        RECT 22.830 119.625 113.450 119.795 ;
        RECT 22.915 118.535 24.125 119.625 ;
        RECT 25.220 118.955 25.475 119.455 ;
        RECT 25.645 119.125 25.975 119.625 ;
        RECT 25.220 118.785 25.970 118.955 ;
        RECT 22.915 117.825 23.435 118.365 ;
        RECT 23.605 117.995 24.125 118.535 ;
        RECT 25.220 117.965 25.570 118.615 ;
        RECT 22.915 117.075 24.125 117.825 ;
        RECT 25.740 117.795 25.970 118.785 ;
        RECT 25.220 117.625 25.970 117.795 ;
        RECT 25.220 117.335 25.475 117.625 ;
        RECT 25.645 117.075 25.975 117.455 ;
        RECT 26.145 117.335 26.315 119.455 ;
        RECT 26.485 118.655 26.810 119.440 ;
        RECT 26.980 119.165 27.230 119.625 ;
        RECT 27.400 119.125 27.650 119.455 ;
        RECT 27.865 119.125 28.545 119.455 ;
        RECT 27.400 118.995 27.570 119.125 ;
        RECT 27.175 118.825 27.570 118.995 ;
        RECT 26.545 117.605 27.005 118.655 ;
        RECT 27.175 117.465 27.345 118.825 ;
        RECT 27.740 118.565 28.205 118.955 ;
        RECT 27.515 117.755 27.865 118.375 ;
        RECT 28.035 117.975 28.205 118.565 ;
        RECT 28.375 118.345 28.545 119.125 ;
        RECT 28.715 119.025 28.885 119.365 ;
        RECT 29.120 119.195 29.450 119.625 ;
        RECT 29.620 119.025 29.790 119.365 ;
        RECT 30.085 119.165 30.455 119.625 ;
        RECT 28.715 118.855 29.790 119.025 ;
        RECT 30.625 118.995 30.795 119.455 ;
        RECT 31.030 119.115 31.900 119.455 ;
        RECT 32.070 119.165 32.320 119.625 ;
        RECT 30.235 118.825 30.795 118.995 ;
        RECT 30.235 118.685 30.405 118.825 ;
        RECT 28.905 118.515 30.405 118.685 ;
        RECT 31.100 118.655 31.560 118.945 ;
        RECT 28.375 118.175 30.065 118.345 ;
        RECT 28.035 117.755 28.390 117.975 ;
        RECT 28.560 117.465 28.730 118.175 ;
        RECT 28.935 117.755 29.725 118.005 ;
        RECT 29.895 117.995 30.065 118.175 ;
        RECT 30.235 117.825 30.405 118.515 ;
        RECT 26.675 117.075 27.005 117.435 ;
        RECT 27.175 117.295 27.670 117.465 ;
        RECT 27.875 117.295 28.730 117.465 ;
        RECT 29.605 117.075 29.935 117.535 ;
        RECT 30.145 117.435 30.405 117.825 ;
        RECT 30.595 118.645 31.560 118.655 ;
        RECT 31.730 118.735 31.900 119.115 ;
        RECT 32.490 119.075 32.660 119.365 ;
        RECT 32.840 119.245 33.170 119.625 ;
        RECT 32.490 118.905 33.290 119.075 ;
        RECT 30.595 118.485 31.270 118.645 ;
        RECT 31.730 118.565 32.950 118.735 ;
        RECT 30.595 117.695 30.805 118.485 ;
        RECT 31.730 118.475 31.900 118.565 ;
        RECT 30.975 117.695 31.325 118.315 ;
        RECT 31.495 118.305 31.900 118.475 ;
        RECT 31.495 117.525 31.665 118.305 ;
        RECT 31.835 117.855 32.055 118.135 ;
        RECT 32.235 118.025 32.775 118.395 ;
        RECT 33.120 118.285 33.290 118.905 ;
        RECT 33.465 118.565 33.635 119.625 ;
        RECT 33.845 118.615 34.135 119.455 ;
        RECT 34.305 118.785 34.475 119.625 ;
        RECT 34.685 118.615 34.935 119.455 ;
        RECT 35.145 118.785 35.315 119.625 ;
        RECT 33.845 118.445 35.570 118.615 ;
        RECT 35.795 118.460 36.085 119.625 ;
        RECT 36.295 118.485 36.525 119.625 ;
        RECT 36.695 118.475 37.025 119.455 ;
        RECT 37.195 118.485 37.405 119.625 ;
        RECT 37.635 118.550 37.905 119.455 ;
        RECT 38.075 118.865 38.405 119.625 ;
        RECT 38.585 118.695 38.755 119.455 ;
        RECT 31.835 117.685 32.365 117.855 ;
        RECT 30.145 117.265 30.495 117.435 ;
        RECT 30.715 117.245 31.665 117.525 ;
        RECT 31.835 117.075 32.025 117.515 ;
        RECT 32.195 117.455 32.365 117.685 ;
        RECT 32.535 117.625 32.775 118.025 ;
        RECT 32.945 118.275 33.290 118.285 ;
        RECT 32.945 118.065 34.975 118.275 ;
        RECT 32.945 117.810 33.270 118.065 ;
        RECT 35.160 117.895 35.570 118.445 ;
        RECT 36.275 118.065 36.605 118.315 ;
        RECT 32.945 117.455 33.265 117.810 ;
        RECT 32.195 117.285 33.265 117.455 ;
        RECT 33.465 117.075 33.635 117.885 ;
        RECT 33.805 117.725 35.570 117.895 ;
        RECT 33.805 117.245 34.135 117.725 ;
        RECT 34.305 117.075 34.475 117.545 ;
        RECT 34.645 117.245 34.975 117.725 ;
        RECT 35.145 117.075 35.315 117.545 ;
        RECT 35.795 117.075 36.085 117.800 ;
        RECT 36.295 117.075 36.525 117.895 ;
        RECT 36.775 117.875 37.025 118.475 ;
        RECT 36.695 117.245 37.025 117.875 ;
        RECT 37.195 117.075 37.405 117.895 ;
        RECT 37.635 117.750 37.805 118.550 ;
        RECT 38.090 118.525 38.755 118.695 ;
        RECT 39.015 118.550 39.285 119.455 ;
        RECT 39.455 118.865 39.785 119.625 ;
        RECT 39.965 118.695 40.135 119.455 ;
        RECT 40.400 118.955 40.655 119.455 ;
        RECT 40.825 119.125 41.155 119.625 ;
        RECT 40.400 118.785 41.150 118.955 ;
        RECT 38.090 118.380 38.260 118.525 ;
        RECT 37.975 118.050 38.260 118.380 ;
        RECT 38.090 117.795 38.260 118.050 ;
        RECT 38.495 117.975 38.825 118.345 ;
        RECT 37.635 117.245 37.895 117.750 ;
        RECT 38.090 117.625 38.755 117.795 ;
        RECT 38.075 117.075 38.405 117.455 ;
        RECT 38.585 117.245 38.755 117.625 ;
        RECT 39.015 117.750 39.185 118.550 ;
        RECT 39.470 118.525 40.135 118.695 ;
        RECT 39.470 118.380 39.640 118.525 ;
        RECT 39.355 118.050 39.640 118.380 ;
        RECT 39.470 117.795 39.640 118.050 ;
        RECT 39.875 117.975 40.205 118.345 ;
        RECT 40.400 117.965 40.750 118.615 ;
        RECT 40.920 117.795 41.150 118.785 ;
        RECT 39.015 117.245 39.275 117.750 ;
        RECT 39.470 117.625 40.135 117.795 ;
        RECT 39.455 117.075 39.785 117.455 ;
        RECT 39.965 117.245 40.135 117.625 ;
        RECT 40.400 117.625 41.150 117.795 ;
        RECT 40.400 117.335 40.655 117.625 ;
        RECT 40.825 117.075 41.155 117.455 ;
        RECT 41.325 117.335 41.495 119.455 ;
        RECT 41.665 118.655 41.990 119.440 ;
        RECT 42.160 119.165 42.410 119.625 ;
        RECT 42.580 119.125 42.830 119.455 ;
        RECT 43.045 119.125 43.725 119.455 ;
        RECT 42.580 118.995 42.750 119.125 ;
        RECT 42.355 118.825 42.750 118.995 ;
        RECT 41.725 117.605 42.185 118.655 ;
        RECT 42.355 117.465 42.525 118.825 ;
        RECT 42.920 118.565 43.385 118.955 ;
        RECT 42.695 117.755 43.045 118.375 ;
        RECT 43.215 117.975 43.385 118.565 ;
        RECT 43.555 118.345 43.725 119.125 ;
        RECT 43.895 119.025 44.065 119.365 ;
        RECT 44.300 119.195 44.630 119.625 ;
        RECT 44.800 119.025 44.970 119.365 ;
        RECT 45.265 119.165 45.635 119.625 ;
        RECT 43.895 118.855 44.970 119.025 ;
        RECT 45.805 118.995 45.975 119.455 ;
        RECT 46.210 119.115 47.080 119.455 ;
        RECT 47.250 119.165 47.500 119.625 ;
        RECT 45.415 118.825 45.975 118.995 ;
        RECT 45.415 118.685 45.585 118.825 ;
        RECT 44.085 118.515 45.585 118.685 ;
        RECT 46.280 118.655 46.740 118.945 ;
        RECT 43.555 118.175 45.245 118.345 ;
        RECT 43.215 117.755 43.570 117.975 ;
        RECT 43.740 117.465 43.910 118.175 ;
        RECT 44.115 117.755 44.905 118.005 ;
        RECT 45.075 117.995 45.245 118.175 ;
        RECT 45.415 117.825 45.585 118.515 ;
        RECT 41.855 117.075 42.185 117.435 ;
        RECT 42.355 117.295 42.850 117.465 ;
        RECT 43.055 117.295 43.910 117.465 ;
        RECT 44.785 117.075 45.115 117.535 ;
        RECT 45.325 117.435 45.585 117.825 ;
        RECT 45.775 118.645 46.740 118.655 ;
        RECT 46.910 118.735 47.080 119.115 ;
        RECT 47.670 119.075 47.840 119.365 ;
        RECT 48.020 119.245 48.350 119.625 ;
        RECT 47.670 118.905 48.470 119.075 ;
        RECT 45.775 118.485 46.450 118.645 ;
        RECT 46.910 118.565 48.130 118.735 ;
        RECT 45.775 117.695 45.985 118.485 ;
        RECT 46.910 118.475 47.080 118.565 ;
        RECT 46.155 117.695 46.505 118.315 ;
        RECT 46.675 118.305 47.080 118.475 ;
        RECT 46.675 117.525 46.845 118.305 ;
        RECT 47.015 117.855 47.235 118.135 ;
        RECT 47.415 118.025 47.955 118.395 ;
        RECT 48.300 118.285 48.470 118.905 ;
        RECT 48.645 118.565 48.815 119.625 ;
        RECT 49.025 118.615 49.315 119.455 ;
        RECT 49.485 118.785 49.655 119.625 ;
        RECT 49.865 118.615 50.115 119.455 ;
        RECT 50.325 118.785 50.495 119.625 ;
        RECT 51.285 118.785 51.455 119.625 ;
        RECT 51.665 118.615 51.915 119.455 ;
        RECT 52.125 118.785 52.295 119.625 ;
        RECT 52.465 118.615 52.755 119.455 ;
        RECT 49.025 118.445 50.750 118.615 ;
        RECT 47.015 117.685 47.545 117.855 ;
        RECT 45.325 117.265 45.675 117.435 ;
        RECT 45.895 117.245 46.845 117.525 ;
        RECT 47.015 117.075 47.205 117.515 ;
        RECT 47.375 117.455 47.545 117.685 ;
        RECT 47.715 117.625 47.955 118.025 ;
        RECT 48.125 118.275 48.470 118.285 ;
        RECT 48.125 118.065 50.155 118.275 ;
        RECT 48.125 117.810 48.450 118.065 ;
        RECT 50.340 117.895 50.750 118.445 ;
        RECT 48.125 117.455 48.445 117.810 ;
        RECT 47.375 117.285 48.445 117.455 ;
        RECT 48.645 117.075 48.815 117.885 ;
        RECT 48.985 117.725 50.750 117.895 ;
        RECT 51.030 118.445 52.755 118.615 ;
        RECT 52.965 118.565 53.135 119.625 ;
        RECT 53.430 119.245 53.760 119.625 ;
        RECT 53.940 119.075 54.110 119.365 ;
        RECT 54.280 119.165 54.530 119.625 ;
        RECT 53.310 118.905 54.110 119.075 ;
        RECT 54.700 119.115 55.570 119.455 ;
        RECT 51.030 117.895 51.440 118.445 ;
        RECT 53.310 118.285 53.480 118.905 ;
        RECT 54.700 118.735 54.870 119.115 ;
        RECT 55.805 118.995 55.975 119.455 ;
        RECT 56.145 119.165 56.515 119.625 ;
        RECT 56.810 119.025 56.980 119.365 ;
        RECT 57.150 119.195 57.480 119.625 ;
        RECT 57.715 119.025 57.885 119.365 ;
        RECT 53.650 118.565 54.870 118.735 ;
        RECT 55.040 118.655 55.500 118.945 ;
        RECT 55.805 118.825 56.365 118.995 ;
        RECT 56.810 118.855 57.885 119.025 ;
        RECT 58.055 119.125 58.735 119.455 ;
        RECT 58.950 119.125 59.200 119.455 ;
        RECT 59.370 119.165 59.620 119.625 ;
        RECT 56.195 118.685 56.365 118.825 ;
        RECT 55.040 118.645 56.005 118.655 ;
        RECT 54.700 118.475 54.870 118.565 ;
        RECT 55.330 118.485 56.005 118.645 ;
        RECT 53.310 118.275 53.655 118.285 ;
        RECT 51.625 118.065 53.655 118.275 ;
        RECT 51.030 117.725 52.795 117.895 ;
        RECT 48.985 117.245 49.315 117.725 ;
        RECT 49.485 117.075 49.655 117.545 ;
        RECT 49.825 117.245 50.155 117.725 ;
        RECT 50.325 117.075 50.495 117.545 ;
        RECT 51.285 117.075 51.455 117.545 ;
        RECT 51.625 117.245 51.955 117.725 ;
        RECT 52.125 117.075 52.295 117.545 ;
        RECT 52.465 117.245 52.795 117.725 ;
        RECT 52.965 117.075 53.135 117.885 ;
        RECT 53.330 117.810 53.655 118.065 ;
        RECT 53.335 117.455 53.655 117.810 ;
        RECT 53.825 118.025 54.365 118.395 ;
        RECT 54.700 118.305 55.105 118.475 ;
        RECT 53.825 117.625 54.065 118.025 ;
        RECT 54.545 117.855 54.765 118.135 ;
        RECT 54.235 117.685 54.765 117.855 ;
        RECT 54.235 117.455 54.405 117.685 ;
        RECT 54.935 117.525 55.105 118.305 ;
        RECT 55.275 117.695 55.625 118.315 ;
        RECT 55.795 117.695 56.005 118.485 ;
        RECT 56.195 118.515 57.695 118.685 ;
        RECT 56.195 117.825 56.365 118.515 ;
        RECT 58.055 118.345 58.225 119.125 ;
        RECT 59.030 118.995 59.200 119.125 ;
        RECT 56.535 118.175 58.225 118.345 ;
        RECT 58.395 118.565 58.860 118.955 ;
        RECT 59.030 118.825 59.425 118.995 ;
        RECT 56.535 117.995 56.705 118.175 ;
        RECT 53.335 117.285 54.405 117.455 ;
        RECT 54.575 117.075 54.765 117.515 ;
        RECT 54.935 117.245 55.885 117.525 ;
        RECT 56.195 117.435 56.455 117.825 ;
        RECT 56.875 117.755 57.665 118.005 ;
        RECT 56.105 117.265 56.455 117.435 ;
        RECT 56.665 117.075 56.995 117.535 ;
        RECT 57.870 117.465 58.040 118.175 ;
        RECT 58.395 117.975 58.565 118.565 ;
        RECT 58.210 117.755 58.565 117.975 ;
        RECT 58.735 117.755 59.085 118.375 ;
        RECT 59.255 117.465 59.425 118.825 ;
        RECT 59.790 118.655 60.115 119.440 ;
        RECT 59.595 117.605 60.055 118.655 ;
        RECT 57.870 117.295 58.725 117.465 ;
        RECT 58.930 117.295 59.425 117.465 ;
        RECT 59.595 117.075 59.925 117.435 ;
        RECT 60.285 117.335 60.455 119.455 ;
        RECT 60.625 119.125 60.955 119.625 ;
        RECT 61.125 118.955 61.380 119.455 ;
        RECT 60.630 118.785 61.380 118.955 ;
        RECT 60.630 117.795 60.860 118.785 ;
        RECT 61.030 117.965 61.380 118.615 ;
        RECT 61.555 118.460 61.845 119.625 ;
        RECT 62.325 118.785 62.495 119.625 ;
        RECT 62.705 118.615 62.955 119.455 ;
        RECT 63.165 118.785 63.335 119.625 ;
        RECT 63.505 118.615 63.795 119.455 ;
        RECT 62.070 118.445 63.795 118.615 ;
        RECT 64.005 118.565 64.175 119.625 ;
        RECT 64.470 119.245 64.800 119.625 ;
        RECT 64.980 119.075 65.150 119.365 ;
        RECT 65.320 119.165 65.570 119.625 ;
        RECT 64.350 118.905 65.150 119.075 ;
        RECT 65.740 119.115 66.610 119.455 ;
        RECT 62.070 117.895 62.480 118.445 ;
        RECT 64.350 118.285 64.520 118.905 ;
        RECT 65.740 118.735 65.910 119.115 ;
        RECT 66.845 118.995 67.015 119.455 ;
        RECT 67.185 119.165 67.555 119.625 ;
        RECT 67.850 119.025 68.020 119.365 ;
        RECT 68.190 119.195 68.520 119.625 ;
        RECT 68.755 119.025 68.925 119.365 ;
        RECT 64.690 118.565 65.910 118.735 ;
        RECT 66.080 118.655 66.540 118.945 ;
        RECT 66.845 118.825 67.405 118.995 ;
        RECT 67.850 118.855 68.925 119.025 ;
        RECT 69.095 119.125 69.775 119.455 ;
        RECT 69.990 119.125 70.240 119.455 ;
        RECT 70.410 119.165 70.660 119.625 ;
        RECT 67.235 118.685 67.405 118.825 ;
        RECT 66.080 118.645 67.045 118.655 ;
        RECT 65.740 118.475 65.910 118.565 ;
        RECT 66.370 118.485 67.045 118.645 ;
        RECT 64.350 118.275 64.695 118.285 ;
        RECT 62.665 118.065 64.695 118.275 ;
        RECT 60.630 117.625 61.380 117.795 ;
        RECT 60.625 117.075 60.955 117.455 ;
        RECT 61.125 117.335 61.380 117.625 ;
        RECT 61.555 117.075 61.845 117.800 ;
        RECT 62.070 117.725 63.835 117.895 ;
        RECT 62.325 117.075 62.495 117.545 ;
        RECT 62.665 117.245 62.995 117.725 ;
        RECT 63.165 117.075 63.335 117.545 ;
        RECT 63.505 117.245 63.835 117.725 ;
        RECT 64.005 117.075 64.175 117.885 ;
        RECT 64.370 117.810 64.695 118.065 ;
        RECT 64.375 117.455 64.695 117.810 ;
        RECT 64.865 118.025 65.405 118.395 ;
        RECT 65.740 118.305 66.145 118.475 ;
        RECT 64.865 117.625 65.105 118.025 ;
        RECT 65.585 117.855 65.805 118.135 ;
        RECT 65.275 117.685 65.805 117.855 ;
        RECT 65.275 117.455 65.445 117.685 ;
        RECT 65.975 117.525 66.145 118.305 ;
        RECT 66.315 117.695 66.665 118.315 ;
        RECT 66.835 117.695 67.045 118.485 ;
        RECT 67.235 118.515 68.735 118.685 ;
        RECT 67.235 117.825 67.405 118.515 ;
        RECT 69.095 118.345 69.265 119.125 ;
        RECT 70.070 118.995 70.240 119.125 ;
        RECT 67.575 118.175 69.265 118.345 ;
        RECT 69.435 118.565 69.900 118.955 ;
        RECT 70.070 118.825 70.465 118.995 ;
        RECT 67.575 117.995 67.745 118.175 ;
        RECT 64.375 117.285 65.445 117.455 ;
        RECT 65.615 117.075 65.805 117.515 ;
        RECT 65.975 117.245 66.925 117.525 ;
        RECT 67.235 117.435 67.495 117.825 ;
        RECT 67.915 117.755 68.705 118.005 ;
        RECT 67.145 117.265 67.495 117.435 ;
        RECT 67.705 117.075 68.035 117.535 ;
        RECT 68.910 117.465 69.080 118.175 ;
        RECT 69.435 117.975 69.605 118.565 ;
        RECT 69.250 117.755 69.605 117.975 ;
        RECT 69.775 117.755 70.125 118.375 ;
        RECT 70.295 117.465 70.465 118.825 ;
        RECT 70.830 118.655 71.155 119.440 ;
        RECT 70.635 117.605 71.095 118.655 ;
        RECT 68.910 117.295 69.765 117.465 ;
        RECT 69.970 117.295 70.465 117.465 ;
        RECT 70.635 117.075 70.965 117.435 ;
        RECT 71.325 117.335 71.495 119.455 ;
        RECT 71.665 119.125 71.995 119.625 ;
        RECT 72.165 118.955 72.420 119.455 ;
        RECT 71.670 118.785 72.420 118.955 ;
        RECT 72.905 118.785 73.075 119.625 ;
        RECT 71.670 117.795 71.900 118.785 ;
        RECT 73.285 118.615 73.535 119.455 ;
        RECT 73.745 118.785 73.915 119.625 ;
        RECT 74.085 118.615 74.375 119.455 ;
        RECT 72.070 117.965 72.420 118.615 ;
        RECT 72.650 118.445 74.375 118.615 ;
        RECT 74.585 118.565 74.755 119.625 ;
        RECT 75.050 119.245 75.380 119.625 ;
        RECT 75.560 119.075 75.730 119.365 ;
        RECT 75.900 119.165 76.150 119.625 ;
        RECT 74.930 118.905 75.730 119.075 ;
        RECT 76.320 119.115 77.190 119.455 ;
        RECT 72.650 117.895 73.060 118.445 ;
        RECT 74.930 118.285 75.100 118.905 ;
        RECT 76.320 118.735 76.490 119.115 ;
        RECT 77.425 118.995 77.595 119.455 ;
        RECT 77.765 119.165 78.135 119.625 ;
        RECT 78.430 119.025 78.600 119.365 ;
        RECT 78.770 119.195 79.100 119.625 ;
        RECT 79.335 119.025 79.505 119.365 ;
        RECT 75.270 118.565 76.490 118.735 ;
        RECT 76.660 118.655 77.120 118.945 ;
        RECT 77.425 118.825 77.985 118.995 ;
        RECT 78.430 118.855 79.505 119.025 ;
        RECT 79.675 119.125 80.355 119.455 ;
        RECT 80.570 119.125 80.820 119.455 ;
        RECT 80.990 119.165 81.240 119.625 ;
        RECT 77.815 118.685 77.985 118.825 ;
        RECT 76.660 118.645 77.625 118.655 ;
        RECT 76.320 118.475 76.490 118.565 ;
        RECT 76.950 118.485 77.625 118.645 ;
        RECT 74.930 118.275 75.275 118.285 ;
        RECT 73.245 118.065 75.275 118.275 ;
        RECT 71.670 117.625 72.420 117.795 ;
        RECT 72.650 117.725 74.415 117.895 ;
        RECT 71.665 117.075 71.995 117.455 ;
        RECT 72.165 117.335 72.420 117.625 ;
        RECT 72.905 117.075 73.075 117.545 ;
        RECT 73.245 117.245 73.575 117.725 ;
        RECT 73.745 117.075 73.915 117.545 ;
        RECT 74.085 117.245 74.415 117.725 ;
        RECT 74.585 117.075 74.755 117.885 ;
        RECT 74.950 117.810 75.275 118.065 ;
        RECT 74.955 117.455 75.275 117.810 ;
        RECT 75.445 118.025 75.985 118.395 ;
        RECT 76.320 118.305 76.725 118.475 ;
        RECT 75.445 117.625 75.685 118.025 ;
        RECT 76.165 117.855 76.385 118.135 ;
        RECT 75.855 117.685 76.385 117.855 ;
        RECT 75.855 117.455 76.025 117.685 ;
        RECT 76.555 117.525 76.725 118.305 ;
        RECT 76.895 117.695 77.245 118.315 ;
        RECT 77.415 117.695 77.625 118.485 ;
        RECT 77.815 118.515 79.315 118.685 ;
        RECT 77.815 117.825 77.985 118.515 ;
        RECT 79.675 118.345 79.845 119.125 ;
        RECT 80.650 118.995 80.820 119.125 ;
        RECT 78.155 118.175 79.845 118.345 ;
        RECT 80.015 118.565 80.480 118.955 ;
        RECT 80.650 118.825 81.045 118.995 ;
        RECT 78.155 117.995 78.325 118.175 ;
        RECT 74.955 117.285 76.025 117.455 ;
        RECT 76.195 117.075 76.385 117.515 ;
        RECT 76.555 117.245 77.505 117.525 ;
        RECT 77.815 117.435 78.075 117.825 ;
        RECT 78.495 117.755 79.285 118.005 ;
        RECT 77.725 117.265 78.075 117.435 ;
        RECT 78.285 117.075 78.615 117.535 ;
        RECT 79.490 117.465 79.660 118.175 ;
        RECT 80.015 117.975 80.185 118.565 ;
        RECT 79.830 117.755 80.185 117.975 ;
        RECT 80.355 117.755 80.705 118.375 ;
        RECT 80.875 117.465 81.045 118.825 ;
        RECT 81.410 118.655 81.735 119.440 ;
        RECT 81.215 117.605 81.675 118.655 ;
        RECT 79.490 117.295 80.345 117.465 ;
        RECT 80.550 117.295 81.045 117.465 ;
        RECT 81.215 117.075 81.545 117.435 ;
        RECT 81.905 117.335 82.075 119.455 ;
        RECT 82.245 119.125 82.575 119.625 ;
        RECT 82.745 118.955 83.000 119.455 ;
        RECT 82.250 118.785 83.000 118.955 ;
        RECT 82.250 117.795 82.480 118.785 ;
        RECT 82.650 117.965 83.000 118.615 ;
        RECT 83.235 118.485 83.445 119.625 ;
        RECT 83.615 118.475 83.945 119.455 ;
        RECT 84.115 118.485 84.345 119.625 ;
        RECT 84.595 118.485 84.825 119.625 ;
        RECT 84.995 118.475 85.325 119.455 ;
        RECT 85.495 118.485 85.705 119.625 ;
        RECT 85.975 118.485 86.205 119.625 ;
        RECT 86.375 118.475 86.705 119.455 ;
        RECT 86.875 118.485 87.085 119.625 ;
        RECT 82.250 117.625 83.000 117.795 ;
        RECT 82.245 117.075 82.575 117.455 ;
        RECT 82.745 117.335 83.000 117.625 ;
        RECT 83.235 117.075 83.445 117.895 ;
        RECT 83.615 117.875 83.865 118.475 ;
        RECT 84.035 118.065 84.365 118.315 ;
        RECT 84.575 118.065 84.905 118.315 ;
        RECT 83.615 117.245 83.945 117.875 ;
        RECT 84.115 117.075 84.345 117.895 ;
        RECT 84.595 117.075 84.825 117.895 ;
        RECT 85.075 117.875 85.325 118.475 ;
        RECT 85.955 118.065 86.285 118.315 ;
        RECT 84.995 117.245 85.325 117.875 ;
        RECT 85.495 117.075 85.705 117.895 ;
        RECT 85.975 117.075 86.205 117.895 ;
        RECT 86.455 117.875 86.705 118.475 ;
        RECT 87.315 118.460 87.605 119.625 ;
        RECT 88.085 118.785 88.255 119.625 ;
        RECT 88.465 118.615 88.715 119.455 ;
        RECT 88.925 118.785 89.095 119.625 ;
        RECT 89.265 118.615 89.555 119.455 ;
        RECT 87.830 118.445 89.555 118.615 ;
        RECT 89.765 118.565 89.935 119.625 ;
        RECT 90.230 119.245 90.560 119.625 ;
        RECT 90.740 119.075 90.910 119.365 ;
        RECT 91.080 119.165 91.330 119.625 ;
        RECT 90.110 118.905 90.910 119.075 ;
        RECT 91.500 119.115 92.370 119.455 ;
        RECT 87.830 117.895 88.240 118.445 ;
        RECT 90.110 118.285 90.280 118.905 ;
        RECT 91.500 118.735 91.670 119.115 ;
        RECT 92.605 118.995 92.775 119.455 ;
        RECT 92.945 119.165 93.315 119.625 ;
        RECT 93.610 119.025 93.780 119.365 ;
        RECT 93.950 119.195 94.280 119.625 ;
        RECT 94.515 119.025 94.685 119.365 ;
        RECT 90.450 118.565 91.670 118.735 ;
        RECT 91.840 118.655 92.300 118.945 ;
        RECT 92.605 118.825 93.165 118.995 ;
        RECT 93.610 118.855 94.685 119.025 ;
        RECT 94.855 119.125 95.535 119.455 ;
        RECT 95.750 119.125 96.000 119.455 ;
        RECT 96.170 119.165 96.420 119.625 ;
        RECT 92.995 118.685 93.165 118.825 ;
        RECT 91.840 118.645 92.805 118.655 ;
        RECT 91.500 118.475 91.670 118.565 ;
        RECT 92.130 118.485 92.805 118.645 ;
        RECT 90.110 118.275 90.455 118.285 ;
        RECT 88.425 118.065 90.455 118.275 ;
        RECT 86.375 117.245 86.705 117.875 ;
        RECT 86.875 117.075 87.085 117.895 ;
        RECT 87.315 117.075 87.605 117.800 ;
        RECT 87.830 117.725 89.595 117.895 ;
        RECT 88.085 117.075 88.255 117.545 ;
        RECT 88.425 117.245 88.755 117.725 ;
        RECT 88.925 117.075 89.095 117.545 ;
        RECT 89.265 117.245 89.595 117.725 ;
        RECT 89.765 117.075 89.935 117.885 ;
        RECT 90.130 117.810 90.455 118.065 ;
        RECT 90.135 117.455 90.455 117.810 ;
        RECT 90.625 118.025 91.165 118.395 ;
        RECT 91.500 118.305 91.905 118.475 ;
        RECT 90.625 117.625 90.865 118.025 ;
        RECT 91.345 117.855 91.565 118.135 ;
        RECT 91.035 117.685 91.565 117.855 ;
        RECT 91.035 117.455 91.205 117.685 ;
        RECT 91.735 117.525 91.905 118.305 ;
        RECT 92.075 117.695 92.425 118.315 ;
        RECT 92.595 117.695 92.805 118.485 ;
        RECT 92.995 118.515 94.495 118.685 ;
        RECT 92.995 117.825 93.165 118.515 ;
        RECT 94.855 118.345 95.025 119.125 ;
        RECT 95.830 118.995 96.000 119.125 ;
        RECT 93.335 118.175 95.025 118.345 ;
        RECT 95.195 118.565 95.660 118.955 ;
        RECT 95.830 118.825 96.225 118.995 ;
        RECT 93.335 117.995 93.505 118.175 ;
        RECT 90.135 117.285 91.205 117.455 ;
        RECT 91.375 117.075 91.565 117.515 ;
        RECT 91.735 117.245 92.685 117.525 ;
        RECT 92.995 117.435 93.255 117.825 ;
        RECT 93.675 117.755 94.465 118.005 ;
        RECT 92.905 117.265 93.255 117.435 ;
        RECT 93.465 117.075 93.795 117.535 ;
        RECT 94.670 117.465 94.840 118.175 ;
        RECT 95.195 117.975 95.365 118.565 ;
        RECT 95.010 117.755 95.365 117.975 ;
        RECT 95.535 117.755 95.885 118.375 ;
        RECT 96.055 117.465 96.225 118.825 ;
        RECT 96.590 118.655 96.915 119.440 ;
        RECT 96.395 117.605 96.855 118.655 ;
        RECT 94.670 117.295 95.525 117.465 ;
        RECT 95.730 117.295 96.225 117.465 ;
        RECT 96.395 117.075 96.725 117.435 ;
        RECT 97.085 117.335 97.255 119.455 ;
        RECT 97.425 119.125 97.755 119.625 ;
        RECT 97.925 118.955 98.180 119.455 ;
        RECT 97.430 118.785 98.180 118.955 ;
        RECT 98.360 118.955 98.615 119.455 ;
        RECT 98.785 119.125 99.115 119.625 ;
        RECT 98.360 118.785 99.110 118.955 ;
        RECT 97.430 117.795 97.660 118.785 ;
        RECT 97.830 117.965 98.180 118.615 ;
        RECT 98.360 117.965 98.710 118.615 ;
        RECT 98.880 117.795 99.110 118.785 ;
        RECT 97.430 117.625 98.180 117.795 ;
        RECT 97.425 117.075 97.755 117.455 ;
        RECT 97.925 117.335 98.180 117.625 ;
        RECT 98.360 117.625 99.110 117.795 ;
        RECT 98.360 117.335 98.615 117.625 ;
        RECT 98.785 117.075 99.115 117.455 ;
        RECT 99.285 117.335 99.455 119.455 ;
        RECT 99.625 118.655 99.950 119.440 ;
        RECT 100.120 119.165 100.370 119.625 ;
        RECT 100.540 119.125 100.790 119.455 ;
        RECT 101.005 119.125 101.685 119.455 ;
        RECT 100.540 118.995 100.710 119.125 ;
        RECT 100.315 118.825 100.710 118.995 ;
        RECT 99.685 117.605 100.145 118.655 ;
        RECT 100.315 117.465 100.485 118.825 ;
        RECT 100.880 118.565 101.345 118.955 ;
        RECT 100.655 117.755 101.005 118.375 ;
        RECT 101.175 117.975 101.345 118.565 ;
        RECT 101.515 118.345 101.685 119.125 ;
        RECT 101.855 119.025 102.025 119.365 ;
        RECT 102.260 119.195 102.590 119.625 ;
        RECT 102.760 119.025 102.930 119.365 ;
        RECT 103.225 119.165 103.595 119.625 ;
        RECT 101.855 118.855 102.930 119.025 ;
        RECT 103.765 118.995 103.935 119.455 ;
        RECT 104.170 119.115 105.040 119.455 ;
        RECT 105.210 119.165 105.460 119.625 ;
        RECT 103.375 118.825 103.935 118.995 ;
        RECT 103.375 118.685 103.545 118.825 ;
        RECT 102.045 118.515 103.545 118.685 ;
        RECT 104.240 118.655 104.700 118.945 ;
        RECT 101.515 118.175 103.205 118.345 ;
        RECT 101.175 117.755 101.530 117.975 ;
        RECT 101.700 117.465 101.870 118.175 ;
        RECT 102.075 117.755 102.865 118.005 ;
        RECT 103.035 117.995 103.205 118.175 ;
        RECT 103.375 117.825 103.545 118.515 ;
        RECT 99.815 117.075 100.145 117.435 ;
        RECT 100.315 117.295 100.810 117.465 ;
        RECT 101.015 117.295 101.870 117.465 ;
        RECT 102.745 117.075 103.075 117.535 ;
        RECT 103.285 117.435 103.545 117.825 ;
        RECT 103.735 118.645 104.700 118.655 ;
        RECT 104.870 118.735 105.040 119.115 ;
        RECT 105.630 119.075 105.800 119.365 ;
        RECT 105.980 119.245 106.310 119.625 ;
        RECT 105.630 118.905 106.430 119.075 ;
        RECT 103.735 118.485 104.410 118.645 ;
        RECT 104.870 118.565 106.090 118.735 ;
        RECT 103.735 117.695 103.945 118.485 ;
        RECT 104.870 118.475 105.040 118.565 ;
        RECT 104.115 117.695 104.465 118.315 ;
        RECT 104.635 118.305 105.040 118.475 ;
        RECT 104.635 117.525 104.805 118.305 ;
        RECT 104.975 117.855 105.195 118.135 ;
        RECT 105.375 118.025 105.915 118.395 ;
        RECT 106.260 118.285 106.430 118.905 ;
        RECT 106.605 118.565 106.775 119.625 ;
        RECT 106.985 118.615 107.275 119.455 ;
        RECT 107.445 118.785 107.615 119.625 ;
        RECT 107.825 118.615 108.075 119.455 ;
        RECT 108.285 118.785 108.455 119.625 ;
        RECT 106.985 118.445 108.710 118.615 ;
        RECT 108.995 118.485 109.205 119.625 ;
        RECT 104.975 117.685 105.505 117.855 ;
        RECT 103.285 117.265 103.635 117.435 ;
        RECT 103.855 117.245 104.805 117.525 ;
        RECT 104.975 117.075 105.165 117.515 ;
        RECT 105.335 117.455 105.505 117.685 ;
        RECT 105.675 117.625 105.915 118.025 ;
        RECT 106.085 118.275 106.430 118.285 ;
        RECT 106.085 118.065 108.115 118.275 ;
        RECT 106.085 117.810 106.410 118.065 ;
        RECT 108.300 117.895 108.710 118.445 ;
        RECT 109.375 118.475 109.705 119.455 ;
        RECT 109.875 118.485 110.105 119.625 ;
        RECT 110.355 118.485 110.585 119.625 ;
        RECT 110.755 118.475 111.085 119.455 ;
        RECT 111.255 118.485 111.465 119.625 ;
        RECT 112.155 118.535 113.365 119.625 ;
        RECT 106.085 117.455 106.405 117.810 ;
        RECT 105.335 117.285 106.405 117.455 ;
        RECT 106.605 117.075 106.775 117.885 ;
        RECT 106.945 117.725 108.710 117.895 ;
        RECT 106.945 117.245 107.275 117.725 ;
        RECT 107.445 117.075 107.615 117.545 ;
        RECT 107.785 117.245 108.115 117.725 ;
        RECT 108.285 117.075 108.455 117.545 ;
        RECT 108.995 117.075 109.205 117.895 ;
        RECT 109.375 117.875 109.625 118.475 ;
        RECT 109.795 118.065 110.125 118.315 ;
        RECT 110.335 118.065 110.665 118.315 ;
        RECT 109.375 117.245 109.705 117.875 ;
        RECT 109.875 117.075 110.105 117.895 ;
        RECT 110.355 117.075 110.585 117.895 ;
        RECT 110.835 117.875 111.085 118.475 ;
        RECT 112.155 117.995 112.675 118.535 ;
        RECT 110.755 117.245 111.085 117.875 ;
        RECT 111.255 117.075 111.465 117.895 ;
        RECT 112.845 117.825 113.365 118.365 ;
        RECT 112.155 117.075 113.365 117.825 ;
        RECT 22.830 116.905 113.450 117.075 ;
        RECT 22.915 116.155 24.125 116.905 ;
        RECT 24.605 116.435 24.775 116.905 ;
        RECT 24.945 116.255 25.275 116.735 ;
        RECT 25.445 116.435 25.615 116.905 ;
        RECT 25.785 116.255 26.115 116.735 ;
        RECT 22.915 115.615 23.435 116.155 ;
        RECT 24.350 116.085 26.115 116.255 ;
        RECT 26.285 116.095 26.455 116.905 ;
        RECT 26.655 116.525 27.725 116.695 ;
        RECT 26.655 116.170 26.975 116.525 ;
        RECT 23.605 115.445 24.125 115.985 ;
        RECT 22.915 114.355 24.125 115.445 ;
        RECT 24.350 115.535 24.760 116.085 ;
        RECT 26.650 115.915 26.975 116.170 ;
        RECT 24.945 115.705 26.975 115.915 ;
        RECT 26.630 115.695 26.975 115.705 ;
        RECT 27.145 115.955 27.385 116.355 ;
        RECT 27.555 116.295 27.725 116.525 ;
        RECT 27.895 116.465 28.085 116.905 ;
        RECT 28.255 116.455 29.205 116.735 ;
        RECT 29.425 116.545 29.775 116.715 ;
        RECT 27.555 116.125 28.085 116.295 ;
        RECT 24.350 115.365 26.075 115.535 ;
        RECT 24.605 114.355 24.775 115.195 ;
        RECT 24.985 114.525 25.235 115.365 ;
        RECT 25.445 114.355 25.615 115.195 ;
        RECT 25.785 114.525 26.075 115.365 ;
        RECT 26.285 114.355 26.455 115.415 ;
        RECT 26.630 115.075 26.800 115.695 ;
        RECT 27.145 115.585 27.685 115.955 ;
        RECT 27.865 115.845 28.085 116.125 ;
        RECT 28.255 115.675 28.425 116.455 ;
        RECT 28.020 115.505 28.425 115.675 ;
        RECT 28.595 115.665 28.945 116.285 ;
        RECT 28.020 115.415 28.190 115.505 ;
        RECT 29.115 115.495 29.325 116.285 ;
        RECT 26.970 115.245 28.190 115.415 ;
        RECT 28.650 115.335 29.325 115.495 ;
        RECT 26.630 114.905 27.430 115.075 ;
        RECT 26.750 114.355 27.080 114.735 ;
        RECT 27.260 114.615 27.430 114.905 ;
        RECT 28.020 114.865 28.190 115.245 ;
        RECT 28.360 115.325 29.325 115.335 ;
        RECT 29.515 116.155 29.775 116.545 ;
        RECT 29.985 116.445 30.315 116.905 ;
        RECT 31.190 116.515 32.045 116.685 ;
        RECT 32.250 116.515 32.745 116.685 ;
        RECT 32.915 116.545 33.245 116.905 ;
        RECT 29.515 115.465 29.685 116.155 ;
        RECT 29.855 115.805 30.025 115.985 ;
        RECT 30.195 115.975 30.985 116.225 ;
        RECT 31.190 115.805 31.360 116.515 ;
        RECT 31.530 116.005 31.885 116.225 ;
        RECT 29.855 115.635 31.545 115.805 ;
        RECT 28.360 115.035 28.820 115.325 ;
        RECT 29.515 115.295 31.015 115.465 ;
        RECT 29.515 115.155 29.685 115.295 ;
        RECT 29.125 114.985 29.685 115.155 ;
        RECT 27.600 114.355 27.850 114.815 ;
        RECT 28.020 114.525 28.890 114.865 ;
        RECT 29.125 114.525 29.295 114.985 ;
        RECT 30.130 114.955 31.205 115.125 ;
        RECT 29.465 114.355 29.835 114.815 ;
        RECT 30.130 114.615 30.300 114.955 ;
        RECT 30.470 114.355 30.800 114.785 ;
        RECT 31.035 114.615 31.205 114.955 ;
        RECT 31.375 114.855 31.545 115.635 ;
        RECT 31.715 115.415 31.885 116.005 ;
        RECT 32.055 115.605 32.405 116.225 ;
        RECT 31.715 115.025 32.180 115.415 ;
        RECT 32.575 115.155 32.745 116.515 ;
        RECT 32.915 115.325 33.375 116.375 ;
        RECT 32.350 114.985 32.745 115.155 ;
        RECT 32.350 114.855 32.520 114.985 ;
        RECT 31.375 114.525 32.055 114.855 ;
        RECT 32.270 114.525 32.520 114.855 ;
        RECT 32.690 114.355 32.940 114.815 ;
        RECT 33.110 114.540 33.435 115.325 ;
        RECT 33.605 114.525 33.775 116.645 ;
        RECT 33.945 116.525 34.275 116.905 ;
        RECT 34.445 116.355 34.700 116.645 ;
        RECT 33.950 116.185 34.700 116.355 ;
        RECT 33.950 115.195 34.180 116.185 ;
        RECT 35.795 116.180 36.085 116.905 ;
        RECT 36.315 116.085 36.525 116.905 ;
        RECT 36.695 116.105 37.025 116.735 ;
        RECT 34.350 115.365 34.700 116.015 ;
        RECT 33.950 115.025 34.700 115.195 ;
        RECT 33.945 114.355 34.275 114.855 ;
        RECT 34.445 114.525 34.700 115.025 ;
        RECT 35.795 114.355 36.085 115.520 ;
        RECT 36.695 115.505 36.945 116.105 ;
        RECT 37.195 116.085 37.425 116.905 ;
        RECT 37.635 116.230 37.895 116.735 ;
        RECT 38.075 116.525 38.405 116.905 ;
        RECT 38.585 116.355 38.755 116.735 ;
        RECT 37.115 115.665 37.445 115.915 ;
        RECT 36.315 114.355 36.525 115.495 ;
        RECT 36.695 114.525 37.025 115.505 ;
        RECT 37.195 114.355 37.425 115.495 ;
        RECT 37.635 115.430 37.805 116.230 ;
        RECT 38.090 116.185 38.755 116.355 ;
        RECT 38.090 115.930 38.260 116.185 ;
        RECT 39.075 116.085 39.285 116.905 ;
        RECT 39.455 116.105 39.785 116.735 ;
        RECT 37.975 115.600 38.260 115.930 ;
        RECT 38.495 115.635 38.825 116.005 ;
        RECT 38.090 115.455 38.260 115.600 ;
        RECT 39.455 115.505 39.705 116.105 ;
        RECT 39.955 116.085 40.185 116.905 ;
        RECT 40.455 116.085 40.665 116.905 ;
        RECT 40.835 116.105 41.165 116.735 ;
        RECT 39.875 115.665 40.205 115.915 ;
        RECT 40.835 115.505 41.085 116.105 ;
        RECT 41.335 116.085 41.565 116.905 ;
        RECT 41.775 116.135 44.365 116.905 ;
        RECT 41.255 115.665 41.585 115.915 ;
        RECT 37.635 114.525 37.905 115.430 ;
        RECT 38.090 115.285 38.755 115.455 ;
        RECT 38.075 114.355 38.405 115.115 ;
        RECT 38.585 114.525 38.755 115.285 ;
        RECT 39.075 114.355 39.285 115.495 ;
        RECT 39.455 114.525 39.785 115.505 ;
        RECT 39.955 114.355 40.185 115.495 ;
        RECT 40.455 114.355 40.665 115.495 ;
        RECT 40.835 114.525 41.165 115.505 ;
        RECT 41.335 114.355 41.565 115.495 ;
        RECT 41.775 115.445 42.985 115.965 ;
        RECT 43.155 115.615 44.365 116.135 ;
        RECT 44.575 116.085 44.805 116.905 ;
        RECT 44.975 116.105 45.305 116.735 ;
        RECT 44.555 115.665 44.885 115.915 ;
        RECT 45.055 115.505 45.305 116.105 ;
        RECT 45.475 116.085 45.685 116.905 ;
        RECT 46.005 116.355 46.175 116.735 ;
        RECT 46.355 116.525 46.685 116.905 ;
        RECT 46.005 116.185 46.670 116.355 ;
        RECT 46.865 116.230 47.125 116.735 ;
        RECT 45.935 115.635 46.265 116.005 ;
        RECT 46.500 115.930 46.670 116.185 ;
        RECT 41.775 114.355 44.365 115.445 ;
        RECT 44.575 114.355 44.805 115.495 ;
        RECT 44.975 114.525 45.305 115.505 ;
        RECT 46.500 115.600 46.785 115.930 ;
        RECT 45.475 114.355 45.685 115.495 ;
        RECT 46.500 115.455 46.670 115.600 ;
        RECT 46.005 115.285 46.670 115.455 ;
        RECT 46.955 115.430 47.125 116.230 ;
        RECT 47.295 116.155 48.505 116.905 ;
        RECT 48.675 116.180 48.965 116.905 ;
        RECT 46.005 114.525 46.175 115.285 ;
        RECT 46.355 114.355 46.685 115.115 ;
        RECT 46.855 114.525 47.125 115.430 ;
        RECT 47.295 115.445 47.815 115.985 ;
        RECT 47.985 115.615 48.505 116.155 ;
        RECT 49.135 116.135 51.725 116.905 ;
        RECT 51.900 116.360 57.245 116.905 ;
        RECT 47.295 114.355 48.505 115.445 ;
        RECT 48.675 114.355 48.965 115.520 ;
        RECT 49.135 115.445 50.345 115.965 ;
        RECT 50.515 115.615 51.725 116.135 ;
        RECT 49.135 114.355 51.725 115.445 ;
        RECT 53.490 114.790 53.840 116.040 ;
        RECT 55.320 115.530 55.660 116.360 ;
        RECT 57.475 116.085 57.685 116.905 ;
        RECT 57.855 116.105 58.185 116.735 ;
        RECT 57.855 115.505 58.105 116.105 ;
        RECT 58.355 116.085 58.585 116.905 ;
        RECT 58.795 116.135 61.385 116.905 ;
        RECT 61.555 116.180 61.845 116.905 ;
        RECT 58.275 115.665 58.605 115.915 ;
        RECT 51.900 114.355 57.245 114.790 ;
        RECT 57.475 114.355 57.685 115.495 ;
        RECT 57.855 114.525 58.185 115.505 ;
        RECT 58.355 114.355 58.585 115.495 ;
        RECT 58.795 115.445 60.005 115.965 ;
        RECT 60.175 115.615 61.385 116.135 ;
        RECT 62.055 116.085 62.285 116.905 ;
        RECT 62.455 116.105 62.785 116.735 ;
        RECT 62.035 115.665 62.365 115.915 ;
        RECT 58.795 114.355 61.385 115.445 ;
        RECT 61.555 114.355 61.845 115.520 ;
        RECT 62.535 115.505 62.785 116.105 ;
        RECT 62.955 116.085 63.165 116.905 ;
        RECT 63.895 116.085 64.125 116.905 ;
        RECT 64.295 116.105 64.625 116.735 ;
        RECT 63.875 115.665 64.205 115.915 ;
        RECT 64.375 115.505 64.625 116.105 ;
        RECT 64.795 116.085 65.005 116.905 ;
        RECT 65.695 116.135 67.365 116.905 ;
        RECT 67.540 116.360 72.885 116.905 ;
        RECT 62.055 114.355 62.285 115.495 ;
        RECT 62.455 114.525 62.785 115.505 ;
        RECT 62.955 114.355 63.165 115.495 ;
        RECT 63.895 114.355 64.125 115.495 ;
        RECT 64.295 114.525 64.625 115.505 ;
        RECT 64.795 114.355 65.005 115.495 ;
        RECT 65.695 115.445 66.445 115.965 ;
        RECT 66.615 115.615 67.365 116.135 ;
        RECT 65.695 114.355 67.365 115.445 ;
        RECT 69.130 114.790 69.480 116.040 ;
        RECT 70.960 115.530 71.300 116.360 ;
        RECT 73.115 116.085 73.325 116.905 ;
        RECT 73.495 116.105 73.825 116.735 ;
        RECT 73.495 115.505 73.745 116.105 ;
        RECT 73.995 116.085 74.225 116.905 ;
        RECT 74.435 116.180 74.725 116.905 ;
        RECT 75.395 116.085 75.625 116.905 ;
        RECT 75.795 116.105 76.125 116.735 ;
        RECT 73.915 115.665 74.245 115.915 ;
        RECT 75.375 115.665 75.705 115.915 ;
        RECT 67.540 114.355 72.885 114.790 ;
        RECT 73.115 114.355 73.325 115.495 ;
        RECT 73.495 114.525 73.825 115.505 ;
        RECT 73.995 114.355 74.225 115.495 ;
        RECT 74.435 114.355 74.725 115.520 ;
        RECT 75.875 115.505 76.125 116.105 ;
        RECT 76.295 116.085 76.505 116.905 ;
        RECT 76.740 116.355 76.995 116.645 ;
        RECT 77.165 116.525 77.495 116.905 ;
        RECT 76.740 116.185 77.490 116.355 ;
        RECT 75.395 114.355 75.625 115.495 ;
        RECT 75.795 114.525 76.125 115.505 ;
        RECT 76.295 114.355 76.505 115.495 ;
        RECT 76.740 115.365 77.090 116.015 ;
        RECT 77.260 115.195 77.490 116.185 ;
        RECT 76.740 115.025 77.490 115.195 ;
        RECT 76.740 114.525 76.995 115.025 ;
        RECT 77.165 114.355 77.495 114.855 ;
        RECT 77.665 114.525 77.835 116.645 ;
        RECT 78.195 116.545 78.525 116.905 ;
        RECT 78.695 116.515 79.190 116.685 ;
        RECT 79.395 116.515 80.250 116.685 ;
        RECT 78.065 115.325 78.525 116.375 ;
        RECT 78.005 114.540 78.330 115.325 ;
        RECT 78.695 115.155 78.865 116.515 ;
        RECT 79.035 115.605 79.385 116.225 ;
        RECT 79.555 116.005 79.910 116.225 ;
        RECT 79.555 115.415 79.725 116.005 ;
        RECT 80.080 115.805 80.250 116.515 ;
        RECT 81.125 116.445 81.455 116.905 ;
        RECT 81.665 116.545 82.015 116.715 ;
        RECT 80.455 115.975 81.245 116.225 ;
        RECT 81.665 116.155 81.925 116.545 ;
        RECT 82.235 116.455 83.185 116.735 ;
        RECT 83.355 116.465 83.545 116.905 ;
        RECT 83.715 116.525 84.785 116.695 ;
        RECT 81.415 115.805 81.585 115.985 ;
        RECT 78.695 114.985 79.090 115.155 ;
        RECT 79.260 115.025 79.725 115.415 ;
        RECT 79.895 115.635 81.585 115.805 ;
        RECT 78.920 114.855 79.090 114.985 ;
        RECT 79.895 114.855 80.065 115.635 ;
        RECT 81.755 115.465 81.925 116.155 ;
        RECT 80.425 115.295 81.925 115.465 ;
        RECT 82.115 115.495 82.325 116.285 ;
        RECT 82.495 115.665 82.845 116.285 ;
        RECT 83.015 115.675 83.185 116.455 ;
        RECT 83.715 116.295 83.885 116.525 ;
        RECT 83.355 116.125 83.885 116.295 ;
        RECT 83.355 115.845 83.575 116.125 ;
        RECT 84.055 115.955 84.295 116.355 ;
        RECT 83.015 115.505 83.420 115.675 ;
        RECT 83.755 115.585 84.295 115.955 ;
        RECT 84.465 116.170 84.785 116.525 ;
        RECT 84.465 115.915 84.790 116.170 ;
        RECT 84.985 116.095 85.155 116.905 ;
        RECT 85.325 116.255 85.655 116.735 ;
        RECT 85.825 116.435 85.995 116.905 ;
        RECT 86.165 116.255 86.495 116.735 ;
        RECT 86.665 116.435 86.835 116.905 ;
        RECT 85.325 116.085 87.090 116.255 ;
        RECT 87.315 116.180 87.605 116.905 ;
        RECT 88.275 116.085 88.505 116.905 ;
        RECT 88.675 116.105 89.005 116.735 ;
        RECT 84.465 115.705 86.495 115.915 ;
        RECT 84.465 115.695 84.810 115.705 ;
        RECT 82.115 115.335 82.790 115.495 ;
        RECT 83.250 115.415 83.420 115.505 ;
        RECT 82.115 115.325 83.080 115.335 ;
        RECT 81.755 115.155 81.925 115.295 ;
        RECT 78.500 114.355 78.750 114.815 ;
        RECT 78.920 114.525 79.170 114.855 ;
        RECT 79.385 114.525 80.065 114.855 ;
        RECT 80.235 114.955 81.310 115.125 ;
        RECT 81.755 114.985 82.315 115.155 ;
        RECT 82.620 115.035 83.080 115.325 ;
        RECT 83.250 115.245 84.470 115.415 ;
        RECT 80.235 114.615 80.405 114.955 ;
        RECT 80.640 114.355 80.970 114.785 ;
        RECT 81.140 114.615 81.310 114.955 ;
        RECT 81.605 114.355 81.975 114.815 ;
        RECT 82.145 114.525 82.315 114.985 ;
        RECT 83.250 114.865 83.420 115.245 ;
        RECT 84.640 115.075 84.810 115.695 ;
        RECT 86.680 115.535 87.090 116.085 ;
        RECT 88.255 115.665 88.585 115.915 ;
        RECT 82.550 114.525 83.420 114.865 ;
        RECT 84.010 114.905 84.810 115.075 ;
        RECT 83.590 114.355 83.840 114.815 ;
        RECT 84.010 114.615 84.180 114.905 ;
        RECT 84.360 114.355 84.690 114.735 ;
        RECT 84.985 114.355 85.155 115.415 ;
        RECT 85.365 115.365 87.090 115.535 ;
        RECT 85.365 114.525 85.655 115.365 ;
        RECT 85.825 114.355 85.995 115.195 ;
        RECT 86.205 114.525 86.455 115.365 ;
        RECT 86.665 114.355 86.835 115.195 ;
        RECT 87.315 114.355 87.605 115.520 ;
        RECT 88.755 115.505 89.005 116.105 ;
        RECT 89.175 116.085 89.385 116.905 ;
        RECT 89.925 116.435 90.095 116.905 ;
        RECT 90.265 116.255 90.595 116.735 ;
        RECT 90.765 116.435 90.935 116.905 ;
        RECT 91.105 116.255 91.435 116.735 ;
        RECT 89.670 116.085 91.435 116.255 ;
        RECT 91.605 116.095 91.775 116.905 ;
        RECT 91.975 116.525 93.045 116.695 ;
        RECT 91.975 116.170 92.295 116.525 ;
        RECT 88.275 114.355 88.505 115.495 ;
        RECT 88.675 114.525 89.005 115.505 ;
        RECT 89.670 115.535 90.080 116.085 ;
        RECT 91.970 115.915 92.295 116.170 ;
        RECT 90.265 115.705 92.295 115.915 ;
        RECT 91.950 115.695 92.295 115.705 ;
        RECT 92.465 115.955 92.705 116.355 ;
        RECT 92.875 116.295 93.045 116.525 ;
        RECT 93.215 116.465 93.405 116.905 ;
        RECT 93.575 116.455 94.525 116.735 ;
        RECT 94.745 116.545 95.095 116.715 ;
        RECT 92.875 116.125 93.405 116.295 ;
        RECT 89.175 114.355 89.385 115.495 ;
        RECT 89.670 115.365 91.395 115.535 ;
        RECT 89.925 114.355 90.095 115.195 ;
        RECT 90.305 114.525 90.555 115.365 ;
        RECT 90.765 114.355 90.935 115.195 ;
        RECT 91.105 114.525 91.395 115.365 ;
        RECT 91.605 114.355 91.775 115.415 ;
        RECT 91.950 115.075 92.120 115.695 ;
        RECT 92.465 115.585 93.005 115.955 ;
        RECT 93.185 115.845 93.405 116.125 ;
        RECT 93.575 115.675 93.745 116.455 ;
        RECT 93.340 115.505 93.745 115.675 ;
        RECT 93.915 115.665 94.265 116.285 ;
        RECT 93.340 115.415 93.510 115.505 ;
        RECT 94.435 115.495 94.645 116.285 ;
        RECT 92.290 115.245 93.510 115.415 ;
        RECT 93.970 115.335 94.645 115.495 ;
        RECT 91.950 114.905 92.750 115.075 ;
        RECT 92.070 114.355 92.400 114.735 ;
        RECT 92.580 114.615 92.750 114.905 ;
        RECT 93.340 114.865 93.510 115.245 ;
        RECT 93.680 115.325 94.645 115.335 ;
        RECT 94.835 116.155 95.095 116.545 ;
        RECT 95.305 116.445 95.635 116.905 ;
        RECT 96.510 116.515 97.365 116.685 ;
        RECT 97.570 116.515 98.065 116.685 ;
        RECT 98.235 116.545 98.565 116.905 ;
        RECT 94.835 115.465 95.005 116.155 ;
        RECT 95.175 115.805 95.345 115.985 ;
        RECT 95.515 115.975 96.305 116.225 ;
        RECT 96.510 115.805 96.680 116.515 ;
        RECT 96.850 116.005 97.205 116.225 ;
        RECT 95.175 115.635 96.865 115.805 ;
        RECT 93.680 115.035 94.140 115.325 ;
        RECT 94.835 115.295 96.335 115.465 ;
        RECT 94.835 115.155 95.005 115.295 ;
        RECT 94.445 114.985 95.005 115.155 ;
        RECT 92.920 114.355 93.170 114.815 ;
        RECT 93.340 114.525 94.210 114.865 ;
        RECT 94.445 114.525 94.615 114.985 ;
        RECT 95.450 114.955 96.525 115.125 ;
        RECT 94.785 114.355 95.155 114.815 ;
        RECT 95.450 114.615 95.620 114.955 ;
        RECT 95.790 114.355 96.120 114.785 ;
        RECT 96.355 114.615 96.525 114.955 ;
        RECT 96.695 114.855 96.865 115.635 ;
        RECT 97.035 115.415 97.205 116.005 ;
        RECT 97.375 115.605 97.725 116.225 ;
        RECT 97.035 115.025 97.500 115.415 ;
        RECT 97.895 115.155 98.065 116.515 ;
        RECT 98.235 115.325 98.695 116.375 ;
        RECT 97.670 114.985 98.065 115.155 ;
        RECT 97.670 114.855 97.840 114.985 ;
        RECT 96.695 114.525 97.375 114.855 ;
        RECT 97.590 114.525 97.840 114.855 ;
        RECT 98.010 114.355 98.260 114.815 ;
        RECT 98.430 114.540 98.755 115.325 ;
        RECT 98.925 114.525 99.095 116.645 ;
        RECT 99.265 116.525 99.595 116.905 ;
        RECT 99.765 116.355 100.020 116.645 ;
        RECT 99.270 116.185 100.020 116.355 ;
        RECT 99.270 115.195 99.500 116.185 ;
        RECT 100.195 116.180 100.485 116.905 ;
        RECT 101.580 116.355 101.835 116.645 ;
        RECT 102.005 116.525 102.335 116.905 ;
        RECT 101.580 116.185 102.330 116.355 ;
        RECT 99.670 115.365 100.020 116.015 ;
        RECT 99.270 115.025 100.020 115.195 ;
        RECT 99.265 114.355 99.595 114.855 ;
        RECT 99.765 114.525 100.020 115.025 ;
        RECT 100.195 114.355 100.485 115.520 ;
        RECT 101.580 115.365 101.930 116.015 ;
        RECT 102.100 115.195 102.330 116.185 ;
        RECT 101.580 115.025 102.330 115.195 ;
        RECT 101.580 114.525 101.835 115.025 ;
        RECT 102.005 114.355 102.335 114.855 ;
        RECT 102.505 114.525 102.675 116.645 ;
        RECT 103.035 116.545 103.365 116.905 ;
        RECT 103.535 116.515 104.030 116.685 ;
        RECT 104.235 116.515 105.090 116.685 ;
        RECT 102.905 115.325 103.365 116.375 ;
        RECT 102.845 114.540 103.170 115.325 ;
        RECT 103.535 115.155 103.705 116.515 ;
        RECT 103.875 115.605 104.225 116.225 ;
        RECT 104.395 116.005 104.750 116.225 ;
        RECT 104.395 115.415 104.565 116.005 ;
        RECT 104.920 115.805 105.090 116.515 ;
        RECT 105.965 116.445 106.295 116.905 ;
        RECT 106.505 116.545 106.855 116.715 ;
        RECT 105.295 115.975 106.085 116.225 ;
        RECT 106.505 116.155 106.765 116.545 ;
        RECT 107.075 116.455 108.025 116.735 ;
        RECT 108.195 116.465 108.385 116.905 ;
        RECT 108.555 116.525 109.625 116.695 ;
        RECT 106.255 115.805 106.425 115.985 ;
        RECT 103.535 114.985 103.930 115.155 ;
        RECT 104.100 115.025 104.565 115.415 ;
        RECT 104.735 115.635 106.425 115.805 ;
        RECT 103.760 114.855 103.930 114.985 ;
        RECT 104.735 114.855 104.905 115.635 ;
        RECT 106.595 115.465 106.765 116.155 ;
        RECT 105.265 115.295 106.765 115.465 ;
        RECT 106.955 115.495 107.165 116.285 ;
        RECT 107.335 115.665 107.685 116.285 ;
        RECT 107.855 115.675 108.025 116.455 ;
        RECT 108.555 116.295 108.725 116.525 ;
        RECT 108.195 116.125 108.725 116.295 ;
        RECT 108.195 115.845 108.415 116.125 ;
        RECT 108.895 115.955 109.135 116.355 ;
        RECT 107.855 115.505 108.260 115.675 ;
        RECT 108.595 115.585 109.135 115.955 ;
        RECT 109.305 116.170 109.625 116.525 ;
        RECT 109.305 115.915 109.630 116.170 ;
        RECT 109.825 116.095 109.995 116.905 ;
        RECT 110.165 116.255 110.495 116.735 ;
        RECT 110.665 116.435 110.835 116.905 ;
        RECT 111.005 116.255 111.335 116.735 ;
        RECT 111.505 116.435 111.675 116.905 ;
        RECT 110.165 116.085 111.930 116.255 ;
        RECT 112.155 116.155 113.365 116.905 ;
        RECT 109.305 115.705 111.335 115.915 ;
        RECT 109.305 115.695 109.650 115.705 ;
        RECT 106.955 115.335 107.630 115.495 ;
        RECT 108.090 115.415 108.260 115.505 ;
        RECT 106.955 115.325 107.920 115.335 ;
        RECT 106.595 115.155 106.765 115.295 ;
        RECT 103.340 114.355 103.590 114.815 ;
        RECT 103.760 114.525 104.010 114.855 ;
        RECT 104.225 114.525 104.905 114.855 ;
        RECT 105.075 114.955 106.150 115.125 ;
        RECT 106.595 114.985 107.155 115.155 ;
        RECT 107.460 115.035 107.920 115.325 ;
        RECT 108.090 115.245 109.310 115.415 ;
        RECT 105.075 114.615 105.245 114.955 ;
        RECT 105.480 114.355 105.810 114.785 ;
        RECT 105.980 114.615 106.150 114.955 ;
        RECT 106.445 114.355 106.815 114.815 ;
        RECT 106.985 114.525 107.155 114.985 ;
        RECT 108.090 114.865 108.260 115.245 ;
        RECT 109.480 115.075 109.650 115.695 ;
        RECT 111.520 115.535 111.930 116.085 ;
        RECT 107.390 114.525 108.260 114.865 ;
        RECT 108.850 114.905 109.650 115.075 ;
        RECT 108.430 114.355 108.680 114.815 ;
        RECT 108.850 114.615 109.020 114.905 ;
        RECT 109.200 114.355 109.530 114.735 ;
        RECT 109.825 114.355 109.995 115.415 ;
        RECT 110.205 115.365 111.930 115.535 ;
        RECT 112.155 115.445 112.675 115.985 ;
        RECT 112.845 115.615 113.365 116.155 ;
        RECT 110.205 114.525 110.495 115.365 ;
        RECT 110.665 114.355 110.835 115.195 ;
        RECT 111.045 114.525 111.295 115.365 ;
        RECT 111.505 114.355 111.675 115.195 ;
        RECT 112.155 114.355 113.365 115.445 ;
        RECT 22.830 114.185 113.450 114.355 ;
        RECT 19.165 66.070 30.165 66.940 ;
        RECT 19.165 54.930 20.835 66.070 ;
        RECT 21.465 65.555 26.465 65.725 ;
        RECT 21.235 55.300 21.405 65.340 ;
        RECT 26.525 55.300 26.695 65.340 ;
        RECT 27.095 54.930 27.265 66.070 ;
        RECT 27.895 65.555 28.895 65.725 ;
        RECT 27.665 55.300 27.835 65.340 ;
        RECT 28.955 55.300 29.125 65.340 ;
        RECT 29.525 54.930 30.165 66.070 ;
        RECT 19.165 52.860 30.165 54.930 ;
        RECT 19.165 49.370 21.005 52.860 ;
        RECT 22.765 52.780 30.165 52.860 ;
        RECT 21.635 52.350 22.135 52.520 ;
        RECT 21.405 50.095 21.575 52.135 ;
        RECT 22.195 50.095 22.365 52.135 ;
        RECT 21.635 49.710 22.135 49.880 ;
        RECT 22.765 49.370 25.085 52.780 ;
        RECT 25.715 52.270 26.215 52.440 ;
        RECT 19.165 48.650 25.085 49.370 ;
        RECT 19.135 48.040 23.045 48.260 ;
        RECT 19.135 45.640 20.855 48.040 ;
        RECT 21.485 47.530 21.985 47.700 ;
        RECT 21.255 46.320 21.425 47.360 ;
        RECT 22.045 46.320 22.215 47.360 ;
        RECT 21.485 45.980 21.985 46.150 ;
        RECT 22.615 45.640 23.045 48.040 ;
        RECT 24.025 46.290 25.085 48.650 ;
        RECT 25.485 47.015 25.655 52.055 ;
        RECT 26.275 47.015 26.445 52.055 ;
        RECT 25.715 46.630 26.215 46.800 ;
        RECT 26.845 46.290 27.015 52.780 ;
        RECT 27.645 52.270 28.145 52.440 ;
        RECT 27.415 47.015 27.585 52.055 ;
        RECT 28.205 47.015 28.375 52.055 ;
        RECT 27.645 46.630 28.145 46.800 ;
        RECT 28.775 46.290 30.165 52.780 ;
        RECT 30.365 66.080 41.365 66.950 ;
        RECT 30.365 54.940 32.035 66.080 ;
        RECT 32.665 65.565 37.665 65.735 ;
        RECT 32.435 55.310 32.605 65.350 ;
        RECT 37.725 55.310 37.895 65.350 ;
        RECT 38.295 54.940 38.465 66.080 ;
        RECT 39.095 65.565 40.095 65.735 ;
        RECT 38.865 55.310 39.035 65.350 ;
        RECT 40.155 55.310 40.325 65.350 ;
        RECT 40.725 54.940 41.365 66.080 ;
        RECT 30.365 52.870 41.365 54.940 ;
        RECT 30.365 49.380 32.205 52.870 ;
        RECT 33.965 52.790 41.365 52.870 ;
        RECT 32.835 52.360 33.335 52.530 ;
        RECT 32.605 50.105 32.775 52.145 ;
        RECT 33.395 50.105 33.565 52.145 ;
        RECT 32.835 49.720 33.335 49.890 ;
        RECT 33.965 49.380 36.285 52.790 ;
        RECT 36.915 52.280 37.415 52.450 ;
        RECT 30.365 48.660 36.285 49.380 ;
        RECT 24.025 45.800 30.165 46.290 ;
        RECT 30.335 48.050 34.245 48.270 ;
        RECT 19.135 45.370 23.045 45.640 ;
        RECT 30.335 45.650 32.055 48.050 ;
        RECT 32.685 47.540 33.185 47.710 ;
        RECT 32.455 46.330 32.625 47.370 ;
        RECT 33.245 46.330 33.415 47.370 ;
        RECT 32.685 45.990 33.185 46.160 ;
        RECT 33.815 45.650 34.245 48.050 ;
        RECT 35.225 46.300 36.285 48.660 ;
        RECT 36.685 47.025 36.855 52.065 ;
        RECT 37.475 47.025 37.645 52.065 ;
        RECT 36.915 46.640 37.415 46.810 ;
        RECT 38.045 46.300 38.215 52.790 ;
        RECT 38.845 52.280 39.345 52.450 ;
        RECT 38.615 47.025 38.785 52.065 ;
        RECT 39.405 47.025 39.575 52.065 ;
        RECT 38.845 46.640 39.345 46.810 ;
        RECT 39.975 46.300 41.365 52.790 ;
        RECT 41.585 66.050 52.585 66.920 ;
        RECT 41.585 54.910 43.255 66.050 ;
        RECT 43.885 65.535 48.885 65.705 ;
        RECT 43.655 55.280 43.825 65.320 ;
        RECT 48.945 55.280 49.115 65.320 ;
        RECT 49.515 54.910 49.685 66.050 ;
        RECT 50.315 65.535 51.315 65.705 ;
        RECT 50.085 55.280 50.255 65.320 ;
        RECT 51.375 55.280 51.545 65.320 ;
        RECT 51.945 54.910 52.585 66.050 ;
        RECT 41.585 52.840 52.585 54.910 ;
        RECT 41.585 49.350 43.425 52.840 ;
        RECT 45.185 52.760 52.585 52.840 ;
        RECT 44.055 52.330 44.555 52.500 ;
        RECT 43.825 50.075 43.995 52.115 ;
        RECT 44.615 50.075 44.785 52.115 ;
        RECT 44.055 49.690 44.555 49.860 ;
        RECT 45.185 49.350 47.505 52.760 ;
        RECT 48.135 52.250 48.635 52.420 ;
        RECT 41.585 48.630 47.505 49.350 ;
        RECT 35.225 45.810 41.365 46.300 ;
        RECT 41.555 48.020 45.465 48.240 ;
        RECT 30.335 45.380 34.245 45.650 ;
        RECT 41.555 45.620 43.275 48.020 ;
        RECT 43.905 47.510 44.405 47.680 ;
        RECT 43.675 46.300 43.845 47.340 ;
        RECT 44.465 46.300 44.635 47.340 ;
        RECT 43.905 45.960 44.405 46.130 ;
        RECT 45.035 45.620 45.465 48.020 ;
        RECT 46.445 46.270 47.505 48.630 ;
        RECT 47.905 46.995 48.075 52.035 ;
        RECT 48.695 46.995 48.865 52.035 ;
        RECT 48.135 46.610 48.635 46.780 ;
        RECT 49.265 46.270 49.435 52.760 ;
        RECT 50.065 52.250 50.565 52.420 ;
        RECT 49.835 46.995 50.005 52.035 ;
        RECT 50.625 46.995 50.795 52.035 ;
        RECT 50.065 46.610 50.565 46.780 ;
        RECT 51.195 46.270 52.585 52.760 ;
        RECT 52.835 66.030 63.835 66.900 ;
        RECT 52.835 54.890 54.505 66.030 ;
        RECT 55.135 65.515 60.135 65.685 ;
        RECT 54.905 55.260 55.075 65.300 ;
        RECT 60.195 55.260 60.365 65.300 ;
        RECT 60.765 54.890 60.935 66.030 ;
        RECT 61.565 65.515 62.565 65.685 ;
        RECT 61.335 55.260 61.505 65.300 ;
        RECT 62.625 55.260 62.795 65.300 ;
        RECT 63.195 54.890 63.835 66.030 ;
        RECT 52.835 52.820 63.835 54.890 ;
        RECT 52.835 49.330 54.675 52.820 ;
        RECT 56.435 52.740 63.835 52.820 ;
        RECT 55.305 52.310 55.805 52.480 ;
        RECT 55.075 50.055 55.245 52.095 ;
        RECT 55.865 50.055 56.035 52.095 ;
        RECT 55.305 49.670 55.805 49.840 ;
        RECT 56.435 49.330 58.755 52.740 ;
        RECT 59.385 52.230 59.885 52.400 ;
        RECT 52.835 48.610 58.755 49.330 ;
        RECT 46.445 45.780 52.585 46.270 ;
        RECT 52.805 48.000 56.715 48.220 ;
        RECT 41.555 45.350 45.465 45.620 ;
        RECT 52.805 45.600 54.525 48.000 ;
        RECT 55.155 47.490 55.655 47.660 ;
        RECT 54.925 46.280 55.095 47.320 ;
        RECT 55.715 46.280 55.885 47.320 ;
        RECT 55.155 45.940 55.655 46.110 ;
        RECT 56.285 45.600 56.715 48.000 ;
        RECT 57.695 46.250 58.755 48.610 ;
        RECT 59.155 46.975 59.325 52.015 ;
        RECT 59.945 46.975 60.115 52.015 ;
        RECT 59.385 46.590 59.885 46.760 ;
        RECT 60.515 46.250 60.685 52.740 ;
        RECT 61.315 52.230 61.815 52.400 ;
        RECT 61.085 46.975 61.255 52.015 ;
        RECT 61.875 46.975 62.045 52.015 ;
        RECT 61.315 46.590 61.815 46.760 ;
        RECT 62.445 46.250 63.835 52.740 ;
        RECT 64.055 66.020 75.055 66.890 ;
        RECT 64.055 54.880 65.725 66.020 ;
        RECT 66.355 65.505 71.355 65.675 ;
        RECT 66.125 55.250 66.295 65.290 ;
        RECT 71.415 55.250 71.585 65.290 ;
        RECT 71.985 54.880 72.155 66.020 ;
        RECT 72.785 65.505 73.785 65.675 ;
        RECT 72.555 55.250 72.725 65.290 ;
        RECT 73.845 55.250 74.015 65.290 ;
        RECT 74.415 54.880 75.055 66.020 ;
        RECT 64.055 52.810 75.055 54.880 ;
        RECT 64.055 49.320 65.895 52.810 ;
        RECT 67.655 52.730 75.055 52.810 ;
        RECT 66.525 52.300 67.025 52.470 ;
        RECT 66.295 50.045 66.465 52.085 ;
        RECT 67.085 50.045 67.255 52.085 ;
        RECT 66.525 49.660 67.025 49.830 ;
        RECT 67.655 49.320 69.975 52.730 ;
        RECT 70.605 52.220 71.105 52.390 ;
        RECT 64.055 48.600 69.975 49.320 ;
        RECT 57.695 45.760 63.835 46.250 ;
        RECT 64.025 47.990 67.935 48.210 ;
        RECT 52.805 45.330 56.715 45.600 ;
        RECT 64.025 45.590 65.745 47.990 ;
        RECT 66.375 47.480 66.875 47.650 ;
        RECT 66.145 46.270 66.315 47.310 ;
        RECT 66.935 46.270 67.105 47.310 ;
        RECT 66.375 45.930 66.875 46.100 ;
        RECT 67.505 45.590 67.935 47.990 ;
        RECT 68.915 46.240 69.975 48.600 ;
        RECT 70.375 46.965 70.545 52.005 ;
        RECT 71.165 46.965 71.335 52.005 ;
        RECT 70.605 46.580 71.105 46.750 ;
        RECT 71.735 46.240 71.905 52.730 ;
        RECT 72.535 52.220 73.035 52.390 ;
        RECT 72.305 46.965 72.475 52.005 ;
        RECT 73.095 46.965 73.265 52.005 ;
        RECT 72.535 46.580 73.035 46.750 ;
        RECT 73.665 46.240 75.055 52.730 ;
        RECT 75.295 66.010 86.295 66.880 ;
        RECT 75.295 54.870 76.965 66.010 ;
        RECT 77.595 65.495 82.595 65.665 ;
        RECT 77.365 55.240 77.535 65.280 ;
        RECT 82.655 55.240 82.825 65.280 ;
        RECT 83.225 54.870 83.395 66.010 ;
        RECT 84.025 65.495 85.025 65.665 ;
        RECT 83.795 55.240 83.965 65.280 ;
        RECT 85.085 55.240 85.255 65.280 ;
        RECT 85.655 54.870 86.295 66.010 ;
        RECT 75.295 52.800 86.295 54.870 ;
        RECT 75.295 49.310 77.135 52.800 ;
        RECT 78.895 52.720 86.295 52.800 ;
        RECT 77.765 52.290 78.265 52.460 ;
        RECT 77.535 50.035 77.705 52.075 ;
        RECT 78.325 50.035 78.495 52.075 ;
        RECT 77.765 49.650 78.265 49.820 ;
        RECT 78.895 49.310 81.215 52.720 ;
        RECT 81.845 52.210 82.345 52.380 ;
        RECT 75.295 48.590 81.215 49.310 ;
        RECT 68.915 45.750 75.055 46.240 ;
        RECT 75.265 47.980 79.175 48.200 ;
        RECT 64.025 45.320 67.935 45.590 ;
        RECT 75.265 45.580 76.985 47.980 ;
        RECT 77.615 47.470 78.115 47.640 ;
        RECT 77.385 46.260 77.555 47.300 ;
        RECT 78.175 46.260 78.345 47.300 ;
        RECT 77.615 45.920 78.115 46.090 ;
        RECT 78.745 45.580 79.175 47.980 ;
        RECT 80.155 46.230 81.215 48.590 ;
        RECT 81.615 46.955 81.785 51.995 ;
        RECT 82.405 46.955 82.575 51.995 ;
        RECT 81.845 46.570 82.345 46.740 ;
        RECT 82.975 46.230 83.145 52.720 ;
        RECT 83.775 52.210 84.275 52.380 ;
        RECT 83.545 46.955 83.715 51.995 ;
        RECT 84.335 46.955 84.505 51.995 ;
        RECT 83.775 46.570 84.275 46.740 ;
        RECT 84.905 46.230 86.295 52.720 ;
        RECT 86.545 66.020 97.545 66.890 ;
        RECT 131.125 66.880 140.025 66.890 ;
        RECT 86.545 54.880 88.215 66.020 ;
        RECT 88.845 65.505 93.845 65.675 ;
        RECT 88.615 55.250 88.785 65.290 ;
        RECT 93.905 55.250 94.075 65.290 ;
        RECT 94.475 54.880 94.645 66.020 ;
        RECT 95.275 65.505 96.275 65.675 ;
        RECT 95.045 55.250 95.215 65.290 ;
        RECT 96.335 55.250 96.505 65.290 ;
        RECT 96.905 54.880 97.545 66.020 ;
        RECT 86.545 52.810 97.545 54.880 ;
        RECT 86.545 49.320 88.385 52.810 ;
        RECT 90.145 52.730 97.545 52.810 ;
        RECT 89.015 52.300 89.515 52.470 ;
        RECT 88.785 50.045 88.955 52.085 ;
        RECT 89.575 50.045 89.745 52.085 ;
        RECT 89.015 49.660 89.515 49.830 ;
        RECT 90.145 49.320 92.465 52.730 ;
        RECT 93.095 52.220 93.595 52.390 ;
        RECT 86.545 48.600 92.465 49.320 ;
        RECT 80.155 45.740 86.295 46.230 ;
        RECT 86.515 47.990 90.425 48.210 ;
        RECT 75.265 45.310 79.175 45.580 ;
        RECT 86.515 45.590 88.235 47.990 ;
        RECT 88.865 47.480 89.365 47.650 ;
        RECT 88.635 46.270 88.805 47.310 ;
        RECT 89.425 46.270 89.595 47.310 ;
        RECT 88.865 45.930 89.365 46.100 ;
        RECT 89.995 45.590 90.425 47.990 ;
        RECT 91.405 46.240 92.465 48.600 ;
        RECT 92.865 46.965 93.035 52.005 ;
        RECT 93.655 46.965 93.825 52.005 ;
        RECT 93.095 46.580 93.595 46.750 ;
        RECT 94.225 46.240 94.395 52.730 ;
        RECT 95.025 52.220 95.525 52.390 ;
        RECT 94.795 46.965 94.965 52.005 ;
        RECT 95.585 46.965 95.755 52.005 ;
        RECT 95.025 46.580 95.525 46.750 ;
        RECT 96.155 46.240 97.545 52.730 ;
        RECT 97.825 66.010 108.825 66.880 ;
        RECT 97.825 54.870 99.495 66.010 ;
        RECT 100.125 65.495 105.125 65.665 ;
        RECT 99.895 55.240 100.065 65.280 ;
        RECT 105.185 55.240 105.355 65.280 ;
        RECT 105.755 54.870 105.925 66.010 ;
        RECT 106.555 65.495 107.555 65.665 ;
        RECT 106.325 55.240 106.495 65.280 ;
        RECT 107.615 55.240 107.785 65.280 ;
        RECT 108.185 54.870 108.825 66.010 ;
        RECT 97.825 52.800 108.825 54.870 ;
        RECT 97.825 49.310 99.665 52.800 ;
        RECT 101.425 52.720 108.825 52.800 ;
        RECT 100.295 52.290 100.795 52.460 ;
        RECT 100.065 50.035 100.235 52.075 ;
        RECT 100.855 50.035 101.025 52.075 ;
        RECT 100.295 49.650 100.795 49.820 ;
        RECT 101.425 49.310 103.745 52.720 ;
        RECT 104.375 52.210 104.875 52.380 ;
        RECT 97.825 48.590 103.745 49.310 ;
        RECT 91.405 45.750 97.545 46.240 ;
        RECT 97.795 47.980 101.705 48.200 ;
        RECT 86.515 45.320 90.425 45.590 ;
        RECT 97.795 45.580 99.515 47.980 ;
        RECT 100.145 47.470 100.645 47.640 ;
        RECT 99.915 46.260 100.085 47.300 ;
        RECT 100.705 46.260 100.875 47.300 ;
        RECT 100.145 45.920 100.645 46.090 ;
        RECT 101.275 45.580 101.705 47.980 ;
        RECT 102.685 46.230 103.745 48.590 ;
        RECT 104.145 46.955 104.315 51.995 ;
        RECT 104.935 46.955 105.105 51.995 ;
        RECT 104.375 46.570 104.875 46.740 ;
        RECT 105.505 46.230 105.675 52.720 ;
        RECT 106.305 52.210 106.805 52.380 ;
        RECT 106.075 46.955 106.245 51.995 ;
        RECT 106.865 46.955 107.035 51.995 ;
        RECT 106.305 46.570 106.805 46.740 ;
        RECT 107.435 46.230 108.825 52.720 ;
        RECT 109.095 66.010 120.095 66.880 ;
        RECT 109.095 54.870 110.765 66.010 ;
        RECT 111.395 65.495 116.395 65.665 ;
        RECT 111.165 55.240 111.335 65.280 ;
        RECT 116.455 55.240 116.625 65.280 ;
        RECT 117.025 54.870 117.195 66.010 ;
        RECT 117.825 65.495 118.825 65.665 ;
        RECT 117.595 55.240 117.765 65.280 ;
        RECT 118.885 55.240 119.055 65.280 ;
        RECT 119.455 54.870 120.095 66.010 ;
        RECT 109.095 52.800 120.095 54.870 ;
        RECT 109.095 49.310 110.935 52.800 ;
        RECT 112.695 52.720 120.095 52.800 ;
        RECT 111.565 52.290 112.065 52.460 ;
        RECT 111.335 50.035 111.505 52.075 ;
        RECT 112.125 50.035 112.295 52.075 ;
        RECT 111.565 49.650 112.065 49.820 ;
        RECT 112.695 49.310 115.015 52.720 ;
        RECT 115.645 52.210 116.145 52.380 ;
        RECT 109.095 48.590 115.015 49.310 ;
        RECT 102.685 45.740 108.825 46.230 ;
        RECT 109.065 47.980 112.975 48.200 ;
        RECT 97.795 45.310 101.705 45.580 ;
        RECT 109.065 45.580 110.785 47.980 ;
        RECT 111.415 47.470 111.915 47.640 ;
        RECT 111.185 46.260 111.355 47.300 ;
        RECT 111.975 46.260 112.145 47.300 ;
        RECT 111.415 45.920 111.915 46.090 ;
        RECT 112.545 45.580 112.975 47.980 ;
        RECT 113.955 46.230 115.015 48.590 ;
        RECT 115.415 46.955 115.585 51.995 ;
        RECT 116.205 46.955 116.375 51.995 ;
        RECT 115.645 46.570 116.145 46.740 ;
        RECT 116.775 46.230 116.945 52.720 ;
        RECT 117.575 52.210 118.075 52.380 ;
        RECT 117.345 46.955 117.515 51.995 ;
        RECT 118.135 46.955 118.305 51.995 ;
        RECT 117.575 46.570 118.075 46.740 ;
        RECT 118.705 46.230 120.095 52.720 ;
        RECT 120.345 66.010 140.025 66.880 ;
        RECT 120.345 54.870 122.015 66.010 ;
        RECT 122.645 65.495 127.645 65.665 ;
        RECT 122.415 55.240 122.585 65.280 ;
        RECT 127.705 55.240 127.875 65.280 ;
        RECT 128.275 54.870 128.445 66.010 ;
        RECT 130.705 65.980 140.025 66.010 ;
        RECT 129.075 65.495 130.075 65.665 ;
        RECT 128.845 55.240 129.015 65.280 ;
        RECT 130.135 55.240 130.305 65.280 ;
        RECT 130.705 54.870 132.765 65.980 ;
        RECT 133.395 65.465 138.395 65.635 ;
        RECT 133.165 55.210 133.335 65.250 ;
        RECT 138.455 55.210 138.625 65.250 ;
        RECT 120.345 54.840 132.765 54.870 ;
        RECT 139.025 54.840 140.025 65.980 ;
        RECT 120.345 54.720 140.025 54.840 ;
        RECT 120.345 53.550 140.035 54.720 ;
        RECT 120.345 52.800 131.345 53.550 ;
        RECT 120.345 49.310 122.185 52.800 ;
        RECT 123.945 52.720 131.345 52.800 ;
        RECT 122.815 52.290 123.315 52.460 ;
        RECT 122.585 50.035 122.755 52.075 ;
        RECT 123.375 50.035 123.545 52.075 ;
        RECT 122.815 49.650 123.315 49.820 ;
        RECT 123.945 49.310 126.265 52.720 ;
        RECT 126.895 52.210 127.395 52.380 ;
        RECT 120.345 48.590 126.265 49.310 ;
        RECT 113.955 45.740 120.095 46.230 ;
        RECT 120.315 47.980 124.225 48.200 ;
        RECT 109.065 45.310 112.975 45.580 ;
        RECT 120.315 45.580 122.035 47.980 ;
        RECT 122.665 47.470 123.165 47.640 ;
        RECT 122.435 46.260 122.605 47.300 ;
        RECT 123.225 46.260 123.395 47.300 ;
        RECT 122.665 45.920 123.165 46.090 ;
        RECT 123.795 45.580 124.225 47.980 ;
        RECT 125.205 46.230 126.265 48.590 ;
        RECT 126.665 46.955 126.835 51.995 ;
        RECT 127.455 46.955 127.625 51.995 ;
        RECT 126.895 46.570 127.395 46.740 ;
        RECT 128.025 46.230 128.195 52.720 ;
        RECT 128.825 52.210 129.325 52.380 ;
        RECT 128.595 46.955 128.765 51.995 ;
        RECT 129.385 46.955 129.555 51.995 ;
        RECT 128.825 46.570 129.325 46.740 ;
        RECT 129.955 46.230 131.345 52.720 ;
        RECT 125.205 45.740 131.345 46.230 ;
        RECT 120.315 45.310 124.225 45.580 ;
        RECT 25.695 39.770 29.605 40.040 ;
        RECT 18.575 39.120 24.715 39.610 ;
        RECT 18.575 32.630 19.965 39.120 ;
        RECT 20.595 38.610 21.095 38.780 ;
        RECT 20.365 33.355 20.535 38.395 ;
        RECT 21.155 33.355 21.325 38.395 ;
        RECT 20.595 32.970 21.095 33.140 ;
        RECT 21.725 32.630 21.895 39.120 ;
        RECT 22.525 38.610 23.025 38.780 ;
        RECT 22.295 33.355 22.465 38.395 ;
        RECT 23.085 33.355 23.255 38.395 ;
        RECT 23.655 36.760 24.715 39.120 ;
        RECT 25.695 37.370 26.125 39.770 ;
        RECT 26.755 39.260 27.255 39.430 ;
        RECT 26.525 38.050 26.695 39.090 ;
        RECT 27.315 38.050 27.485 39.090 ;
        RECT 26.755 37.710 27.255 37.880 ;
        RECT 27.885 37.370 29.605 39.770 ;
        RECT 36.975 39.770 40.885 40.040 ;
        RECT 25.695 37.150 29.605 37.370 ;
        RECT 29.855 39.120 35.995 39.610 ;
        RECT 23.655 36.040 29.575 36.760 ;
        RECT 22.525 32.970 23.025 33.140 ;
        RECT 23.655 32.630 25.975 36.040 ;
        RECT 26.605 35.530 27.105 35.700 ;
        RECT 26.375 33.275 26.545 35.315 ;
        RECT 27.165 33.275 27.335 35.315 ;
        RECT 26.605 32.890 27.105 33.060 ;
        RECT 18.575 32.550 25.975 32.630 ;
        RECT 27.735 32.550 29.575 36.040 ;
        RECT 18.575 30.480 29.575 32.550 ;
        RECT 18.575 19.340 19.215 30.480 ;
        RECT 19.615 20.070 19.785 30.110 ;
        RECT 20.905 20.070 21.075 30.110 ;
        RECT 19.845 19.685 20.845 19.855 ;
        RECT 21.475 19.340 21.645 30.480 ;
        RECT 22.045 20.070 22.215 30.110 ;
        RECT 27.335 20.070 27.505 30.110 ;
        RECT 22.275 19.685 27.275 19.855 ;
        RECT 27.905 19.340 29.575 30.480 ;
        RECT 18.575 18.470 29.575 19.340 ;
        RECT 29.855 32.630 31.245 39.120 ;
        RECT 31.875 38.610 32.375 38.780 ;
        RECT 31.645 33.355 31.815 38.395 ;
        RECT 32.435 33.355 32.605 38.395 ;
        RECT 31.875 32.970 32.375 33.140 ;
        RECT 33.005 32.630 33.175 39.120 ;
        RECT 33.805 38.610 34.305 38.780 ;
        RECT 33.575 33.355 33.745 38.395 ;
        RECT 34.365 33.355 34.535 38.395 ;
        RECT 34.935 36.760 35.995 39.120 ;
        RECT 36.975 37.370 37.405 39.770 ;
        RECT 38.035 39.260 38.535 39.430 ;
        RECT 37.805 38.050 37.975 39.090 ;
        RECT 38.595 38.050 38.765 39.090 ;
        RECT 38.035 37.710 38.535 37.880 ;
        RECT 39.165 37.370 40.885 39.770 ;
        RECT 48.265 39.750 52.175 40.020 ;
        RECT 36.975 37.150 40.885 37.370 ;
        RECT 41.145 39.100 47.285 39.590 ;
        RECT 34.935 36.040 40.855 36.760 ;
        RECT 33.805 32.970 34.305 33.140 ;
        RECT 34.935 32.630 37.255 36.040 ;
        RECT 37.885 35.530 38.385 35.700 ;
        RECT 37.655 33.275 37.825 35.315 ;
        RECT 38.445 33.275 38.615 35.315 ;
        RECT 37.885 32.890 38.385 33.060 ;
        RECT 29.855 32.550 37.255 32.630 ;
        RECT 39.015 32.550 40.855 36.040 ;
        RECT 29.855 30.480 40.855 32.550 ;
        RECT 29.855 19.340 30.495 30.480 ;
        RECT 30.895 20.070 31.065 30.110 ;
        RECT 32.185 20.070 32.355 30.110 ;
        RECT 31.125 19.685 32.125 19.855 ;
        RECT 32.755 19.340 32.925 30.480 ;
        RECT 33.325 20.070 33.495 30.110 ;
        RECT 38.615 20.070 38.785 30.110 ;
        RECT 33.555 19.685 38.555 19.855 ;
        RECT 39.185 19.340 40.855 30.480 ;
        RECT 29.855 18.470 40.855 19.340 ;
        RECT 41.145 32.610 42.535 39.100 ;
        RECT 43.165 38.590 43.665 38.760 ;
        RECT 42.935 33.335 43.105 38.375 ;
        RECT 43.725 33.335 43.895 38.375 ;
        RECT 43.165 32.950 43.665 33.120 ;
        RECT 44.295 32.610 44.465 39.100 ;
        RECT 45.095 38.590 45.595 38.760 ;
        RECT 44.865 33.335 45.035 38.375 ;
        RECT 45.655 33.335 45.825 38.375 ;
        RECT 46.225 36.740 47.285 39.100 ;
        RECT 48.265 37.350 48.695 39.750 ;
        RECT 49.325 39.240 49.825 39.410 ;
        RECT 49.095 38.030 49.265 39.070 ;
        RECT 49.885 38.030 50.055 39.070 ;
        RECT 49.325 37.690 49.825 37.860 ;
        RECT 50.455 37.350 52.175 39.750 ;
        RECT 59.485 39.750 63.395 40.020 ;
        RECT 48.265 37.130 52.175 37.350 ;
        RECT 52.365 39.100 58.505 39.590 ;
        RECT 46.225 36.020 52.145 36.740 ;
        RECT 45.095 32.950 45.595 33.120 ;
        RECT 46.225 32.610 48.545 36.020 ;
        RECT 49.175 35.510 49.675 35.680 ;
        RECT 48.945 33.255 49.115 35.295 ;
        RECT 49.735 33.255 49.905 35.295 ;
        RECT 49.175 32.870 49.675 33.040 ;
        RECT 41.145 32.530 48.545 32.610 ;
        RECT 50.305 32.530 52.145 36.020 ;
        RECT 41.145 30.460 52.145 32.530 ;
        RECT 41.145 19.320 41.785 30.460 ;
        RECT 42.185 20.050 42.355 30.090 ;
        RECT 43.475 20.050 43.645 30.090 ;
        RECT 42.415 19.665 43.415 19.835 ;
        RECT 44.045 19.320 44.215 30.460 ;
        RECT 44.615 20.050 44.785 30.090 ;
        RECT 49.905 20.050 50.075 30.090 ;
        RECT 44.845 19.665 49.845 19.835 ;
        RECT 50.475 19.320 52.145 30.460 ;
        RECT 41.145 18.450 52.145 19.320 ;
        RECT 52.365 32.610 53.755 39.100 ;
        RECT 54.385 38.590 54.885 38.760 ;
        RECT 54.155 33.335 54.325 38.375 ;
        RECT 54.945 33.335 55.115 38.375 ;
        RECT 54.385 32.950 54.885 33.120 ;
        RECT 55.515 32.610 55.685 39.100 ;
        RECT 56.315 38.590 56.815 38.760 ;
        RECT 56.085 33.335 56.255 38.375 ;
        RECT 56.875 33.335 57.045 38.375 ;
        RECT 57.445 36.740 58.505 39.100 ;
        RECT 59.485 37.350 59.915 39.750 ;
        RECT 60.545 39.240 61.045 39.410 ;
        RECT 60.315 38.030 60.485 39.070 ;
        RECT 61.105 38.030 61.275 39.070 ;
        RECT 60.545 37.690 61.045 37.860 ;
        RECT 61.675 37.350 63.395 39.750 ;
        RECT 70.685 39.750 74.595 40.020 ;
        RECT 59.485 37.130 63.395 37.350 ;
        RECT 63.565 39.100 69.705 39.590 ;
        RECT 57.445 36.020 63.365 36.740 ;
        RECT 56.315 32.950 56.815 33.120 ;
        RECT 57.445 32.610 59.765 36.020 ;
        RECT 60.395 35.510 60.895 35.680 ;
        RECT 60.165 33.255 60.335 35.295 ;
        RECT 60.955 33.255 61.125 35.295 ;
        RECT 60.395 32.870 60.895 33.040 ;
        RECT 52.365 32.530 59.765 32.610 ;
        RECT 61.525 32.530 63.365 36.020 ;
        RECT 52.365 30.460 63.365 32.530 ;
        RECT 52.365 19.320 53.005 30.460 ;
        RECT 53.405 20.050 53.575 30.090 ;
        RECT 54.695 20.050 54.865 30.090 ;
        RECT 53.635 19.665 54.635 19.835 ;
        RECT 55.265 19.320 55.435 30.460 ;
        RECT 55.835 20.050 56.005 30.090 ;
        RECT 61.125 20.050 61.295 30.090 ;
        RECT 56.065 19.665 61.065 19.835 ;
        RECT 61.695 19.320 63.365 30.460 ;
        RECT 52.365 18.450 63.365 19.320 ;
        RECT 63.565 32.610 64.955 39.100 ;
        RECT 65.585 38.590 66.085 38.760 ;
        RECT 65.355 33.335 65.525 38.375 ;
        RECT 66.145 33.335 66.315 38.375 ;
        RECT 65.585 32.950 66.085 33.120 ;
        RECT 66.715 32.610 66.885 39.100 ;
        RECT 67.515 38.590 68.015 38.760 ;
        RECT 67.285 33.335 67.455 38.375 ;
        RECT 68.075 33.335 68.245 38.375 ;
        RECT 68.645 36.740 69.705 39.100 ;
        RECT 70.685 37.350 71.115 39.750 ;
        RECT 71.745 39.240 72.245 39.410 ;
        RECT 71.515 38.030 71.685 39.070 ;
        RECT 72.305 38.030 72.475 39.070 ;
        RECT 71.745 37.690 72.245 37.860 ;
        RECT 72.875 37.350 74.595 39.750 ;
        RECT 81.975 39.740 85.885 40.010 ;
        RECT 70.685 37.130 74.595 37.350 ;
        RECT 74.855 39.090 80.995 39.580 ;
        RECT 68.645 36.020 74.565 36.740 ;
        RECT 67.515 32.950 68.015 33.120 ;
        RECT 68.645 32.610 70.965 36.020 ;
        RECT 71.595 35.510 72.095 35.680 ;
        RECT 71.365 33.255 71.535 35.295 ;
        RECT 72.155 33.255 72.325 35.295 ;
        RECT 71.595 32.870 72.095 33.040 ;
        RECT 63.565 32.530 70.965 32.610 ;
        RECT 72.725 32.530 74.565 36.020 ;
        RECT 63.565 30.460 74.565 32.530 ;
        RECT 63.565 19.320 64.205 30.460 ;
        RECT 64.605 20.050 64.775 30.090 ;
        RECT 65.895 20.050 66.065 30.090 ;
        RECT 64.835 19.665 65.835 19.835 ;
        RECT 66.465 19.320 66.635 30.460 ;
        RECT 67.035 20.050 67.205 30.090 ;
        RECT 72.325 20.050 72.495 30.090 ;
        RECT 67.265 19.665 72.265 19.835 ;
        RECT 72.895 19.320 74.565 30.460 ;
        RECT 63.565 18.450 74.565 19.320 ;
        RECT 74.855 32.600 76.245 39.090 ;
        RECT 76.875 38.580 77.375 38.750 ;
        RECT 76.645 33.325 76.815 38.365 ;
        RECT 77.435 33.325 77.605 38.365 ;
        RECT 76.875 32.940 77.375 33.110 ;
        RECT 78.005 32.600 78.175 39.090 ;
        RECT 78.805 38.580 79.305 38.750 ;
        RECT 78.575 33.325 78.745 38.365 ;
        RECT 79.365 33.325 79.535 38.365 ;
        RECT 79.935 36.730 80.995 39.090 ;
        RECT 81.975 37.340 82.405 39.740 ;
        RECT 83.035 39.230 83.535 39.400 ;
        RECT 82.805 38.020 82.975 39.060 ;
        RECT 83.595 38.020 83.765 39.060 ;
        RECT 83.035 37.680 83.535 37.850 ;
        RECT 84.165 37.340 85.885 39.740 ;
        RECT 93.215 39.760 97.125 40.030 ;
        RECT 81.975 37.120 85.885 37.340 ;
        RECT 86.095 39.110 92.235 39.600 ;
        RECT 79.935 36.010 85.855 36.730 ;
        RECT 78.805 32.940 79.305 33.110 ;
        RECT 79.935 32.600 82.255 36.010 ;
        RECT 82.885 35.500 83.385 35.670 ;
        RECT 82.655 33.245 82.825 35.285 ;
        RECT 83.445 33.245 83.615 35.285 ;
        RECT 82.885 32.860 83.385 33.030 ;
        RECT 74.855 32.520 82.255 32.600 ;
        RECT 84.015 32.520 85.855 36.010 ;
        RECT 74.855 30.450 85.855 32.520 ;
        RECT 74.855 19.310 75.495 30.450 ;
        RECT 75.895 20.040 76.065 30.080 ;
        RECT 77.185 20.040 77.355 30.080 ;
        RECT 76.125 19.655 77.125 19.825 ;
        RECT 77.755 19.310 77.925 30.450 ;
        RECT 78.325 20.040 78.495 30.080 ;
        RECT 83.615 20.040 83.785 30.080 ;
        RECT 78.555 19.655 83.555 19.825 ;
        RECT 84.185 19.310 85.855 30.450 ;
        RECT 74.855 18.440 85.855 19.310 ;
        RECT 86.095 32.620 87.485 39.110 ;
        RECT 88.115 38.600 88.615 38.770 ;
        RECT 87.885 33.345 88.055 38.385 ;
        RECT 88.675 33.345 88.845 38.385 ;
        RECT 88.115 32.960 88.615 33.130 ;
        RECT 89.245 32.620 89.415 39.110 ;
        RECT 90.045 38.600 90.545 38.770 ;
        RECT 89.815 33.345 89.985 38.385 ;
        RECT 90.605 33.345 90.775 38.385 ;
        RECT 91.175 36.750 92.235 39.110 ;
        RECT 93.215 37.360 93.645 39.760 ;
        RECT 94.275 39.250 94.775 39.420 ;
        RECT 94.045 38.040 94.215 39.080 ;
        RECT 94.835 38.040 95.005 39.080 ;
        RECT 94.275 37.700 94.775 37.870 ;
        RECT 95.405 37.360 97.125 39.760 ;
        RECT 104.425 39.780 108.335 40.050 ;
        RECT 93.215 37.140 97.125 37.360 ;
        RECT 97.305 39.130 103.445 39.620 ;
        RECT 91.175 36.030 97.095 36.750 ;
        RECT 90.045 32.960 90.545 33.130 ;
        RECT 91.175 32.620 93.495 36.030 ;
        RECT 94.125 35.520 94.625 35.690 ;
        RECT 93.895 33.265 94.065 35.305 ;
        RECT 94.685 33.265 94.855 35.305 ;
        RECT 94.125 32.880 94.625 33.050 ;
        RECT 86.095 32.540 93.495 32.620 ;
        RECT 95.255 32.540 97.095 36.030 ;
        RECT 86.095 30.470 97.095 32.540 ;
        RECT 86.095 19.330 86.735 30.470 ;
        RECT 87.135 20.060 87.305 30.100 ;
        RECT 88.425 20.060 88.595 30.100 ;
        RECT 87.365 19.675 88.365 19.845 ;
        RECT 88.995 19.330 89.165 30.470 ;
        RECT 89.565 20.060 89.735 30.100 ;
        RECT 94.855 20.060 95.025 30.100 ;
        RECT 89.795 19.675 94.795 19.845 ;
        RECT 95.425 19.330 97.095 30.470 ;
        RECT 86.095 18.460 97.095 19.330 ;
        RECT 97.305 32.640 98.695 39.130 ;
        RECT 99.325 38.620 99.825 38.790 ;
        RECT 99.095 33.365 99.265 38.405 ;
        RECT 99.885 33.365 100.055 38.405 ;
        RECT 99.325 32.980 99.825 33.150 ;
        RECT 100.455 32.640 100.625 39.130 ;
        RECT 101.255 38.620 101.755 38.790 ;
        RECT 101.025 33.365 101.195 38.405 ;
        RECT 101.815 33.365 101.985 38.405 ;
        RECT 102.385 36.770 103.445 39.130 ;
        RECT 104.425 37.380 104.855 39.780 ;
        RECT 105.485 39.270 105.985 39.440 ;
        RECT 105.255 38.060 105.425 39.100 ;
        RECT 106.045 38.060 106.215 39.100 ;
        RECT 105.485 37.720 105.985 37.890 ;
        RECT 106.615 37.380 108.335 39.780 ;
        RECT 115.625 39.820 119.535 40.090 ;
        RECT 104.425 37.160 108.335 37.380 ;
        RECT 108.505 39.170 114.645 39.660 ;
        RECT 102.385 36.050 108.305 36.770 ;
        RECT 101.255 32.980 101.755 33.150 ;
        RECT 102.385 32.640 104.705 36.050 ;
        RECT 105.335 35.540 105.835 35.710 ;
        RECT 105.105 33.285 105.275 35.325 ;
        RECT 105.895 33.285 106.065 35.325 ;
        RECT 105.335 32.900 105.835 33.070 ;
        RECT 97.305 32.560 104.705 32.640 ;
        RECT 106.465 32.560 108.305 36.050 ;
        RECT 97.305 30.490 108.305 32.560 ;
        RECT 97.305 19.350 97.945 30.490 ;
        RECT 98.345 20.080 98.515 30.120 ;
        RECT 99.635 20.080 99.805 30.120 ;
        RECT 98.575 19.695 99.575 19.865 ;
        RECT 100.205 19.350 100.375 30.490 ;
        RECT 100.775 20.080 100.945 30.120 ;
        RECT 106.065 20.080 106.235 30.120 ;
        RECT 101.005 19.695 106.005 19.865 ;
        RECT 106.635 19.350 108.305 30.490 ;
        RECT 97.305 18.480 108.305 19.350 ;
        RECT 108.505 32.680 109.895 39.170 ;
        RECT 110.525 38.660 111.025 38.830 ;
        RECT 110.295 33.405 110.465 38.445 ;
        RECT 111.085 33.405 111.255 38.445 ;
        RECT 110.525 33.020 111.025 33.190 ;
        RECT 111.655 32.680 111.825 39.170 ;
        RECT 112.455 38.660 112.955 38.830 ;
        RECT 112.225 33.405 112.395 38.445 ;
        RECT 113.015 33.405 113.185 38.445 ;
        RECT 113.585 36.810 114.645 39.170 ;
        RECT 115.625 37.420 116.055 39.820 ;
        RECT 116.685 39.310 117.185 39.480 ;
        RECT 116.455 38.100 116.625 39.140 ;
        RECT 117.245 38.100 117.415 39.140 ;
        RECT 116.685 37.760 117.185 37.930 ;
        RECT 117.815 37.420 119.535 39.820 ;
        RECT 126.835 39.840 130.745 40.110 ;
        RECT 115.625 37.200 119.535 37.420 ;
        RECT 119.715 39.190 125.855 39.680 ;
        RECT 113.585 36.090 119.505 36.810 ;
        RECT 112.455 33.020 112.955 33.190 ;
        RECT 113.585 32.680 115.905 36.090 ;
        RECT 116.535 35.580 117.035 35.750 ;
        RECT 116.305 33.325 116.475 35.365 ;
        RECT 117.095 33.325 117.265 35.365 ;
        RECT 116.535 32.940 117.035 33.110 ;
        RECT 108.505 32.600 115.905 32.680 ;
        RECT 117.665 32.600 119.505 36.090 ;
        RECT 108.505 30.530 119.505 32.600 ;
        RECT 108.505 19.390 109.145 30.530 ;
        RECT 109.545 20.120 109.715 30.160 ;
        RECT 110.835 20.120 111.005 30.160 ;
        RECT 109.775 19.735 110.775 19.905 ;
        RECT 111.405 19.390 111.575 30.530 ;
        RECT 111.975 20.120 112.145 30.160 ;
        RECT 117.265 20.120 117.435 30.160 ;
        RECT 112.205 19.735 117.205 19.905 ;
        RECT 117.835 19.390 119.505 30.530 ;
        RECT 108.505 18.520 119.505 19.390 ;
        RECT 119.715 32.700 121.105 39.190 ;
        RECT 121.735 38.680 122.235 38.850 ;
        RECT 121.505 33.425 121.675 38.465 ;
        RECT 122.295 33.425 122.465 38.465 ;
        RECT 121.735 33.040 122.235 33.210 ;
        RECT 122.865 32.700 123.035 39.190 ;
        RECT 123.665 38.680 124.165 38.850 ;
        RECT 123.435 33.425 123.605 38.465 ;
        RECT 124.225 33.425 124.395 38.465 ;
        RECT 124.795 36.830 125.855 39.190 ;
        RECT 126.835 37.440 127.265 39.840 ;
        RECT 127.895 39.330 128.395 39.500 ;
        RECT 127.665 38.120 127.835 39.160 ;
        RECT 128.455 38.120 128.625 39.160 ;
        RECT 127.895 37.780 128.395 37.950 ;
        RECT 129.025 37.440 130.745 39.840 ;
        RECT 126.835 37.220 130.745 37.440 ;
        RECT 124.795 36.110 130.715 36.830 ;
        RECT 123.665 33.040 124.165 33.210 ;
        RECT 124.795 32.700 127.115 36.110 ;
        RECT 127.745 35.600 128.245 35.770 ;
        RECT 127.515 33.345 127.685 35.385 ;
        RECT 128.305 33.345 128.475 35.385 ;
        RECT 127.745 32.960 128.245 33.130 ;
        RECT 119.715 32.620 127.115 32.700 ;
        RECT 128.875 32.620 130.715 36.110 ;
        RECT 119.715 31.140 130.715 32.620 ;
        RECT 119.715 30.550 139.465 31.140 ;
        RECT 119.715 19.410 120.355 30.550 ;
        RECT 120.755 20.140 120.925 30.180 ;
        RECT 122.045 20.140 122.215 30.180 ;
        RECT 120.985 19.755 121.985 19.925 ;
        RECT 122.615 19.410 122.785 30.550 ;
        RECT 129.045 30.520 139.465 30.550 ;
        RECT 123.185 20.140 123.355 30.180 ;
        RECT 128.475 20.140 128.645 30.180 ;
        RECT 123.415 19.755 128.415 19.925 ;
        RECT 129.045 19.410 132.075 30.520 ;
        RECT 132.475 20.110 132.645 30.150 ;
        RECT 137.765 20.110 137.935 30.150 ;
        RECT 132.705 19.725 137.705 19.895 ;
        RECT 119.715 19.380 132.075 19.410 ;
        RECT 138.335 19.380 139.465 30.520 ;
        RECT 119.715 18.540 139.465 19.380 ;
        RECT 131.925 18.520 139.465 18.540 ;
      LAYER met1 ;
        RECT 135.340 223.880 136.790 225.180 ;
        RECT 59.700 204.950 60.020 205.010 ;
        RECT 75.800 204.950 76.120 205.010 ;
        RECT 59.700 204.810 76.120 204.950 ;
        RECT 59.700 204.750 60.020 204.810 ;
        RECT 75.800 204.750 76.120 204.810 ;
        RECT 22.830 203.790 113.450 204.270 ;
        RECT 63.315 203.590 63.605 203.635 ;
        RECT 64.775 203.590 65.065 203.635 ;
        RECT 63.315 203.450 65.065 203.590 ;
        RECT 63.315 203.405 63.605 203.450 ;
        RECT 64.775 203.405 65.065 203.450 ;
        RECT 65.680 203.590 66.000 203.650 ;
        RECT 68.440 203.590 68.760 203.650 ;
        RECT 65.680 203.450 68.760 203.590 ;
        RECT 65.680 203.390 66.000 203.450 ;
        RECT 68.440 203.390 68.760 203.450 ;
        RECT 72.120 203.590 72.440 203.650 ;
        RECT 80.860 203.590 81.180 203.650 ;
        RECT 72.120 203.450 81.180 203.590 ;
        RECT 72.120 203.390 72.440 203.450 ;
        RECT 80.860 203.390 81.180 203.450 ;
        RECT 64.315 203.250 64.605 203.295 ;
        RECT 67.980 203.250 68.300 203.310 ;
        RECT 70.280 203.250 70.600 203.310 ;
        RECT 64.315 203.110 68.300 203.250 ;
        RECT 64.315 203.065 64.605 203.110 ;
        RECT 67.980 203.050 68.300 203.110 ;
        RECT 68.530 203.110 73.270 203.250 ;
        RECT 59.700 202.710 60.020 202.970 ;
        RECT 61.095 202.910 61.385 202.955 ;
        RECT 61.095 202.770 62.690 202.910 ;
        RECT 61.095 202.725 61.385 202.770 ;
        RECT 58.780 202.230 59.100 202.290 ;
        RECT 62.550 202.275 62.690 202.770 ;
        RECT 65.680 202.710 66.000 202.970 ;
        RECT 66.140 202.710 66.460 202.970 ;
        RECT 66.615 202.910 66.905 202.955 ;
        RECT 68.530 202.910 68.670 203.110 ;
        RECT 70.280 203.050 70.600 203.110 ;
        RECT 66.615 202.770 68.670 202.910 ;
        RECT 66.615 202.725 66.905 202.770 ;
        RECT 68.900 202.710 69.220 202.970 ;
        RECT 73.130 202.955 73.270 203.110 ;
        RECT 96.130 203.110 99.030 203.250 ;
        RECT 70.755 202.910 71.045 202.955 ;
        RECT 71.215 202.910 71.505 202.955 ;
        RECT 70.755 202.770 71.505 202.910 ;
        RECT 70.755 202.725 71.045 202.770 ;
        RECT 71.215 202.725 71.505 202.770 ;
        RECT 71.675 202.910 71.965 202.955 ;
        RECT 71.675 202.770 72.350 202.910 ;
        RECT 71.675 202.725 71.965 202.770 ;
        RECT 67.060 202.570 67.380 202.630 ;
        RECT 70.830 202.570 70.970 202.725 ;
        RECT 67.060 202.430 70.970 202.570 ;
        RECT 67.060 202.370 67.380 202.430 ;
        RECT 59.255 202.230 59.545 202.275 ;
        RECT 58.780 202.090 59.545 202.230 ;
        RECT 58.780 202.030 59.100 202.090 ;
        RECT 59.255 202.045 59.545 202.090 ;
        RECT 62.475 202.045 62.765 202.275 ;
        RECT 66.140 202.230 66.460 202.290 ;
        RECT 71.675 202.230 71.965 202.275 ;
        RECT 66.140 202.090 71.965 202.230 ;
        RECT 66.140 202.030 66.460 202.090 ;
        RECT 71.675 202.045 71.965 202.090 ;
        RECT 72.210 202.230 72.350 202.770 ;
        RECT 73.055 202.725 73.345 202.955 ;
        RECT 75.800 202.910 76.120 202.970 ;
        RECT 96.130 202.955 96.270 203.110 ;
        RECT 77.195 202.910 77.485 202.955 ;
        RECT 75.800 202.770 77.485 202.910 ;
        RECT 75.800 202.710 76.120 202.770 ;
        RECT 77.195 202.725 77.485 202.770 ;
        RECT 77.655 202.725 77.945 202.955 ;
        RECT 96.055 202.725 96.345 202.955 ;
        RECT 96.960 202.910 97.280 202.970 ;
        RECT 98.890 202.955 99.030 203.110 ;
        RECT 97.435 202.910 97.725 202.955 ;
        RECT 96.960 202.770 97.725 202.910 ;
        RECT 75.340 202.570 75.660 202.630 ;
        RECT 77.730 202.570 77.870 202.725 ;
        RECT 96.960 202.710 97.280 202.770 ;
        RECT 97.435 202.725 97.725 202.770 ;
        RECT 98.815 202.910 99.105 202.955 ;
        RECT 101.560 202.910 101.880 202.970 ;
        RECT 98.815 202.770 101.880 202.910 ;
        RECT 98.815 202.725 99.105 202.770 ;
        RECT 101.560 202.710 101.880 202.770 ;
        RECT 75.340 202.430 77.870 202.570 ;
        RECT 102.955 202.570 103.245 202.615 ;
        RECT 104.320 202.570 104.640 202.630 ;
        RECT 102.955 202.430 104.640 202.570 ;
        RECT 75.340 202.370 75.660 202.430 ;
        RECT 102.955 202.385 103.245 202.430 ;
        RECT 104.320 202.370 104.640 202.430 ;
        RECT 79.940 202.230 80.260 202.290 ;
        RECT 72.210 202.090 80.260 202.230 ;
        RECT 56.020 201.890 56.340 201.950 ;
        RECT 60.175 201.890 60.465 201.935 ;
        RECT 56.020 201.750 60.465 201.890 ;
        RECT 56.020 201.690 56.340 201.750 ;
        RECT 60.175 201.705 60.465 201.750 ;
        RECT 63.395 201.890 63.685 201.935 ;
        RECT 66.230 201.890 66.370 202.030 ;
        RECT 63.395 201.750 66.370 201.890 ;
        RECT 63.395 201.705 63.685 201.750 ;
        RECT 67.980 201.690 68.300 201.950 ;
        RECT 68.440 201.890 68.760 201.950 ;
        RECT 69.820 201.890 70.140 201.950 ;
        RECT 70.295 201.890 70.585 201.935 ;
        RECT 72.210 201.890 72.350 202.090 ;
        RECT 79.940 202.030 80.260 202.090 ;
        RECT 68.440 201.750 72.350 201.890 ;
        RECT 74.880 201.890 75.200 201.950 ;
        RECT 75.355 201.890 75.645 201.935 ;
        RECT 74.880 201.750 75.645 201.890 ;
        RECT 68.440 201.690 68.760 201.750 ;
        RECT 69.820 201.690 70.140 201.750 ;
        RECT 70.295 201.705 70.585 201.750 ;
        RECT 74.880 201.690 75.200 201.750 ;
        RECT 75.355 201.705 75.645 201.750 ;
        RECT 76.720 201.690 77.040 201.950 ;
        RECT 78.575 201.890 78.865 201.935 ;
        RECT 79.480 201.890 79.800 201.950 ;
        RECT 78.575 201.750 79.800 201.890 ;
        RECT 78.575 201.705 78.865 201.750 ;
        RECT 79.480 201.690 79.800 201.750 ;
        RECT 95.580 201.690 95.900 201.950 ;
        RECT 98.340 201.690 98.660 201.950 ;
        RECT 99.260 201.690 99.580 201.950 ;
        RECT 101.100 201.690 101.420 201.950 ;
        RECT 105.715 201.890 106.005 201.935 ;
        RECT 106.620 201.890 106.940 201.950 ;
        RECT 105.715 201.750 106.940 201.890 ;
        RECT 105.715 201.705 106.005 201.750 ;
        RECT 106.620 201.690 106.940 201.750 ;
        RECT 22.830 201.070 113.450 201.550 ;
        RECT 67.520 200.870 67.840 200.930 ;
        RECT 70.295 200.870 70.585 200.915 ;
        RECT 67.520 200.730 70.585 200.870 ;
        RECT 67.520 200.670 67.840 200.730 ;
        RECT 70.295 200.685 70.585 200.730 ;
        RECT 75.800 200.870 76.120 200.930 ;
        RECT 75.800 200.730 88.910 200.870 ;
        RECT 75.800 200.670 76.120 200.730 ;
        RECT 53.225 200.530 53.515 200.575 ;
        RECT 55.115 200.530 55.405 200.575 ;
        RECT 58.235 200.530 58.525 200.575 ;
        RECT 53.225 200.390 58.525 200.530 ;
        RECT 53.225 200.345 53.515 200.390 ;
        RECT 55.115 200.345 55.405 200.390 ;
        RECT 58.235 200.345 58.525 200.390 ;
        RECT 63.855 200.345 64.145 200.575 ;
        RECT 73.615 200.530 73.905 200.575 ;
        RECT 76.735 200.530 77.025 200.575 ;
        RECT 78.625 200.530 78.915 200.575 ;
        RECT 73.615 200.390 78.915 200.530 ;
        RECT 73.615 200.345 73.905 200.390 ;
        RECT 76.735 200.345 77.025 200.390 ;
        RECT 78.625 200.345 78.915 200.390 ;
        RECT 53.735 200.190 54.025 200.235 ;
        RECT 63.930 200.190 64.070 200.345 ;
        RECT 79.480 200.330 79.800 200.590 ;
        RECT 80.860 200.530 81.180 200.590 ;
        RECT 80.860 200.390 86.150 200.530 ;
        RECT 80.860 200.330 81.180 200.390 ;
        RECT 53.735 200.050 64.070 200.190 ;
        RECT 53.735 200.005 54.025 200.050 ;
        RECT 66.140 199.990 66.460 200.250 ;
        RECT 70.755 200.005 71.045 200.235 ;
        RECT 78.115 200.190 78.405 200.235 ;
        RECT 79.570 200.190 79.710 200.330 ;
        RECT 78.115 200.050 79.710 200.190 ;
        RECT 80.400 200.190 80.720 200.250 ;
        RECT 81.335 200.190 81.625 200.235 ;
        RECT 80.400 200.050 81.625 200.190 ;
        RECT 78.115 200.005 78.405 200.050 ;
        RECT 52.340 199.650 52.660 199.910 ;
        RECT 52.820 199.850 53.110 199.895 ;
        RECT 54.655 199.850 54.945 199.895 ;
        RECT 58.235 199.850 58.525 199.895 ;
        RECT 52.820 199.710 58.525 199.850 ;
        RECT 52.820 199.665 53.110 199.710 ;
        RECT 54.655 199.665 54.945 199.710 ;
        RECT 58.235 199.665 58.525 199.710 ;
        RECT 59.240 199.870 59.560 199.910 ;
        RECT 59.240 199.650 59.605 199.870 ;
        RECT 65.680 199.650 66.000 199.910 ;
        RECT 67.060 199.650 67.380 199.910 ;
        RECT 68.440 199.850 68.760 199.910 ;
        RECT 69.360 199.895 69.680 199.910 ;
        RECT 68.915 199.850 69.205 199.895 ;
        RECT 68.440 199.710 69.205 199.850 ;
        RECT 68.440 199.650 68.760 199.710 ;
        RECT 68.915 199.665 69.205 199.710 ;
        RECT 69.360 199.850 69.790 199.895 ;
        RECT 70.830 199.850 70.970 200.005 ;
        RECT 80.400 199.990 80.720 200.050 ;
        RECT 81.335 200.005 81.625 200.050 ;
        RECT 69.360 199.710 70.970 199.850 ;
        RECT 69.360 199.665 69.790 199.710 ;
        RECT 69.360 199.650 69.680 199.665 ;
        RECT 59.315 199.555 59.605 199.650 ;
        RECT 72.535 199.555 72.825 199.870 ;
        RECT 73.615 199.850 73.905 199.895 ;
        RECT 77.195 199.850 77.485 199.895 ;
        RECT 79.030 199.850 79.320 199.895 ;
        RECT 73.615 199.710 79.320 199.850 ;
        RECT 73.615 199.665 73.905 199.710 ;
        RECT 77.195 199.665 77.485 199.710 ;
        RECT 79.030 199.665 79.320 199.710 ;
        RECT 79.495 199.665 79.785 199.895 ;
        RECT 79.940 199.850 80.260 199.910 ;
        RECT 86.010 199.895 86.150 200.390 ;
        RECT 88.770 200.190 88.910 200.730 ;
        RECT 96.960 200.670 97.280 200.930 ;
        RECT 97.435 200.870 97.725 200.915 ;
        RECT 98.800 200.870 99.120 200.930 ;
        RECT 102.940 200.870 103.260 200.930 ;
        RECT 97.435 200.730 103.260 200.870 ;
        RECT 97.435 200.685 97.725 200.730 ;
        RECT 98.800 200.670 99.120 200.730 ;
        RECT 102.940 200.670 103.260 200.730 ;
        RECT 100.295 200.530 100.585 200.575 ;
        RECT 103.415 200.530 103.705 200.575 ;
        RECT 105.305 200.530 105.595 200.575 ;
        RECT 100.295 200.390 105.595 200.530 ;
        RECT 100.295 200.345 100.585 200.390 ;
        RECT 103.415 200.345 103.705 200.390 ;
        RECT 105.305 200.345 105.595 200.390 ;
        RECT 107.095 200.345 107.385 200.575 ;
        RECT 101.560 200.190 101.880 200.250 ;
        RECT 88.770 200.050 101.880 200.190 ;
        RECT 88.770 199.895 88.910 200.050 ;
        RECT 101.560 199.990 101.880 200.050 ;
        RECT 104.795 200.190 105.085 200.235 ;
        RECT 107.170 200.190 107.310 200.345 ;
        RECT 104.795 200.050 107.310 200.190 ;
        RECT 104.795 200.005 105.085 200.050 ;
        RECT 81.795 199.850 82.085 199.895 ;
        RECT 79.940 199.710 82.085 199.850 ;
        RECT 56.015 199.510 56.665 199.555 ;
        RECT 59.315 199.510 59.905 199.555 ;
        RECT 56.015 199.370 59.905 199.510 ;
        RECT 56.015 199.325 56.665 199.370 ;
        RECT 59.615 199.325 59.905 199.370 ;
        RECT 72.235 199.510 72.825 199.555 ;
        RECT 75.475 199.510 76.125 199.555 ;
        RECT 76.720 199.510 77.040 199.570 ;
        RECT 72.235 199.370 77.040 199.510 ;
        RECT 79.570 199.510 79.710 199.665 ;
        RECT 79.940 199.650 80.260 199.710 ;
        RECT 81.795 199.665 82.085 199.710 ;
        RECT 85.935 199.665 86.225 199.895 ;
        RECT 88.695 199.665 88.985 199.895 ;
        RECT 90.535 199.850 90.825 199.895 ;
        RECT 90.980 199.850 91.300 199.910 ;
        RECT 90.535 199.710 91.300 199.850 ;
        RECT 90.535 199.665 90.825 199.710 ;
        RECT 90.980 199.650 91.300 199.710 ;
        RECT 94.215 199.850 94.505 199.895 ;
        RECT 97.420 199.850 97.740 199.910 ;
        RECT 94.215 199.710 97.740 199.850 ;
        RECT 94.215 199.665 94.505 199.710 ;
        RECT 97.420 199.650 97.740 199.710 ;
        RECT 87.300 199.510 87.620 199.570 ;
        RECT 99.215 199.555 99.505 199.870 ;
        RECT 100.295 199.850 100.585 199.895 ;
        RECT 103.875 199.850 104.165 199.895 ;
        RECT 105.710 199.850 106.000 199.895 ;
        RECT 100.295 199.710 106.000 199.850 ;
        RECT 100.295 199.665 100.585 199.710 ;
        RECT 103.875 199.665 104.165 199.710 ;
        RECT 105.710 199.665 106.000 199.710 ;
        RECT 106.175 199.665 106.465 199.895 ;
        RECT 106.620 199.850 106.940 199.910 ;
        RECT 108.015 199.850 108.305 199.895 ;
        RECT 106.620 199.710 108.305 199.850 ;
        RECT 79.570 199.370 87.620 199.510 ;
        RECT 72.235 199.325 72.525 199.370 ;
        RECT 75.475 199.325 76.125 199.370 ;
        RECT 76.720 199.310 77.040 199.370 ;
        RECT 87.300 199.310 87.620 199.370 ;
        RECT 98.915 199.510 99.505 199.555 ;
        RECT 101.100 199.510 101.420 199.570 ;
        RECT 102.155 199.510 102.805 199.555 ;
        RECT 98.915 199.370 102.805 199.510 ;
        RECT 98.915 199.325 99.205 199.370 ;
        RECT 101.100 199.310 101.420 199.370 ;
        RECT 102.155 199.325 102.805 199.370 ;
        RECT 105.240 199.510 105.560 199.570 ;
        RECT 106.250 199.510 106.390 199.665 ;
        RECT 106.620 199.650 106.940 199.710 ;
        RECT 108.015 199.665 108.305 199.710 ;
        RECT 105.240 199.370 106.390 199.510 ;
        RECT 105.240 199.310 105.560 199.370 ;
        RECT 61.095 199.170 61.385 199.215 ;
        RECT 65.220 199.170 65.540 199.230 ;
        RECT 61.095 199.030 65.540 199.170 ;
        RECT 61.095 198.985 61.385 199.030 ;
        RECT 65.220 198.970 65.540 199.030 ;
        RECT 68.455 199.170 68.745 199.215 ;
        RECT 70.740 199.170 71.060 199.230 ;
        RECT 68.455 199.030 71.060 199.170 ;
        RECT 68.455 198.985 68.745 199.030 ;
        RECT 70.740 198.970 71.060 199.030 ;
        RECT 79.940 198.970 80.260 199.230 ;
        RECT 86.380 198.970 86.700 199.230 ;
        RECT 89.155 199.170 89.445 199.215 ;
        RECT 89.600 199.170 89.920 199.230 ;
        RECT 89.155 199.030 89.920 199.170 ;
        RECT 89.155 198.985 89.445 199.030 ;
        RECT 89.600 198.970 89.920 199.030 ;
        RECT 93.295 199.170 93.585 199.215 ;
        RECT 99.720 199.170 100.040 199.230 ;
        RECT 93.295 199.030 100.040 199.170 ;
        RECT 93.295 198.985 93.585 199.030 ;
        RECT 99.720 198.970 100.040 199.030 ;
        RECT 22.830 198.350 113.450 198.830 ;
        RECT 65.680 198.150 66.000 198.210 ;
        RECT 68.455 198.150 68.745 198.195 ;
        RECT 65.680 198.010 68.745 198.150 ;
        RECT 65.680 197.950 66.000 198.010 ;
        RECT 68.455 197.965 68.745 198.010 ;
        RECT 69.375 198.150 69.665 198.195 ;
        RECT 69.820 198.150 70.140 198.210 ;
        RECT 69.375 198.010 70.140 198.150 ;
        RECT 69.375 197.965 69.665 198.010 ;
        RECT 69.820 197.950 70.140 198.010 ;
        RECT 75.340 197.950 75.660 198.210 ;
        RECT 80.400 198.150 80.720 198.210 ;
        RECT 78.650 198.010 80.720 198.150 ;
        RECT 56.020 197.610 56.340 197.870 ;
        RECT 58.780 197.855 59.100 197.870 ;
        RECT 58.315 197.810 59.100 197.855 ;
        RECT 61.915 197.810 62.205 197.855 ;
        RECT 58.315 197.670 62.205 197.810 ;
        RECT 58.315 197.625 59.100 197.670 ;
        RECT 58.780 197.610 59.100 197.625 ;
        RECT 61.615 197.625 62.205 197.670 ;
        RECT 67.980 197.810 68.300 197.870 ;
        RECT 76.115 197.810 76.405 197.855 ;
        RECT 67.980 197.670 76.405 197.810 ;
        RECT 46.360 197.470 46.680 197.530 ;
        RECT 50.055 197.470 50.345 197.515 ;
        RECT 46.360 197.330 50.345 197.470 ;
        RECT 46.360 197.270 46.680 197.330 ;
        RECT 50.055 197.285 50.345 197.330 ;
        RECT 52.340 197.470 52.660 197.530 ;
        RECT 54.655 197.470 54.945 197.515 ;
        RECT 52.340 197.330 54.945 197.470 ;
        RECT 52.340 197.270 52.660 197.330 ;
        RECT 54.655 197.285 54.945 197.330 ;
        RECT 55.120 197.470 55.410 197.515 ;
        RECT 56.955 197.470 57.245 197.515 ;
        RECT 60.535 197.470 60.825 197.515 ;
        RECT 55.120 197.330 60.825 197.470 ;
        RECT 55.120 197.285 55.410 197.330 ;
        RECT 56.955 197.285 57.245 197.330 ;
        RECT 60.535 197.285 60.825 197.330 ;
        RECT 61.615 197.310 61.905 197.625 ;
        RECT 67.980 197.610 68.300 197.670 ;
        RECT 76.115 197.625 76.405 197.670 ;
        RECT 77.195 197.810 77.485 197.855 ;
        RECT 78.650 197.810 78.790 198.010 ;
        RECT 80.400 197.950 80.720 198.010 ;
        RECT 104.320 197.950 104.640 198.210 ;
        RECT 77.195 197.670 78.790 197.810 ;
        RECT 79.135 197.810 79.425 197.855 ;
        RECT 81.780 197.810 82.100 197.870 ;
        RECT 82.375 197.810 83.025 197.855 ;
        RECT 79.135 197.670 83.025 197.810 ;
        RECT 77.195 197.625 77.485 197.670 ;
        RECT 79.135 197.625 79.725 197.670 ;
        RECT 54.730 197.130 54.870 197.285 ;
        RECT 65.220 197.270 65.540 197.530 ;
        RECT 70.295 197.470 70.585 197.515 ;
        RECT 70.740 197.470 71.060 197.530 ;
        RECT 70.295 197.330 71.060 197.470 ;
        RECT 70.295 197.285 70.585 197.330 ;
        RECT 70.740 197.270 71.060 197.330 ;
        RECT 79.435 197.310 79.725 197.625 ;
        RECT 81.780 197.610 82.100 197.670 ;
        RECT 82.375 197.625 83.025 197.670 ;
        RECT 85.015 197.810 85.305 197.855 ;
        RECT 86.380 197.810 86.700 197.870 ;
        RECT 95.580 197.855 95.900 197.870 ;
        RECT 85.015 197.670 86.700 197.810 ;
        RECT 85.015 197.625 85.305 197.670 ;
        RECT 86.380 197.610 86.700 197.670 ;
        RECT 92.475 197.810 92.765 197.855 ;
        RECT 95.580 197.810 96.365 197.855 ;
        RECT 92.475 197.670 96.365 197.810 ;
        RECT 92.475 197.625 93.065 197.670 ;
        RECT 80.515 197.470 80.805 197.515 ;
        RECT 84.095 197.470 84.385 197.515 ;
        RECT 85.930 197.470 86.220 197.515 ;
        RECT 80.515 197.330 86.220 197.470 ;
        RECT 80.515 197.285 80.805 197.330 ;
        RECT 84.095 197.285 84.385 197.330 ;
        RECT 85.930 197.285 86.220 197.330 ;
        RECT 92.775 197.310 93.065 197.625 ;
        RECT 95.580 197.625 96.365 197.670 ;
        RECT 95.580 197.610 95.900 197.625 ;
        RECT 98.340 197.610 98.660 197.870 ;
        RECT 99.720 197.810 100.040 197.870 ;
        RECT 102.495 197.810 102.785 197.855 ;
        RECT 99.720 197.670 102.785 197.810 ;
        RECT 99.720 197.610 100.040 197.670 ;
        RECT 102.495 197.625 102.785 197.670 ;
        RECT 93.855 197.470 94.145 197.515 ;
        RECT 97.435 197.470 97.725 197.515 ;
        RECT 99.270 197.470 99.560 197.515 ;
        RECT 93.855 197.330 99.560 197.470 ;
        RECT 93.855 197.285 94.145 197.330 ;
        RECT 97.435 197.285 97.725 197.330 ;
        RECT 99.270 197.285 99.560 197.330 ;
        RECT 100.640 197.470 100.960 197.530 ;
        RECT 104.795 197.470 105.085 197.515 ;
        RECT 100.640 197.330 105.085 197.470 ;
        RECT 100.640 197.270 100.960 197.330 ;
        RECT 104.795 197.285 105.085 197.330 ;
        RECT 108.015 197.470 108.305 197.515 ;
        RECT 109.395 197.470 109.685 197.515 ;
        RECT 108.015 197.330 109.685 197.470 ;
        RECT 108.015 197.285 108.305 197.330 ;
        RECT 109.395 197.285 109.685 197.330 ;
        RECT 110.775 197.285 111.065 197.515 ;
        RECT 61.080 197.130 61.400 197.190 ;
        RECT 54.730 196.990 61.400 197.130 ;
        RECT 61.080 196.930 61.400 196.990 ;
        RECT 64.775 197.130 65.065 197.175 ;
        RECT 67.060 197.130 67.380 197.190 ;
        RECT 67.980 197.130 68.300 197.190 ;
        RECT 64.775 196.990 68.300 197.130 ;
        RECT 64.775 196.945 65.065 196.990 ;
        RECT 67.060 196.930 67.380 196.990 ;
        RECT 67.980 196.930 68.300 196.990 ;
        RECT 68.440 197.130 68.760 197.190 ;
        RECT 71.215 197.130 71.505 197.175 ;
        RECT 77.655 197.130 77.945 197.175 ;
        RECT 68.440 196.990 77.945 197.130 ;
        RECT 68.440 196.930 68.760 196.990 ;
        RECT 71.215 196.945 71.505 196.990 ;
        RECT 77.655 196.945 77.945 196.990 ;
        RECT 86.395 197.130 86.685 197.175 ;
        RECT 87.300 197.130 87.620 197.190 ;
        RECT 86.395 196.990 87.620 197.130 ;
        RECT 86.395 196.945 86.685 196.990 ;
        RECT 87.300 196.930 87.620 196.990 ;
        RECT 87.775 197.130 88.065 197.175 ;
        RECT 89.140 197.130 89.460 197.190 ;
        RECT 87.775 196.990 89.460 197.130 ;
        RECT 87.775 196.945 88.065 196.990 ;
        RECT 89.140 196.930 89.460 196.990 ;
        RECT 99.720 196.930 100.040 197.190 ;
        RECT 101.100 196.930 101.420 197.190 ;
        RECT 102.035 197.130 102.325 197.175 ;
        RECT 102.940 197.130 103.260 197.190 ;
        RECT 102.035 196.990 103.260 197.130 ;
        RECT 102.035 196.945 102.325 196.990 ;
        RECT 102.940 196.930 103.260 196.990 ;
        RECT 104.320 197.130 104.640 197.190 ;
        RECT 110.850 197.130 110.990 197.285 ;
        RECT 104.320 196.990 110.990 197.130 ;
        RECT 104.320 196.930 104.640 196.990 ;
        RECT 55.525 196.790 55.815 196.835 ;
        RECT 57.415 196.790 57.705 196.835 ;
        RECT 60.535 196.790 60.825 196.835 ;
        RECT 55.525 196.650 60.825 196.790 ;
        RECT 55.525 196.605 55.815 196.650 ;
        RECT 57.415 196.605 57.705 196.650 ;
        RECT 60.535 196.605 60.825 196.650 ;
        RECT 80.515 196.790 80.805 196.835 ;
        RECT 83.635 196.790 83.925 196.835 ;
        RECT 85.525 196.790 85.815 196.835 ;
        RECT 80.515 196.650 85.815 196.790 ;
        RECT 80.515 196.605 80.805 196.650 ;
        RECT 83.635 196.605 83.925 196.650 ;
        RECT 85.525 196.605 85.815 196.650 ;
        RECT 93.855 196.790 94.145 196.835 ;
        RECT 96.975 196.790 97.265 196.835 ;
        RECT 98.865 196.790 99.155 196.835 ;
        RECT 93.855 196.650 99.155 196.790 ;
        RECT 93.855 196.605 94.145 196.650 ;
        RECT 96.975 196.605 97.265 196.650 ;
        RECT 98.865 196.605 99.155 196.650 ;
        RECT 46.820 196.450 47.140 196.510 ;
        RECT 49.135 196.450 49.425 196.495 ;
        RECT 46.820 196.310 49.425 196.450 ;
        RECT 46.820 196.250 47.140 196.310 ;
        RECT 49.135 196.265 49.425 196.310 ;
        RECT 73.040 196.450 73.360 196.510 ;
        RECT 73.975 196.450 74.265 196.495 ;
        RECT 73.040 196.310 74.265 196.450 ;
        RECT 73.040 196.250 73.360 196.310 ;
        RECT 73.975 196.265 74.265 196.310 ;
        RECT 76.275 196.450 76.565 196.495 ;
        RECT 76.720 196.450 77.040 196.510 ;
        RECT 76.275 196.310 77.040 196.450 ;
        RECT 76.275 196.265 76.565 196.310 ;
        RECT 76.720 196.250 77.040 196.310 ;
        RECT 90.520 196.250 90.840 196.510 ;
        RECT 90.980 196.250 91.300 196.510 ;
        RECT 101.560 196.450 101.880 196.510 ;
        RECT 105.700 196.450 106.020 196.510 ;
        RECT 101.560 196.310 106.020 196.450 ;
        RECT 101.560 196.250 101.880 196.310 ;
        RECT 105.700 196.250 106.020 196.310 ;
        RECT 107.080 196.450 107.400 196.510 ;
        RECT 108.475 196.450 108.765 196.495 ;
        RECT 107.080 196.310 108.765 196.450 ;
        RECT 107.080 196.250 107.400 196.310 ;
        RECT 108.475 196.265 108.765 196.310 ;
        RECT 109.840 196.250 110.160 196.510 ;
        RECT 22.830 195.630 113.450 196.110 ;
        RECT 46.360 195.230 46.680 195.490 ;
        RECT 59.240 195.230 59.560 195.490 ;
        RECT 64.775 195.430 65.065 195.475 ;
        RECT 65.220 195.430 65.540 195.490 ;
        RECT 64.775 195.290 65.540 195.430 ;
        RECT 64.775 195.245 65.065 195.290 ;
        RECT 65.220 195.230 65.540 195.290 ;
        RECT 65.695 195.430 65.985 195.475 ;
        RECT 68.900 195.430 69.220 195.490 ;
        RECT 65.695 195.290 69.220 195.430 ;
        RECT 65.695 195.245 65.985 195.290 ;
        RECT 68.900 195.230 69.220 195.290 ;
        RECT 70.740 195.230 71.060 195.490 ;
        RECT 80.400 195.230 80.720 195.490 ;
        RECT 81.780 195.230 82.100 195.490 ;
        RECT 98.800 195.430 99.120 195.490 ;
        RECT 105.240 195.430 105.560 195.490 ;
        RECT 87.390 195.290 99.120 195.430 ;
        RECT 35.320 194.890 35.640 195.150 ;
        RECT 66.615 195.090 66.905 195.135 ;
        RECT 69.820 195.090 70.140 195.150 ;
        RECT 66.615 194.950 70.140 195.090 ;
        RECT 66.615 194.905 66.905 194.950 ;
        RECT 69.820 194.890 70.140 194.950 ;
        RECT 73.615 195.090 73.905 195.135 ;
        RECT 76.735 195.090 77.025 195.135 ;
        RECT 78.625 195.090 78.915 195.135 ;
        RECT 79.940 195.090 80.260 195.150 ;
        RECT 73.615 194.950 78.915 195.090 ;
        RECT 73.615 194.905 73.905 194.950 ;
        RECT 76.735 194.905 77.025 194.950 ;
        RECT 78.625 194.905 78.915 194.950 ;
        RECT 79.110 194.950 80.260 195.090 ;
        RECT 31.195 194.750 31.485 194.795 ;
        RECT 36.240 194.750 36.560 194.810 ;
        RECT 31.195 194.610 36.560 194.750 ;
        RECT 31.195 194.565 31.485 194.610 ;
        RECT 36.240 194.550 36.560 194.610 ;
        RECT 50.055 194.750 50.345 194.795 ;
        RECT 53.260 194.750 53.580 194.810 ;
        RECT 50.055 194.610 53.580 194.750 ;
        RECT 50.055 194.565 50.345 194.610 ;
        RECT 53.260 194.550 53.580 194.610 ;
        RECT 68.440 194.750 68.760 194.810 ;
        RECT 69.375 194.750 69.665 194.795 ;
        RECT 68.440 194.610 69.665 194.750 ;
        RECT 68.440 194.550 68.760 194.610 ;
        RECT 69.375 194.565 69.665 194.610 ;
        RECT 78.115 194.750 78.405 194.795 ;
        RECT 79.110 194.750 79.250 194.950 ;
        RECT 79.940 194.890 80.260 194.950 ;
        RECT 78.115 194.610 79.250 194.750 ;
        RECT 79.495 194.750 79.785 194.795 ;
        RECT 84.095 194.750 84.385 194.795 ;
        RECT 87.390 194.750 87.530 195.290 ;
        RECT 98.800 195.230 99.120 195.290 ;
        RECT 100.730 195.290 105.560 195.430 ;
        RECT 90.635 195.090 90.925 195.135 ;
        RECT 93.755 195.090 94.045 195.135 ;
        RECT 95.645 195.090 95.935 195.135 ;
        RECT 90.635 194.950 95.935 195.090 ;
        RECT 90.635 194.905 90.925 194.950 ;
        RECT 93.755 194.905 94.045 194.950 ;
        RECT 95.645 194.905 95.935 194.950 ;
        RECT 79.495 194.610 83.850 194.750 ;
        RECT 78.115 194.565 78.405 194.610 ;
        RECT 79.495 194.565 79.785 194.610 ;
        RECT 30.260 194.410 30.580 194.470 ;
        RECT 30.735 194.410 31.025 194.455 ;
        RECT 30.260 194.270 31.025 194.410 ;
        RECT 30.260 194.210 30.580 194.270 ;
        RECT 30.735 194.225 31.025 194.270 ;
        RECT 32.100 194.210 32.420 194.470 ;
        RECT 33.035 194.225 33.325 194.455 ;
        RECT 33.110 194.070 33.250 194.225 ;
        RECT 33.480 194.210 33.800 194.470 ;
        RECT 33.955 194.410 34.245 194.455 ;
        RECT 35.320 194.410 35.640 194.470 ;
        RECT 33.955 194.270 35.640 194.410 ;
        RECT 33.955 194.225 34.245 194.270 ;
        RECT 35.320 194.210 35.640 194.270 ;
        RECT 38.095 194.410 38.385 194.455 ;
        RECT 39.460 194.410 39.780 194.470 ;
        RECT 38.095 194.270 39.780 194.410 ;
        RECT 38.095 194.225 38.385 194.270 ;
        RECT 39.460 194.210 39.780 194.270 ;
        RECT 43.600 194.210 43.920 194.470 ;
        RECT 45.900 194.410 46.220 194.470 ;
        RECT 46.835 194.410 47.125 194.455 ;
        RECT 45.900 194.270 47.125 194.410 ;
        RECT 45.900 194.210 46.220 194.270 ;
        RECT 46.835 194.225 47.125 194.270 ;
        RECT 50.960 194.410 51.280 194.470 ;
        RECT 51.435 194.410 51.725 194.455 ;
        RECT 50.960 194.270 51.725 194.410 ;
        RECT 50.960 194.210 51.280 194.270 ;
        RECT 51.435 194.225 51.725 194.270 ;
        RECT 51.895 194.410 52.185 194.455 ;
        RECT 56.940 194.410 57.260 194.470 ;
        RECT 51.895 194.270 57.260 194.410 ;
        RECT 51.895 194.225 52.185 194.270 ;
        RECT 56.940 194.210 57.260 194.270 ;
        RECT 59.700 194.210 60.020 194.470 ;
        RECT 62.935 194.225 63.225 194.455 ;
        RECT 64.775 194.410 65.065 194.455 ;
        RECT 70.280 194.410 70.600 194.470 ;
        RECT 64.775 194.270 70.600 194.410 ;
        RECT 64.775 194.225 65.065 194.270 ;
        RECT 35.780 194.070 36.100 194.130 ;
        RECT 33.110 193.930 36.100 194.070 ;
        RECT 35.780 193.870 36.100 193.930 ;
        RECT 40.855 194.070 41.145 194.115 ;
        RECT 42.220 194.070 42.540 194.130 ;
        RECT 40.855 193.930 42.540 194.070 ;
        RECT 63.010 194.070 63.150 194.225 ;
        RECT 70.280 194.210 70.600 194.270 ;
        RECT 66.140 194.070 66.460 194.130 ;
        RECT 63.010 193.930 66.460 194.070 ;
        RECT 40.855 193.885 41.145 193.930 ;
        RECT 42.220 193.870 42.540 193.930 ;
        RECT 66.140 193.870 66.460 193.930 ;
        RECT 66.615 194.070 66.905 194.115 ;
        RECT 67.980 194.070 68.300 194.130 ;
        RECT 66.615 193.930 68.300 194.070 ;
        RECT 66.615 193.885 66.905 193.930 ;
        RECT 67.980 193.870 68.300 193.930 ;
        RECT 68.440 194.070 68.760 194.130 ;
        RECT 72.535 194.115 72.825 194.430 ;
        RECT 73.615 194.410 73.905 194.455 ;
        RECT 77.195 194.410 77.485 194.455 ;
        RECT 79.030 194.410 79.320 194.455 ;
        RECT 73.615 194.270 79.320 194.410 ;
        RECT 73.615 194.225 73.905 194.270 ;
        RECT 77.195 194.225 77.485 194.270 ;
        RECT 79.030 194.225 79.320 194.270 ;
        RECT 79.940 194.210 80.260 194.470 ;
        RECT 80.860 194.210 81.180 194.470 ;
        RECT 82.255 194.410 82.545 194.455 ;
        RECT 81.410 194.270 82.545 194.410 ;
        RECT 83.710 194.410 83.850 194.610 ;
        RECT 84.095 194.610 87.530 194.750 ;
        RECT 87.775 194.750 88.065 194.795 ;
        RECT 89.140 194.750 89.460 194.810 ;
        RECT 87.775 194.610 89.460 194.750 ;
        RECT 84.095 194.565 84.385 194.610 ;
        RECT 87.775 194.565 88.065 194.610 ;
        RECT 89.140 194.550 89.460 194.610 ;
        RECT 96.960 194.550 97.280 194.810 ;
        RECT 100.730 194.795 100.870 195.290 ;
        RECT 105.240 195.230 105.560 195.290 ;
        RECT 105.700 195.430 106.020 195.490 ;
        RECT 105.700 195.290 110.530 195.430 ;
        RECT 105.700 195.230 106.020 195.290 ;
        RECT 101.525 195.090 101.815 195.135 ;
        RECT 103.415 195.090 103.705 195.135 ;
        RECT 106.535 195.090 106.825 195.135 ;
        RECT 109.840 195.090 110.160 195.150 ;
        RECT 101.525 194.950 106.825 195.090 ;
        RECT 101.525 194.905 101.815 194.950 ;
        RECT 103.415 194.905 103.705 194.950 ;
        RECT 106.535 194.905 106.825 194.950 ;
        RECT 109.470 194.950 110.160 195.090 ;
        RECT 100.655 194.565 100.945 194.795 ;
        RECT 102.035 194.750 102.325 194.795 ;
        RECT 109.470 194.750 109.610 194.950 ;
        RECT 109.840 194.890 110.160 194.950 ;
        RECT 110.390 194.750 110.530 195.290 ;
        RECT 102.035 194.610 109.610 194.750 ;
        RECT 109.930 194.610 110.530 194.750 ;
        RECT 102.035 194.565 102.325 194.610 ;
        RECT 87.300 194.410 87.620 194.470 ;
        RECT 89.600 194.430 89.920 194.470 ;
        RECT 83.710 194.270 87.620 194.410 ;
        RECT 72.235 194.070 72.825 194.115 ;
        RECT 74.880 194.070 75.200 194.130 ;
        RECT 75.475 194.070 76.125 194.115 ;
        RECT 81.410 194.070 81.550 194.270 ;
        RECT 82.255 194.225 82.545 194.270 ;
        RECT 87.300 194.210 87.620 194.270 ;
        RECT 89.555 194.210 89.920 194.430 ;
        RECT 90.635 194.410 90.925 194.455 ;
        RECT 94.215 194.410 94.505 194.455 ;
        RECT 96.050 194.410 96.340 194.455 ;
        RECT 90.635 194.270 96.340 194.410 ;
        RECT 90.635 194.225 90.925 194.270 ;
        RECT 94.215 194.225 94.505 194.270 ;
        RECT 96.050 194.225 96.340 194.270 ;
        RECT 96.515 194.410 96.805 194.455 ;
        RECT 98.340 194.410 98.660 194.470 ;
        RECT 99.720 194.410 100.040 194.470 ;
        RECT 96.515 194.270 100.040 194.410 ;
        RECT 96.515 194.225 96.805 194.270 ;
        RECT 98.340 194.210 98.660 194.270 ;
        RECT 99.720 194.210 100.040 194.270 ;
        RECT 100.180 194.210 100.500 194.470 ;
        RECT 109.930 194.455 110.070 194.610 ;
        RECT 101.120 194.410 101.410 194.455 ;
        RECT 102.955 194.410 103.245 194.455 ;
        RECT 106.535 194.410 106.825 194.455 ;
        RECT 101.120 194.270 106.825 194.410 ;
        RECT 101.120 194.225 101.410 194.270 ;
        RECT 102.955 194.225 103.245 194.270 ;
        RECT 106.535 194.225 106.825 194.270 ;
        RECT 89.555 194.115 89.845 194.210 ;
        RECT 68.440 193.930 70.510 194.070 ;
        RECT 68.440 193.870 68.760 193.930 ;
        RECT 35.320 193.730 35.640 193.790 ;
        RECT 52.340 193.730 52.660 193.790 ;
        RECT 35.320 193.590 52.660 193.730 ;
        RECT 35.320 193.530 35.640 193.590 ;
        RECT 52.340 193.530 52.660 193.590 ;
        RECT 68.915 193.730 69.205 193.775 ;
        RECT 69.360 193.730 69.680 193.790 ;
        RECT 70.370 193.775 70.510 193.930 ;
        RECT 72.235 193.930 76.125 194.070 ;
        RECT 72.235 193.885 72.525 193.930 ;
        RECT 74.880 193.870 75.200 193.930 ;
        RECT 75.475 193.885 76.125 193.930 ;
        RECT 76.350 193.930 81.550 194.070 ;
        RECT 89.255 194.070 89.845 194.115 ;
        RECT 92.495 194.070 93.145 194.115 ;
        RECT 89.255 193.930 93.145 194.070 ;
        RECT 76.350 193.790 76.490 193.930 ;
        RECT 89.255 193.885 89.545 193.930 ;
        RECT 92.495 193.885 93.145 193.930 ;
        RECT 94.660 194.070 94.980 194.130 ;
        RECT 107.615 194.115 107.905 194.430 ;
        RECT 109.855 194.225 110.145 194.455 ;
        RECT 110.315 194.225 110.605 194.455 ;
        RECT 95.135 194.070 95.425 194.115 ;
        RECT 94.660 193.930 95.425 194.070 ;
        RECT 94.660 193.870 94.980 193.930 ;
        RECT 95.135 193.885 95.425 193.930 ;
        RECT 104.315 194.070 104.965 194.115 ;
        RECT 107.615 194.070 108.205 194.115 ;
        RECT 110.390 194.070 110.530 194.225 ;
        RECT 104.315 193.930 110.530 194.070 ;
        RECT 104.315 193.885 104.965 193.930 ;
        RECT 107.915 193.885 108.205 193.930 ;
        RECT 68.915 193.590 69.680 193.730 ;
        RECT 68.915 193.545 69.205 193.590 ;
        RECT 69.360 193.530 69.680 193.590 ;
        RECT 70.295 193.545 70.585 193.775 ;
        RECT 76.260 193.530 76.580 193.790 ;
        RECT 79.480 193.730 79.800 193.790 ;
        RECT 80.860 193.730 81.180 193.790 ;
        RECT 79.480 193.590 81.180 193.730 ;
        RECT 79.480 193.530 79.800 193.590 ;
        RECT 80.860 193.530 81.180 193.590 ;
        RECT 86.855 193.730 87.145 193.775 ;
        RECT 102.480 193.730 102.800 193.790 ;
        RECT 86.855 193.590 102.800 193.730 ;
        RECT 86.855 193.545 87.145 193.590 ;
        RECT 102.480 193.530 102.800 193.590 ;
        RECT 109.395 193.730 109.685 193.775 ;
        RECT 111.680 193.730 112.000 193.790 ;
        RECT 109.395 193.590 112.000 193.730 ;
        RECT 109.395 193.545 109.685 193.590 ;
        RECT 111.680 193.530 112.000 193.590 ;
        RECT 22.830 192.910 113.450 193.390 ;
        RECT 35.335 192.710 35.625 192.755 ;
        RECT 39.000 192.710 39.320 192.770 ;
        RECT 35.335 192.570 39.320 192.710 ;
        RECT 35.335 192.525 35.625 192.570 ;
        RECT 39.000 192.510 39.320 192.570 ;
        RECT 68.915 192.710 69.205 192.755 ;
        RECT 70.280 192.710 70.600 192.770 ;
        RECT 68.915 192.570 70.600 192.710 ;
        RECT 68.915 192.525 69.205 192.570 ;
        RECT 70.280 192.510 70.600 192.570 ;
        RECT 76.720 192.710 77.040 192.770 ;
        RECT 77.655 192.710 77.945 192.755 ;
        RECT 79.940 192.710 80.260 192.770 ;
        RECT 76.720 192.570 77.945 192.710 ;
        RECT 76.720 192.510 77.040 192.570 ;
        RECT 77.655 192.525 77.945 192.570 ;
        RECT 78.650 192.570 80.260 192.710 ;
        RECT 40.955 192.370 41.245 192.415 ;
        RECT 41.760 192.370 42.080 192.430 ;
        RECT 44.195 192.370 44.845 192.415 ;
        RECT 40.955 192.230 44.845 192.370 ;
        RECT 40.955 192.185 41.545 192.230 ;
        RECT 27.500 192.030 27.820 192.090 ;
        RECT 30.260 192.030 30.580 192.090 ;
        RECT 27.500 191.890 30.580 192.030 ;
        RECT 27.500 191.830 27.820 191.890 ;
        RECT 30.260 191.830 30.580 191.890 ;
        RECT 30.720 191.830 31.040 192.090 ;
        RECT 35.320 192.030 35.640 192.090 ;
        RECT 37.175 192.030 37.465 192.075 ;
        RECT 35.320 191.890 37.465 192.030 ;
        RECT 35.320 191.830 35.640 191.890 ;
        RECT 37.175 191.845 37.465 191.890 ;
        RECT 37.620 191.830 37.940 192.090 ;
        RECT 38.095 192.030 38.385 192.075 ;
        RECT 38.540 192.030 38.860 192.090 ;
        RECT 38.095 191.890 38.860 192.030 ;
        RECT 38.095 191.845 38.385 191.890 ;
        RECT 38.540 191.830 38.860 191.890 ;
        RECT 39.015 191.845 39.305 192.075 ;
        RECT 41.255 191.870 41.545 192.185 ;
        RECT 41.760 192.170 42.080 192.230 ;
        RECT 44.195 192.185 44.845 192.230 ;
        RECT 46.820 192.170 47.140 192.430 ;
        RECT 69.360 192.170 69.680 192.430 ;
        RECT 73.040 192.170 73.360 192.430 ;
        RECT 76.260 192.170 76.580 192.430 ;
        RECT 42.335 192.030 42.625 192.075 ;
        RECT 45.915 192.030 46.205 192.075 ;
        RECT 47.750 192.030 48.040 192.075 ;
        RECT 42.335 191.890 48.040 192.030 ;
        RECT 42.335 191.845 42.625 191.890 ;
        RECT 45.915 191.845 46.205 191.890 ;
        RECT 47.750 191.845 48.040 191.890 ;
        RECT 50.975 192.030 51.265 192.075 ;
        RECT 51.420 192.030 51.740 192.090 ;
        RECT 50.975 191.890 51.740 192.030 ;
        RECT 50.975 191.845 51.265 191.890 ;
        RECT 32.575 191.690 32.865 191.735 ;
        RECT 35.780 191.690 36.100 191.750 ;
        RECT 39.090 191.690 39.230 191.845 ;
        RECT 51.420 191.830 51.740 191.890 ;
        RECT 56.035 192.030 56.325 192.075 ;
        RECT 56.940 192.030 57.260 192.090 ;
        RECT 60.620 192.030 60.940 192.090 ;
        RECT 56.035 191.890 60.940 192.030 ;
        RECT 56.035 191.845 56.325 191.890 ;
        RECT 56.940 191.830 57.260 191.890 ;
        RECT 60.620 191.830 60.940 191.890 ;
        RECT 65.680 192.030 66.000 192.090 ;
        RECT 73.960 192.030 74.280 192.090 ;
        RECT 78.650 192.075 78.790 192.570 ;
        RECT 79.940 192.510 80.260 192.570 ;
        RECT 84.555 192.710 84.845 192.755 ;
        RECT 86.380 192.710 86.700 192.770 ;
        RECT 84.555 192.570 86.700 192.710 ;
        RECT 84.555 192.525 84.845 192.570 ;
        RECT 86.380 192.510 86.700 192.570 ;
        RECT 86.840 192.710 87.160 192.770 ;
        RECT 90.075 192.710 90.365 192.755 ;
        RECT 86.840 192.570 90.365 192.710 ;
        RECT 86.840 192.510 87.160 192.570 ;
        RECT 90.075 192.525 90.365 192.570 ;
        RECT 91.915 192.525 92.205 192.755 ;
        RECT 93.295 192.710 93.585 192.755 ;
        RECT 94.660 192.710 94.980 192.770 ;
        RECT 93.295 192.570 94.980 192.710 ;
        RECT 93.295 192.525 93.585 192.570 ;
        RECT 79.480 192.370 79.800 192.430 ;
        RECT 79.110 192.230 79.800 192.370 ;
        RECT 74.895 192.030 75.185 192.075 ;
        RECT 65.680 191.890 75.185 192.030 ;
        RECT 65.680 191.830 66.000 191.890 ;
        RECT 73.960 191.830 74.280 191.890 ;
        RECT 74.895 191.845 75.185 191.890 ;
        RECT 78.575 191.845 78.865 192.075 ;
        RECT 32.575 191.550 36.100 191.690 ;
        RECT 32.575 191.505 32.865 191.550 ;
        RECT 35.780 191.490 36.100 191.550 ;
        RECT 38.630 191.550 39.230 191.690 ;
        RECT 43.140 191.690 43.460 191.750 ;
        RECT 48.215 191.690 48.505 191.735 ;
        RECT 43.140 191.550 48.505 191.690 ;
        RECT 32.100 191.350 32.420 191.410 ;
        RECT 34.400 191.350 34.720 191.410 ;
        RECT 38.630 191.350 38.770 191.550 ;
        RECT 43.140 191.490 43.460 191.550 ;
        RECT 48.215 191.505 48.505 191.550 ;
        RECT 51.880 191.490 52.200 191.750 ;
        RECT 70.740 191.690 71.060 191.750 ;
        RECT 78.650 191.690 78.790 191.845 ;
        RECT 70.740 191.550 78.790 191.690 ;
        RECT 70.740 191.490 71.060 191.550 ;
        RECT 32.100 191.210 38.770 191.350 ;
        RECT 42.335 191.350 42.625 191.395 ;
        RECT 45.455 191.350 45.745 191.395 ;
        RECT 47.345 191.350 47.635 191.395 ;
        RECT 79.110 191.350 79.250 192.230 ;
        RECT 79.480 192.170 79.800 192.230 ;
        RECT 80.400 192.370 80.720 192.430 ;
        RECT 82.255 192.370 82.545 192.415 ;
        RECT 85.920 192.370 86.240 192.430 ;
        RECT 80.400 192.230 86.240 192.370 ;
        RECT 80.400 192.170 80.720 192.230 ;
        RECT 82.255 192.185 82.545 192.230 ;
        RECT 85.920 192.170 86.240 192.230 ;
        RECT 82.715 192.030 83.005 192.075 ;
        RECT 79.570 191.890 83.005 192.030 ;
        RECT 79.570 191.750 79.710 191.890 ;
        RECT 82.715 191.845 83.005 191.890 ;
        RECT 86.380 191.830 86.700 192.090 ;
        RECT 86.840 192.030 87.160 192.090 ;
        RECT 87.775 192.030 88.065 192.075 ;
        RECT 86.840 191.890 88.065 192.030 ;
        RECT 91.990 192.030 92.130 192.525 ;
        RECT 94.660 192.510 94.980 192.570 ;
        RECT 97.420 192.510 97.740 192.770 ;
        RECT 102.480 192.510 102.800 192.770 ;
        RECT 104.320 192.510 104.640 192.770 ;
        RECT 92.375 192.030 92.665 192.075 ;
        RECT 95.595 192.030 95.885 192.075 ;
        RECT 91.990 191.890 92.665 192.030 ;
        RECT 86.840 191.830 87.160 191.890 ;
        RECT 87.775 191.845 88.065 191.890 ;
        RECT 92.375 191.845 92.665 191.890 ;
        RECT 92.910 191.890 95.885 192.030 ;
        RECT 79.480 191.490 79.800 191.750 ;
        RECT 81.320 191.690 81.640 191.750 ;
        RECT 88.680 191.690 89.000 191.750 ;
        RECT 81.320 191.550 89.000 191.690 ;
        RECT 81.320 191.490 81.640 191.550 ;
        RECT 88.680 191.490 89.000 191.550 ;
        RECT 89.615 191.690 89.905 191.735 ;
        RECT 90.520 191.690 90.840 191.750 ;
        RECT 92.910 191.690 93.050 191.890 ;
        RECT 95.595 191.845 95.885 191.890 ;
        RECT 98.815 192.030 99.105 192.075 ;
        RECT 104.795 192.030 105.085 192.075 ;
        RECT 98.815 191.890 105.085 192.030 ;
        RECT 98.815 191.845 99.105 191.890 ;
        RECT 104.795 191.845 105.085 191.890 ;
        RECT 89.615 191.550 93.050 191.690 ;
        RECT 89.615 191.505 89.905 191.550 ;
        RECT 90.520 191.490 90.840 191.550 ;
        RECT 94.200 191.490 94.520 191.750 ;
        RECT 95.135 191.690 95.425 191.735 ;
        RECT 96.500 191.690 96.820 191.750 ;
        RECT 95.135 191.550 96.820 191.690 ;
        RECT 95.135 191.505 95.425 191.550 ;
        RECT 87.315 191.350 87.605 191.395 ;
        RECT 42.335 191.210 47.635 191.350 ;
        RECT 32.100 191.150 32.420 191.210 ;
        RECT 34.400 191.150 34.720 191.210 ;
        RECT 42.335 191.165 42.625 191.210 ;
        RECT 45.455 191.165 45.745 191.210 ;
        RECT 47.345 191.165 47.635 191.210 ;
        RECT 73.590 191.210 79.250 191.350 ;
        RECT 85.090 191.210 87.605 191.350 ;
        RECT 29.815 191.010 30.105 191.055 ;
        RECT 30.260 191.010 30.580 191.070 ;
        RECT 29.815 190.870 30.580 191.010 ;
        RECT 29.815 190.825 30.105 190.870 ;
        RECT 30.260 190.810 30.580 190.870 ;
        RECT 31.640 190.810 31.960 191.070 ;
        RECT 35.320 191.010 35.640 191.070 ;
        RECT 35.795 191.010 36.085 191.055 ;
        RECT 35.320 190.870 36.085 191.010 ;
        RECT 35.320 190.810 35.640 190.870 ;
        RECT 35.795 190.825 36.085 190.870 ;
        RECT 39.460 190.810 39.780 191.070 ;
        RECT 44.520 191.010 44.840 191.070 ;
        RECT 50.055 191.010 50.345 191.055 ;
        RECT 44.520 190.870 50.345 191.010 ;
        RECT 44.520 190.810 44.840 190.870 ;
        RECT 50.055 190.825 50.345 190.870 ;
        RECT 54.640 190.810 54.960 191.070 ;
        RECT 55.575 191.010 55.865 191.055 ;
        RECT 56.020 191.010 56.340 191.070 ;
        RECT 55.575 190.870 56.340 191.010 ;
        RECT 55.575 190.825 55.865 190.870 ;
        RECT 56.020 190.810 56.340 190.870 ;
        RECT 66.140 191.010 66.460 191.070 ;
        RECT 72.120 191.010 72.440 191.070 ;
        RECT 73.590 191.055 73.730 191.210 ;
        RECT 73.515 191.010 73.805 191.055 ;
        RECT 66.140 190.870 73.805 191.010 ;
        RECT 66.140 190.810 66.460 190.870 ;
        RECT 72.120 190.810 72.440 190.870 ;
        RECT 73.515 190.825 73.805 190.870 ;
        RECT 83.160 191.010 83.480 191.070 ;
        RECT 85.090 191.010 85.230 191.210 ;
        RECT 87.315 191.165 87.605 191.210 ;
        RECT 90.980 191.350 91.300 191.410 ;
        RECT 95.210 191.350 95.350 191.505 ;
        RECT 96.500 191.490 96.820 191.550 ;
        RECT 101.100 191.490 101.420 191.750 ;
        RECT 102.020 191.490 102.340 191.750 ;
        RECT 104.320 191.690 104.640 191.750 ;
        RECT 107.555 191.690 107.845 191.735 ;
        RECT 104.320 191.550 107.845 191.690 ;
        RECT 104.320 191.490 104.640 191.550 ;
        RECT 107.555 191.505 107.845 191.550 ;
        RECT 111.680 191.490 112.000 191.750 ;
        RECT 90.980 191.210 95.350 191.350 ;
        RECT 102.110 191.350 102.250 191.490 ;
        RECT 108.475 191.350 108.765 191.395 ;
        RECT 102.110 191.210 108.765 191.350 ;
        RECT 90.980 191.150 91.300 191.210 ;
        RECT 108.475 191.165 108.765 191.210 ;
        RECT 83.160 190.870 85.230 191.010 ;
        RECT 83.160 190.810 83.480 190.870 ;
        RECT 85.460 190.810 85.780 191.070 ;
        RECT 99.735 191.010 100.025 191.055 ;
        RECT 102.480 191.010 102.800 191.070 ;
        RECT 99.735 190.870 102.800 191.010 ;
        RECT 99.735 190.825 100.025 190.870 ;
        RECT 102.480 190.810 102.800 190.870 ;
        RECT 22.830 190.190 113.450 190.670 ;
        RECT 28.435 189.990 28.725 190.035 ;
        RECT 30.720 189.990 31.040 190.050 ;
        RECT 28.435 189.850 31.040 189.990 ;
        RECT 28.435 189.805 28.725 189.850 ;
        RECT 30.720 189.790 31.040 189.850 ;
        RECT 34.400 189.990 34.720 190.050 ;
        RECT 35.320 189.990 35.640 190.050 ;
        RECT 39.460 189.990 39.780 190.050 ;
        RECT 34.400 189.850 35.640 189.990 ;
        RECT 34.400 189.790 34.720 189.850 ;
        RECT 35.320 189.790 35.640 189.850 ;
        RECT 36.790 189.850 39.780 189.990 ;
        RECT 36.255 189.650 36.545 189.695 ;
        RECT 31.730 189.510 36.545 189.650 ;
        RECT 31.730 189.355 31.870 189.510 ;
        RECT 36.255 189.465 36.545 189.510 ;
        RECT 31.655 189.125 31.945 189.355 ;
        RECT 32.100 189.110 32.420 189.370 ;
        RECT 36.790 189.310 36.930 189.850 ;
        RECT 39.460 189.790 39.780 189.850 ;
        RECT 41.760 189.990 42.080 190.050 ;
        RECT 42.235 189.990 42.525 190.035 ;
        RECT 51.880 189.990 52.200 190.050 ;
        RECT 52.355 189.990 52.645 190.035 ;
        RECT 41.760 189.850 42.525 189.990 ;
        RECT 41.760 189.790 42.080 189.850 ;
        RECT 42.235 189.805 42.525 189.850 ;
        RECT 43.690 189.850 52.645 189.990 ;
        RECT 37.620 189.650 37.940 189.710 ;
        RECT 43.690 189.650 43.830 189.850 ;
        RECT 51.880 189.790 52.200 189.850 ;
        RECT 52.355 189.805 52.645 189.850 ;
        RECT 100.640 189.790 100.960 190.050 ;
        RECT 37.620 189.510 43.830 189.650 ;
        RECT 44.025 189.650 44.315 189.695 ;
        RECT 45.915 189.650 46.205 189.695 ;
        RECT 49.035 189.650 49.325 189.695 ;
        RECT 44.025 189.510 49.325 189.650 ;
        RECT 37.620 189.450 37.940 189.510 ;
        RECT 44.025 189.465 44.315 189.510 ;
        RECT 45.915 189.465 46.205 189.510 ;
        RECT 49.035 189.465 49.325 189.510 ;
        RECT 55.215 189.650 55.505 189.695 ;
        RECT 58.335 189.650 58.625 189.695 ;
        RECT 60.225 189.650 60.515 189.695 ;
        RECT 55.215 189.510 60.515 189.650 ;
        RECT 55.215 189.465 55.505 189.510 ;
        RECT 58.335 189.465 58.625 189.510 ;
        RECT 60.225 189.465 60.515 189.510 ;
        RECT 69.820 189.650 70.140 189.710 ;
        RECT 81.750 189.650 82.040 189.695 ;
        RECT 84.530 189.650 84.820 189.695 ;
        RECT 86.390 189.650 86.680 189.695 ;
        RECT 101.100 189.650 101.420 189.710 ;
        RECT 69.820 189.510 72.810 189.650 ;
        RECT 69.820 189.450 70.140 189.510 ;
        RECT 34.490 189.170 36.930 189.310 ;
        RECT 38.080 189.310 38.400 189.370 ;
        RECT 39.015 189.310 39.305 189.355 ;
        RECT 38.080 189.170 39.305 189.310 ;
        RECT 24.755 188.970 25.045 189.015 ;
        RECT 26.580 188.970 26.900 189.030 ;
        RECT 24.755 188.830 26.900 188.970 ;
        RECT 24.755 188.785 25.045 188.830 ;
        RECT 26.580 188.770 26.900 188.830 ;
        RECT 33.480 188.770 33.800 189.030 ;
        RECT 33.940 188.770 34.260 189.030 ;
        RECT 34.490 189.015 34.630 189.170 ;
        RECT 38.080 189.110 38.400 189.170 ;
        RECT 39.015 189.125 39.305 189.170 ;
        RECT 43.140 189.110 43.460 189.370 ;
        RECT 44.520 189.110 44.840 189.370 ;
        RECT 50.500 189.310 50.820 189.370 ;
        RECT 59.715 189.310 60.005 189.355 ;
        RECT 50.500 189.170 60.005 189.310 ;
        RECT 50.500 189.110 50.820 189.170 ;
        RECT 59.715 189.125 60.005 189.170 ;
        RECT 61.080 189.110 61.400 189.370 ;
        RECT 67.980 189.310 68.300 189.370 ;
        RECT 68.455 189.310 68.745 189.355 ;
        RECT 67.980 189.170 68.745 189.310 ;
        RECT 67.980 189.110 68.300 189.170 ;
        RECT 68.455 189.125 68.745 189.170 ;
        RECT 68.915 189.310 69.205 189.355 ;
        RECT 69.910 189.310 70.050 189.450 ;
        RECT 70.740 189.310 71.060 189.370 ;
        RECT 72.670 189.355 72.810 189.510 ;
        RECT 81.750 189.510 86.680 189.650 ;
        RECT 81.750 189.465 82.040 189.510 ;
        RECT 84.530 189.465 84.820 189.510 ;
        RECT 86.390 189.465 86.680 189.510 ;
        RECT 97.510 189.510 101.420 189.650 ;
        RECT 71.675 189.310 71.965 189.355 ;
        RECT 68.915 189.170 70.050 189.310 ;
        RECT 70.370 189.170 71.965 189.310 ;
        RECT 68.915 189.125 69.205 189.170 ;
        RECT 34.415 188.785 34.705 189.015 ;
        RECT 35.335 188.970 35.625 189.015 ;
        RECT 36.700 188.970 37.020 189.030 ;
        RECT 35.335 188.830 37.020 188.970 ;
        RECT 35.335 188.785 35.625 188.830 ;
        RECT 36.700 188.770 37.020 188.830 ;
        RECT 40.380 188.770 40.700 189.030 ;
        RECT 41.775 188.785 42.065 189.015 ;
        RECT 43.620 188.970 43.910 189.015 ;
        RECT 45.455 188.970 45.745 189.015 ;
        RECT 49.035 188.970 49.325 189.015 ;
        RECT 43.620 188.830 49.325 188.970 ;
        RECT 43.620 188.785 43.910 188.830 ;
        RECT 45.455 188.785 45.745 188.830 ;
        RECT 49.035 188.785 49.325 188.830 ;
        RECT 26.670 188.630 26.810 188.770 ;
        RECT 38.540 188.630 38.860 188.690 ;
        RECT 26.670 188.490 38.860 188.630 ;
        RECT 41.850 188.630 41.990 188.785 ;
        RECT 44.520 188.630 44.840 188.690 ;
        RECT 50.115 188.675 50.405 188.990 ;
        RECT 41.850 188.490 44.840 188.630 ;
        RECT 38.540 188.430 38.860 188.490 ;
        RECT 44.520 188.430 44.840 188.490 ;
        RECT 46.815 188.630 47.465 188.675 ;
        RECT 50.115 188.630 50.705 188.675 ;
        RECT 50.960 188.630 51.280 188.690 ;
        RECT 54.135 188.675 54.425 188.990 ;
        RECT 55.215 188.970 55.505 189.015 ;
        RECT 58.795 188.970 59.085 189.015 ;
        RECT 60.630 188.970 60.920 189.015 ;
        RECT 55.215 188.830 60.920 188.970 ;
        RECT 69.375 188.955 69.665 189.015 ;
        RECT 55.215 188.785 55.505 188.830 ;
        RECT 58.795 188.785 59.085 188.830 ;
        RECT 60.630 188.785 60.920 188.830 ;
        RECT 68.990 188.815 69.665 188.955 ;
        RECT 46.815 188.490 51.280 188.630 ;
        RECT 46.815 188.445 47.465 188.490 ;
        RECT 50.415 188.445 50.705 188.490 ;
        RECT 50.960 188.430 51.280 188.490 ;
        RECT 53.835 188.630 54.425 188.675 ;
        RECT 56.020 188.630 56.340 188.690 ;
        RECT 57.075 188.630 57.725 188.675 ;
        RECT 53.835 188.490 57.725 188.630 ;
        RECT 53.835 188.445 54.125 188.490 ;
        RECT 56.020 188.430 56.340 188.490 ;
        RECT 57.075 188.445 57.725 188.490 ;
        RECT 67.535 188.630 67.825 188.675 ;
        RECT 68.440 188.630 68.760 188.690 ;
        RECT 67.535 188.490 68.760 188.630 ;
        RECT 68.990 188.630 69.130 188.815 ;
        RECT 69.375 188.785 69.665 188.815 ;
        RECT 69.925 188.970 70.215 189.015 ;
        RECT 70.370 188.970 70.510 189.170 ;
        RECT 70.740 189.110 71.060 189.170 ;
        RECT 71.675 189.125 71.965 189.170 ;
        RECT 72.595 189.125 72.885 189.355 ;
        RECT 85.015 189.310 85.305 189.355 ;
        RECT 85.460 189.310 85.780 189.370 ;
        RECT 85.015 189.170 85.780 189.310 ;
        RECT 85.015 189.125 85.305 189.170 ;
        RECT 85.460 189.110 85.780 189.170 ;
        RECT 88.680 189.310 89.000 189.370 ;
        RECT 92.375 189.310 92.665 189.355 ;
        RECT 94.200 189.310 94.520 189.370 ;
        RECT 97.510 189.355 97.650 189.510 ;
        RECT 101.100 189.450 101.420 189.510 ;
        RECT 103.975 189.650 104.265 189.695 ;
        RECT 107.095 189.650 107.385 189.695 ;
        RECT 108.985 189.650 109.275 189.695 ;
        RECT 103.975 189.510 109.275 189.650 ;
        RECT 103.975 189.465 104.265 189.510 ;
        RECT 107.095 189.465 107.385 189.510 ;
        RECT 108.985 189.465 109.275 189.510 ;
        RECT 97.435 189.310 97.725 189.355 ;
        RECT 100.180 189.310 100.500 189.370 ;
        RECT 88.680 189.170 97.725 189.310 ;
        RECT 88.680 189.110 89.000 189.170 ;
        RECT 92.375 189.125 92.665 189.170 ;
        RECT 94.200 189.110 94.520 189.170 ;
        RECT 97.435 189.125 97.725 189.170 ;
        RECT 98.430 189.170 100.500 189.310 ;
        RECT 69.925 188.830 70.510 188.970 ;
        RECT 69.925 188.785 70.215 188.830 ;
        RECT 71.200 188.770 71.520 189.030 ;
        RECT 72.120 188.770 72.440 189.030 ;
        RECT 73.960 188.770 74.280 189.030 ;
        RECT 81.750 188.970 82.040 189.015 ;
        RECT 86.855 188.970 87.145 189.015 ;
        RECT 87.300 188.970 87.620 189.030 ;
        RECT 81.750 188.830 84.285 188.970 ;
        RECT 81.750 188.785 82.040 188.830 ;
        RECT 72.210 188.630 72.350 188.770 ;
        RECT 68.990 188.490 72.350 188.630 ;
        RECT 73.040 188.630 73.360 188.690 ;
        RECT 73.515 188.630 73.805 188.675 ;
        RECT 73.040 188.490 73.805 188.630 ;
        RECT 67.535 188.445 67.825 188.490 ;
        RECT 68.440 188.430 68.760 188.490 ;
        RECT 73.040 188.430 73.360 188.490 ;
        RECT 73.515 188.445 73.805 188.490 ;
        RECT 75.355 188.630 75.645 188.675 ;
        RECT 75.800 188.630 76.120 188.690 ;
        RECT 83.160 188.675 83.480 188.690 ;
        RECT 75.355 188.490 76.120 188.630 ;
        RECT 75.355 188.445 75.645 188.490 ;
        RECT 75.800 188.430 76.120 188.490 ;
        RECT 79.890 188.630 80.180 188.675 ;
        RECT 83.150 188.630 83.480 188.675 ;
        RECT 79.890 188.490 83.480 188.630 ;
        RECT 79.890 188.445 80.180 188.490 ;
        RECT 83.150 188.445 83.480 188.490 ;
        RECT 84.070 188.675 84.285 188.830 ;
        RECT 86.855 188.830 87.620 188.970 ;
        RECT 86.855 188.785 87.145 188.830 ;
        RECT 87.300 188.770 87.620 188.830 ;
        RECT 87.760 188.770 88.080 189.030 ;
        RECT 90.995 188.970 91.285 189.015 ;
        RECT 93.295 188.970 93.585 189.015 ;
        RECT 90.995 188.830 93.585 188.970 ;
        RECT 90.995 188.785 91.285 188.830 ;
        RECT 93.295 188.785 93.585 188.830 ;
        RECT 93.755 188.970 94.045 189.015 ;
        RECT 98.430 188.970 98.570 189.170 ;
        RECT 100.180 189.110 100.500 189.170 ;
        RECT 93.755 188.830 98.570 188.970 ;
        RECT 98.815 188.970 99.105 189.015 ;
        RECT 102.020 188.970 102.340 189.030 ;
        RECT 98.815 188.830 102.340 188.970 ;
        RECT 93.755 188.785 94.045 188.830 ;
        RECT 98.815 188.785 99.105 188.830 ;
        RECT 102.020 188.770 102.340 188.830 ;
        RECT 84.070 188.630 84.360 188.675 ;
        RECT 85.930 188.630 86.220 188.675 ;
        RECT 84.070 188.490 86.220 188.630 ;
        RECT 84.070 188.445 84.360 188.490 ;
        RECT 85.930 188.445 86.220 188.490 ;
        RECT 99.260 188.630 99.580 188.690 ;
        RECT 102.895 188.675 103.185 188.990 ;
        RECT 103.975 188.970 104.265 189.015 ;
        RECT 107.555 188.970 107.845 189.015 ;
        RECT 109.390 188.970 109.680 189.015 ;
        RECT 103.975 188.830 109.680 188.970 ;
        RECT 103.975 188.785 104.265 188.830 ;
        RECT 107.555 188.785 107.845 188.830 ;
        RECT 109.390 188.785 109.680 188.830 ;
        RECT 109.855 188.970 110.145 189.015 ;
        RECT 110.300 188.970 110.620 189.030 ;
        RECT 109.855 188.830 110.620 188.970 ;
        RECT 109.855 188.785 110.145 188.830 ;
        RECT 110.300 188.770 110.620 188.830 ;
        RECT 111.220 188.770 111.540 189.030 ;
        RECT 102.595 188.630 103.185 188.675 ;
        RECT 105.835 188.630 106.485 188.675 ;
        RECT 99.260 188.490 106.485 188.630 ;
        RECT 83.160 188.430 83.480 188.445 ;
        RECT 99.260 188.430 99.580 188.490 ;
        RECT 102.595 188.445 102.885 188.490 ;
        RECT 105.835 188.445 106.485 188.490 ;
        RECT 107.080 188.630 107.400 188.690 ;
        RECT 108.475 188.630 108.765 188.675 ;
        RECT 107.080 188.490 108.765 188.630 ;
        RECT 107.080 188.430 107.400 188.490 ;
        RECT 108.475 188.445 108.765 188.490 ;
        RECT 27.515 188.290 27.805 188.335 ;
        RECT 28.420 188.290 28.740 188.350 ;
        RECT 27.515 188.150 28.740 188.290 ;
        RECT 27.515 188.105 27.805 188.150 ;
        RECT 28.420 188.090 28.740 188.150 ;
        RECT 29.800 188.290 30.120 188.350 ;
        RECT 33.480 188.290 33.800 188.350 ;
        RECT 34.860 188.290 35.180 188.350 ;
        RECT 29.800 188.150 35.180 188.290 ;
        RECT 29.800 188.090 30.120 188.150 ;
        RECT 33.480 188.090 33.800 188.150 ;
        RECT 34.860 188.090 35.180 188.150 ;
        RECT 38.095 188.290 38.385 188.335 ;
        RECT 39.000 188.290 39.320 188.350 ;
        RECT 38.095 188.150 39.320 188.290 ;
        RECT 38.095 188.105 38.385 188.150 ;
        RECT 39.000 188.090 39.320 188.150 ;
        RECT 41.315 188.290 41.605 188.335 ;
        RECT 41.760 188.290 42.080 188.350 ;
        RECT 41.315 188.150 42.080 188.290 ;
        RECT 41.315 188.105 41.605 188.150 ;
        RECT 41.760 188.090 42.080 188.150 ;
        RECT 45.900 188.290 46.220 188.350 ;
        RECT 51.895 188.290 52.185 188.335 ;
        RECT 45.900 188.150 52.185 188.290 ;
        RECT 45.900 188.090 46.220 188.150 ;
        RECT 51.895 188.105 52.185 188.150 ;
        RECT 67.980 188.290 68.300 188.350 ;
        RECT 70.280 188.290 70.600 188.350 ;
        RECT 71.200 188.290 71.520 188.350 ;
        RECT 67.980 188.150 71.520 188.290 ;
        RECT 67.980 188.090 68.300 188.150 ;
        RECT 70.280 188.090 70.600 188.150 ;
        RECT 71.200 188.090 71.520 188.150 ;
        RECT 77.885 188.290 78.175 188.335 ;
        RECT 80.400 188.290 80.720 188.350 ;
        RECT 77.885 188.150 80.720 188.290 ;
        RECT 77.885 188.105 78.175 188.150 ;
        RECT 80.400 188.090 80.720 188.150 ;
        RECT 95.595 188.290 95.885 188.335 ;
        RECT 96.040 188.290 96.360 188.350 ;
        RECT 95.595 188.150 96.360 188.290 ;
        RECT 95.595 188.105 95.885 188.150 ;
        RECT 96.040 188.090 96.360 188.150 ;
        RECT 98.355 188.290 98.645 188.335 ;
        RECT 101.100 188.290 101.420 188.350 ;
        RECT 98.355 188.150 101.420 188.290 ;
        RECT 98.355 188.105 98.645 188.150 ;
        RECT 101.100 188.090 101.420 188.150 ;
        RECT 110.315 188.290 110.605 188.335 ;
        RECT 110.760 188.290 111.080 188.350 ;
        RECT 110.315 188.150 111.080 188.290 ;
        RECT 110.315 188.105 110.605 188.150 ;
        RECT 110.760 188.090 111.080 188.150 ;
        RECT 22.830 187.470 113.450 187.950 ;
        RECT 26.580 187.070 26.900 187.330 ;
        RECT 35.780 187.070 36.100 187.330 ;
        RECT 41.300 187.270 41.620 187.330 ;
        RECT 50.500 187.270 50.820 187.330 ;
        RECT 50.975 187.270 51.265 187.315 ;
        RECT 41.300 187.130 45.210 187.270 ;
        RECT 41.300 187.070 41.620 187.130 ;
        RECT 28.075 186.930 28.365 186.975 ;
        RECT 30.260 186.930 30.580 186.990 ;
        RECT 31.315 186.930 31.965 186.975 ;
        RECT 28.075 186.790 31.965 186.930 ;
        RECT 28.075 186.745 28.665 186.790 ;
        RECT 28.375 186.430 28.665 186.745 ;
        RECT 30.260 186.730 30.580 186.790 ;
        RECT 31.315 186.745 31.965 186.790 ;
        RECT 36.240 186.930 36.560 186.990 ;
        RECT 37.275 186.930 37.565 186.975 ;
        RECT 40.515 186.930 41.165 186.975 ;
        RECT 36.240 186.790 41.165 186.930 ;
        RECT 36.240 186.730 36.560 186.790 ;
        RECT 37.275 186.745 37.865 186.790 ;
        RECT 40.515 186.745 41.165 186.790 ;
        RECT 41.760 186.930 42.080 186.990 ;
        RECT 43.155 186.930 43.445 186.975 ;
        RECT 41.760 186.790 43.445 186.930 ;
        RECT 29.455 186.590 29.745 186.635 ;
        RECT 33.035 186.590 33.325 186.635 ;
        RECT 34.870 186.590 35.160 186.635 ;
        RECT 29.455 186.450 35.160 186.590 ;
        RECT 29.455 186.405 29.745 186.450 ;
        RECT 33.035 186.405 33.325 186.450 ;
        RECT 34.870 186.405 35.160 186.450 ;
        RECT 37.575 186.430 37.865 186.745 ;
        RECT 41.760 186.730 42.080 186.790 ;
        RECT 43.155 186.745 43.445 186.790 ;
        RECT 45.070 186.930 45.210 187.130 ;
        RECT 50.500 187.130 51.265 187.270 ;
        RECT 50.500 187.070 50.820 187.130 ;
        RECT 50.975 187.085 51.265 187.130 ;
        RECT 51.420 187.070 51.740 187.330 ;
        RECT 52.340 187.270 52.660 187.330 ;
        RECT 66.140 187.270 66.460 187.330 ;
        RECT 52.340 187.130 69.590 187.270 ;
        RECT 52.340 187.070 52.660 187.130 ;
        RECT 66.140 187.070 66.460 187.130 ;
        RECT 51.880 186.930 52.200 186.990 ;
        RECT 45.070 186.790 52.200 186.930 ;
        RECT 45.070 186.635 45.210 186.790 ;
        RECT 51.880 186.730 52.200 186.790 ;
        RECT 53.275 186.930 53.565 186.975 ;
        RECT 54.640 186.930 54.960 186.990 ;
        RECT 57.875 186.930 58.165 186.975 ;
        RECT 67.535 186.930 67.825 186.975 ;
        RECT 67.980 186.930 68.300 186.990 ;
        RECT 53.275 186.790 58.165 186.930 ;
        RECT 53.275 186.745 53.565 186.790 ;
        RECT 54.640 186.730 54.960 186.790 ;
        RECT 57.875 186.745 58.165 186.790 ;
        RECT 65.310 186.790 68.300 186.930 ;
        RECT 69.450 186.930 69.590 187.130 ;
        RECT 69.820 187.070 70.140 187.330 ;
        RECT 70.295 187.270 70.585 187.315 ;
        RECT 70.740 187.270 71.060 187.330 ;
        RECT 88.680 187.270 89.000 187.330 ;
        RECT 70.295 187.130 71.060 187.270 ;
        RECT 70.295 187.085 70.585 187.130 ;
        RECT 70.740 187.070 71.060 187.130 ;
        RECT 75.890 187.130 89.000 187.270 ;
        RECT 75.890 186.930 76.030 187.130 ;
        RECT 88.680 187.070 89.000 187.130 ;
        RECT 95.120 187.270 95.440 187.330 ;
        RECT 96.960 187.270 97.280 187.330 ;
        RECT 101.575 187.270 101.865 187.315 ;
        RECT 95.120 187.130 101.865 187.270 ;
        RECT 95.120 187.070 95.440 187.130 ;
        RECT 96.960 187.070 97.280 187.130 ;
        RECT 101.575 187.085 101.865 187.130 ;
        RECT 102.480 187.270 102.800 187.330 ;
        RECT 109.840 187.270 110.160 187.330 ;
        RECT 111.235 187.270 111.525 187.315 ;
        RECT 102.480 187.130 109.150 187.270 ;
        RECT 102.480 187.070 102.800 187.130 ;
        RECT 109.010 186.975 109.150 187.130 ;
        RECT 109.840 187.130 111.525 187.270 ;
        RECT 109.840 187.070 110.160 187.130 ;
        RECT 111.235 187.085 111.525 187.130 ;
        RECT 69.450 186.790 76.030 186.930 ;
        RECT 76.275 186.930 76.565 186.975 ;
        RECT 79.430 186.930 79.720 186.975 ;
        RECT 82.690 186.930 82.980 186.975 ;
        RECT 76.275 186.790 82.980 186.930 ;
        RECT 38.655 186.590 38.945 186.635 ;
        RECT 42.235 186.590 42.525 186.635 ;
        RECT 44.070 186.590 44.360 186.635 ;
        RECT 38.655 186.450 44.360 186.590 ;
        RECT 38.655 186.405 38.945 186.450 ;
        RECT 42.235 186.405 42.525 186.450 ;
        RECT 44.070 186.405 44.360 186.450 ;
        RECT 44.995 186.405 45.285 186.635 ;
        RECT 45.900 186.390 46.220 186.650 ;
        RECT 46.360 186.390 46.680 186.650 ;
        RECT 46.835 186.405 47.125 186.635 ;
        RECT 50.055 186.405 50.345 186.635 ;
        RECT 56.480 186.590 56.800 186.650 ;
        RECT 57.415 186.590 57.705 186.635 ;
        RECT 56.480 186.450 57.705 186.590 ;
        RECT 31.640 186.250 31.960 186.310 ;
        RECT 33.955 186.250 34.245 186.295 ;
        RECT 31.640 186.110 34.245 186.250 ;
        RECT 31.640 186.050 31.960 186.110 ;
        RECT 33.955 186.065 34.245 186.110 ;
        RECT 35.320 186.250 35.640 186.310 ;
        RECT 43.140 186.250 43.460 186.310 ;
        RECT 44.535 186.250 44.825 186.295 ;
        RECT 46.910 186.250 47.050 186.405 ;
        RECT 35.320 186.110 44.825 186.250 ;
        RECT 35.320 186.050 35.640 186.110 ;
        RECT 43.140 186.050 43.460 186.110 ;
        RECT 44.535 186.065 44.825 186.110 ;
        RECT 46.450 186.110 47.050 186.250 ;
        RECT 29.455 185.910 29.745 185.955 ;
        RECT 32.575 185.910 32.865 185.955 ;
        RECT 34.465 185.910 34.755 185.955 ;
        RECT 29.455 185.770 34.755 185.910 ;
        RECT 29.455 185.725 29.745 185.770 ;
        RECT 32.575 185.725 32.865 185.770 ;
        RECT 34.465 185.725 34.755 185.770 ;
        RECT 38.655 185.910 38.945 185.955 ;
        RECT 41.775 185.910 42.065 185.955 ;
        RECT 43.665 185.910 43.955 185.955 ;
        RECT 38.655 185.770 43.955 185.910 ;
        RECT 38.655 185.725 38.945 185.770 ;
        RECT 41.775 185.725 42.065 185.770 ;
        RECT 43.665 185.725 43.955 185.770 ;
        RECT 42.680 185.570 43.000 185.630 ;
        RECT 46.450 185.570 46.590 186.110 ;
        RECT 50.130 185.910 50.270 186.405 ;
        RECT 56.480 186.390 56.800 186.450 ;
        RECT 57.415 186.405 57.705 186.450 ;
        RECT 60.620 186.390 60.940 186.650 ;
        RECT 62.935 186.405 63.225 186.635 ;
        RECT 53.260 186.250 53.580 186.310 ;
        RECT 53.735 186.250 54.025 186.295 ;
        RECT 53.260 186.110 54.025 186.250 ;
        RECT 53.260 186.050 53.580 186.110 ;
        RECT 53.735 186.065 54.025 186.110 ;
        RECT 54.640 186.250 54.960 186.310 ;
        RECT 58.335 186.250 58.625 186.295 ;
        RECT 63.010 186.250 63.150 186.405 ;
        RECT 64.760 186.390 65.080 186.650 ;
        RECT 65.310 186.635 65.450 186.790 ;
        RECT 67.535 186.745 67.825 186.790 ;
        RECT 67.980 186.730 68.300 186.790 ;
        RECT 76.275 186.745 76.565 186.790 ;
        RECT 79.430 186.745 79.720 186.790 ;
        RECT 82.690 186.745 82.980 186.790 ;
        RECT 83.610 186.930 83.900 186.975 ;
        RECT 85.470 186.930 85.760 186.975 ;
        RECT 83.610 186.790 85.760 186.930 ;
        RECT 83.610 186.745 83.900 186.790 ;
        RECT 85.470 186.745 85.760 186.790 ;
        RECT 87.315 186.930 87.605 186.975 ;
        RECT 89.715 186.930 90.005 186.975 ;
        RECT 92.955 186.930 93.605 186.975 ;
        RECT 87.315 186.790 88.910 186.930 ;
        RECT 87.315 186.745 87.605 186.790 ;
        RECT 65.235 186.405 65.525 186.635 ;
        RECT 66.155 186.590 66.445 186.635 ;
        RECT 69.820 186.590 70.140 186.650 ;
        RECT 66.155 186.450 70.140 186.590 ;
        RECT 66.155 186.405 66.445 186.450 ;
        RECT 69.820 186.390 70.140 186.450 ;
        RECT 71.660 186.590 71.980 186.650 ;
        RECT 72.135 186.590 72.425 186.635 ;
        RECT 74.420 186.590 74.740 186.650 ;
        RECT 71.660 186.450 74.740 186.590 ;
        RECT 71.660 186.390 71.980 186.450 ;
        RECT 72.135 186.405 72.425 186.450 ;
        RECT 74.420 186.390 74.740 186.450 ;
        RECT 75.800 186.390 76.120 186.650 ;
        RECT 81.290 186.590 81.580 186.635 ;
        RECT 83.610 186.590 83.825 186.745 ;
        RECT 86.840 186.590 87.160 186.650 ;
        RECT 81.290 186.450 83.825 186.590 ;
        RECT 84.170 186.450 87.160 186.590 ;
        RECT 88.770 186.590 88.910 186.790 ;
        RECT 89.715 186.790 93.605 186.930 ;
        RECT 89.715 186.745 90.305 186.790 ;
        RECT 92.955 186.745 93.605 186.790 ;
        RECT 99.275 186.930 99.565 186.975 ;
        RECT 103.055 186.930 103.345 186.975 ;
        RECT 106.295 186.930 106.945 186.975 ;
        RECT 99.275 186.790 106.945 186.930 ;
        RECT 99.275 186.745 99.565 186.790 ;
        RECT 103.055 186.745 103.645 186.790 ;
        RECT 106.295 186.745 106.945 186.790 ;
        RECT 108.935 186.745 109.225 186.975 ;
        RECT 90.015 186.590 90.305 186.745 ;
        RECT 88.770 186.450 90.305 186.590 ;
        RECT 81.290 186.405 81.580 186.450 ;
        RECT 54.640 186.110 58.625 186.250 ;
        RECT 54.640 186.050 54.960 186.110 ;
        RECT 58.335 186.065 58.625 186.110 ;
        RECT 59.790 186.110 63.150 186.250 ;
        RECT 65.695 186.250 65.985 186.295 ;
        RECT 70.740 186.250 71.060 186.310 ;
        RECT 65.695 186.110 71.060 186.250 ;
        RECT 75.890 186.250 76.030 186.390 ;
        RECT 84.170 186.250 84.310 186.450 ;
        RECT 86.840 186.390 87.160 186.450 ;
        RECT 90.015 186.430 90.305 186.450 ;
        RECT 91.095 186.590 91.385 186.635 ;
        RECT 94.675 186.590 94.965 186.635 ;
        RECT 96.510 186.590 96.800 186.635 ;
        RECT 91.095 186.450 96.800 186.590 ;
        RECT 91.095 186.405 91.385 186.450 ;
        RECT 94.675 186.405 94.965 186.450 ;
        RECT 96.510 186.405 96.800 186.450 ;
        RECT 97.435 186.590 97.725 186.635 ;
        RECT 98.815 186.590 99.105 186.635 ;
        RECT 99.720 186.590 100.040 186.650 ;
        RECT 97.435 186.450 100.040 186.590 ;
        RECT 97.435 186.405 97.725 186.450 ;
        RECT 98.815 186.405 99.105 186.450 ;
        RECT 99.720 186.390 100.040 186.450 ;
        RECT 103.355 186.430 103.645 186.745 ;
        RECT 104.435 186.590 104.725 186.635 ;
        RECT 108.015 186.590 108.305 186.635 ;
        RECT 109.850 186.590 110.140 186.635 ;
        RECT 104.435 186.450 110.140 186.590 ;
        RECT 104.435 186.405 104.725 186.450 ;
        RECT 108.015 186.405 108.305 186.450 ;
        RECT 109.850 186.405 110.140 186.450 ;
        RECT 110.775 186.405 111.065 186.635 ;
        RECT 75.890 186.110 84.310 186.250 ;
        RECT 55.575 185.910 55.865 185.955 ;
        RECT 59.790 185.910 59.930 186.110 ;
        RECT 65.695 186.065 65.985 186.110 ;
        RECT 70.740 186.050 71.060 186.110 ;
        RECT 84.540 186.050 84.860 186.310 ;
        RECT 86.395 186.250 86.685 186.295 ;
        RECT 87.300 186.250 87.620 186.310 ;
        RECT 96.975 186.250 97.265 186.295 ;
        RECT 105.240 186.250 105.560 186.310 ;
        RECT 110.300 186.250 110.620 186.310 ;
        RECT 86.395 186.110 110.620 186.250 ;
        RECT 86.395 186.065 86.685 186.110 ;
        RECT 87.300 186.050 87.620 186.110 ;
        RECT 96.975 186.065 97.265 186.110 ;
        RECT 105.240 186.050 105.560 186.110 ;
        RECT 110.300 186.050 110.620 186.110 ;
        RECT 50.130 185.770 55.865 185.910 ;
        RECT 55.575 185.725 55.865 185.770 ;
        RECT 58.870 185.770 59.930 185.910 ;
        RECT 58.870 185.630 59.010 185.770 ;
        RECT 60.160 185.710 60.480 185.970 ;
        RECT 66.600 185.910 66.920 185.970 ;
        RECT 67.535 185.910 67.825 185.955 ;
        RECT 75.340 185.910 75.660 185.970 ;
        RECT 66.600 185.770 67.825 185.910 ;
        RECT 66.600 185.710 66.920 185.770 ;
        RECT 67.535 185.725 67.825 185.770 ;
        RECT 68.070 185.770 75.660 185.910 ;
        RECT 42.680 185.430 46.590 185.570 ;
        RECT 48.215 185.570 48.505 185.615 ;
        RECT 55.100 185.570 55.420 185.630 ;
        RECT 48.215 185.430 55.420 185.570 ;
        RECT 42.680 185.370 43.000 185.430 ;
        RECT 48.215 185.385 48.505 185.430 ;
        RECT 55.100 185.370 55.420 185.430 ;
        RECT 58.780 185.370 59.100 185.630 ;
        RECT 59.700 185.570 60.020 185.630 ;
        RECT 62.015 185.570 62.305 185.615 ;
        RECT 59.700 185.430 62.305 185.570 ;
        RECT 59.700 185.370 60.020 185.430 ;
        RECT 62.015 185.385 62.305 185.430 ;
        RECT 63.840 185.370 64.160 185.630 ;
        RECT 65.220 185.570 65.540 185.630 ;
        RECT 68.070 185.570 68.210 185.770 ;
        RECT 75.340 185.710 75.660 185.770 ;
        RECT 81.290 185.910 81.580 185.955 ;
        RECT 84.070 185.910 84.360 185.955 ;
        RECT 85.930 185.910 86.220 185.955 ;
        RECT 81.290 185.770 86.220 185.910 ;
        RECT 81.290 185.725 81.580 185.770 ;
        RECT 84.070 185.725 84.360 185.770 ;
        RECT 85.930 185.725 86.220 185.770 ;
        RECT 91.095 185.910 91.385 185.955 ;
        RECT 94.215 185.910 94.505 185.955 ;
        RECT 96.105 185.910 96.395 185.955 ;
        RECT 91.095 185.770 96.395 185.910 ;
        RECT 91.095 185.725 91.385 185.770 ;
        RECT 94.215 185.725 94.505 185.770 ;
        RECT 96.105 185.725 96.395 185.770 ;
        RECT 97.880 185.710 98.200 185.970 ;
        RECT 104.435 185.910 104.725 185.955 ;
        RECT 107.555 185.910 107.845 185.955 ;
        RECT 109.445 185.910 109.735 185.955 ;
        RECT 104.435 185.770 109.735 185.910 ;
        RECT 104.435 185.725 104.725 185.770 ;
        RECT 107.555 185.725 107.845 185.770 ;
        RECT 109.445 185.725 109.735 185.770 ;
        RECT 65.220 185.430 68.210 185.570 ;
        RECT 65.220 185.370 65.540 185.430 ;
        RECT 71.200 185.370 71.520 185.630 ;
        RECT 73.515 185.570 73.805 185.615 ;
        RECT 76.720 185.570 77.040 185.630 ;
        RECT 73.515 185.430 77.040 185.570 ;
        RECT 73.515 185.385 73.805 185.430 ;
        RECT 76.720 185.370 77.040 185.430 ;
        RECT 77.425 185.570 77.715 185.615 ;
        RECT 79.480 185.570 79.800 185.630 ;
        RECT 77.425 185.430 79.800 185.570 ;
        RECT 77.425 185.385 77.715 185.430 ;
        RECT 79.480 185.370 79.800 185.430 ;
        RECT 86.380 185.570 86.700 185.630 ;
        RECT 87.760 185.570 88.080 185.630 ;
        RECT 88.235 185.570 88.525 185.615 ;
        RECT 86.380 185.430 88.525 185.570 ;
        RECT 86.380 185.370 86.700 185.430 ;
        RECT 87.760 185.370 88.080 185.430 ;
        RECT 88.235 185.385 88.525 185.430 ;
        RECT 95.690 185.570 95.980 185.615 ;
        RECT 99.260 185.570 99.580 185.630 ;
        RECT 95.690 185.430 99.580 185.570 ;
        RECT 95.690 185.385 95.980 185.430 ;
        RECT 99.260 185.370 99.580 185.430 ;
        RECT 99.720 185.570 100.040 185.630 ;
        RECT 102.020 185.570 102.340 185.630 ;
        RECT 110.850 185.570 110.990 186.405 ;
        RECT 99.720 185.430 110.990 185.570 ;
        RECT 99.720 185.370 100.040 185.430 ;
        RECT 102.020 185.370 102.340 185.430 ;
        RECT 22.830 184.750 113.450 185.230 ;
        RECT 40.380 184.350 40.700 184.610 ;
        RECT 43.600 184.550 43.920 184.610 ;
        RECT 46.835 184.550 47.125 184.595 ;
        RECT 41.850 184.410 43.370 184.550 ;
        RECT 29.455 184.210 29.745 184.255 ;
        RECT 32.575 184.210 32.865 184.255 ;
        RECT 34.465 184.210 34.755 184.255 ;
        RECT 41.850 184.210 41.990 184.410 ;
        RECT 29.455 184.070 34.755 184.210 ;
        RECT 29.455 184.025 29.745 184.070 ;
        RECT 32.575 184.025 32.865 184.070 ;
        RECT 34.465 184.025 34.755 184.070 ;
        RECT 38.170 184.070 41.990 184.210 ;
        RECT 26.580 183.670 26.900 183.930 ;
        RECT 35.320 183.670 35.640 183.930 ;
        RECT 26.135 183.530 26.425 183.575 ;
        RECT 27.500 183.530 27.820 183.590 ;
        RECT 26.135 183.390 27.820 183.530 ;
        RECT 26.135 183.345 26.425 183.390 ;
        RECT 27.500 183.330 27.820 183.390 ;
        RECT 28.375 183.235 28.665 183.550 ;
        RECT 29.455 183.530 29.745 183.575 ;
        RECT 33.035 183.530 33.325 183.575 ;
        RECT 34.870 183.530 35.160 183.575 ;
        RECT 29.455 183.390 35.160 183.530 ;
        RECT 29.455 183.345 29.745 183.390 ;
        RECT 33.035 183.345 33.325 183.390 ;
        RECT 34.870 183.345 35.160 183.390 ;
        RECT 36.700 183.330 37.020 183.590 ;
        RECT 37.620 183.330 37.940 183.590 ;
        RECT 38.170 183.575 38.310 184.070 ;
        RECT 42.220 184.010 42.540 184.270 ;
        RECT 43.230 184.210 43.370 184.410 ;
        RECT 43.600 184.410 47.125 184.550 ;
        RECT 43.600 184.350 43.920 184.410 ;
        RECT 46.835 184.365 47.125 184.410 ;
        RECT 56.020 184.550 56.340 184.610 ;
        RECT 62.475 184.550 62.765 184.595 ;
        RECT 56.020 184.410 62.765 184.550 ;
        RECT 56.020 184.350 56.340 184.410 ;
        RECT 62.475 184.365 62.765 184.410 ;
        RECT 65.220 184.350 65.540 184.610 ;
        RECT 66.140 184.550 66.460 184.610 ;
        RECT 66.615 184.550 66.905 184.595 ;
        RECT 66.140 184.410 66.905 184.550 ;
        RECT 66.140 184.350 66.460 184.410 ;
        RECT 66.615 184.365 66.905 184.410 ;
        RECT 70.740 184.550 71.060 184.610 ;
        RECT 70.740 184.410 71.890 184.550 ;
        RECT 70.740 184.350 71.060 184.410 ;
        RECT 46.360 184.210 46.680 184.270 ;
        RECT 52.800 184.210 53.120 184.270 ;
        RECT 43.230 184.070 53.120 184.210 ;
        RECT 46.360 184.010 46.680 184.070 ;
        RECT 52.800 184.010 53.120 184.070 ;
        RECT 55.215 184.210 55.505 184.255 ;
        RECT 58.335 184.210 58.625 184.255 ;
        RECT 60.225 184.210 60.515 184.255 ;
        RECT 55.215 184.070 60.515 184.210 ;
        RECT 55.215 184.025 55.505 184.070 ;
        RECT 58.335 184.025 58.625 184.070 ;
        RECT 60.225 184.025 60.515 184.070 ;
        RECT 69.820 184.210 70.140 184.270 ;
        RECT 69.820 184.070 71.430 184.210 ;
        RECT 69.820 184.010 70.140 184.070 ;
        RECT 38.095 183.345 38.385 183.575 ;
        RECT 25.675 183.190 25.965 183.235 ;
        RECT 28.075 183.190 28.665 183.235 ;
        RECT 31.315 183.190 31.965 183.235 ;
        RECT 25.675 183.050 31.965 183.190 ;
        RECT 25.675 183.005 25.965 183.050 ;
        RECT 28.075 183.005 28.365 183.050 ;
        RECT 31.315 183.005 31.965 183.050 ;
        RECT 33.955 183.005 34.245 183.235 ;
        RECT 38.170 183.190 38.310 183.345 ;
        RECT 38.540 183.330 38.860 183.590 ;
        RECT 42.310 183.575 42.450 184.010 ;
        RECT 42.695 183.870 42.985 183.915 ;
        RECT 43.140 183.870 43.460 183.930 ;
        RECT 42.695 183.730 43.460 183.870 ;
        RECT 42.695 183.685 42.985 183.730 ;
        RECT 43.140 183.670 43.460 183.730 ;
        RECT 43.600 183.870 43.920 183.930 ;
        RECT 49.595 183.870 49.885 183.915 ;
        RECT 54.640 183.870 54.960 183.930 ;
        RECT 56.020 183.870 56.340 183.930 ;
        RECT 43.600 183.730 56.340 183.870 ;
        RECT 43.600 183.670 43.920 183.730 ;
        RECT 49.595 183.685 49.885 183.730 ;
        RECT 54.640 183.670 54.960 183.730 ;
        RECT 56.020 183.670 56.340 183.730 ;
        RECT 59.700 183.670 60.020 183.930 ;
        RECT 61.080 183.670 61.400 183.930 ;
        RECT 68.900 183.870 69.220 183.930 ;
        RECT 71.290 183.915 71.430 184.070 ;
        RECT 71.750 183.915 71.890 184.410 ;
        RECT 74.420 184.350 74.740 184.610 ;
        RECT 84.540 184.550 84.860 184.610 ;
        RECT 85.935 184.550 86.225 184.595 ;
        RECT 92.820 184.550 93.140 184.610 ;
        RECT 84.540 184.410 86.225 184.550 ;
        RECT 84.540 184.350 84.860 184.410 ;
        RECT 85.935 184.365 86.225 184.410 ;
        RECT 89.690 184.410 99.030 184.550 ;
        RECT 79.955 184.210 80.245 184.255 ;
        RECT 79.955 184.070 87.070 184.210 ;
        RECT 79.955 184.025 80.245 184.070 ;
        RECT 67.610 183.730 70.050 183.870 ;
        RECT 42.235 183.345 42.525 183.575 ;
        RECT 48.675 183.530 48.965 183.575 ;
        RECT 53.260 183.530 53.580 183.590 ;
        RECT 48.675 183.390 53.580 183.530 ;
        RECT 48.675 183.345 48.965 183.390 ;
        RECT 53.260 183.330 53.580 183.390 ;
        RECT 34.950 183.050 38.310 183.190 ;
        RECT 39.460 183.190 39.780 183.250 ;
        RECT 54.135 183.235 54.425 183.550 ;
        RECT 55.215 183.530 55.505 183.575 ;
        RECT 58.795 183.530 59.085 183.575 ;
        RECT 60.630 183.530 60.920 183.575 ;
        RECT 55.215 183.390 60.920 183.530 ;
        RECT 55.215 183.345 55.505 183.390 ;
        RECT 58.795 183.345 59.085 183.390 ;
        RECT 60.630 183.345 60.920 183.390 ;
        RECT 63.855 183.530 64.145 183.575 ;
        RECT 64.300 183.530 64.620 183.590 ;
        RECT 63.855 183.390 64.620 183.530 ;
        RECT 63.855 183.345 64.145 183.390 ;
        RECT 64.300 183.330 64.620 183.390 ;
        RECT 64.760 183.330 65.080 183.590 ;
        RECT 67.610 183.575 67.750 183.730 ;
        RECT 68.900 183.670 69.220 183.730 ;
        RECT 69.910 183.590 70.050 183.730 ;
        RECT 71.215 183.685 71.505 183.915 ;
        RECT 71.675 183.685 71.965 183.915 ;
        RECT 72.120 183.670 72.440 183.930 ;
        RECT 72.580 183.870 72.900 183.930 ;
        RECT 74.895 183.870 75.185 183.915 ;
        RECT 72.580 183.730 75.185 183.870 ;
        RECT 72.580 183.670 72.900 183.730 ;
        RECT 74.895 183.685 75.185 183.730 ;
        RECT 75.340 183.670 75.660 183.930 ;
        RECT 76.720 183.870 77.040 183.930 ;
        RECT 80.875 183.870 81.165 183.915 ;
        RECT 81.320 183.870 81.640 183.930 ;
        RECT 86.380 183.870 86.700 183.930 ;
        RECT 76.720 183.730 81.640 183.870 ;
        RECT 76.720 183.670 77.040 183.730 ;
        RECT 80.875 183.685 81.165 183.730 ;
        RECT 81.320 183.670 81.640 183.730 ;
        RECT 82.330 183.730 86.700 183.870 ;
        RECT 67.535 183.345 67.825 183.575 ;
        RECT 67.980 183.530 68.300 183.590 ;
        RECT 69.375 183.530 69.665 183.575 ;
        RECT 67.980 183.390 69.665 183.530 ;
        RECT 67.980 183.330 68.300 183.390 ;
        RECT 69.375 183.345 69.665 183.390 ;
        RECT 49.135 183.190 49.425 183.235 ;
        RECT 39.460 183.050 49.425 183.190 ;
        RECT 26.120 182.850 26.440 182.910 ;
        RECT 34.030 182.850 34.170 183.005 ;
        RECT 34.950 182.910 35.090 183.050 ;
        RECT 39.460 182.990 39.780 183.050 ;
        RECT 49.135 183.005 49.425 183.050 ;
        RECT 53.835 183.190 54.425 183.235 ;
        RECT 57.075 183.190 57.725 183.235 ;
        RECT 60.160 183.190 60.480 183.250 ;
        RECT 53.835 183.050 60.480 183.190 ;
        RECT 69.450 183.190 69.590 183.345 ;
        RECT 69.820 183.330 70.140 183.590 ;
        RECT 70.740 183.330 71.060 183.590 ;
        RECT 73.500 183.330 73.820 183.590 ;
        RECT 82.330 183.575 82.470 183.730 ;
        RECT 86.380 183.670 86.700 183.730 ;
        RECT 73.975 183.345 74.265 183.575 ;
        RECT 82.255 183.530 82.545 183.575 ;
        RECT 77.270 183.390 82.545 183.530 ;
        RECT 73.040 183.190 73.360 183.250 ;
        RECT 74.050 183.190 74.190 183.345 ;
        RECT 69.450 183.050 74.190 183.190 ;
        RECT 53.835 183.005 54.125 183.050 ;
        RECT 57.075 183.005 57.725 183.050 ;
        RECT 60.160 182.990 60.480 183.050 ;
        RECT 73.040 182.990 73.360 183.050 ;
        RECT 26.120 182.710 34.170 182.850 ;
        RECT 26.120 182.650 26.440 182.710 ;
        RECT 34.860 182.650 35.180 182.910 ;
        RECT 39.920 182.650 40.240 182.910 ;
        RECT 52.340 182.650 52.660 182.910 ;
        RECT 52.800 182.850 53.120 182.910 ;
        RECT 59.700 182.850 60.020 182.910 ;
        RECT 68.455 182.850 68.745 182.895 ;
        RECT 70.740 182.850 71.060 182.910 ;
        RECT 52.800 182.710 71.060 182.850 ;
        RECT 52.800 182.650 53.120 182.710 ;
        RECT 59.700 182.650 60.020 182.710 ;
        RECT 68.455 182.665 68.745 182.710 ;
        RECT 70.740 182.650 71.060 182.710 ;
        RECT 71.660 182.850 71.980 182.910 ;
        RECT 77.270 182.850 77.410 183.390 ;
        RECT 82.255 183.345 82.545 183.390 ;
        RECT 84.540 183.330 84.860 183.590 ;
        RECT 86.930 183.575 87.070 184.070 ;
        RECT 89.690 183.590 89.830 184.410 ;
        RECT 92.820 184.350 93.140 184.410 ;
        RECT 90.060 184.210 90.380 184.270 ;
        RECT 98.890 184.210 99.030 184.410 ;
        RECT 99.260 184.350 99.580 184.610 ;
        RECT 99.810 184.410 102.710 184.550 ;
        RECT 99.810 184.210 99.950 184.410 ;
        RECT 90.060 184.070 95.810 184.210 ;
        RECT 98.890 184.070 99.950 184.210 ;
        RECT 100.180 184.210 100.500 184.270 ;
        RECT 100.180 184.070 102.250 184.210 ;
        RECT 90.060 184.010 90.380 184.070 ;
        RECT 95.120 183.870 95.440 183.930 ;
        RECT 95.670 183.915 95.810 184.070 ;
        RECT 100.180 184.010 100.500 184.070 ;
        RECT 90.150 183.730 95.440 183.870 ;
        RECT 86.855 183.345 87.145 183.575 ;
        RECT 88.680 183.530 89.000 183.590 ;
        RECT 89.155 183.530 89.445 183.575 ;
        RECT 88.680 183.390 89.445 183.530 ;
        RECT 88.680 183.330 89.000 183.390 ;
        RECT 89.155 183.345 89.445 183.390 ;
        RECT 77.655 183.190 77.945 183.235 ;
        RECT 79.480 183.190 79.800 183.250 ;
        RECT 77.655 183.050 79.800 183.190 ;
        RECT 89.230 183.190 89.370 183.345 ;
        RECT 89.600 183.330 89.920 183.590 ;
        RECT 90.150 183.575 90.290 183.730 ;
        RECT 95.120 183.670 95.440 183.730 ;
        RECT 95.595 183.685 95.885 183.915 ;
        RECT 96.500 183.870 96.820 183.930 ;
        RECT 96.500 183.730 100.870 183.870 ;
        RECT 96.500 183.670 96.820 183.730 ;
        RECT 90.075 183.345 90.365 183.575 ;
        RECT 90.995 183.530 91.285 183.575 ;
        RECT 91.440 183.530 91.760 183.590 ;
        RECT 90.995 183.390 91.760 183.530 ;
        RECT 90.995 183.345 91.285 183.390 ;
        RECT 91.440 183.330 91.760 183.390 ;
        RECT 92.375 183.345 92.665 183.575 ;
        RECT 90.520 183.190 90.840 183.250 ;
        RECT 89.230 183.050 90.840 183.190 ;
        RECT 92.450 183.190 92.590 183.345 ;
        RECT 92.820 183.330 93.140 183.590 ;
        RECT 93.280 183.330 93.600 183.590 ;
        RECT 96.040 183.530 96.360 183.590 ;
        RECT 100.195 183.530 100.485 183.575 ;
        RECT 96.040 183.390 100.485 183.530 ;
        RECT 100.730 183.530 100.870 183.730 ;
        RECT 101.560 183.670 101.880 183.930 ;
        RECT 102.110 183.915 102.250 184.070 ;
        RECT 102.035 183.685 102.325 183.915 ;
        RECT 102.570 183.870 102.710 184.410 ;
        RECT 104.320 184.350 104.640 184.610 ;
        RECT 102.940 184.210 103.260 184.270 ;
        RECT 107.080 184.210 107.400 184.270 ;
        RECT 111.680 184.210 112.000 184.270 ;
        RECT 102.940 184.070 107.400 184.210 ;
        RECT 102.940 184.010 103.260 184.070 ;
        RECT 107.080 184.010 107.400 184.070 ;
        RECT 110.850 184.070 112.000 184.210 ;
        RECT 102.570 183.730 110.530 183.870 ;
        RECT 106.710 183.590 106.850 183.730 ;
        RECT 100.730 183.390 105.240 183.530 ;
        RECT 96.040 183.330 96.360 183.390 ;
        RECT 100.195 183.345 100.485 183.390 ;
        RECT 101.100 183.190 101.420 183.250 ;
        RECT 102.495 183.190 102.785 183.235 ;
        RECT 92.450 183.050 102.785 183.190 ;
        RECT 105.100 183.190 105.240 183.390 ;
        RECT 106.160 183.330 106.480 183.590 ;
        RECT 106.620 183.330 106.940 183.590 ;
        RECT 107.080 183.330 107.400 183.590 ;
        RECT 108.015 183.530 108.305 183.575 ;
        RECT 108.920 183.530 109.240 183.590 ;
        RECT 110.390 183.575 110.530 183.730 ;
        RECT 110.850 183.575 110.990 184.070 ;
        RECT 111.680 184.010 112.000 184.070 ;
        RECT 108.015 183.390 109.240 183.530 ;
        RECT 108.015 183.345 108.305 183.390 ;
        RECT 108.920 183.330 109.240 183.390 ;
        RECT 109.855 183.345 110.145 183.575 ;
        RECT 110.315 183.345 110.605 183.575 ;
        RECT 110.775 183.345 111.065 183.575 ;
        RECT 111.695 183.345 111.985 183.575 ;
        RECT 106.250 183.190 106.390 183.330 ;
        RECT 109.930 183.190 110.070 183.345 ;
        RECT 105.100 183.050 105.470 183.190 ;
        RECT 106.250 183.050 110.070 183.190 ;
        RECT 77.655 183.005 77.945 183.050 ;
        RECT 79.480 182.990 79.800 183.050 ;
        RECT 90.520 182.990 90.840 183.050 ;
        RECT 101.100 182.990 101.420 183.050 ;
        RECT 102.495 183.005 102.785 183.050 ;
        RECT 71.660 182.710 77.410 182.850 ;
        RECT 78.100 182.850 78.420 182.910 ;
        RECT 81.795 182.850 82.085 182.895 ;
        RECT 78.100 182.710 82.085 182.850 ;
        RECT 71.660 182.650 71.980 182.710 ;
        RECT 78.100 182.650 78.420 182.710 ;
        RECT 81.795 182.665 82.085 182.710 ;
        RECT 84.080 182.650 84.400 182.910 ;
        RECT 85.475 182.850 85.765 182.895 ;
        RECT 85.920 182.850 86.240 182.910 ;
        RECT 85.475 182.710 86.240 182.850 ;
        RECT 85.475 182.665 85.765 182.710 ;
        RECT 85.920 182.650 86.240 182.710 ;
        RECT 87.775 182.850 88.065 182.895 ;
        RECT 88.680 182.850 89.000 182.910 ;
        RECT 87.775 182.710 89.000 182.850 ;
        RECT 90.610 182.850 90.750 182.990 ;
        RECT 93.280 182.850 93.600 182.910 ;
        RECT 90.610 182.710 93.600 182.850 ;
        RECT 87.775 182.665 88.065 182.710 ;
        RECT 88.680 182.650 89.000 182.710 ;
        RECT 93.280 182.650 93.600 182.710 ;
        RECT 94.675 182.850 94.965 182.895 ;
        RECT 96.500 182.850 96.820 182.910 ;
        RECT 94.675 182.710 96.820 182.850 ;
        RECT 94.675 182.665 94.965 182.710 ;
        RECT 96.500 182.650 96.820 182.710 ;
        RECT 98.355 182.850 98.645 182.895 ;
        RECT 99.720 182.850 100.040 182.910 ;
        RECT 98.355 182.710 100.040 182.850 ;
        RECT 98.355 182.665 98.645 182.710 ;
        RECT 99.720 182.650 100.040 182.710 ;
        RECT 100.640 182.850 100.960 182.910 ;
        RECT 104.795 182.850 105.085 182.895 ;
        RECT 100.640 182.710 105.085 182.850 ;
        RECT 105.330 182.850 105.470 183.050 ;
        RECT 107.080 182.850 107.400 182.910 ;
        RECT 105.330 182.710 107.400 182.850 ;
        RECT 100.640 182.650 100.960 182.710 ;
        RECT 104.795 182.665 105.085 182.710 ;
        RECT 107.080 182.650 107.400 182.710 ;
        RECT 108.460 182.650 108.780 182.910 ;
        RECT 108.920 182.850 109.240 182.910 ;
        RECT 111.770 182.850 111.910 183.345 ;
        RECT 108.920 182.710 111.910 182.850 ;
        RECT 108.920 182.650 109.240 182.710 ;
        RECT 22.830 182.030 113.450 182.510 ;
        RECT 26.120 181.630 26.440 181.890 ;
        RECT 26.595 181.645 26.885 181.875 ;
        RECT 25.215 181.150 25.505 181.195 ;
        RECT 26.670 181.150 26.810 181.645 ;
        RECT 28.420 181.630 28.740 181.890 ;
        RECT 28.880 181.830 29.200 181.890 ;
        RECT 28.880 181.690 34.170 181.830 ;
        RECT 28.880 181.630 29.200 181.690 ;
        RECT 31.660 181.490 31.950 181.535 ;
        RECT 33.520 181.490 33.810 181.535 ;
        RECT 31.660 181.350 33.810 181.490 ;
        RECT 34.030 181.490 34.170 181.690 ;
        RECT 42.680 181.630 43.000 181.890 ;
        RECT 48.215 181.830 48.505 181.875 ;
        RECT 56.480 181.830 56.800 181.890 ;
        RECT 48.215 181.690 56.800 181.830 ;
        RECT 48.215 181.645 48.505 181.690 ;
        RECT 56.480 181.630 56.800 181.690 ;
        RECT 58.780 181.630 59.100 181.890 ;
        RECT 69.835 181.830 70.125 181.875 ;
        RECT 60.250 181.690 70.125 181.830 ;
        RECT 34.440 181.490 34.730 181.535 ;
        RECT 37.700 181.490 37.990 181.535 ;
        RECT 34.030 181.350 37.990 181.490 ;
        RECT 31.660 181.305 31.950 181.350 ;
        RECT 33.520 181.305 33.810 181.350 ;
        RECT 34.440 181.305 34.730 181.350 ;
        RECT 37.700 181.305 37.990 181.350 ;
        RECT 38.540 181.490 38.860 181.550 ;
        RECT 42.770 181.490 42.910 181.630 ;
        RECT 57.400 181.490 57.720 181.550 ;
        RECT 60.250 181.490 60.390 181.690 ;
        RECT 69.835 181.645 70.125 181.690 ;
        RECT 70.740 181.830 71.060 181.890 ;
        RECT 72.120 181.830 72.440 181.890 ;
        RECT 70.740 181.690 72.440 181.830 ;
        RECT 38.540 181.350 60.390 181.490 ;
        RECT 60.735 181.490 61.025 181.535 ;
        RECT 62.920 181.490 63.240 181.550 ;
        RECT 63.975 181.490 64.625 181.535 ;
        RECT 60.735 181.350 64.625 181.490 ;
        RECT 25.215 181.010 26.810 181.150 ;
        RECT 32.100 181.150 32.420 181.210 ;
        RECT 32.575 181.150 32.865 181.195 ;
        RECT 32.100 181.010 32.865 181.150 ;
        RECT 33.595 181.150 33.810 181.305 ;
        RECT 38.540 181.290 38.860 181.350 ;
        RECT 35.840 181.150 36.130 181.195 ;
        RECT 33.595 181.010 36.130 181.150 ;
        RECT 25.215 180.965 25.505 181.010 ;
        RECT 32.100 180.950 32.420 181.010 ;
        RECT 32.575 180.965 32.865 181.010 ;
        RECT 35.840 180.965 36.130 181.010 ;
        RECT 36.700 181.150 37.020 181.210 ;
        RECT 41.300 181.150 41.620 181.210 ;
        RECT 36.700 181.010 41.620 181.150 ;
        RECT 36.700 180.950 37.020 181.010 ;
        RECT 41.300 180.950 41.620 181.010 ;
        RECT 41.760 181.150 42.080 181.210 ;
        RECT 43.230 181.195 43.370 181.350 ;
        RECT 42.235 181.150 42.525 181.195 ;
        RECT 41.760 181.010 42.525 181.150 ;
        RECT 41.760 180.950 42.080 181.010 ;
        RECT 42.235 180.965 42.525 181.010 ;
        RECT 42.695 180.965 42.985 181.195 ;
        RECT 43.155 180.965 43.445 181.195 ;
        RECT 49.580 181.150 49.900 181.210 ;
        RECT 44.610 181.010 49.900 181.150 ;
        RECT 28.420 180.810 28.740 180.870 ;
        RECT 28.895 180.810 29.185 180.855 ;
        RECT 28.420 180.670 29.185 180.810 ;
        RECT 28.420 180.610 28.740 180.670 ;
        RECT 28.895 180.625 29.185 180.670 ;
        RECT 29.815 180.810 30.105 180.855 ;
        RECT 30.260 180.810 30.580 180.870 ;
        RECT 29.815 180.670 30.580 180.810 ;
        RECT 29.815 180.625 30.105 180.670 ;
        RECT 30.260 180.610 30.580 180.670 ;
        RECT 30.735 180.810 31.025 180.855 ;
        RECT 35.320 180.810 35.640 180.870 ;
        RECT 42.770 180.810 42.910 180.965 ;
        RECT 44.610 180.855 44.750 181.010 ;
        RECT 49.580 180.950 49.900 181.010 ;
        RECT 50.040 180.950 50.360 181.210 ;
        RECT 51.435 181.150 51.725 181.195 ;
        RECT 51.880 181.150 52.200 181.210 ;
        RECT 51.435 181.010 52.200 181.150 ;
        RECT 51.435 180.965 51.725 181.010 ;
        RECT 51.880 180.950 52.200 181.010 ;
        RECT 52.340 180.950 52.660 181.210 ;
        RECT 52.800 180.950 53.120 181.210 ;
        RECT 53.350 181.195 53.490 181.350 ;
        RECT 57.400 181.290 57.720 181.350 ;
        RECT 60.735 181.305 61.325 181.350 ;
        RECT 53.275 180.965 53.565 181.195 ;
        RECT 56.940 180.950 57.260 181.210 ;
        RECT 61.035 180.990 61.325 181.305 ;
        RECT 62.920 181.290 63.240 181.350 ;
        RECT 63.975 181.305 64.625 181.350 ;
        RECT 69.910 181.490 70.050 181.645 ;
        RECT 70.740 181.630 71.060 181.690 ;
        RECT 72.120 181.630 72.440 181.690 ;
        RECT 78.100 181.630 78.420 181.890 ;
        RECT 90.980 181.830 91.300 181.890 ;
        RECT 97.895 181.830 98.185 181.875 ;
        RECT 100.655 181.830 100.945 181.875 ;
        RECT 106.160 181.830 106.480 181.890 ;
        RECT 90.980 181.690 100.945 181.830 ;
        RECT 90.980 181.630 91.300 181.690 ;
        RECT 97.895 181.645 98.185 181.690 ;
        RECT 100.655 181.645 100.945 181.690 ;
        RECT 101.190 181.690 106.480 181.830 ;
        RECT 73.975 181.490 74.265 181.535 ;
        RECT 75.340 181.490 75.660 181.550 ;
        RECT 83.620 181.535 83.940 181.550 ;
        RECT 69.910 181.350 72.810 181.490 ;
        RECT 62.115 181.150 62.405 181.195 ;
        RECT 65.695 181.150 65.985 181.195 ;
        RECT 67.530 181.150 67.820 181.195 ;
        RECT 62.115 181.010 67.820 181.150 ;
        RECT 62.115 180.965 62.405 181.010 ;
        RECT 65.695 180.965 65.985 181.010 ;
        RECT 67.530 180.965 67.820 181.010 ;
        RECT 68.900 180.950 69.220 181.210 ;
        RECT 30.735 180.670 35.640 180.810 ;
        RECT 30.735 180.625 31.025 180.670 ;
        RECT 35.320 180.610 35.640 180.670 ;
        RECT 36.330 180.670 42.910 180.810 ;
        RECT 31.200 180.470 31.490 180.515 ;
        RECT 33.060 180.470 33.350 180.515 ;
        RECT 35.840 180.470 36.130 180.515 ;
        RECT 31.200 180.330 36.130 180.470 ;
        RECT 31.200 180.285 31.490 180.330 ;
        RECT 33.060 180.285 33.350 180.330 ;
        RECT 35.840 180.285 36.130 180.330 ;
        RECT 29.340 180.130 29.660 180.190 ;
        RECT 34.860 180.130 35.180 180.190 ;
        RECT 36.330 180.130 36.470 180.670 ;
        RECT 44.535 180.625 44.825 180.855 ;
        RECT 45.455 180.810 45.745 180.855 ;
        RECT 52.430 180.810 52.570 180.950 ;
        RECT 45.455 180.670 52.570 180.810 ;
        RECT 45.455 180.625 45.745 180.670 ;
        RECT 54.640 180.610 54.960 180.870 ;
        RECT 56.020 180.810 56.340 180.870 ;
        RECT 58.320 180.810 58.640 180.870 ;
        RECT 56.020 180.670 58.640 180.810 ;
        RECT 56.020 180.610 56.340 180.670 ;
        RECT 58.320 180.610 58.640 180.670 ;
        RECT 61.540 180.810 61.860 180.870 ;
        RECT 67.995 180.810 68.285 180.855 ;
        RECT 61.540 180.670 68.285 180.810 ;
        RECT 61.540 180.610 61.860 180.670 ;
        RECT 67.995 180.625 68.285 180.670 ;
        RECT 62.115 180.470 62.405 180.515 ;
        RECT 65.235 180.470 65.525 180.515 ;
        RECT 67.125 180.470 67.415 180.515 ;
        RECT 62.115 180.330 67.415 180.470 ;
        RECT 69.910 180.470 70.050 181.350 ;
        RECT 70.740 180.950 71.060 181.210 ;
        RECT 71.660 180.950 71.980 181.210 ;
        RECT 72.120 180.950 72.440 181.210 ;
        RECT 72.670 181.195 72.810 181.350 ;
        RECT 73.975 181.350 75.660 181.490 ;
        RECT 73.975 181.305 74.265 181.350 ;
        RECT 75.340 181.290 75.660 181.350 ;
        RECT 80.055 181.490 80.345 181.535 ;
        RECT 83.295 181.490 83.945 181.535 ;
        RECT 80.055 181.350 83.945 181.490 ;
        RECT 80.055 181.305 80.645 181.350 ;
        RECT 83.295 181.305 83.945 181.350 ;
        RECT 72.595 181.150 72.885 181.195 ;
        RECT 74.420 181.150 74.740 181.210 ;
        RECT 72.595 181.010 74.740 181.150 ;
        RECT 72.595 180.965 72.885 181.010 ;
        RECT 74.420 180.950 74.740 181.010 ;
        RECT 74.970 181.010 80.170 181.150 ;
        RECT 70.280 180.810 70.600 180.870 ;
        RECT 74.970 180.810 75.110 181.010 ;
        RECT 70.280 180.670 75.110 180.810 ;
        RECT 75.355 180.810 75.645 180.855 ;
        RECT 76.260 180.810 76.580 180.870 ;
        RECT 78.575 180.810 78.865 180.855 ;
        RECT 75.355 180.670 78.865 180.810 ;
        RECT 80.030 180.810 80.170 181.010 ;
        RECT 80.355 180.990 80.645 181.305 ;
        RECT 83.620 181.290 83.940 181.305 ;
        RECT 85.920 181.290 86.240 181.550 ;
        RECT 91.440 181.490 91.760 181.550 ;
        RECT 101.190 181.490 101.330 181.690 ;
        RECT 88.310 181.350 91.760 181.490 ;
        RECT 88.310 181.195 88.450 181.350 ;
        RECT 91.440 181.290 91.760 181.350 ;
        RECT 94.750 181.350 101.330 181.490 ;
        RECT 81.435 181.150 81.725 181.195 ;
        RECT 85.015 181.150 85.305 181.195 ;
        RECT 86.850 181.150 87.140 181.195 ;
        RECT 88.235 181.150 88.525 181.195 ;
        RECT 81.435 181.010 87.140 181.150 ;
        RECT 81.435 180.965 81.725 181.010 ;
        RECT 85.015 180.965 85.305 181.010 ;
        RECT 86.850 180.965 87.140 181.010 ;
        RECT 87.850 181.010 88.525 181.150 ;
        RECT 80.030 180.670 87.070 180.810 ;
        RECT 70.280 180.610 70.600 180.670 ;
        RECT 75.355 180.625 75.645 180.670 ;
        RECT 76.260 180.610 76.580 180.670 ;
        RECT 78.575 180.625 78.865 180.670 ;
        RECT 71.660 180.470 71.980 180.530 ;
        RECT 69.910 180.330 71.980 180.470 ;
        RECT 62.115 180.285 62.405 180.330 ;
        RECT 65.235 180.285 65.525 180.330 ;
        RECT 67.125 180.285 67.415 180.330 ;
        RECT 71.660 180.270 71.980 180.330 ;
        RECT 81.435 180.470 81.725 180.515 ;
        RECT 84.555 180.470 84.845 180.515 ;
        RECT 86.445 180.470 86.735 180.515 ;
        RECT 81.435 180.330 86.735 180.470 ;
        RECT 86.930 180.470 87.070 180.670 ;
        RECT 87.300 180.610 87.620 180.870 ;
        RECT 87.850 180.470 87.990 181.010 ;
        RECT 88.235 180.965 88.525 181.010 ;
        RECT 89.140 180.950 89.460 181.210 ;
        RECT 89.600 180.950 89.920 181.210 ;
        RECT 90.075 181.150 90.365 181.195 ;
        RECT 90.520 181.150 90.840 181.210 ;
        RECT 94.750 181.150 94.890 181.350 ;
        RECT 104.320 181.290 104.640 181.550 ;
        RECT 90.075 181.010 94.890 181.150 ;
        RECT 95.120 181.150 95.440 181.210 ;
        RECT 105.790 181.195 105.930 181.690 ;
        RECT 106.160 181.630 106.480 181.690 ;
        RECT 106.620 181.630 106.940 181.890 ;
        RECT 111.220 181.630 111.540 181.890 ;
        RECT 106.710 181.490 106.850 181.630 ;
        RECT 106.250 181.350 106.850 181.490 ;
        RECT 106.250 181.195 106.390 181.350 ;
        RECT 103.415 181.150 103.705 181.195 ;
        RECT 95.120 181.010 103.705 181.150 ;
        RECT 90.075 180.965 90.365 181.010 ;
        RECT 90.520 180.950 90.840 181.010 ;
        RECT 95.120 180.950 95.440 181.010 ;
        RECT 103.415 180.965 103.705 181.010 ;
        RECT 105.715 180.965 106.005 181.195 ;
        RECT 106.175 180.965 106.465 181.195 ;
        RECT 106.635 181.150 106.925 181.195 ;
        RECT 107.080 181.150 107.400 181.210 ;
        RECT 106.635 181.010 107.400 181.150 ;
        RECT 106.635 180.965 106.925 181.010 ;
        RECT 107.080 180.950 107.400 181.010 ;
        RECT 107.555 181.150 107.845 181.195 ;
        RECT 108.920 181.150 109.240 181.210 ;
        RECT 107.555 181.010 109.240 181.150 ;
        RECT 107.555 180.965 107.845 181.010 ;
        RECT 108.920 180.950 109.240 181.010 ;
        RECT 89.690 180.810 89.830 180.950 ;
        RECT 86.930 180.330 87.990 180.470 ;
        RECT 88.310 180.670 89.830 180.810 ;
        RECT 91.455 180.810 91.745 180.855 ;
        RECT 91.900 180.810 92.220 180.870 ;
        RECT 91.455 180.670 92.220 180.810 ;
        RECT 81.435 180.285 81.725 180.330 ;
        RECT 84.555 180.285 84.845 180.330 ;
        RECT 86.445 180.285 86.735 180.330 ;
        RECT 29.340 179.990 36.470 180.130 ;
        RECT 39.460 180.175 39.780 180.190 ;
        RECT 29.340 179.930 29.660 179.990 ;
        RECT 34.860 179.930 35.180 179.990 ;
        RECT 39.460 179.945 39.995 180.175 ;
        RECT 50.975 180.130 51.265 180.175 ;
        RECT 51.880 180.130 52.200 180.190 ;
        RECT 50.975 179.990 52.200 180.130 ;
        RECT 50.975 179.945 51.265 179.990 ;
        RECT 39.460 179.930 39.780 179.945 ;
        RECT 51.880 179.930 52.200 179.990 ;
        RECT 57.860 180.130 58.180 180.190 ;
        RECT 59.255 180.130 59.545 180.175 ;
        RECT 60.160 180.130 60.480 180.190 ;
        RECT 57.860 179.990 60.480 180.130 ;
        RECT 57.860 179.930 58.180 179.990 ;
        RECT 59.255 179.945 59.545 179.990 ;
        RECT 60.160 179.930 60.480 179.990 ;
        RECT 64.760 180.130 65.080 180.190 ;
        RECT 66.680 180.130 66.970 180.175 ;
        RECT 64.760 179.990 66.970 180.130 ;
        RECT 64.760 179.930 65.080 179.990 ;
        RECT 66.680 179.945 66.970 179.990 ;
        RECT 69.820 180.130 70.140 180.190 ;
        RECT 88.310 180.130 88.450 180.670 ;
        RECT 91.455 180.625 91.745 180.670 ;
        RECT 91.900 180.610 92.220 180.670 ;
        RECT 92.835 180.810 93.125 180.855 ;
        RECT 95.580 180.810 95.900 180.870 ;
        RECT 92.835 180.670 95.900 180.810 ;
        RECT 92.835 180.625 93.125 180.670 ;
        RECT 95.580 180.610 95.900 180.670 ;
        RECT 96.515 180.625 96.805 180.855 ;
        RECT 97.435 180.810 97.725 180.855 ;
        RECT 108.015 180.810 108.305 180.855 ;
        RECT 97.435 180.670 98.110 180.810 ;
        RECT 97.435 180.625 97.725 180.670 ;
        RECT 94.660 180.470 94.980 180.530 ;
        RECT 96.590 180.470 96.730 180.625 ;
        RECT 94.660 180.330 96.730 180.470 ;
        RECT 94.660 180.270 94.980 180.330 ;
        RECT 69.820 179.990 88.450 180.130 ;
        RECT 95.595 180.130 95.885 180.175 ;
        RECT 97.420 180.130 97.740 180.190 ;
        RECT 95.595 179.990 97.740 180.130 ;
        RECT 97.970 180.130 98.110 180.670 ;
        RECT 99.810 180.670 108.305 180.810 ;
        RECT 99.810 180.515 99.950 180.670 ;
        RECT 108.015 180.625 108.305 180.670 ;
        RECT 99.735 180.285 100.025 180.515 ;
        RECT 103.400 180.130 103.720 180.190 ;
        RECT 97.970 179.990 103.720 180.130 ;
        RECT 69.820 179.930 70.140 179.990 ;
        RECT 95.595 179.945 95.885 179.990 ;
        RECT 97.420 179.930 97.740 179.990 ;
        RECT 103.400 179.930 103.720 179.990 ;
        RECT 22.830 179.310 113.450 179.790 ;
        RECT 31.180 178.910 31.500 179.170 ;
        RECT 38.540 179.110 38.860 179.170 ;
        RECT 36.790 178.970 38.860 179.110 ;
        RECT 36.790 178.770 36.930 178.970 ;
        RECT 38.540 178.910 38.860 178.970 ;
        RECT 39.920 179.110 40.240 179.170 ;
        RECT 43.140 179.110 43.460 179.170 ;
        RECT 50.040 179.110 50.360 179.170 ;
        RECT 39.920 178.970 43.460 179.110 ;
        RECT 39.920 178.910 40.240 178.970 ;
        RECT 43.140 178.910 43.460 178.970 ;
        RECT 46.910 178.970 50.360 179.110 ;
        RECT 41.760 178.770 42.080 178.830 ;
        RECT 29.890 178.630 36.930 178.770 ;
        RECT 37.250 178.630 42.080 178.770 ;
        RECT 24.755 178.430 25.045 178.475 ;
        RECT 26.580 178.430 26.900 178.490 ;
        RECT 24.755 178.290 29.110 178.430 ;
        RECT 24.755 178.245 25.045 178.290 ;
        RECT 26.580 178.230 26.900 178.290 ;
        RECT 27.960 177.890 28.280 178.150 ;
        RECT 28.970 178.135 29.110 178.290 ;
        RECT 28.895 177.905 29.185 178.135 ;
        RECT 29.340 177.890 29.660 178.150 ;
        RECT 29.890 178.135 30.030 178.630 ;
        RECT 30.260 178.430 30.580 178.490 ;
        RECT 37.250 178.475 37.390 178.630 ;
        RECT 41.760 178.570 42.080 178.630 ;
        RECT 44.075 178.770 44.365 178.815 ;
        RECT 46.910 178.770 47.050 178.970 ;
        RECT 50.040 178.910 50.360 178.970 ;
        RECT 62.475 179.110 62.765 179.155 ;
        RECT 62.920 179.110 63.240 179.170 ;
        RECT 62.475 178.970 63.240 179.110 ;
        RECT 62.475 178.925 62.765 178.970 ;
        RECT 62.920 178.910 63.240 178.970 ;
        RECT 64.760 178.910 65.080 179.170 ;
        RECT 67.060 179.110 67.380 179.170 ;
        RECT 69.820 179.110 70.140 179.170 ;
        RECT 67.060 178.970 70.140 179.110 ;
        RECT 67.060 178.910 67.380 178.970 ;
        RECT 69.820 178.910 70.140 178.970 ;
        RECT 72.120 179.110 72.440 179.170 ;
        RECT 75.800 179.110 76.120 179.170 ;
        RECT 72.120 178.970 80.170 179.110 ;
        RECT 72.120 178.910 72.440 178.970 ;
        RECT 75.800 178.910 76.120 178.970 ;
        RECT 44.075 178.630 47.050 178.770 ;
        RECT 47.395 178.770 47.685 178.815 ;
        RECT 50.515 178.770 50.805 178.815 ;
        RECT 52.405 178.770 52.695 178.815 ;
        RECT 47.395 178.630 52.695 178.770 ;
        RECT 44.075 178.585 44.365 178.630 ;
        RECT 47.395 178.585 47.685 178.630 ;
        RECT 50.515 178.585 50.805 178.630 ;
        RECT 52.405 178.585 52.695 178.630 ;
        RECT 56.940 178.770 57.260 178.830 ;
        RECT 61.095 178.770 61.385 178.815 ;
        RECT 61.540 178.770 61.860 178.830 ;
        RECT 56.940 178.630 59.010 178.770 ;
        RECT 56.940 178.570 57.260 178.630 ;
        RECT 34.415 178.430 34.705 178.475 ;
        RECT 30.260 178.290 34.705 178.430 ;
        RECT 30.260 178.230 30.580 178.290 ;
        RECT 34.415 178.245 34.705 178.290 ;
        RECT 37.175 178.245 37.465 178.475 ;
        RECT 40.855 178.430 41.145 178.475 ;
        RECT 43.600 178.430 43.920 178.490 ;
        RECT 39.550 178.290 43.920 178.430 ;
        RECT 29.815 177.905 30.105 178.135 ;
        RECT 31.640 178.090 31.960 178.150 ;
        RECT 33.955 178.090 34.245 178.135 ;
        RECT 31.640 177.950 34.245 178.090 ;
        RECT 34.490 178.090 34.630 178.245 ;
        RECT 38.080 178.090 38.400 178.150 ;
        RECT 39.550 178.090 39.690 178.290 ;
        RECT 40.855 178.245 41.145 178.290 ;
        RECT 43.600 178.230 43.920 178.290 ;
        RECT 51.880 178.230 52.200 178.490 ;
        RECT 54.195 178.430 54.485 178.475 ;
        RECT 57.860 178.430 58.180 178.490 ;
        RECT 54.195 178.290 58.180 178.430 ;
        RECT 54.195 178.245 54.485 178.290 ;
        RECT 57.860 178.230 58.180 178.290 ;
        RECT 58.320 178.230 58.640 178.490 ;
        RECT 58.870 178.475 59.010 178.630 ;
        RECT 61.095 178.630 61.860 178.770 ;
        RECT 61.095 178.585 61.385 178.630 ;
        RECT 61.540 178.570 61.860 178.630 ;
        RECT 62.000 178.770 62.320 178.830 ;
        RECT 68.915 178.770 69.205 178.815 ;
        RECT 70.740 178.770 71.060 178.830 ;
        RECT 79.480 178.770 79.800 178.830 ;
        RECT 62.000 178.630 71.060 178.770 ;
        RECT 62.000 178.570 62.320 178.630 ;
        RECT 68.915 178.585 69.205 178.630 ;
        RECT 70.740 178.570 71.060 178.630 ;
        RECT 72.670 178.630 79.800 178.770 ;
        RECT 58.795 178.245 59.085 178.475 ;
        RECT 65.220 178.430 65.540 178.490 ;
        RECT 65.220 178.290 70.050 178.430 ;
        RECT 65.220 178.230 65.540 178.290 ;
        RECT 69.910 178.150 70.050 178.290 ;
        RECT 34.490 177.950 39.690 178.090 ;
        RECT 39.935 178.090 40.225 178.135 ;
        RECT 41.775 178.090 42.065 178.135 ;
        RECT 39.935 177.950 42.065 178.090 ;
        RECT 31.640 177.890 31.960 177.950 ;
        RECT 33.955 177.905 34.245 177.950 ;
        RECT 27.515 177.750 27.805 177.795 ;
        RECT 28.420 177.750 28.740 177.810 ;
        RECT 33.495 177.750 33.785 177.795 ;
        RECT 27.515 177.610 33.785 177.750 ;
        RECT 34.030 177.750 34.170 177.905 ;
        RECT 38.080 177.890 38.400 177.950 ;
        RECT 39.935 177.905 40.225 177.950 ;
        RECT 41.775 177.905 42.065 177.950 ;
        RECT 39.460 177.750 39.780 177.810 ;
        RECT 42.235 177.750 42.525 177.795 ;
        RECT 34.030 177.610 42.525 177.750 ;
        RECT 27.515 177.565 27.805 177.610 ;
        RECT 28.420 177.550 28.740 177.610 ;
        RECT 33.495 177.565 33.785 177.610 ;
        RECT 39.460 177.550 39.780 177.610 ;
        RECT 42.235 177.565 42.525 177.610 ;
        RECT 43.600 177.750 43.920 177.810 ;
        RECT 46.315 177.795 46.605 178.110 ;
        RECT 47.395 178.090 47.685 178.135 ;
        RECT 50.975 178.090 51.265 178.135 ;
        RECT 52.810 178.090 53.100 178.135 ;
        RECT 47.395 177.950 53.100 178.090 ;
        RECT 47.395 177.905 47.685 177.950 ;
        RECT 50.975 177.905 51.265 177.950 ;
        RECT 52.810 177.905 53.100 177.950 ;
        RECT 53.275 178.090 53.565 178.135 ;
        RECT 56.940 178.090 57.260 178.150 ;
        RECT 60.620 178.090 60.940 178.150 ;
        RECT 62.935 178.090 63.225 178.135 ;
        RECT 53.275 177.950 60.390 178.090 ;
        RECT 53.275 177.905 53.565 177.950 ;
        RECT 56.940 177.890 57.260 177.950 ;
        RECT 46.015 177.750 46.605 177.795 ;
        RECT 49.255 177.750 49.905 177.795 ;
        RECT 60.250 177.750 60.390 177.950 ;
        RECT 60.620 177.950 63.225 178.090 ;
        RECT 60.620 177.890 60.940 177.950 ;
        RECT 62.935 177.905 63.225 177.950 ;
        RECT 63.855 178.090 64.145 178.135 ;
        RECT 64.760 178.090 65.080 178.150 ;
        RECT 63.855 177.950 65.080 178.090 ;
        RECT 63.855 177.905 64.145 177.950 ;
        RECT 64.760 177.890 65.080 177.950 ;
        RECT 67.980 177.890 68.300 178.150 ;
        RECT 69.820 177.890 70.140 178.150 ;
        RECT 71.660 177.890 71.980 178.150 ;
        RECT 72.120 177.890 72.440 178.150 ;
        RECT 72.670 178.135 72.810 178.630 ;
        RECT 79.480 178.570 79.800 178.630 ;
        RECT 80.030 178.430 80.170 178.970 ;
        RECT 84.540 178.910 84.860 179.170 ;
        RECT 95.580 178.910 95.900 179.170 ;
        RECT 110.300 179.110 110.620 179.170 ;
        RECT 110.300 178.970 111.910 179.110 ;
        RECT 110.300 178.910 110.620 178.970 ;
        RECT 83.620 178.770 83.940 178.830 ;
        RECT 85.475 178.770 85.765 178.815 ;
        RECT 105.815 178.770 106.105 178.815 ;
        RECT 108.935 178.770 109.225 178.815 ;
        RECT 110.825 178.770 111.115 178.815 ;
        RECT 83.620 178.630 85.765 178.770 ;
        RECT 83.620 178.570 83.940 178.630 ;
        RECT 85.475 178.585 85.765 178.630 ;
        RECT 90.150 178.630 101.790 178.770 ;
        RECT 75.430 178.290 79.250 178.430 ;
        RECT 72.595 177.905 72.885 178.135 ;
        RECT 73.515 177.905 73.805 178.135 ;
        RECT 74.420 178.090 74.740 178.150 ;
        RECT 75.430 178.135 75.570 178.290 ;
        RECT 75.355 178.090 75.645 178.135 ;
        RECT 74.420 177.950 75.645 178.090 ;
        RECT 61.080 177.750 61.400 177.810 ;
        RECT 43.600 177.610 49.905 177.750 ;
        RECT 43.600 177.550 43.920 177.610 ;
        RECT 46.015 177.565 46.305 177.610 ;
        RECT 49.255 177.565 49.905 177.610 ;
        RECT 50.130 177.610 56.940 177.750 ;
        RECT 60.250 177.610 61.400 177.750 ;
        RECT 26.580 177.410 26.900 177.470 ;
        RECT 31.655 177.410 31.945 177.455 ;
        RECT 26.580 177.270 31.945 177.410 ;
        RECT 26.580 177.210 26.900 177.270 ;
        RECT 31.655 177.225 31.945 177.270 ;
        RECT 41.760 177.410 42.080 177.470 ;
        RECT 44.535 177.410 44.825 177.455 ;
        RECT 50.130 177.410 50.270 177.610 ;
        RECT 41.760 177.270 50.270 177.410 ;
        RECT 56.800 177.410 56.940 177.610 ;
        RECT 61.080 177.550 61.400 177.610 ;
        RECT 70.740 177.750 71.060 177.810 ;
        RECT 73.590 177.750 73.730 177.905 ;
        RECT 74.420 177.890 74.740 177.950 ;
        RECT 75.355 177.905 75.645 177.950 ;
        RECT 75.800 177.890 76.120 178.150 ;
        RECT 76.260 177.890 76.580 178.150 ;
        RECT 79.110 178.135 79.250 178.290 ;
        RECT 79.570 178.290 80.170 178.430 ;
        RECT 81.795 178.430 82.085 178.475 ;
        RECT 84.080 178.430 84.400 178.490 ;
        RECT 81.795 178.290 84.400 178.430 ;
        RECT 79.570 178.135 79.710 178.290 ;
        RECT 81.795 178.245 82.085 178.290 ;
        RECT 84.080 178.230 84.400 178.290 ;
        RECT 77.195 177.905 77.485 178.135 ;
        RECT 79.035 177.905 79.325 178.135 ;
        RECT 79.495 177.905 79.785 178.135 ;
        RECT 79.955 178.090 80.245 178.135 ;
        RECT 80.400 178.090 80.720 178.150 ;
        RECT 79.955 177.950 80.720 178.090 ;
        RECT 79.955 177.905 80.245 177.950 ;
        RECT 77.270 177.750 77.410 177.905 ;
        RECT 80.400 177.890 80.720 177.950 ;
        RECT 80.875 177.905 81.165 178.135 ;
        RECT 85.935 178.090 86.225 178.135 ;
        RECT 86.380 178.090 86.700 178.150 ;
        RECT 87.760 178.090 88.080 178.150 ;
        RECT 90.150 178.090 90.290 178.630 ;
        RECT 97.895 178.430 98.185 178.475 ;
        RECT 90.610 178.290 98.185 178.430 ;
        RECT 90.610 178.150 90.750 178.290 ;
        RECT 97.895 178.245 98.185 178.290 ;
        RECT 98.355 178.245 98.645 178.475 ;
        RECT 85.935 177.950 90.290 178.090 ;
        RECT 85.935 177.905 86.225 177.950 ;
        RECT 80.950 177.750 81.090 177.905 ;
        RECT 86.380 177.890 86.700 177.950 ;
        RECT 87.760 177.890 88.080 177.950 ;
        RECT 90.520 177.890 90.840 178.150 ;
        RECT 93.755 178.090 94.045 178.135 ;
        RECT 91.070 177.950 94.045 178.090 ;
        RECT 70.740 177.610 81.090 177.750 ;
        RECT 85.000 177.750 85.320 177.810 ;
        RECT 91.070 177.750 91.210 177.950 ;
        RECT 93.755 177.905 94.045 177.950 ;
        RECT 94.660 178.090 94.980 178.150 ;
        RECT 98.430 178.090 98.570 178.245 ;
        RECT 94.660 177.950 98.570 178.090 ;
        RECT 94.660 177.890 94.980 177.950 ;
        RECT 100.180 177.890 100.500 178.150 ;
        RECT 101.650 178.135 101.790 178.630 ;
        RECT 105.815 178.630 111.115 178.770 ;
        RECT 105.815 178.585 106.105 178.630 ;
        RECT 108.935 178.585 109.225 178.630 ;
        RECT 110.825 178.585 111.115 178.630 ;
        RECT 111.770 178.475 111.910 178.970 ;
        RECT 111.695 178.245 111.985 178.475 ;
        RECT 101.575 178.090 101.865 178.135 ;
        RECT 102.020 178.090 102.340 178.150 ;
        RECT 101.575 177.950 102.340 178.090 ;
        RECT 101.575 177.905 101.865 177.950 ;
        RECT 102.020 177.890 102.340 177.950 ;
        RECT 85.000 177.610 91.210 177.750 ;
        RECT 93.295 177.750 93.585 177.795 ;
        RECT 96.040 177.750 96.360 177.810 ;
        RECT 93.295 177.610 96.360 177.750 ;
        RECT 70.740 177.550 71.060 177.610 ;
        RECT 85.000 177.550 85.320 177.610 ;
        RECT 93.295 177.565 93.585 177.610 ;
        RECT 96.040 177.550 96.360 177.610 ;
        RECT 97.880 177.750 98.200 177.810 ;
        RECT 104.735 177.795 105.025 178.110 ;
        RECT 105.815 178.090 106.105 178.135 ;
        RECT 109.395 178.090 109.685 178.135 ;
        RECT 111.230 178.090 111.520 178.135 ;
        RECT 105.815 177.950 111.520 178.090 ;
        RECT 105.815 177.905 106.105 177.950 ;
        RECT 109.395 177.905 109.685 177.950 ;
        RECT 111.230 177.905 111.520 177.950 ;
        RECT 104.435 177.750 105.025 177.795 ;
        RECT 107.675 177.750 108.325 177.795 ;
        RECT 97.880 177.610 108.325 177.750 ;
        RECT 97.880 177.550 98.200 177.610 ;
        RECT 104.435 177.565 104.725 177.610 ;
        RECT 107.675 177.565 108.325 177.610 ;
        RECT 110.315 177.750 110.605 177.795 ;
        RECT 110.760 177.750 111.080 177.810 ;
        RECT 110.315 177.610 111.080 177.750 ;
        RECT 110.315 177.565 110.605 177.610 ;
        RECT 110.760 177.550 111.080 177.610 ;
        RECT 59.255 177.410 59.545 177.455 ;
        RECT 56.800 177.270 59.545 177.410 ;
        RECT 41.760 177.210 42.080 177.270 ;
        RECT 44.535 177.225 44.825 177.270 ;
        RECT 59.255 177.225 59.545 177.270 ;
        RECT 68.900 177.410 69.220 177.470 ;
        RECT 70.295 177.410 70.585 177.455 ;
        RECT 68.900 177.270 70.585 177.410 ;
        RECT 68.900 177.210 69.220 177.270 ;
        RECT 70.295 177.225 70.585 177.270 ;
        RECT 73.960 177.210 74.280 177.470 ;
        RECT 74.880 177.410 75.200 177.470 ;
        RECT 77.655 177.410 77.945 177.455 ;
        RECT 74.880 177.270 77.945 177.410 ;
        RECT 74.880 177.210 75.200 177.270 ;
        RECT 77.655 177.225 77.945 177.270 ;
        RECT 88.220 177.210 88.540 177.470 ;
        RECT 94.675 177.410 94.965 177.455 ;
        RECT 96.960 177.410 97.280 177.470 ;
        RECT 94.675 177.270 97.280 177.410 ;
        RECT 94.675 177.225 94.965 177.270 ;
        RECT 96.960 177.210 97.280 177.270 ;
        RECT 97.435 177.410 97.725 177.455 ;
        RECT 99.720 177.410 100.040 177.470 ;
        RECT 97.435 177.270 100.040 177.410 ;
        RECT 97.435 177.225 97.725 177.270 ;
        RECT 99.720 177.210 100.040 177.270 ;
        RECT 101.100 177.210 101.420 177.470 ;
        RECT 102.020 177.210 102.340 177.470 ;
        RECT 102.955 177.410 103.245 177.455 ;
        RECT 103.400 177.410 103.720 177.470 ;
        RECT 102.955 177.270 103.720 177.410 ;
        RECT 102.955 177.225 103.245 177.270 ;
        RECT 103.400 177.210 103.720 177.270 ;
        RECT 22.830 176.590 113.450 177.070 ;
        RECT 28.435 176.390 28.725 176.435 ;
        RECT 28.880 176.390 29.200 176.450 ;
        RECT 35.780 176.390 36.100 176.450 ;
        RECT 41.760 176.390 42.080 176.450 ;
        RECT 28.435 176.250 29.200 176.390 ;
        RECT 28.435 176.205 28.725 176.250 ;
        RECT 28.880 176.190 29.200 176.250 ;
        RECT 32.650 176.250 42.080 176.390 ;
        RECT 32.650 175.770 32.790 176.250 ;
        RECT 35.780 176.190 36.100 176.250 ;
        RECT 41.760 176.190 42.080 176.250 ;
        RECT 42.235 176.205 42.525 176.435 ;
        RECT 42.680 176.390 43.000 176.450 ;
        RECT 42.680 176.250 64.530 176.390 ;
        RECT 33.480 176.050 33.800 176.110 ;
        RECT 34.515 176.050 34.805 176.095 ;
        RECT 37.755 176.050 38.405 176.095 ;
        RECT 33.480 175.910 38.405 176.050 ;
        RECT 33.480 175.850 33.800 175.910 ;
        RECT 34.515 175.865 35.105 175.910 ;
        RECT 37.755 175.865 38.405 175.910 ;
        RECT 40.395 176.050 40.685 176.095 ;
        RECT 42.310 176.050 42.450 176.205 ;
        RECT 42.680 176.190 43.000 176.250 ;
        RECT 40.395 175.910 42.450 176.050 ;
        RECT 52.340 176.050 52.660 176.110 ;
        RECT 62.000 176.050 62.320 176.110 ;
        RECT 52.340 175.910 62.320 176.050 ;
        RECT 64.390 176.050 64.530 176.250 ;
        RECT 64.760 176.190 65.080 176.450 ;
        RECT 68.455 176.390 68.745 176.435 ;
        RECT 70.280 176.390 70.600 176.450 ;
        RECT 68.455 176.250 70.600 176.390 ;
        RECT 68.455 176.205 68.745 176.250 ;
        RECT 68.530 176.050 68.670 176.205 ;
        RECT 70.280 176.190 70.600 176.250 ;
        RECT 89.615 176.390 89.905 176.435 ;
        RECT 95.120 176.390 95.440 176.450 ;
        RECT 89.615 176.250 95.440 176.390 ;
        RECT 89.615 176.205 89.905 176.250 ;
        RECT 95.120 176.190 95.440 176.250 ;
        RECT 88.220 176.050 88.540 176.110 ;
        RECT 91.095 176.050 91.385 176.095 ;
        RECT 94.335 176.050 94.985 176.095 ;
        RECT 64.390 175.910 68.670 176.050 ;
        RECT 69.450 175.910 70.510 176.050 ;
        RECT 40.395 175.865 40.685 175.910 ;
        RECT 26.580 175.510 26.900 175.770 ;
        RECT 27.960 175.510 28.280 175.770 ;
        RECT 29.800 175.710 30.120 175.770 ;
        RECT 30.735 175.710 31.025 175.755 ;
        RECT 29.800 175.570 31.025 175.710 ;
        RECT 29.800 175.510 30.120 175.570 ;
        RECT 30.735 175.525 31.025 175.570 ;
        RECT 31.195 175.525 31.485 175.755 ;
        RECT 31.270 175.370 31.410 175.525 ;
        RECT 31.640 175.510 31.960 175.770 ;
        RECT 32.560 175.510 32.880 175.770 ;
        RECT 34.815 175.550 35.105 175.865 ;
        RECT 52.340 175.850 52.660 175.910 ;
        RECT 35.895 175.710 36.185 175.755 ;
        RECT 39.475 175.710 39.765 175.755 ;
        RECT 41.310 175.710 41.600 175.755 ;
        RECT 35.895 175.570 41.600 175.710 ;
        RECT 35.895 175.525 36.185 175.570 ;
        RECT 39.475 175.525 39.765 175.570 ;
        RECT 41.310 175.525 41.600 175.570 ;
        RECT 42.680 175.710 43.000 175.770 ;
        RECT 43.155 175.710 43.445 175.755 ;
        RECT 42.680 175.570 43.445 175.710 ;
        RECT 42.680 175.510 43.000 175.570 ;
        RECT 43.155 175.525 43.445 175.570 ;
        RECT 44.520 175.510 44.840 175.770 ;
        RECT 44.980 175.510 45.300 175.770 ;
        RECT 45.900 175.510 46.220 175.770 ;
        RECT 46.360 175.510 46.680 175.770 ;
        RECT 46.820 175.510 47.140 175.770 ;
        RECT 49.580 175.710 49.900 175.770 ;
        RECT 50.055 175.710 50.345 175.755 ;
        RECT 49.580 175.570 50.345 175.710 ;
        RECT 49.580 175.510 49.900 175.570 ;
        RECT 50.055 175.525 50.345 175.570 ;
        RECT 50.500 175.510 50.820 175.770 ;
        RECT 55.115 175.710 55.405 175.755 ;
        RECT 56.940 175.710 57.260 175.770 ;
        RECT 55.115 175.570 57.260 175.710 ;
        RECT 55.115 175.525 55.405 175.570 ;
        RECT 56.940 175.510 57.260 175.570 ;
        RECT 57.400 175.710 57.720 175.770 ;
        RECT 59.255 175.710 59.545 175.755 ;
        RECT 57.400 175.570 59.545 175.710 ;
        RECT 57.400 175.510 57.720 175.570 ;
        RECT 59.255 175.525 59.545 175.570 ;
        RECT 59.700 175.510 60.020 175.770 ;
        RECT 60.160 175.510 60.480 175.770 ;
        RECT 61.170 175.755 61.310 175.910 ;
        RECT 62.000 175.850 62.320 175.910 ;
        RECT 61.095 175.525 61.385 175.755 ;
        RECT 61.540 175.510 61.860 175.770 ;
        RECT 69.450 175.755 69.590 175.910 ;
        RECT 70.370 175.770 70.510 175.910 ;
        RECT 88.220 175.910 94.985 176.050 ;
        RECT 88.220 175.850 88.540 175.910 ;
        RECT 91.095 175.865 91.685 175.910 ;
        RECT 94.335 175.865 94.985 175.910 ;
        RECT 69.375 175.525 69.665 175.755 ;
        RECT 69.835 175.525 70.125 175.755 ;
        RECT 70.280 175.710 70.600 175.770 ;
        RECT 71.675 175.710 71.965 175.755 ;
        RECT 70.280 175.570 71.965 175.710 ;
        RECT 35.320 175.370 35.640 175.430 ;
        RECT 41.775 175.370 42.065 175.415 ;
        RECT 67.060 175.370 67.380 175.430 ;
        RECT 31.270 175.230 32.790 175.370 ;
        RECT 27.515 175.030 27.805 175.075 ;
        RECT 32.100 175.030 32.420 175.090 ;
        RECT 27.515 174.890 32.420 175.030 ;
        RECT 32.650 175.030 32.790 175.230 ;
        RECT 35.320 175.230 42.065 175.370 ;
        RECT 35.320 175.170 35.640 175.230 ;
        RECT 41.775 175.185 42.065 175.230 ;
        RECT 42.310 175.230 67.380 175.370 ;
        RECT 35.895 175.030 36.185 175.075 ;
        RECT 39.015 175.030 39.305 175.075 ;
        RECT 40.905 175.030 41.195 175.075 ;
        RECT 32.650 174.890 35.550 175.030 ;
        RECT 27.515 174.845 27.805 174.890 ;
        RECT 32.100 174.830 32.420 174.890 ;
        RECT 29.355 174.690 29.645 174.735 ;
        RECT 30.720 174.690 31.040 174.750 ;
        RECT 29.355 174.550 31.040 174.690 ;
        RECT 29.355 174.505 29.645 174.550 ;
        RECT 30.720 174.490 31.040 174.550 ;
        RECT 33.035 174.690 33.325 174.735 ;
        RECT 34.860 174.690 35.180 174.750 ;
        RECT 33.035 174.550 35.180 174.690 ;
        RECT 35.410 174.690 35.550 174.890 ;
        RECT 35.895 174.890 41.195 175.030 ;
        RECT 35.895 174.845 36.185 174.890 ;
        RECT 39.015 174.845 39.305 174.890 ;
        RECT 40.905 174.845 41.195 174.890 ;
        RECT 37.160 174.690 37.480 174.750 ;
        RECT 42.310 174.690 42.450 175.230 ;
        RECT 67.060 175.170 67.380 175.230 ;
        RECT 68.440 175.370 68.760 175.430 ;
        RECT 69.910 175.370 70.050 175.525 ;
        RECT 70.280 175.510 70.600 175.570 ;
        RECT 71.675 175.525 71.965 175.570 ;
        RECT 74.420 175.710 74.740 175.770 ;
        RECT 77.195 175.710 77.485 175.755 ;
        RECT 74.420 175.570 77.485 175.710 ;
        RECT 74.420 175.510 74.740 175.570 ;
        RECT 77.195 175.525 77.485 175.570 ;
        RECT 78.575 175.710 78.865 175.755 ;
        RECT 79.955 175.710 80.245 175.755 ;
        RECT 78.575 175.570 80.245 175.710 ;
        RECT 78.575 175.525 78.865 175.570 ;
        RECT 79.955 175.525 80.245 175.570 ;
        RECT 68.440 175.230 70.050 175.370 ;
        RECT 71.215 175.370 71.505 175.415 ;
        RECT 72.580 175.370 72.900 175.430 ;
        RECT 71.215 175.230 72.900 175.370 ;
        RECT 80.030 175.370 80.170 175.525 ;
        RECT 80.400 175.510 80.720 175.770 ;
        RECT 91.395 175.550 91.685 175.865 ;
        RECT 96.960 175.850 97.280 176.110 ;
        RECT 97.420 176.050 97.740 176.110 ;
        RECT 101.100 176.050 101.420 176.110 ;
        RECT 104.335 176.050 104.625 176.095 ;
        RECT 97.420 175.910 99.950 176.050 ;
        RECT 97.420 175.850 97.740 175.910 ;
        RECT 92.475 175.710 92.765 175.755 ;
        RECT 96.055 175.710 96.345 175.755 ;
        RECT 97.890 175.710 98.180 175.755 ;
        RECT 92.475 175.570 98.180 175.710 ;
        RECT 92.475 175.525 92.765 175.570 ;
        RECT 96.055 175.525 96.345 175.570 ;
        RECT 97.890 175.525 98.180 175.570 ;
        RECT 98.340 175.510 98.660 175.770 ;
        RECT 99.810 175.755 99.950 175.910 ;
        RECT 101.100 175.910 104.625 176.050 ;
        RECT 101.100 175.850 101.420 175.910 ;
        RECT 104.335 175.865 104.625 175.910 ;
        RECT 106.615 176.050 107.265 176.095 ;
        RECT 110.215 176.050 110.505 176.095 ;
        RECT 106.615 175.910 110.505 176.050 ;
        RECT 106.615 175.865 107.265 175.910 ;
        RECT 109.915 175.865 110.505 175.910 ;
        RECT 109.915 175.770 110.205 175.865 ;
        RECT 99.735 175.525 100.025 175.755 ;
        RECT 101.560 175.510 101.880 175.770 ;
        RECT 103.420 175.710 103.710 175.755 ;
        RECT 105.255 175.710 105.545 175.755 ;
        RECT 108.835 175.710 109.125 175.755 ;
        RECT 103.420 175.570 109.125 175.710 ;
        RECT 103.420 175.525 103.710 175.570 ;
        RECT 105.255 175.525 105.545 175.570 ;
        RECT 108.835 175.525 109.125 175.570 ;
        RECT 109.840 175.550 110.205 175.770 ;
        RECT 109.840 175.510 110.160 175.550 ;
        RECT 88.220 175.370 88.540 175.430 ;
        RECT 80.030 175.230 88.540 175.370 ;
        RECT 98.430 175.370 98.570 175.510 ;
        RECT 102.940 175.370 103.260 175.430 ;
        RECT 98.430 175.230 103.260 175.370 ;
        RECT 68.440 175.170 68.760 175.230 ;
        RECT 71.215 175.185 71.505 175.230 ;
        RECT 72.580 175.170 72.900 175.230 ;
        RECT 88.220 175.170 88.540 175.230 ;
        RECT 102.940 175.170 103.260 175.230 ;
        RECT 45.440 175.030 45.760 175.090 ;
        RECT 48.215 175.030 48.505 175.075 ;
        RECT 45.440 174.890 48.505 175.030 ;
        RECT 45.440 174.830 45.760 174.890 ;
        RECT 48.215 174.845 48.505 174.890 ;
        RECT 67.520 175.030 67.840 175.090 ;
        RECT 70.280 175.030 70.600 175.090 ;
        RECT 67.520 174.890 70.600 175.030 ;
        RECT 67.520 174.830 67.840 174.890 ;
        RECT 70.280 174.830 70.600 174.890 ;
        RECT 72.120 175.030 72.440 175.090 ;
        RECT 78.115 175.030 78.405 175.075 ;
        RECT 72.120 174.890 78.405 175.030 ;
        RECT 72.120 174.830 72.440 174.890 ;
        RECT 78.115 174.845 78.405 174.890 ;
        RECT 92.475 175.030 92.765 175.075 ;
        RECT 95.595 175.030 95.885 175.075 ;
        RECT 97.485 175.030 97.775 175.075 ;
        RECT 92.475 174.890 97.775 175.030 ;
        RECT 92.475 174.845 92.765 174.890 ;
        RECT 95.595 174.845 95.885 174.890 ;
        RECT 97.485 174.845 97.775 174.890 ;
        RECT 103.825 175.030 104.115 175.075 ;
        RECT 105.715 175.030 106.005 175.075 ;
        RECT 108.835 175.030 109.125 175.075 ;
        RECT 103.825 174.890 109.125 175.030 ;
        RECT 103.825 174.845 104.115 174.890 ;
        RECT 105.715 174.845 106.005 174.890 ;
        RECT 108.835 174.845 109.125 174.890 ;
        RECT 35.410 174.550 42.450 174.690 ;
        RECT 33.035 174.505 33.325 174.550 ;
        RECT 34.860 174.490 35.180 174.550 ;
        RECT 37.160 174.490 37.480 174.550 ;
        RECT 44.060 174.490 44.380 174.750 ;
        RECT 46.820 174.690 47.140 174.750 ;
        RECT 49.135 174.690 49.425 174.735 ;
        RECT 46.820 174.550 49.425 174.690 ;
        RECT 46.820 174.490 47.140 174.550 ;
        RECT 49.135 174.505 49.425 174.550 ;
        RECT 50.960 174.490 51.280 174.750 ;
        RECT 57.875 174.690 58.165 174.735 ;
        RECT 58.320 174.690 58.640 174.750 ;
        RECT 57.875 174.550 58.640 174.690 ;
        RECT 57.875 174.505 58.165 174.550 ;
        RECT 58.320 174.490 58.640 174.550 ;
        RECT 69.820 174.690 70.140 174.750 ;
        RECT 70.755 174.690 71.045 174.735 ;
        RECT 69.820 174.550 71.045 174.690 ;
        RECT 69.820 174.490 70.140 174.550 ;
        RECT 70.755 174.505 71.045 174.550 ;
        RECT 73.960 174.690 74.280 174.750 ;
        RECT 76.275 174.690 76.565 174.735 ;
        RECT 73.960 174.550 76.565 174.690 ;
        RECT 73.960 174.490 74.280 174.550 ;
        RECT 76.275 174.505 76.565 174.550 ;
        RECT 79.480 174.490 79.800 174.750 ;
        RECT 86.840 174.490 87.160 174.750 ;
        RECT 98.800 174.490 99.120 174.750 ;
        RECT 102.495 174.690 102.785 174.735 ;
        RECT 104.320 174.690 104.640 174.750 ;
        RECT 102.495 174.550 104.640 174.690 ;
        RECT 102.495 174.505 102.785 174.550 ;
        RECT 104.320 174.490 104.640 174.550 ;
        RECT 110.760 174.690 111.080 174.750 ;
        RECT 111.695 174.690 111.985 174.735 ;
        RECT 110.760 174.550 111.985 174.690 ;
        RECT 135.635 174.550 136.775 223.880 ;
        RECT 138.130 223.810 139.580 225.110 ;
        RECT 143.180 223.840 144.630 225.140 ;
        RECT 110.760 174.490 111.080 174.550 ;
        RECT 111.695 174.505 111.985 174.550 ;
        RECT 22.830 173.870 113.450 174.350 ;
        RECT 27.960 173.670 28.280 173.730 ;
        RECT 44.520 173.670 44.840 173.730 ;
        RECT 50.500 173.670 50.820 173.730 ;
        RECT 27.960 173.530 50.820 173.670 ;
        RECT 27.960 173.470 28.280 173.530 ;
        RECT 44.520 173.470 44.840 173.530 ;
        RECT 50.500 173.470 50.820 173.530 ;
        RECT 90.060 173.670 90.380 173.730 ;
        RECT 90.060 173.530 91.670 173.670 ;
        RECT 90.060 173.470 90.380 173.530 ;
        RECT 27.515 173.330 27.805 173.375 ;
        RECT 33.480 173.330 33.800 173.390 ;
        RECT 27.515 173.190 33.800 173.330 ;
        RECT 27.515 173.145 27.805 173.190 ;
        RECT 33.480 173.130 33.800 173.190 ;
        RECT 33.940 173.330 34.260 173.390 ;
        RECT 56.480 173.330 56.800 173.390 ;
        RECT 62.475 173.330 62.765 173.375 ;
        RECT 33.940 173.190 62.765 173.330 ;
        RECT 33.940 173.130 34.260 173.190 ;
        RECT 56.480 173.130 56.800 173.190 ;
        RECT 62.475 173.145 62.765 173.190 ;
        RECT 64.760 173.330 65.080 173.390 ;
        RECT 65.680 173.330 66.000 173.390 ;
        RECT 64.760 173.190 66.000 173.330 ;
        RECT 64.760 173.130 65.080 173.190 ;
        RECT 65.680 173.130 66.000 173.190 ;
        RECT 70.710 173.330 71.000 173.375 ;
        RECT 73.490 173.330 73.780 173.375 ;
        RECT 75.350 173.330 75.640 173.375 ;
        RECT 70.710 173.190 75.640 173.330 ;
        RECT 70.710 173.145 71.000 173.190 ;
        RECT 73.490 173.145 73.780 173.190 ;
        RECT 75.350 173.145 75.640 173.190 ;
        RECT 89.140 173.330 89.460 173.390 ;
        RECT 90.150 173.330 90.290 173.470 ;
        RECT 89.140 173.190 90.290 173.330 ;
        RECT 90.520 173.330 90.840 173.390 ;
        RECT 90.995 173.330 91.285 173.375 ;
        RECT 90.520 173.190 91.285 173.330 ;
        RECT 91.530 173.330 91.670 173.530 ;
        RECT 135.580 173.430 136.830 174.550 ;
        RECT 135.635 173.420 136.775 173.430 ;
        RECT 93.855 173.330 94.145 173.375 ;
        RECT 96.975 173.330 97.265 173.375 ;
        RECT 98.865 173.330 99.155 173.375 ;
        RECT 91.530 173.190 93.510 173.330 ;
        RECT 89.140 173.130 89.460 173.190 ;
        RECT 90.520 173.130 90.840 173.190 ;
        RECT 90.995 173.145 91.285 173.190 ;
        RECT 28.895 172.990 29.185 173.035 ;
        RECT 34.860 172.990 35.180 173.050 ;
        RECT 25.290 172.850 27.730 172.990 ;
        RECT 25.290 172.695 25.430 172.850 ;
        RECT 25.215 172.465 25.505 172.695 ;
        RECT 25.660 172.450 25.980 172.710 ;
        RECT 27.055 172.465 27.345 172.695 ;
        RECT 27.590 172.650 27.730 172.850 ;
        RECT 28.895 172.850 35.180 172.990 ;
        RECT 28.895 172.805 29.185 172.850 ;
        RECT 34.860 172.790 35.180 172.850 ;
        RECT 35.320 172.990 35.640 173.050 ;
        RECT 36.255 172.990 36.545 173.035 ;
        RECT 60.620 172.990 60.940 173.050 ;
        RECT 66.600 172.990 66.920 173.050 ;
        RECT 35.320 172.850 36.545 172.990 ;
        RECT 35.320 172.790 35.640 172.850 ;
        RECT 36.255 172.805 36.545 172.850 ;
        RECT 46.450 172.850 66.920 172.990 ;
        RECT 29.800 172.650 30.120 172.710 ;
        RECT 27.590 172.510 30.120 172.650 ;
        RECT 27.130 172.310 27.270 172.465 ;
        RECT 29.800 172.450 30.120 172.510 ;
        RECT 31.640 172.450 31.960 172.710 ;
        RECT 32.115 172.650 32.405 172.695 ;
        RECT 32.560 172.650 32.880 172.710 ;
        RECT 32.115 172.510 32.880 172.650 ;
        RECT 32.115 172.465 32.405 172.510 ;
        RECT 32.560 172.450 32.880 172.510 ;
        RECT 33.035 172.465 33.325 172.695 ;
        RECT 33.495 172.465 33.785 172.695 ;
        RECT 33.955 172.650 34.245 172.695 ;
        RECT 37.620 172.650 37.940 172.710 ;
        RECT 33.955 172.510 37.940 172.650 ;
        RECT 33.955 172.465 34.245 172.510 ;
        RECT 27.960 172.310 28.280 172.370 ;
        RECT 27.130 172.170 28.280 172.310 ;
        RECT 27.960 172.110 28.280 172.170 ;
        RECT 28.880 172.310 29.200 172.370 ;
        RECT 33.110 172.310 33.250 172.465 ;
        RECT 28.880 172.170 33.250 172.310 ;
        RECT 33.570 172.310 33.710 172.465 ;
        RECT 37.620 172.450 37.940 172.510 ;
        RECT 43.600 172.650 43.920 172.710 ;
        RECT 46.450 172.695 46.590 172.850 ;
        RECT 60.620 172.790 60.940 172.850 ;
        RECT 66.600 172.790 66.920 172.850 ;
        RECT 73.960 172.790 74.280 173.050 ;
        RECT 88.235 172.990 88.525 173.035 ;
        RECT 93.370 172.990 93.510 173.190 ;
        RECT 93.855 173.190 99.155 173.330 ;
        RECT 93.855 173.145 94.145 173.190 ;
        RECT 96.975 173.145 97.265 173.190 ;
        RECT 98.865 173.145 99.155 173.190 ;
        RECT 103.055 173.330 103.345 173.375 ;
        RECT 106.175 173.330 106.465 173.375 ;
        RECT 108.065 173.330 108.355 173.375 ;
        RECT 103.055 173.190 108.355 173.330 ;
        RECT 103.055 173.145 103.345 173.190 ;
        RECT 106.175 173.145 106.465 173.190 ;
        RECT 108.065 173.145 108.355 173.190 ;
        RECT 100.195 172.990 100.485 173.035 ;
        RECT 88.235 172.850 93.050 172.990 ;
        RECT 93.370 172.850 100.485 172.990 ;
        RECT 88.235 172.805 88.525 172.850 ;
        RECT 45.915 172.650 46.205 172.695 ;
        RECT 43.600 172.510 46.205 172.650 ;
        RECT 43.600 172.450 43.920 172.510 ;
        RECT 45.915 172.465 46.205 172.510 ;
        RECT 46.375 172.465 46.665 172.695 ;
        RECT 50.500 172.650 50.820 172.710 ;
        RECT 51.880 172.650 52.200 172.710 ;
        RECT 60.160 172.650 60.480 172.710 ;
        RECT 50.500 172.510 60.480 172.650 ;
        RECT 50.500 172.450 50.820 172.510 ;
        RECT 51.880 172.450 52.200 172.510 ;
        RECT 60.160 172.450 60.480 172.510 ;
        RECT 63.395 172.650 63.685 172.695 ;
        RECT 65.220 172.650 65.540 172.710 ;
        RECT 63.395 172.510 65.540 172.650 ;
        RECT 63.395 172.465 63.685 172.510 ;
        RECT 65.220 172.450 65.540 172.510 ;
        RECT 70.710 172.650 71.000 172.695 ;
        RECT 75.815 172.650 76.105 172.695 ;
        RECT 83.620 172.650 83.940 172.710 ;
        RECT 85.935 172.650 86.225 172.695 ;
        RECT 86.840 172.650 87.160 172.710 ;
        RECT 70.710 172.510 73.245 172.650 ;
        RECT 70.710 172.465 71.000 172.510 ;
        RECT 37.160 172.310 37.480 172.370 ;
        RECT 44.520 172.310 44.840 172.370 ;
        RECT 33.570 172.170 44.840 172.310 ;
        RECT 28.880 172.110 29.200 172.170 ;
        RECT 37.160 172.110 37.480 172.170 ;
        RECT 44.520 172.110 44.840 172.170 ;
        RECT 44.995 172.310 45.285 172.355 ;
        RECT 46.820 172.310 47.140 172.370 ;
        RECT 44.995 172.170 47.140 172.310 ;
        RECT 44.995 172.125 45.285 172.170 ;
        RECT 46.820 172.110 47.140 172.170 ;
        RECT 55.575 172.310 55.865 172.355 ;
        RECT 56.940 172.310 57.260 172.370 ;
        RECT 55.575 172.170 57.260 172.310 ;
        RECT 55.575 172.125 55.865 172.170 ;
        RECT 56.940 172.110 57.260 172.170 ;
        RECT 65.680 172.110 66.000 172.370 ;
        RECT 72.120 172.355 72.440 172.370 ;
        RECT 68.850 172.310 69.140 172.355 ;
        RECT 72.110 172.310 72.440 172.355 ;
        RECT 68.850 172.170 72.440 172.310 ;
        RECT 68.850 172.125 69.140 172.170 ;
        RECT 72.110 172.125 72.440 172.170 ;
        RECT 73.030 172.355 73.245 172.510 ;
        RECT 75.815 172.510 87.160 172.650 ;
        RECT 75.815 172.465 76.105 172.510 ;
        RECT 83.620 172.450 83.940 172.510 ;
        RECT 85.935 172.465 86.225 172.510 ;
        RECT 86.840 172.450 87.160 172.510 ;
        RECT 87.760 172.450 88.080 172.710 ;
        RECT 89.155 172.650 89.445 172.695 ;
        RECT 92.910 172.670 93.050 172.850 ;
        RECT 100.195 172.805 100.485 172.850 ;
        RECT 102.480 172.990 102.800 173.050 ;
        RECT 107.555 172.990 107.845 173.035 ;
        RECT 102.480 172.850 107.845 172.990 ;
        RECT 102.480 172.790 102.800 172.850 ;
        RECT 107.555 172.805 107.845 172.850 ;
        RECT 88.310 172.510 89.445 172.650 ;
        RECT 73.030 172.310 73.320 172.355 ;
        RECT 74.890 172.310 75.180 172.355 ;
        RECT 73.030 172.170 75.180 172.310 ;
        RECT 73.030 172.125 73.320 172.170 ;
        RECT 74.890 172.125 75.180 172.170 ;
        RECT 72.120 172.110 72.440 172.125 ;
        RECT 24.755 171.970 25.045 172.015 ;
        RECT 25.200 171.970 25.520 172.030 ;
        RECT 24.755 171.830 25.520 171.970 ;
        RECT 24.755 171.785 25.045 171.830 ;
        RECT 25.200 171.770 25.520 171.830 ;
        RECT 26.595 171.970 26.885 172.015 ;
        RECT 32.100 171.970 32.420 172.030 ;
        RECT 26.595 171.830 32.420 171.970 ;
        RECT 26.595 171.785 26.885 171.830 ;
        RECT 32.100 171.770 32.420 171.830 ;
        RECT 35.335 171.970 35.625 172.015 ;
        RECT 42.220 171.970 42.540 172.030 ;
        RECT 35.335 171.830 42.540 171.970 ;
        RECT 35.335 171.785 35.625 171.830 ;
        RECT 42.220 171.770 42.540 171.830 ;
        RECT 43.600 171.970 43.920 172.030 ;
        RECT 59.240 171.970 59.560 172.030 ;
        RECT 43.600 171.830 59.560 171.970 ;
        RECT 43.600 171.770 43.920 171.830 ;
        RECT 59.240 171.770 59.560 171.830 ;
        RECT 60.620 171.770 60.940 172.030 ;
        RECT 66.845 171.970 67.135 172.015 ;
        RECT 71.660 171.970 71.980 172.030 ;
        RECT 66.845 171.830 71.980 171.970 ;
        RECT 86.930 171.970 87.070 172.450 ;
        RECT 88.310 172.370 88.450 172.510 ;
        RECT 89.155 172.465 89.445 172.510 ;
        RECT 88.220 172.110 88.540 172.370 ;
        RECT 89.615 172.310 89.905 172.355 ;
        RECT 90.060 172.310 90.380 172.370 ;
        RECT 92.775 172.355 93.065 172.670 ;
        RECT 93.855 172.650 94.145 172.695 ;
        RECT 97.435 172.650 97.725 172.695 ;
        RECT 99.270 172.650 99.560 172.695 ;
        RECT 93.855 172.510 99.560 172.650 ;
        RECT 93.855 172.465 94.145 172.510 ;
        RECT 97.435 172.465 97.725 172.510 ;
        RECT 99.270 172.465 99.560 172.510 ;
        RECT 99.735 172.465 100.025 172.695 ;
        RECT 102.020 172.670 102.340 172.710 ;
        RECT 89.615 172.170 90.380 172.310 ;
        RECT 89.615 172.125 89.905 172.170 ;
        RECT 90.060 172.110 90.380 172.170 ;
        RECT 92.475 172.310 93.065 172.355 ;
        RECT 95.715 172.310 96.365 172.355 ;
        RECT 92.475 172.170 96.365 172.310 ;
        RECT 92.475 172.125 92.765 172.170 ;
        RECT 95.715 172.125 96.365 172.170 ;
        RECT 98.355 172.310 98.645 172.355 ;
        RECT 98.800 172.310 99.120 172.370 ;
        RECT 98.355 172.170 99.120 172.310 ;
        RECT 98.355 172.125 98.645 172.170 ;
        RECT 98.800 172.110 99.120 172.170 ;
        RECT 99.810 171.970 99.950 172.465 ;
        RECT 101.975 172.450 102.340 172.670 ;
        RECT 103.055 172.650 103.345 172.695 ;
        RECT 106.635 172.650 106.925 172.695 ;
        RECT 108.470 172.650 108.760 172.695 ;
        RECT 103.055 172.510 108.760 172.650 ;
        RECT 103.055 172.465 103.345 172.510 ;
        RECT 106.635 172.465 106.925 172.510 ;
        RECT 108.470 172.465 108.760 172.510 ;
        RECT 108.935 172.650 109.225 172.695 ;
        RECT 111.220 172.650 111.540 172.710 ;
        RECT 108.935 172.510 111.540 172.650 ;
        RECT 108.935 172.465 109.225 172.510 ;
        RECT 101.975 172.355 102.265 172.450 ;
        RECT 101.675 172.310 102.265 172.355 ;
        RECT 104.915 172.310 105.565 172.355 ;
        RECT 101.675 172.170 105.565 172.310 ;
        RECT 101.675 172.125 101.965 172.170 ;
        RECT 104.915 172.125 105.565 172.170 ;
        RECT 86.930 171.830 99.950 171.970 ;
        RECT 102.940 171.970 103.260 172.030 ;
        RECT 109.010 171.970 109.150 172.465 ;
        RECT 111.220 172.450 111.540 172.510 ;
        RECT 111.680 172.450 112.000 172.710 ;
        RECT 110.300 172.110 110.620 172.370 ;
        RECT 133.700 172.190 134.930 172.680 ;
        RECT 102.940 171.830 109.150 171.970 ;
        RECT 133.700 171.930 136.690 172.190 ;
        RECT 138.330 171.930 139.470 223.810 ;
        RECT 66.845 171.785 67.135 171.830 ;
        RECT 71.660 171.770 71.980 171.830 ;
        RECT 102.940 171.770 103.260 171.830 ;
        RECT 22.830 171.150 113.450 171.630 ;
        RECT 35.780 170.950 36.100 171.010 ;
        RECT 31.270 170.810 36.100 170.950 ;
        RECT 27.450 170.610 27.740 170.655 ;
        RECT 30.710 170.610 31.000 170.655 ;
        RECT 31.270 170.610 31.410 170.810 ;
        RECT 35.780 170.750 36.100 170.810 ;
        RECT 36.240 170.950 36.560 171.010 ;
        RECT 44.980 170.950 45.300 171.010 ;
        RECT 36.240 170.810 45.300 170.950 ;
        RECT 36.240 170.750 36.560 170.810 ;
        RECT 44.980 170.750 45.300 170.810 ;
        RECT 52.340 170.950 52.660 171.010 ;
        RECT 69.820 170.950 70.140 171.010 ;
        RECT 52.340 170.810 59.470 170.950 ;
        RECT 52.340 170.750 52.660 170.810 ;
        RECT 44.060 170.655 44.380 170.670 ;
        RECT 27.450 170.470 31.410 170.610 ;
        RECT 31.630 170.610 31.920 170.655 ;
        RECT 33.490 170.610 33.780 170.655 ;
        RECT 31.630 170.470 33.780 170.610 ;
        RECT 27.450 170.425 27.740 170.470 ;
        RECT 30.710 170.425 31.000 170.470 ;
        RECT 31.630 170.425 31.920 170.470 ;
        RECT 33.490 170.425 33.780 170.470 ;
        RECT 40.955 170.610 41.245 170.655 ;
        RECT 44.060 170.610 44.845 170.655 ;
        RECT 40.955 170.470 44.845 170.610 ;
        RECT 40.955 170.425 41.545 170.470 ;
        RECT 29.310 170.270 29.600 170.315 ;
        RECT 31.630 170.270 31.845 170.425 ;
        RECT 29.310 170.130 31.845 170.270 ;
        RECT 32.100 170.270 32.420 170.330 ;
        RECT 32.575 170.270 32.865 170.315 ;
        RECT 32.100 170.130 32.865 170.270 ;
        RECT 29.310 170.085 29.600 170.130 ;
        RECT 32.100 170.070 32.420 170.130 ;
        RECT 32.575 170.085 32.865 170.130 ;
        RECT 35.795 170.270 36.085 170.315 ;
        RECT 36.240 170.270 36.560 170.330 ;
        RECT 35.795 170.130 36.560 170.270 ;
        RECT 35.795 170.085 36.085 170.130 ;
        RECT 36.240 170.070 36.560 170.130 ;
        RECT 36.700 170.070 37.020 170.330 ;
        RECT 37.160 170.070 37.480 170.330 ;
        RECT 37.620 170.270 37.940 170.330 ;
        RECT 40.380 170.270 40.700 170.330 ;
        RECT 37.620 170.130 40.700 170.270 ;
        RECT 37.620 170.070 37.940 170.130 ;
        RECT 40.380 170.070 40.700 170.130 ;
        RECT 41.255 170.110 41.545 170.425 ;
        RECT 44.060 170.425 44.845 170.470 ;
        RECT 46.835 170.610 47.125 170.655 ;
        RECT 47.280 170.610 47.600 170.670 ;
        RECT 46.835 170.470 47.600 170.610 ;
        RECT 46.835 170.425 47.125 170.470 ;
        RECT 44.060 170.410 44.380 170.425 ;
        RECT 47.280 170.410 47.600 170.470 ;
        RECT 50.615 170.610 50.905 170.655 ;
        RECT 53.855 170.610 54.505 170.655 ;
        RECT 50.615 170.470 54.505 170.610 ;
        RECT 50.615 170.425 51.205 170.470 ;
        RECT 53.855 170.425 54.505 170.470 ;
        RECT 56.940 170.610 57.260 170.670 ;
        RECT 56.940 170.470 58.090 170.610 ;
        RECT 50.915 170.330 51.205 170.425 ;
        RECT 56.940 170.410 57.260 170.470 ;
        RECT 42.335 170.270 42.625 170.315 ;
        RECT 45.915 170.270 46.205 170.315 ;
        RECT 47.750 170.270 48.040 170.315 ;
        RECT 42.335 170.130 48.040 170.270 ;
        RECT 42.335 170.085 42.625 170.130 ;
        RECT 45.915 170.085 46.205 170.130 ;
        RECT 47.750 170.085 48.040 170.130 ;
        RECT 50.915 170.110 51.280 170.330 ;
        RECT 57.950 170.315 58.090 170.470 ;
        RECT 59.330 170.315 59.470 170.810 ;
        RECT 62.550 170.810 70.140 170.950 ;
        RECT 62.550 170.655 62.690 170.810 ;
        RECT 69.820 170.750 70.140 170.810 ;
        RECT 73.975 170.950 74.265 170.995 ;
        RECT 74.420 170.950 74.740 171.010 ;
        RECT 88.220 170.950 88.540 171.010 ;
        RECT 73.975 170.810 74.740 170.950 ;
        RECT 73.975 170.765 74.265 170.810 ;
        RECT 74.420 170.750 74.740 170.810 ;
        RECT 74.970 170.810 87.990 170.950 ;
        RECT 62.475 170.425 62.765 170.655 ;
        RECT 74.970 170.610 75.110 170.810 ;
        RECT 69.450 170.470 75.110 170.610 ;
        RECT 77.130 170.610 77.420 170.655 ;
        RECT 79.480 170.610 79.800 170.670 ;
        RECT 80.390 170.610 80.680 170.655 ;
        RECT 77.130 170.470 80.680 170.610 ;
        RECT 50.960 170.070 51.280 170.110 ;
        RECT 51.995 170.270 52.285 170.315 ;
        RECT 55.575 170.270 55.865 170.315 ;
        RECT 57.410 170.270 57.700 170.315 ;
        RECT 51.995 170.130 57.700 170.270 ;
        RECT 51.995 170.085 52.285 170.130 ;
        RECT 55.575 170.085 55.865 170.130 ;
        RECT 57.410 170.085 57.700 170.130 ;
        RECT 57.875 170.085 58.165 170.315 ;
        RECT 59.255 170.085 59.545 170.315 ;
        RECT 60.160 170.270 60.480 170.330 ;
        RECT 64.315 170.270 64.605 170.315 ;
        RECT 60.160 170.130 64.605 170.270 ;
        RECT 29.800 169.930 30.120 169.990 ;
        RECT 33.020 169.930 33.340 169.990 ;
        RECT 29.800 169.790 33.340 169.930 ;
        RECT 29.800 169.730 30.120 169.790 ;
        RECT 33.020 169.730 33.340 169.790 ;
        RECT 34.415 169.930 34.705 169.975 ;
        RECT 35.320 169.930 35.640 169.990 ;
        RECT 48.215 169.930 48.505 169.975 ;
        RECT 34.415 169.790 48.505 169.930 ;
        RECT 34.415 169.745 34.705 169.790 ;
        RECT 35.320 169.730 35.640 169.790 ;
        RECT 48.215 169.745 48.505 169.790 ;
        RECT 50.500 169.930 50.820 169.990 ;
        RECT 56.495 169.930 56.785 169.975 ;
        RECT 50.500 169.790 56.785 169.930 ;
        RECT 50.500 169.730 50.820 169.790 ;
        RECT 56.495 169.745 56.785 169.790 ;
        RECT 29.310 169.590 29.600 169.635 ;
        RECT 32.090 169.590 32.380 169.635 ;
        RECT 33.950 169.590 34.240 169.635 ;
        RECT 39.920 169.590 40.240 169.650 ;
        RECT 42.335 169.590 42.625 169.635 ;
        RECT 45.455 169.590 45.745 169.635 ;
        RECT 47.345 169.590 47.635 169.635 ;
        RECT 29.310 169.450 34.240 169.590 ;
        RECT 29.310 169.405 29.600 169.450 ;
        RECT 32.090 169.405 32.380 169.450 ;
        RECT 33.950 169.405 34.240 169.450 ;
        RECT 34.490 169.450 41.990 169.590 ;
        RECT 25.445 169.250 25.735 169.295 ;
        RECT 32.560 169.250 32.880 169.310 ;
        RECT 25.445 169.110 32.880 169.250 ;
        RECT 25.445 169.065 25.735 169.110 ;
        RECT 32.560 169.050 32.880 169.110 ;
        RECT 33.020 169.250 33.340 169.310 ;
        RECT 34.490 169.250 34.630 169.450 ;
        RECT 39.920 169.390 40.240 169.450 ;
        RECT 33.020 169.110 34.630 169.250 ;
        RECT 33.020 169.050 33.340 169.110 ;
        RECT 39.000 169.050 39.320 169.310 ;
        RECT 39.475 169.250 39.765 169.295 ;
        RECT 41.300 169.250 41.620 169.310 ;
        RECT 39.475 169.110 41.620 169.250 ;
        RECT 41.850 169.250 41.990 169.450 ;
        RECT 42.335 169.450 47.635 169.590 ;
        RECT 42.335 169.405 42.625 169.450 ;
        RECT 45.455 169.405 45.745 169.450 ;
        RECT 47.345 169.405 47.635 169.450 ;
        RECT 51.995 169.590 52.285 169.635 ;
        RECT 55.115 169.590 55.405 169.635 ;
        RECT 57.005 169.590 57.295 169.635 ;
        RECT 51.995 169.450 57.295 169.590 ;
        RECT 57.950 169.590 58.090 170.085 ;
        RECT 60.160 170.070 60.480 170.130 ;
        RECT 64.315 170.085 64.605 170.130 ;
        RECT 65.680 170.270 66.000 170.330 ;
        RECT 69.450 170.315 69.590 170.470 ;
        RECT 77.130 170.425 77.420 170.470 ;
        RECT 79.480 170.410 79.800 170.470 ;
        RECT 80.390 170.425 80.680 170.470 ;
        RECT 81.310 170.610 81.600 170.655 ;
        RECT 83.170 170.610 83.460 170.655 ;
        RECT 81.310 170.470 83.460 170.610 ;
        RECT 81.310 170.425 81.600 170.470 ;
        RECT 83.170 170.425 83.460 170.470 ;
        RECT 69.375 170.270 69.665 170.315 ;
        RECT 65.680 170.130 69.665 170.270 ;
        RECT 65.680 170.070 66.000 170.130 ;
        RECT 69.375 170.085 69.665 170.130 ;
        RECT 72.135 170.270 72.425 170.315 ;
        RECT 73.500 170.270 73.820 170.330 ;
        RECT 72.135 170.130 73.820 170.270 ;
        RECT 72.135 170.085 72.425 170.130 ;
        RECT 73.500 170.070 73.820 170.130 ;
        RECT 78.990 170.270 79.280 170.315 ;
        RECT 81.310 170.270 81.525 170.425 ;
        RECT 78.990 170.130 81.525 170.270 ;
        RECT 87.850 170.270 87.990 170.810 ;
        RECT 88.220 170.810 94.890 170.950 ;
        RECT 88.220 170.750 88.540 170.810 ;
        RECT 91.440 170.610 91.760 170.670 ;
        RECT 93.755 170.610 94.045 170.655 ;
        RECT 91.440 170.470 94.045 170.610 ;
        RECT 94.750 170.610 94.890 170.810 ;
        RECT 96.040 170.750 96.360 171.010 ;
        RECT 99.720 170.950 100.040 171.010 ;
        RECT 102.955 170.950 103.245 170.995 ;
        RECT 99.720 170.810 103.245 170.950 ;
        RECT 99.720 170.750 100.040 170.810 ;
        RECT 102.955 170.765 103.245 170.810 ;
        RECT 133.700 170.790 139.470 171.930 ;
        RECT 99.275 170.610 99.565 170.655 ;
        RECT 112.140 170.610 112.460 170.670 ;
        RECT 94.750 170.470 99.030 170.610 ;
        RECT 91.440 170.410 91.760 170.470 ;
        RECT 93.755 170.425 94.045 170.470 ;
        RECT 97.880 170.270 98.200 170.330 ;
        RECT 98.355 170.270 98.645 170.315 ;
        RECT 87.850 170.130 98.645 170.270 ;
        RECT 98.890 170.270 99.030 170.470 ;
        RECT 99.275 170.470 112.460 170.610 ;
        RECT 99.275 170.425 99.565 170.470 ;
        RECT 112.140 170.410 112.460 170.470 ;
        RECT 133.700 170.600 136.690 170.790 ;
        RECT 101.100 170.270 101.420 170.330 ;
        RECT 98.890 170.130 101.420 170.270 ;
        RECT 78.990 170.085 79.280 170.130 ;
        RECT 97.880 170.070 98.200 170.130 ;
        RECT 98.355 170.085 98.645 170.130 ;
        RECT 101.100 170.070 101.420 170.130 ;
        RECT 102.495 170.270 102.785 170.315 ;
        RECT 102.940 170.270 103.260 170.330 ;
        RECT 104.795 170.270 105.085 170.315 ;
        RECT 102.495 170.130 105.085 170.270 ;
        RECT 102.495 170.085 102.785 170.130 ;
        RECT 102.940 170.070 103.260 170.130 ;
        RECT 104.795 170.085 105.085 170.130 ;
        RECT 111.220 170.070 111.540 170.330 ;
        RECT 133.700 170.120 134.930 170.600 ;
        RECT 59.700 169.930 60.020 169.990 ;
        RECT 64.760 169.930 65.080 169.990 ;
        RECT 59.700 169.790 65.080 169.930 ;
        RECT 59.700 169.730 60.020 169.790 ;
        RECT 64.760 169.730 65.080 169.790 ;
        RECT 66.600 169.930 66.920 169.990 ;
        RECT 67.995 169.930 68.285 169.975 ;
        RECT 66.600 169.790 68.285 169.930 ;
        RECT 66.600 169.730 66.920 169.790 ;
        RECT 67.995 169.745 68.285 169.790 ;
        RECT 70.740 169.730 71.060 169.990 ;
        RECT 71.660 169.730 71.980 169.990 ;
        RECT 75.800 169.930 76.120 169.990 ;
        RECT 82.255 169.930 82.545 169.975 ;
        RECT 75.800 169.790 82.545 169.930 ;
        RECT 75.800 169.730 76.120 169.790 ;
        RECT 82.255 169.745 82.545 169.790 ;
        RECT 84.095 169.930 84.385 169.975 ;
        RECT 85.460 169.930 85.780 169.990 ;
        RECT 84.095 169.790 85.780 169.930 ;
        RECT 84.095 169.745 84.385 169.790 ;
        RECT 85.460 169.730 85.780 169.790 ;
        RECT 94.660 169.930 94.980 169.990 ;
        RECT 95.135 169.930 95.425 169.975 ;
        RECT 94.660 169.790 95.425 169.930 ;
        RECT 94.660 169.730 94.980 169.790 ;
        RECT 95.135 169.745 95.425 169.790 ;
        RECT 61.080 169.590 61.400 169.650 ;
        RECT 57.950 169.450 61.400 169.590 ;
        RECT 51.995 169.405 52.285 169.450 ;
        RECT 55.115 169.405 55.405 169.450 ;
        RECT 57.005 169.405 57.295 169.450 ;
        RECT 61.080 169.390 61.400 169.450 ;
        RECT 63.380 169.590 63.700 169.650 ;
        RECT 78.990 169.590 79.280 169.635 ;
        RECT 81.770 169.590 82.060 169.635 ;
        RECT 83.630 169.590 83.920 169.635 ;
        RECT 95.210 169.590 95.350 169.745 ;
        RECT 95.580 169.730 95.900 169.990 ;
        RECT 102.020 169.930 102.340 169.990 ;
        RECT 103.415 169.930 103.705 169.975 ;
        RECT 96.130 169.790 103.705 169.930 ;
        RECT 96.130 169.590 96.270 169.790 ;
        RECT 102.020 169.730 102.340 169.790 ;
        RECT 103.415 169.745 103.705 169.790 ;
        RECT 105.240 169.930 105.560 169.990 ;
        RECT 107.555 169.930 107.845 169.975 ;
        RECT 110.760 169.930 111.080 169.990 ;
        RECT 105.240 169.790 111.080 169.930 ;
        RECT 105.240 169.730 105.560 169.790 ;
        RECT 107.555 169.745 107.845 169.790 ;
        RECT 110.760 169.730 111.080 169.790 ;
        RECT 63.380 169.450 78.790 169.590 ;
        RECT 63.380 169.390 63.700 169.450 ;
        RECT 43.600 169.250 43.920 169.310 ;
        RECT 41.850 169.110 43.920 169.250 ;
        RECT 39.475 169.065 39.765 169.110 ;
        RECT 41.300 169.050 41.620 169.110 ;
        RECT 43.600 169.050 43.920 169.110 ;
        RECT 44.060 169.250 44.380 169.310 ;
        RECT 49.135 169.250 49.425 169.295 ;
        RECT 53.720 169.250 54.040 169.310 ;
        RECT 44.060 169.110 54.040 169.250 ;
        RECT 44.060 169.050 44.380 169.110 ;
        RECT 49.135 169.065 49.425 169.110 ;
        RECT 53.720 169.050 54.040 169.110 ;
        RECT 59.700 169.250 60.020 169.310 ;
        RECT 60.175 169.250 60.465 169.295 ;
        RECT 59.700 169.110 60.465 169.250 ;
        RECT 59.700 169.050 60.020 169.110 ;
        RECT 60.175 169.065 60.465 169.110 ;
        RECT 62.000 169.050 62.320 169.310 ;
        RECT 73.500 169.250 73.820 169.310 ;
        RECT 75.125 169.250 75.415 169.295 ;
        RECT 73.500 169.110 75.415 169.250 ;
        RECT 78.650 169.250 78.790 169.450 ;
        RECT 78.990 169.450 83.920 169.590 ;
        RECT 78.990 169.405 79.280 169.450 ;
        RECT 81.770 169.405 82.060 169.450 ;
        RECT 83.630 169.405 83.920 169.450 ;
        RECT 84.630 169.450 96.270 169.590 ;
        RECT 83.160 169.250 83.480 169.310 ;
        RECT 78.650 169.110 83.480 169.250 ;
        RECT 73.500 169.050 73.820 169.110 ;
        RECT 75.125 169.065 75.415 169.110 ;
        RECT 83.160 169.050 83.480 169.110 ;
        RECT 84.080 169.250 84.400 169.310 ;
        RECT 84.630 169.250 84.770 169.450 ;
        RECT 84.080 169.110 84.770 169.250 ;
        RECT 85.460 169.250 85.780 169.310 ;
        RECT 87.315 169.250 87.605 169.295 ;
        RECT 89.600 169.250 89.920 169.310 ;
        RECT 85.460 169.110 89.920 169.250 ;
        RECT 84.080 169.050 84.400 169.110 ;
        RECT 85.460 169.050 85.780 169.110 ;
        RECT 87.315 169.065 87.605 169.110 ;
        RECT 89.600 169.050 89.920 169.110 ;
        RECT 97.420 169.250 97.740 169.310 ;
        RECT 97.895 169.250 98.185 169.295 ;
        RECT 97.420 169.110 98.185 169.250 ;
        RECT 97.420 169.050 97.740 169.110 ;
        RECT 97.895 169.065 98.185 169.110 ;
        RECT 98.800 169.250 99.120 169.310 ;
        RECT 100.655 169.250 100.945 169.295 ;
        RECT 98.800 169.110 100.945 169.250 ;
        RECT 98.800 169.050 99.120 169.110 ;
        RECT 100.655 169.065 100.945 169.110 ;
        RECT 101.100 169.250 101.420 169.310 ;
        RECT 110.300 169.250 110.620 169.310 ;
        RECT 101.100 169.110 110.620 169.250 ;
        RECT 101.100 169.050 101.420 169.110 ;
        RECT 110.300 169.050 110.620 169.110 ;
        RECT 22.830 168.430 113.450 168.910 ;
        RECT 24.295 168.230 24.585 168.275 ;
        RECT 25.660 168.230 25.980 168.290 ;
        RECT 24.295 168.090 25.980 168.230 ;
        RECT 24.295 168.045 24.585 168.090 ;
        RECT 25.660 168.030 25.980 168.090 ;
        RECT 31.640 168.230 31.960 168.290 ;
        RECT 37.620 168.230 37.940 168.290 ;
        RECT 31.640 168.090 37.940 168.230 ;
        RECT 31.640 168.030 31.960 168.090 ;
        RECT 37.620 168.030 37.940 168.090 ;
        RECT 38.540 168.230 38.860 168.290 ;
        RECT 49.135 168.230 49.425 168.275 ;
        RECT 49.580 168.230 49.900 168.290 ;
        RECT 38.540 168.090 45.670 168.230 ;
        RECT 38.540 168.030 38.860 168.090 ;
        RECT 39.935 167.890 40.225 167.935 ;
        RECT 42.680 167.890 43.000 167.950 ;
        RECT 39.935 167.750 43.000 167.890 ;
        RECT 39.935 167.705 40.225 167.750 ;
        RECT 42.680 167.690 43.000 167.750 ;
        RECT 27.515 167.550 27.805 167.595 ;
        RECT 29.340 167.550 29.660 167.610 ;
        RECT 36.715 167.550 37.005 167.595 ;
        RECT 27.515 167.410 37.005 167.550 ;
        RECT 27.515 167.365 27.805 167.410 ;
        RECT 29.340 167.350 29.660 167.410 ;
        RECT 36.715 167.365 37.005 167.410 ;
        RECT 41.300 167.550 41.620 167.610 ;
        RECT 42.235 167.550 42.525 167.595 ;
        RECT 45.530 167.550 45.670 168.090 ;
        RECT 49.135 168.090 49.900 168.230 ;
        RECT 49.135 168.045 49.425 168.090 ;
        RECT 49.580 168.030 49.900 168.090 ;
        RECT 50.500 168.030 50.820 168.290 ;
        RECT 63.380 168.230 63.700 168.290 ;
        RECT 51.050 168.090 63.700 168.230 ;
        RECT 46.360 167.890 46.680 167.950 ;
        RECT 51.050 167.890 51.190 168.090 ;
        RECT 63.380 168.030 63.700 168.090 ;
        RECT 67.980 168.030 68.300 168.290 ;
        RECT 70.740 168.230 71.060 168.290 ;
        RECT 71.215 168.230 71.505 168.275 ;
        RECT 88.005 168.230 88.295 168.275 ;
        RECT 92.360 168.230 92.680 168.290 ;
        RECT 95.580 168.230 95.900 168.290 ;
        RECT 70.740 168.090 71.505 168.230 ;
        RECT 70.740 168.030 71.060 168.090 ;
        RECT 71.215 168.045 71.505 168.090 ;
        RECT 85.090 168.090 95.900 168.230 ;
        RECT 46.360 167.750 51.190 167.890 ;
        RECT 55.215 167.890 55.505 167.935 ;
        RECT 58.335 167.890 58.625 167.935 ;
        RECT 60.225 167.890 60.515 167.935 ;
        RECT 70.280 167.890 70.600 167.950 ;
        RECT 55.215 167.750 60.515 167.890 ;
        RECT 46.360 167.690 46.680 167.750 ;
        RECT 55.215 167.705 55.505 167.750 ;
        RECT 58.335 167.705 58.625 167.750 ;
        RECT 60.225 167.705 60.515 167.750 ;
        RECT 64.390 167.750 70.600 167.890 ;
        RECT 45.915 167.550 46.205 167.595 ;
        RECT 50.040 167.550 50.360 167.610 ;
        RECT 41.300 167.410 42.910 167.550 ;
        RECT 45.530 167.410 50.360 167.550 ;
        RECT 26.120 167.210 26.440 167.270 ;
        RECT 28.880 167.210 29.200 167.270 ;
        RECT 29.815 167.210 30.105 167.255 ;
        RECT 26.120 167.070 30.105 167.210 ;
        RECT 26.120 167.010 26.440 167.070 ;
        RECT 28.880 167.010 29.200 167.070 ;
        RECT 29.815 167.025 30.105 167.070 ;
        RECT 34.875 167.210 35.165 167.255 ;
        RECT 35.320 167.210 35.640 167.270 ;
        RECT 34.875 167.070 35.640 167.210 ;
        RECT 36.790 167.210 36.930 167.365 ;
        RECT 41.300 167.350 41.620 167.410 ;
        RECT 42.235 167.365 42.525 167.410 ;
        RECT 42.770 167.270 42.910 167.410 ;
        RECT 45.915 167.365 46.205 167.410 ;
        RECT 50.040 167.350 50.360 167.410 ;
        RECT 59.700 167.350 60.020 167.610 ;
        RECT 61.080 167.350 61.400 167.610 ;
        RECT 38.540 167.210 38.860 167.270 ;
        RECT 36.790 167.070 38.860 167.210 ;
        RECT 34.875 167.025 35.165 167.070 ;
        RECT 35.320 167.010 35.640 167.070 ;
        RECT 38.540 167.010 38.860 167.070 ;
        RECT 39.920 167.210 40.240 167.270 ;
        RECT 40.395 167.210 40.685 167.255 ;
        RECT 39.920 167.070 40.685 167.210 ;
        RECT 39.920 167.010 40.240 167.070 ;
        RECT 40.395 167.025 40.685 167.070 ;
        RECT 42.680 167.010 43.000 167.270 ;
        RECT 47.295 167.210 47.585 167.255 ;
        RECT 43.230 167.070 47.585 167.210 ;
        RECT 26.595 166.870 26.885 166.915 ;
        RECT 32.560 166.870 32.880 166.930 ;
        RECT 38.095 166.870 38.385 166.915 ;
        RECT 26.595 166.730 38.385 166.870 ;
        RECT 26.595 166.685 26.885 166.730 ;
        RECT 32.560 166.670 32.880 166.730 ;
        RECT 38.095 166.685 38.385 166.730 ;
        RECT 40.855 166.870 41.145 166.915 ;
        RECT 41.300 166.870 41.620 166.930 ;
        RECT 43.230 166.870 43.370 167.070 ;
        RECT 47.295 167.025 47.585 167.070 ;
        RECT 47.740 167.210 48.060 167.270 ;
        RECT 49.595 167.210 49.885 167.255 ;
        RECT 47.740 167.070 49.885 167.210 ;
        RECT 47.740 167.010 48.060 167.070 ;
        RECT 49.595 167.025 49.885 167.070 ;
        RECT 50.975 167.210 51.265 167.255 ;
        RECT 51.880 167.210 52.200 167.270 ;
        RECT 64.390 167.255 64.530 167.750 ;
        RECT 70.280 167.690 70.600 167.750 ;
        RECT 66.155 167.550 66.445 167.595 ;
        RECT 64.850 167.410 66.445 167.550 ;
        RECT 71.290 167.550 71.430 168.045 ;
        RECT 82.715 167.890 83.005 167.935 ;
        RECT 82.715 167.750 84.770 167.890 ;
        RECT 82.715 167.705 83.005 167.750 ;
        RECT 84.630 167.610 84.770 167.750 ;
        RECT 77.195 167.550 77.485 167.595 ;
        RECT 78.560 167.550 78.880 167.610 ;
        RECT 79.955 167.550 80.245 167.595 ;
        RECT 84.080 167.550 84.400 167.610 ;
        RECT 71.290 167.410 84.400 167.550 ;
        RECT 50.975 167.070 52.200 167.210 ;
        RECT 50.975 167.025 51.265 167.070 ;
        RECT 51.880 167.010 52.200 167.070 ;
        RECT 40.855 166.730 41.620 166.870 ;
        RECT 40.855 166.685 41.145 166.730 ;
        RECT 41.300 166.670 41.620 166.730 ;
        RECT 41.850 166.730 43.370 166.870 ;
        RECT 44.995 166.870 45.285 166.915 ;
        RECT 46.820 166.870 47.140 166.930 ;
        RECT 54.135 166.915 54.425 167.230 ;
        RECT 55.215 167.210 55.505 167.255 ;
        RECT 58.795 167.210 59.085 167.255 ;
        RECT 60.630 167.210 60.920 167.255 ;
        RECT 55.215 167.070 60.920 167.210 ;
        RECT 55.215 167.025 55.505 167.070 ;
        RECT 58.795 167.025 59.085 167.070 ;
        RECT 60.630 167.025 60.920 167.070 ;
        RECT 64.315 167.025 64.605 167.255 ;
        RECT 44.995 166.730 47.140 166.870 ;
        RECT 27.500 166.530 27.820 166.590 ;
        RECT 30.275 166.530 30.565 166.575 ;
        RECT 27.500 166.390 30.565 166.530 ;
        RECT 27.500 166.330 27.820 166.390 ;
        RECT 30.275 166.345 30.565 166.390 ;
        RECT 32.115 166.530 32.405 166.575 ;
        RECT 34.860 166.530 35.180 166.590 ;
        RECT 32.115 166.390 35.180 166.530 ;
        RECT 32.115 166.345 32.405 166.390 ;
        RECT 34.860 166.330 35.180 166.390 ;
        RECT 37.620 166.530 37.940 166.590 ;
        RECT 41.850 166.530 41.990 166.730 ;
        RECT 44.995 166.685 45.285 166.730 ;
        RECT 46.820 166.670 47.140 166.730 ;
        RECT 51.435 166.870 51.725 166.915 ;
        RECT 53.835 166.870 54.425 166.915 ;
        RECT 57.075 166.870 57.725 166.915 ;
        RECT 51.435 166.730 57.725 166.870 ;
        RECT 51.435 166.685 51.725 166.730 ;
        RECT 53.835 166.685 54.125 166.730 ;
        RECT 57.075 166.685 57.725 166.730 ;
        RECT 59.700 166.870 60.020 166.930 ;
        RECT 64.850 166.870 64.990 167.410 ;
        RECT 66.155 167.365 66.445 167.410 ;
        RECT 77.195 167.365 77.485 167.410 ;
        RECT 78.560 167.350 78.880 167.410 ;
        RECT 79.955 167.365 80.245 167.410 ;
        RECT 84.080 167.350 84.400 167.410 ;
        RECT 84.540 167.350 84.860 167.610 ;
        RECT 65.680 167.210 66.000 167.270 ;
        RECT 67.075 167.210 67.365 167.255 ;
        RECT 65.680 167.070 67.365 167.210 ;
        RECT 65.680 167.010 66.000 167.070 ;
        RECT 67.075 167.025 67.365 167.070 ;
        RECT 68.440 167.210 68.760 167.270 ;
        RECT 68.915 167.210 69.205 167.255 ;
        RECT 68.440 167.070 69.205 167.210 ;
        RECT 68.440 167.010 68.760 167.070 ;
        RECT 68.915 167.025 69.205 167.070 ;
        RECT 69.820 167.010 70.140 167.270 ;
        RECT 70.280 167.210 70.600 167.270 ;
        RECT 72.135 167.210 72.425 167.255 ;
        RECT 70.280 167.070 72.425 167.210 ;
        RECT 70.280 167.010 70.600 167.070 ;
        RECT 72.135 167.025 72.425 167.070 ;
        RECT 73.500 167.210 73.820 167.270 ;
        RECT 85.090 167.255 85.230 168.090 ;
        RECT 88.005 168.045 88.295 168.090 ;
        RECT 92.360 168.030 92.680 168.090 ;
        RECT 95.580 168.030 95.900 168.090 ;
        RECT 100.180 168.230 100.500 168.290 ;
        RECT 105.715 168.230 106.005 168.275 ;
        RECT 100.180 168.090 106.005 168.230 ;
        RECT 100.180 168.030 100.500 168.090 ;
        RECT 105.715 168.045 106.005 168.090 ;
        RECT 91.870 167.890 92.160 167.935 ;
        RECT 94.650 167.890 94.940 167.935 ;
        RECT 96.510 167.890 96.800 167.935 ;
        RECT 91.870 167.750 96.800 167.890 ;
        RECT 91.870 167.705 92.160 167.750 ;
        RECT 94.650 167.705 94.940 167.750 ;
        RECT 96.510 167.705 96.800 167.750 ;
        RECT 105.255 167.890 105.545 167.935 ;
        RECT 105.255 167.750 108.690 167.890 ;
        RECT 105.255 167.705 105.545 167.750 ;
        RECT 89.600 167.550 89.920 167.610 ;
        RECT 89.600 167.410 94.890 167.550 ;
        RECT 89.600 167.350 89.920 167.410 ;
        RECT 76.735 167.210 77.025 167.255 ;
        RECT 80.875 167.210 81.165 167.255 ;
        RECT 73.500 167.070 77.025 167.210 ;
        RECT 73.500 167.010 73.820 167.070 ;
        RECT 76.735 167.025 77.025 167.070 ;
        RECT 77.270 167.070 81.165 167.210 ;
        RECT 59.700 166.730 64.990 166.870 ;
        RECT 71.660 166.870 71.980 166.930 ;
        RECT 77.270 166.870 77.410 167.070 ;
        RECT 80.875 167.025 81.165 167.070 ;
        RECT 85.015 167.025 85.305 167.255 ;
        RECT 90.980 167.210 91.300 167.270 ;
        RECT 89.690 167.070 91.300 167.210 ;
        RECT 71.660 166.730 77.410 166.870 ;
        RECT 79.480 166.870 79.800 166.930 ;
        RECT 84.555 166.870 84.845 166.915 ;
        RECT 89.690 166.870 89.830 167.070 ;
        RECT 90.980 167.010 91.300 167.070 ;
        RECT 91.870 167.210 92.160 167.255 ;
        RECT 94.750 167.210 94.890 167.410 ;
        RECT 95.120 167.350 95.440 167.610 ;
        RECT 96.975 167.550 97.265 167.595 ;
        RECT 97.880 167.550 98.200 167.610 ;
        RECT 96.975 167.410 98.200 167.550 ;
        RECT 96.975 167.365 97.265 167.410 ;
        RECT 97.050 167.210 97.190 167.365 ;
        RECT 97.880 167.350 98.200 167.410 ;
        RECT 102.020 167.350 102.340 167.610 ;
        RECT 102.940 167.350 103.260 167.610 ;
        RECT 108.550 167.595 108.690 167.750 ;
        RECT 108.475 167.365 108.765 167.595 ;
        RECT 91.870 167.070 94.405 167.210 ;
        RECT 94.750 167.070 97.190 167.210 ;
        RECT 98.355 167.210 98.645 167.255 ;
        RECT 99.260 167.210 99.580 167.270 ;
        RECT 98.355 167.070 99.580 167.210 ;
        RECT 91.870 167.025 92.160 167.070 ;
        RECT 90.060 166.915 90.380 166.930 ;
        RECT 94.190 166.915 94.405 167.070 ;
        RECT 98.355 167.025 98.645 167.070 ;
        RECT 99.260 167.010 99.580 167.070 ;
        RECT 111.680 167.010 112.000 167.270 ;
        RECT 79.480 166.730 84.845 166.870 ;
        RECT 59.700 166.670 60.020 166.730 ;
        RECT 71.660 166.670 71.980 166.730 ;
        RECT 79.480 166.670 79.800 166.730 ;
        RECT 84.555 166.685 84.845 166.730 ;
        RECT 85.090 166.730 89.830 166.870 ;
        RECT 90.010 166.870 90.380 166.915 ;
        RECT 93.270 166.870 93.560 166.915 ;
        RECT 90.010 166.730 93.560 166.870 ;
        RECT 37.620 166.390 41.990 166.530 ;
        RECT 43.600 166.530 43.920 166.590 ;
        RECT 52.355 166.530 52.645 166.575 ;
        RECT 52.800 166.530 53.120 166.590 ;
        RECT 43.600 166.390 53.120 166.530 ;
        RECT 37.620 166.330 37.940 166.390 ;
        RECT 43.600 166.330 43.920 166.390 ;
        RECT 52.355 166.345 52.645 166.390 ;
        RECT 52.800 166.330 53.120 166.390 ;
        RECT 72.120 166.530 72.440 166.590 ;
        RECT 73.055 166.530 73.345 166.575 ;
        RECT 72.120 166.390 73.345 166.530 ;
        RECT 72.120 166.330 72.440 166.390 ;
        RECT 73.055 166.345 73.345 166.390 ;
        RECT 74.435 166.530 74.725 166.575 ;
        RECT 74.880 166.530 75.200 166.590 ;
        RECT 74.435 166.390 75.200 166.530 ;
        RECT 74.435 166.345 74.725 166.390 ;
        RECT 74.880 166.330 75.200 166.390 ;
        RECT 76.275 166.530 76.565 166.575 ;
        RECT 76.720 166.530 77.040 166.590 ;
        RECT 76.275 166.390 77.040 166.530 ;
        RECT 76.275 166.345 76.565 166.390 ;
        RECT 76.720 166.330 77.040 166.390 ;
        RECT 80.415 166.530 80.705 166.575 ;
        RECT 85.090 166.530 85.230 166.730 ;
        RECT 90.010 166.685 90.380 166.730 ;
        RECT 93.270 166.685 93.560 166.730 ;
        RECT 94.190 166.870 94.480 166.915 ;
        RECT 96.050 166.870 96.340 166.915 ;
        RECT 94.190 166.730 96.340 166.870 ;
        RECT 94.190 166.685 94.480 166.730 ;
        RECT 96.050 166.685 96.340 166.730 ;
        RECT 101.115 166.870 101.405 166.915 ;
        RECT 102.940 166.870 103.260 166.930 ;
        RECT 101.115 166.730 103.260 166.870 ;
        RECT 101.115 166.685 101.405 166.730 ;
        RECT 90.060 166.670 90.380 166.685 ;
        RECT 102.940 166.670 103.260 166.730 ;
        RECT 106.620 166.870 106.940 166.930 ;
        RECT 110.315 166.870 110.605 166.915 ;
        RECT 106.620 166.730 110.605 166.870 ;
        RECT 106.620 166.670 106.940 166.730 ;
        RECT 110.315 166.685 110.605 166.730 ;
        RECT 80.415 166.390 85.230 166.530 ;
        RECT 85.920 166.530 86.240 166.590 ;
        RECT 86.855 166.530 87.145 166.575 ;
        RECT 85.920 166.390 87.145 166.530 ;
        RECT 80.415 166.345 80.705 166.390 ;
        RECT 85.920 166.330 86.240 166.390 ;
        RECT 86.855 166.345 87.145 166.390 ;
        RECT 99.720 166.530 100.040 166.590 ;
        RECT 103.400 166.530 103.720 166.590 ;
        RECT 99.720 166.390 103.720 166.530 ;
        RECT 99.720 166.330 100.040 166.390 ;
        RECT 103.400 166.330 103.720 166.390 ;
        RECT 22.830 165.710 113.450 166.190 ;
        RECT 40.855 165.510 41.145 165.555 ;
        RECT 47.740 165.510 48.060 165.570 ;
        RECT 40.855 165.370 48.060 165.510 ;
        RECT 40.855 165.325 41.145 165.370 ;
        RECT 47.740 165.310 48.060 165.370 ;
        RECT 48.215 165.510 48.505 165.555 ;
        RECT 52.340 165.510 52.660 165.570 ;
        RECT 48.215 165.370 52.660 165.510 ;
        RECT 48.215 165.325 48.505 165.370 ;
        RECT 52.340 165.310 52.660 165.370 ;
        RECT 53.720 165.310 54.040 165.570 ;
        RECT 62.000 165.510 62.320 165.570 ;
        RECT 60.250 165.370 62.320 165.510 ;
        RECT 25.200 165.170 25.520 165.230 ;
        RECT 26.530 165.170 26.820 165.215 ;
        RECT 29.790 165.170 30.080 165.215 ;
        RECT 25.200 165.030 30.080 165.170 ;
        RECT 25.200 164.970 25.520 165.030 ;
        RECT 26.530 164.985 26.820 165.030 ;
        RECT 29.790 164.985 30.080 165.030 ;
        RECT 30.710 165.170 31.000 165.215 ;
        RECT 32.570 165.170 32.860 165.215 ;
        RECT 30.710 165.030 32.860 165.170 ;
        RECT 30.710 164.985 31.000 165.030 ;
        RECT 32.570 164.985 32.860 165.030 ;
        RECT 44.535 165.170 44.825 165.215 ;
        RECT 53.275 165.170 53.565 165.215 ;
        RECT 44.535 165.030 53.565 165.170 ;
        RECT 44.535 164.985 44.825 165.030 ;
        RECT 53.275 164.985 53.565 165.030 ;
        RECT 28.390 164.830 28.680 164.875 ;
        RECT 30.710 164.830 30.925 164.985 ;
        RECT 28.390 164.690 30.925 164.830 ;
        RECT 34.415 164.830 34.705 164.875 ;
        RECT 41.775 164.830 42.065 164.875 ;
        RECT 43.600 164.830 43.920 164.890 ;
        RECT 34.415 164.690 41.530 164.830 ;
        RECT 28.390 164.645 28.680 164.690 ;
        RECT 34.415 164.645 34.705 164.690 ;
        RECT 24.525 164.490 24.815 164.535 ;
        RECT 26.120 164.490 26.440 164.550 ;
        RECT 24.525 164.350 26.440 164.490 ;
        RECT 24.525 164.305 24.815 164.350 ;
        RECT 26.120 164.290 26.440 164.350 ;
        RECT 31.640 164.290 31.960 164.550 ;
        RECT 33.495 164.490 33.785 164.535 ;
        RECT 35.320 164.490 35.640 164.550 ;
        RECT 33.495 164.350 35.640 164.490 ;
        RECT 33.495 164.305 33.785 164.350 ;
        RECT 35.320 164.290 35.640 164.350 ;
        RECT 38.095 164.305 38.385 164.535 ;
        RECT 41.390 164.490 41.530 164.690 ;
        RECT 41.775 164.690 43.920 164.830 ;
        RECT 41.775 164.645 42.065 164.690 ;
        RECT 43.600 164.630 43.920 164.690 ;
        RECT 46.820 164.830 47.140 164.890 ;
        RECT 57.415 164.830 57.705 164.875 ;
        RECT 46.820 164.690 57.705 164.830 ;
        RECT 46.820 164.630 47.140 164.690 ;
        RECT 57.415 164.645 57.705 164.690 ;
        RECT 44.060 164.490 44.380 164.550 ;
        RECT 41.390 164.350 44.380 164.490 ;
        RECT 28.390 164.150 28.680 164.195 ;
        RECT 31.170 164.150 31.460 164.195 ;
        RECT 33.030 164.150 33.320 164.195 ;
        RECT 28.390 164.010 33.320 164.150 ;
        RECT 38.170 164.150 38.310 164.305 ;
        RECT 44.060 164.290 44.380 164.350 ;
        RECT 45.455 164.490 45.745 164.535 ;
        RECT 50.960 164.490 51.280 164.550 ;
        RECT 45.455 164.350 51.280 164.490 ;
        RECT 45.455 164.305 45.745 164.350 ;
        RECT 50.960 164.290 51.280 164.350 ;
        RECT 53.260 164.490 53.580 164.550 ;
        RECT 54.195 164.490 54.485 164.535 ;
        RECT 56.035 164.490 56.325 164.535 ;
        RECT 53.260 164.350 56.325 164.490 ;
        RECT 53.260 164.290 53.580 164.350 ;
        RECT 54.195 164.305 54.485 164.350 ;
        RECT 56.035 164.305 56.325 164.350 ;
        RECT 51.435 164.150 51.725 164.195 ;
        RECT 38.170 164.010 51.725 164.150 ;
        RECT 56.110 164.150 56.250 164.305 ;
        RECT 56.940 164.290 57.260 164.550 ;
        RECT 60.250 164.490 60.390 165.370 ;
        RECT 62.000 165.310 62.320 165.370 ;
        RECT 67.520 165.510 67.840 165.570 ;
        RECT 69.835 165.510 70.125 165.555 ;
        RECT 67.520 165.370 70.125 165.510 ;
        RECT 67.520 165.310 67.840 165.370 ;
        RECT 69.835 165.325 70.125 165.370 ;
        RECT 75.800 165.310 76.120 165.570 ;
        RECT 93.740 165.510 94.060 165.570 ;
        RECT 90.150 165.370 94.060 165.510 ;
        RECT 60.620 165.170 60.940 165.230 ;
        RECT 61.195 165.170 61.485 165.215 ;
        RECT 64.435 165.170 65.085 165.215 ;
        RECT 60.620 165.030 65.085 165.170 ;
        RECT 60.620 164.970 60.940 165.030 ;
        RECT 61.195 164.985 61.785 165.030 ;
        RECT 64.435 164.985 65.085 165.030 ;
        RECT 61.495 164.670 61.785 164.985 ;
        RECT 67.060 164.970 67.380 165.230 ;
        RECT 71.200 165.170 71.520 165.230 ;
        RECT 68.990 165.030 71.520 165.170 ;
        RECT 68.990 164.875 69.130 165.030 ;
        RECT 71.200 164.970 71.520 165.030 ;
        RECT 82.650 165.170 82.940 165.215 ;
        RECT 85.000 165.170 85.320 165.230 ;
        RECT 85.910 165.170 86.200 165.215 ;
        RECT 82.650 165.030 86.200 165.170 ;
        RECT 82.650 164.985 82.940 165.030 ;
        RECT 85.000 164.970 85.320 165.030 ;
        RECT 85.910 164.985 86.200 165.030 ;
        RECT 86.830 165.170 87.120 165.215 ;
        RECT 88.690 165.170 88.980 165.215 ;
        RECT 86.830 165.030 88.980 165.170 ;
        RECT 86.830 164.985 87.120 165.030 ;
        RECT 88.690 164.985 88.980 165.030 ;
        RECT 62.575 164.830 62.865 164.875 ;
        RECT 66.155 164.830 66.445 164.875 ;
        RECT 67.990 164.830 68.280 164.875 ;
        RECT 62.575 164.690 68.280 164.830 ;
        RECT 62.575 164.645 62.865 164.690 ;
        RECT 66.155 164.645 66.445 164.690 ;
        RECT 67.990 164.645 68.280 164.690 ;
        RECT 68.915 164.645 69.205 164.875 ;
        RECT 70.740 164.630 71.060 164.890 ;
        RECT 71.660 164.630 71.980 164.890 ;
        RECT 72.120 164.630 72.440 164.890 ;
        RECT 72.580 164.630 72.900 164.890 ;
        RECT 74.880 164.630 75.200 164.890 ;
        RECT 76.720 164.830 77.040 164.890 ;
        RECT 77.655 164.830 77.945 164.875 ;
        RECT 76.720 164.690 77.945 164.830 ;
        RECT 76.720 164.630 77.040 164.690 ;
        RECT 77.655 164.645 77.945 164.690 ;
        RECT 78.115 164.830 78.405 164.875 ;
        RECT 79.480 164.830 79.800 164.890 ;
        RECT 80.645 164.830 80.935 164.875 ;
        RECT 78.115 164.690 80.935 164.830 ;
        RECT 78.115 164.645 78.405 164.690 ;
        RECT 79.480 164.630 79.800 164.690 ;
        RECT 80.645 164.645 80.935 164.690 ;
        RECT 84.510 164.830 84.800 164.875 ;
        RECT 86.830 164.830 87.045 164.985 ;
        RECT 84.510 164.690 87.045 164.830 ;
        RECT 84.510 164.645 84.800 164.690 ;
        RECT 89.140 164.630 89.460 164.890 ;
        RECT 89.600 164.630 89.920 164.890 ;
        RECT 90.150 164.875 90.290 165.370 ;
        RECT 93.740 165.310 94.060 165.370 ;
        RECT 95.120 165.510 95.440 165.570 ;
        RECT 97.435 165.510 97.725 165.555 ;
        RECT 95.120 165.370 97.725 165.510 ;
        RECT 95.120 165.310 95.440 165.370 ;
        RECT 97.435 165.325 97.725 165.370 ;
        RECT 99.735 165.510 100.025 165.555 ;
        RECT 102.480 165.510 102.800 165.570 ;
        RECT 99.735 165.370 102.800 165.510 ;
        RECT 135.580 165.470 136.830 166.590 ;
        RECT 99.735 165.325 100.025 165.370 ;
        RECT 102.480 165.310 102.800 165.370 ;
        RECT 90.520 165.170 90.840 165.230 ;
        RECT 103.400 165.170 103.720 165.230 ;
        RECT 103.975 165.170 104.265 165.215 ;
        RECT 107.215 165.170 107.865 165.215 ;
        RECT 90.520 165.030 94.890 165.170 ;
        RECT 90.520 164.970 90.840 165.030 ;
        RECT 90.075 164.645 90.365 164.875 ;
        RECT 90.995 164.645 91.285 164.875 ;
        RECT 91.455 164.645 91.745 164.875 ;
        RECT 91.915 164.830 92.205 164.875 ;
        RECT 92.360 164.830 92.680 164.890 ;
        RECT 91.915 164.690 92.680 164.830 ;
        RECT 91.915 164.645 92.205 164.690 ;
        RECT 60.620 164.490 60.940 164.550 ;
        RECT 59.435 164.350 60.940 164.490 ;
        RECT 59.435 164.150 59.575 164.350 ;
        RECT 60.620 164.290 60.940 164.350 ;
        RECT 61.080 164.490 61.400 164.550 ;
        RECT 68.455 164.490 68.745 164.535 ;
        RECT 72.210 164.490 72.350 164.630 ;
        RECT 61.080 164.350 68.745 164.490 ;
        RECT 61.080 164.290 61.400 164.350 ;
        RECT 68.455 164.305 68.745 164.350 ;
        RECT 71.750 164.350 72.350 164.490 ;
        RECT 77.195 164.490 77.485 164.535 ;
        RECT 78.560 164.490 78.880 164.550 ;
        RECT 77.195 164.350 78.880 164.490 ;
        RECT 71.750 164.210 71.890 164.350 ;
        RECT 77.195 164.305 77.485 164.350 ;
        RECT 78.560 164.290 78.880 164.350 ;
        RECT 87.760 164.290 88.080 164.550 ;
        RECT 89.230 164.490 89.370 164.630 ;
        RECT 91.070 164.490 91.210 164.645 ;
        RECT 89.230 164.350 91.210 164.490 ;
        RECT 91.530 164.490 91.670 164.645 ;
        RECT 92.360 164.630 92.680 164.690 ;
        RECT 93.740 164.630 94.060 164.890 ;
        RECT 94.750 164.875 94.890 165.030 ;
        RECT 103.400 165.030 107.865 165.170 ;
        RECT 103.400 164.970 103.720 165.030 ;
        RECT 103.975 164.985 104.565 165.030 ;
        RECT 107.215 164.985 107.865 165.030 ;
        RECT 94.675 164.645 94.965 164.875 ;
        RECT 95.135 164.645 95.425 164.875 ;
        RECT 95.595 164.645 95.885 164.875 ;
        RECT 97.420 164.830 97.740 164.890 ;
        RECT 98.355 164.830 98.645 164.875 ;
        RECT 97.420 164.690 98.645 164.830 ;
        RECT 95.210 164.490 95.350 164.645 ;
        RECT 91.530 164.350 95.350 164.490 ;
        RECT 56.110 164.010 59.575 164.150 ;
        RECT 59.715 164.150 60.005 164.195 ;
        RECT 62.575 164.150 62.865 164.195 ;
        RECT 65.695 164.150 65.985 164.195 ;
        RECT 67.585 164.150 67.875 164.195 ;
        RECT 59.715 164.010 61.770 164.150 ;
        RECT 28.390 163.965 28.680 164.010 ;
        RECT 31.170 163.965 31.460 164.010 ;
        RECT 33.030 163.965 33.320 164.010 ;
        RECT 51.435 163.965 51.725 164.010 ;
        RECT 59.715 163.965 60.005 164.010 ;
        RECT 37.175 163.810 37.465 163.855 ;
        RECT 50.500 163.810 50.820 163.870 ;
        RECT 37.175 163.670 50.820 163.810 ;
        RECT 37.175 163.625 37.465 163.670 ;
        RECT 50.500 163.610 50.820 163.670 ;
        RECT 59.255 163.810 59.545 163.855 ;
        RECT 61.080 163.810 61.400 163.870 ;
        RECT 59.255 163.670 61.400 163.810 ;
        RECT 61.630 163.810 61.770 164.010 ;
        RECT 62.575 164.010 67.875 164.150 ;
        RECT 62.575 163.965 62.865 164.010 ;
        RECT 65.695 163.965 65.985 164.010 ;
        RECT 67.585 163.965 67.875 164.010 ;
        RECT 71.660 163.950 71.980 164.210 ;
        RECT 82.700 164.150 83.020 164.210 ;
        RECT 72.210 164.010 83.020 164.150 ;
        RECT 64.300 163.810 64.620 163.870 ;
        RECT 61.630 163.670 64.620 163.810 ;
        RECT 59.255 163.625 59.545 163.670 ;
        RECT 61.080 163.610 61.400 163.670 ;
        RECT 64.300 163.610 64.620 163.670 ;
        RECT 67.980 163.810 68.300 163.870 ;
        RECT 72.210 163.810 72.350 164.010 ;
        RECT 82.700 163.950 83.020 164.010 ;
        RECT 84.510 164.150 84.800 164.195 ;
        RECT 87.290 164.150 87.580 164.195 ;
        RECT 89.150 164.150 89.440 164.195 ;
        RECT 84.510 164.010 89.440 164.150 ;
        RECT 84.510 163.965 84.800 164.010 ;
        RECT 87.290 163.965 87.580 164.010 ;
        RECT 89.150 163.965 89.440 164.010 ;
        RECT 67.980 163.670 72.350 163.810 ;
        RECT 72.580 163.810 72.900 163.870 ;
        RECT 73.975 163.810 74.265 163.855 ;
        RECT 72.580 163.670 74.265 163.810 ;
        RECT 67.980 163.610 68.300 163.670 ;
        RECT 72.580 163.610 72.900 163.670 ;
        RECT 73.975 163.625 74.265 163.670 ;
        RECT 79.940 163.610 80.260 163.870 ;
        RECT 83.160 163.810 83.480 163.870 ;
        RECT 90.980 163.810 91.300 163.870 ;
        RECT 91.530 163.810 91.670 164.350 ;
        RECT 94.200 164.150 94.520 164.210 ;
        RECT 95.670 164.150 95.810 164.645 ;
        RECT 97.420 164.630 97.740 164.690 ;
        RECT 98.355 164.645 98.645 164.690 ;
        RECT 98.800 164.630 99.120 164.890 ;
        RECT 101.100 164.630 101.420 164.890 ;
        RECT 104.275 164.670 104.565 164.985 ;
        RECT 105.355 164.830 105.645 164.875 ;
        RECT 108.935 164.830 109.225 164.875 ;
        RECT 110.770 164.830 111.060 164.875 ;
        RECT 105.355 164.690 111.060 164.830 ;
        RECT 105.355 164.645 105.645 164.690 ;
        RECT 108.935 164.645 109.225 164.690 ;
        RECT 110.770 164.645 111.060 164.690 ;
        RECT 111.220 164.630 111.540 164.890 ;
        RECT 109.840 164.290 110.160 164.550 ;
        RECT 97.880 164.150 98.200 164.210 ;
        RECT 94.200 164.010 98.200 164.150 ;
        RECT 94.200 163.950 94.520 164.010 ;
        RECT 97.880 163.950 98.200 164.010 ;
        RECT 98.800 164.150 99.120 164.210 ;
        RECT 102.495 164.150 102.785 164.195 ;
        RECT 98.800 164.010 102.785 164.150 ;
        RECT 98.800 163.950 99.120 164.010 ;
        RECT 102.495 163.965 102.785 164.010 ;
        RECT 105.355 164.150 105.645 164.195 ;
        RECT 108.475 164.150 108.765 164.195 ;
        RECT 110.365 164.150 110.655 164.195 ;
        RECT 105.355 164.010 110.655 164.150 ;
        RECT 105.355 163.965 105.645 164.010 ;
        RECT 108.475 163.965 108.765 164.010 ;
        RECT 110.365 163.965 110.655 164.010 ;
        RECT 83.160 163.670 91.670 163.810 ;
        RECT 93.295 163.810 93.585 163.855 ;
        RECT 96.040 163.810 96.360 163.870 ;
        RECT 93.295 163.670 96.360 163.810 ;
        RECT 83.160 163.610 83.480 163.670 ;
        RECT 90.980 163.610 91.300 163.670 ;
        RECT 93.295 163.625 93.585 163.670 ;
        RECT 96.040 163.610 96.360 163.670 ;
        RECT 96.960 163.610 97.280 163.870 ;
        RECT 101.575 163.810 101.865 163.855 ;
        RECT 106.160 163.810 106.480 163.870 ;
        RECT 101.575 163.670 106.480 163.810 ;
        RECT 101.575 163.625 101.865 163.670 ;
        RECT 106.160 163.610 106.480 163.670 ;
        RECT 22.830 162.990 113.450 163.470 ;
        RECT 31.640 162.790 31.960 162.850 ;
        RECT 33.955 162.790 34.245 162.835 ;
        RECT 31.640 162.650 34.245 162.790 ;
        RECT 31.640 162.590 31.960 162.650 ;
        RECT 33.955 162.605 34.245 162.650 ;
        RECT 35.780 162.790 36.100 162.850 ;
        RECT 36.715 162.790 37.005 162.835 ;
        RECT 35.780 162.650 37.005 162.790 ;
        RECT 35.780 162.590 36.100 162.650 ;
        RECT 36.715 162.605 37.005 162.650 ;
        RECT 39.245 162.790 39.535 162.835 ;
        RECT 40.840 162.790 41.160 162.850 ;
        RECT 46.820 162.790 47.140 162.850 ;
        RECT 50.960 162.790 51.280 162.850 ;
        RECT 57.415 162.790 57.705 162.835 ;
        RECT 39.245 162.650 48.430 162.790 ;
        RECT 39.245 162.605 39.535 162.650 ;
        RECT 40.840 162.590 41.160 162.650 ;
        RECT 46.820 162.590 47.140 162.650 ;
        RECT 28.390 162.450 28.680 162.495 ;
        RECT 31.170 162.450 31.460 162.495 ;
        RECT 33.030 162.450 33.320 162.495 ;
        RECT 28.390 162.310 33.320 162.450 ;
        RECT 28.390 162.265 28.680 162.310 ;
        RECT 31.170 162.265 31.460 162.310 ;
        RECT 33.030 162.265 33.320 162.310 ;
        RECT 43.110 162.450 43.400 162.495 ;
        RECT 45.890 162.450 46.180 162.495 ;
        RECT 47.750 162.450 48.040 162.495 ;
        RECT 43.110 162.310 48.040 162.450 ;
        RECT 43.110 162.265 43.400 162.310 ;
        RECT 45.890 162.265 46.180 162.310 ;
        RECT 47.750 162.265 48.040 162.310 ;
        RECT 30.260 162.110 30.580 162.170 ;
        RECT 31.655 162.110 31.945 162.155 ;
        RECT 30.260 161.970 31.945 162.110 ;
        RECT 30.260 161.910 30.580 161.970 ;
        RECT 31.655 161.925 31.945 161.970 ;
        RECT 33.495 162.110 33.785 162.155 ;
        RECT 35.320 162.110 35.640 162.170 ;
        RECT 38.080 162.110 38.400 162.170 ;
        RECT 33.495 161.970 46.130 162.110 ;
        RECT 33.495 161.925 33.785 161.970 ;
        RECT 35.320 161.910 35.640 161.970 ;
        RECT 38.080 161.910 38.400 161.970 ;
        RECT 28.390 161.770 28.680 161.815 ;
        RECT 28.390 161.630 30.925 161.770 ;
        RECT 28.390 161.585 28.680 161.630 ;
        RECT 26.530 161.430 26.820 161.475 ;
        RECT 28.880 161.430 29.200 161.490 ;
        RECT 30.710 161.475 30.925 161.630 ;
        RECT 34.860 161.570 35.180 161.830 ;
        RECT 37.175 161.585 37.465 161.815 ;
        RECT 29.790 161.430 30.080 161.475 ;
        RECT 26.530 161.290 30.080 161.430 ;
        RECT 26.530 161.245 26.820 161.290 ;
        RECT 28.880 161.230 29.200 161.290 ;
        RECT 29.790 161.245 30.080 161.290 ;
        RECT 30.710 161.430 31.000 161.475 ;
        RECT 32.570 161.430 32.860 161.475 ;
        RECT 30.710 161.290 32.860 161.430 ;
        RECT 30.710 161.245 31.000 161.290 ;
        RECT 32.570 161.245 32.860 161.290 ;
        RECT 35.320 161.430 35.640 161.490 ;
        RECT 37.250 161.430 37.390 161.585 ;
        RECT 38.540 161.570 38.860 161.830 ;
        RECT 43.110 161.770 43.400 161.815 ;
        RECT 45.990 161.770 46.130 161.970 ;
        RECT 46.360 161.910 46.680 162.170 ;
        RECT 48.290 162.110 48.430 162.650 ;
        RECT 50.960 162.650 57.705 162.790 ;
        RECT 50.960 162.590 51.280 162.650 ;
        RECT 57.415 162.605 57.705 162.650 ;
        RECT 66.615 162.790 66.905 162.835 ;
        RECT 67.060 162.790 67.380 162.850 ;
        RECT 79.480 162.790 79.800 162.850 ;
        RECT 66.615 162.650 67.380 162.790 ;
        RECT 66.615 162.605 66.905 162.650 ;
        RECT 67.060 162.590 67.380 162.650 ;
        RECT 68.070 162.650 79.800 162.790 ;
        RECT 50.040 162.450 50.360 162.510 ;
        RECT 53.260 162.450 53.580 162.510 ;
        RECT 64.300 162.450 64.620 162.510 ;
        RECT 50.040 162.310 53.580 162.450 ;
        RECT 50.040 162.250 50.360 162.310 ;
        RECT 51.510 162.155 51.650 162.310 ;
        RECT 53.260 162.250 53.580 162.310 ;
        RECT 60.250 162.310 64.620 162.450 ;
        RECT 50.975 162.110 51.265 162.155 ;
        RECT 48.290 161.970 51.265 162.110 ;
        RECT 50.975 161.925 51.265 161.970 ;
        RECT 51.435 161.925 51.725 162.155 ;
        RECT 54.195 162.110 54.485 162.155 ;
        RECT 60.250 162.110 60.390 162.310 ;
        RECT 64.300 162.250 64.620 162.310 ;
        RECT 64.760 162.450 65.080 162.510 ;
        RECT 64.760 162.310 67.750 162.450 ;
        RECT 64.760 162.250 65.080 162.310 ;
        RECT 54.195 161.970 60.390 162.110 ;
        RECT 54.195 161.925 54.485 161.970 ;
        RECT 60.620 161.910 60.940 162.170 ;
        RECT 61.080 162.110 61.400 162.170 ;
        RECT 61.080 161.970 65.910 162.110 ;
        RECT 61.080 161.910 61.400 161.970 ;
        RECT 48.215 161.770 48.505 161.815 ;
        RECT 43.110 161.630 45.645 161.770 ;
        RECT 45.990 161.630 48.505 161.770 ;
        RECT 43.110 161.585 43.400 161.630 ;
        RECT 39.920 161.430 40.240 161.490 ;
        RECT 41.300 161.475 41.620 161.490 ;
        RECT 45.430 161.475 45.645 161.630 ;
        RECT 48.215 161.585 48.505 161.630 ;
        RECT 50.500 161.570 50.820 161.830 ;
        RECT 56.940 161.770 57.260 161.830 ;
        RECT 59.255 161.770 59.545 161.815 ;
        RECT 56.940 161.630 59.545 161.770 ;
        RECT 56.940 161.570 57.260 161.630 ;
        RECT 59.255 161.585 59.545 161.630 ;
        RECT 63.395 161.585 63.685 161.815 ;
        RECT 63.855 161.585 64.145 161.815 ;
        RECT 35.320 161.290 40.240 161.430 ;
        RECT 35.320 161.230 35.640 161.290 ;
        RECT 39.920 161.230 40.240 161.290 ;
        RECT 41.250 161.430 41.620 161.475 ;
        RECT 44.510 161.430 44.800 161.475 ;
        RECT 41.250 161.290 44.800 161.430 ;
        RECT 41.250 161.245 41.620 161.290 ;
        RECT 44.510 161.245 44.800 161.290 ;
        RECT 45.430 161.430 45.720 161.475 ;
        RECT 47.290 161.430 47.580 161.475 ;
        RECT 45.430 161.290 47.580 161.430 ;
        RECT 45.430 161.245 45.720 161.290 ;
        RECT 47.290 161.245 47.580 161.290 ;
        RECT 57.400 161.430 57.720 161.490 ;
        RECT 63.470 161.430 63.610 161.585 ;
        RECT 57.400 161.290 63.610 161.430 ;
        RECT 63.930 161.430 64.070 161.585 ;
        RECT 64.300 161.570 64.620 161.830 ;
        RECT 65.220 161.570 65.540 161.830 ;
        RECT 65.770 161.815 65.910 161.970 ;
        RECT 65.695 161.585 65.985 161.815 ;
        RECT 67.075 161.585 67.365 161.815 ;
        RECT 64.760 161.430 65.080 161.490 ;
        RECT 63.930 161.290 65.080 161.430 ;
        RECT 65.310 161.430 65.450 161.570 ;
        RECT 67.150 161.430 67.290 161.585 ;
        RECT 65.310 161.290 67.290 161.430 ;
        RECT 67.610 161.430 67.750 162.310 ;
        RECT 68.070 161.815 68.210 162.650 ;
        RECT 79.480 162.590 79.800 162.650 ;
        RECT 82.700 162.790 83.020 162.850 ;
        RECT 84.555 162.790 84.845 162.835 ;
        RECT 85.000 162.790 85.320 162.850 ;
        RECT 82.700 162.650 84.310 162.790 ;
        RECT 82.700 162.590 83.020 162.650 ;
        RECT 71.660 162.450 71.980 162.510 ;
        RECT 78.530 162.450 78.820 162.495 ;
        RECT 81.310 162.450 81.600 162.495 ;
        RECT 83.170 162.450 83.460 162.495 ;
        RECT 68.530 162.310 72.810 162.450 ;
        RECT 68.530 161.815 68.670 162.310 ;
        RECT 71.660 162.250 71.980 162.310 ;
        RECT 68.990 161.970 72.350 162.110 ;
        RECT 68.990 161.815 69.130 161.970 ;
        RECT 72.210 161.830 72.350 161.970 ;
        RECT 67.995 161.585 68.285 161.815 ;
        RECT 68.455 161.585 68.745 161.815 ;
        RECT 68.915 161.585 69.205 161.815 ;
        RECT 68.530 161.430 68.670 161.585 ;
        RECT 67.610 161.290 68.670 161.430 ;
        RECT 41.300 161.230 41.620 161.245 ;
        RECT 57.400 161.230 57.720 161.290 ;
        RECT 24.525 161.090 24.815 161.135 ;
        RECT 27.500 161.090 27.820 161.150 ;
        RECT 24.525 160.950 27.820 161.090 ;
        RECT 24.525 160.905 24.815 160.950 ;
        RECT 27.500 160.890 27.820 160.950 ;
        RECT 36.700 161.090 37.020 161.150 ;
        RECT 37.635 161.090 37.925 161.135 ;
        RECT 36.700 160.950 37.925 161.090 ;
        RECT 36.700 160.890 37.020 160.950 ;
        RECT 37.635 160.905 37.925 160.950 ;
        RECT 43.600 161.090 43.920 161.150 ;
        RECT 48.675 161.090 48.965 161.135 ;
        RECT 43.600 160.950 48.965 161.090 ;
        RECT 43.600 160.890 43.920 160.950 ;
        RECT 48.675 160.905 48.965 160.950 ;
        RECT 52.800 161.090 53.120 161.150 ;
        RECT 59.715 161.090 60.005 161.135 ;
        RECT 52.800 160.950 60.005 161.090 ;
        RECT 52.800 160.890 53.120 160.950 ;
        RECT 59.715 160.905 60.005 160.950 ;
        RECT 62.000 160.890 62.320 161.150 ;
        RECT 63.470 161.090 63.610 161.290 ;
        RECT 64.760 161.230 65.080 161.290 ;
        RECT 68.990 161.090 69.130 161.585 ;
        RECT 70.740 161.570 71.060 161.830 ;
        RECT 72.120 161.570 72.440 161.830 ;
        RECT 72.670 161.815 72.810 162.310 ;
        RECT 78.530 162.310 83.460 162.450 ;
        RECT 78.530 162.265 78.820 162.310 ;
        RECT 81.310 162.265 81.600 162.310 ;
        RECT 83.170 162.265 83.460 162.310 ;
        RECT 74.665 162.110 74.955 162.155 ;
        RECT 76.720 162.110 77.040 162.170 ;
        RECT 73.130 161.970 77.040 162.110 ;
        RECT 73.130 161.815 73.270 161.970 ;
        RECT 74.665 161.925 74.955 161.970 ;
        RECT 76.720 161.910 77.040 161.970 ;
        RECT 83.620 161.910 83.940 162.170 ;
        RECT 84.170 162.110 84.310 162.650 ;
        RECT 84.555 162.650 85.320 162.790 ;
        RECT 84.555 162.605 84.845 162.650 ;
        RECT 85.000 162.590 85.320 162.650 ;
        RECT 86.855 162.790 87.145 162.835 ;
        RECT 87.760 162.790 88.080 162.850 ;
        RECT 92.360 162.790 92.680 162.850 ;
        RECT 94.200 162.790 94.520 162.850 ;
        RECT 86.855 162.650 88.080 162.790 ;
        RECT 86.855 162.605 87.145 162.650 ;
        RECT 87.760 162.590 88.080 162.650 ;
        RECT 90.150 162.650 94.520 162.790 ;
        RECT 90.150 162.110 90.290 162.650 ;
        RECT 92.360 162.590 92.680 162.650 ;
        RECT 94.200 162.590 94.520 162.650 ;
        RECT 101.575 162.790 101.865 162.835 ;
        RECT 103.400 162.790 103.720 162.850 ;
        RECT 101.575 162.650 103.720 162.790 ;
        RECT 101.575 162.605 101.865 162.650 ;
        RECT 103.400 162.590 103.720 162.650 ;
        RECT 90.520 162.450 90.840 162.510 ;
        RECT 96.515 162.450 96.805 162.495 ;
        RECT 90.520 162.310 96.805 162.450 ;
        RECT 90.520 162.250 90.840 162.310 ;
        RECT 96.515 162.265 96.805 162.310 ;
        RECT 98.340 162.450 98.660 162.510 ;
        RECT 102.960 162.450 103.250 162.495 ;
        RECT 104.820 162.450 105.110 162.495 ;
        RECT 107.600 162.450 107.890 162.495 ;
        RECT 98.340 162.310 102.710 162.450 ;
        RECT 98.340 162.250 98.660 162.310 ;
        RECT 102.570 162.155 102.710 162.310 ;
        RECT 102.960 162.310 107.890 162.450 ;
        RECT 102.960 162.265 103.250 162.310 ;
        RECT 104.820 162.265 105.110 162.310 ;
        RECT 107.600 162.265 107.890 162.310 ;
        RECT 84.170 161.970 90.750 162.110 ;
        RECT 72.595 161.585 72.885 161.815 ;
        RECT 73.055 161.585 73.345 161.815 ;
        RECT 73.975 161.585 74.265 161.815 ;
        RECT 78.530 161.770 78.820 161.815 ;
        RECT 78.530 161.630 81.065 161.770 ;
        RECT 78.530 161.585 78.820 161.630 ;
        RECT 70.830 161.430 70.970 161.570 ;
        RECT 74.050 161.430 74.190 161.585 ;
        RECT 70.830 161.290 74.190 161.430 ;
        RECT 76.670 161.430 76.960 161.475 ;
        RECT 79.020 161.430 79.340 161.490 ;
        RECT 80.850 161.475 81.065 161.630 ;
        RECT 81.780 161.570 82.100 161.830 ;
        RECT 85.015 161.595 85.305 161.825 ;
        RECT 79.930 161.430 80.220 161.475 ;
        RECT 76.670 161.290 80.220 161.430 ;
        RECT 76.670 161.245 76.960 161.290 ;
        RECT 79.020 161.230 79.340 161.290 ;
        RECT 79.930 161.245 80.220 161.290 ;
        RECT 80.850 161.430 81.140 161.475 ;
        RECT 82.710 161.430 83.000 161.475 ;
        RECT 80.850 161.290 83.000 161.430 ;
        RECT 80.850 161.245 81.140 161.290 ;
        RECT 82.710 161.245 83.000 161.290 ;
        RECT 83.160 161.430 83.480 161.490 ;
        RECT 85.090 161.430 85.230 161.595 ;
        RECT 85.920 161.570 86.240 161.830 ;
        RECT 90.610 161.815 90.750 161.970 ;
        RECT 91.070 161.970 98.570 162.110 ;
        RECT 91.070 161.830 91.210 161.970 ;
        RECT 94.750 161.830 94.890 161.970 ;
        RECT 90.535 161.585 90.825 161.815 ;
        RECT 90.980 161.570 91.300 161.830 ;
        RECT 91.455 161.770 91.745 161.815 ;
        RECT 91.900 161.770 92.220 161.830 ;
        RECT 91.455 161.630 92.220 161.770 ;
        RECT 91.455 161.585 91.745 161.630 ;
        RECT 91.900 161.570 92.220 161.630 ;
        RECT 92.375 161.770 92.665 161.815 ;
        RECT 93.740 161.770 94.060 161.830 ;
        RECT 92.375 161.630 94.060 161.770 ;
        RECT 92.375 161.585 92.665 161.630 ;
        RECT 88.220 161.430 88.540 161.490 ;
        RECT 92.450 161.430 92.590 161.585 ;
        RECT 93.740 161.570 94.060 161.630 ;
        RECT 94.200 161.570 94.520 161.830 ;
        RECT 94.660 161.570 94.980 161.830 ;
        RECT 95.120 161.570 95.440 161.830 ;
        RECT 96.055 161.585 96.345 161.815 ;
        RECT 83.160 161.290 88.540 161.430 ;
        RECT 83.160 161.230 83.480 161.290 ;
        RECT 88.220 161.230 88.540 161.290 ;
        RECT 88.770 161.290 92.590 161.430 ;
        RECT 93.830 161.430 93.970 161.570 ;
        RECT 96.130 161.430 96.270 161.585 ;
        RECT 97.880 161.570 98.200 161.830 ;
        RECT 98.430 161.815 98.570 161.970 ;
        RECT 102.495 161.925 102.785 162.155 ;
        RECT 104.320 161.910 104.640 162.170 ;
        RECT 98.355 161.585 98.645 161.815 ;
        RECT 98.815 161.770 99.105 161.815 ;
        RECT 99.260 161.770 99.580 161.830 ;
        RECT 98.815 161.630 99.580 161.770 ;
        RECT 98.815 161.585 99.105 161.630 ;
        RECT 99.260 161.570 99.580 161.630 ;
        RECT 99.735 161.585 100.025 161.815 ;
        RECT 96.500 161.430 96.820 161.490 ;
        RECT 99.810 161.430 99.950 161.585 ;
        RECT 101.100 161.570 101.420 161.830 ;
        RECT 107.600 161.770 107.890 161.815 ;
        RECT 105.355 161.630 107.890 161.770 ;
        RECT 105.355 161.475 105.570 161.630 ;
        RECT 107.600 161.585 107.890 161.630 ;
        RECT 93.830 161.290 99.950 161.430 ;
        RECT 103.420 161.430 103.710 161.475 ;
        RECT 105.280 161.430 105.570 161.475 ;
        RECT 103.420 161.290 105.570 161.430 ;
        RECT 63.470 160.950 69.130 161.090 ;
        RECT 70.280 160.890 70.600 161.150 ;
        RECT 70.755 161.090 71.045 161.135 ;
        RECT 73.040 161.090 73.360 161.150 ;
        RECT 70.755 160.950 73.360 161.090 ;
        RECT 70.755 160.905 71.045 160.950 ;
        RECT 73.040 160.890 73.360 160.950 ;
        RECT 78.560 161.090 78.880 161.150 ;
        RECT 88.770 161.090 88.910 161.290 ;
        RECT 96.500 161.230 96.820 161.290 ;
        RECT 103.420 161.245 103.710 161.290 ;
        RECT 105.280 161.245 105.570 161.290 ;
        RECT 106.160 161.475 106.480 161.490 ;
        RECT 106.160 161.430 106.490 161.475 ;
        RECT 109.460 161.430 109.750 161.475 ;
        RECT 106.160 161.290 109.750 161.430 ;
        RECT 106.160 161.245 106.490 161.290 ;
        RECT 109.460 161.245 109.750 161.290 ;
        RECT 106.160 161.230 106.480 161.245 ;
        RECT 78.560 160.950 88.910 161.090 ;
        RECT 89.155 161.090 89.445 161.135 ;
        RECT 90.980 161.090 91.300 161.150 ;
        RECT 89.155 160.950 91.300 161.090 ;
        RECT 78.560 160.890 78.880 160.950 ;
        RECT 89.155 160.905 89.445 160.950 ;
        RECT 90.980 160.890 91.300 160.950 ;
        RECT 91.900 161.090 92.220 161.150 ;
        RECT 92.835 161.090 93.125 161.135 ;
        RECT 91.900 160.950 93.125 161.090 ;
        RECT 91.900 160.890 92.220 160.950 ;
        RECT 92.835 160.905 93.125 160.950 ;
        RECT 108.000 161.090 108.320 161.150 ;
        RECT 111.465 161.090 111.755 161.135 ;
        RECT 108.000 160.950 111.755 161.090 ;
        RECT 108.000 160.890 108.320 160.950 ;
        RECT 111.465 160.905 111.755 160.950 ;
        RECT 22.830 160.270 113.450 160.750 ;
        RECT 38.540 160.070 38.860 160.130 ;
        RECT 39.015 160.070 39.305 160.115 ;
        RECT 38.540 159.930 39.305 160.070 ;
        RECT 38.540 159.870 38.860 159.930 ;
        RECT 39.015 159.885 39.305 159.930 ;
        RECT 40.840 159.870 41.160 160.130 ;
        RECT 44.535 160.070 44.825 160.115 ;
        RECT 46.360 160.070 46.680 160.130 ;
        RECT 44.535 159.930 46.680 160.070 ;
        RECT 44.535 159.885 44.825 159.930 ;
        RECT 46.360 159.870 46.680 159.930 ;
        RECT 46.820 160.070 47.140 160.130 ;
        RECT 52.800 160.070 53.120 160.130 ;
        RECT 69.375 160.070 69.665 160.115 ;
        RECT 70.740 160.070 71.060 160.130 ;
        RECT 46.820 159.930 51.650 160.070 ;
        RECT 46.820 159.870 47.140 159.930 ;
        RECT 26.595 159.730 26.885 159.775 ;
        RECT 27.500 159.730 27.820 159.790 ;
        RECT 31.640 159.775 31.960 159.790 ;
        RECT 26.595 159.590 27.820 159.730 ;
        RECT 26.595 159.545 26.885 159.590 ;
        RECT 27.500 159.530 27.820 159.590 ;
        RECT 31.590 159.730 31.960 159.775 ;
        RECT 34.850 159.730 35.140 159.775 ;
        RECT 31.590 159.590 35.140 159.730 ;
        RECT 31.590 159.545 31.960 159.590 ;
        RECT 34.850 159.545 35.140 159.590 ;
        RECT 35.770 159.730 36.060 159.775 ;
        RECT 37.630 159.730 37.920 159.775 ;
        RECT 35.770 159.590 37.920 159.730 ;
        RECT 35.770 159.545 36.060 159.590 ;
        RECT 37.630 159.545 37.920 159.590 ;
        RECT 44.060 159.730 44.380 159.790 ;
        RECT 51.510 159.730 51.650 159.930 ;
        RECT 52.800 159.930 54.410 160.070 ;
        RECT 52.800 159.870 53.120 159.930 ;
        RECT 44.060 159.590 46.130 159.730 ;
        RECT 31.640 159.530 31.960 159.545 ;
        RECT 27.055 159.205 27.345 159.435 ;
        RECT 33.450 159.390 33.740 159.435 ;
        RECT 35.770 159.390 35.985 159.545 ;
        RECT 44.060 159.530 44.380 159.590 ;
        RECT 33.450 159.250 35.985 159.390 ;
        RECT 33.450 159.205 33.740 159.250 ;
        RECT 26.135 158.865 26.425 159.095 ;
        RECT 27.130 159.050 27.270 159.205 ;
        RECT 36.700 159.190 37.020 159.450 ;
        RECT 38.080 159.390 38.400 159.450 ;
        RECT 38.555 159.390 38.845 159.435 ;
        RECT 38.080 159.250 38.845 159.390 ;
        RECT 38.080 159.190 38.400 159.250 ;
        RECT 38.555 159.205 38.845 159.250 ;
        RECT 40.380 159.390 40.700 159.450 ;
        RECT 40.380 159.250 43.370 159.390 ;
        RECT 40.380 159.190 40.700 159.250 ;
        RECT 29.585 159.050 29.875 159.095 ;
        RECT 41.300 159.050 41.620 159.110 ;
        RECT 27.130 158.910 41.620 159.050 ;
        RECT 29.585 158.865 29.875 158.910 ;
        RECT 26.210 158.710 26.350 158.865 ;
        RECT 41.300 158.850 41.620 158.910 ;
        RECT 41.775 158.865 42.065 159.095 ;
        RECT 43.230 159.050 43.370 159.250 ;
        RECT 43.600 159.190 43.920 159.450 ;
        RECT 44.980 159.190 45.300 159.450 ;
        RECT 45.990 159.435 46.130 159.590 ;
        RECT 46.910 159.590 51.190 159.730 ;
        RECT 51.510 159.590 53.950 159.730 ;
        RECT 45.915 159.205 46.205 159.435 ;
        RECT 46.360 159.190 46.680 159.450 ;
        RECT 46.910 159.435 47.050 159.590 ;
        RECT 46.835 159.205 47.125 159.435 ;
        RECT 50.040 159.390 50.360 159.450 ;
        RECT 50.515 159.390 50.805 159.435 ;
        RECT 50.040 159.250 50.805 159.390 ;
        RECT 51.050 159.390 51.190 159.590 ;
        RECT 53.810 159.435 53.950 159.590 ;
        RECT 54.270 159.435 54.410 159.930 ;
        RECT 65.310 159.930 71.060 160.070 ;
        RECT 65.310 159.790 65.450 159.930 ;
        RECT 69.375 159.885 69.665 159.930 ;
        RECT 70.740 159.870 71.060 159.930 ;
        RECT 80.875 160.070 81.165 160.115 ;
        RECT 81.780 160.070 82.100 160.130 ;
        RECT 80.875 159.930 82.100 160.070 ;
        RECT 80.875 159.885 81.165 159.930 ;
        RECT 81.780 159.870 82.100 159.930 ;
        RECT 82.700 160.070 83.020 160.130 ;
        RECT 93.740 160.070 94.060 160.130 ;
        RECT 97.880 160.070 98.200 160.130 ;
        RECT 82.700 159.930 94.060 160.070 ;
        RECT 82.700 159.870 83.020 159.930 ;
        RECT 93.740 159.870 94.060 159.930 ;
        RECT 94.290 159.930 98.200 160.070 ;
        RECT 65.220 159.730 65.540 159.790 ;
        RECT 55.650 159.590 65.540 159.730 ;
        RECT 55.650 159.450 55.790 159.590 ;
        RECT 65.220 159.530 65.540 159.590 ;
        RECT 67.980 159.530 68.300 159.790 ;
        RECT 70.830 159.730 70.970 159.870 ;
        RECT 70.830 159.590 74.190 159.730 ;
        RECT 53.275 159.405 53.565 159.435 ;
        RECT 52.430 159.390 53.565 159.405 ;
        RECT 51.050 159.265 53.565 159.390 ;
        RECT 51.050 159.250 52.570 159.265 ;
        RECT 46.910 159.050 47.050 159.205 ;
        RECT 50.040 159.190 50.360 159.250 ;
        RECT 50.515 159.205 50.805 159.250 ;
        RECT 43.230 158.910 47.050 159.050 ;
        RECT 33.450 158.710 33.740 158.755 ;
        RECT 36.230 158.710 36.520 158.755 ;
        RECT 38.090 158.710 38.380 158.755 ;
        RECT 41.850 158.710 41.990 158.865 ;
        RECT 26.210 158.570 30.030 158.710 ;
        RECT 29.890 158.430 30.030 158.570 ;
        RECT 33.450 158.570 38.380 158.710 ;
        RECT 33.450 158.525 33.740 158.570 ;
        RECT 36.230 158.525 36.520 158.570 ;
        RECT 38.090 158.525 38.380 158.570 ;
        RECT 41.390 158.570 41.990 158.710 ;
        RECT 44.980 158.710 45.300 158.770 ;
        RECT 51.895 158.710 52.185 158.755 ;
        RECT 44.980 158.570 52.185 158.710 ;
        RECT 52.890 158.710 53.030 159.265 ;
        RECT 53.275 159.205 53.565 159.265 ;
        RECT 53.735 159.205 54.025 159.435 ;
        RECT 54.195 159.205 54.485 159.435 ;
        RECT 55.115 159.390 55.405 159.435 ;
        RECT 55.560 159.390 55.880 159.450 ;
        RECT 55.115 159.250 55.880 159.390 ;
        RECT 55.115 159.205 55.405 159.250 ;
        RECT 53.810 159.050 53.950 159.205 ;
        RECT 55.560 159.190 55.880 159.250 ;
        RECT 56.480 159.190 56.800 159.450 ;
        RECT 56.955 159.205 57.245 159.435 ;
        RECT 57.030 159.050 57.170 159.205 ;
        RECT 57.400 159.190 57.720 159.450 ;
        RECT 65.680 159.390 66.000 159.450 ;
        RECT 68.455 159.390 68.745 159.435 ;
        RECT 70.740 159.390 71.060 159.450 ;
        RECT 65.680 159.250 71.060 159.390 ;
        RECT 65.680 159.190 66.000 159.250 ;
        RECT 68.455 159.205 68.745 159.250 ;
        RECT 70.740 159.190 71.060 159.250 ;
        RECT 72.120 159.190 72.440 159.450 ;
        RECT 72.595 159.205 72.885 159.435 ;
        RECT 73.055 159.390 73.345 159.435 ;
        RECT 73.500 159.390 73.820 159.450 ;
        RECT 74.050 159.435 74.190 159.590 ;
        RECT 79.020 159.530 79.340 159.790 ;
        RECT 83.160 159.730 83.480 159.790 ;
        RECT 79.570 159.590 83.480 159.730 ;
        RECT 73.055 159.250 73.820 159.390 ;
        RECT 73.055 159.205 73.345 159.250 ;
        RECT 64.760 159.050 65.080 159.110 ;
        RECT 53.810 158.910 65.080 159.050 ;
        RECT 64.760 158.850 65.080 158.910 ;
        RECT 71.660 159.050 71.980 159.110 ;
        RECT 72.670 159.050 72.810 159.205 ;
        RECT 73.500 159.190 73.820 159.250 ;
        RECT 73.975 159.205 74.265 159.435 ;
        RECT 74.880 159.190 75.200 159.450 ;
        RECT 79.570 159.435 79.710 159.590 ;
        RECT 83.160 159.530 83.480 159.590 ;
        RECT 84.195 159.730 84.485 159.775 ;
        RECT 87.435 159.730 88.085 159.775 ;
        RECT 84.195 159.590 88.085 159.730 ;
        RECT 84.195 159.545 84.785 159.590 ;
        RECT 87.435 159.545 88.085 159.590 ;
        RECT 78.115 159.390 78.405 159.435 ;
        RECT 79.495 159.390 79.785 159.435 ;
        RECT 78.115 159.250 79.785 159.390 ;
        RECT 78.115 159.205 78.405 159.250 ;
        RECT 79.495 159.205 79.785 159.250 ;
        RECT 79.940 159.190 80.260 159.450 ;
        RECT 81.335 159.390 81.625 159.435 ;
        RECT 82.240 159.390 82.560 159.450 ;
        RECT 81.335 159.250 82.560 159.390 ;
        RECT 81.335 159.205 81.625 159.250 ;
        RECT 82.240 159.190 82.560 159.250 ;
        RECT 84.495 159.230 84.785 159.545 ;
        RECT 90.060 159.530 90.380 159.790 ;
        RECT 94.290 159.435 94.430 159.930 ;
        RECT 97.880 159.870 98.200 159.930 ;
        RECT 103.400 159.870 103.720 160.130 ;
        RECT 105.240 160.070 105.560 160.130 ;
        RECT 104.410 159.930 105.560 160.070 ;
        RECT 104.410 159.730 104.550 159.930 ;
        RECT 105.240 159.870 105.560 159.930 ;
        RECT 105.700 160.070 106.020 160.130 ;
        RECT 108.000 160.070 108.320 160.130 ;
        RECT 105.700 159.930 108.320 160.070 ;
        RECT 105.700 159.870 106.020 159.930 ;
        RECT 108.000 159.870 108.320 159.930 ;
        RECT 109.840 159.870 110.160 160.130 ;
        RECT 107.555 159.730 107.845 159.775 ;
        RECT 95.210 159.590 104.550 159.730 ;
        RECT 105.100 159.590 107.845 159.730 ;
        RECT 85.575 159.390 85.865 159.435 ;
        RECT 89.155 159.390 89.445 159.435 ;
        RECT 90.990 159.390 91.280 159.435 ;
        RECT 85.575 159.250 91.280 159.390 ;
        RECT 71.660 158.910 72.810 159.050 ;
        RECT 77.655 159.050 77.945 159.095 ;
        RECT 84.630 159.050 84.770 159.230 ;
        RECT 85.575 159.205 85.865 159.250 ;
        RECT 89.155 159.205 89.445 159.250 ;
        RECT 90.990 159.205 91.280 159.250 ;
        RECT 94.215 159.205 94.505 159.435 ;
        RECT 94.660 159.190 94.980 159.450 ;
        RECT 95.210 159.435 95.350 159.590 ;
        RECT 95.135 159.205 95.425 159.435 ;
        RECT 96.055 159.390 96.345 159.435 ;
        RECT 96.500 159.390 96.820 159.450 ;
        RECT 96.055 159.250 96.820 159.390 ;
        RECT 96.055 159.205 96.345 159.250 ;
        RECT 96.500 159.190 96.820 159.250 ;
        RECT 97.880 159.190 98.200 159.450 ;
        RECT 98.355 159.205 98.645 159.435 ;
        RECT 77.655 158.910 84.770 159.050 ;
        RECT 89.600 159.050 89.920 159.110 ;
        RECT 91.455 159.050 91.745 159.095 ;
        RECT 89.600 158.910 91.745 159.050 ;
        RECT 98.430 159.050 98.570 159.205 ;
        RECT 98.800 159.190 99.120 159.450 ;
        RECT 99.720 159.190 100.040 159.450 ;
        RECT 102.940 159.390 103.260 159.450 ;
        RECT 105.100 159.390 105.240 159.590 ;
        RECT 107.555 159.545 107.845 159.590 ;
        RECT 102.940 159.250 105.240 159.390 ;
        RECT 110.300 159.390 110.620 159.450 ;
        RECT 110.775 159.390 111.065 159.435 ;
        RECT 110.300 159.250 111.065 159.390 ;
        RECT 102.940 159.190 103.260 159.250 ;
        RECT 110.300 159.190 110.620 159.250 ;
        RECT 110.775 159.205 111.065 159.250 ;
        RECT 100.180 159.050 100.500 159.110 ;
        RECT 98.430 158.910 100.500 159.050 ;
        RECT 71.660 158.850 71.980 158.910 ;
        RECT 77.655 158.865 77.945 158.910 ;
        RECT 89.600 158.850 89.920 158.910 ;
        RECT 91.455 158.865 91.745 158.910 ;
        RECT 100.180 158.850 100.500 158.910 ;
        RECT 102.495 159.050 102.785 159.095 ;
        RECT 103.860 159.050 104.180 159.110 ;
        RECT 108.475 159.050 108.765 159.095 ;
        RECT 102.495 158.910 108.765 159.050 ;
        RECT 102.495 158.865 102.785 158.910 ;
        RECT 103.860 158.850 104.180 158.910 ;
        RECT 108.475 158.865 108.765 158.910 ;
        RECT 57.400 158.710 57.720 158.770 ;
        RECT 52.890 158.570 57.720 158.710 ;
        RECT 28.895 158.370 29.185 158.415 ;
        RECT 29.340 158.370 29.660 158.430 ;
        RECT 28.895 158.230 29.660 158.370 ;
        RECT 28.895 158.185 29.185 158.230 ;
        RECT 29.340 158.170 29.660 158.230 ;
        RECT 29.800 158.370 30.120 158.430 ;
        RECT 41.390 158.370 41.530 158.570 ;
        RECT 44.980 158.510 45.300 158.570 ;
        RECT 51.895 158.525 52.185 158.570 ;
        RECT 57.400 158.510 57.720 158.570 ;
        RECT 61.540 158.510 61.860 158.770 ;
        RECT 62.460 158.710 62.780 158.770 ;
        RECT 75.815 158.710 76.105 158.755 ;
        RECT 78.560 158.710 78.880 158.770 ;
        RECT 62.460 158.570 78.880 158.710 ;
        RECT 62.460 158.510 62.780 158.570 ;
        RECT 75.815 158.525 76.105 158.570 ;
        RECT 78.560 158.510 78.880 158.570 ;
        RECT 85.575 158.710 85.865 158.755 ;
        RECT 88.695 158.710 88.985 158.755 ;
        RECT 90.585 158.710 90.875 158.755 ;
        RECT 85.575 158.570 90.875 158.710 ;
        RECT 85.575 158.525 85.865 158.570 ;
        RECT 88.695 158.525 88.985 158.570 ;
        RECT 90.585 158.525 90.875 158.570 ;
        RECT 95.580 158.710 95.900 158.770 ;
        RECT 97.880 158.710 98.200 158.770 ;
        RECT 95.580 158.570 98.200 158.710 ;
        RECT 95.580 158.510 95.900 158.570 ;
        RECT 97.880 158.510 98.200 158.570 ;
        RECT 101.560 158.710 101.880 158.770 ;
        RECT 105.715 158.710 106.005 158.755 ;
        RECT 101.560 158.570 106.005 158.710 ;
        RECT 101.560 158.510 101.880 158.570 ;
        RECT 105.715 158.525 106.005 158.570 ;
        RECT 29.800 158.230 41.530 158.370 ;
        RECT 44.520 158.370 44.840 158.430 ;
        RECT 46.360 158.370 46.680 158.430 ;
        RECT 44.520 158.230 46.680 158.370 ;
        RECT 29.800 158.170 30.120 158.230 ;
        RECT 44.520 158.170 44.840 158.230 ;
        RECT 46.360 158.170 46.680 158.230 ;
        RECT 48.215 158.370 48.505 158.415 ;
        RECT 49.580 158.370 49.900 158.430 ;
        RECT 48.215 158.230 49.900 158.370 ;
        RECT 48.215 158.185 48.505 158.230 ;
        RECT 49.580 158.170 49.900 158.230 ;
        RECT 51.420 158.170 51.740 158.430 ;
        RECT 58.780 158.170 59.100 158.430 ;
        RECT 70.755 158.370 71.045 158.415 ;
        RECT 71.660 158.370 71.980 158.430 ;
        RECT 70.755 158.230 71.980 158.370 ;
        RECT 70.755 158.185 71.045 158.230 ;
        RECT 71.660 158.170 71.980 158.230 ;
        RECT 82.255 158.370 82.545 158.415 ;
        RECT 84.540 158.370 84.860 158.430 ;
        RECT 82.255 158.230 84.860 158.370 ;
        RECT 82.255 158.185 82.545 158.230 ;
        RECT 84.540 158.170 84.860 158.230 ;
        RECT 92.835 158.370 93.125 158.415 ;
        RECT 94.660 158.370 94.980 158.430 ;
        RECT 92.835 158.230 94.980 158.370 ;
        RECT 92.835 158.185 93.125 158.230 ;
        RECT 94.660 158.170 94.980 158.230 ;
        RECT 96.500 158.170 96.820 158.430 ;
        RECT 105.240 158.170 105.560 158.430 ;
        RECT 22.830 157.550 113.450 158.030 ;
        RECT 28.435 157.350 28.725 157.395 ;
        RECT 28.880 157.350 29.200 157.410 ;
        RECT 28.435 157.210 29.200 157.350 ;
        RECT 28.435 157.165 28.725 157.210 ;
        RECT 28.880 157.150 29.200 157.210 ;
        RECT 30.260 157.150 30.580 157.410 ;
        RECT 31.195 157.350 31.485 157.395 ;
        RECT 31.640 157.350 31.960 157.410 ;
        RECT 31.195 157.210 31.960 157.350 ;
        RECT 31.195 157.165 31.485 157.210 ;
        RECT 31.640 157.150 31.960 157.210 ;
        RECT 33.480 157.350 33.800 157.410 ;
        RECT 57.400 157.350 57.720 157.410 ;
        RECT 63.855 157.350 64.145 157.395 ;
        RECT 33.480 157.210 39.230 157.350 ;
        RECT 33.480 157.150 33.800 157.210 ;
        RECT 35.320 157.010 35.640 157.070 ;
        RECT 30.810 156.870 35.640 157.010 ;
        RECT 30.810 156.670 30.950 156.870 ;
        RECT 35.320 156.810 35.640 156.870 ;
        RECT 39.090 156.730 39.230 157.210 ;
        RECT 57.400 157.210 64.145 157.350 ;
        RECT 57.400 157.150 57.720 157.210 ;
        RECT 63.855 157.165 64.145 157.210 ;
        RECT 71.200 157.150 71.520 157.410 ;
        RECT 74.435 157.350 74.725 157.395 ;
        RECT 71.750 157.210 74.725 157.350 ;
        RECT 45.900 157.010 46.220 157.070 ;
        RECT 40.930 156.870 46.220 157.010 ;
        RECT 28.970 156.530 30.950 156.670 ;
        RECT 28.970 156.375 29.110 156.530 ;
        RECT 28.895 156.145 29.185 156.375 ;
        RECT 29.340 156.130 29.660 156.390 ;
        RECT 30.810 156.375 30.950 156.530 ;
        RECT 31.180 156.670 31.500 156.730 ;
        RECT 38.540 156.670 38.860 156.730 ;
        RECT 31.180 156.530 38.860 156.670 ;
        RECT 31.180 156.470 31.500 156.530 ;
        RECT 38.540 156.470 38.860 156.530 ;
        RECT 39.000 156.670 39.320 156.730 ;
        RECT 40.930 156.670 41.070 156.870 ;
        RECT 45.900 156.810 46.220 156.870 ;
        RECT 50.470 157.010 50.760 157.055 ;
        RECT 53.250 157.010 53.540 157.055 ;
        RECT 55.110 157.010 55.400 157.055 ;
        RECT 50.470 156.870 55.400 157.010 ;
        RECT 50.470 156.825 50.760 156.870 ;
        RECT 53.250 156.825 53.540 156.870 ;
        RECT 55.110 156.825 55.400 156.870 ;
        RECT 56.480 157.010 56.800 157.070 ;
        RECT 71.750 157.010 71.890 157.210 ;
        RECT 74.435 157.165 74.725 157.210 ;
        RECT 73.960 157.010 74.280 157.070 ;
        RECT 56.480 156.870 71.890 157.010 ;
        RECT 72.210 156.870 74.280 157.010 ;
        RECT 74.510 157.010 74.650 157.165 ;
        RECT 88.220 157.150 88.540 157.410 ;
        RECT 92.360 157.150 92.680 157.410 ;
        RECT 98.340 157.350 98.660 157.410 ;
        RECT 99.260 157.350 99.580 157.410 ;
        RECT 92.910 157.210 99.580 157.350 ;
        RECT 92.910 157.010 93.050 157.210 ;
        RECT 98.340 157.150 98.660 157.210 ;
        RECT 99.260 157.150 99.580 157.210 ;
        RECT 110.300 157.150 110.620 157.410 ;
        RECT 74.510 156.870 93.050 157.010 ;
        RECT 56.480 156.810 56.800 156.870 ;
        RECT 46.820 156.670 47.140 156.730 ;
        RECT 50.960 156.670 51.280 156.730 ;
        RECT 39.000 156.530 41.070 156.670 ;
        RECT 43.690 156.530 47.140 156.670 ;
        RECT 39.000 156.470 39.320 156.530 ;
        RECT 30.735 156.145 31.025 156.375 ;
        RECT 32.115 156.145 32.405 156.375 ;
        RECT 32.560 156.330 32.880 156.390 ;
        RECT 33.035 156.330 33.325 156.375 ;
        RECT 32.560 156.190 33.325 156.330 ;
        RECT 32.190 155.990 32.330 156.145 ;
        RECT 32.560 156.130 32.880 156.190 ;
        RECT 33.035 156.145 33.325 156.190 ;
        RECT 33.480 156.130 33.800 156.390 ;
        RECT 33.955 156.330 34.245 156.375 ;
        RECT 39.460 156.330 39.780 156.390 ;
        RECT 40.470 156.375 40.610 156.530 ;
        RECT 39.935 156.330 40.225 156.375 ;
        RECT 33.955 156.190 40.225 156.330 ;
        RECT 33.955 156.145 34.245 156.190 ;
        RECT 39.460 156.130 39.780 156.190 ;
        RECT 39.935 156.145 40.225 156.190 ;
        RECT 40.395 156.145 40.685 156.375 ;
        RECT 40.855 156.330 41.145 156.375 ;
        RECT 41.300 156.330 41.620 156.390 ;
        RECT 40.855 156.190 41.620 156.330 ;
        RECT 40.855 156.145 41.145 156.190 ;
        RECT 41.300 156.130 41.620 156.190 ;
        RECT 41.760 156.130 42.080 156.390 ;
        RECT 43.690 156.330 43.830 156.530 ;
        RECT 46.820 156.470 47.140 156.530 ;
        RECT 49.670 156.530 51.280 156.670 ;
        RECT 43.975 156.330 44.265 156.375 ;
        RECT 43.690 156.190 44.265 156.330 ;
        RECT 43.975 156.145 44.265 156.190 ;
        RECT 44.520 156.130 44.840 156.390 ;
        RECT 44.995 156.130 45.285 156.360 ;
        RECT 45.900 156.330 46.220 156.390 ;
        RECT 49.670 156.330 49.810 156.530 ;
        RECT 50.960 156.470 51.280 156.530 ;
        RECT 51.420 156.670 51.740 156.730 ;
        RECT 53.735 156.670 54.025 156.715 ;
        RECT 51.420 156.530 54.025 156.670 ;
        RECT 51.420 156.470 51.740 156.530 ;
        RECT 53.735 156.485 54.025 156.530 ;
        RECT 54.180 156.670 54.500 156.730 ;
        RECT 68.440 156.670 68.760 156.730 ;
        RECT 71.200 156.670 71.520 156.730 ;
        RECT 72.210 156.715 72.350 156.870 ;
        RECT 73.960 156.810 74.280 156.870 ;
        RECT 54.180 156.530 60.390 156.670 ;
        RECT 54.180 156.470 54.500 156.530 ;
        RECT 45.900 156.190 49.810 156.330 ;
        RECT 50.470 156.330 50.760 156.375 ;
        RECT 50.470 156.190 53.005 156.330 ;
        RECT 45.900 156.130 46.220 156.190 ;
        RECT 50.470 156.145 50.760 156.190 ;
        RECT 41.850 155.990 41.990 156.130 ;
        RECT 32.190 155.850 41.990 155.990 ;
        RECT 45.070 155.990 45.210 156.130 ;
        RECT 52.790 156.035 53.005 156.190 ;
        RECT 55.560 156.130 55.880 156.390 ;
        RECT 56.035 156.330 56.325 156.375 ;
        RECT 56.800 156.330 56.940 156.530 ;
        RECT 60.250 156.390 60.390 156.530 ;
        RECT 64.850 156.530 68.760 156.670 ;
        RECT 56.035 156.190 56.940 156.330 ;
        RECT 56.035 156.145 56.325 156.190 ;
        RECT 57.400 156.130 57.720 156.390 ;
        RECT 60.160 156.330 60.480 156.390 ;
        RECT 64.850 156.375 64.990 156.530 ;
        RECT 68.440 156.470 68.760 156.530 ;
        RECT 68.990 156.530 71.520 156.670 ;
        RECT 62.935 156.330 63.225 156.375 ;
        RECT 60.160 156.190 63.225 156.330 ;
        RECT 60.160 156.130 60.480 156.190 ;
        RECT 62.935 156.145 63.225 156.190 ;
        RECT 64.775 156.145 65.065 156.375 ;
        RECT 65.235 156.330 65.525 156.375 ;
        RECT 65.680 156.330 66.000 156.390 ;
        RECT 68.990 156.375 69.130 156.530 ;
        RECT 71.200 156.470 71.520 156.530 ;
        RECT 72.135 156.485 72.425 156.715 ;
        RECT 72.595 156.670 72.885 156.715 ;
        RECT 74.880 156.670 75.200 156.730 ;
        RECT 72.595 156.530 75.200 156.670 ;
        RECT 72.595 156.485 72.885 156.530 ;
        RECT 65.235 156.190 66.000 156.330 ;
        RECT 65.235 156.145 65.525 156.190 ;
        RECT 65.680 156.130 66.000 156.190 ;
        RECT 67.075 156.145 67.365 156.375 ;
        RECT 68.915 156.145 69.205 156.375 ;
        RECT 69.360 156.330 69.680 156.390 ;
        RECT 70.755 156.330 71.045 156.375 ;
        RECT 73.515 156.330 73.805 156.375 ;
        RECT 69.360 156.190 73.805 156.330 ;
        RECT 48.610 155.990 48.900 156.035 ;
        RECT 51.870 155.990 52.160 156.035 ;
        RECT 52.790 155.990 53.080 156.035 ;
        RECT 54.650 155.990 54.940 156.035 ;
        RECT 62.475 155.990 62.765 156.035 ;
        RECT 45.070 155.850 46.130 155.990 ;
        RECT 45.990 155.710 46.130 155.850 ;
        RECT 48.610 155.850 52.570 155.990 ;
        RECT 48.610 155.805 48.900 155.850 ;
        RECT 51.870 155.805 52.160 155.850 ;
        RECT 35.335 155.650 35.625 155.695 ;
        RECT 35.780 155.650 36.100 155.710 ;
        RECT 35.335 155.510 36.100 155.650 ;
        RECT 35.335 155.465 35.625 155.510 ;
        RECT 35.780 155.450 36.100 155.510 ;
        RECT 38.555 155.650 38.845 155.695 ;
        RECT 39.920 155.650 40.240 155.710 ;
        RECT 38.555 155.510 40.240 155.650 ;
        RECT 38.555 155.465 38.845 155.510 ;
        RECT 39.920 155.450 40.240 155.510 ;
        RECT 42.680 155.450 43.000 155.710 ;
        RECT 45.900 155.650 46.220 155.710 ;
        RECT 46.605 155.650 46.895 155.695 ;
        RECT 45.900 155.510 46.895 155.650 ;
        RECT 52.430 155.650 52.570 155.850 ;
        RECT 52.790 155.850 54.940 155.990 ;
        RECT 52.790 155.805 53.080 155.850 ;
        RECT 54.650 155.805 54.940 155.850 ;
        RECT 55.190 155.850 62.765 155.990 ;
        RECT 67.150 155.990 67.290 156.145 ;
        RECT 69.360 156.130 69.680 156.190 ;
        RECT 70.755 156.145 71.045 156.190 ;
        RECT 73.515 156.145 73.805 156.190 ;
        RECT 69.450 155.990 69.590 156.130 ;
        RECT 67.150 155.850 69.590 155.990 ;
        RECT 71.200 155.990 71.520 156.050 ;
        RECT 74.050 155.990 74.190 156.530 ;
        RECT 74.880 156.470 75.200 156.530 ;
        RECT 79.495 156.670 79.785 156.715 ;
        RECT 82.700 156.670 83.020 156.730 ;
        RECT 79.495 156.530 83.020 156.670 ;
        RECT 79.495 156.485 79.785 156.530 ;
        RECT 82.700 156.470 83.020 156.530 ;
        RECT 83.635 156.670 83.925 156.715 ;
        RECT 85.000 156.670 85.320 156.730 ;
        RECT 83.635 156.530 85.320 156.670 ;
        RECT 83.635 156.485 83.925 156.530 ;
        RECT 85.000 156.470 85.320 156.530 ;
        RECT 87.300 156.670 87.620 156.730 ;
        RECT 88.695 156.670 88.985 156.715 ;
        RECT 90.520 156.670 90.840 156.730 ;
        RECT 87.300 156.530 88.985 156.670 ;
        RECT 87.300 156.470 87.620 156.530 ;
        RECT 88.695 156.485 88.985 156.530 ;
        RECT 89.690 156.530 90.840 156.670 ;
        RECT 77.655 156.330 77.945 156.375 ;
        RECT 79.940 156.330 80.260 156.390 ;
        RECT 77.655 156.190 80.260 156.330 ;
        RECT 77.655 156.145 77.945 156.190 ;
        RECT 79.940 156.130 80.260 156.190 ;
        RECT 82.255 156.330 82.545 156.375 ;
        RECT 84.095 156.330 84.385 156.375 ;
        RECT 82.255 156.190 84.385 156.330 ;
        RECT 82.255 156.145 82.545 156.190 ;
        RECT 84.095 156.145 84.385 156.190 ;
        RECT 88.235 156.330 88.525 156.375 ;
        RECT 89.140 156.330 89.460 156.390 ;
        RECT 89.690 156.375 89.830 156.530 ;
        RECT 90.520 156.470 90.840 156.530 ;
        RECT 91.440 156.470 91.760 156.730 ;
        RECT 88.235 156.190 89.460 156.330 ;
        RECT 88.235 156.145 88.525 156.190 ;
        RECT 89.140 156.130 89.460 156.190 ;
        RECT 89.615 156.145 89.905 156.375 ;
        RECT 92.360 156.130 92.680 156.390 ;
        RECT 92.910 156.330 93.050 156.870 ;
        RECT 93.280 157.010 93.600 157.070 ;
        RECT 95.580 157.010 95.900 157.070 ;
        RECT 96.500 157.010 96.820 157.070 ;
        RECT 103.400 157.010 103.720 157.070 ;
        RECT 93.280 156.870 95.900 157.010 ;
        RECT 93.280 156.810 93.600 156.870 ;
        RECT 95.580 156.810 95.900 156.870 ;
        RECT 96.130 156.870 103.720 157.010 ;
        RECT 93.740 156.670 94.060 156.730 ;
        RECT 96.130 156.670 96.270 156.870 ;
        RECT 96.500 156.810 96.820 156.870 ;
        RECT 103.400 156.810 103.720 156.870 ;
        RECT 106.635 157.010 106.925 157.055 ;
        RECT 106.635 156.870 111.910 157.010 ;
        RECT 106.635 156.825 106.925 156.870 ;
        RECT 93.740 156.530 96.270 156.670 ;
        RECT 97.510 156.530 101.330 156.670 ;
        RECT 93.740 156.470 94.060 156.530 ;
        RECT 94.905 156.330 95.195 156.375 ;
        RECT 92.910 156.190 95.195 156.330 ;
        RECT 94.905 156.145 95.195 156.190 ;
        RECT 95.595 156.145 95.885 156.375 ;
        RECT 96.055 156.330 96.345 156.375 ;
        RECT 96.500 156.330 96.820 156.390 ;
        RECT 96.055 156.190 96.820 156.330 ;
        RECT 96.055 156.145 96.345 156.190 ;
        RECT 71.200 155.850 74.190 155.990 ;
        RECT 90.995 155.990 91.285 156.035 ;
        RECT 93.755 155.990 94.045 156.035 ;
        RECT 90.995 155.850 94.045 155.990 ;
        RECT 95.670 155.990 95.810 156.145 ;
        RECT 96.500 156.130 96.820 156.190 ;
        RECT 97.035 156.315 97.325 156.375 ;
        RECT 97.510 156.315 97.650 156.530 ;
        RECT 97.035 156.175 97.650 156.315 ;
        RECT 97.035 156.145 97.325 156.175 ;
        RECT 99.260 156.130 99.580 156.390 ;
        RECT 99.720 156.130 100.040 156.390 ;
        RECT 101.190 156.375 101.330 156.530 ;
        RECT 103.860 156.470 104.180 156.730 ;
        RECT 105.240 156.670 105.560 156.730 ;
        RECT 107.095 156.670 107.385 156.715 ;
        RECT 105.240 156.530 107.385 156.670 ;
        RECT 105.240 156.470 105.560 156.530 ;
        RECT 107.095 156.485 107.385 156.530 ;
        RECT 100.195 156.145 100.485 156.375 ;
        RECT 101.115 156.330 101.405 156.375 ;
        RECT 101.560 156.330 101.880 156.390 ;
        RECT 101.115 156.190 101.880 156.330 ;
        RECT 101.115 156.145 101.405 156.190 ;
        RECT 99.810 155.990 99.950 156.130 ;
        RECT 95.670 155.850 99.950 155.990 ;
        RECT 100.270 155.990 100.410 156.145 ;
        RECT 101.560 156.130 101.880 156.190 ;
        RECT 104.795 156.330 105.085 156.375 ;
        RECT 105.700 156.330 106.020 156.390 ;
        RECT 111.770 156.375 111.910 156.870 ;
        RECT 104.795 156.190 106.020 156.330 ;
        RECT 104.795 156.145 105.085 156.190 ;
        RECT 104.870 155.990 105.010 156.145 ;
        RECT 105.700 156.130 106.020 156.190 ;
        RECT 111.695 156.145 111.985 156.375 ;
        RECT 100.270 155.850 105.010 155.990 ;
        RECT 55.190 155.650 55.330 155.850 ;
        RECT 62.475 155.805 62.765 155.850 ;
        RECT 71.200 155.790 71.520 155.850 ;
        RECT 90.995 155.805 91.285 155.850 ;
        RECT 93.755 155.805 94.045 155.850 ;
        RECT 52.430 155.510 55.330 155.650 ;
        RECT 56.495 155.650 56.785 155.695 ;
        RECT 56.940 155.650 57.260 155.710 ;
        RECT 56.495 155.510 57.260 155.650 ;
        RECT 45.900 155.450 46.220 155.510 ;
        RECT 46.605 155.465 46.895 155.510 ;
        RECT 56.495 155.465 56.785 155.510 ;
        RECT 56.940 155.450 57.260 155.510 ;
        RECT 60.635 155.650 60.925 155.695 ;
        RECT 64.760 155.650 65.080 155.710 ;
        RECT 60.635 155.510 65.080 155.650 ;
        RECT 60.635 155.465 60.925 155.510 ;
        RECT 64.760 155.450 65.080 155.510 ;
        RECT 65.680 155.650 66.000 155.710 ;
        RECT 66.155 155.650 66.445 155.695 ;
        RECT 65.680 155.510 66.445 155.650 ;
        RECT 65.680 155.450 66.000 155.510 ;
        RECT 66.155 155.465 66.445 155.510 ;
        RECT 67.980 155.450 68.300 155.710 ;
        RECT 69.820 155.450 70.140 155.710 ;
        RECT 72.120 155.650 72.440 155.710 ;
        RECT 72.595 155.650 72.885 155.695 ;
        RECT 72.120 155.510 72.885 155.650 ;
        RECT 72.120 155.450 72.440 155.510 ;
        RECT 72.595 155.465 72.885 155.510 ;
        RECT 78.100 155.450 78.420 155.710 ;
        RECT 83.620 155.650 83.940 155.710 ;
        RECT 84.555 155.650 84.845 155.695 ;
        RECT 83.620 155.510 84.845 155.650 ;
        RECT 83.620 155.450 83.940 155.510 ;
        RECT 84.555 155.465 84.845 155.510 ;
        RECT 86.395 155.650 86.685 155.695 ;
        RECT 87.760 155.650 88.080 155.710 ;
        RECT 86.395 155.510 88.080 155.650 ;
        RECT 86.395 155.465 86.685 155.510 ;
        RECT 87.760 155.450 88.080 155.510 ;
        RECT 90.520 155.450 90.840 155.710 ;
        RECT 91.900 155.650 92.220 155.710 ;
        RECT 93.295 155.650 93.585 155.695 ;
        RECT 91.900 155.510 93.585 155.650 ;
        RECT 91.900 155.450 92.220 155.510 ;
        RECT 93.295 155.465 93.585 155.510 ;
        RECT 95.120 155.650 95.440 155.710 ;
        RECT 97.895 155.650 98.185 155.695 ;
        RECT 95.120 155.510 98.185 155.650 ;
        RECT 95.120 155.450 95.440 155.510 ;
        RECT 97.895 155.465 98.185 155.510 ;
        RECT 104.320 155.450 104.640 155.710 ;
        RECT 109.840 155.650 110.160 155.710 ;
        RECT 110.775 155.650 111.065 155.695 ;
        RECT 109.840 155.510 111.065 155.650 ;
        RECT 109.840 155.450 110.160 155.510 ;
        RECT 110.775 155.465 111.065 155.510 ;
        RECT 22.830 154.830 113.450 155.310 ;
        RECT 35.320 154.430 35.640 154.690 ;
        RECT 40.840 154.630 41.160 154.690 ;
        RECT 37.710 154.490 41.160 154.630 ;
        RECT 27.500 154.290 27.820 154.350 ;
        RECT 37.710 154.335 37.850 154.490 ;
        RECT 40.840 154.430 41.160 154.490 ;
        RECT 45.900 154.430 46.220 154.690 ;
        RECT 73.515 154.630 73.805 154.675 ;
        RECT 85.000 154.630 85.320 154.690 ;
        RECT 46.450 154.490 64.070 154.630 ;
        RECT 27.500 154.150 36.010 154.290 ;
        RECT 27.500 154.090 27.820 154.150 ;
        RECT 26.120 153.950 26.440 154.010 ;
        RECT 26.595 153.950 26.885 153.995 ;
        RECT 26.120 153.810 26.885 153.950 ;
        RECT 26.120 153.750 26.440 153.810 ;
        RECT 26.595 153.765 26.885 153.810 ;
        RECT 29.800 153.750 30.120 154.010 ;
        RECT 28.895 153.425 29.185 153.655 ;
        RECT 28.970 153.270 29.110 153.425 ;
        RECT 29.340 153.410 29.660 153.670 ;
        RECT 35.870 153.270 36.010 154.150 ;
        RECT 37.635 154.105 37.925 154.335 ;
        RECT 38.095 154.105 38.385 154.335 ;
        RECT 38.540 154.290 38.860 154.350 ;
        RECT 41.775 154.290 42.065 154.335 ;
        RECT 38.540 154.150 42.065 154.290 ;
        RECT 36.255 153.950 36.545 153.995 ;
        RECT 38.170 153.950 38.310 154.105 ;
        RECT 38.540 154.090 38.860 154.150 ;
        RECT 41.775 154.105 42.065 154.150 ;
        RECT 42.680 154.290 43.000 154.350 ;
        RECT 46.450 154.290 46.590 154.490 ;
        RECT 42.680 154.150 46.590 154.290 ;
        RECT 48.200 154.290 48.520 154.350 ;
        RECT 50.040 154.290 50.360 154.350 ;
        RECT 56.020 154.290 56.340 154.350 ;
        RECT 56.940 154.335 57.260 154.350 ;
        RECT 48.200 154.150 50.360 154.290 ;
        RECT 42.680 154.090 43.000 154.150 ;
        RECT 36.255 153.810 38.310 153.950 ;
        RECT 36.255 153.765 36.545 153.810 ;
        RECT 39.460 153.750 39.780 154.010 ;
        RECT 39.935 153.765 40.225 153.995 ;
        RECT 40.395 153.765 40.685 153.995 ;
        RECT 36.700 153.410 37.020 153.670 ;
        RECT 39.000 153.610 39.320 153.670 ;
        RECT 40.010 153.610 40.150 153.765 ;
        RECT 39.000 153.470 40.150 153.610 ;
        RECT 39.000 153.410 39.320 153.470 ;
        RECT 40.470 153.270 40.610 153.765 ;
        RECT 41.300 153.750 41.620 154.010 ;
        RECT 43.230 153.995 43.370 154.150 ;
        RECT 48.200 154.090 48.520 154.150 ;
        RECT 50.040 154.090 50.360 154.150 ;
        RECT 50.590 154.150 56.340 154.290 ;
        RECT 43.155 153.765 43.445 153.995 ;
        RECT 46.360 153.750 46.680 154.010 ;
        RECT 46.820 153.950 47.140 154.010 ;
        RECT 50.590 153.995 50.730 154.150 ;
        RECT 56.020 154.090 56.340 154.150 ;
        RECT 56.890 154.290 57.260 154.335 ;
        RECT 60.150 154.290 60.440 154.335 ;
        RECT 56.890 154.150 60.440 154.290 ;
        RECT 56.890 154.105 57.260 154.150 ;
        RECT 60.150 154.105 60.440 154.150 ;
        RECT 61.070 154.290 61.360 154.335 ;
        RECT 62.930 154.290 63.220 154.335 ;
        RECT 61.070 154.150 63.220 154.290 ;
        RECT 63.930 154.290 64.070 154.490 ;
        RECT 65.770 154.490 68.670 154.630 ;
        RECT 65.770 154.335 65.910 154.490 ;
        RECT 63.930 154.150 65.450 154.290 ;
        RECT 61.070 154.105 61.360 154.150 ;
        RECT 62.930 154.105 63.220 154.150 ;
        RECT 56.940 154.090 57.260 154.105 ;
        RECT 50.515 153.950 50.805 153.995 ;
        RECT 46.820 153.810 50.805 153.950 ;
        RECT 46.820 153.750 47.140 153.810 ;
        RECT 50.515 153.765 50.805 153.810 ;
        RECT 50.960 153.750 51.280 154.010 ;
        RECT 51.435 153.950 51.725 153.995 ;
        RECT 52.355 153.950 52.645 153.995 ;
        RECT 52.800 153.950 53.120 154.010 ;
        RECT 51.435 153.810 52.110 153.950 ;
        RECT 51.435 153.765 51.725 153.810 ;
        RECT 42.220 153.410 42.540 153.670 ;
        RECT 45.455 153.610 45.745 153.655 ;
        RECT 45.455 153.470 50.730 153.610 ;
        RECT 45.455 153.425 45.745 153.470 ;
        RECT 50.590 153.330 50.730 153.470 ;
        RECT 28.970 153.130 35.550 153.270 ;
        RECT 35.870 153.130 40.610 153.270 ;
        RECT 27.040 152.730 27.360 152.990 ;
        RECT 31.655 152.930 31.945 152.975 ;
        RECT 32.560 152.930 32.880 152.990 ;
        RECT 31.655 152.790 32.880 152.930 ;
        RECT 35.410 152.930 35.550 153.130 ;
        RECT 44.060 153.070 44.380 153.330 ;
        RECT 48.200 153.070 48.520 153.330 ;
        RECT 50.500 153.070 50.820 153.330 ;
        RECT 51.970 153.270 52.110 153.810 ;
        RECT 52.355 153.810 53.120 153.950 ;
        RECT 52.355 153.765 52.645 153.810 ;
        RECT 52.800 153.750 53.120 153.810 ;
        RECT 53.260 153.750 53.580 154.010 ;
        RECT 58.750 153.950 59.040 153.995 ;
        RECT 61.070 153.950 61.285 154.105 ;
        RECT 65.310 153.995 65.450 154.150 ;
        RECT 65.695 154.105 65.985 154.335 ;
        RECT 67.535 154.290 67.825 154.335 ;
        RECT 66.230 154.150 67.825 154.290 ;
        RECT 66.230 154.010 66.370 154.150 ;
        RECT 67.535 154.105 67.825 154.150 ;
        RECT 68.530 154.010 68.670 154.490 ;
        RECT 73.515 154.490 85.320 154.630 ;
        RECT 73.515 154.445 73.805 154.490 ;
        RECT 85.000 154.430 85.320 154.490 ;
        RECT 88.695 154.630 88.985 154.675 ;
        RECT 90.060 154.630 90.380 154.690 ;
        RECT 88.695 154.490 90.380 154.630 ;
        RECT 88.695 154.445 88.985 154.490 ;
        RECT 90.060 154.430 90.380 154.490 ;
        RECT 91.900 154.630 92.220 154.690 ;
        RECT 106.160 154.630 106.480 154.690 ;
        RECT 91.900 154.490 106.480 154.630 ;
        RECT 91.900 154.430 92.220 154.490 ;
        RECT 106.160 154.430 106.480 154.490 ;
        RECT 69.375 154.290 69.665 154.335 ;
        RECT 72.120 154.290 72.440 154.350 ;
        RECT 69.375 154.150 72.440 154.290 ;
        RECT 69.375 154.105 69.665 154.150 ;
        RECT 72.120 154.090 72.440 154.150 ;
        RECT 78.100 154.290 78.420 154.350 ;
        RECT 79.430 154.290 79.720 154.335 ;
        RECT 82.690 154.290 82.980 154.335 ;
        RECT 78.100 154.150 82.980 154.290 ;
        RECT 78.100 154.090 78.420 154.150 ;
        RECT 79.430 154.105 79.720 154.150 ;
        RECT 82.690 154.105 82.980 154.150 ;
        RECT 83.610 154.290 83.900 154.335 ;
        RECT 85.470 154.290 85.760 154.335 ;
        RECT 94.660 154.290 94.980 154.350 ;
        RECT 83.610 154.150 85.760 154.290 ;
        RECT 83.610 154.105 83.900 154.150 ;
        RECT 85.470 154.105 85.760 154.150 ;
        RECT 93.830 154.150 94.980 154.290 ;
        RECT 58.750 153.810 61.285 153.950 ;
        RECT 62.015 153.950 62.305 153.995 ;
        RECT 62.015 153.810 64.530 153.950 ;
        RECT 58.750 153.765 59.040 153.810 ;
        RECT 62.015 153.765 62.305 153.810 ;
        RECT 55.560 153.610 55.880 153.670 ;
        RECT 59.240 153.610 59.560 153.670 ;
        RECT 63.855 153.610 64.145 153.655 ;
        RECT 55.560 153.470 64.145 153.610 ;
        RECT 55.560 153.410 55.880 153.470 ;
        RECT 59.240 153.410 59.560 153.470 ;
        RECT 63.855 153.425 64.145 153.470 ;
        RECT 54.885 153.270 55.175 153.315 ;
        RECT 57.400 153.270 57.720 153.330 ;
        RECT 64.390 153.315 64.530 153.810 ;
        RECT 65.235 153.765 65.525 153.995 ;
        RECT 66.140 153.750 66.460 154.010 ;
        RECT 67.075 153.765 67.365 153.995 ;
        RECT 68.440 153.950 68.760 154.010 ;
        RECT 73.960 153.950 74.280 154.010 ;
        RECT 68.440 153.810 74.280 153.950 ;
        RECT 64.760 153.610 65.080 153.670 ;
        RECT 67.150 153.610 67.290 153.765 ;
        RECT 68.440 153.750 68.760 153.810 ;
        RECT 73.960 153.750 74.280 153.810 ;
        RECT 81.290 153.950 81.580 153.995 ;
        RECT 83.610 153.950 83.825 154.105 ;
        RECT 81.290 153.810 83.825 153.950 ;
        RECT 81.290 153.765 81.580 153.810 ;
        RECT 84.540 153.750 84.860 154.010 ;
        RECT 87.760 153.750 88.080 154.010 ;
        RECT 93.830 153.995 93.970 154.150 ;
        RECT 94.660 154.090 94.980 154.150 ;
        RECT 95.120 154.090 95.440 154.350 ;
        RECT 100.640 154.290 100.960 154.350 ;
        RECT 95.670 154.150 100.960 154.290 ;
        RECT 93.755 153.765 94.045 153.995 ;
        RECT 94.215 153.950 94.505 153.995 ;
        RECT 95.670 153.950 95.810 154.150 ;
        RECT 100.640 154.090 100.960 154.150 ;
        RECT 101.575 154.290 101.865 154.335 ;
        RECT 104.730 154.290 105.020 154.335 ;
        RECT 107.990 154.290 108.280 154.335 ;
        RECT 101.575 154.150 108.280 154.290 ;
        RECT 101.575 154.105 101.865 154.150 ;
        RECT 104.730 154.105 105.020 154.150 ;
        RECT 107.990 154.105 108.280 154.150 ;
        RECT 108.910 154.290 109.200 154.335 ;
        RECT 110.770 154.290 111.060 154.335 ;
        RECT 108.910 154.150 111.060 154.290 ;
        RECT 108.910 154.105 109.200 154.150 ;
        RECT 110.770 154.105 111.060 154.150 ;
        RECT 94.215 153.810 95.810 153.950 ;
        RECT 96.040 153.950 96.360 154.010 ;
        RECT 96.515 153.950 96.805 153.995 ;
        RECT 96.040 153.810 96.805 153.950 ;
        RECT 94.215 153.765 94.505 153.810 ;
        RECT 96.040 153.750 96.360 153.810 ;
        RECT 96.515 153.765 96.805 153.810 ;
        RECT 97.880 153.750 98.200 154.010 ;
        RECT 101.100 153.750 101.420 154.010 ;
        RECT 106.590 153.950 106.880 153.995 ;
        RECT 108.910 153.950 109.125 154.105 ;
        RECT 106.590 153.810 109.125 153.950 ;
        RECT 106.590 153.765 106.880 153.810 ;
        RECT 109.840 153.750 110.160 154.010 ;
        RECT 111.220 153.950 111.540 154.010 ;
        RECT 111.695 153.950 111.985 153.995 ;
        RECT 111.220 153.810 111.985 153.950 ;
        RECT 111.220 153.750 111.540 153.810 ;
        RECT 111.695 153.765 111.985 153.810 ;
        RECT 64.760 153.470 67.290 153.610 ;
        RECT 64.760 153.410 65.080 153.470 ;
        RECT 86.380 153.410 86.700 153.670 ;
        RECT 97.435 153.610 97.725 153.655 ;
        RECT 98.340 153.610 98.660 153.670 ;
        RECT 97.435 153.470 98.660 153.610 ;
        RECT 97.435 153.425 97.725 153.470 ;
        RECT 98.340 153.410 98.660 153.470 ;
        RECT 51.970 153.130 57.720 153.270 ;
        RECT 54.885 153.085 55.175 153.130 ;
        RECT 57.400 153.070 57.720 153.130 ;
        RECT 58.750 153.270 59.040 153.315 ;
        RECT 61.530 153.270 61.820 153.315 ;
        RECT 63.390 153.270 63.680 153.315 ;
        RECT 58.750 153.130 63.680 153.270 ;
        RECT 58.750 153.085 59.040 153.130 ;
        RECT 61.530 153.085 61.820 153.130 ;
        RECT 63.390 153.085 63.680 153.130 ;
        RECT 64.315 153.085 64.605 153.315 ;
        RECT 67.520 153.270 67.840 153.330 ;
        RECT 81.290 153.270 81.580 153.315 ;
        RECT 84.070 153.270 84.360 153.315 ;
        RECT 85.930 153.270 86.220 153.315 ;
        RECT 94.200 153.270 94.520 153.330 ;
        RECT 67.520 153.130 81.090 153.270 ;
        RECT 67.520 153.070 67.840 153.130 ;
        RECT 36.700 152.930 37.020 152.990 ;
        RECT 35.410 152.790 37.020 152.930 ;
        RECT 31.655 152.745 31.945 152.790 ;
        RECT 32.560 152.730 32.880 152.790 ;
        RECT 36.700 152.730 37.020 152.790 ;
        RECT 37.620 152.730 37.940 152.990 ;
        RECT 42.680 152.730 43.000 152.990 ;
        RECT 43.140 152.930 43.460 152.990 ;
        RECT 49.135 152.930 49.425 152.975 ;
        RECT 43.140 152.790 49.425 152.930 ;
        RECT 43.140 152.730 43.460 152.790 ;
        RECT 49.135 152.745 49.425 152.790 ;
        RECT 54.195 152.930 54.485 152.975 ;
        RECT 56.020 152.930 56.340 152.990 ;
        RECT 54.195 152.790 56.340 152.930 ;
        RECT 54.195 152.745 54.485 152.790 ;
        RECT 56.020 152.730 56.340 152.790 ;
        RECT 77.425 152.930 77.715 152.975 ;
        RECT 79.480 152.930 79.800 152.990 ;
        RECT 77.425 152.790 79.800 152.930 ;
        RECT 80.950 152.930 81.090 153.130 ;
        RECT 81.290 153.130 86.220 153.270 ;
        RECT 81.290 153.085 81.580 153.130 ;
        RECT 84.070 153.085 84.360 153.130 ;
        RECT 85.930 153.085 86.220 153.130 ;
        RECT 91.070 153.130 94.520 153.270 ;
        RECT 89.600 152.930 89.920 152.990 ;
        RECT 91.070 152.930 91.210 153.130 ;
        RECT 94.200 153.070 94.520 153.130 ;
        RECT 106.590 153.270 106.880 153.315 ;
        RECT 109.370 153.270 109.660 153.315 ;
        RECT 111.230 153.270 111.520 153.315 ;
        RECT 106.590 153.130 111.520 153.270 ;
        RECT 106.590 153.085 106.880 153.130 ;
        RECT 109.370 153.085 109.660 153.130 ;
        RECT 111.230 153.085 111.520 153.130 ;
        RECT 80.950 152.790 91.210 152.930 ;
        RECT 91.440 152.930 91.760 152.990 ;
        RECT 92.835 152.930 93.125 152.975 ;
        RECT 91.440 152.790 93.125 152.930 ;
        RECT 77.425 152.745 77.715 152.790 ;
        RECT 79.480 152.730 79.800 152.790 ;
        RECT 89.600 152.730 89.920 152.790 ;
        RECT 91.440 152.730 91.760 152.790 ;
        RECT 92.835 152.745 93.125 152.790 ;
        RECT 95.120 152.730 95.440 152.990 ;
        RECT 95.580 152.730 95.900 152.990 ;
        RECT 97.895 152.930 98.185 152.975 ;
        RECT 98.340 152.930 98.660 152.990 ;
        RECT 97.895 152.790 98.660 152.930 ;
        RECT 97.895 152.745 98.185 152.790 ;
        RECT 98.340 152.730 98.660 152.790 ;
        RECT 102.725 152.930 103.015 152.975 ;
        RECT 104.320 152.930 104.640 152.990 ;
        RECT 102.725 152.790 104.640 152.930 ;
        RECT 102.725 152.745 103.015 152.790 ;
        RECT 104.320 152.730 104.640 152.790 ;
        RECT 22.830 152.110 113.450 152.590 ;
        RECT 30.260 151.910 30.580 151.970 ;
        RECT 30.260 151.770 36.010 151.910 ;
        RECT 30.260 151.710 30.580 151.770 ;
        RECT 28.850 151.570 29.140 151.615 ;
        RECT 31.630 151.570 31.920 151.615 ;
        RECT 33.490 151.570 33.780 151.615 ;
        RECT 28.850 151.430 33.780 151.570 ;
        RECT 28.850 151.385 29.140 151.430 ;
        RECT 31.630 151.385 31.920 151.430 ;
        RECT 33.490 151.385 33.780 151.430 ;
        RECT 24.985 151.230 25.275 151.275 ;
        RECT 29.340 151.230 29.660 151.290 ;
        RECT 24.985 151.090 29.660 151.230 ;
        RECT 24.985 151.045 25.275 151.090 ;
        RECT 29.340 151.030 29.660 151.090 ;
        RECT 32.560 151.230 32.880 151.290 ;
        RECT 35.870 151.230 36.010 151.770 ;
        RECT 38.540 151.710 38.860 151.970 ;
        RECT 40.840 151.710 41.160 151.970 ;
        RECT 41.300 151.710 41.620 151.970 ;
        RECT 44.520 151.710 44.840 151.970 ;
        RECT 50.960 151.910 51.280 151.970 ;
        RECT 47.370 151.770 51.280 151.910 ;
        RECT 40.930 151.570 41.070 151.710 ;
        RECT 41.775 151.570 42.065 151.615 ;
        RECT 40.930 151.430 42.065 151.570 ;
        RECT 41.775 151.385 42.065 151.430 ;
        RECT 43.600 151.570 43.920 151.630 ;
        RECT 44.610 151.570 44.750 151.710 ;
        RECT 47.370 151.570 47.510 151.770 ;
        RECT 50.960 151.710 51.280 151.770 ;
        RECT 53.260 151.710 53.580 151.970 ;
        RECT 61.540 151.910 61.860 151.970 ;
        RECT 65.680 151.910 66.000 151.970 ;
        RECT 61.540 151.770 70.510 151.910 ;
        RECT 61.540 151.710 61.860 151.770 ;
        RECT 65.680 151.710 66.000 151.770 ;
        RECT 43.600 151.430 47.510 151.570 ;
        RECT 43.600 151.370 43.920 151.430 ;
        RECT 37.635 151.230 37.925 151.275 ;
        RECT 32.560 151.090 35.550 151.230 ;
        RECT 35.870 151.090 37.925 151.230 ;
        RECT 32.560 151.030 32.880 151.090 ;
        RECT 28.850 150.890 29.140 150.935 ;
        RECT 28.850 150.750 31.385 150.890 ;
        RECT 28.850 150.705 29.140 150.750 ;
        RECT 27.040 150.595 27.360 150.610 ;
        RECT 31.170 150.595 31.385 150.750 ;
        RECT 32.100 150.690 32.420 150.950 ;
        RECT 33.955 150.890 34.245 150.935 ;
        RECT 34.860 150.890 35.180 150.950 ;
        RECT 35.410 150.935 35.550 151.090 ;
        RECT 37.635 151.045 37.925 151.090 ;
        RECT 40.380 151.030 40.700 151.290 ;
        RECT 43.230 151.090 47.050 151.230 ;
        RECT 33.955 150.750 35.180 150.890 ;
        RECT 33.955 150.705 34.245 150.750 ;
        RECT 34.860 150.690 35.180 150.750 ;
        RECT 35.335 150.705 35.625 150.935 ;
        RECT 35.780 150.890 36.100 150.950 ;
        RECT 37.175 150.890 37.465 150.935 ;
        RECT 35.780 150.750 37.465 150.890 ;
        RECT 35.780 150.690 36.100 150.750 ;
        RECT 37.175 150.705 37.465 150.750 ;
        RECT 39.920 150.690 40.240 150.950 ;
        RECT 43.230 150.935 43.370 151.090 ;
        RECT 46.910 150.950 47.050 151.090 ;
        RECT 43.155 150.705 43.445 150.935 ;
        RECT 43.600 150.690 43.920 150.950 ;
        RECT 44.060 150.690 44.380 150.950 ;
        RECT 44.995 150.890 45.285 150.935 ;
        RECT 44.995 150.750 46.590 150.890 ;
        RECT 44.995 150.705 45.285 150.750 ;
        RECT 26.990 150.550 27.360 150.595 ;
        RECT 30.250 150.550 30.540 150.595 ;
        RECT 26.990 150.410 30.540 150.550 ;
        RECT 26.990 150.365 27.360 150.410 ;
        RECT 30.250 150.365 30.540 150.410 ;
        RECT 31.170 150.550 31.460 150.595 ;
        RECT 33.030 150.550 33.320 150.595 ;
        RECT 31.170 150.410 33.320 150.550 ;
        RECT 31.170 150.365 31.460 150.410 ;
        RECT 33.030 150.365 33.320 150.410 ;
        RECT 38.555 150.550 38.845 150.595 ;
        RECT 41.315 150.550 41.605 150.595 ;
        RECT 45.455 150.550 45.745 150.595 ;
        RECT 38.555 150.410 41.070 150.550 ;
        RECT 38.555 150.365 38.845 150.410 ;
        RECT 27.040 150.350 27.360 150.365 ;
        RECT 31.640 150.210 31.960 150.270 ;
        RECT 34.415 150.210 34.705 150.255 ;
        RECT 31.640 150.070 34.705 150.210 ;
        RECT 31.640 150.010 31.960 150.070 ;
        RECT 34.415 150.025 34.705 150.070 ;
        RECT 36.240 150.010 36.560 150.270 ;
        RECT 39.000 150.010 39.320 150.270 ;
        RECT 40.930 150.210 41.070 150.410 ;
        RECT 41.315 150.410 45.745 150.550 ;
        RECT 41.315 150.365 41.605 150.410 ;
        RECT 45.455 150.365 45.745 150.410 ;
        RECT 43.140 150.210 43.460 150.270 ;
        RECT 40.930 150.070 43.460 150.210 ;
        RECT 46.450 150.210 46.590 150.750 ;
        RECT 46.820 150.690 47.140 150.950 ;
        RECT 47.370 150.935 47.510 151.430 ;
        RECT 48.200 151.570 48.520 151.630 ;
        RECT 54.180 151.570 54.500 151.630 ;
        RECT 48.200 151.430 54.500 151.570 ;
        RECT 48.200 151.370 48.520 151.430 ;
        RECT 54.180 151.370 54.500 151.430 ;
        RECT 61.095 151.570 61.385 151.615 ;
        RECT 64.300 151.570 64.620 151.630 ;
        RECT 61.095 151.430 64.620 151.570 ;
        RECT 61.095 151.385 61.385 151.430 ;
        RECT 64.300 151.370 64.620 151.430 ;
        RECT 64.875 151.570 65.165 151.615 ;
        RECT 67.995 151.570 68.285 151.615 ;
        RECT 69.885 151.570 70.175 151.615 ;
        RECT 64.875 151.430 70.175 151.570 ;
        RECT 70.370 151.570 70.510 151.770 ;
        RECT 73.500 151.710 73.820 151.970 ;
        RECT 82.240 151.710 82.560 151.970 ;
        RECT 96.975 151.910 97.265 151.955 ;
        RECT 97.880 151.910 98.200 151.970 ;
        RECT 96.975 151.770 98.200 151.910 ;
        RECT 96.975 151.725 97.265 151.770 ;
        RECT 97.880 151.710 98.200 151.770 ;
        RECT 73.960 151.570 74.280 151.630 ;
        RECT 101.560 151.570 101.880 151.630 ;
        RECT 70.370 151.430 76.950 151.570 ;
        RECT 64.875 151.385 65.165 151.430 ;
        RECT 67.995 151.385 68.285 151.430 ;
        RECT 69.885 151.385 70.175 151.430 ;
        RECT 73.960 151.370 74.280 151.430 ;
        RECT 50.500 151.030 50.820 151.290 ;
        RECT 58.335 151.230 58.625 151.275 ;
        RECT 62.015 151.230 62.305 151.275 ;
        RECT 56.570 151.090 62.305 151.230 ;
        RECT 47.295 150.705 47.585 150.935 ;
        RECT 47.755 150.705 48.045 150.935 ;
        RECT 48.660 150.890 48.980 150.950 ;
        RECT 51.880 150.890 52.200 150.950 ;
        RECT 56.570 150.935 56.710 151.090 ;
        RECT 58.335 151.045 58.625 151.090 ;
        RECT 62.015 151.045 62.305 151.090 ;
        RECT 73.055 151.230 73.345 151.275 ;
        RECT 74.420 151.230 74.740 151.290 ;
        RECT 73.055 151.090 74.740 151.230 ;
        RECT 73.055 151.045 73.345 151.090 ;
        RECT 74.420 151.030 74.740 151.090 ;
        RECT 48.660 150.750 52.200 150.890 ;
        RECT 47.830 150.550 47.970 150.705 ;
        RECT 48.660 150.690 48.980 150.750 ;
        RECT 51.880 150.690 52.200 150.750 ;
        RECT 55.575 150.705 55.865 150.935 ;
        RECT 56.035 150.705 56.325 150.935 ;
        RECT 56.495 150.705 56.785 150.935 ;
        RECT 57.415 150.890 57.705 150.935 ;
        RECT 61.540 150.890 61.860 150.950 ;
        RECT 57.415 150.750 61.860 150.890 ;
        RECT 57.415 150.705 57.705 150.750 ;
        RECT 51.435 150.550 51.725 150.595 ;
        RECT 52.340 150.550 52.660 150.610 ;
        RECT 47.830 150.410 52.660 150.550 ;
        RECT 51.435 150.365 51.725 150.410 ;
        RECT 52.340 150.350 52.660 150.410 ;
        RECT 48.660 150.210 48.980 150.270 ;
        RECT 46.450 150.070 48.980 150.210 ;
        RECT 43.140 150.010 43.460 150.070 ;
        RECT 48.660 150.010 48.980 150.070 ;
        RECT 49.580 150.210 49.900 150.270 ;
        RECT 50.975 150.210 51.265 150.255 ;
        RECT 49.580 150.070 51.265 150.210 ;
        RECT 49.580 150.010 49.900 150.070 ;
        RECT 50.975 150.025 51.265 150.070 ;
        RECT 51.880 150.210 52.200 150.270 ;
        RECT 54.195 150.210 54.485 150.255 ;
        RECT 51.880 150.070 54.485 150.210 ;
        RECT 55.650 150.210 55.790 150.705 ;
        RECT 56.110 150.550 56.250 150.705 ;
        RECT 61.540 150.690 61.860 150.750 ;
        RECT 60.620 150.550 60.940 150.610 ;
        RECT 56.110 150.410 60.940 150.550 ;
        RECT 60.620 150.350 60.940 150.410 ;
        RECT 61.080 150.550 61.400 150.610 ;
        RECT 63.795 150.595 64.085 150.910 ;
        RECT 64.875 150.890 65.165 150.935 ;
        RECT 68.455 150.890 68.745 150.935 ;
        RECT 70.290 150.890 70.580 150.935 ;
        RECT 64.875 150.750 70.580 150.890 ;
        RECT 64.875 150.705 65.165 150.750 ;
        RECT 68.455 150.705 68.745 150.750 ;
        RECT 70.290 150.705 70.580 150.750 ;
        RECT 70.740 150.690 71.060 150.950 ;
        RECT 72.135 150.890 72.425 150.935 ;
        RECT 72.580 150.890 72.900 150.950 ;
        RECT 75.355 150.890 75.645 150.935 ;
        RECT 72.135 150.750 72.900 150.890 ;
        RECT 72.135 150.705 72.425 150.750 ;
        RECT 72.580 150.690 72.900 150.750 ;
        RECT 73.130 150.750 75.645 150.890 ;
        RECT 63.495 150.550 64.085 150.595 ;
        RECT 66.735 150.550 67.385 150.595 ;
        RECT 61.080 150.410 67.385 150.550 ;
        RECT 61.080 150.350 61.400 150.410 ;
        RECT 63.495 150.365 63.785 150.410 ;
        RECT 66.735 150.365 67.385 150.410 ;
        RECT 69.360 150.350 69.680 150.610 ;
        RECT 73.130 150.550 73.270 150.750 ;
        RECT 75.355 150.705 75.645 150.750 ;
        RECT 75.800 150.690 76.120 150.950 ;
        RECT 76.275 150.705 76.565 150.935 ;
        RECT 76.810 150.890 76.950 151.430 ;
        RECT 79.110 151.430 85.690 151.570 ;
        RECT 79.110 151.275 79.250 151.430 ;
        RECT 85.550 151.290 85.690 151.430 ;
        RECT 93.830 151.430 101.880 151.570 ;
        RECT 79.035 151.045 79.325 151.275 ;
        RECT 79.495 151.230 79.785 151.275 ;
        RECT 79.495 151.090 84.310 151.230 ;
        RECT 79.495 151.045 79.785 151.090 ;
        RECT 77.195 150.890 77.485 150.935 ;
        RECT 76.810 150.750 77.485 150.890 ;
        RECT 77.195 150.705 77.485 150.750 ;
        RECT 78.560 150.890 78.880 150.950 ;
        RECT 79.570 150.890 79.710 151.045 ;
        RECT 84.170 150.935 84.310 151.090 ;
        RECT 85.460 151.030 85.780 151.290 ;
        RECT 78.560 150.750 79.710 150.890 ;
        RECT 70.600 150.410 73.270 150.550 ;
        RECT 73.515 150.550 73.805 150.595 ;
        RECT 73.975 150.550 74.265 150.595 ;
        RECT 73.515 150.410 74.265 150.550 ;
        RECT 76.350 150.550 76.490 150.705 ;
        RECT 78.560 150.690 78.880 150.750 ;
        RECT 84.095 150.705 84.385 150.935 ;
        RECT 91.900 150.890 92.220 150.950 ;
        RECT 93.830 150.935 93.970 151.430 ;
        RECT 101.560 151.370 101.880 151.430 ;
        RECT 94.200 151.230 94.520 151.290 ;
        RECT 97.435 151.230 97.725 151.275 ;
        RECT 97.880 151.230 98.200 151.290 ;
        RECT 100.180 151.230 100.500 151.290 ;
        RECT 101.650 151.230 101.790 151.370 ;
        RECT 94.200 151.090 97.190 151.230 ;
        RECT 94.200 151.030 94.520 151.090 ;
        RECT 95.210 150.935 95.350 151.090 ;
        RECT 93.755 150.890 94.045 150.935 ;
        RECT 91.900 150.750 94.045 150.890 ;
        RECT 91.900 150.690 92.220 150.750 ;
        RECT 93.755 150.705 94.045 150.750 ;
        RECT 94.675 150.705 94.965 150.935 ;
        RECT 95.135 150.705 95.425 150.935 ;
        RECT 95.595 150.705 95.885 150.935 ;
        RECT 97.050 150.890 97.190 151.090 ;
        RECT 97.435 151.090 98.200 151.230 ;
        RECT 97.435 151.045 97.725 151.090 ;
        RECT 97.880 151.030 98.200 151.090 ;
        RECT 98.430 151.090 100.500 151.230 ;
        RECT 98.430 150.890 98.570 151.090 ;
        RECT 97.050 150.750 98.570 150.890 ;
        RECT 79.480 150.550 79.800 150.610 ;
        RECT 83.620 150.550 83.940 150.610 ;
        RECT 84.555 150.550 84.845 150.595 ;
        RECT 76.350 150.410 84.845 150.550 ;
        RECT 57.400 150.210 57.720 150.270 ;
        RECT 55.650 150.070 57.720 150.210 ;
        RECT 51.880 150.010 52.200 150.070 ;
        RECT 54.195 150.025 54.485 150.070 ;
        RECT 57.400 150.010 57.720 150.070 ;
        RECT 67.980 150.210 68.300 150.270 ;
        RECT 70.600 150.210 70.740 150.410 ;
        RECT 73.515 150.365 73.805 150.410 ;
        RECT 73.975 150.365 74.265 150.410 ;
        RECT 79.480 150.350 79.800 150.410 ;
        RECT 83.620 150.350 83.940 150.410 ;
        RECT 84.555 150.365 84.845 150.410 ;
        RECT 67.980 150.070 70.740 150.210 ;
        RECT 67.980 150.010 68.300 150.070 ;
        RECT 71.200 150.010 71.520 150.270 ;
        RECT 79.955 150.210 80.245 150.255 ;
        RECT 80.860 150.210 81.180 150.270 ;
        RECT 79.955 150.070 81.180 150.210 ;
        RECT 79.955 150.025 80.245 150.070 ;
        RECT 80.860 150.010 81.180 150.070 ;
        RECT 81.795 150.210 82.085 150.255 ;
        RECT 87.760 150.210 88.080 150.270 ;
        RECT 81.795 150.070 88.080 150.210 ;
        RECT 94.750 150.210 94.890 150.705 ;
        RECT 95.670 150.550 95.810 150.705 ;
        RECT 98.800 150.690 99.120 150.950 ;
        RECT 99.350 150.935 99.490 151.090 ;
        RECT 100.180 151.030 100.500 151.090 ;
        RECT 100.730 151.090 101.790 151.230 ;
        RECT 100.730 150.935 100.870 151.090 ;
        RECT 103.860 151.030 104.180 151.290 ;
        RECT 99.275 150.705 99.565 150.935 ;
        RECT 99.735 150.705 100.025 150.935 ;
        RECT 100.655 150.705 100.945 150.935 ;
        RECT 101.100 150.890 101.420 150.950 ;
        RECT 101.575 150.890 101.865 150.935 ;
        RECT 101.100 150.750 101.865 150.890 ;
        RECT 96.040 150.550 96.360 150.610 ;
        RECT 98.890 150.550 99.030 150.690 ;
        RECT 95.670 150.410 99.030 150.550 ;
        RECT 99.810 150.550 99.950 150.705 ;
        RECT 101.100 150.690 101.420 150.750 ;
        RECT 101.575 150.705 101.865 150.750 ;
        RECT 102.020 150.890 102.340 150.950 ;
        RECT 104.320 150.890 104.640 150.950 ;
        RECT 104.795 150.890 105.085 150.935 ;
        RECT 108.015 150.890 108.305 150.935 ;
        RECT 102.020 150.750 105.085 150.890 ;
        RECT 102.020 150.690 102.340 150.750 ;
        RECT 104.320 150.690 104.640 150.750 ;
        RECT 104.795 150.705 105.085 150.750 ;
        RECT 106.710 150.750 108.305 150.890 ;
        RECT 99.810 150.410 104.090 150.550 ;
        RECT 96.040 150.350 96.360 150.410 ;
        RECT 103.950 150.270 104.090 150.410 ;
        RECT 101.560 150.210 101.880 150.270 ;
        RECT 94.750 150.070 101.880 150.210 ;
        RECT 81.795 150.025 82.085 150.070 ;
        RECT 87.760 150.010 88.080 150.070 ;
        RECT 101.560 150.010 101.880 150.070 ;
        RECT 102.020 150.010 102.340 150.270 ;
        RECT 103.860 150.210 104.180 150.270 ;
        RECT 106.710 150.255 106.850 150.750 ;
        RECT 108.015 150.705 108.305 150.750 ;
        RECT 104.335 150.210 104.625 150.255 ;
        RECT 103.860 150.070 104.625 150.210 ;
        RECT 103.860 150.010 104.180 150.070 ;
        RECT 104.335 150.025 104.625 150.070 ;
        RECT 106.635 150.025 106.925 150.255 ;
        RECT 108.935 150.210 109.225 150.255 ;
        RECT 109.840 150.210 110.160 150.270 ;
        RECT 108.935 150.070 110.160 150.210 ;
        RECT 108.935 150.025 109.225 150.070 ;
        RECT 109.840 150.010 110.160 150.070 ;
        RECT 22.830 149.390 113.450 149.870 ;
        RECT 29.340 149.190 29.660 149.250 ;
        RECT 35.795 149.190 36.085 149.235 ;
        RECT 39.920 149.190 40.240 149.250 ;
        RECT 29.340 149.050 40.240 149.190 ;
        RECT 29.340 148.990 29.660 149.050 ;
        RECT 35.795 149.005 36.085 149.050 ;
        RECT 39.920 148.990 40.240 149.050 ;
        RECT 40.395 149.190 40.685 149.235 ;
        RECT 41.300 149.190 41.620 149.250 ;
        RECT 40.395 149.050 41.620 149.190 ;
        RECT 40.395 149.005 40.685 149.050 ;
        RECT 41.300 148.990 41.620 149.050 ;
        RECT 42.680 148.990 43.000 149.250 ;
        RECT 44.060 149.190 44.380 149.250 ;
        RECT 46.360 149.190 46.680 149.250 ;
        RECT 49.580 149.235 49.900 149.250 ;
        RECT 49.365 149.190 49.900 149.235 ;
        RECT 44.060 149.050 49.900 149.190 ;
        RECT 44.060 148.990 44.380 149.050 ;
        RECT 46.360 148.990 46.680 149.050 ;
        RECT 49.365 149.005 49.900 149.050 ;
        RECT 49.580 148.990 49.900 149.005 ;
        RECT 61.080 148.990 61.400 149.250 ;
        RECT 65.695 149.005 65.985 149.235 ;
        RECT 67.075 149.190 67.365 149.235 ;
        RECT 69.360 149.190 69.680 149.250 ;
        RECT 67.075 149.050 69.680 149.190 ;
        RECT 67.075 149.005 67.365 149.050 ;
        RECT 25.200 148.850 25.520 148.910 ;
        RECT 26.530 148.850 26.820 148.895 ;
        RECT 29.790 148.850 30.080 148.895 ;
        RECT 25.200 148.710 30.080 148.850 ;
        RECT 25.200 148.650 25.520 148.710 ;
        RECT 26.530 148.665 26.820 148.710 ;
        RECT 29.790 148.665 30.080 148.710 ;
        RECT 30.710 148.850 31.000 148.895 ;
        RECT 32.570 148.850 32.860 148.895 ;
        RECT 47.755 148.850 48.045 148.895 ;
        RECT 51.370 148.850 51.660 148.895 ;
        RECT 54.630 148.850 54.920 148.895 ;
        RECT 30.710 148.710 32.860 148.850 ;
        RECT 30.710 148.665 31.000 148.710 ;
        RECT 32.570 148.665 32.860 148.710 ;
        RECT 36.330 148.710 39.230 148.850 ;
        RECT 28.390 148.510 28.680 148.555 ;
        RECT 30.710 148.510 30.925 148.665 ;
        RECT 28.390 148.370 30.925 148.510 ;
        RECT 28.390 148.325 28.680 148.370 ;
        RECT 31.640 148.310 31.960 148.570 ;
        RECT 35.320 148.510 35.640 148.570 ;
        RECT 36.330 148.555 36.470 148.710 ;
        RECT 36.255 148.510 36.545 148.555 ;
        RECT 38.555 148.510 38.845 148.555 ;
        RECT 35.320 148.370 36.545 148.510 ;
        RECT 35.320 148.310 35.640 148.370 ;
        RECT 36.255 148.325 36.545 148.370 ;
        RECT 37.250 148.370 38.845 148.510 ;
        RECT 33.495 148.170 33.785 148.215 ;
        RECT 34.860 148.170 35.180 148.230 ;
        RECT 33.495 148.030 35.180 148.170 ;
        RECT 33.495 147.985 33.785 148.030 ;
        RECT 34.860 147.970 35.180 148.030 ;
        RECT 36.700 147.970 37.020 148.230 ;
        RECT 28.390 147.830 28.680 147.875 ;
        RECT 31.170 147.830 31.460 147.875 ;
        RECT 33.030 147.830 33.320 147.875 ;
        RECT 28.390 147.690 33.320 147.830 ;
        RECT 28.390 147.645 28.680 147.690 ;
        RECT 31.170 147.645 31.460 147.690 ;
        RECT 33.030 147.645 33.320 147.690 ;
        RECT 34.400 147.830 34.720 147.890 ;
        RECT 37.250 147.830 37.390 148.370 ;
        RECT 38.555 148.325 38.845 148.370 ;
        RECT 39.090 148.170 39.230 148.710 ;
        RECT 39.550 148.710 41.990 148.850 ;
        RECT 39.550 148.570 39.690 148.710 ;
        RECT 39.460 148.310 39.780 148.570 ;
        RECT 39.920 148.510 40.240 148.570 ;
        RECT 41.850 148.555 41.990 148.710 ;
        RECT 47.755 148.710 54.920 148.850 ;
        RECT 47.755 148.665 48.045 148.710 ;
        RECT 51.370 148.665 51.660 148.710 ;
        RECT 54.630 148.665 54.920 148.710 ;
        RECT 55.550 148.850 55.840 148.895 ;
        RECT 57.410 148.850 57.700 148.895 ;
        RECT 55.550 148.710 57.700 148.850 ;
        RECT 55.550 148.665 55.840 148.710 ;
        RECT 57.410 148.665 57.700 148.710 ;
        RECT 57.860 148.850 58.180 148.910 ;
        RECT 63.855 148.850 64.145 148.895 ;
        RECT 57.860 148.710 64.145 148.850 ;
        RECT 40.855 148.510 41.145 148.555 ;
        RECT 39.920 148.370 41.145 148.510 ;
        RECT 39.920 148.310 40.240 148.370 ;
        RECT 40.855 148.325 41.145 148.370 ;
        RECT 41.775 148.510 42.065 148.555 ;
        RECT 44.075 148.510 44.365 148.555 ;
        RECT 47.295 148.510 47.585 148.555 ;
        RECT 48.200 148.510 48.520 148.570 ;
        RECT 49.580 148.510 49.900 148.570 ;
        RECT 41.775 148.370 47.050 148.510 ;
        RECT 41.775 148.325 42.065 148.370 ;
        RECT 44.075 148.325 44.365 148.370 ;
        RECT 44.995 148.170 45.285 148.215 ;
        RECT 39.090 148.030 45.285 148.170 ;
        RECT 46.910 148.170 47.050 148.370 ;
        RECT 47.295 148.370 49.900 148.510 ;
        RECT 47.295 148.325 47.585 148.370 ;
        RECT 48.200 148.310 48.520 148.370 ;
        RECT 49.580 148.310 49.900 148.370 ;
        RECT 53.230 148.510 53.520 148.555 ;
        RECT 55.550 148.510 55.765 148.665 ;
        RECT 57.860 148.650 58.180 148.710 ;
        RECT 63.855 148.665 64.145 148.710 ;
        RECT 53.230 148.370 55.765 148.510 ;
        RECT 56.020 148.510 56.340 148.570 ;
        RECT 56.495 148.510 56.785 148.555 ;
        RECT 56.020 148.370 56.785 148.510 ;
        RECT 53.230 148.325 53.520 148.370 ;
        RECT 56.020 148.310 56.340 148.370 ;
        RECT 56.495 148.325 56.785 148.370 ;
        RECT 56.940 148.510 57.260 148.570 ;
        RECT 58.335 148.510 58.625 148.555 ;
        RECT 59.240 148.510 59.560 148.570 ;
        RECT 56.940 148.370 59.560 148.510 ;
        RECT 56.940 148.310 57.260 148.370 ;
        RECT 58.335 148.325 58.625 148.370 ;
        RECT 59.240 148.310 59.560 148.370 ;
        RECT 59.700 148.510 60.020 148.570 ;
        RECT 60.635 148.510 60.925 148.555 ;
        RECT 65.770 148.510 65.910 149.005 ;
        RECT 69.360 148.990 69.680 149.050 ;
        RECT 69.820 149.190 70.140 149.250 ;
        RECT 69.820 149.050 72.810 149.190 ;
        RECT 69.820 148.990 70.140 149.050 ;
        RECT 67.995 148.850 68.285 148.895 ;
        RECT 70.755 148.850 71.045 148.895 ;
        RECT 67.995 148.710 71.045 148.850 ;
        RECT 67.995 148.665 68.285 148.710 ;
        RECT 70.755 148.665 71.045 148.710 ;
        RECT 72.670 148.850 72.810 149.050 ;
        RECT 86.855 149.005 87.145 149.235 ;
        RECT 93.280 149.190 93.600 149.250 ;
        RECT 96.040 149.190 96.360 149.250 ;
        RECT 93.280 149.050 96.360 149.190 ;
        RECT 75.800 148.850 76.120 148.910 ;
        RECT 72.670 148.710 76.120 148.850 ;
        RECT 66.155 148.510 66.445 148.555 ;
        RECT 59.700 148.370 60.925 148.510 ;
        RECT 59.700 148.310 60.020 148.370 ;
        RECT 60.635 148.325 60.925 148.370 ;
        RECT 61.170 148.370 64.530 148.510 ;
        RECT 65.770 148.370 66.445 148.510 ;
        RECT 61.170 148.170 61.310 148.370 ;
        RECT 46.910 148.030 61.310 148.170 ;
        RECT 44.995 147.985 45.285 148.030 ;
        RECT 62.935 147.985 63.225 148.215 ;
        RECT 63.395 148.170 63.685 148.215 ;
        RECT 63.840 148.170 64.160 148.230 ;
        RECT 63.395 148.030 64.160 148.170 ;
        RECT 64.390 148.170 64.530 148.370 ;
        RECT 66.155 148.325 66.445 148.370 ;
        RECT 68.900 148.310 69.220 148.570 ;
        RECT 69.375 148.510 69.665 148.555 ;
        RECT 71.660 148.510 71.980 148.570 ;
        RECT 72.670 148.555 72.810 148.710 ;
        RECT 75.800 148.650 76.120 148.710 ;
        RECT 76.275 148.850 76.565 148.895 ;
        RECT 79.430 148.850 79.720 148.895 ;
        RECT 82.690 148.850 82.980 148.895 ;
        RECT 76.275 148.710 82.980 148.850 ;
        RECT 76.275 148.665 76.565 148.710 ;
        RECT 79.430 148.665 79.720 148.710 ;
        RECT 82.690 148.665 82.980 148.710 ;
        RECT 83.610 148.850 83.900 148.895 ;
        RECT 85.470 148.850 85.760 148.895 ;
        RECT 86.930 148.850 87.070 149.005 ;
        RECT 93.280 148.990 93.600 149.050 ;
        RECT 96.040 148.990 96.360 149.050 ;
        RECT 83.610 148.710 85.760 148.850 ;
        RECT 83.610 148.665 83.900 148.710 ;
        RECT 85.470 148.665 85.760 148.710 ;
        RECT 86.010 148.710 87.070 148.850 ;
        RECT 89.155 148.850 89.445 148.895 ;
        RECT 91.915 148.850 92.205 148.895 ;
        RECT 89.155 148.710 92.205 148.850 ;
        RECT 69.375 148.370 71.980 148.510 ;
        RECT 69.375 148.325 69.665 148.370 ;
        RECT 71.660 148.310 71.980 148.370 ;
        RECT 72.135 148.325 72.425 148.555 ;
        RECT 72.595 148.325 72.885 148.555 ;
        RECT 73.055 148.325 73.345 148.555 ;
        RECT 73.975 148.510 74.265 148.555 ;
        RECT 74.420 148.510 74.740 148.570 ;
        RECT 73.975 148.370 74.740 148.510 ;
        RECT 73.975 148.325 74.265 148.370 ;
        RECT 67.520 148.170 67.840 148.230 ;
        RECT 64.390 148.030 67.840 148.170 ;
        RECT 63.395 147.985 63.685 148.030 ;
        RECT 34.400 147.690 37.390 147.830 ;
        RECT 53.230 147.830 53.520 147.875 ;
        RECT 56.010 147.830 56.300 147.875 ;
        RECT 57.870 147.830 58.160 147.875 ;
        RECT 53.230 147.690 58.160 147.830 ;
        RECT 63.010 147.830 63.150 147.985 ;
        RECT 63.840 147.970 64.160 148.030 ;
        RECT 67.520 147.970 67.840 148.030 ;
        RECT 67.980 148.170 68.300 148.230 ;
        RECT 72.210 148.170 72.350 148.325 ;
        RECT 67.980 148.030 69.590 148.170 ;
        RECT 67.980 147.970 68.300 148.030 ;
        RECT 69.450 147.890 69.590 148.030 ;
        RECT 70.600 148.030 72.350 148.170 ;
        RECT 73.130 148.170 73.270 148.325 ;
        RECT 74.420 148.310 74.740 148.370 ;
        RECT 76.735 148.510 77.025 148.555 ;
        RECT 79.940 148.510 80.260 148.570 ;
        RECT 81.290 148.510 81.580 148.555 ;
        RECT 83.610 148.510 83.825 148.665 ;
        RECT 76.735 148.370 81.090 148.510 ;
        RECT 76.735 148.325 77.025 148.370 ;
        RECT 79.940 148.310 80.260 148.370 ;
        RECT 77.425 148.170 77.715 148.215 ;
        RECT 78.560 148.170 78.880 148.230 ;
        RECT 73.130 148.030 78.880 148.170 ;
        RECT 80.950 148.170 81.090 148.370 ;
        RECT 81.290 148.370 83.825 148.510 ;
        RECT 84.555 148.510 84.845 148.555 ;
        RECT 86.010 148.510 86.150 148.710 ;
        RECT 89.155 148.665 89.445 148.710 ;
        RECT 91.915 148.665 92.205 148.710 ;
        RECT 92.360 148.850 92.680 148.910 ;
        RECT 95.595 148.850 95.885 148.895 ;
        RECT 97.880 148.850 98.200 148.910 ;
        RECT 92.360 148.710 95.350 148.850 ;
        RECT 92.360 148.650 92.680 148.710 ;
        RECT 84.555 148.370 86.150 148.510 ;
        RECT 81.290 148.325 81.580 148.370 ;
        RECT 84.555 148.325 84.845 148.370 ;
        RECT 86.380 148.310 86.700 148.570 ;
        RECT 87.760 148.310 88.080 148.570 ;
        RECT 88.680 148.510 89.000 148.570 ;
        RECT 90.075 148.510 90.365 148.555 ;
        RECT 88.680 148.370 90.365 148.510 ;
        RECT 88.680 148.310 89.000 148.370 ;
        RECT 90.075 148.325 90.365 148.370 ;
        RECT 90.535 148.510 90.825 148.555 ;
        RECT 90.980 148.510 91.300 148.570 ;
        RECT 90.535 148.370 91.300 148.510 ;
        RECT 90.535 148.325 90.825 148.370 ;
        RECT 90.980 148.310 91.300 148.370 ;
        RECT 93.280 148.310 93.600 148.570 ;
        RECT 93.755 148.325 94.045 148.555 ;
        RECT 83.620 148.170 83.940 148.230 ;
        RECT 80.950 148.030 83.940 148.170 ;
        RECT 64.300 147.830 64.620 147.890 ;
        RECT 66.140 147.830 66.460 147.890 ;
        RECT 63.010 147.690 66.460 147.830 ;
        RECT 34.400 147.630 34.720 147.690 ;
        RECT 53.230 147.645 53.520 147.690 ;
        RECT 56.010 147.645 56.300 147.690 ;
        RECT 57.870 147.645 58.160 147.690 ;
        RECT 64.300 147.630 64.620 147.690 ;
        RECT 66.140 147.630 66.460 147.690 ;
        RECT 69.360 147.830 69.680 147.890 ;
        RECT 70.600 147.830 70.740 148.030 ;
        RECT 77.425 147.985 77.715 148.030 ;
        RECT 78.560 147.970 78.880 148.030 ;
        RECT 83.620 147.970 83.940 148.030 ;
        RECT 69.360 147.690 70.740 147.830 ;
        RECT 81.290 147.830 81.580 147.875 ;
        RECT 84.070 147.830 84.360 147.875 ;
        RECT 85.930 147.830 86.220 147.875 ;
        RECT 81.290 147.690 86.220 147.830 ;
        RECT 86.470 147.830 86.610 148.310 ;
        RECT 89.600 148.170 89.920 148.230 ;
        RECT 93.830 148.170 93.970 148.325 ;
        RECT 94.200 148.310 94.520 148.570 ;
        RECT 95.210 148.555 95.350 148.710 ;
        RECT 95.595 148.710 98.200 148.850 ;
        RECT 95.595 148.665 95.885 148.710 ;
        RECT 97.880 148.650 98.200 148.710 ;
        RECT 102.020 148.850 102.340 148.910 ;
        RECT 104.730 148.850 105.020 148.895 ;
        RECT 107.990 148.850 108.280 148.895 ;
        RECT 102.020 148.710 108.280 148.850 ;
        RECT 102.020 148.650 102.340 148.710 ;
        RECT 104.730 148.665 105.020 148.710 ;
        RECT 107.990 148.665 108.280 148.710 ;
        RECT 108.910 148.850 109.200 148.895 ;
        RECT 110.770 148.850 111.060 148.895 ;
        RECT 108.910 148.710 111.060 148.850 ;
        RECT 108.910 148.665 109.200 148.710 ;
        RECT 110.770 148.665 111.060 148.710 ;
        RECT 95.135 148.325 95.425 148.555 ;
        RECT 96.040 148.510 96.360 148.570 ;
        RECT 96.975 148.510 97.265 148.555 ;
        RECT 96.040 148.370 97.265 148.510 ;
        RECT 96.040 148.310 96.360 148.370 ;
        RECT 96.975 148.325 97.265 148.370 ;
        RECT 106.590 148.510 106.880 148.555 ;
        RECT 108.910 148.510 109.125 148.665 ;
        RECT 106.590 148.370 109.125 148.510 ;
        RECT 106.590 148.325 106.880 148.370 ;
        RECT 109.840 148.310 110.160 148.570 ;
        RECT 111.220 148.510 111.540 148.570 ;
        RECT 111.695 148.510 111.985 148.555 ;
        RECT 111.220 148.370 111.985 148.510 ;
        RECT 111.220 148.310 111.540 148.370 ;
        RECT 111.695 148.325 111.985 148.370 ;
        RECT 89.600 148.030 93.970 148.170 ;
        RECT 96.515 148.170 96.805 148.215 ;
        RECT 97.420 148.170 97.740 148.230 ;
        RECT 96.515 148.030 97.740 148.170 ;
        RECT 89.600 147.970 89.920 148.030 ;
        RECT 96.515 147.985 96.805 148.030 ;
        RECT 97.420 147.970 97.740 148.030 ;
        RECT 90.060 147.830 90.380 147.890 ;
        RECT 86.470 147.690 90.380 147.830 ;
        RECT 69.360 147.630 69.680 147.690 ;
        RECT 81.290 147.645 81.580 147.690 ;
        RECT 84.070 147.645 84.360 147.690 ;
        RECT 85.930 147.645 86.220 147.690 ;
        RECT 90.060 147.630 90.380 147.690 ;
        RECT 106.590 147.830 106.880 147.875 ;
        RECT 109.370 147.830 109.660 147.875 ;
        RECT 111.230 147.830 111.520 147.875 ;
        RECT 106.590 147.690 111.520 147.830 ;
        RECT 106.590 147.645 106.880 147.690 ;
        RECT 109.370 147.645 109.660 147.690 ;
        RECT 111.230 147.645 111.520 147.690 ;
        RECT 24.525 147.490 24.815 147.535 ;
        RECT 29.800 147.490 30.120 147.550 ;
        RECT 24.525 147.350 30.120 147.490 ;
        RECT 24.525 147.305 24.815 147.350 ;
        RECT 29.800 147.290 30.120 147.350 ;
        RECT 30.260 147.490 30.580 147.550 ;
        RECT 33.955 147.490 34.245 147.535 ;
        RECT 30.260 147.350 34.245 147.490 ;
        RECT 30.260 147.290 30.580 147.350 ;
        RECT 33.955 147.305 34.245 147.350 ;
        RECT 37.620 147.490 37.940 147.550 ;
        RECT 43.155 147.490 43.445 147.535 ;
        RECT 37.620 147.350 43.445 147.490 ;
        RECT 37.620 147.290 37.940 147.350 ;
        RECT 43.155 147.305 43.445 147.350 ;
        RECT 67.060 147.490 67.380 147.550 ;
        RECT 67.995 147.490 68.285 147.535 ;
        RECT 67.060 147.350 68.285 147.490 ;
        RECT 67.060 147.290 67.380 147.350 ;
        RECT 67.995 147.305 68.285 147.350 ;
        RECT 69.820 147.490 70.140 147.550 ;
        RECT 70.295 147.490 70.585 147.535 ;
        RECT 69.820 147.350 70.585 147.490 ;
        RECT 69.820 147.290 70.140 147.350 ;
        RECT 70.295 147.305 70.585 147.350 ;
        RECT 89.600 147.290 89.920 147.550 ;
        RECT 91.440 147.290 91.760 147.550 ;
        RECT 96.960 147.290 97.280 147.550 ;
        RECT 97.880 147.290 98.200 147.550 ;
        RECT 102.725 147.490 103.015 147.535 ;
        RECT 103.860 147.490 104.180 147.550 ;
        RECT 102.725 147.350 104.180 147.490 ;
        RECT 102.725 147.305 103.015 147.350 ;
        RECT 103.860 147.290 104.180 147.350 ;
        RECT 22.830 146.670 113.450 147.150 ;
        RECT 25.200 146.270 25.520 146.530 ;
        RECT 30.720 146.470 31.040 146.530 ;
        RECT 34.400 146.470 34.720 146.530 ;
        RECT 35.320 146.515 35.640 146.530 ;
        RECT 30.720 146.330 34.720 146.470 ;
        RECT 30.720 146.270 31.040 146.330 ;
        RECT 34.400 146.270 34.720 146.330 ;
        RECT 35.105 146.285 35.640 146.515 ;
        RECT 35.320 146.270 35.640 146.285 ;
        RECT 38.540 146.270 38.860 146.530 ;
        RECT 48.215 146.470 48.505 146.515 ;
        RECT 51.895 146.470 52.185 146.515 ;
        RECT 57.415 146.470 57.705 146.515 ;
        RECT 48.215 146.330 52.185 146.470 ;
        RECT 48.215 146.285 48.505 146.330 ;
        RECT 51.895 146.285 52.185 146.330 ;
        RECT 54.730 146.330 57.705 146.470 ;
        RECT 26.600 146.130 26.890 146.175 ;
        RECT 28.460 146.130 28.750 146.175 ;
        RECT 31.240 146.130 31.530 146.175 ;
        RECT 26.600 145.990 31.530 146.130 ;
        RECT 26.600 145.945 26.890 145.990 ;
        RECT 28.460 145.945 28.750 145.990 ;
        RECT 31.240 145.945 31.530 145.990 ;
        RECT 35.780 146.130 36.100 146.190 ;
        RECT 54.730 146.130 54.870 146.330 ;
        RECT 57.415 146.285 57.705 146.330 ;
        RECT 59.715 146.470 60.005 146.515 ;
        RECT 60.160 146.470 60.480 146.530 ;
        RECT 59.715 146.330 60.480 146.470 ;
        RECT 59.715 146.285 60.005 146.330 ;
        RECT 60.160 146.270 60.480 146.330 ;
        RECT 89.600 146.270 89.920 146.530 ;
        RECT 96.975 146.470 97.265 146.515 ;
        RECT 98.340 146.470 98.660 146.530 ;
        RECT 96.975 146.330 98.660 146.470 ;
        RECT 96.975 146.285 97.265 146.330 ;
        RECT 98.340 146.270 98.660 146.330 ;
        RECT 35.780 145.990 41.990 146.130 ;
        RECT 35.780 145.930 36.100 145.990 ;
        RECT 27.975 145.790 28.265 145.835 ;
        RECT 29.340 145.790 29.660 145.850 ;
        RECT 27.975 145.650 29.660 145.790 ;
        RECT 27.975 145.605 28.265 145.650 ;
        RECT 29.340 145.590 29.660 145.650 ;
        RECT 29.800 145.790 30.120 145.850 ;
        RECT 41.850 145.835 41.990 145.990 ;
        RECT 52.430 145.990 54.870 146.130 ;
        RECT 56.020 146.130 56.340 146.190 ;
        RECT 64.300 146.130 64.620 146.190 ;
        RECT 66.140 146.130 66.460 146.190 ;
        RECT 56.020 145.990 66.460 146.130 ;
        RECT 36.715 145.790 37.005 145.835 ;
        RECT 41.315 145.790 41.605 145.835 ;
        RECT 29.800 145.650 41.605 145.790 ;
        RECT 29.800 145.590 30.120 145.650 ;
        RECT 36.715 145.605 37.005 145.650 ;
        RECT 41.315 145.605 41.605 145.650 ;
        RECT 41.775 145.605 42.065 145.835 ;
        RECT 46.375 145.790 46.665 145.835 ;
        RECT 52.430 145.790 52.570 145.990 ;
        RECT 56.020 145.930 56.340 145.990 ;
        RECT 43.230 145.650 46.665 145.790 ;
        RECT 25.660 145.250 25.980 145.510 ;
        RECT 26.135 145.265 26.425 145.495 ;
        RECT 31.240 145.450 31.530 145.495 ;
        RECT 28.995 145.310 31.530 145.450 ;
        RECT 26.210 144.770 26.350 145.265 ;
        RECT 28.995 145.155 29.210 145.310 ;
        RECT 31.240 145.265 31.530 145.310 ;
        RECT 37.635 145.450 37.925 145.495 ;
        RECT 39.460 145.450 39.780 145.510 ;
        RECT 43.230 145.450 43.370 145.650 ;
        RECT 46.375 145.605 46.665 145.650 ;
        RECT 46.910 145.650 52.570 145.790 ;
        RECT 37.635 145.310 39.780 145.450 ;
        RECT 37.635 145.265 37.925 145.310 ;
        RECT 39.460 145.250 39.780 145.310 ;
        RECT 40.930 145.310 43.370 145.450 ;
        RECT 27.060 145.110 27.350 145.155 ;
        RECT 28.920 145.110 29.210 145.155 ;
        RECT 27.060 144.970 29.210 145.110 ;
        RECT 27.060 144.925 27.350 144.970 ;
        RECT 28.920 144.925 29.210 144.970 ;
        RECT 29.800 145.155 30.120 145.170 ;
        RECT 29.800 145.110 30.130 145.155 ;
        RECT 33.100 145.110 33.390 145.155 ;
        RECT 29.800 144.970 33.390 145.110 ;
        RECT 29.800 144.925 30.130 144.970 ;
        RECT 33.100 144.925 33.390 144.970 ;
        RECT 29.800 144.910 30.120 144.925 ;
        RECT 40.930 144.830 41.070 145.310 ;
        RECT 44.060 145.250 44.380 145.510 ;
        RECT 44.995 145.265 45.285 145.495 ;
        RECT 45.915 145.450 46.205 145.495 ;
        RECT 46.910 145.450 47.050 145.650 ;
        RECT 52.800 145.590 53.120 145.850 ;
        RECT 58.320 145.590 58.640 145.850 ;
        RECT 63.010 145.835 63.150 145.990 ;
        RECT 64.300 145.930 64.620 145.990 ;
        RECT 66.140 145.930 66.460 145.990 ;
        RECT 71.660 146.130 71.980 146.190 ;
        RECT 78.100 146.130 78.420 146.190 ;
        RECT 85.460 146.130 85.780 146.190 ;
        RECT 103.400 146.130 103.720 146.190 ;
        RECT 71.660 145.990 80.170 146.130 ;
        RECT 71.660 145.930 71.980 145.990 ;
        RECT 78.100 145.930 78.420 145.990 ;
        RECT 62.935 145.605 63.225 145.835 ;
        RECT 69.360 145.790 69.680 145.850 ;
        RECT 63.470 145.650 76.490 145.790 ;
        RECT 45.915 145.310 47.050 145.450 ;
        RECT 45.915 145.265 46.205 145.310 ;
        RECT 47.295 145.265 47.585 145.495 ;
        RECT 45.070 145.110 45.210 145.265 ;
        RECT 47.370 145.110 47.510 145.265 ;
        RECT 51.880 145.250 52.200 145.510 ;
        RECT 53.275 145.450 53.565 145.495 ;
        RECT 53.720 145.450 54.040 145.510 ;
        RECT 53.275 145.310 54.040 145.450 ;
        RECT 53.275 145.265 53.565 145.310 ;
        RECT 53.720 145.250 54.040 145.310 ;
        RECT 58.780 145.250 59.100 145.510 ;
        RECT 63.470 145.450 63.610 145.650 ;
        RECT 69.360 145.590 69.680 145.650 ;
        RECT 59.330 145.310 63.610 145.450 ;
        RECT 45.070 144.970 56.940 145.110 ;
        RECT 52.430 144.830 52.570 144.970 ;
        RECT 34.860 144.770 35.180 144.830 ;
        RECT 26.210 144.630 35.180 144.770 ;
        RECT 34.860 144.570 35.180 144.630 ;
        RECT 36.240 144.770 36.560 144.830 ;
        RECT 39.015 144.770 39.305 144.815 ;
        RECT 36.240 144.630 39.305 144.770 ;
        RECT 36.240 144.570 36.560 144.630 ;
        RECT 39.015 144.585 39.305 144.630 ;
        RECT 40.840 144.570 41.160 144.830 ;
        RECT 52.340 144.570 52.660 144.830 ;
        RECT 54.195 144.770 54.485 144.815 ;
        RECT 55.100 144.770 55.420 144.830 ;
        RECT 54.195 144.630 55.420 144.770 ;
        RECT 56.800 144.770 56.940 144.970 ;
        RECT 57.400 144.910 57.720 145.170 ;
        RECT 57.860 145.110 58.180 145.170 ;
        RECT 59.330 145.110 59.470 145.310 ;
        RECT 63.840 145.250 64.160 145.510 ;
        RECT 66.600 145.250 66.920 145.510 ;
        RECT 67.995 145.265 68.285 145.495 ;
        RECT 64.760 145.110 65.080 145.170 ;
        RECT 68.070 145.110 68.210 145.265 ;
        RECT 74.420 145.250 74.740 145.510 ;
        RECT 75.355 145.265 75.645 145.495 ;
        RECT 57.860 144.970 59.470 145.110 ;
        RECT 59.790 144.970 65.080 145.110 ;
        RECT 57.860 144.910 58.180 144.970 ;
        RECT 59.790 144.770 59.930 144.970 ;
        RECT 64.760 144.910 65.080 144.970 ;
        RECT 65.770 144.970 68.210 145.110 ;
        RECT 75.430 145.110 75.570 145.265 ;
        RECT 75.800 145.250 76.120 145.510 ;
        RECT 76.350 145.495 76.490 145.650 ;
        RECT 76.275 145.265 76.565 145.495 ;
        RECT 80.030 145.450 80.170 145.990 ;
        RECT 80.490 145.990 103.720 146.130 ;
        RECT 80.490 145.835 80.630 145.990 ;
        RECT 85.460 145.930 85.780 145.990 ;
        RECT 91.070 145.835 91.210 145.990 ;
        RECT 80.415 145.605 80.705 145.835 ;
        RECT 90.995 145.605 91.285 145.835 ;
        RECT 94.215 145.790 94.505 145.835 ;
        RECT 94.660 145.790 94.980 145.850 ;
        RECT 103.030 145.835 103.170 145.990 ;
        RECT 103.400 145.930 103.720 145.990 ;
        RECT 94.215 145.650 94.980 145.790 ;
        RECT 94.215 145.605 94.505 145.650 ;
        RECT 94.660 145.590 94.980 145.650 ;
        RECT 95.210 145.650 98.110 145.790 ;
        RECT 80.860 145.450 81.180 145.510 ;
        RECT 83.635 145.450 83.925 145.495 ;
        RECT 80.030 145.310 81.180 145.450 ;
        RECT 80.860 145.250 81.180 145.310 ;
        RECT 83.250 145.310 83.925 145.450 ;
        RECT 81.320 145.110 81.640 145.170 ;
        RECT 75.430 144.970 81.640 145.110 ;
        RECT 56.800 144.630 59.930 144.770 ;
        RECT 63.395 144.770 63.685 144.815 ;
        RECT 65.220 144.770 65.540 144.830 ;
        RECT 65.770 144.815 65.910 144.970 ;
        RECT 81.320 144.910 81.640 144.970 ;
        RECT 63.395 144.630 65.540 144.770 ;
        RECT 54.195 144.585 54.485 144.630 ;
        RECT 55.100 144.570 55.420 144.630 ;
        RECT 63.395 144.585 63.685 144.630 ;
        RECT 65.220 144.570 65.540 144.630 ;
        RECT 65.695 144.585 65.985 144.815 ;
        RECT 67.075 144.770 67.365 144.815 ;
        RECT 67.520 144.770 67.840 144.830 ;
        RECT 67.075 144.630 67.840 144.770 ;
        RECT 67.075 144.585 67.365 144.630 ;
        RECT 67.520 144.570 67.840 144.630 ;
        RECT 67.980 144.770 68.300 144.830 ;
        RECT 68.915 144.770 69.205 144.815 ;
        RECT 67.980 144.630 69.205 144.770 ;
        RECT 67.980 144.570 68.300 144.630 ;
        RECT 68.915 144.585 69.205 144.630 ;
        RECT 74.880 144.770 75.200 144.830 ;
        RECT 83.250 144.815 83.390 145.310 ;
        RECT 83.635 145.265 83.925 145.310 ;
        RECT 87.760 145.250 88.080 145.510 ;
        RECT 88.680 145.450 89.000 145.510 ;
        RECT 95.210 145.495 95.350 145.650 ;
        RECT 95.135 145.450 95.425 145.495 ;
        RECT 88.680 145.310 95.425 145.450 ;
        RECT 88.680 145.250 89.000 145.310 ;
        RECT 95.135 145.265 95.425 145.310 ;
        RECT 96.055 145.450 96.345 145.495 ;
        RECT 96.500 145.450 96.820 145.510 ;
        RECT 96.055 145.310 96.820 145.450 ;
        RECT 96.055 145.265 96.345 145.310 ;
        RECT 96.500 145.250 96.820 145.310 ;
        RECT 97.420 145.450 97.740 145.510 ;
        RECT 97.970 145.495 98.110 145.650 ;
        RECT 102.955 145.605 103.245 145.835 ;
        RECT 97.895 145.450 98.185 145.495 ;
        RECT 97.420 145.310 98.185 145.450 ;
        RECT 97.420 145.250 97.740 145.310 ;
        RECT 97.895 145.265 98.185 145.310 ;
        RECT 98.800 145.250 99.120 145.510 ;
        RECT 103.860 145.250 104.180 145.510 ;
        RECT 107.555 145.450 107.845 145.495 ;
        RECT 105.790 145.310 107.845 145.450 ;
        RECT 91.915 145.110 92.205 145.155 ;
        RECT 94.200 145.110 94.520 145.170 ;
        RECT 91.915 144.970 103.630 145.110 ;
        RECT 91.915 144.925 92.205 144.970 ;
        RECT 94.200 144.910 94.520 144.970 ;
        RECT 103.490 144.830 103.630 144.970 ;
        RECT 77.655 144.770 77.945 144.815 ;
        RECT 74.880 144.630 77.945 144.770 ;
        RECT 74.880 144.570 75.200 144.630 ;
        RECT 77.655 144.585 77.945 144.630 ;
        RECT 83.175 144.585 83.465 144.815 ;
        RECT 84.540 144.570 84.860 144.830 ;
        RECT 90.980 144.770 91.300 144.830 ;
        RECT 91.455 144.770 91.745 144.815 ;
        RECT 90.980 144.630 91.745 144.770 ;
        RECT 90.980 144.570 91.300 144.630 ;
        RECT 91.455 144.585 91.745 144.630 ;
        RECT 93.755 144.770 94.045 144.815 ;
        RECT 94.660 144.770 94.980 144.830 ;
        RECT 93.755 144.630 94.980 144.770 ;
        RECT 93.755 144.585 94.045 144.630 ;
        RECT 94.660 144.570 94.980 144.630 ;
        RECT 103.400 144.570 103.720 144.830 ;
        RECT 105.790 144.815 105.930 145.310 ;
        RECT 107.555 145.265 107.845 145.310 ;
        RECT 105.715 144.585 106.005 144.815 ;
        RECT 108.475 144.770 108.765 144.815 ;
        RECT 109.380 144.770 109.700 144.830 ;
        RECT 108.475 144.630 109.700 144.770 ;
        RECT 108.475 144.585 108.765 144.630 ;
        RECT 109.380 144.570 109.700 144.630 ;
        RECT 22.830 143.950 113.450 144.430 ;
        RECT 29.340 143.550 29.660 143.810 ;
        RECT 32.115 143.750 32.405 143.795 ;
        RECT 30.390 143.610 32.405 143.750 ;
        RECT 27.055 143.410 27.345 143.455 ;
        RECT 29.800 143.410 30.120 143.470 ;
        RECT 27.055 143.270 30.120 143.410 ;
        RECT 27.055 143.225 27.345 143.270 ;
        RECT 29.800 143.210 30.120 143.270 ;
        RECT 26.120 143.070 26.440 143.130 ;
        RECT 26.595 143.070 26.885 143.115 ;
        RECT 27.500 143.070 27.820 143.130 ;
        RECT 26.120 142.930 27.820 143.070 ;
        RECT 26.120 142.870 26.440 142.930 ;
        RECT 26.595 142.885 26.885 142.930 ;
        RECT 27.500 142.870 27.820 142.930 ;
        RECT 27.975 142.885 28.265 143.115 ;
        RECT 28.420 143.070 28.740 143.130 ;
        RECT 30.390 143.115 30.530 143.610 ;
        RECT 32.115 143.565 32.405 143.610 ;
        RECT 33.955 143.750 34.245 143.795 ;
        RECT 35.320 143.750 35.640 143.810 ;
        RECT 40.840 143.750 41.160 143.810 ;
        RECT 45.225 143.750 45.515 143.795 ;
        RECT 33.955 143.610 35.640 143.750 ;
        RECT 33.955 143.565 34.245 143.610 ;
        RECT 35.320 143.550 35.640 143.610 ;
        RECT 36.790 143.610 39.690 143.750 ;
        RECT 36.790 143.410 36.930 143.610 ;
        RECT 34.490 143.270 36.930 143.410 ;
        RECT 37.180 143.410 37.470 143.455 ;
        RECT 39.040 143.410 39.330 143.455 ;
        RECT 37.180 143.270 39.330 143.410 ;
        RECT 39.550 143.410 39.690 143.610 ;
        RECT 40.840 143.610 45.515 143.750 ;
        RECT 40.840 143.550 41.160 143.610 ;
        RECT 45.225 143.565 45.515 143.610 ;
        RECT 45.900 143.750 46.220 143.810 ;
        RECT 49.580 143.750 49.900 143.810 ;
        RECT 45.900 143.610 49.900 143.750 ;
        RECT 45.900 143.550 46.220 143.610 ;
        RECT 49.580 143.550 49.900 143.610 ;
        RECT 52.355 143.750 52.645 143.795 ;
        RECT 53.720 143.750 54.040 143.810 ;
        RECT 52.355 143.610 54.040 143.750 ;
        RECT 52.355 143.565 52.645 143.610 ;
        RECT 53.720 143.550 54.040 143.610 ;
        RECT 56.955 143.750 57.245 143.795 ;
        RECT 57.400 143.750 57.720 143.810 ;
        RECT 56.955 143.610 57.720 143.750 ;
        RECT 56.955 143.565 57.245 143.610 ;
        RECT 57.400 143.550 57.720 143.610 ;
        RECT 58.320 143.750 58.640 143.810 ;
        RECT 62.000 143.750 62.320 143.810 ;
        RECT 58.320 143.610 62.320 143.750 ;
        RECT 58.320 143.550 58.640 143.610 ;
        RECT 62.000 143.550 62.320 143.610 ;
        RECT 70.280 143.750 70.600 143.810 ;
        RECT 78.100 143.795 78.420 143.810 ;
        RECT 70.280 143.610 76.490 143.750 ;
        RECT 70.280 143.550 70.600 143.610 ;
        RECT 39.960 143.410 40.250 143.455 ;
        RECT 43.220 143.410 43.510 143.455 ;
        RECT 39.550 143.270 43.510 143.410 ;
        RECT 28.420 142.930 30.030 143.070 ;
        RECT 28.050 142.730 28.190 142.885 ;
        RECT 28.420 142.870 28.740 142.930 ;
        RECT 29.340 142.730 29.660 142.790 ;
        RECT 28.050 142.590 29.660 142.730 ;
        RECT 29.890 142.730 30.030 142.930 ;
        RECT 30.275 142.885 30.565 143.115 ;
        RECT 30.735 142.885 31.025 143.115 ;
        RECT 31.195 143.070 31.485 143.115 ;
        RECT 34.490 143.070 34.630 143.270 ;
        RECT 37.180 143.225 37.470 143.270 ;
        RECT 39.040 143.225 39.330 143.270 ;
        RECT 39.960 143.225 40.250 143.270 ;
        RECT 43.220 143.225 43.510 143.270 ;
        RECT 46.360 143.410 46.680 143.470 ;
        RECT 48.215 143.410 48.505 143.455 ;
        RECT 61.080 143.410 61.400 143.470 ;
        RECT 46.360 143.270 48.505 143.410 ;
        RECT 31.195 142.930 34.630 143.070 ;
        RECT 34.860 143.070 35.180 143.130 ;
        RECT 36.255 143.070 36.545 143.115 ;
        RECT 34.860 142.930 36.545 143.070 ;
        RECT 39.115 143.070 39.330 143.225 ;
        RECT 46.360 143.210 46.680 143.270 ;
        RECT 48.215 143.225 48.505 143.270 ;
        RECT 59.790 143.270 61.400 143.410 ;
        RECT 41.360 143.070 41.650 143.115 ;
        RECT 39.115 142.930 41.650 143.070 ;
        RECT 31.195 142.885 31.485 142.930 ;
        RECT 30.770 142.730 30.910 142.885 ;
        RECT 34.860 142.870 35.180 142.930 ;
        RECT 36.255 142.885 36.545 142.930 ;
        RECT 41.360 142.885 41.650 142.930 ;
        RECT 45.440 143.070 45.760 143.130 ;
        RECT 46.835 143.070 47.125 143.115 ;
        RECT 45.440 142.930 47.125 143.070 ;
        RECT 45.440 142.870 45.760 142.930 ;
        RECT 46.835 142.885 47.125 142.930 ;
        RECT 47.280 142.870 47.600 143.130 ;
        RECT 49.135 143.070 49.425 143.115 ;
        RECT 49.580 143.070 49.900 143.130 ;
        RECT 49.135 142.930 49.900 143.070 ;
        RECT 49.135 142.885 49.425 142.930 ;
        RECT 49.580 142.870 49.900 142.930 ;
        RECT 50.500 143.070 50.820 143.130 ;
        RECT 56.020 143.070 56.340 143.130 ;
        RECT 50.500 142.930 56.340 143.070 ;
        RECT 50.500 142.870 50.820 142.930 ;
        RECT 29.890 142.590 30.910 142.730 ;
        RECT 29.340 142.530 29.660 142.590 ;
        RECT 34.400 142.530 34.720 142.790 ;
        RECT 35.320 142.530 35.640 142.790 ;
        RECT 35.780 142.730 36.100 142.790 ;
        RECT 38.095 142.730 38.385 142.775 ;
        RECT 35.780 142.590 38.385 142.730 ;
        RECT 35.780 142.530 36.100 142.590 ;
        RECT 38.095 142.545 38.385 142.590 ;
        RECT 52.800 142.530 53.120 142.790 ;
        RECT 53.350 142.775 53.490 142.930 ;
        RECT 56.020 142.870 56.340 142.930 ;
        RECT 57.860 143.085 58.180 143.130 ;
        RECT 58.335 143.085 58.625 143.115 ;
        RECT 57.860 142.945 58.625 143.085 ;
        RECT 57.860 142.870 58.180 142.945 ;
        RECT 58.335 142.885 58.625 142.945 ;
        RECT 58.780 142.870 59.100 143.130 ;
        RECT 59.360 143.085 59.650 143.130 ;
        RECT 59.790 143.085 59.930 143.270 ;
        RECT 61.080 143.210 61.400 143.270 ;
        RECT 62.870 143.410 63.160 143.455 ;
        RECT 63.380 143.410 63.700 143.470 ;
        RECT 66.130 143.410 66.420 143.455 ;
        RECT 62.870 143.270 66.420 143.410 ;
        RECT 62.870 143.225 63.160 143.270 ;
        RECT 63.380 143.210 63.700 143.270 ;
        RECT 66.130 143.225 66.420 143.270 ;
        RECT 67.050 143.410 67.340 143.455 ;
        RECT 68.910 143.410 69.200 143.455 ;
        RECT 67.050 143.270 69.200 143.410 ;
        RECT 67.050 143.225 67.340 143.270 ;
        RECT 68.910 143.225 69.200 143.270 ;
        RECT 69.360 143.410 69.680 143.470 ;
        RECT 69.360 143.270 73.730 143.410 ;
        RECT 59.360 142.945 59.930 143.085 ;
        RECT 60.175 143.070 60.465 143.115 ;
        RECT 61.540 143.070 61.860 143.130 ;
        RECT 59.360 142.900 59.650 142.945 ;
        RECT 60.175 142.930 61.860 143.070 ;
        RECT 60.175 142.885 60.465 142.930 ;
        RECT 61.540 142.870 61.860 142.930 ;
        RECT 64.730 143.070 65.020 143.115 ;
        RECT 67.050 143.070 67.265 143.225 ;
        RECT 69.360 143.210 69.680 143.270 ;
        RECT 64.730 142.930 67.265 143.070 ;
        RECT 64.730 142.885 65.020 142.930 ;
        RECT 67.980 142.870 68.300 143.130 ;
        RECT 69.835 143.070 70.125 143.115 ;
        RECT 70.280 143.070 70.600 143.130 ;
        RECT 69.835 142.930 70.600 143.070 ;
        RECT 69.835 142.885 70.125 142.930 ;
        RECT 70.280 142.870 70.600 142.930 ;
        RECT 70.755 143.020 71.045 143.115 ;
        RECT 70.755 142.885 71.430 143.020 ;
        RECT 70.830 142.880 71.430 142.885 ;
        RECT 53.275 142.545 53.565 142.775 ;
        RECT 60.620 142.730 60.940 142.790 ;
        RECT 60.620 142.590 70.740 142.730 ;
        RECT 60.620 142.530 60.940 142.590 ;
        RECT 28.895 142.390 29.185 142.435 ;
        RECT 32.100 142.390 32.420 142.450 ;
        RECT 28.895 142.250 32.420 142.390 ;
        RECT 28.895 142.205 29.185 142.250 ;
        RECT 32.100 142.190 32.420 142.250 ;
        RECT 36.720 142.390 37.010 142.435 ;
        RECT 38.580 142.390 38.870 142.435 ;
        RECT 41.360 142.390 41.650 142.435 ;
        RECT 36.720 142.250 41.650 142.390 ;
        RECT 36.720 142.205 37.010 142.250 ;
        RECT 38.580 142.205 38.870 142.250 ;
        RECT 41.360 142.205 41.650 142.250 ;
        RECT 42.680 142.390 43.000 142.450 ;
        RECT 58.780 142.390 59.100 142.450 ;
        RECT 60.710 142.390 60.850 142.530 ;
        RECT 42.680 142.250 47.050 142.390 ;
        RECT 42.680 142.190 43.000 142.250 ;
        RECT 30.720 142.050 31.040 142.110 ;
        RECT 34.400 142.050 34.720 142.110 ;
        RECT 30.720 141.910 34.720 142.050 ;
        RECT 30.720 141.850 31.040 141.910 ;
        RECT 34.400 141.850 34.720 141.910 ;
        RECT 45.440 142.050 45.760 142.110 ;
        RECT 46.910 142.095 47.050 142.250 ;
        RECT 58.780 142.250 60.850 142.390 ;
        RECT 64.730 142.390 65.020 142.435 ;
        RECT 67.510 142.390 67.800 142.435 ;
        RECT 69.370 142.390 69.660 142.435 ;
        RECT 64.730 142.250 69.660 142.390 ;
        RECT 58.780 142.190 59.100 142.250 ;
        RECT 64.730 142.205 65.020 142.250 ;
        RECT 67.510 142.205 67.800 142.250 ;
        RECT 69.370 142.205 69.660 142.250 ;
        RECT 45.915 142.050 46.205 142.095 ;
        RECT 45.440 141.910 46.205 142.050 ;
        RECT 45.440 141.850 45.760 141.910 ;
        RECT 45.915 141.865 46.205 141.910 ;
        RECT 46.835 141.865 47.125 142.095 ;
        RECT 49.580 141.850 49.900 142.110 ;
        RECT 50.515 142.050 50.805 142.095 ;
        RECT 51.880 142.050 52.200 142.110 ;
        RECT 61.080 142.095 61.400 142.110 ;
        RECT 50.515 141.910 52.200 142.050 ;
        RECT 50.515 141.865 50.805 141.910 ;
        RECT 51.880 141.850 52.200 141.910 ;
        RECT 60.865 142.050 61.400 142.095 ;
        RECT 65.220 142.050 65.540 142.110 ;
        RECT 60.865 141.910 65.540 142.050 ;
        RECT 70.600 142.050 70.740 142.590 ;
        RECT 71.290 142.390 71.430 142.880 ;
        RECT 71.660 142.870 71.980 143.130 ;
        RECT 72.120 142.870 72.440 143.130 ;
        RECT 72.595 143.060 72.885 143.115 ;
        RECT 73.590 143.070 73.730 143.270 ;
        RECT 74.880 143.210 75.200 143.470 ;
        RECT 76.350 143.115 76.490 143.610 ;
        RECT 77.885 143.565 78.420 143.795 ;
        RECT 78.100 143.550 78.420 143.565 ;
        RECT 81.320 143.750 81.640 143.810 ;
        RECT 87.545 143.750 87.835 143.795 ;
        RECT 90.980 143.750 91.300 143.810 ;
        RECT 81.320 143.610 91.300 143.750 ;
        RECT 81.320 143.550 81.640 143.610 ;
        RECT 87.545 143.565 87.835 143.610 ;
        RECT 90.980 143.550 91.300 143.610 ;
        RECT 96.960 143.550 97.280 143.810 ;
        RECT 102.265 143.750 102.555 143.795 ;
        RECT 103.400 143.750 103.720 143.810 ;
        RECT 102.265 143.610 103.720 143.750 ;
        RECT 102.265 143.565 102.555 143.610 ;
        RECT 103.400 143.550 103.720 143.610 ;
        RECT 83.160 143.455 83.480 143.470 ;
        RECT 89.600 143.455 89.920 143.470 ;
        RECT 79.890 143.410 80.180 143.455 ;
        RECT 83.150 143.410 83.480 143.455 ;
        RECT 79.890 143.270 83.480 143.410 ;
        RECT 79.890 143.225 80.180 143.270 ;
        RECT 83.150 143.225 83.480 143.270 ;
        RECT 83.160 143.210 83.480 143.225 ;
        RECT 84.070 143.410 84.360 143.455 ;
        RECT 85.930 143.410 86.220 143.455 ;
        RECT 84.070 143.270 86.220 143.410 ;
        RECT 84.070 143.225 84.360 143.270 ;
        RECT 85.930 143.225 86.220 143.270 ;
        RECT 89.550 143.410 89.920 143.455 ;
        RECT 92.810 143.410 93.100 143.455 ;
        RECT 89.550 143.270 93.100 143.410 ;
        RECT 89.550 143.225 89.920 143.270 ;
        RECT 92.810 143.225 93.100 143.270 ;
        RECT 93.730 143.410 94.020 143.455 ;
        RECT 95.590 143.410 95.880 143.455 ;
        RECT 93.730 143.270 95.880 143.410 ;
        RECT 93.730 143.225 94.020 143.270 ;
        RECT 95.590 143.225 95.880 143.270 ;
        RECT 101.115 143.410 101.405 143.455 ;
        RECT 104.270 143.410 104.560 143.455 ;
        RECT 107.530 143.410 107.820 143.455 ;
        RECT 101.115 143.270 107.820 143.410 ;
        RECT 101.115 143.225 101.405 143.270 ;
        RECT 104.270 143.225 104.560 143.270 ;
        RECT 107.530 143.225 107.820 143.270 ;
        RECT 108.450 143.410 108.740 143.455 ;
        RECT 110.310 143.410 110.600 143.455 ;
        RECT 108.450 143.270 110.600 143.410 ;
        RECT 108.450 143.225 108.740 143.270 ;
        RECT 110.310 143.225 110.600 143.270 ;
        RECT 73.130 143.060 73.730 143.070 ;
        RECT 72.595 142.930 73.730 143.060 ;
        RECT 72.595 142.920 73.270 142.930 ;
        RECT 72.595 142.885 72.885 142.920 ;
        RECT 76.275 142.885 76.565 143.115 ;
        RECT 81.750 143.070 82.040 143.115 ;
        RECT 84.070 143.070 84.285 143.225 ;
        RECT 89.600 143.210 89.920 143.225 ;
        RECT 81.750 142.930 84.285 143.070 ;
        RECT 84.540 143.070 84.860 143.130 ;
        RECT 85.015 143.070 85.305 143.115 ;
        RECT 84.540 142.930 85.305 143.070 ;
        RECT 81.750 142.885 82.040 142.930 ;
        RECT 84.540 142.870 84.860 142.930 ;
        RECT 85.015 142.885 85.305 142.930 ;
        RECT 91.410 143.070 91.700 143.115 ;
        RECT 93.730 143.070 93.945 143.225 ;
        RECT 91.410 142.930 93.945 143.070 ;
        RECT 97.420 143.070 97.740 143.130 ;
        RECT 97.895 143.070 98.185 143.115 ;
        RECT 97.420 142.930 98.185 143.070 ;
        RECT 91.410 142.885 91.700 142.930 ;
        RECT 97.420 142.870 97.740 142.930 ;
        RECT 97.895 142.885 98.185 142.930 ;
        RECT 100.655 143.070 100.945 143.115 ;
        RECT 106.130 143.070 106.420 143.115 ;
        RECT 108.450 143.070 108.665 143.225 ;
        RECT 100.655 142.930 105.240 143.070 ;
        RECT 100.655 142.885 100.945 142.930 ;
        RECT 75.340 142.530 75.660 142.790 ;
        RECT 85.460 142.730 85.780 142.790 ;
        RECT 86.855 142.730 87.145 142.775 ;
        RECT 85.460 142.590 87.145 142.730 ;
        RECT 85.460 142.530 85.780 142.590 ;
        RECT 86.855 142.545 87.145 142.590 ;
        RECT 94.675 142.730 94.965 142.775 ;
        RECT 95.580 142.730 95.900 142.790 ;
        RECT 94.675 142.590 95.900 142.730 ;
        RECT 94.675 142.545 94.965 142.590 ;
        RECT 95.580 142.530 95.900 142.590 ;
        RECT 96.515 142.545 96.805 142.775 ;
        RECT 98.815 142.545 99.105 142.775 ;
        RECT 105.100 142.730 105.240 142.930 ;
        RECT 106.130 142.930 108.665 143.070 ;
        RECT 106.130 142.885 106.420 142.930 ;
        RECT 109.380 142.870 109.700 143.130 ;
        RECT 105.700 142.730 106.020 142.790 ;
        RECT 106.620 142.730 106.940 142.790 ;
        RECT 105.100 142.590 106.940 142.730 ;
        RECT 71.660 142.390 71.980 142.450 ;
        RECT 75.800 142.390 76.120 142.450 ;
        RECT 71.290 142.250 71.980 142.390 ;
        RECT 71.660 142.190 71.980 142.250 ;
        RECT 73.130 142.250 76.120 142.390 ;
        RECT 72.120 142.050 72.440 142.110 ;
        RECT 73.130 142.050 73.270 142.250 ;
        RECT 75.800 142.190 76.120 142.250 ;
        RECT 81.750 142.390 82.040 142.435 ;
        RECT 84.530 142.390 84.820 142.435 ;
        RECT 86.390 142.390 86.680 142.435 ;
        RECT 81.750 142.250 86.680 142.390 ;
        RECT 81.750 142.205 82.040 142.250 ;
        RECT 84.530 142.205 84.820 142.250 ;
        RECT 86.390 142.205 86.680 142.250 ;
        RECT 91.410 142.390 91.700 142.435 ;
        RECT 94.190 142.390 94.480 142.435 ;
        RECT 96.050 142.390 96.340 142.435 ;
        RECT 91.410 142.250 96.340 142.390 ;
        RECT 91.410 142.205 91.700 142.250 ;
        RECT 94.190 142.205 94.480 142.250 ;
        RECT 96.050 142.205 96.340 142.250 ;
        RECT 70.600 141.910 73.270 142.050 ;
        RECT 60.865 141.865 61.400 141.910 ;
        RECT 61.080 141.850 61.400 141.865 ;
        RECT 65.220 141.850 65.540 141.910 ;
        RECT 72.120 141.850 72.440 141.910 ;
        RECT 73.960 141.850 74.280 142.110 ;
        RECT 74.880 141.850 75.200 142.110 ;
        RECT 76.720 142.050 77.040 142.110 ;
        RECT 77.195 142.050 77.485 142.095 ;
        RECT 76.720 141.910 77.485 142.050 ;
        RECT 76.720 141.850 77.040 141.910 ;
        RECT 77.195 141.865 77.485 141.910 ;
        RECT 93.740 142.050 94.060 142.110 ;
        RECT 96.590 142.050 96.730 142.545 ;
        RECT 97.420 142.390 97.740 142.450 ;
        RECT 98.890 142.390 99.030 142.545 ;
        RECT 105.700 142.530 106.020 142.590 ;
        RECT 106.620 142.530 106.940 142.590 ;
        RECT 111.220 142.530 111.540 142.790 ;
        RECT 97.420 142.250 99.030 142.390 ;
        RECT 106.130 142.390 106.420 142.435 ;
        RECT 108.910 142.390 109.200 142.435 ;
        RECT 110.770 142.390 111.060 142.435 ;
        RECT 106.130 142.250 111.060 142.390 ;
        RECT 97.420 142.190 97.740 142.250 ;
        RECT 106.130 142.205 106.420 142.250 ;
        RECT 108.910 142.205 109.200 142.250 ;
        RECT 110.770 142.205 111.060 142.250 ;
        RECT 101.100 142.050 101.420 142.110 ;
        RECT 93.740 141.910 101.420 142.050 ;
        RECT 93.740 141.850 94.060 141.910 ;
        RECT 101.100 141.850 101.420 141.910 ;
        RECT 22.830 141.230 113.450 141.710 ;
        RECT 135.635 141.220 136.775 165.470 ;
        RECT 34.415 141.030 34.705 141.075 ;
        RECT 35.320 141.030 35.640 141.090 ;
        RECT 34.415 140.890 35.640 141.030 ;
        RECT 34.415 140.845 34.705 140.890 ;
        RECT 26.595 140.690 26.885 140.735 ;
        RECT 28.420 140.690 28.740 140.750 ;
        RECT 26.595 140.550 28.740 140.690 ;
        RECT 26.595 140.505 26.885 140.550 ;
        RECT 28.420 140.490 28.740 140.550 ;
        RECT 31.640 140.350 31.960 140.410 ;
        RECT 32.115 140.350 32.405 140.395 ;
        RECT 34.490 140.350 34.630 140.845 ;
        RECT 35.320 140.830 35.640 140.890 ;
        RECT 47.525 141.030 47.815 141.075 ;
        RECT 52.800 141.030 53.120 141.090 ;
        RECT 47.525 140.890 53.120 141.030 ;
        RECT 47.525 140.845 47.815 140.890 ;
        RECT 52.800 140.830 53.120 140.890 ;
        RECT 54.640 141.030 54.960 141.090 ;
        RECT 58.335 141.030 58.625 141.075 ;
        RECT 58.780 141.030 59.100 141.090 ;
        RECT 54.640 140.890 57.630 141.030 ;
        RECT 54.640 140.830 54.960 140.890 ;
        RECT 51.390 140.690 51.680 140.735 ;
        RECT 54.170 140.690 54.460 140.735 ;
        RECT 56.030 140.690 56.320 140.735 ;
        RECT 51.390 140.550 56.320 140.690 ;
        RECT 51.390 140.505 51.680 140.550 ;
        RECT 54.170 140.505 54.460 140.550 ;
        RECT 56.030 140.505 56.320 140.550 ;
        RECT 31.640 140.210 34.630 140.350 ;
        RECT 34.950 140.210 54.410 140.350 ;
        RECT 31.640 140.150 31.960 140.210 ;
        RECT 32.115 140.165 32.405 140.210 ;
        RECT 26.120 139.810 26.440 140.070 ;
        RECT 34.950 140.055 35.090 140.210 ;
        RECT 28.435 140.010 28.725 140.055 ;
        RECT 28.435 139.870 29.110 140.010 ;
        RECT 28.435 139.825 28.725 139.870 ;
        RECT 26.580 139.330 26.900 139.390 ;
        RECT 28.970 139.375 29.110 139.870 ;
        RECT 34.875 139.825 35.165 140.055 ;
        RECT 35.320 140.010 35.640 140.070 ;
        RECT 45.915 140.010 46.205 140.055 ;
        RECT 35.320 139.870 46.205 140.010 ;
        RECT 35.320 139.810 35.640 139.870 ;
        RECT 45.915 139.825 46.205 139.870 ;
        RECT 51.390 140.010 51.680 140.055 ;
        RECT 54.270 140.010 54.410 140.210 ;
        RECT 54.640 140.150 54.960 140.410 ;
        RECT 56.495 140.350 56.785 140.395 ;
        RECT 56.940 140.350 57.260 140.410 ;
        RECT 57.490 140.395 57.630 140.890 ;
        RECT 58.335 140.890 59.100 141.030 ;
        RECT 58.335 140.845 58.625 140.890 ;
        RECT 58.780 140.830 59.100 140.890 ;
        RECT 59.240 140.830 59.560 141.090 ;
        RECT 63.380 140.830 63.700 141.090 ;
        RECT 64.760 140.830 65.080 141.090 ;
        RECT 73.500 141.030 73.820 141.090 ;
        RECT 81.335 141.030 81.625 141.075 ;
        RECT 73.500 140.890 81.625 141.030 ;
        RECT 73.500 140.830 73.820 140.890 ;
        RECT 81.335 140.845 81.625 140.890 ;
        RECT 83.160 141.030 83.480 141.090 ;
        RECT 84.095 141.030 84.385 141.075 ;
        RECT 83.160 140.890 84.385 141.030 ;
        RECT 83.160 140.830 83.480 140.890 ;
        RECT 84.095 140.845 84.385 140.890 ;
        RECT 86.855 141.030 87.145 141.075 ;
        RECT 88.220 141.030 88.540 141.090 ;
        RECT 86.855 140.890 88.540 141.030 ;
        RECT 86.855 140.845 87.145 140.890 ;
        RECT 88.220 140.830 88.540 140.890 ;
        RECT 90.060 141.030 90.380 141.090 ;
        RECT 93.740 141.030 94.060 141.090 ;
        RECT 94.215 141.030 94.505 141.075 ;
        RECT 90.060 140.890 94.505 141.030 ;
        RECT 90.060 140.830 90.380 140.890 ;
        RECT 93.740 140.830 94.060 140.890 ;
        RECT 94.215 140.845 94.505 140.890 ;
        RECT 95.120 141.030 95.440 141.090 ;
        RECT 96.975 141.030 97.265 141.075 ;
        RECT 95.120 140.890 97.265 141.030 ;
        RECT 95.120 140.830 95.440 140.890 ;
        RECT 96.975 140.845 97.265 140.890 ;
        RECT 67.520 140.690 67.840 140.750 ;
        RECT 88.680 140.690 89.000 140.750 ;
        RECT 67.520 140.550 89.000 140.690 ;
        RECT 67.520 140.490 67.840 140.550 ;
        RECT 56.495 140.210 57.260 140.350 ;
        RECT 56.495 140.165 56.785 140.210 ;
        RECT 56.940 140.150 57.260 140.210 ;
        RECT 57.415 140.165 57.705 140.395 ;
        RECT 66.155 140.350 66.445 140.395 ;
        RECT 67.995 140.350 68.285 140.395 ;
        RECT 68.440 140.350 68.760 140.410 ;
        RECT 57.950 140.210 67.750 140.350 ;
        RECT 57.950 140.010 58.090 140.210 ;
        RECT 66.155 140.165 66.445 140.210 ;
        RECT 51.390 139.870 53.925 140.010 ;
        RECT 54.270 139.870 58.090 140.010 ;
        RECT 51.390 139.825 51.680 139.870 ;
        RECT 30.720 139.470 31.040 139.730 ;
        RECT 49.580 139.715 49.900 139.730 ;
        RECT 53.710 139.715 53.925 139.870 ;
        RECT 58.320 139.810 58.640 140.070 ;
        RECT 59.700 140.010 60.020 140.070 ;
        RECT 62.935 140.010 63.225 140.055 ;
        RECT 59.700 139.870 63.225 140.010 ;
        RECT 59.700 139.810 60.020 139.870 ;
        RECT 62.935 139.825 63.225 139.870 ;
        RECT 65.235 140.010 65.525 140.055 ;
        RECT 66.600 140.010 66.920 140.070 ;
        RECT 67.075 140.010 67.365 140.055 ;
        RECT 65.235 139.870 67.365 140.010 ;
        RECT 67.610 140.010 67.750 140.210 ;
        RECT 67.995 140.210 68.760 140.350 ;
        RECT 67.995 140.165 68.285 140.210 ;
        RECT 68.440 140.150 68.760 140.210 ;
        RECT 70.740 140.350 71.060 140.410 ;
        RECT 72.135 140.350 72.425 140.395 ;
        RECT 70.740 140.210 72.425 140.350 ;
        RECT 70.740 140.150 71.060 140.210 ;
        RECT 72.135 140.165 72.425 140.210 ;
        RECT 80.490 140.210 82.470 140.350 ;
        RECT 68.915 140.010 69.205 140.055 ;
        RECT 67.610 139.870 69.205 140.010 ;
        RECT 65.235 139.825 65.525 139.870 ;
        RECT 66.600 139.810 66.920 139.870 ;
        RECT 67.075 139.825 67.365 139.870 ;
        RECT 68.915 139.825 69.205 139.870 ;
        RECT 69.820 140.010 70.140 140.070 ;
        RECT 80.490 140.010 80.630 140.210 ;
        RECT 69.820 139.870 80.630 140.010 ;
        RECT 69.820 139.810 70.140 139.870 ;
        RECT 80.860 139.810 81.180 140.070 ;
        RECT 82.330 140.055 82.470 140.210 ;
        RECT 85.015 140.165 85.305 140.395 ;
        RECT 82.255 139.825 82.545 140.055 ;
        RECT 82.700 139.810 83.020 140.070 ;
        RECT 84.540 139.810 84.860 140.070 ;
        RECT 49.530 139.670 49.900 139.715 ;
        RECT 52.790 139.670 53.080 139.715 ;
        RECT 49.530 139.530 53.080 139.670 ;
        RECT 49.530 139.485 49.900 139.530 ;
        RECT 52.790 139.485 53.080 139.530 ;
        RECT 53.710 139.670 54.000 139.715 ;
        RECT 55.570 139.670 55.860 139.715 ;
        RECT 53.710 139.530 55.860 139.670 ;
        RECT 53.710 139.485 54.000 139.530 ;
        RECT 55.570 139.485 55.860 139.530 ;
        RECT 56.955 139.670 57.245 139.715 ;
        RECT 58.780 139.670 59.100 139.730 ;
        RECT 56.955 139.530 59.100 139.670 ;
        RECT 56.955 139.485 57.245 139.530 ;
        RECT 49.580 139.470 49.900 139.485 ;
        RECT 58.780 139.470 59.100 139.530 ;
        RECT 70.755 139.670 71.045 139.715 ;
        RECT 73.500 139.670 73.820 139.730 ;
        RECT 70.755 139.530 73.820 139.670 ;
        RECT 70.755 139.485 71.045 139.530 ;
        RECT 73.500 139.470 73.820 139.530 ;
        RECT 27.515 139.330 27.805 139.375 ;
        RECT 26.580 139.190 27.805 139.330 ;
        RECT 26.580 139.130 26.900 139.190 ;
        RECT 27.515 139.145 27.805 139.190 ;
        RECT 28.895 139.145 29.185 139.375 ;
        RECT 30.260 139.330 30.580 139.390 ;
        RECT 31.195 139.330 31.485 139.375 ;
        RECT 30.260 139.190 31.485 139.330 ;
        RECT 85.090 139.330 85.230 140.165 ;
        RECT 86.010 140.055 86.150 140.550 ;
        RECT 88.680 140.490 89.000 140.550 ;
        RECT 104.750 140.690 105.040 140.735 ;
        RECT 107.530 140.690 107.820 140.735 ;
        RECT 109.390 140.690 109.680 140.735 ;
        RECT 104.750 140.550 109.680 140.690 ;
        RECT 104.750 140.505 105.040 140.550 ;
        RECT 107.530 140.505 107.820 140.550 ;
        RECT 109.390 140.505 109.680 140.550 ;
        RECT 101.100 140.350 101.420 140.410 ;
        RECT 101.100 140.210 107.770 140.350 ;
        RECT 101.100 140.150 101.420 140.210 ;
        RECT 85.935 139.825 86.225 140.055 ;
        RECT 96.960 140.010 97.280 140.070 ;
        RECT 97.895 140.010 98.185 140.055 ;
        RECT 96.960 139.870 98.185 140.010 ;
        RECT 96.960 139.810 97.280 139.870 ;
        RECT 97.895 139.825 98.185 139.870 ;
        RECT 98.815 140.010 99.105 140.055 ;
        RECT 102.020 140.010 102.340 140.070 ;
        RECT 98.815 139.870 102.340 140.010 ;
        RECT 98.815 139.825 99.105 139.870 ;
        RECT 102.020 139.810 102.340 139.870 ;
        RECT 104.750 140.010 105.040 140.055 ;
        RECT 107.630 140.010 107.770 140.210 ;
        RECT 108.000 140.150 108.320 140.410 ;
        RECT 135.580 140.230 136.830 141.220 ;
        RECT 135.635 140.155 136.775 140.230 ;
        RECT 109.855 140.010 110.145 140.055 ;
        RECT 111.220 140.010 111.540 140.070 ;
        RECT 104.750 139.870 107.285 140.010 ;
        RECT 107.630 139.870 111.540 140.010 ;
        RECT 104.750 139.825 105.040 139.870 ;
        RECT 87.300 139.670 87.620 139.730 ;
        RECT 87.775 139.670 88.065 139.715 ;
        RECT 100.885 139.670 101.175 139.715 ;
        RECT 87.300 139.530 88.065 139.670 ;
        RECT 87.300 139.470 87.620 139.530 ;
        RECT 87.775 139.485 88.065 139.530 ;
        RECT 98.430 139.530 101.175 139.670 ;
        RECT 98.430 139.390 98.570 139.530 ;
        RECT 100.885 139.485 101.175 139.530 ;
        RECT 102.890 139.670 103.180 139.715 ;
        RECT 104.320 139.670 104.640 139.730 ;
        RECT 107.070 139.715 107.285 139.870 ;
        RECT 109.855 139.825 110.145 139.870 ;
        RECT 111.220 139.810 111.540 139.870 ;
        RECT 106.150 139.670 106.440 139.715 ;
        RECT 102.890 139.530 106.440 139.670 ;
        RECT 102.890 139.485 103.180 139.530 ;
        RECT 104.320 139.470 104.640 139.530 ;
        RECT 106.150 139.485 106.440 139.530 ;
        RECT 107.070 139.670 107.360 139.715 ;
        RECT 108.930 139.670 109.220 139.715 ;
        RECT 107.070 139.530 109.220 139.670 ;
        RECT 107.070 139.485 107.360 139.530 ;
        RECT 108.930 139.485 109.220 139.530 ;
        RECT 98.340 139.330 98.660 139.390 ;
        RECT 85.090 139.190 98.660 139.330 ;
        RECT 30.260 139.130 30.580 139.190 ;
        RECT 31.195 139.145 31.485 139.190 ;
        RECT 98.340 139.130 98.660 139.190 ;
        RECT 132.510 139.190 135.210 140.010 ;
        RECT 143.370 139.390 144.510 223.840 ;
        RECT 137.240 139.380 144.510 139.390 ;
        RECT 136.210 139.190 144.510 139.380 ;
        RECT 22.830 138.510 113.450 138.990 ;
        RECT 132.510 138.530 144.510 139.190 ;
        RECT 30.720 138.310 31.040 138.370 ;
        RECT 33.725 138.310 34.015 138.355 ;
        RECT 30.720 138.170 34.015 138.310 ;
        RECT 30.720 138.110 31.040 138.170 ;
        RECT 33.725 138.125 34.015 138.170 ;
        RECT 35.335 138.310 35.625 138.355 ;
        RECT 35.780 138.310 36.100 138.370 ;
        RECT 35.335 138.170 36.100 138.310 ;
        RECT 35.335 138.125 35.625 138.170 ;
        RECT 35.780 138.110 36.100 138.170 ;
        RECT 44.995 138.310 45.285 138.355 ;
        RECT 46.360 138.310 46.680 138.370 ;
        RECT 44.995 138.170 46.680 138.310 ;
        RECT 44.995 138.125 45.285 138.170 ;
        RECT 46.360 138.110 46.680 138.170 ;
        RECT 56.495 138.310 56.785 138.355 ;
        RECT 56.940 138.310 57.260 138.370 ;
        RECT 56.495 138.170 57.260 138.310 ;
        RECT 56.495 138.125 56.785 138.170 ;
        RECT 56.940 138.110 57.260 138.170 ;
        RECT 58.780 138.110 59.100 138.370 ;
        RECT 64.315 138.310 64.605 138.355 ;
        RECT 65.220 138.310 65.540 138.370 ;
        RECT 64.315 138.170 65.540 138.310 ;
        RECT 64.315 138.125 64.605 138.170 ;
        RECT 65.220 138.110 65.540 138.170 ;
        RECT 67.060 138.110 67.380 138.370 ;
        RECT 71.660 138.310 71.980 138.370 ;
        RECT 77.195 138.310 77.485 138.355 ;
        RECT 68.530 138.170 77.485 138.310 ;
        RECT 28.420 138.015 28.740 138.030 ;
        RECT 25.680 137.970 25.970 138.015 ;
        RECT 27.540 137.970 27.830 138.015 ;
        RECT 25.680 137.830 27.830 137.970 ;
        RECT 25.680 137.785 25.970 137.830 ;
        RECT 27.540 137.785 27.830 137.830 ;
        RECT 24.755 137.630 25.045 137.675 ;
        RECT 25.200 137.630 25.520 137.690 ;
        RECT 24.755 137.490 25.520 137.630 ;
        RECT 24.755 137.445 25.045 137.490 ;
        RECT 25.200 137.430 25.520 137.490 ;
        RECT 26.580 137.430 26.900 137.690 ;
        RECT 27.615 137.630 27.830 137.785 ;
        RECT 28.420 137.970 28.750 138.015 ;
        RECT 31.720 137.970 32.010 138.015 ;
        RECT 28.420 137.830 32.010 137.970 ;
        RECT 28.420 137.785 28.750 137.830 ;
        RECT 31.720 137.785 32.010 137.830 ;
        RECT 44.520 137.970 44.840 138.030 ;
        RECT 49.135 137.970 49.425 138.015 ;
        RECT 64.760 137.970 65.080 138.030 ;
        RECT 44.520 137.830 49.425 137.970 ;
        RECT 28.420 137.770 28.740 137.785 ;
        RECT 44.520 137.770 44.840 137.830 ;
        RECT 49.135 137.785 49.425 137.830 ;
        RECT 56.800 137.830 61.770 137.970 ;
        RECT 29.860 137.630 30.150 137.675 ;
        RECT 27.615 137.490 30.150 137.630 ;
        RECT 29.860 137.445 30.150 137.490 ;
        RECT 34.415 137.630 34.705 137.675 ;
        RECT 35.780 137.630 36.100 137.690 ;
        RECT 34.415 137.490 36.100 137.630 ;
        RECT 34.415 137.445 34.705 137.490 ;
        RECT 35.780 137.430 36.100 137.490 ;
        RECT 46.375 137.445 46.665 137.675 ;
        RECT 46.835 137.445 47.125 137.675 ;
        RECT 34.860 137.290 35.180 137.350 ;
        RECT 36.255 137.290 36.545 137.335 ;
        RECT 34.860 137.150 36.545 137.290 ;
        RECT 34.860 137.090 35.180 137.150 ;
        RECT 36.255 137.105 36.545 137.150 ;
        RECT 25.220 136.950 25.510 136.995 ;
        RECT 27.080 136.950 27.370 136.995 ;
        RECT 29.860 136.950 30.150 136.995 ;
        RECT 25.220 136.810 30.150 136.950 ;
        RECT 46.450 136.950 46.590 137.445 ;
        RECT 46.910 137.290 47.050 137.445 ;
        RECT 47.280 137.430 47.600 137.690 ;
        RECT 48.215 137.630 48.505 137.675 ;
        RECT 49.580 137.630 49.900 137.690 ;
        RECT 56.800 137.630 56.940 137.830 ;
        RECT 58.870 137.690 59.010 137.830 ;
        RECT 61.630 137.690 61.770 137.830 ;
        RECT 64.760 137.830 68.210 137.970 ;
        RECT 64.760 137.770 65.080 137.830 ;
        RECT 48.215 137.490 56.940 137.630 ;
        RECT 48.215 137.445 48.505 137.490 ;
        RECT 49.580 137.430 49.900 137.490 ;
        RECT 58.780 137.430 59.100 137.690 ;
        RECT 60.175 137.445 60.465 137.675 ;
        RECT 50.500 137.290 50.820 137.350 ;
        RECT 46.910 137.150 50.820 137.290 ;
        RECT 50.500 137.090 50.820 137.150 ;
        RECT 57.860 137.290 58.180 137.350 ;
        RECT 60.250 137.290 60.390 137.445 ;
        RECT 60.620 137.430 60.940 137.690 ;
        RECT 61.095 137.445 61.385 137.675 ;
        RECT 61.540 137.630 61.860 137.690 ;
        RECT 62.015 137.630 62.305 137.675 ;
        RECT 65.220 137.630 65.540 137.690 ;
        RECT 66.140 137.630 66.460 137.690 ;
        RECT 68.070 137.675 68.210 137.830 ;
        RECT 68.530 137.675 68.670 138.170 ;
        RECT 71.660 138.110 71.980 138.170 ;
        RECT 77.195 138.125 77.485 138.170 ;
        RECT 82.715 138.310 83.005 138.355 ;
        RECT 93.985 138.310 94.275 138.355 ;
        RECT 82.715 138.170 94.275 138.310 ;
        RECT 82.715 138.125 83.005 138.170 ;
        RECT 93.985 138.125 94.275 138.170 ;
        RECT 73.960 137.770 74.280 138.030 ;
        RECT 84.540 137.970 84.860 138.030 ;
        RECT 85.460 137.970 85.780 138.030 ;
        RECT 88.680 138.015 89.000 138.030 ;
        RECT 84.540 137.830 85.780 137.970 ;
        RECT 84.540 137.770 84.860 137.830 ;
        RECT 85.460 137.770 85.780 137.830 ;
        RECT 85.940 137.970 86.230 138.015 ;
        RECT 87.800 137.970 88.090 138.015 ;
        RECT 85.940 137.830 88.090 137.970 ;
        RECT 85.940 137.785 86.230 137.830 ;
        RECT 87.800 137.785 88.090 137.830 ;
        RECT 67.995 137.630 68.285 137.675 ;
        RECT 61.540 137.490 62.305 137.630 ;
        RECT 57.860 137.150 60.390 137.290 ;
        RECT 57.860 137.090 58.180 137.150 ;
        RECT 50.960 136.950 51.280 137.010 ;
        RECT 46.450 136.810 51.280 136.950 ;
        RECT 61.170 136.950 61.310 137.445 ;
        RECT 61.540 137.430 61.860 137.490 ;
        RECT 62.015 137.445 62.305 137.490 ;
        RECT 63.470 137.490 66.460 137.630 ;
        RECT 63.470 137.335 63.610 137.490 ;
        RECT 65.220 137.430 65.540 137.490 ;
        RECT 66.140 137.430 66.460 137.490 ;
        RECT 67.610 137.490 68.285 137.630 ;
        RECT 67.610 137.350 67.750 137.490 ;
        RECT 67.995 137.445 68.285 137.490 ;
        RECT 68.455 137.445 68.745 137.675 ;
        RECT 69.820 137.630 70.140 137.690 ;
        RECT 70.295 137.630 70.585 137.675 ;
        RECT 68.990 137.490 70.585 137.630 ;
        RECT 63.395 137.105 63.685 137.335 ;
        RECT 63.855 137.290 64.145 137.335 ;
        RECT 64.760 137.290 65.080 137.350 ;
        RECT 63.855 137.150 65.080 137.290 ;
        RECT 63.855 137.105 64.145 137.150 ;
        RECT 63.930 136.950 64.070 137.105 ;
        RECT 64.760 137.090 65.080 137.150 ;
        RECT 67.520 137.290 67.840 137.350 ;
        RECT 68.990 137.290 69.130 137.490 ;
        RECT 69.820 137.430 70.140 137.490 ;
        RECT 70.295 137.445 70.585 137.490 ;
        RECT 72.580 137.430 72.900 137.690 ;
        RECT 73.040 137.430 73.360 137.690 ;
        RECT 76.260 137.630 76.580 137.690 ;
        RECT 77.655 137.630 77.945 137.675 ;
        RECT 82.255 137.630 82.545 137.675 ;
        RECT 82.700 137.630 83.020 137.690 ;
        RECT 76.260 137.490 83.020 137.630 ;
        RECT 87.875 137.630 88.090 137.785 ;
        RECT 88.680 137.970 89.010 138.015 ;
        RECT 91.980 137.970 92.270 138.015 ;
        RECT 88.680 137.830 92.270 137.970 ;
        RECT 94.060 137.970 94.200 138.125 ;
        RECT 95.580 138.110 95.900 138.370 ;
        RECT 97.895 138.310 98.185 138.355 ;
        RECT 98.340 138.310 98.660 138.370 ;
        RECT 97.895 138.170 98.660 138.310 ;
        RECT 97.895 138.125 98.185 138.170 ;
        RECT 98.340 138.110 98.660 138.170 ;
        RECT 99.735 138.125 100.025 138.355 ;
        RECT 107.095 138.310 107.385 138.355 ;
        RECT 108.000 138.310 108.320 138.370 ;
        RECT 107.095 138.170 108.320 138.310 ;
        RECT 132.510 138.190 135.210 138.530 ;
        RECT 136.210 138.250 144.510 138.530 ;
        RECT 136.210 138.240 138.350 138.250 ;
        RECT 107.095 138.125 107.385 138.170 ;
        RECT 96.500 137.970 96.820 138.030 ;
        RECT 97.435 137.970 97.725 138.015 ;
        RECT 94.060 137.830 97.725 137.970 ;
        RECT 88.680 137.785 89.010 137.830 ;
        RECT 91.980 137.785 92.270 137.830 ;
        RECT 88.680 137.770 89.000 137.785 ;
        RECT 96.500 137.770 96.820 137.830 ;
        RECT 97.435 137.785 97.725 137.830 ;
        RECT 90.120 137.630 90.410 137.675 ;
        RECT 87.875 137.490 90.410 137.630 ;
        RECT 76.260 137.430 76.580 137.490 ;
        RECT 77.655 137.445 77.945 137.490 ;
        RECT 82.255 137.445 82.545 137.490 ;
        RECT 82.700 137.430 83.020 137.490 ;
        RECT 90.120 137.445 90.410 137.490 ;
        RECT 94.660 137.430 94.980 137.690 ;
        RECT 98.430 137.630 98.570 138.110 ;
        RECT 99.810 137.970 99.950 138.125 ;
        RECT 108.000 138.110 108.320 138.170 ;
        RECT 99.810 137.830 106.390 137.970 ;
        RECT 102.035 137.630 102.325 137.675 ;
        RECT 98.430 137.490 102.325 137.630 ;
        RECT 102.035 137.445 102.325 137.490 ;
        RECT 102.480 137.430 102.800 137.690 ;
        RECT 104.320 137.630 104.640 137.690 ;
        RECT 105.255 137.630 105.545 137.675 ;
        RECT 104.320 137.490 105.545 137.630 ;
        RECT 104.320 137.430 104.640 137.490 ;
        RECT 105.255 137.445 105.545 137.490 ;
        RECT 105.700 137.430 106.020 137.690 ;
        RECT 106.250 137.675 106.390 137.830 ;
        RECT 106.175 137.445 106.465 137.675 ;
        RECT 107.555 137.445 107.845 137.675 ;
        RECT 67.520 137.150 69.130 137.290 ;
        RECT 67.520 137.090 67.840 137.150 ;
        RECT 69.375 137.105 69.665 137.335 ;
        RECT 71.215 137.290 71.505 137.335 ;
        RECT 74.880 137.290 75.200 137.350 ;
        RECT 71.215 137.150 75.200 137.290 ;
        RECT 71.215 137.105 71.505 137.150 ;
        RECT 61.170 136.810 64.070 136.950 ;
        RECT 68.900 136.950 69.220 137.010 ;
        RECT 69.450 136.950 69.590 137.105 ;
        RECT 74.880 137.090 75.200 137.150 ;
        RECT 76.735 137.290 77.025 137.335 ;
        RECT 81.335 137.290 81.625 137.335 ;
        RECT 84.540 137.290 84.860 137.350 ;
        RECT 76.735 137.150 84.860 137.290 ;
        RECT 76.735 137.105 77.025 137.150 ;
        RECT 81.335 137.105 81.625 137.150 ;
        RECT 68.900 136.810 69.590 136.950 ;
        RECT 71.675 136.950 71.965 136.995 ;
        RECT 72.120 136.950 72.440 137.010 ;
        RECT 71.675 136.810 72.440 136.950 ;
        RECT 25.220 136.765 25.510 136.810 ;
        RECT 27.080 136.765 27.370 136.810 ;
        RECT 29.860 136.765 30.150 136.810 ;
        RECT 50.960 136.750 51.280 136.810 ;
        RECT 68.900 136.750 69.220 136.810 ;
        RECT 71.675 136.765 71.965 136.810 ;
        RECT 72.120 136.750 72.440 136.810 ;
        RECT 73.500 136.950 73.820 137.010 ;
        RECT 76.810 136.950 76.950 137.105 ;
        RECT 84.540 137.090 84.860 137.150 ;
        RECT 85.000 137.090 85.320 137.350 ;
        RECT 86.855 137.290 87.145 137.335 ;
        RECT 89.600 137.290 89.920 137.350 ;
        RECT 86.855 137.150 89.920 137.290 ;
        RECT 86.855 137.105 87.145 137.150 ;
        RECT 89.600 137.090 89.920 137.150 ;
        RECT 96.500 137.290 96.820 137.350 ;
        RECT 101.115 137.290 101.405 137.335 ;
        RECT 107.630 137.290 107.770 137.445 ;
        RECT 96.500 137.150 101.405 137.290 ;
        RECT 96.500 137.090 96.820 137.150 ;
        RECT 101.115 137.105 101.405 137.150 ;
        RECT 105.100 137.150 107.770 137.290 ;
        RECT 73.500 136.810 76.950 136.950 ;
        RECT 85.480 136.950 85.770 136.995 ;
        RECT 87.340 136.950 87.630 136.995 ;
        RECT 90.120 136.950 90.410 136.995 ;
        RECT 85.480 136.810 90.410 136.950 ;
        RECT 73.500 136.750 73.820 136.810 ;
        RECT 85.480 136.765 85.770 136.810 ;
        RECT 87.340 136.765 87.630 136.810 ;
        RECT 90.120 136.765 90.410 136.810 ;
        RECT 104.335 136.950 104.625 136.995 ;
        RECT 105.100 136.950 105.240 137.150 ;
        RECT 104.335 136.810 105.240 136.950 ;
        RECT 104.335 136.765 104.625 136.810 ;
        RECT 47.280 136.610 47.600 136.670 ;
        RECT 53.720 136.610 54.040 136.670 ;
        RECT 47.280 136.470 54.040 136.610 ;
        RECT 47.280 136.410 47.600 136.470 ;
        RECT 53.720 136.410 54.040 136.470 ;
        RECT 66.140 136.410 66.460 136.670 ;
        RECT 69.820 136.610 70.140 136.670 ;
        RECT 72.595 136.610 72.885 136.655 ;
        RECT 69.820 136.470 72.885 136.610 ;
        RECT 69.820 136.410 70.140 136.470 ;
        RECT 72.595 136.425 72.885 136.470 ;
        RECT 79.495 136.610 79.785 136.655 ;
        RECT 79.940 136.610 80.260 136.670 ;
        RECT 79.495 136.470 80.260 136.610 ;
        RECT 79.495 136.425 79.785 136.470 ;
        RECT 79.940 136.410 80.260 136.470 ;
        RECT 84.555 136.610 84.845 136.655 ;
        RECT 90.980 136.610 91.300 136.670 ;
        RECT 84.555 136.470 91.300 136.610 ;
        RECT 84.555 136.425 84.845 136.470 ;
        RECT 90.980 136.410 91.300 136.470 ;
        RECT 108.475 136.610 108.765 136.655 ;
        RECT 109.840 136.610 110.160 136.670 ;
        RECT 108.475 136.470 110.160 136.610 ;
        RECT 108.475 136.425 108.765 136.470 ;
        RECT 109.840 136.410 110.160 136.470 ;
        RECT 22.830 135.790 113.450 136.270 ;
        RECT 35.335 135.590 35.625 135.635 ;
        RECT 42.680 135.590 43.000 135.650 ;
        RECT 35.335 135.450 43.000 135.590 ;
        RECT 35.335 135.405 35.625 135.450 ;
        RECT 42.680 135.390 43.000 135.450 ;
        RECT 44.060 135.590 44.380 135.650 ;
        RECT 45.225 135.590 45.515 135.635 ;
        RECT 44.060 135.450 45.515 135.590 ;
        RECT 44.060 135.390 44.380 135.450 ;
        RECT 45.225 135.405 45.515 135.450 ;
        RECT 46.820 135.390 47.140 135.650 ;
        RECT 56.495 135.590 56.785 135.635 ;
        RECT 60.620 135.590 60.940 135.650 ;
        RECT 48.290 135.450 56.785 135.590 ;
        RECT 27.960 135.250 28.280 135.310 ;
        RECT 28.435 135.250 28.725 135.295 ;
        RECT 27.960 135.110 28.725 135.250 ;
        RECT 27.960 135.050 28.280 135.110 ;
        RECT 28.435 135.065 28.725 135.110 ;
        RECT 36.720 135.250 37.010 135.295 ;
        RECT 38.580 135.250 38.870 135.295 ;
        RECT 41.360 135.250 41.650 135.295 ;
        RECT 36.720 135.110 41.650 135.250 ;
        RECT 36.720 135.065 37.010 135.110 ;
        RECT 38.580 135.065 38.870 135.110 ;
        RECT 41.360 135.065 41.650 135.110 ;
        RECT 25.290 134.770 26.350 134.910 ;
        RECT 25.290 134.615 25.430 134.770 ;
        RECT 26.210 134.630 26.350 134.770 ;
        RECT 31.640 134.710 31.960 134.970 ;
        RECT 43.600 134.910 43.920 134.970 ;
        RECT 46.375 134.910 46.665 134.955 ;
        RECT 43.600 134.770 46.665 134.910 ;
        RECT 43.600 134.710 43.920 134.770 ;
        RECT 46.375 134.725 46.665 134.770 ;
        RECT 25.215 134.385 25.505 134.615 ;
        RECT 25.675 134.385 25.965 134.615 ;
        RECT 26.120 134.570 26.440 134.630 ;
        RECT 27.055 134.570 27.345 134.615 ;
        RECT 26.120 134.430 27.345 134.570 ;
        RECT 25.750 134.230 25.890 134.385 ;
        RECT 26.120 134.370 26.440 134.430 ;
        RECT 27.055 134.385 27.345 134.430 ;
        RECT 30.720 134.370 31.040 134.630 ;
        RECT 33.495 134.385 33.785 134.615 ;
        RECT 34.415 134.385 34.705 134.615 ;
        RECT 34.860 134.570 35.180 134.630 ;
        RECT 36.255 134.570 36.545 134.615 ;
        RECT 34.860 134.430 36.545 134.570 ;
        RECT 28.420 134.230 28.740 134.290 ;
        RECT 25.750 134.090 28.740 134.230 ;
        RECT 28.420 134.030 28.740 134.090 ;
        RECT 30.260 134.230 30.580 134.290 ;
        RECT 33.570 134.230 33.710 134.385 ;
        RECT 30.260 134.090 33.710 134.230 ;
        RECT 34.490 134.230 34.630 134.385 ;
        RECT 34.860 134.370 35.180 134.430 ;
        RECT 36.255 134.385 36.545 134.430 ;
        RECT 37.620 134.570 37.940 134.630 ;
        RECT 38.095 134.570 38.385 134.615 ;
        RECT 41.360 134.570 41.650 134.615 ;
        RECT 37.620 134.430 38.385 134.570 ;
        RECT 37.620 134.370 37.940 134.430 ;
        RECT 38.095 134.385 38.385 134.430 ;
        RECT 39.115 134.430 41.650 134.570 ;
        RECT 35.320 134.230 35.640 134.290 ;
        RECT 39.115 134.275 39.330 134.430 ;
        RECT 41.360 134.385 41.650 134.430 ;
        RECT 44.980 134.570 45.300 134.630 ;
        RECT 47.295 134.570 47.585 134.615 ;
        RECT 44.980 134.430 47.585 134.570 ;
        RECT 44.980 134.370 45.300 134.430 ;
        RECT 47.295 134.385 47.585 134.430 ;
        RECT 34.490 134.090 35.640 134.230 ;
        RECT 30.260 134.030 30.580 134.090 ;
        RECT 35.320 134.030 35.640 134.090 ;
        RECT 37.180 134.230 37.470 134.275 ;
        RECT 39.040 134.230 39.330 134.275 ;
        RECT 39.960 134.230 40.250 134.275 ;
        RECT 43.220 134.230 43.510 134.275 ;
        RECT 37.180 134.090 39.330 134.230 ;
        RECT 37.180 134.045 37.470 134.090 ;
        RECT 39.040 134.045 39.330 134.090 ;
        RECT 39.550 134.090 43.510 134.230 ;
        RECT 24.755 133.890 25.045 133.935 ;
        RECT 25.660 133.890 25.980 133.950 ;
        RECT 24.755 133.750 25.980 133.890 ;
        RECT 24.755 133.705 25.045 133.750 ;
        RECT 25.660 133.690 25.980 133.750 ;
        RECT 26.595 133.890 26.885 133.935 ;
        RECT 27.040 133.890 27.360 133.950 ;
        RECT 26.595 133.750 27.360 133.890 ;
        RECT 26.595 133.705 26.885 133.750 ;
        RECT 27.040 133.690 27.360 133.750 ;
        RECT 27.515 133.890 27.805 133.935 ;
        RECT 39.550 133.890 39.690 134.090 ;
        RECT 39.960 134.045 40.250 134.090 ;
        RECT 43.220 134.045 43.510 134.090 ;
        RECT 45.915 134.230 46.205 134.275 ;
        RECT 48.290 134.230 48.430 135.450 ;
        RECT 56.495 135.405 56.785 135.450 ;
        RECT 58.410 135.450 60.940 135.590 ;
        RECT 49.580 135.050 49.900 135.310 ;
        RECT 50.500 135.050 50.820 135.310 ;
        RECT 49.670 134.910 49.810 135.050 ;
        RECT 50.590 134.910 50.730 135.050 ;
        RECT 58.410 134.910 58.550 135.450 ;
        RECT 60.620 135.390 60.940 135.450 ;
        RECT 62.245 135.590 62.535 135.635 ;
        RECT 64.760 135.590 65.080 135.650 ;
        RECT 62.245 135.450 65.080 135.590 ;
        RECT 62.245 135.405 62.535 135.450 ;
        RECT 64.760 135.390 65.080 135.450 ;
        RECT 75.585 135.590 75.875 135.635 ;
        RECT 76.260 135.590 76.580 135.650 ;
        RECT 75.585 135.450 76.580 135.590 ;
        RECT 75.585 135.405 75.875 135.450 ;
        RECT 76.260 135.390 76.580 135.450 ;
        RECT 86.395 135.590 86.685 135.635 ;
        RECT 88.680 135.590 89.000 135.650 ;
        RECT 86.395 135.450 89.000 135.590 ;
        RECT 86.395 135.405 86.685 135.450 ;
        RECT 88.680 135.390 89.000 135.450 ;
        RECT 89.140 135.390 89.460 135.650 ;
        RECT 89.600 135.590 89.920 135.650 ;
        RECT 102.480 135.635 102.800 135.650 ;
        RECT 90.075 135.590 90.365 135.635 ;
        RECT 89.600 135.450 90.365 135.590 ;
        RECT 89.600 135.390 89.920 135.450 ;
        RECT 90.075 135.405 90.365 135.450 ;
        RECT 102.265 135.405 102.800 135.635 ;
        RECT 102.480 135.390 102.800 135.405 ;
        RECT 58.780 135.050 59.100 135.310 ;
        RECT 59.700 135.050 60.020 135.310 ;
        RECT 66.110 135.250 66.400 135.295 ;
        RECT 68.890 135.250 69.180 135.295 ;
        RECT 70.750 135.250 71.040 135.295 ;
        RECT 66.110 135.110 71.040 135.250 ;
        RECT 66.110 135.065 66.400 135.110 ;
        RECT 68.890 135.065 69.180 135.110 ;
        RECT 70.750 135.065 71.040 135.110 ;
        RECT 79.450 135.250 79.740 135.295 ;
        RECT 82.230 135.250 82.520 135.295 ;
        RECT 84.090 135.250 84.380 135.295 ;
        RECT 79.450 135.110 84.380 135.250 ;
        RECT 79.450 135.065 79.740 135.110 ;
        RECT 82.230 135.065 82.520 135.110 ;
        RECT 84.090 135.065 84.380 135.110 ;
        RECT 96.010 135.250 96.300 135.295 ;
        RECT 98.790 135.250 99.080 135.295 ;
        RECT 100.650 135.250 100.940 135.295 ;
        RECT 96.010 135.110 100.940 135.250 ;
        RECT 96.010 135.065 96.300 135.110 ;
        RECT 98.790 135.065 99.080 135.110 ;
        RECT 100.650 135.065 100.940 135.110 ;
        RECT 106.130 135.250 106.420 135.295 ;
        RECT 108.910 135.250 109.200 135.295 ;
        RECT 110.770 135.250 111.060 135.295 ;
        RECT 106.130 135.110 111.060 135.250 ;
        RECT 106.130 135.065 106.420 135.110 ;
        RECT 108.910 135.065 109.200 135.110 ;
        RECT 110.770 135.065 111.060 135.110 ;
        RECT 48.750 134.770 49.810 134.910 ;
        RECT 50.130 134.770 58.550 134.910 ;
        RECT 58.870 134.910 59.010 135.050 ;
        RECT 59.790 134.910 59.930 135.050 ;
        RECT 60.620 134.910 60.940 134.970 ;
        RECT 58.870 134.770 59.470 134.910 ;
        RECT 59.790 134.770 60.940 134.910 ;
        RECT 48.750 134.615 48.890 134.770 ;
        RECT 50.130 134.615 50.270 134.770 ;
        RECT 48.675 134.385 48.965 134.615 ;
        RECT 49.595 134.385 49.885 134.615 ;
        RECT 50.055 134.385 50.345 134.615 ;
        RECT 50.515 134.570 50.805 134.615 ;
        RECT 50.960 134.570 51.280 134.630 ;
        RECT 50.515 134.430 51.280 134.570 ;
        RECT 50.515 134.385 50.805 134.430 ;
        RECT 45.915 134.090 48.430 134.230 ;
        RECT 45.915 134.045 46.205 134.090 ;
        RECT 27.515 133.750 39.690 133.890 ;
        RECT 46.360 133.890 46.680 133.950 ;
        RECT 48.215 133.890 48.505 133.935 ;
        RECT 46.360 133.750 48.505 133.890 ;
        RECT 49.670 133.890 49.810 134.385 ;
        RECT 50.960 134.370 51.280 134.430 ;
        RECT 55.575 134.570 55.865 134.615 ;
        RECT 56.940 134.570 57.260 134.630 ;
        RECT 55.575 134.430 57.260 134.570 ;
        RECT 55.575 134.385 55.865 134.430 ;
        RECT 56.940 134.370 57.260 134.430 ;
        RECT 57.860 134.370 58.180 134.630 ;
        RECT 58.410 134.615 58.550 134.770 ;
        RECT 58.335 134.385 58.625 134.615 ;
        RECT 58.795 134.385 59.085 134.615 ;
        RECT 59.330 134.570 59.470 134.770 ;
        RECT 60.250 134.615 60.390 134.770 ;
        RECT 60.620 134.710 60.940 134.770 ;
        RECT 72.670 134.770 82.470 134.910 ;
        RECT 59.715 134.570 60.005 134.615 ;
        RECT 59.330 134.430 60.005 134.570 ;
        RECT 59.715 134.385 60.005 134.430 ;
        RECT 60.175 134.385 60.465 134.615 ;
        RECT 66.110 134.570 66.400 134.615 ;
        RECT 66.110 134.430 68.645 134.570 ;
        RECT 66.110 134.385 66.400 134.430 ;
        RECT 51.050 134.230 51.190 134.370 ;
        RECT 57.950 134.230 58.090 134.370 ;
        RECT 51.050 134.090 58.090 134.230 ;
        RECT 58.870 134.230 59.010 134.385 ;
        RECT 68.430 134.275 68.645 134.430 ;
        RECT 69.360 134.370 69.680 134.630 ;
        RECT 70.740 134.570 71.060 134.630 ;
        RECT 72.670 134.615 72.810 134.770 ;
        RECT 71.215 134.570 71.505 134.615 ;
        RECT 72.595 134.570 72.885 134.615 ;
        RECT 70.740 134.430 72.885 134.570 ;
        RECT 70.740 134.370 71.060 134.430 ;
        RECT 71.215 134.385 71.505 134.430 ;
        RECT 72.595 134.385 72.885 134.430 ;
        RECT 79.450 134.570 79.740 134.615 ;
        RECT 82.330 134.570 82.470 134.770 ;
        RECT 82.700 134.710 83.020 134.970 ;
        RECT 91.900 134.955 92.220 134.970 ;
        RECT 91.900 134.910 92.435 134.955 ;
        RECT 97.420 134.910 97.740 134.970 ;
        RECT 91.900 134.770 97.740 134.910 ;
        RECT 91.900 134.725 92.435 134.770 ;
        RECT 91.900 134.710 92.220 134.725 ;
        RECT 97.420 134.710 97.740 134.770 ;
        RECT 101.100 134.710 101.420 134.970 ;
        RECT 109.395 134.910 109.685 134.955 ;
        RECT 109.840 134.910 110.160 134.970 ;
        RECT 109.395 134.770 110.160 134.910 ;
        RECT 109.395 134.725 109.685 134.770 ;
        RECT 109.840 134.710 110.160 134.770 ;
        RECT 111.220 134.710 111.540 134.970 ;
        RECT 84.555 134.570 84.845 134.615 ;
        RECT 85.000 134.570 85.320 134.630 ;
        RECT 79.450 134.430 81.985 134.570 ;
        RECT 82.330 134.430 85.320 134.570 ;
        RECT 79.450 134.385 79.740 134.430 ;
        RECT 60.635 134.230 60.925 134.275 ;
        RECT 64.250 134.230 64.540 134.275 ;
        RECT 67.510 134.230 67.800 134.275 ;
        RECT 58.870 134.090 59.930 134.230 ;
        RECT 59.790 133.950 59.930 134.090 ;
        RECT 60.635 134.090 67.800 134.230 ;
        RECT 60.635 134.045 60.925 134.090 ;
        RECT 64.250 134.045 64.540 134.090 ;
        RECT 67.510 134.045 67.800 134.090 ;
        RECT 68.430 134.230 68.720 134.275 ;
        RECT 70.290 134.230 70.580 134.275 ;
        RECT 68.430 134.090 70.580 134.230 ;
        RECT 68.430 134.045 68.720 134.090 ;
        RECT 70.290 134.045 70.580 134.090 ;
        RECT 74.420 134.230 74.740 134.290 ;
        RECT 81.770 134.275 81.985 134.430 ;
        RECT 84.555 134.385 84.845 134.430 ;
        RECT 85.000 134.370 85.320 134.430 ;
        RECT 85.460 134.570 85.780 134.630 ;
        RECT 85.935 134.570 86.225 134.615 ;
        RECT 88.680 134.570 89.000 134.630 ;
        RECT 85.460 134.430 89.000 134.570 ;
        RECT 85.460 134.370 85.780 134.430 ;
        RECT 85.935 134.385 86.225 134.430 ;
        RECT 88.680 134.370 89.000 134.430 ;
        RECT 90.980 134.370 91.300 134.630 ;
        RECT 96.010 134.570 96.300 134.615 ;
        RECT 96.010 134.430 98.545 134.570 ;
        RECT 96.010 134.385 96.300 134.430 ;
        RECT 77.590 134.230 77.880 134.275 ;
        RECT 80.850 134.230 81.140 134.275 ;
        RECT 74.420 134.090 81.140 134.230 ;
        RECT 74.420 134.030 74.740 134.090 ;
        RECT 77.590 134.045 77.880 134.090 ;
        RECT 80.850 134.045 81.140 134.090 ;
        RECT 81.770 134.230 82.060 134.275 ;
        RECT 83.630 134.230 83.920 134.275 ;
        RECT 81.770 134.090 83.920 134.230 ;
        RECT 81.770 134.045 82.060 134.090 ;
        RECT 83.630 134.045 83.920 134.090 ;
        RECT 94.150 134.230 94.440 134.275 ;
        RECT 95.120 134.230 95.440 134.290 ;
        RECT 98.330 134.275 98.545 134.430 ;
        RECT 99.260 134.370 99.580 134.630 ;
        RECT 106.130 134.570 106.420 134.615 ;
        RECT 106.130 134.430 108.665 134.570 ;
        RECT 135.660 134.480 136.800 134.510 ;
        RECT 106.130 134.385 106.420 134.430 ;
        RECT 97.410 134.230 97.700 134.275 ;
        RECT 94.150 134.090 97.700 134.230 ;
        RECT 94.150 134.045 94.440 134.090 ;
        RECT 95.120 134.030 95.440 134.090 ;
        RECT 97.410 134.045 97.700 134.090 ;
        RECT 98.330 134.230 98.620 134.275 ;
        RECT 100.190 134.230 100.480 134.275 ;
        RECT 98.330 134.090 100.480 134.230 ;
        RECT 98.330 134.045 98.620 134.090 ;
        RECT 100.190 134.045 100.480 134.090 ;
        RECT 104.270 134.230 104.560 134.275 ;
        RECT 105.700 134.230 106.020 134.290 ;
        RECT 108.450 134.275 108.665 134.430 ;
        RECT 107.530 134.230 107.820 134.275 ;
        RECT 104.270 134.090 107.820 134.230 ;
        RECT 104.270 134.045 104.560 134.090 ;
        RECT 105.700 134.030 106.020 134.090 ;
        RECT 107.530 134.045 107.820 134.090 ;
        RECT 108.450 134.230 108.740 134.275 ;
        RECT 110.310 134.230 110.600 134.275 ;
        RECT 108.450 134.090 110.600 134.230 ;
        RECT 108.450 134.045 108.740 134.090 ;
        RECT 110.310 134.045 110.600 134.090 ;
        RECT 50.960 133.890 51.280 133.950 ;
        RECT 49.670 133.750 51.280 133.890 ;
        RECT 27.515 133.705 27.805 133.750 ;
        RECT 46.360 133.690 46.680 133.750 ;
        RECT 48.215 133.705 48.505 133.750 ;
        RECT 50.960 133.690 51.280 133.750 ;
        RECT 51.420 133.890 51.740 133.950 ;
        RECT 51.895 133.890 52.185 133.935 ;
        RECT 51.420 133.750 52.185 133.890 ;
        RECT 51.420 133.690 51.740 133.750 ;
        RECT 51.895 133.705 52.185 133.750 ;
        RECT 59.700 133.690 60.020 133.950 ;
        RECT 22.830 133.070 113.450 133.550 ;
        RECT 135.590 133.400 136.850 134.480 ;
        RECT 37.160 132.870 37.480 132.930 ;
        RECT 38.095 132.870 38.385 132.915 ;
        RECT 37.160 132.730 38.385 132.870 ;
        RECT 37.160 132.670 37.480 132.730 ;
        RECT 38.095 132.685 38.385 132.730 ;
        RECT 42.695 132.685 42.985 132.915 ;
        RECT 25.660 132.530 25.980 132.590 ;
        RECT 26.530 132.530 26.820 132.575 ;
        RECT 29.790 132.530 30.080 132.575 ;
        RECT 25.660 132.390 30.080 132.530 ;
        RECT 25.660 132.330 25.980 132.390 ;
        RECT 26.530 132.345 26.820 132.390 ;
        RECT 29.790 132.345 30.080 132.390 ;
        RECT 30.710 132.530 31.000 132.575 ;
        RECT 32.570 132.530 32.860 132.575 ;
        RECT 30.710 132.390 32.860 132.530 ;
        RECT 30.710 132.345 31.000 132.390 ;
        RECT 32.570 132.345 32.860 132.390 ;
        RECT 38.540 132.530 38.860 132.590 ;
        RECT 42.770 132.530 42.910 132.685 ;
        RECT 44.520 132.670 44.840 132.930 ;
        RECT 49.135 132.870 49.425 132.915 ;
        RECT 49.580 132.870 49.900 132.930 ;
        RECT 49.135 132.730 49.900 132.870 ;
        RECT 49.135 132.685 49.425 132.730 ;
        RECT 49.580 132.670 49.900 132.730 ;
        RECT 50.960 132.870 51.280 132.930 ;
        RECT 52.815 132.870 53.105 132.915 ;
        RECT 54.180 132.870 54.500 132.930 ;
        RECT 50.960 132.730 52.570 132.870 ;
        RECT 50.960 132.670 51.280 132.730 ;
        RECT 44.060 132.530 44.380 132.590 ;
        RECT 44.995 132.530 45.285 132.575 ;
        RECT 47.295 132.530 47.585 132.575 ;
        RECT 38.540 132.390 42.910 132.530 ;
        RECT 43.690 132.390 45.285 132.530 ;
        RECT 28.390 132.190 28.680 132.235 ;
        RECT 30.710 132.190 30.925 132.345 ;
        RECT 38.540 132.330 38.860 132.390 ;
        RECT 28.390 132.050 30.925 132.190 ;
        RECT 28.390 132.005 28.680 132.050 ;
        RECT 31.640 131.990 31.960 132.250 ;
        RECT 32.100 132.190 32.420 132.250 ;
        RECT 36.240 132.190 36.560 132.250 ;
        RECT 39.920 132.190 40.240 132.250 ;
        RECT 32.100 132.050 35.550 132.190 ;
        RECT 32.100 131.990 32.420 132.050 ;
        RECT 25.200 131.850 25.520 131.910 ;
        RECT 33.495 131.850 33.785 131.895 ;
        RECT 34.860 131.850 35.180 131.910 ;
        RECT 35.410 131.895 35.550 132.050 ;
        RECT 36.240 132.050 40.240 132.190 ;
        RECT 36.240 131.990 36.560 132.050 ;
        RECT 39.920 131.990 40.240 132.050 ;
        RECT 40.395 132.190 40.685 132.235 ;
        RECT 43.690 132.190 43.830 132.390 ;
        RECT 44.060 132.330 44.380 132.390 ;
        RECT 44.995 132.345 45.285 132.390 ;
        RECT 45.530 132.390 47.585 132.530 ;
        RECT 45.530 132.190 45.670 132.390 ;
        RECT 47.295 132.345 47.585 132.390 ;
        RECT 51.420 132.330 51.740 132.590 ;
        RECT 52.430 132.530 52.570 132.730 ;
        RECT 52.815 132.730 54.500 132.870 ;
        RECT 52.815 132.685 53.105 132.730 ;
        RECT 54.180 132.670 54.500 132.730 ;
        RECT 56.940 132.670 57.260 132.930 ;
        RECT 63.855 132.870 64.145 132.915 ;
        RECT 64.760 132.870 65.080 132.930 ;
        RECT 63.855 132.730 65.080 132.870 ;
        RECT 63.855 132.685 64.145 132.730 ;
        RECT 64.760 132.670 65.080 132.730 ;
        RECT 67.535 132.870 67.825 132.915 ;
        RECT 69.360 132.870 69.680 132.930 ;
        RECT 67.535 132.730 69.680 132.870 ;
        RECT 67.535 132.685 67.825 132.730 ;
        RECT 69.360 132.670 69.680 132.730 ;
        RECT 69.820 132.670 70.140 132.930 ;
        RECT 71.660 132.870 71.980 132.930 ;
        RECT 72.135 132.870 72.425 132.915 ;
        RECT 71.660 132.730 72.425 132.870 ;
        RECT 71.660 132.670 71.980 132.730 ;
        RECT 72.135 132.685 72.425 132.730 ;
        RECT 73.975 132.685 74.265 132.915 ;
        RECT 55.115 132.530 55.405 132.575 ;
        RECT 58.795 132.530 59.085 132.575 ;
        RECT 52.430 132.390 59.085 132.530 ;
        RECT 55.115 132.345 55.405 132.390 ;
        RECT 58.795 132.345 59.085 132.390 ;
        RECT 40.395 132.050 43.830 132.190 ;
        RECT 44.150 132.050 45.670 132.190 ;
        RECT 40.395 132.005 40.685 132.050 ;
        RECT 25.200 131.710 35.180 131.850 ;
        RECT 25.200 131.650 25.520 131.710 ;
        RECT 33.495 131.665 33.785 131.710 ;
        RECT 34.860 131.650 35.180 131.710 ;
        RECT 35.335 131.665 35.625 131.895 ;
        RECT 35.795 131.850 36.085 131.895 ;
        RECT 35.795 131.710 40.610 131.850 ;
        RECT 35.795 131.665 36.085 131.710 ;
        RECT 28.390 131.510 28.680 131.555 ;
        RECT 31.170 131.510 31.460 131.555 ;
        RECT 33.030 131.510 33.320 131.555 ;
        RECT 28.390 131.370 33.320 131.510 ;
        RECT 35.410 131.510 35.550 131.665 ;
        RECT 40.470 131.570 40.610 131.710 ;
        RECT 40.840 131.650 41.160 131.910 ;
        RECT 41.315 131.665 41.605 131.895 ;
        RECT 43.600 131.850 43.920 131.910 ;
        RECT 44.150 131.850 44.290 132.050 ;
        RECT 46.835 132.005 47.125 132.235 ;
        RECT 45.455 131.850 45.745 131.895 ;
        RECT 43.600 131.710 44.290 131.850 ;
        RECT 44.610 131.710 45.745 131.850 ;
        RECT 46.910 131.850 47.050 132.005 ;
        RECT 50.040 131.990 50.360 132.250 ;
        RECT 51.880 131.990 52.200 132.250 ;
        RECT 53.720 132.190 54.040 132.250 ;
        RECT 54.655 132.190 54.945 132.235 ;
        RECT 53.720 132.050 54.945 132.190 ;
        RECT 53.720 131.990 54.040 132.050 ;
        RECT 54.655 132.005 54.945 132.050 ;
        RECT 59.255 132.190 59.545 132.235 ;
        RECT 59.700 132.190 60.020 132.250 ;
        RECT 66.140 132.190 66.460 132.250 ;
        RECT 66.615 132.190 66.905 132.235 ;
        RECT 59.255 132.050 63.610 132.190 ;
        RECT 59.255 132.005 59.545 132.050 ;
        RECT 59.700 131.990 60.020 132.050 ;
        RECT 63.470 131.910 63.610 132.050 ;
        RECT 66.140 132.050 66.905 132.190 ;
        RECT 66.140 131.990 66.460 132.050 ;
        RECT 66.615 132.005 66.905 132.050 ;
        RECT 67.520 132.190 67.840 132.250 ;
        RECT 68.915 132.190 69.205 132.235 ;
        RECT 73.500 132.190 73.820 132.250 ;
        RECT 67.520 132.050 69.205 132.190 ;
        RECT 67.520 131.990 67.840 132.050 ;
        RECT 68.915 132.005 69.205 132.050 ;
        RECT 71.290 132.050 73.820 132.190 ;
        RECT 74.050 132.190 74.190 132.685 ;
        RECT 79.020 132.670 79.340 132.930 ;
        RECT 81.795 132.870 82.085 132.915 ;
        RECT 82.700 132.870 83.020 132.930 ;
        RECT 81.795 132.730 83.020 132.870 ;
        RECT 81.795 132.685 82.085 132.730 ;
        RECT 82.700 132.670 83.020 132.730 ;
        RECT 88.680 132.870 89.000 132.930 ;
        RECT 88.680 132.730 94.890 132.870 ;
        RECT 88.680 132.670 89.000 132.730 ;
        RECT 76.260 132.530 76.580 132.590 ;
        RECT 77.195 132.530 77.485 132.575 ;
        RECT 76.260 132.390 77.485 132.530 ;
        RECT 76.260 132.330 76.580 132.390 ;
        RECT 77.195 132.345 77.485 132.390 ;
        RECT 79.940 132.530 80.260 132.590 ;
        RECT 87.250 132.530 87.540 132.575 ;
        RECT 88.220 132.530 88.540 132.590 ;
        RECT 90.510 132.530 90.800 132.575 ;
        RECT 79.940 132.390 81.090 132.530 ;
        RECT 79.940 132.330 80.260 132.390 ;
        RECT 80.950 132.235 81.090 132.390 ;
        RECT 87.250 132.390 90.800 132.530 ;
        RECT 87.250 132.345 87.540 132.390 ;
        RECT 88.220 132.330 88.540 132.390 ;
        RECT 90.510 132.345 90.800 132.390 ;
        RECT 91.430 132.530 91.720 132.575 ;
        RECT 93.290 132.530 93.580 132.575 ;
        RECT 91.430 132.390 93.580 132.530 ;
        RECT 91.430 132.345 91.720 132.390 ;
        RECT 93.290 132.345 93.580 132.390 ;
        RECT 94.750 132.530 94.890 132.730 ;
        RECT 95.120 132.670 95.440 132.930 ;
        RECT 97.420 132.870 97.740 132.930 ;
        RECT 97.895 132.870 98.185 132.915 ;
        RECT 97.420 132.730 98.185 132.870 ;
        RECT 97.420 132.670 97.740 132.730 ;
        RECT 97.895 132.685 98.185 132.730 ;
        RECT 101.100 132.530 101.420 132.590 ;
        RECT 102.890 132.530 103.180 132.575 ;
        RECT 104.320 132.530 104.640 132.590 ;
        RECT 106.150 132.530 106.440 132.575 ;
        RECT 94.750 132.390 98.110 132.530 ;
        RECT 80.415 132.190 80.705 132.235 ;
        RECT 74.050 132.050 80.705 132.190 ;
        RECT 47.280 131.850 47.600 131.910 ;
        RECT 46.910 131.710 47.600 131.850 ;
        RECT 35.410 131.370 40.150 131.510 ;
        RECT 28.390 131.325 28.680 131.370 ;
        RECT 31.170 131.325 31.460 131.370 ;
        RECT 33.030 131.325 33.320 131.370 ;
        RECT 24.525 131.170 24.815 131.215 ;
        RECT 30.260 131.170 30.580 131.230 ;
        RECT 24.525 131.030 30.580 131.170 ;
        RECT 24.525 130.985 24.815 131.030 ;
        RECT 30.260 130.970 30.580 131.030 ;
        RECT 38.080 131.170 38.400 131.230 ;
        RECT 38.555 131.170 38.845 131.215 ;
        RECT 38.080 131.030 38.845 131.170 ;
        RECT 40.010 131.170 40.150 131.370 ;
        RECT 40.380 131.310 40.700 131.570 ;
        RECT 41.390 131.510 41.530 131.665 ;
        RECT 43.600 131.650 43.920 131.710 ;
        RECT 44.610 131.510 44.750 131.710 ;
        RECT 45.455 131.665 45.745 131.710 ;
        RECT 47.280 131.650 47.600 131.710 ;
        RECT 50.975 131.665 51.265 131.895 ;
        RECT 54.195 131.850 54.485 131.895 ;
        RECT 58.335 131.850 58.625 131.895 ;
        RECT 62.935 131.850 63.225 131.895 ;
        RECT 54.195 131.710 63.225 131.850 ;
        RECT 54.195 131.665 54.485 131.710 ;
        RECT 58.335 131.665 58.625 131.710 ;
        RECT 62.935 131.665 63.225 131.710 ;
        RECT 41.390 131.370 44.750 131.510 ;
        RECT 51.050 131.510 51.190 131.665 ;
        RECT 55.560 131.510 55.880 131.570 ;
        RECT 51.050 131.370 55.880 131.510 ;
        RECT 63.010 131.510 63.150 131.665 ;
        RECT 63.380 131.650 63.700 131.910 ;
        RECT 71.290 131.895 71.430 132.050 ;
        RECT 73.500 131.990 73.820 132.050 ;
        RECT 80.415 132.005 80.705 132.050 ;
        RECT 80.875 132.005 81.165 132.235 ;
        RECT 83.635 132.005 83.925 132.235 ;
        RECT 84.095 132.190 84.385 132.235 ;
        RECT 85.460 132.190 85.780 132.250 ;
        RECT 84.095 132.050 85.780 132.190 ;
        RECT 84.095 132.005 84.385 132.050 ;
        RECT 67.995 131.665 68.285 131.895 ;
        RECT 71.215 131.665 71.505 131.895 ;
        RECT 71.675 131.850 71.965 131.895 ;
        RECT 75.800 131.850 76.120 131.910 ;
        RECT 71.675 131.710 76.120 131.850 ;
        RECT 71.675 131.665 71.965 131.710 ;
        RECT 65.220 131.510 65.540 131.570 ;
        RECT 63.010 131.370 65.540 131.510 ;
        RECT 68.070 131.510 68.210 131.665 ;
        RECT 71.750 131.510 71.890 131.665 ;
        RECT 75.800 131.650 76.120 131.710 ;
        RECT 76.275 131.665 76.565 131.895 ;
        RECT 76.735 131.665 77.025 131.895 ;
        RECT 81.320 131.850 81.640 131.910 ;
        RECT 83.710 131.850 83.850 132.005 ;
        RECT 85.460 131.990 85.780 132.050 ;
        RECT 89.110 132.190 89.400 132.235 ;
        RECT 91.430 132.190 91.645 132.345 ;
        RECT 94.750 132.235 94.890 132.390 ;
        RECT 89.110 132.050 91.645 132.190 ;
        RECT 89.110 132.005 89.400 132.050 ;
        RECT 94.675 132.005 94.965 132.235 ;
        RECT 97.970 132.190 98.110 132.390 ;
        RECT 101.100 132.390 102.250 132.530 ;
        RECT 101.100 132.330 101.420 132.390 ;
        RECT 97.970 132.050 101.790 132.190 ;
        RECT 81.320 131.710 83.850 131.850 ;
        RECT 68.070 131.370 71.890 131.510 ;
        RECT 73.500 131.510 73.820 131.570 ;
        RECT 76.350 131.510 76.490 131.665 ;
        RECT 73.500 131.370 76.490 131.510 ;
        RECT 76.810 131.510 76.950 131.665 ;
        RECT 81.320 131.650 81.640 131.710 ;
        RECT 92.360 131.650 92.680 131.910 ;
        RECT 94.200 131.650 94.520 131.910 ;
        RECT 96.500 131.850 96.820 131.910 ;
        RECT 96.130 131.710 96.820 131.850 ;
        RECT 83.620 131.510 83.940 131.570 ;
        RECT 76.810 131.370 83.940 131.510 ;
        RECT 41.390 131.170 41.530 131.370 ;
        RECT 55.560 131.310 55.880 131.370 ;
        RECT 65.220 131.310 65.540 131.370 ;
        RECT 73.500 131.310 73.820 131.370 ;
        RECT 40.010 131.030 41.530 131.170 ;
        RECT 38.080 130.970 38.400 131.030 ;
        RECT 38.555 130.985 38.845 131.030 ;
        RECT 50.040 130.970 50.360 131.230 ;
        RECT 61.095 131.170 61.385 131.215 ;
        RECT 61.540 131.170 61.860 131.230 ;
        RECT 61.095 131.030 61.860 131.170 ;
        RECT 61.095 130.985 61.385 131.030 ;
        RECT 61.540 130.970 61.860 131.030 ;
        RECT 65.695 131.170 65.985 131.215 ;
        RECT 66.140 131.170 66.460 131.230 ;
        RECT 65.695 131.030 66.460 131.170 ;
        RECT 65.695 130.985 65.985 131.030 ;
        RECT 66.140 130.970 66.460 131.030 ;
        RECT 68.900 131.170 69.220 131.230 ;
        RECT 76.810 131.170 76.950 131.370 ;
        RECT 83.620 131.310 83.940 131.370 ;
        RECT 84.540 131.510 84.860 131.570 ;
        RECT 85.245 131.510 85.535 131.555 ;
        RECT 87.760 131.510 88.080 131.570 ;
        RECT 84.540 131.370 88.080 131.510 ;
        RECT 84.540 131.310 84.860 131.370 ;
        RECT 85.245 131.325 85.535 131.370 ;
        RECT 87.760 131.310 88.080 131.370 ;
        RECT 89.110 131.510 89.400 131.555 ;
        RECT 91.890 131.510 92.180 131.555 ;
        RECT 93.750 131.510 94.040 131.555 ;
        RECT 89.110 131.370 94.040 131.510 ;
        RECT 89.110 131.325 89.400 131.370 ;
        RECT 91.890 131.325 92.180 131.370 ;
        RECT 93.750 131.325 94.040 131.370 ;
        RECT 68.900 131.030 76.950 131.170 ;
        RECT 79.495 131.170 79.785 131.215 ;
        RECT 79.940 131.170 80.260 131.230 ;
        RECT 79.495 131.030 80.260 131.170 ;
        RECT 68.900 130.970 69.220 131.030 ;
        RECT 79.495 130.985 79.785 131.030 ;
        RECT 79.940 130.970 80.260 131.030 ;
        RECT 90.980 131.170 91.300 131.230 ;
        RECT 96.130 131.170 96.270 131.710 ;
        RECT 96.500 131.650 96.820 131.710 ;
        RECT 97.435 131.850 97.725 131.895 ;
        RECT 98.800 131.850 99.120 131.910 ;
        RECT 100.885 131.850 101.175 131.895 ;
        RECT 97.435 131.710 101.175 131.850 ;
        RECT 97.435 131.665 97.725 131.710 ;
        RECT 98.800 131.650 99.120 131.710 ;
        RECT 100.885 131.665 101.175 131.710 ;
        RECT 90.980 131.030 96.270 131.170 ;
        RECT 98.340 131.170 98.660 131.230 ;
        RECT 99.735 131.170 100.025 131.215 ;
        RECT 98.340 131.030 100.025 131.170 ;
        RECT 101.650 131.170 101.790 132.050 ;
        RECT 102.110 131.850 102.250 132.390 ;
        RECT 102.890 132.390 106.440 132.530 ;
        RECT 102.890 132.345 103.180 132.390 ;
        RECT 104.320 132.330 104.640 132.390 ;
        RECT 106.150 132.345 106.440 132.390 ;
        RECT 107.070 132.530 107.360 132.575 ;
        RECT 108.930 132.530 109.220 132.575 ;
        RECT 107.070 132.390 109.220 132.530 ;
        RECT 107.070 132.345 107.360 132.390 ;
        RECT 108.930 132.345 109.220 132.390 ;
        RECT 104.750 132.190 105.040 132.235 ;
        RECT 107.070 132.190 107.285 132.345 ;
        RECT 104.750 132.050 107.285 132.190 ;
        RECT 107.540 132.190 107.860 132.250 ;
        RECT 108.015 132.190 108.305 132.235 ;
        RECT 107.540 132.050 108.305 132.190 ;
        RECT 104.750 132.005 105.040 132.050 ;
        RECT 107.540 131.990 107.860 132.050 ;
        RECT 108.015 132.005 108.305 132.050 ;
        RECT 109.855 131.850 110.145 131.895 ;
        RECT 102.110 131.710 110.145 131.850 ;
        RECT 109.855 131.665 110.145 131.710 ;
        RECT 104.750 131.510 105.040 131.555 ;
        RECT 107.530 131.510 107.820 131.555 ;
        RECT 109.390 131.510 109.680 131.555 ;
        RECT 104.750 131.370 109.680 131.510 ;
        RECT 104.750 131.325 105.040 131.370 ;
        RECT 107.530 131.325 107.820 131.370 ;
        RECT 109.390 131.325 109.680 131.370 ;
        RECT 105.240 131.170 105.560 131.230 ;
        RECT 101.650 131.030 105.560 131.170 ;
        RECT 90.980 130.970 91.300 131.030 ;
        RECT 98.340 130.970 98.660 131.030 ;
        RECT 99.735 130.985 100.025 131.030 ;
        RECT 105.240 130.970 105.560 131.030 ;
        RECT 22.830 130.350 113.450 130.830 ;
        RECT 37.175 130.150 37.465 130.195 ;
        RECT 37.620 130.150 37.940 130.210 ;
        RECT 40.840 130.150 41.160 130.210 ;
        RECT 37.175 130.010 37.940 130.150 ;
        RECT 37.175 129.965 37.465 130.010 ;
        RECT 37.620 129.950 37.940 130.010 ;
        RECT 38.170 130.010 41.160 130.150 ;
        RECT 25.680 129.810 25.970 129.855 ;
        RECT 27.540 129.810 27.830 129.855 ;
        RECT 30.320 129.810 30.610 129.855 ;
        RECT 25.680 129.670 30.610 129.810 ;
        RECT 25.680 129.625 25.970 129.670 ;
        RECT 27.540 129.625 27.830 129.670 ;
        RECT 30.320 129.625 30.610 129.670 ;
        RECT 35.320 129.810 35.640 129.870 ;
        RECT 38.170 129.810 38.310 130.010 ;
        RECT 40.840 129.950 41.160 130.010 ;
        RECT 41.760 130.150 42.080 130.210 ;
        RECT 44.520 130.150 44.840 130.210 ;
        RECT 47.985 130.150 48.275 130.195 ;
        RECT 41.760 130.010 48.275 130.150 ;
        RECT 41.760 129.950 42.080 130.010 ;
        RECT 44.520 129.950 44.840 130.010 ;
        RECT 47.985 129.965 48.275 130.010 ;
        RECT 50.960 130.150 51.280 130.210 ;
        RECT 52.125 130.150 52.415 130.195 ;
        RECT 50.960 130.010 52.415 130.150 ;
        RECT 50.960 129.950 51.280 130.010 ;
        RECT 52.125 129.965 52.415 130.010 ;
        RECT 62.245 130.150 62.535 130.195 ;
        RECT 63.380 130.150 63.700 130.210 ;
        RECT 62.245 130.010 63.700 130.150 ;
        RECT 62.245 129.965 62.535 130.010 ;
        RECT 63.380 129.950 63.700 130.010 ;
        RECT 65.680 130.150 66.000 130.210 ;
        RECT 81.320 130.150 81.640 130.210 ;
        RECT 65.680 130.010 81.640 130.150 ;
        RECT 65.680 129.950 66.000 130.010 ;
        RECT 81.320 129.950 81.640 130.010 ;
        RECT 85.090 130.010 87.990 130.150 ;
        RECT 35.320 129.670 38.310 129.810 ;
        RECT 39.480 129.810 39.770 129.855 ;
        RECT 41.340 129.810 41.630 129.855 ;
        RECT 44.120 129.810 44.410 129.855 ;
        RECT 39.480 129.670 44.410 129.810 ;
        RECT 35.320 129.610 35.640 129.670 ;
        RECT 39.480 129.625 39.770 129.670 ;
        RECT 41.340 129.625 41.630 129.670 ;
        RECT 44.120 129.625 44.410 129.670 ;
        RECT 46.820 129.810 47.140 129.870 ;
        RECT 71.660 129.855 71.980 129.870 ;
        RECT 49.135 129.810 49.425 129.855 ;
        RECT 46.820 129.670 49.425 129.810 ;
        RECT 46.820 129.610 47.140 129.670 ;
        RECT 49.135 129.625 49.425 129.670 ;
        RECT 55.990 129.810 56.280 129.855 ;
        RECT 58.770 129.810 59.060 129.855 ;
        RECT 60.630 129.810 60.920 129.855 ;
        RECT 55.990 129.670 60.920 129.810 ;
        RECT 55.990 129.625 56.280 129.670 ;
        RECT 58.770 129.625 59.060 129.670 ;
        RECT 60.630 129.625 60.920 129.670 ;
        RECT 66.110 129.810 66.400 129.855 ;
        RECT 68.890 129.810 69.180 129.855 ;
        RECT 70.750 129.810 71.040 129.855 ;
        RECT 66.110 129.670 71.040 129.810 ;
        RECT 66.110 129.625 66.400 129.670 ;
        RECT 68.890 129.625 69.180 129.670 ;
        RECT 70.750 129.625 71.040 129.670 ;
        RECT 71.660 129.625 72.195 129.855 ;
        RECT 75.770 129.810 76.060 129.855 ;
        RECT 78.550 129.810 78.840 129.855 ;
        RECT 80.410 129.810 80.700 129.855 ;
        RECT 75.770 129.670 80.700 129.810 ;
        RECT 75.770 129.625 76.060 129.670 ;
        RECT 78.550 129.625 78.840 129.670 ;
        RECT 80.410 129.625 80.700 129.670 ;
        RECT 71.660 129.610 71.980 129.625 ;
        RECT 27.040 129.270 27.360 129.530 ;
        RECT 34.860 129.470 35.180 129.530 ;
        RECT 39.015 129.470 39.305 129.515 ;
        RECT 34.860 129.330 39.305 129.470 ;
        RECT 34.860 129.270 35.180 129.330 ;
        RECT 39.015 129.285 39.305 129.330 ;
        RECT 39.920 129.470 40.240 129.530 ;
        RECT 50.975 129.470 51.265 129.515 ;
        RECT 39.920 129.330 51.265 129.470 ;
        RECT 39.920 129.270 40.240 129.330 ;
        RECT 50.975 129.285 51.265 129.330 ;
        RECT 57.400 129.470 57.720 129.530 ;
        RECT 59.255 129.470 59.545 129.515 ;
        RECT 59.700 129.470 60.020 129.530 ;
        RECT 79.035 129.470 79.325 129.515 ;
        RECT 79.940 129.470 80.260 129.530 ;
        RECT 57.400 129.330 59.010 129.470 ;
        RECT 57.400 129.270 57.720 129.330 ;
        RECT 25.200 128.930 25.520 129.190 ;
        RECT 30.320 129.130 30.610 129.175 ;
        RECT 28.075 128.990 30.610 129.130 ;
        RECT 28.075 128.835 28.290 128.990 ;
        RECT 30.320 128.945 30.610 128.990 ;
        RECT 38.080 128.930 38.400 129.190 ;
        RECT 39.460 129.130 39.780 129.190 ;
        RECT 40.855 129.130 41.145 129.175 ;
        RECT 44.120 129.130 44.410 129.175 ;
        RECT 39.460 128.990 41.145 129.130 ;
        RECT 39.460 128.930 39.780 128.990 ;
        RECT 40.855 128.945 41.145 128.990 ;
        RECT 41.875 128.990 44.410 129.130 ;
        RECT 26.140 128.790 26.430 128.835 ;
        RECT 28.000 128.790 28.290 128.835 ;
        RECT 28.920 128.790 29.210 128.835 ;
        RECT 32.180 128.790 32.470 128.835 ;
        RECT 26.140 128.650 28.290 128.790 ;
        RECT 26.140 128.605 26.430 128.650 ;
        RECT 28.000 128.605 28.290 128.650 ;
        RECT 28.510 128.650 32.470 128.790 ;
        RECT 24.740 128.450 25.060 128.510 ;
        RECT 28.510 128.450 28.650 128.650 ;
        RECT 28.920 128.605 29.210 128.650 ;
        RECT 32.180 128.605 32.470 128.650 ;
        RECT 34.185 128.790 34.475 128.835 ;
        RECT 35.320 128.790 35.640 128.850 ;
        RECT 41.875 128.835 42.090 128.990 ;
        RECT 44.120 128.945 44.410 128.990 ;
        RECT 44.980 129.130 45.300 129.190 ;
        RECT 50.055 129.130 50.345 129.175 ;
        RECT 52.340 129.130 52.660 129.190 ;
        RECT 44.980 128.990 52.660 129.130 ;
        RECT 44.980 128.930 45.300 128.990 ;
        RECT 50.055 128.945 50.345 128.990 ;
        RECT 52.340 128.930 52.660 128.990 ;
        RECT 55.990 129.130 56.280 129.175 ;
        RECT 58.870 129.130 59.010 129.330 ;
        RECT 59.255 129.330 60.020 129.470 ;
        RECT 59.255 129.285 59.545 129.330 ;
        RECT 59.700 129.270 60.020 129.330 ;
        RECT 71.290 129.330 78.790 129.470 ;
        RECT 61.095 129.130 61.385 129.175 ;
        RECT 55.990 128.990 58.525 129.130 ;
        RECT 58.870 128.990 61.385 129.130 ;
        RECT 55.990 128.945 56.280 128.990 ;
        RECT 58.310 128.835 58.525 128.990 ;
        RECT 61.095 128.945 61.385 128.990 ;
        RECT 66.110 129.130 66.400 129.175 ;
        RECT 66.110 128.990 68.645 129.130 ;
        RECT 66.110 128.945 66.400 128.990 ;
        RECT 34.185 128.650 35.640 128.790 ;
        RECT 34.185 128.605 34.475 128.650 ;
        RECT 35.320 128.590 35.640 128.650 ;
        RECT 39.940 128.790 40.230 128.835 ;
        RECT 41.800 128.790 42.090 128.835 ;
        RECT 42.720 128.790 43.010 128.835 ;
        RECT 45.980 128.790 46.270 128.835 ;
        RECT 39.940 128.650 42.090 128.790 ;
        RECT 39.940 128.605 40.230 128.650 ;
        RECT 41.800 128.605 42.090 128.650 ;
        RECT 42.310 128.650 46.270 128.790 ;
        RECT 24.740 128.310 28.650 128.450 ;
        RECT 31.180 128.450 31.500 128.510 ;
        RECT 42.310 128.450 42.450 128.650 ;
        RECT 42.720 128.605 43.010 128.650 ;
        RECT 45.980 128.605 46.270 128.650 ;
        RECT 54.130 128.790 54.420 128.835 ;
        RECT 57.390 128.790 57.680 128.835 ;
        RECT 58.310 128.790 58.600 128.835 ;
        RECT 60.170 128.790 60.460 128.835 ;
        RECT 54.130 128.650 58.090 128.790 ;
        RECT 54.130 128.605 54.420 128.650 ;
        RECT 57.390 128.605 57.680 128.650 ;
        RECT 31.180 128.310 42.450 128.450 ;
        RECT 57.950 128.450 58.090 128.650 ;
        RECT 58.310 128.650 60.460 128.790 ;
        RECT 58.310 128.605 58.600 128.650 ;
        RECT 60.170 128.605 60.460 128.650 ;
        RECT 64.250 128.790 64.540 128.835 ;
        RECT 64.760 128.790 65.080 128.850 ;
        RECT 68.430 128.835 68.645 128.990 ;
        RECT 69.360 128.930 69.680 129.190 ;
        RECT 70.740 129.130 71.060 129.190 ;
        RECT 71.290 129.175 71.430 129.330 ;
        RECT 71.215 129.130 71.505 129.175 ;
        RECT 70.740 128.990 71.505 129.130 ;
        RECT 70.740 128.930 71.060 128.990 ;
        RECT 71.215 128.945 71.505 128.990 ;
        RECT 75.770 129.130 76.060 129.175 ;
        RECT 78.650 129.130 78.790 129.330 ;
        RECT 79.035 129.330 80.260 129.470 ;
        RECT 79.035 129.285 79.325 129.330 ;
        RECT 79.940 129.270 80.260 129.330 ;
        RECT 80.875 129.130 81.165 129.175 ;
        RECT 75.770 128.990 78.305 129.130 ;
        RECT 78.650 128.990 81.165 129.130 ;
        RECT 81.410 129.130 81.550 129.950 ;
        RECT 85.090 129.870 85.230 130.010 ;
        RECT 85.000 129.810 85.320 129.870 ;
        RECT 84.170 129.670 85.320 129.810 ;
        RECT 84.170 129.515 84.310 129.670 ;
        RECT 85.000 129.610 85.320 129.670 ;
        RECT 86.855 129.625 87.145 129.855 ;
        RECT 87.850 129.810 87.990 130.010 ;
        RECT 88.220 129.950 88.540 130.210 ;
        RECT 92.360 130.150 92.680 130.210 ;
        RECT 95.135 130.150 95.425 130.195 ;
        RECT 92.360 130.010 95.425 130.150 ;
        RECT 92.360 129.950 92.680 130.010 ;
        RECT 95.135 129.965 95.425 130.010 ;
        RECT 99.260 129.950 99.580 130.210 ;
        RECT 104.320 129.950 104.640 130.210 ;
        RECT 105.700 129.950 106.020 130.210 ;
        RECT 107.080 130.150 107.400 130.210 ;
        RECT 107.555 130.150 107.845 130.195 ;
        RECT 107.080 130.010 107.845 130.150 ;
        RECT 107.080 129.950 107.400 130.010 ;
        RECT 107.555 129.965 107.845 130.010 ;
        RECT 90.980 129.810 91.300 129.870 ;
        RECT 87.850 129.670 91.670 129.810 ;
        RECT 84.095 129.285 84.385 129.515 ;
        RECT 84.540 129.270 84.860 129.530 ;
        RECT 86.930 129.470 87.070 129.625 ;
        RECT 90.980 129.610 91.300 129.670 ;
        RECT 91.530 129.515 91.670 129.670 ;
        RECT 94.675 129.625 94.965 129.855 ;
        RECT 103.415 129.810 103.705 129.855 ;
        RECT 103.415 129.670 105.240 129.810 ;
        RECT 103.415 129.625 103.705 129.670 ;
        RECT 86.930 129.330 89.370 129.470 ;
        RECT 89.230 129.175 89.370 129.330 ;
        RECT 91.455 129.285 91.745 129.515 ;
        RECT 92.360 129.270 92.680 129.530 ;
        RECT 82.255 129.130 82.545 129.175 ;
        RECT 87.775 129.130 88.065 129.175 ;
        RECT 81.410 128.990 88.065 129.130 ;
        RECT 75.770 128.945 76.060 128.990 ;
        RECT 78.090 128.835 78.305 128.990 ;
        RECT 80.875 128.945 81.165 128.990 ;
        RECT 82.255 128.945 82.545 128.990 ;
        RECT 87.775 128.945 88.065 128.990 ;
        RECT 89.155 128.945 89.445 129.175 ;
        RECT 94.750 129.130 94.890 129.625 ;
        RECT 96.500 129.470 96.820 129.530 ;
        RECT 100.195 129.470 100.485 129.515 ;
        RECT 96.500 129.330 100.485 129.470 ;
        RECT 96.500 129.270 96.820 129.330 ;
        RECT 100.195 129.285 100.485 129.330 ;
        RECT 101.115 129.470 101.405 129.515 ;
        RECT 102.480 129.470 102.800 129.530 ;
        RECT 101.115 129.330 102.800 129.470 ;
        RECT 105.100 129.470 105.240 129.670 ;
        RECT 105.100 129.330 106.850 129.470 ;
        RECT 101.115 129.285 101.405 129.330 ;
        RECT 102.480 129.270 102.800 129.330 ;
        RECT 96.055 129.130 96.345 129.175 ;
        RECT 94.750 128.990 96.345 129.130 ;
        RECT 96.055 128.945 96.345 128.990 ;
        RECT 67.510 128.790 67.800 128.835 ;
        RECT 64.250 128.650 67.800 128.790 ;
        RECT 64.250 128.605 64.540 128.650 ;
        RECT 64.760 128.590 65.080 128.650 ;
        RECT 67.510 128.605 67.800 128.650 ;
        RECT 68.430 128.790 68.720 128.835 ;
        RECT 70.290 128.790 70.580 128.835 ;
        RECT 73.910 128.790 74.200 128.835 ;
        RECT 77.170 128.790 77.460 128.835 ;
        RECT 68.430 128.650 70.580 128.790 ;
        RECT 68.430 128.605 68.720 128.650 ;
        RECT 70.290 128.605 70.580 128.650 ;
        RECT 70.830 128.650 77.460 128.790 ;
        RECT 70.830 128.510 70.970 128.650 ;
        RECT 73.910 128.605 74.200 128.650 ;
        RECT 77.170 128.605 77.460 128.650 ;
        RECT 78.090 128.790 78.380 128.835 ;
        RECT 79.950 128.790 80.240 128.835 ;
        RECT 78.090 128.650 80.240 128.790 ;
        RECT 80.950 128.790 81.090 128.945 ;
        RECT 98.340 128.930 98.660 129.190 ;
        RECT 98.800 129.130 99.120 129.190 ;
        RECT 101.575 129.130 101.865 129.175 ;
        RECT 98.800 128.990 101.865 129.130 ;
        RECT 98.800 128.930 99.120 128.990 ;
        RECT 101.575 128.945 101.865 128.990 ;
        RECT 103.875 129.130 104.165 129.175 ;
        RECT 105.240 129.130 105.560 129.190 ;
        RECT 106.710 129.175 106.850 129.330 ;
        RECT 103.875 128.990 105.560 129.130 ;
        RECT 103.875 128.945 104.165 128.990 ;
        RECT 105.240 128.930 105.560 128.990 ;
        RECT 106.635 128.945 106.925 129.175 ;
        RECT 84.080 128.790 84.400 128.850 ;
        RECT 80.950 128.650 84.400 128.790 ;
        RECT 78.090 128.605 78.380 128.650 ;
        RECT 79.950 128.605 80.240 128.650 ;
        RECT 84.080 128.590 84.400 128.650 ;
        RECT 88.220 128.790 88.540 128.850 ;
        RECT 92.835 128.790 93.125 128.835 ;
        RECT 88.220 128.650 93.125 128.790 ;
        RECT 88.220 128.590 88.540 128.650 ;
        RECT 92.835 128.605 93.125 128.650 ;
        RECT 94.200 128.790 94.520 128.850 ;
        RECT 101.100 128.790 101.420 128.850 ;
        RECT 94.200 128.650 101.420 128.790 ;
        RECT 94.200 128.590 94.520 128.650 ;
        RECT 101.100 128.590 101.420 128.650 ;
        RECT 59.240 128.450 59.560 128.510 ;
        RECT 57.950 128.310 59.560 128.450 ;
        RECT 24.740 128.250 25.060 128.310 ;
        RECT 31.180 128.250 31.500 128.310 ;
        RECT 59.240 128.250 59.560 128.310 ;
        RECT 70.740 128.250 71.060 128.510 ;
        RECT 80.400 128.450 80.720 128.510 ;
        RECT 81.795 128.450 82.085 128.495 ;
        RECT 80.400 128.310 82.085 128.450 ;
        RECT 80.400 128.250 80.720 128.310 ;
        RECT 81.795 128.265 82.085 128.310 ;
        RECT 83.620 128.450 83.940 128.510 ;
        RECT 85.015 128.450 85.305 128.495 ;
        RECT 83.620 128.310 85.305 128.450 ;
        RECT 83.620 128.250 83.940 128.310 ;
        RECT 85.015 128.265 85.305 128.310 ;
        RECT 90.075 128.450 90.365 128.495 ;
        RECT 91.900 128.450 92.220 128.510 ;
        RECT 90.075 128.310 92.220 128.450 ;
        RECT 90.075 128.265 90.365 128.310 ;
        RECT 91.900 128.250 92.220 128.310 ;
        RECT 22.830 127.630 113.450 128.110 ;
        RECT 24.740 127.230 25.060 127.490 ;
        RECT 27.975 127.245 28.265 127.475 ;
        RECT 28.050 127.090 28.190 127.245 ;
        RECT 28.420 127.230 28.740 127.490 ;
        RECT 30.735 127.430 31.025 127.475 ;
        RECT 32.805 127.430 33.095 127.475 ;
        RECT 36.240 127.430 36.560 127.490 ;
        RECT 43.600 127.430 43.920 127.490 ;
        RECT 30.735 127.290 36.560 127.430 ;
        RECT 30.735 127.245 31.025 127.290 ;
        RECT 32.805 127.245 33.095 127.290 ;
        RECT 36.240 127.230 36.560 127.290 ;
        RECT 38.630 127.290 43.920 127.430 ;
        RECT 31.640 127.090 31.960 127.150 ;
        RECT 28.050 126.950 31.960 127.090 ;
        RECT 31.640 126.890 31.960 126.950 ;
        RECT 34.810 127.090 35.100 127.135 ;
        RECT 38.070 127.090 38.360 127.135 ;
        RECT 38.630 127.090 38.770 127.290 ;
        RECT 43.600 127.230 43.920 127.290 ;
        RECT 49.365 127.430 49.655 127.475 ;
        RECT 53.720 127.430 54.040 127.490 ;
        RECT 49.365 127.290 54.040 127.430 ;
        RECT 49.365 127.245 49.655 127.290 ;
        RECT 53.720 127.230 54.040 127.290 ;
        RECT 59.240 127.230 59.560 127.490 ;
        RECT 59.700 127.430 60.020 127.490 ;
        RECT 60.635 127.430 60.925 127.475 ;
        RECT 59.700 127.290 60.925 127.430 ;
        RECT 59.700 127.230 60.020 127.290 ;
        RECT 60.635 127.245 60.925 127.290 ;
        RECT 64.315 127.430 64.605 127.475 ;
        RECT 64.760 127.430 65.080 127.490 ;
        RECT 64.315 127.290 65.080 127.430 ;
        RECT 64.315 127.245 64.605 127.290 ;
        RECT 64.760 127.230 65.080 127.290 ;
        RECT 67.075 127.430 67.365 127.475 ;
        RECT 69.360 127.430 69.680 127.490 ;
        RECT 67.075 127.290 69.680 127.430 ;
        RECT 67.075 127.245 67.365 127.290 ;
        RECT 69.360 127.230 69.680 127.290 ;
        RECT 70.740 127.230 71.060 127.490 ;
        RECT 72.135 127.430 72.425 127.475 ;
        RECT 74.420 127.430 74.740 127.490 ;
        RECT 72.135 127.290 74.740 127.430 ;
        RECT 72.135 127.245 72.425 127.290 ;
        RECT 74.420 127.230 74.740 127.290 ;
        RECT 75.125 127.430 75.415 127.475 ;
        RECT 76.260 127.430 76.580 127.490 ;
        RECT 75.125 127.290 76.580 127.430 ;
        RECT 75.125 127.245 75.415 127.290 ;
        RECT 76.260 127.230 76.580 127.290 ;
        RECT 83.620 127.430 83.940 127.490 ;
        RECT 84.785 127.430 85.075 127.475 ;
        RECT 83.620 127.290 85.075 127.430 ;
        RECT 83.620 127.230 83.940 127.290 ;
        RECT 84.785 127.245 85.075 127.290 ;
        RECT 34.810 126.950 38.770 127.090 ;
        RECT 38.990 127.090 39.280 127.135 ;
        RECT 40.850 127.090 41.140 127.135 ;
        RECT 38.990 126.950 41.140 127.090 ;
        RECT 34.810 126.905 35.100 126.950 ;
        RECT 38.070 126.905 38.360 126.950 ;
        RECT 38.990 126.905 39.280 126.950 ;
        RECT 40.850 126.905 41.140 126.950 ;
        RECT 44.060 127.090 44.380 127.150 ;
        RECT 45.455 127.090 45.745 127.135 ;
        RECT 44.060 126.950 45.745 127.090 ;
        RECT 25.215 126.750 25.505 126.795 ;
        RECT 25.660 126.750 25.980 126.810 ;
        RECT 25.215 126.610 25.980 126.750 ;
        RECT 25.215 126.565 25.505 126.610 ;
        RECT 25.660 126.550 25.980 126.610 ;
        RECT 27.055 126.750 27.345 126.795 ;
        RECT 27.960 126.750 28.280 126.810 ;
        RECT 27.055 126.610 28.280 126.750 ;
        RECT 27.055 126.565 27.345 126.610 ;
        RECT 27.960 126.550 28.280 126.610 ;
        RECT 30.275 126.750 30.565 126.795 ;
        RECT 30.720 126.750 31.040 126.810 ;
        RECT 35.320 126.750 35.640 126.810 ;
        RECT 30.275 126.610 35.640 126.750 ;
        RECT 30.275 126.565 30.565 126.610 ;
        RECT 30.720 126.550 31.040 126.610 ;
        RECT 35.320 126.550 35.640 126.610 ;
        RECT 36.670 126.750 36.960 126.795 ;
        RECT 38.990 126.750 39.205 126.905 ;
        RECT 44.060 126.890 44.380 126.950 ;
        RECT 45.455 126.905 45.745 126.950 ;
        RECT 47.755 127.090 48.045 127.135 ;
        RECT 51.370 127.090 51.660 127.135 ;
        RECT 54.630 127.090 54.920 127.135 ;
        RECT 47.755 126.950 54.920 127.090 ;
        RECT 47.755 126.905 48.045 126.950 ;
        RECT 51.370 126.905 51.660 126.950 ;
        RECT 54.630 126.905 54.920 126.950 ;
        RECT 55.550 127.090 55.840 127.135 ;
        RECT 57.410 127.090 57.700 127.135 ;
        RECT 55.550 126.950 57.700 127.090 ;
        RECT 55.550 126.905 55.840 126.950 ;
        RECT 57.410 126.905 57.700 126.950 ;
        RECT 65.680 127.090 66.000 127.150 ;
        RECT 80.400 127.135 80.720 127.150 ;
        RECT 77.130 127.090 77.420 127.135 ;
        RECT 80.390 127.090 80.720 127.135 ;
        RECT 65.680 126.950 70.510 127.090 ;
        RECT 36.670 126.610 39.205 126.750 ;
        RECT 36.670 126.565 36.960 126.610 ;
        RECT 39.920 126.550 40.240 126.810 ;
        RECT 41.300 126.750 41.620 126.810 ;
        RECT 43.155 126.750 43.445 126.795 ;
        RECT 44.980 126.750 45.300 126.810 ;
        RECT 41.300 126.610 45.300 126.750 ;
        RECT 41.300 126.550 41.620 126.610 ;
        RECT 43.155 126.565 43.445 126.610 ;
        RECT 44.980 126.550 45.300 126.610 ;
        RECT 45.900 126.750 46.220 126.810 ;
        RECT 46.820 126.750 47.140 126.810 ;
        RECT 47.295 126.750 47.585 126.795 ;
        RECT 45.900 126.610 47.585 126.750 ;
        RECT 45.900 126.550 46.220 126.610 ;
        RECT 46.820 126.550 47.140 126.610 ;
        RECT 47.295 126.565 47.585 126.610 ;
        RECT 53.230 126.750 53.520 126.795 ;
        RECT 55.550 126.750 55.765 126.905 ;
        RECT 65.680 126.890 66.000 126.950 ;
        RECT 53.230 126.610 55.765 126.750 ;
        RECT 59.715 126.750 60.005 126.795 ;
        RECT 60.620 126.750 60.940 126.810 ;
        RECT 59.715 126.610 60.940 126.750 ;
        RECT 53.230 126.565 53.520 126.610 ;
        RECT 59.715 126.565 60.005 126.610 ;
        RECT 60.620 126.550 60.940 126.610 ;
        RECT 61.540 126.550 61.860 126.810 ;
        RECT 63.855 126.565 64.145 126.795 ;
        RECT 26.135 126.410 26.425 126.455 ;
        RECT 31.180 126.410 31.500 126.470 ;
        RECT 26.135 126.270 31.500 126.410 ;
        RECT 26.135 126.225 26.425 126.270 ;
        RECT 31.180 126.210 31.500 126.270 ;
        RECT 31.655 126.410 31.945 126.455 ;
        RECT 32.100 126.410 32.420 126.470 ;
        RECT 31.655 126.270 32.420 126.410 ;
        RECT 31.655 126.225 31.945 126.270 ;
        RECT 32.100 126.210 32.420 126.270 ;
        RECT 37.620 126.410 37.940 126.470 ;
        RECT 41.775 126.410 42.065 126.455 ;
        RECT 37.620 126.270 42.065 126.410 ;
        RECT 37.620 126.210 37.940 126.270 ;
        RECT 41.775 126.225 42.065 126.270 ;
        RECT 42.235 126.225 42.525 126.455 ;
        RECT 44.075 126.410 44.365 126.455 ;
        RECT 50.040 126.410 50.360 126.470 ;
        RECT 44.075 126.270 50.360 126.410 ;
        RECT 44.075 126.225 44.365 126.270 ;
        RECT 36.670 126.070 36.960 126.115 ;
        RECT 39.450 126.070 39.740 126.115 ;
        RECT 41.310 126.070 41.600 126.115 ;
        RECT 36.670 125.930 41.600 126.070 ;
        RECT 36.670 125.885 36.960 125.930 ;
        RECT 39.450 125.885 39.740 125.930 ;
        RECT 41.310 125.885 41.600 125.930 ;
        RECT 35.320 125.730 35.640 125.790 ;
        RECT 42.310 125.730 42.450 126.225 ;
        RECT 50.040 126.210 50.360 126.270 ;
        RECT 56.480 126.210 56.800 126.470 ;
        RECT 57.400 126.410 57.720 126.470 ;
        RECT 58.335 126.410 58.625 126.455 ;
        RECT 57.400 126.270 58.625 126.410 ;
        RECT 60.710 126.410 60.850 126.550 ;
        RECT 63.930 126.410 64.070 126.565 ;
        RECT 66.140 126.550 66.460 126.810 ;
        RECT 70.370 126.795 70.510 126.950 ;
        RECT 77.130 126.950 80.720 127.090 ;
        RECT 77.130 126.905 77.420 126.950 ;
        RECT 80.390 126.905 80.720 126.950 ;
        RECT 80.400 126.890 80.720 126.905 ;
        RECT 81.310 127.090 81.600 127.135 ;
        RECT 83.170 127.090 83.460 127.135 ;
        RECT 81.310 126.950 83.460 127.090 ;
        RECT 81.310 126.905 81.600 126.950 ;
        RECT 83.170 126.905 83.460 126.950 ;
        RECT 85.460 127.090 85.780 127.150 ;
        RECT 86.790 127.090 87.080 127.135 ;
        RECT 90.050 127.090 90.340 127.135 ;
        RECT 85.460 126.950 90.340 127.090 ;
        RECT 70.295 126.750 70.585 126.795 ;
        RECT 71.675 126.750 71.965 126.795 ;
        RECT 70.295 126.610 71.965 126.750 ;
        RECT 70.295 126.565 70.585 126.610 ;
        RECT 71.675 126.565 71.965 126.610 ;
        RECT 78.990 126.750 79.280 126.795 ;
        RECT 81.310 126.750 81.525 126.905 ;
        RECT 85.460 126.890 85.780 126.950 ;
        RECT 86.790 126.905 87.080 126.950 ;
        RECT 90.050 126.905 90.340 126.950 ;
        RECT 90.970 127.090 91.260 127.135 ;
        RECT 92.830 127.090 93.120 127.135 ;
        RECT 90.970 126.950 93.120 127.090 ;
        RECT 90.970 126.905 91.260 126.950 ;
        RECT 92.830 126.905 93.120 126.950 ;
        RECT 78.990 126.610 81.525 126.750 ;
        RECT 78.990 126.565 79.280 126.610 ;
        RECT 84.080 126.550 84.400 126.810 ;
        RECT 88.650 126.750 88.940 126.795 ;
        RECT 90.970 126.750 91.185 126.905 ;
        RECT 88.650 126.610 91.185 126.750 ;
        RECT 88.650 126.565 88.940 126.610 ;
        RECT 91.900 126.550 92.220 126.810 ;
        RECT 93.755 126.750 94.045 126.795 ;
        RECT 94.660 126.750 94.980 126.810 ;
        RECT 93.755 126.610 94.980 126.750 ;
        RECT 93.755 126.565 94.045 126.610 ;
        RECT 94.660 126.550 94.980 126.610 ;
        RECT 106.160 126.550 106.480 126.810 ;
        RECT 106.620 126.750 106.940 126.810 ;
        RECT 109.855 126.750 110.145 126.795 ;
        RECT 106.620 126.610 110.145 126.750 ;
        RECT 106.620 126.550 106.940 126.610 ;
        RECT 109.855 126.565 110.145 126.610 ;
        RECT 111.680 126.550 112.000 126.810 ;
        RECT 60.710 126.270 64.070 126.410 ;
        RECT 79.940 126.410 80.260 126.470 ;
        RECT 82.255 126.410 82.545 126.455 ;
        RECT 79.940 126.270 82.545 126.410 ;
        RECT 57.400 126.210 57.720 126.270 ;
        RECT 58.335 126.225 58.625 126.270 ;
        RECT 79.940 126.210 80.260 126.270 ;
        RECT 82.255 126.225 82.545 126.270 ;
        RECT 88.310 126.270 110.990 126.410 ;
        RECT 53.230 126.070 53.520 126.115 ;
        RECT 56.010 126.070 56.300 126.115 ;
        RECT 57.870 126.070 58.160 126.115 ;
        RECT 53.230 125.930 58.160 126.070 ;
        RECT 53.230 125.885 53.520 125.930 ;
        RECT 56.010 125.885 56.300 125.930 ;
        RECT 57.870 125.885 58.160 125.930 ;
        RECT 78.990 126.070 79.280 126.115 ;
        RECT 81.770 126.070 82.060 126.115 ;
        RECT 83.630 126.070 83.920 126.115 ;
        RECT 78.990 125.930 83.920 126.070 ;
        RECT 78.990 125.885 79.280 125.930 ;
        RECT 81.770 125.885 82.060 125.930 ;
        RECT 83.630 125.885 83.920 125.930 ;
        RECT 35.320 125.590 42.450 125.730 ;
        RECT 73.960 125.730 74.280 125.790 ;
        RECT 88.310 125.730 88.450 126.270 ;
        RECT 88.650 126.070 88.940 126.115 ;
        RECT 91.430 126.070 91.720 126.115 ;
        RECT 93.290 126.070 93.580 126.115 ;
        RECT 88.650 125.930 93.580 126.070 ;
        RECT 88.650 125.885 88.940 125.930 ;
        RECT 91.430 125.885 91.720 125.930 ;
        RECT 93.290 125.885 93.580 125.930 ;
        RECT 102.940 126.070 103.260 126.130 ;
        RECT 110.850 126.115 110.990 126.270 ;
        RECT 108.935 126.070 109.225 126.115 ;
        RECT 102.940 125.930 109.225 126.070 ;
        RECT 102.940 125.870 103.260 125.930 ;
        RECT 108.935 125.885 109.225 125.930 ;
        RECT 110.775 125.885 111.065 126.115 ;
        RECT 73.960 125.590 88.450 125.730 ;
        RECT 35.320 125.530 35.640 125.590 ;
        RECT 73.960 125.530 74.280 125.590 ;
        RECT 106.620 125.530 106.940 125.790 ;
        RECT 22.830 124.910 113.450 125.390 ;
        RECT 39.460 124.510 39.780 124.770 ;
        RECT 42.220 124.510 42.540 124.770 ;
        RECT 56.035 124.710 56.325 124.755 ;
        RECT 56.480 124.710 56.800 124.770 ;
        RECT 56.035 124.570 56.800 124.710 ;
        RECT 56.035 124.525 56.325 124.570 ;
        RECT 56.480 124.510 56.800 124.570 ;
        RECT 79.940 124.510 80.260 124.770 ;
        RECT 106.160 124.710 106.480 124.770 ;
        RECT 100.270 124.570 106.480 124.710 ;
        RECT 28.535 124.370 28.825 124.415 ;
        RECT 31.655 124.370 31.945 124.415 ;
        RECT 33.545 124.370 33.835 124.415 ;
        RECT 28.535 124.230 33.835 124.370 ;
        RECT 28.535 124.185 28.825 124.230 ;
        RECT 31.655 124.185 31.945 124.230 ;
        RECT 33.545 124.185 33.835 124.230 ;
        RECT 38.095 124.370 38.385 124.415 ;
        RECT 39.920 124.370 40.240 124.430 ;
        RECT 38.095 124.230 40.240 124.370 ;
        RECT 38.095 124.185 38.385 124.230 ;
        RECT 39.920 124.170 40.240 124.230 ;
        RECT 46.935 124.370 47.225 124.415 ;
        RECT 50.055 124.370 50.345 124.415 ;
        RECT 51.945 124.370 52.235 124.415 ;
        RECT 46.935 124.230 52.235 124.370 ;
        RECT 46.935 124.185 47.225 124.230 ;
        RECT 50.055 124.185 50.345 124.230 ;
        RECT 51.945 124.185 52.235 124.230 ;
        RECT 96.055 124.370 96.345 124.415 ;
        RECT 99.720 124.370 100.040 124.430 ;
        RECT 96.055 124.230 100.040 124.370 ;
        RECT 96.055 124.185 96.345 124.230 ;
        RECT 99.720 124.170 100.040 124.230 ;
        RECT 34.415 124.030 34.705 124.075 ;
        RECT 34.860 124.030 35.180 124.090 ;
        RECT 37.620 124.030 37.940 124.090 ;
        RECT 34.415 123.890 37.940 124.030 ;
        RECT 34.415 123.845 34.705 123.890 ;
        RECT 34.860 123.830 35.180 123.890 ;
        RECT 37.620 123.830 37.940 123.890 ;
        RECT 40.380 123.830 40.700 124.090 ;
        RECT 48.200 124.030 48.520 124.090 ;
        RECT 52.815 124.030 53.105 124.075 ;
        RECT 57.400 124.030 57.720 124.090 ;
        RECT 61.080 124.030 61.400 124.090 ;
        RECT 48.200 123.890 61.400 124.030 ;
        RECT 48.200 123.830 48.520 123.890 ;
        RECT 52.815 123.845 53.105 123.890 ;
        RECT 57.400 123.830 57.720 123.890 ;
        RECT 61.080 123.830 61.400 123.890 ;
        RECT 90.520 124.030 90.840 124.090 ;
        RECT 90.520 123.890 96.730 124.030 ;
        RECT 90.520 123.830 90.840 123.890 ;
        RECT 20.140 123.350 20.460 123.410 ;
        RECT 24.295 123.350 24.585 123.395 ;
        RECT 20.140 123.210 24.585 123.350 ;
        RECT 20.140 123.150 20.460 123.210 ;
        RECT 24.295 123.165 24.585 123.210 ;
        RECT 26.120 123.350 26.440 123.410 ;
        RECT 27.455 123.395 27.745 123.710 ;
        RECT 28.535 123.690 28.825 123.735 ;
        RECT 32.115 123.690 32.405 123.735 ;
        RECT 33.950 123.690 34.240 123.735 ;
        RECT 28.535 123.550 34.240 123.690 ;
        RECT 28.535 123.505 28.825 123.550 ;
        RECT 32.115 123.505 32.405 123.550 ;
        RECT 33.950 123.505 34.240 123.550 ;
        RECT 37.160 123.490 37.480 123.750 ;
        RECT 38.540 123.490 38.860 123.750 ;
        RECT 41.300 123.490 41.620 123.750 ;
        RECT 27.155 123.350 27.745 123.395 ;
        RECT 30.395 123.350 31.045 123.395 ;
        RECT 26.120 123.210 31.045 123.350 ;
        RECT 26.120 123.150 26.440 123.210 ;
        RECT 27.155 123.165 27.445 123.210 ;
        RECT 30.395 123.165 31.045 123.210 ;
        RECT 33.035 123.165 33.325 123.395 ;
        RECT 42.695 123.350 42.985 123.395 ;
        RECT 44.060 123.350 44.380 123.410 ;
        RECT 42.695 123.210 44.380 123.350 ;
        RECT 42.695 123.165 42.985 123.210 ;
        RECT 25.660 123.010 25.980 123.070 ;
        RECT 33.110 123.010 33.250 123.165 ;
        RECT 44.060 123.150 44.380 123.210 ;
        RECT 44.980 123.350 45.300 123.410 ;
        RECT 45.855 123.395 46.145 123.710 ;
        RECT 46.935 123.690 47.225 123.735 ;
        RECT 50.515 123.690 50.805 123.735 ;
        RECT 52.350 123.690 52.640 123.735 ;
        RECT 46.935 123.550 52.640 123.690 ;
        RECT 46.935 123.505 47.225 123.550 ;
        RECT 50.515 123.505 50.805 123.550 ;
        RECT 52.350 123.505 52.640 123.550 ;
        RECT 56.940 123.490 57.260 123.750 ;
        RECT 58.780 123.490 59.100 123.750 ;
        RECT 60.160 123.690 60.480 123.750 ;
        RECT 63.855 123.690 64.145 123.735 ;
        RECT 60.160 123.550 64.145 123.690 ;
        RECT 60.160 123.490 60.480 123.550 ;
        RECT 63.855 123.505 64.145 123.550 ;
        RECT 70.280 123.690 70.600 123.750 ;
        RECT 74.895 123.690 75.185 123.735 ;
        RECT 70.280 123.550 75.185 123.690 ;
        RECT 70.280 123.490 70.600 123.550 ;
        RECT 74.895 123.505 75.185 123.550 ;
        RECT 76.275 123.505 76.565 123.735 ;
        RECT 79.035 123.690 79.325 123.735 ;
        RECT 79.480 123.690 79.800 123.750 ;
        RECT 79.035 123.550 79.800 123.690 ;
        RECT 79.035 123.505 79.325 123.550 ;
        RECT 45.555 123.350 46.145 123.395 ;
        RECT 48.795 123.350 49.445 123.395 ;
        RECT 44.980 123.210 49.445 123.350 ;
        RECT 44.980 123.150 45.300 123.210 ;
        RECT 45.555 123.165 45.845 123.210 ;
        RECT 48.795 123.165 49.445 123.210 ;
        RECT 51.420 123.150 51.740 123.410 ;
        RECT 76.350 123.350 76.490 123.505 ;
        RECT 79.480 123.490 79.800 123.550 ;
        RECT 91.440 123.690 91.760 123.750 ;
        RECT 92.835 123.690 93.125 123.735 ;
        RECT 91.440 123.550 93.125 123.690 ;
        RECT 91.440 123.490 91.760 123.550 ;
        RECT 92.835 123.505 93.125 123.550 ;
        RECT 95.135 123.690 95.425 123.735 ;
        RECT 96.040 123.690 96.360 123.750 ;
        RECT 96.590 123.735 96.730 123.890 ;
        RECT 100.270 123.735 100.410 124.570 ;
        RECT 106.160 124.510 106.480 124.570 ;
        RECT 102.445 124.370 102.735 124.415 ;
        RECT 104.335 124.370 104.625 124.415 ;
        RECT 107.455 124.370 107.745 124.415 ;
        RECT 102.445 124.230 107.745 124.370 ;
        RECT 102.445 124.185 102.735 124.230 ;
        RECT 104.335 124.185 104.625 124.230 ;
        RECT 107.455 124.185 107.745 124.230 ;
        RECT 101.100 124.030 101.420 124.090 ;
        RECT 101.575 124.030 101.865 124.075 ;
        RECT 101.100 123.890 101.865 124.030 ;
        RECT 101.100 123.830 101.420 123.890 ;
        RECT 101.575 123.845 101.865 123.890 ;
        RECT 102.940 123.830 103.260 124.090 ;
        RECT 95.135 123.550 96.360 123.690 ;
        RECT 95.135 123.505 95.425 123.550 ;
        RECT 96.040 123.490 96.360 123.550 ;
        RECT 96.515 123.505 96.805 123.735 ;
        RECT 97.895 123.505 98.185 123.735 ;
        RECT 100.195 123.505 100.485 123.735 ;
        RECT 102.040 123.690 102.330 123.735 ;
        RECT 103.875 123.690 104.165 123.735 ;
        RECT 107.455 123.690 107.745 123.735 ;
        RECT 102.040 123.550 107.745 123.690 ;
        RECT 102.040 123.505 102.330 123.550 ;
        RECT 103.875 123.505 104.165 123.550 ;
        RECT 107.455 123.505 107.745 123.550 ;
        RECT 56.800 123.210 76.490 123.350 ;
        RECT 77.655 123.350 77.945 123.395 ;
        RECT 79.940 123.350 80.260 123.410 ;
        RECT 77.655 123.210 80.260 123.350 ;
        RECT 25.660 122.870 33.250 123.010 ;
        RECT 46.820 123.010 47.140 123.070 ;
        RECT 55.560 123.010 55.880 123.070 ;
        RECT 56.800 123.010 56.940 123.210 ;
        RECT 77.655 123.165 77.945 123.210 ;
        RECT 79.940 123.150 80.260 123.210 ;
        RECT 95.580 123.350 95.900 123.410 ;
        RECT 97.970 123.350 98.110 123.505 ;
        RECT 95.580 123.210 98.110 123.350 ;
        RECT 105.235 123.350 105.885 123.395 ;
        RECT 106.620 123.350 106.940 123.410 ;
        RECT 108.535 123.395 108.825 123.710 ;
        RECT 108.535 123.350 109.125 123.395 ;
        RECT 105.235 123.210 109.125 123.350 ;
        RECT 95.580 123.150 95.900 123.210 ;
        RECT 105.235 123.165 105.885 123.210 ;
        RECT 106.620 123.150 106.940 123.210 ;
        RECT 108.835 123.165 109.125 123.210 ;
        RECT 111.695 123.350 111.985 123.395 ;
        RECT 116.280 123.350 116.600 123.410 ;
        RECT 111.695 123.210 116.600 123.350 ;
        RECT 111.695 123.165 111.985 123.210 ;
        RECT 116.280 123.150 116.600 123.210 ;
        RECT 46.820 122.870 56.940 123.010 ;
        RECT 25.660 122.810 25.980 122.870 ;
        RECT 46.820 122.810 47.140 122.870 ;
        RECT 55.560 122.810 55.880 122.870 ;
        RECT 59.700 122.810 60.020 123.070 ;
        RECT 64.775 123.010 65.065 123.055 ;
        RECT 67.060 123.010 67.380 123.070 ;
        RECT 64.775 122.870 67.380 123.010 ;
        RECT 64.775 122.825 65.065 122.870 ;
        RECT 67.060 122.810 67.380 122.870 ;
        RECT 75.815 123.010 76.105 123.055 ;
        RECT 83.620 123.010 83.940 123.070 ;
        RECT 75.815 122.870 83.940 123.010 ;
        RECT 75.815 122.825 76.105 122.870 ;
        RECT 83.620 122.810 83.940 122.870 ;
        RECT 93.755 123.010 94.045 123.055 ;
        RECT 96.500 123.010 96.820 123.070 ;
        RECT 93.755 122.870 96.820 123.010 ;
        RECT 93.755 122.825 94.045 122.870 ;
        RECT 96.500 122.810 96.820 122.870 ;
        RECT 97.420 122.810 97.740 123.070 ;
        RECT 98.800 122.810 99.120 123.070 ;
        RECT 100.655 123.010 100.945 123.055 ;
        RECT 102.020 123.010 102.340 123.070 ;
        RECT 100.655 122.870 102.340 123.010 ;
        RECT 100.655 122.825 100.945 122.870 ;
        RECT 102.020 122.810 102.340 122.870 ;
        RECT 22.830 122.190 113.450 122.670 ;
        RECT 25.215 121.990 25.505 122.035 ;
        RECT 25.660 121.990 25.980 122.050 ;
        RECT 25.215 121.850 25.980 121.990 ;
        RECT 25.215 121.805 25.505 121.850 ;
        RECT 25.660 121.790 25.980 121.850 ;
        RECT 26.120 121.790 26.440 122.050 ;
        RECT 50.975 121.990 51.265 122.035 ;
        RECT 51.420 121.990 51.740 122.050 ;
        RECT 50.975 121.850 51.740 121.990 ;
        RECT 50.975 121.805 51.265 121.850 ;
        RECT 51.420 121.790 51.740 121.850 ;
        RECT 55.100 121.990 55.420 122.050 ;
        RECT 69.360 121.990 69.680 122.050 ;
        RECT 73.515 121.990 73.805 122.035 ;
        RECT 55.100 121.850 69.130 121.990 ;
        RECT 55.100 121.790 55.420 121.850 ;
        RECT 30.375 121.650 30.665 121.695 ;
        RECT 33.615 121.650 34.265 121.695 ;
        RECT 35.780 121.650 36.100 121.710 ;
        RECT 30.375 121.510 36.100 121.650 ;
        RECT 30.375 121.465 30.965 121.510 ;
        RECT 33.615 121.465 34.265 121.510 ;
        RECT 24.280 121.110 24.600 121.370 ;
        RECT 26.580 121.110 26.900 121.370 ;
        RECT 30.675 121.150 30.965 121.465 ;
        RECT 35.780 121.450 36.100 121.510 ;
        RECT 38.095 121.465 38.385 121.695 ;
        RECT 39.920 121.650 40.240 121.710 ;
        RECT 40.955 121.650 41.245 121.695 ;
        RECT 44.195 121.650 44.845 121.695 ;
        RECT 39.920 121.510 44.845 121.650 ;
        RECT 31.755 121.310 32.045 121.355 ;
        RECT 35.335 121.310 35.625 121.355 ;
        RECT 37.170 121.310 37.460 121.355 ;
        RECT 31.755 121.170 37.460 121.310 ;
        RECT 31.755 121.125 32.045 121.170 ;
        RECT 35.335 121.125 35.625 121.170 ;
        RECT 37.170 121.125 37.460 121.170 ;
        RECT 37.620 121.110 37.940 121.370 ;
        RECT 38.170 121.310 38.310 121.465 ;
        RECT 39.920 121.450 40.240 121.510 ;
        RECT 40.955 121.465 41.545 121.510 ;
        RECT 44.195 121.465 44.845 121.510 ;
        RECT 46.360 121.650 46.680 121.710 ;
        RECT 61.195 121.650 61.485 121.695 ;
        RECT 62.000 121.650 62.320 121.710 ;
        RECT 64.435 121.650 65.085 121.695 ;
        RECT 46.360 121.510 55.330 121.650 ;
        RECT 40.380 121.310 40.700 121.370 ;
        RECT 38.170 121.170 40.700 121.310 ;
        RECT 40.380 121.110 40.700 121.170 ;
        RECT 41.255 121.150 41.545 121.465 ;
        RECT 46.360 121.450 46.680 121.510 ;
        RECT 42.335 121.310 42.625 121.355 ;
        RECT 45.915 121.310 46.205 121.355 ;
        RECT 47.750 121.310 48.040 121.355 ;
        RECT 42.335 121.170 48.040 121.310 ;
        RECT 42.335 121.125 42.625 121.170 ;
        RECT 45.915 121.125 46.205 121.170 ;
        RECT 47.750 121.125 48.040 121.170 ;
        RECT 48.200 121.110 48.520 121.370 ;
        RECT 49.580 121.310 49.900 121.370 ;
        RECT 55.190 121.355 55.330 121.510 ;
        RECT 61.195 121.510 65.085 121.650 ;
        RECT 61.195 121.465 61.785 121.510 ;
        RECT 50.055 121.310 50.345 121.355 ;
        RECT 49.580 121.170 50.345 121.310 ;
        RECT 49.580 121.110 49.900 121.170 ;
        RECT 50.055 121.125 50.345 121.170 ;
        RECT 52.815 121.125 53.105 121.355 ;
        RECT 55.115 121.125 55.405 121.355 ;
        RECT 27.515 120.970 27.805 121.015 ;
        RECT 30.260 120.970 30.580 121.030 ;
        RECT 27.515 120.830 30.580 120.970 ;
        RECT 27.515 120.785 27.805 120.830 ;
        RECT 30.260 120.770 30.580 120.830 ;
        RECT 36.255 120.970 36.545 121.015 ;
        RECT 38.080 120.970 38.400 121.030 ;
        RECT 36.255 120.830 38.400 120.970 ;
        RECT 36.255 120.785 36.545 120.830 ;
        RECT 38.080 120.770 38.400 120.830 ;
        RECT 46.820 120.770 47.140 121.030 ;
        RECT 52.890 120.970 53.030 121.125 ;
        RECT 55.560 121.110 55.880 121.370 ;
        RECT 61.495 121.150 61.785 121.465 ;
        RECT 62.000 121.450 62.320 121.510 ;
        RECT 64.435 121.465 65.085 121.510 ;
        RECT 67.060 121.450 67.380 121.710 ;
        RECT 68.990 121.355 69.130 121.850 ;
        RECT 69.360 121.850 73.805 121.990 ;
        RECT 69.360 121.790 69.680 121.850 ;
        RECT 73.515 121.805 73.805 121.850 ;
        RECT 76.720 121.990 77.040 122.050 ;
        RECT 76.720 121.850 86.610 121.990 ;
        RECT 76.720 121.790 77.040 121.850 ;
        RECT 72.120 121.650 72.440 121.710 ;
        RECT 70.370 121.510 72.440 121.650 ;
        RECT 70.370 121.355 70.510 121.510 ;
        RECT 72.120 121.450 72.440 121.510 ;
        RECT 75.800 121.650 76.120 121.710 ;
        RECT 77.755 121.650 78.045 121.695 ;
        RECT 80.995 121.650 81.645 121.695 ;
        RECT 75.800 121.510 81.645 121.650 ;
        RECT 75.800 121.450 76.120 121.510 ;
        RECT 77.755 121.465 78.345 121.510 ;
        RECT 80.995 121.465 81.645 121.510 ;
        RECT 62.575 121.310 62.865 121.355 ;
        RECT 66.155 121.310 66.445 121.355 ;
        RECT 67.990 121.310 68.280 121.355 ;
        RECT 62.575 121.170 68.280 121.310 ;
        RECT 62.575 121.125 62.865 121.170 ;
        RECT 66.155 121.125 66.445 121.170 ;
        RECT 67.990 121.125 68.280 121.170 ;
        RECT 68.915 121.125 69.205 121.355 ;
        RECT 70.295 121.125 70.585 121.355 ;
        RECT 71.200 121.310 71.520 121.370 ;
        RECT 71.675 121.310 71.965 121.355 ;
        RECT 71.200 121.170 71.965 121.310 ;
        RECT 71.200 121.110 71.520 121.170 ;
        RECT 71.675 121.125 71.965 121.170 ;
        RECT 73.960 121.110 74.280 121.370 ;
        RECT 78.055 121.150 78.345 121.465 ;
        RECT 83.620 121.450 83.940 121.710 ;
        RECT 84.080 121.650 84.400 121.710 ;
        RECT 84.080 121.510 85.230 121.650 ;
        RECT 84.080 121.450 84.400 121.510 ;
        RECT 85.090 121.355 85.230 121.510 ;
        RECT 86.470 121.355 86.610 121.850 ;
        RECT 88.680 121.650 89.000 121.710 ;
        RECT 90.635 121.650 90.925 121.695 ;
        RECT 93.875 121.650 94.525 121.695 ;
        RECT 88.680 121.510 94.525 121.650 ;
        RECT 88.680 121.450 89.000 121.510 ;
        RECT 90.635 121.465 91.225 121.510 ;
        RECT 93.875 121.465 94.525 121.510 ;
        RECT 79.135 121.310 79.425 121.355 ;
        RECT 82.715 121.310 83.005 121.355 ;
        RECT 84.550 121.310 84.840 121.355 ;
        RECT 79.135 121.170 84.840 121.310 ;
        RECT 79.135 121.125 79.425 121.170 ;
        RECT 82.715 121.125 83.005 121.170 ;
        RECT 84.550 121.125 84.840 121.170 ;
        RECT 85.015 121.125 85.305 121.355 ;
        RECT 86.395 121.125 86.685 121.355 ;
        RECT 90.935 121.150 91.225 121.465 ;
        RECT 96.500 121.450 96.820 121.710 ;
        RECT 97.880 121.450 98.200 121.710 ;
        RECT 98.800 121.650 99.120 121.710 ;
        RECT 102.955 121.650 103.245 121.695 ;
        RECT 98.800 121.510 103.245 121.650 ;
        RECT 98.800 121.450 99.120 121.510 ;
        RECT 102.955 121.465 103.245 121.510 ;
        RECT 105.235 121.650 105.885 121.695 ;
        RECT 108.835 121.650 109.125 121.695 ;
        RECT 109.840 121.650 110.160 121.710 ;
        RECT 105.235 121.510 110.160 121.650 ;
        RECT 105.235 121.465 105.885 121.510 ;
        RECT 108.535 121.465 109.125 121.510 ;
        RECT 92.015 121.310 92.305 121.355 ;
        RECT 95.595 121.310 95.885 121.355 ;
        RECT 97.430 121.310 97.720 121.355 ;
        RECT 92.015 121.170 97.720 121.310 ;
        RECT 97.970 121.310 98.110 121.450 ;
        RECT 99.275 121.310 99.565 121.355 ;
        RECT 97.970 121.170 99.565 121.310 ;
        RECT 92.015 121.125 92.305 121.170 ;
        RECT 95.595 121.125 95.885 121.170 ;
        RECT 97.430 121.125 97.720 121.170 ;
        RECT 99.275 121.125 99.565 121.170 ;
        RECT 101.100 121.310 101.420 121.370 ;
        RECT 101.575 121.310 101.865 121.355 ;
        RECT 101.100 121.170 101.865 121.310 ;
        RECT 101.100 121.110 101.420 121.170 ;
        RECT 101.575 121.125 101.865 121.170 ;
        RECT 102.040 121.310 102.330 121.355 ;
        RECT 103.875 121.310 104.165 121.355 ;
        RECT 107.455 121.310 107.745 121.355 ;
        RECT 102.040 121.170 107.745 121.310 ;
        RECT 102.040 121.125 102.330 121.170 ;
        RECT 103.875 121.125 104.165 121.170 ;
        RECT 107.455 121.125 107.745 121.170 ;
        RECT 108.535 121.150 108.825 121.465 ;
        RECT 109.840 121.450 110.160 121.510 ;
        RECT 56.940 120.970 57.260 121.030 ;
        RECT 52.890 120.830 57.260 120.970 ;
        RECT 56.940 120.770 57.260 120.830 ;
        RECT 58.335 120.970 58.625 121.015 ;
        RECT 60.620 120.970 60.940 121.030 ;
        RECT 58.335 120.830 60.940 120.970 ;
        RECT 58.335 120.785 58.625 120.830 ;
        RECT 60.620 120.770 60.940 120.830 ;
        RECT 61.080 120.970 61.400 121.030 ;
        RECT 68.455 120.970 68.745 121.015 ;
        RECT 61.080 120.830 68.745 120.970 ;
        RECT 61.080 120.770 61.400 120.830 ;
        RECT 68.455 120.785 68.745 120.830 ;
        RECT 74.895 120.970 75.185 121.015 ;
        RECT 75.340 120.970 75.660 121.030 ;
        RECT 74.895 120.830 75.660 120.970 ;
        RECT 74.895 120.785 75.185 120.830 ;
        RECT 75.340 120.770 75.660 120.830 ;
        RECT 87.775 120.785 88.065 121.015 ;
        RECT 97.880 120.970 98.200 121.030 ;
        RECT 101.190 120.970 101.330 121.110 ;
        RECT 97.880 120.830 101.330 120.970 ;
        RECT 106.160 120.970 106.480 121.030 ;
        RECT 111.695 120.970 111.985 121.015 ;
        RECT 106.160 120.830 111.985 120.970 ;
        RECT 31.755 120.630 32.045 120.675 ;
        RECT 34.875 120.630 35.165 120.675 ;
        RECT 36.765 120.630 37.055 120.675 ;
        RECT 31.755 120.490 37.055 120.630 ;
        RECT 31.755 120.445 32.045 120.490 ;
        RECT 34.875 120.445 35.165 120.490 ;
        RECT 36.765 120.445 37.055 120.490 ;
        RECT 42.335 120.630 42.625 120.675 ;
        RECT 45.455 120.630 45.745 120.675 ;
        RECT 47.345 120.630 47.635 120.675 ;
        RECT 42.335 120.490 47.635 120.630 ;
        RECT 42.335 120.445 42.625 120.490 ;
        RECT 45.455 120.445 45.745 120.490 ;
        RECT 47.345 120.445 47.635 120.490 ;
        RECT 62.575 120.630 62.865 120.675 ;
        RECT 65.695 120.630 65.985 120.675 ;
        RECT 67.585 120.630 67.875 120.675 ;
        RECT 62.575 120.490 67.875 120.630 ;
        RECT 62.575 120.445 62.865 120.490 ;
        RECT 65.695 120.445 65.985 120.490 ;
        RECT 67.585 120.445 67.875 120.490 ;
        RECT 79.135 120.630 79.425 120.675 ;
        RECT 82.255 120.630 82.545 120.675 ;
        RECT 84.145 120.630 84.435 120.675 ;
        RECT 79.135 120.490 84.435 120.630 ;
        RECT 87.850 120.630 87.990 120.785 ;
        RECT 97.880 120.770 98.200 120.830 ;
        RECT 106.160 120.770 106.480 120.830 ;
        RECT 111.695 120.785 111.985 120.830 ;
        RECT 90.980 120.630 91.300 120.690 ;
        RECT 87.850 120.490 91.300 120.630 ;
        RECT 79.135 120.445 79.425 120.490 ;
        RECT 82.255 120.445 82.545 120.490 ;
        RECT 84.145 120.445 84.435 120.490 ;
        RECT 90.980 120.430 91.300 120.490 ;
        RECT 92.015 120.630 92.305 120.675 ;
        RECT 95.135 120.630 95.425 120.675 ;
        RECT 97.025 120.630 97.315 120.675 ;
        RECT 92.015 120.490 97.315 120.630 ;
        RECT 92.015 120.445 92.305 120.490 ;
        RECT 95.135 120.445 95.425 120.490 ;
        RECT 97.025 120.445 97.315 120.490 ;
        RECT 102.445 120.630 102.735 120.675 ;
        RECT 104.335 120.630 104.625 120.675 ;
        RECT 107.455 120.630 107.745 120.675 ;
        RECT 102.445 120.490 107.745 120.630 ;
        RECT 102.445 120.445 102.735 120.490 ;
        RECT 104.335 120.445 104.625 120.490 ;
        RECT 107.455 120.445 107.745 120.490 ;
        RECT 49.580 120.290 49.900 120.350 ;
        RECT 52.355 120.290 52.645 120.335 ;
        RECT 49.580 120.150 52.645 120.290 ;
        RECT 49.580 120.090 49.900 120.150 ;
        RECT 52.355 120.105 52.645 120.150 ;
        RECT 54.180 120.090 54.500 120.350 ;
        RECT 69.835 120.290 70.125 120.335 ;
        RECT 70.740 120.290 71.060 120.350 ;
        RECT 69.835 120.150 71.060 120.290 ;
        RECT 69.835 120.105 70.125 120.150 ;
        RECT 70.740 120.090 71.060 120.150 ;
        RECT 71.200 120.090 71.520 120.350 ;
        RECT 72.580 120.090 72.900 120.350 ;
        RECT 87.300 120.090 87.620 120.350 ;
        RECT 98.340 120.090 98.660 120.350 ;
        RECT 22.830 119.470 113.450 119.950 ;
        RECT 37.635 119.270 37.925 119.315 ;
        RECT 38.080 119.270 38.400 119.330 ;
        RECT 106.620 119.270 106.940 119.330 ;
        RECT 37.635 119.130 38.400 119.270 ;
        RECT 37.635 119.085 37.925 119.130 ;
        RECT 38.080 119.070 38.400 119.130 ;
        RECT 86.010 119.130 106.940 119.270 ;
        RECT 26.085 118.930 26.375 118.975 ;
        RECT 27.975 118.930 28.265 118.975 ;
        RECT 31.095 118.930 31.385 118.975 ;
        RECT 26.085 118.790 31.385 118.930 ;
        RECT 26.085 118.745 26.375 118.790 ;
        RECT 27.975 118.745 28.265 118.790 ;
        RECT 31.095 118.745 31.385 118.790 ;
        RECT 36.715 118.930 37.005 118.975 ;
        RECT 39.920 118.930 40.240 118.990 ;
        RECT 36.715 118.790 40.240 118.930 ;
        RECT 36.715 118.745 37.005 118.790 ;
        RECT 39.920 118.730 40.240 118.790 ;
        RECT 41.265 118.930 41.555 118.975 ;
        RECT 43.155 118.930 43.445 118.975 ;
        RECT 46.275 118.930 46.565 118.975 ;
        RECT 54.180 118.930 54.500 118.990 ;
        RECT 41.265 118.790 46.565 118.930 ;
        RECT 41.265 118.745 41.555 118.790 ;
        RECT 43.155 118.745 43.445 118.790 ;
        RECT 46.275 118.745 46.565 118.790 ;
        RECT 50.130 118.790 54.500 118.930 ;
        RECT 26.580 118.590 26.900 118.650 ;
        RECT 37.620 118.590 37.940 118.650 ;
        RECT 40.395 118.590 40.685 118.635 ;
        RECT 26.580 118.450 36.470 118.590 ;
        RECT 26.580 118.390 26.900 118.450 ;
        RECT 25.200 118.050 25.520 118.310 ;
        RECT 36.330 118.295 36.470 118.450 ;
        RECT 37.620 118.450 40.685 118.590 ;
        RECT 37.620 118.390 37.940 118.450 ;
        RECT 40.395 118.405 40.685 118.450 ;
        RECT 41.775 118.590 42.065 118.635 ;
        RECT 50.130 118.590 50.270 118.790 ;
        RECT 54.180 118.730 54.500 118.790 ;
        RECT 55.215 118.930 55.505 118.975 ;
        RECT 58.335 118.930 58.625 118.975 ;
        RECT 60.225 118.930 60.515 118.975 ;
        RECT 55.215 118.790 60.515 118.930 ;
        RECT 55.215 118.745 55.505 118.790 ;
        RECT 58.335 118.745 58.625 118.790 ;
        RECT 60.225 118.745 60.515 118.790 ;
        RECT 66.255 118.930 66.545 118.975 ;
        RECT 69.375 118.930 69.665 118.975 ;
        RECT 71.265 118.930 71.555 118.975 ;
        RECT 66.255 118.790 71.555 118.930 ;
        RECT 66.255 118.745 66.545 118.790 ;
        RECT 69.375 118.745 69.665 118.790 ;
        RECT 71.265 118.745 71.555 118.790 ;
        RECT 76.835 118.930 77.125 118.975 ;
        RECT 79.955 118.930 80.245 118.975 ;
        RECT 81.845 118.930 82.135 118.975 ;
        RECT 84.080 118.930 84.400 118.990 ;
        RECT 76.835 118.790 82.135 118.930 ;
        RECT 76.835 118.745 77.125 118.790 ;
        RECT 79.955 118.745 80.245 118.790 ;
        RECT 81.845 118.745 82.135 118.790 ;
        RECT 82.790 118.790 84.400 118.930 ;
        RECT 41.775 118.450 50.270 118.590 ;
        RECT 41.775 118.405 42.065 118.450 ;
        RECT 50.500 118.390 50.820 118.650 ;
        RECT 59.700 118.390 60.020 118.650 ;
        RECT 70.740 118.390 71.060 118.650 ;
        RECT 72.580 118.590 72.900 118.650 ;
        RECT 81.335 118.590 81.625 118.635 ;
        RECT 72.580 118.450 81.625 118.590 ;
        RECT 72.580 118.390 72.900 118.450 ;
        RECT 81.335 118.405 81.625 118.450 ;
        RECT 25.680 118.250 25.970 118.295 ;
        RECT 27.515 118.250 27.805 118.295 ;
        RECT 31.095 118.250 31.385 118.295 ;
        RECT 25.680 118.110 31.385 118.250 ;
        RECT 25.680 118.065 25.970 118.110 ;
        RECT 27.515 118.065 27.805 118.110 ;
        RECT 31.095 118.065 31.385 118.110 ;
        RECT 32.175 117.955 32.465 118.270 ;
        RECT 36.255 118.250 36.545 118.295 ;
        RECT 37.160 118.250 37.480 118.310 ;
        RECT 36.255 118.110 37.480 118.250 ;
        RECT 36.255 118.065 36.545 118.110 ;
        RECT 37.160 118.050 37.480 118.110 ;
        RECT 38.540 118.050 38.860 118.310 ;
        RECT 39.000 118.250 39.320 118.310 ;
        RECT 39.935 118.250 40.225 118.295 ;
        RECT 39.000 118.110 40.225 118.250 ;
        RECT 39.000 118.050 39.320 118.110 ;
        RECT 39.935 118.065 40.225 118.110 ;
        RECT 40.860 118.250 41.150 118.295 ;
        RECT 42.695 118.250 42.985 118.295 ;
        RECT 46.275 118.250 46.565 118.295 ;
        RECT 40.860 118.110 46.565 118.250 ;
        RECT 40.860 118.065 41.150 118.110 ;
        RECT 42.695 118.065 42.985 118.110 ;
        RECT 46.275 118.065 46.565 118.110 ;
        RECT 26.595 117.725 26.885 117.955 ;
        RECT 28.875 117.910 29.525 117.955 ;
        RECT 32.175 117.910 32.765 117.955 ;
        RECT 34.860 117.910 35.180 117.970 ;
        RECT 28.875 117.770 35.180 117.910 ;
        RECT 28.875 117.725 29.525 117.770 ;
        RECT 32.475 117.725 32.765 117.770 ;
        RECT 26.670 117.570 26.810 117.725 ;
        RECT 34.860 117.710 35.180 117.770 ;
        RECT 35.320 117.710 35.640 117.970 ;
        RECT 47.355 117.955 47.645 118.270 ;
        RECT 44.055 117.910 44.705 117.955 ;
        RECT 47.355 117.910 47.945 117.955 ;
        RECT 49.580 117.910 49.900 117.970 ;
        RECT 54.135 117.955 54.425 118.270 ;
        RECT 55.215 118.250 55.505 118.295 ;
        RECT 58.795 118.250 59.085 118.295 ;
        RECT 60.630 118.250 60.920 118.295 ;
        RECT 55.215 118.110 60.920 118.250 ;
        RECT 55.215 118.065 55.505 118.110 ;
        RECT 58.795 118.065 59.085 118.110 ;
        RECT 60.630 118.065 60.920 118.110 ;
        RECT 61.080 118.050 61.400 118.310 ;
        RECT 65.220 118.270 65.540 118.310 ;
        RECT 82.790 118.295 82.930 118.790 ;
        RECT 84.080 118.730 84.400 118.790 ;
        RECT 65.175 118.050 65.540 118.270 ;
        RECT 66.255 118.250 66.545 118.295 ;
        RECT 69.835 118.250 70.125 118.295 ;
        RECT 71.670 118.250 71.960 118.295 ;
        RECT 66.255 118.110 71.960 118.250 ;
        RECT 66.255 118.065 66.545 118.110 ;
        RECT 69.835 118.065 70.125 118.110 ;
        RECT 71.670 118.065 71.960 118.110 ;
        RECT 72.135 118.065 72.425 118.295 ;
        RECT 57.400 117.955 57.720 117.970 ;
        RECT 65.175 117.955 65.465 118.050 ;
        RECT 44.055 117.770 49.900 117.910 ;
        RECT 44.055 117.725 44.705 117.770 ;
        RECT 47.655 117.725 47.945 117.770 ;
        RECT 49.580 117.710 49.900 117.770 ;
        RECT 50.975 117.725 51.265 117.955 ;
        RECT 53.835 117.910 54.425 117.955 ;
        RECT 57.075 117.910 57.725 117.955 ;
        RECT 53.835 117.770 57.725 117.910 ;
        RECT 53.835 117.725 54.125 117.770 ;
        RECT 57.075 117.725 57.725 117.770 ;
        RECT 62.015 117.725 62.305 117.955 ;
        RECT 64.875 117.910 65.465 117.955 ;
        RECT 68.115 117.910 68.765 117.955 ;
        RECT 64.875 117.770 68.765 117.910 ;
        RECT 64.875 117.725 65.165 117.770 ;
        RECT 68.115 117.725 68.765 117.770 ;
        RECT 39.015 117.570 39.305 117.615 ;
        RECT 26.670 117.430 39.305 117.570 ;
        RECT 51.050 117.570 51.190 117.725 ;
        RECT 57.400 117.710 57.720 117.725 ;
        RECT 55.560 117.570 55.880 117.630 ;
        RECT 51.050 117.430 55.880 117.570 ;
        RECT 62.090 117.570 62.230 117.725 ;
        RECT 65.680 117.570 66.000 117.630 ;
        RECT 62.090 117.430 66.000 117.570 ;
        RECT 72.210 117.570 72.350 118.065 ;
        RECT 72.580 117.710 72.900 117.970 ;
        RECT 73.500 117.910 73.820 117.970 ;
        RECT 75.755 117.955 76.045 118.270 ;
        RECT 76.835 118.250 77.125 118.295 ;
        RECT 80.415 118.250 80.705 118.295 ;
        RECT 82.250 118.250 82.540 118.295 ;
        RECT 76.835 118.110 82.540 118.250 ;
        RECT 76.835 118.065 77.125 118.110 ;
        RECT 80.415 118.065 80.705 118.110 ;
        RECT 82.250 118.065 82.540 118.110 ;
        RECT 82.715 118.065 83.005 118.295 ;
        RECT 84.080 118.250 84.400 118.310 ;
        RECT 86.010 118.295 86.150 119.130 ;
        RECT 106.620 119.070 106.940 119.130 ;
        RECT 109.395 119.270 109.685 119.315 ;
        RECT 109.840 119.270 110.160 119.330 ;
        RECT 109.395 119.130 110.160 119.270 ;
        RECT 109.395 119.085 109.685 119.130 ;
        RECT 109.840 119.070 110.160 119.130 ;
        RECT 92.015 118.930 92.305 118.975 ;
        RECT 95.135 118.930 95.425 118.975 ;
        RECT 97.025 118.930 97.315 118.975 ;
        RECT 92.015 118.790 97.315 118.930 ;
        RECT 92.015 118.745 92.305 118.790 ;
        RECT 95.135 118.745 95.425 118.790 ;
        RECT 97.025 118.745 97.315 118.790 ;
        RECT 99.225 118.930 99.515 118.975 ;
        RECT 101.115 118.930 101.405 118.975 ;
        RECT 104.235 118.930 104.525 118.975 ;
        RECT 99.225 118.790 104.525 118.930 ;
        RECT 99.225 118.745 99.515 118.790 ;
        RECT 101.115 118.745 101.405 118.790 ;
        RECT 104.235 118.745 104.525 118.790 ;
        RECT 87.300 118.590 87.620 118.650 ;
        RECT 96.515 118.590 96.805 118.635 ;
        RECT 87.300 118.450 96.805 118.590 ;
        RECT 87.300 118.390 87.620 118.450 ;
        RECT 96.515 118.405 96.805 118.450 ;
        RECT 97.880 118.590 98.200 118.650 ;
        RECT 98.355 118.590 98.645 118.635 ;
        RECT 97.880 118.450 98.645 118.590 ;
        RECT 97.880 118.390 98.200 118.450 ;
        RECT 98.355 118.405 98.645 118.450 ;
        RECT 99.720 118.390 100.040 118.650 ;
        RECT 84.555 118.250 84.845 118.295 ;
        RECT 85.935 118.250 86.225 118.295 ;
        RECT 84.080 118.110 86.225 118.250 ;
        RECT 75.455 117.910 76.045 117.955 ;
        RECT 78.695 117.910 79.345 117.955 ;
        RECT 73.500 117.770 79.345 117.910 ;
        RECT 73.500 117.710 73.820 117.770 ;
        RECT 75.455 117.725 75.745 117.770 ;
        RECT 78.695 117.725 79.345 117.770 ;
        RECT 76.720 117.570 77.040 117.630 ;
        RECT 82.790 117.570 82.930 118.065 ;
        RECT 84.080 118.050 84.400 118.110 ;
        RECT 84.555 118.065 84.845 118.110 ;
        RECT 85.935 118.065 86.225 118.110 ;
        RECT 86.840 118.250 87.160 118.310 ;
        RECT 87.775 118.250 88.065 118.295 ;
        RECT 86.840 118.110 88.065 118.250 ;
        RECT 86.840 118.050 87.160 118.110 ;
        RECT 87.775 118.065 88.065 118.110 ;
        RECT 90.935 117.955 91.225 118.270 ;
        RECT 92.015 118.250 92.305 118.295 ;
        RECT 95.595 118.250 95.885 118.295 ;
        RECT 97.430 118.250 97.720 118.295 ;
        RECT 92.015 118.110 97.720 118.250 ;
        RECT 92.015 118.065 92.305 118.110 ;
        RECT 95.595 118.065 95.885 118.110 ;
        RECT 97.430 118.065 97.720 118.110 ;
        RECT 98.820 118.250 99.110 118.295 ;
        RECT 100.655 118.250 100.945 118.295 ;
        RECT 104.235 118.250 104.525 118.295 ;
        RECT 98.820 118.110 104.525 118.250 ;
        RECT 98.820 118.065 99.110 118.110 ;
        RECT 100.655 118.065 100.945 118.110 ;
        RECT 104.235 118.065 104.525 118.110 ;
        RECT 102.020 117.955 102.340 117.970 ;
        RECT 105.315 117.955 105.605 118.270 ;
        RECT 106.620 118.250 106.940 118.310 ;
        RECT 109.855 118.250 110.145 118.295 ;
        RECT 110.315 118.250 110.605 118.295 ;
        RECT 106.620 118.110 110.605 118.250 ;
        RECT 106.620 118.050 106.940 118.110 ;
        RECT 109.855 118.065 110.145 118.110 ;
        RECT 110.315 118.065 110.605 118.110 ;
        RECT 86.395 117.910 86.685 117.955 ;
        RECT 90.635 117.910 91.225 117.955 ;
        RECT 93.875 117.910 94.525 117.955 ;
        RECT 86.395 117.770 94.525 117.910 ;
        RECT 86.395 117.725 86.685 117.770 ;
        RECT 90.635 117.725 90.925 117.770 ;
        RECT 93.875 117.725 94.525 117.770 ;
        RECT 102.015 117.910 102.665 117.955 ;
        RECT 105.315 117.910 105.905 117.955 ;
        RECT 102.015 117.770 105.905 117.910 ;
        RECT 102.015 117.725 102.665 117.770 ;
        RECT 105.615 117.725 105.905 117.770 ;
        RECT 108.475 117.725 108.765 117.955 ;
        RECT 102.020 117.710 102.340 117.725 ;
        RECT 72.210 117.430 82.930 117.570 ;
        RECT 39.015 117.385 39.305 117.430 ;
        RECT 55.560 117.370 55.880 117.430 ;
        RECT 65.680 117.370 66.000 117.430 ;
        RECT 76.720 117.370 77.040 117.430 ;
        RECT 83.620 117.370 83.940 117.630 ;
        RECT 85.000 117.370 85.320 117.630 ;
        RECT 101.100 117.570 101.420 117.630 ;
        RECT 108.550 117.570 108.690 117.725 ;
        RECT 101.100 117.430 108.690 117.570 ;
        RECT 101.100 117.370 101.420 117.430 ;
        RECT 110.760 117.370 111.080 117.630 ;
        RECT 22.830 116.750 113.450 117.230 ;
        RECT 34.860 116.550 35.180 116.610 ;
        RECT 36.715 116.550 37.005 116.595 ;
        RECT 34.860 116.410 37.005 116.550 ;
        RECT 34.860 116.350 35.180 116.410 ;
        RECT 36.715 116.365 37.005 116.410 ;
        RECT 37.635 116.365 37.925 116.595 ;
        RECT 27.155 116.210 27.445 116.255 ;
        RECT 30.395 116.210 31.045 116.255 ;
        RECT 27.155 116.070 31.045 116.210 ;
        RECT 27.155 116.025 27.745 116.070 ;
        RECT 30.395 116.025 31.045 116.070 ;
        RECT 33.035 116.210 33.325 116.255 ;
        RECT 37.710 116.210 37.850 116.365 ;
        RECT 44.980 116.350 45.300 116.610 ;
        RECT 46.820 116.350 47.140 116.610 ;
        RECT 57.400 116.550 57.720 116.610 ;
        RECT 57.875 116.550 58.165 116.595 ;
        RECT 57.400 116.410 58.165 116.550 ;
        RECT 57.400 116.350 57.720 116.410 ;
        RECT 57.875 116.365 58.165 116.410 ;
        RECT 62.000 116.550 62.320 116.610 ;
        RECT 62.475 116.550 62.765 116.595 ;
        RECT 62.000 116.410 62.765 116.550 ;
        RECT 62.000 116.350 62.320 116.410 ;
        RECT 62.475 116.365 62.765 116.410 ;
        RECT 64.315 116.550 64.605 116.595 ;
        RECT 65.220 116.550 65.540 116.610 ;
        RECT 64.315 116.410 65.540 116.550 ;
        RECT 64.315 116.365 64.605 116.410 ;
        RECT 65.220 116.350 65.540 116.410 ;
        RECT 73.500 116.350 73.820 116.610 ;
        RECT 75.800 116.350 76.120 116.610 ;
        RECT 88.680 116.350 89.000 116.610 ;
        RECT 97.420 116.550 97.740 116.610 ;
        RECT 97.420 116.410 103.170 116.550 ;
        RECT 97.420 116.350 97.740 116.410 ;
        RECT 56.940 116.210 57.260 116.270 ;
        RECT 33.035 116.070 37.850 116.210 ;
        RECT 44.610 116.070 57.260 116.210 ;
        RECT 33.035 116.025 33.325 116.070 ;
        RECT 27.455 115.710 27.745 116.025 ;
        RECT 28.535 115.870 28.825 115.915 ;
        RECT 32.115 115.870 32.405 115.915 ;
        RECT 33.950 115.870 34.240 115.915 ;
        RECT 28.535 115.730 34.240 115.870 ;
        RECT 24.295 115.530 24.585 115.575 ;
        RECT 25.200 115.530 25.520 115.590 ;
        RECT 24.295 115.390 25.520 115.530 ;
        RECT 27.590 115.530 27.730 115.710 ;
        RECT 28.535 115.685 28.825 115.730 ;
        RECT 32.115 115.685 32.405 115.730 ;
        RECT 33.950 115.685 34.240 115.730 ;
        RECT 37.160 115.870 37.480 115.930 ;
        RECT 37.160 115.730 38.310 115.870 ;
        RECT 37.160 115.670 37.480 115.730 ;
        RECT 34.415 115.530 34.705 115.575 ;
        RECT 37.620 115.530 37.940 115.590 ;
        RECT 27.590 115.390 34.170 115.530 ;
        RECT 24.295 115.345 24.585 115.390 ;
        RECT 25.200 115.330 25.520 115.390 ;
        RECT 28.535 115.190 28.825 115.235 ;
        RECT 31.655 115.190 31.945 115.235 ;
        RECT 33.545 115.190 33.835 115.235 ;
        RECT 28.535 115.050 33.835 115.190 ;
        RECT 34.030 115.190 34.170 115.390 ;
        RECT 34.415 115.390 37.940 115.530 ;
        RECT 38.170 115.530 38.310 115.730 ;
        RECT 38.540 115.670 38.860 115.930 ;
        RECT 44.610 115.915 44.750 116.070 ;
        RECT 56.800 116.010 57.260 116.070 ;
        RECT 71.200 116.210 71.520 116.270 ;
        RECT 78.115 116.210 78.405 116.255 ;
        RECT 71.200 116.070 78.405 116.210 ;
        RECT 71.200 116.010 71.520 116.070 ;
        RECT 78.115 116.025 78.405 116.070 ;
        RECT 80.395 116.210 81.045 116.255 ;
        RECT 83.995 116.210 84.285 116.255 ;
        RECT 80.395 116.070 84.285 116.210 ;
        RECT 80.395 116.025 81.045 116.070 ;
        RECT 83.695 116.025 84.285 116.070 ;
        RECT 85.000 116.210 85.320 116.270 ;
        RECT 92.475 116.210 92.765 116.255 ;
        RECT 95.715 116.210 96.365 116.255 ;
        RECT 85.000 116.070 96.365 116.210 ;
        RECT 39.935 115.870 40.225 115.915 ;
        RECT 41.315 115.870 41.605 115.915 ;
        RECT 44.535 115.870 44.825 115.915 ;
        RECT 39.935 115.730 44.825 115.870 ;
        RECT 39.935 115.685 40.225 115.730 ;
        RECT 41.315 115.685 41.605 115.730 ;
        RECT 44.535 115.685 44.825 115.730 ;
        RECT 45.440 115.870 45.760 115.930 ;
        RECT 45.915 115.870 46.205 115.915 ;
        RECT 45.440 115.730 46.205 115.870 ;
        RECT 56.800 115.870 56.940 116.010 ;
        RECT 83.695 115.930 83.985 116.025 ;
        RECT 85.000 116.010 85.320 116.070 ;
        RECT 92.475 116.025 93.065 116.070 ;
        RECT 95.715 116.025 96.365 116.070 ;
        RECT 58.335 115.870 58.625 115.915 ;
        RECT 62.015 115.870 62.305 115.915 ;
        RECT 63.855 115.870 64.145 115.915 ;
        RECT 56.800 115.730 64.145 115.870 ;
        RECT 40.010 115.530 40.150 115.685 ;
        RECT 45.440 115.670 45.760 115.730 ;
        RECT 45.915 115.685 46.205 115.730 ;
        RECT 58.335 115.685 58.625 115.730 ;
        RECT 62.015 115.685 62.305 115.730 ;
        RECT 63.855 115.685 64.145 115.730 ;
        RECT 73.975 115.870 74.265 115.915 ;
        RECT 75.355 115.870 75.645 115.915 ;
        RECT 73.975 115.730 75.645 115.870 ;
        RECT 73.975 115.685 74.265 115.730 ;
        RECT 75.355 115.685 75.645 115.730 ;
        RECT 38.170 115.390 40.150 115.530 ;
        RECT 34.415 115.345 34.705 115.390 ;
        RECT 37.620 115.330 37.940 115.390 ;
        RECT 40.855 115.190 41.145 115.235 ;
        RECT 34.030 115.050 41.145 115.190 ;
        RECT 28.535 115.005 28.825 115.050 ;
        RECT 31.655 115.005 31.945 115.050 ;
        RECT 33.545 115.005 33.835 115.050 ;
        RECT 40.855 115.005 41.145 115.050 ;
        RECT 35.780 114.850 36.100 114.910 ;
        RECT 39.475 114.850 39.765 114.895 ;
        RECT 35.780 114.710 39.765 114.850 ;
        RECT 75.430 114.850 75.570 115.685 ;
        RECT 76.720 115.670 77.040 115.930 ;
        RECT 77.200 115.870 77.490 115.915 ;
        RECT 79.035 115.870 79.325 115.915 ;
        RECT 82.615 115.870 82.905 115.915 ;
        RECT 77.200 115.730 82.905 115.870 ;
        RECT 77.200 115.685 77.490 115.730 ;
        RECT 79.035 115.685 79.325 115.730 ;
        RECT 82.615 115.685 82.905 115.730 ;
        RECT 83.620 115.710 83.985 115.930 ;
        RECT 84.540 115.870 84.860 115.930 ;
        RECT 88.235 115.870 88.525 115.915 ;
        RECT 84.540 115.730 88.525 115.870 ;
        RECT 83.620 115.670 83.940 115.710 ;
        RECT 84.540 115.670 84.860 115.730 ;
        RECT 88.235 115.685 88.525 115.730 ;
        RECT 92.775 115.710 93.065 116.025 ;
        RECT 98.340 116.010 98.660 116.270 ;
        RECT 103.030 116.255 103.170 116.410 ;
        RECT 102.955 116.025 103.245 116.255 ;
        RECT 105.235 116.210 105.885 116.255 ;
        RECT 108.835 116.210 109.125 116.255 ;
        RECT 110.760 116.210 111.080 116.270 ;
        RECT 105.235 116.070 111.080 116.210 ;
        RECT 105.235 116.025 105.885 116.070 ;
        RECT 108.535 116.025 109.125 116.070 ;
        RECT 93.855 115.870 94.145 115.915 ;
        RECT 97.435 115.870 97.725 115.915 ;
        RECT 99.270 115.870 99.560 115.915 ;
        RECT 93.855 115.730 99.560 115.870 ;
        RECT 93.855 115.685 94.145 115.730 ;
        RECT 97.435 115.685 97.725 115.730 ;
        RECT 99.270 115.685 99.560 115.730 ;
        RECT 102.040 115.870 102.330 115.915 ;
        RECT 103.875 115.870 104.165 115.915 ;
        RECT 107.455 115.870 107.745 115.915 ;
        RECT 102.040 115.730 107.745 115.870 ;
        RECT 102.040 115.685 102.330 115.730 ;
        RECT 103.875 115.685 104.165 115.730 ;
        RECT 107.455 115.685 107.745 115.730 ;
        RECT 108.535 115.710 108.825 116.025 ;
        RECT 110.760 116.010 111.080 116.070 ;
        RECT 80.860 115.530 81.180 115.590 ;
        RECT 86.855 115.530 87.145 115.575 ;
        RECT 80.860 115.390 87.145 115.530 ;
        RECT 80.860 115.330 81.180 115.390 ;
        RECT 86.855 115.345 87.145 115.390 ;
        RECT 89.615 115.530 89.905 115.575 ;
        RECT 96.040 115.530 96.360 115.590 ;
        RECT 89.615 115.390 96.360 115.530 ;
        RECT 89.615 115.345 89.905 115.390 ;
        RECT 96.040 115.330 96.360 115.390 ;
        RECT 97.880 115.530 98.200 115.590 ;
        RECT 99.735 115.530 100.025 115.575 ;
        RECT 101.575 115.530 101.865 115.575 ;
        RECT 97.880 115.390 101.865 115.530 ;
        RECT 97.880 115.330 98.200 115.390 ;
        RECT 99.735 115.345 100.025 115.390 ;
        RECT 101.575 115.345 101.865 115.390 ;
        RECT 111.680 115.330 112.000 115.590 ;
        RECT 77.605 115.190 77.895 115.235 ;
        RECT 79.495 115.190 79.785 115.235 ;
        RECT 82.615 115.190 82.905 115.235 ;
        RECT 77.605 115.050 82.905 115.190 ;
        RECT 77.605 115.005 77.895 115.050 ;
        RECT 79.495 115.005 79.785 115.050 ;
        RECT 82.615 115.005 82.905 115.050 ;
        RECT 93.855 115.190 94.145 115.235 ;
        RECT 96.975 115.190 97.265 115.235 ;
        RECT 98.865 115.190 99.155 115.235 ;
        RECT 93.855 115.050 99.155 115.190 ;
        RECT 93.855 115.005 94.145 115.050 ;
        RECT 96.975 115.005 97.265 115.050 ;
        RECT 98.865 115.005 99.155 115.050 ;
        RECT 102.445 115.190 102.735 115.235 ;
        RECT 104.335 115.190 104.625 115.235 ;
        RECT 107.455 115.190 107.745 115.235 ;
        RECT 102.445 115.050 107.745 115.190 ;
        RECT 102.445 115.005 102.735 115.050 ;
        RECT 104.335 115.005 104.625 115.050 ;
        RECT 107.455 115.005 107.745 115.050 ;
        RECT 79.940 114.850 80.260 114.910 ;
        RECT 84.080 114.850 84.400 114.910 ;
        RECT 75.430 114.710 84.400 114.850 ;
        RECT 35.780 114.650 36.100 114.710 ;
        RECT 39.475 114.665 39.765 114.710 ;
        RECT 79.940 114.650 80.260 114.710 ;
        RECT 84.080 114.650 84.400 114.710 ;
        RECT 22.830 114.030 113.450 114.510 ;
        RECT 135.660 106.690 136.800 133.400 ;
        RECT 133.100 106.600 136.850 106.690 ;
        RECT 129.700 105.630 136.850 106.600 ;
        RECT 133.100 105.500 136.850 105.630 ;
        RECT 133.330 76.630 136.060 77.830 ;
        RECT 137.920 77.810 143.450 77.960 ;
        RECT 21.115 74.380 23.065 74.390 ;
        RECT 19.415 73.240 23.065 74.380 ;
        RECT 19.415 73.230 21.125 73.240 ;
        RECT 28.135 73.230 30.305 74.410 ;
        RECT 32.315 74.390 34.265 74.400 ;
        RECT 30.615 73.250 34.265 74.390 ;
        RECT 30.615 73.240 32.325 73.250 ;
        RECT 39.425 73.200 41.595 74.380 ;
        RECT 43.535 74.360 45.485 74.370 ;
        RECT 41.835 73.220 45.485 74.360 ;
        RECT 54.785 74.340 56.735 74.350 ;
        RECT 41.835 73.210 43.545 73.220 ;
        RECT 3.910 73.080 6.100 73.190 ;
        RECT 50.005 73.140 52.175 74.320 ;
        RECT 53.085 73.200 56.735 74.340 ;
        RECT 53.085 73.190 54.795 73.200 ;
        RECT 61.425 73.170 63.595 74.350 ;
        RECT 66.005 74.330 67.955 74.340 ;
        RECT 64.305 73.190 67.955 74.330 ;
        RECT 64.305 73.180 66.015 73.190 ;
        RECT 72.535 73.180 74.705 74.360 ;
        RECT 77.245 74.320 79.195 74.330 ;
        RECT 75.545 73.180 79.195 74.320 ;
        RECT 75.545 73.170 77.255 73.180 ;
        RECT 83.805 73.170 85.975 74.350 ;
        RECT 88.495 74.330 90.445 74.340 ;
        RECT 86.795 73.190 90.445 74.330 ;
        RECT 99.775 74.320 101.725 74.330 ;
        RECT 86.795 73.180 88.505 73.190 ;
        RECT 94.995 73.110 97.165 74.290 ;
        RECT 98.075 73.180 101.725 74.320 ;
        RECT 98.075 73.170 99.785 73.180 ;
        RECT 106.405 73.160 108.575 74.340 ;
        RECT 111.045 74.320 112.995 74.330 ;
        RECT 109.345 73.180 112.995 74.320 ;
        RECT 109.345 73.170 111.055 73.180 ;
        RECT 117.605 73.160 119.775 74.340 ;
        RECT 122.295 74.320 124.245 74.330 ;
        RECT 120.595 73.180 124.245 74.320 ;
        RECT 129.455 73.240 131.625 74.420 ;
        RECT 120.595 73.170 122.305 73.180 ;
        RECT 3.910 72.820 12.240 73.080 ;
        RECT 29.635 72.840 43.235 72.850 ;
        RECT 18.435 72.820 43.235 72.840 ;
        RECT 3.910 72.800 54.455 72.820 ;
        RECT 3.910 72.790 65.705 72.800 ;
        RECT 133.960 72.790 135.640 76.630 ;
        RECT 137.190 76.610 143.450 77.810 ;
        RECT 137.920 75.460 143.450 76.610 ;
        RECT 3.910 72.780 76.925 72.790 ;
        RECT 85.815 72.780 99.415 72.790 ;
        RECT 132.085 72.780 140.600 72.790 ;
        RECT 3.910 71.700 140.600 72.780 ;
        RECT 3.910 71.690 32.035 71.700 ;
        RECT 3.910 71.670 19.135 71.690 ;
        RECT 40.855 71.670 140.600 71.700 ;
        RECT 3.910 71.500 12.240 71.670 ;
        RECT 52.105 71.650 140.600 71.670 ;
        RECT 63.325 71.640 140.600 71.650 ;
        RECT 74.565 71.630 88.165 71.640 ;
        RECT 97.095 71.630 133.215 71.640 ;
        RECT 3.910 71.370 6.100 71.500 ;
        RECT 10.800 71.180 11.950 71.500 ;
        RECT 10.800 69.480 11.915 71.180 ;
        RECT 29.635 71.170 43.285 71.180 ;
        RECT 15.510 71.155 17.040 71.160 ;
        RECT 18.435 71.155 43.285 71.170 ;
        RECT 12.285 71.150 43.285 71.155 ;
        RECT 12.285 71.130 54.505 71.150 ;
        RECT 141.810 71.140 143.230 75.460 ;
        RECT 12.285 71.120 65.755 71.130 ;
        RECT 12.285 71.110 76.975 71.120 ;
        RECT 85.815 71.110 99.465 71.120 ;
        RECT 140.220 71.110 143.240 71.140 ;
        RECT 12.285 70.030 143.240 71.110 ;
        RECT 12.285 70.020 32.085 70.030 ;
        RECT 12.285 70.005 19.375 70.020 ;
        RECT 10.800 13.800 11.950 69.480 ;
        RECT 12.320 15.450 13.470 70.005 ;
        RECT 15.510 68.660 17.040 70.005 ;
        RECT 40.855 70.000 143.240 70.030 ;
        RECT 52.105 69.980 143.240 70.000 ;
        RECT 63.325 69.970 143.240 69.980 ;
        RECT 74.565 69.960 88.215 69.970 ;
        RECT 97.095 69.960 143.240 69.970 ;
        RECT 140.220 69.910 143.240 69.960 ;
        RECT 29.645 69.670 43.315 69.680 ;
        RECT 18.445 69.650 43.315 69.670 ;
        RECT 18.445 69.630 54.535 69.650 ;
        RECT 18.445 69.620 65.785 69.630 ;
        RECT 139.590 69.620 150.610 69.640 ;
        RECT 18.445 69.610 77.005 69.620 ;
        RECT 85.825 69.610 99.495 69.620 ;
        RECT 132.155 69.610 150.610 69.620 ;
        RECT 18.445 69.570 150.610 69.610 ;
        RECT 18.445 68.530 150.740 69.570 ;
        RECT 18.445 68.520 32.115 68.530 ;
        RECT 40.865 68.500 150.740 68.530 ;
        RECT 52.115 68.490 143.320 68.500 ;
        RECT 52.115 68.480 140.670 68.490 ;
        RECT 63.335 68.470 140.670 68.480 ;
        RECT 74.575 68.460 88.245 68.470 ;
        RECT 97.105 68.460 133.295 68.470 ;
        RECT 141.080 68.450 142.300 68.490 ;
        RECT 149.360 68.470 150.740 68.500 ;
        RECT 29.655 68.100 43.325 68.110 ;
        RECT 13.950 68.080 43.325 68.100 ;
        RECT 13.950 68.060 54.545 68.080 ;
        RECT 13.950 68.050 65.795 68.060 ;
        RECT 13.950 68.040 77.015 68.050 ;
        RECT 85.835 68.040 99.505 68.050 ;
        RECT 139.530 68.040 143.320 68.060 ;
        RECT 13.950 66.960 152.870 68.040 ;
        RECT 13.950 66.950 32.125 66.960 ;
        RECT 13.950 18.530 15.100 66.950 ;
        RECT 40.875 66.930 152.870 66.960 ;
        RECT 52.125 66.910 152.870 66.930 ;
        RECT 63.345 66.900 152.870 66.910 ;
        RECT 74.585 66.890 88.255 66.900 ;
        RECT 97.115 66.890 143.320 66.900 ;
        RECT 141.030 66.770 142.490 66.890 ;
        RECT 21.405 65.510 26.555 65.790 ;
        RECT 27.815 65.490 28.965 65.800 ;
        RECT 32.605 65.520 37.755 65.800 ;
        RECT 39.015 65.500 40.165 65.810 ;
        RECT 43.825 65.490 48.975 65.770 ;
        RECT 50.235 65.470 51.385 65.780 ;
        RECT 149.460 65.760 150.600 65.780 ;
        RECT 55.075 65.470 60.225 65.750 ;
        RECT 61.485 65.450 62.635 65.760 ;
        RECT 66.295 65.460 71.445 65.740 ;
        RECT 72.705 65.440 73.855 65.750 ;
        RECT 77.535 65.450 82.685 65.730 ;
        RECT 83.945 65.430 85.095 65.740 ;
        RECT 88.785 65.460 93.935 65.740 ;
        RECT 95.195 65.440 96.345 65.750 ;
        RECT 100.065 65.450 105.215 65.730 ;
        RECT 106.475 65.430 107.625 65.740 ;
        RECT 111.335 65.450 116.485 65.730 ;
        RECT 117.745 65.430 118.895 65.740 ;
        RECT 122.585 65.450 127.735 65.730 ;
        RECT 128.995 65.430 130.145 65.740 ;
        RECT 133.315 65.430 138.455 65.690 ;
        RECT 21.205 65.140 21.435 65.320 ;
        RECT 26.495 65.190 26.725 65.320 ;
        RECT 21.125 55.220 21.485 65.140 ;
        RECT 26.435 55.240 26.805 65.190 ;
        RECT 27.635 65.150 27.865 65.320 ;
        RECT 27.565 55.200 27.935 65.150 ;
        RECT 28.925 65.140 29.155 65.320 ;
        RECT 32.405 65.150 32.635 65.330 ;
        RECT 37.695 65.200 37.925 65.330 ;
        RECT 28.835 55.250 29.255 65.140 ;
        RECT 32.325 55.230 32.685 65.150 ;
        RECT 37.635 55.250 38.005 65.200 ;
        RECT 38.835 65.160 39.065 65.330 ;
        RECT 38.765 55.210 39.135 65.160 ;
        RECT 40.125 65.150 40.355 65.330 ;
        RECT 40.035 55.260 40.455 65.150 ;
        RECT 43.625 65.120 43.855 65.300 ;
        RECT 48.915 65.170 49.145 65.300 ;
        RECT 43.545 55.200 43.905 65.120 ;
        RECT 48.855 55.220 49.225 65.170 ;
        RECT 50.055 65.130 50.285 65.300 ;
        RECT 49.985 55.180 50.355 65.130 ;
        RECT 51.345 65.120 51.575 65.300 ;
        RECT 51.255 55.230 51.675 65.120 ;
        RECT 54.875 65.100 55.105 65.280 ;
        RECT 60.165 65.150 60.395 65.280 ;
        RECT 54.795 55.180 55.155 65.100 ;
        RECT 60.105 55.200 60.475 65.150 ;
        RECT 61.305 65.110 61.535 65.280 ;
        RECT 61.235 55.160 61.605 65.110 ;
        RECT 62.595 65.100 62.825 65.280 ;
        RECT 62.505 55.210 62.925 65.100 ;
        RECT 66.095 65.090 66.325 65.270 ;
        RECT 71.385 65.140 71.615 65.270 ;
        RECT 66.015 55.170 66.375 65.090 ;
        RECT 71.325 55.190 71.695 65.140 ;
        RECT 72.525 65.100 72.755 65.270 ;
        RECT 72.455 55.150 72.825 65.100 ;
        RECT 73.815 65.090 74.045 65.270 ;
        RECT 73.725 55.200 74.145 65.090 ;
        RECT 77.335 65.080 77.565 65.260 ;
        RECT 82.625 65.130 82.855 65.260 ;
        RECT 77.255 55.160 77.615 65.080 ;
        RECT 82.565 55.180 82.935 65.130 ;
        RECT 83.765 65.090 83.995 65.260 ;
        RECT 83.695 55.140 84.065 65.090 ;
        RECT 85.055 65.080 85.285 65.260 ;
        RECT 88.585 65.090 88.815 65.270 ;
        RECT 93.875 65.140 94.105 65.270 ;
        RECT 84.965 55.190 85.385 65.080 ;
        RECT 88.505 55.170 88.865 65.090 ;
        RECT 93.815 55.190 94.185 65.140 ;
        RECT 95.015 65.100 95.245 65.270 ;
        RECT 94.945 55.150 95.315 65.100 ;
        RECT 96.305 65.090 96.535 65.270 ;
        RECT 96.215 55.200 96.635 65.090 ;
        RECT 99.865 65.080 100.095 65.260 ;
        RECT 105.155 65.130 105.385 65.260 ;
        RECT 99.785 55.160 100.145 65.080 ;
        RECT 105.095 55.180 105.465 65.130 ;
        RECT 106.295 65.090 106.525 65.260 ;
        RECT 106.225 55.140 106.595 65.090 ;
        RECT 107.585 65.080 107.815 65.260 ;
        RECT 111.135 65.080 111.365 65.260 ;
        RECT 116.425 65.130 116.655 65.260 ;
        RECT 107.495 55.190 107.915 65.080 ;
        RECT 111.055 55.160 111.415 65.080 ;
        RECT 116.365 55.180 116.735 65.130 ;
        RECT 117.565 65.090 117.795 65.260 ;
        RECT 117.495 55.140 117.865 65.090 ;
        RECT 118.855 65.080 119.085 65.260 ;
        RECT 122.385 65.080 122.615 65.260 ;
        RECT 127.675 65.130 127.905 65.260 ;
        RECT 118.765 55.190 119.185 65.080 ;
        RECT 122.305 55.160 122.665 65.080 ;
        RECT 127.615 55.180 127.985 65.130 ;
        RECT 128.815 65.090 129.045 65.260 ;
        RECT 128.745 55.140 129.115 65.090 ;
        RECT 130.105 65.080 130.335 65.260 ;
        RECT 133.135 65.130 133.365 65.230 ;
        RECT 130.015 55.190 130.435 65.080 ;
        RECT 133.005 55.240 133.405 65.130 ;
        RECT 138.425 65.100 138.655 65.230 ;
        RECT 133.135 55.230 133.365 55.240 ;
        RECT 138.345 55.130 138.725 65.100 ;
        RECT 149.340 64.660 150.720 65.760 ;
        RECT 20.815 54.230 25.555 54.530 ;
        RECT 32.015 54.240 36.755 54.540 ;
        RECT 43.235 54.210 47.975 54.510 ;
        RECT 54.485 54.190 59.225 54.490 ;
        RECT 65.705 54.180 70.445 54.480 ;
        RECT 76.945 54.170 81.685 54.470 ;
        RECT 88.195 54.180 92.935 54.480 ;
        RECT 99.475 54.170 104.215 54.470 ;
        RECT 110.745 54.170 115.485 54.470 ;
        RECT 121.995 54.170 126.735 54.470 ;
        RECT 21.655 52.320 22.115 52.550 ;
        RECT 25.625 52.280 26.255 52.560 ;
        RECT 25.735 52.240 26.195 52.280 ;
        RECT 27.665 52.240 28.125 52.470 ;
        RECT 32.855 52.330 33.315 52.560 ;
        RECT 36.825 52.290 37.455 52.570 ;
        RECT 36.935 52.250 37.395 52.290 ;
        RECT 38.865 52.250 39.325 52.480 ;
        RECT 44.075 52.300 44.535 52.530 ;
        RECT 48.045 52.260 48.675 52.540 ;
        RECT 48.155 52.220 48.615 52.260 ;
        RECT 50.085 52.220 50.545 52.450 ;
        RECT 55.325 52.280 55.785 52.510 ;
        RECT 59.295 52.240 59.925 52.520 ;
        RECT 59.405 52.200 59.865 52.240 ;
        RECT 61.335 52.200 61.795 52.430 ;
        RECT 66.545 52.270 67.005 52.500 ;
        RECT 70.515 52.230 71.145 52.510 ;
        RECT 70.625 52.190 71.085 52.230 ;
        RECT 72.555 52.190 73.015 52.420 ;
        RECT 77.785 52.260 78.245 52.490 ;
        RECT 81.755 52.220 82.385 52.500 ;
        RECT 81.865 52.180 82.325 52.220 ;
        RECT 83.795 52.180 84.255 52.410 ;
        RECT 89.035 52.270 89.495 52.500 ;
        RECT 93.005 52.230 93.635 52.510 ;
        RECT 93.115 52.190 93.575 52.230 ;
        RECT 95.045 52.190 95.505 52.420 ;
        RECT 100.315 52.260 100.775 52.490 ;
        RECT 104.285 52.220 104.915 52.500 ;
        RECT 104.395 52.180 104.855 52.220 ;
        RECT 106.325 52.180 106.785 52.410 ;
        RECT 111.585 52.260 112.045 52.490 ;
        RECT 115.555 52.220 116.185 52.500 ;
        RECT 115.665 52.180 116.125 52.220 ;
        RECT 117.595 52.180 118.055 52.410 ;
        RECT 122.835 52.260 123.295 52.490 ;
        RECT 126.805 52.220 127.435 52.500 ;
        RECT 126.915 52.180 127.375 52.220 ;
        RECT 128.845 52.180 129.305 52.410 ;
        RECT 21.375 52.010 21.605 52.115 ;
        RECT 21.245 50.290 21.615 52.010 ;
        RECT 22.165 51.890 22.395 52.115 ;
        RECT 25.455 51.980 25.685 52.035 ;
        RECT 21.375 50.115 21.605 50.290 ;
        RECT 22.155 50.210 22.525 51.890 ;
        RECT 22.165 50.115 22.395 50.210 ;
        RECT 21.525 49.670 22.245 49.930 ;
        RECT 19.295 46.650 20.065 47.720 ;
        RECT 21.385 47.490 22.105 47.750 ;
        RECT 21.225 47.200 21.455 47.340 ;
        RECT 21.085 46.430 21.475 47.200 ;
        RECT 22.015 47.190 22.245 47.340 ;
        RECT 22.005 46.450 22.375 47.190 ;
        RECT 25.305 47.010 25.735 51.980 ;
        RECT 26.245 51.970 26.475 52.035 ;
        RECT 27.385 51.970 27.615 52.035 ;
        RECT 26.185 46.970 26.585 51.970 ;
        RECT 27.265 46.970 27.665 51.970 ;
        RECT 28.175 51.940 28.405 52.035 ;
        RECT 32.575 52.020 32.805 52.125 ;
        RECT 28.115 46.970 28.545 51.940 ;
        RECT 32.445 50.300 32.815 52.020 ;
        RECT 33.365 51.900 33.595 52.125 ;
        RECT 36.655 51.990 36.885 52.045 ;
        RECT 32.575 50.125 32.805 50.300 ;
        RECT 33.355 50.220 33.725 51.900 ;
        RECT 33.365 50.125 33.595 50.220 ;
        RECT 32.725 49.680 33.445 49.940 ;
        RECT 25.735 46.600 26.195 46.830 ;
        RECT 27.665 46.710 28.125 46.830 ;
        RECT 27.515 46.600 28.125 46.710 ;
        RECT 30.495 46.660 31.265 47.730 ;
        RECT 32.585 47.500 33.305 47.760 ;
        RECT 32.425 47.210 32.655 47.350 ;
        RECT 21.225 46.340 21.455 46.430 ;
        RECT 22.015 46.340 22.245 46.450 ;
        RECT 27.515 46.430 28.095 46.600 ;
        RECT 32.285 46.440 32.675 47.210 ;
        RECT 33.215 47.200 33.445 47.350 ;
        RECT 33.205 46.460 33.575 47.200 ;
        RECT 36.505 47.020 36.935 51.990 ;
        RECT 37.445 51.980 37.675 52.045 ;
        RECT 38.585 51.980 38.815 52.045 ;
        RECT 37.385 46.980 37.785 51.980 ;
        RECT 38.465 46.980 38.865 51.980 ;
        RECT 39.375 51.950 39.605 52.045 ;
        RECT 43.795 51.990 44.025 52.095 ;
        RECT 39.315 46.980 39.745 51.950 ;
        RECT 43.665 50.270 44.035 51.990 ;
        RECT 44.585 51.870 44.815 52.095 ;
        RECT 47.875 51.960 48.105 52.015 ;
        RECT 43.795 50.095 44.025 50.270 ;
        RECT 44.575 50.190 44.945 51.870 ;
        RECT 44.585 50.095 44.815 50.190 ;
        RECT 43.945 49.650 44.665 49.910 ;
        RECT 36.935 46.610 37.395 46.840 ;
        RECT 38.865 46.720 39.325 46.840 ;
        RECT 38.715 46.610 39.325 46.720 ;
        RECT 41.715 46.630 42.485 47.700 ;
        RECT 43.805 47.470 44.525 47.730 ;
        RECT 43.645 47.180 43.875 47.320 ;
        RECT 32.425 46.350 32.655 46.440 ;
        RECT 33.215 46.350 33.445 46.460 ;
        RECT 38.715 46.440 39.295 46.610 ;
        RECT 43.505 46.410 43.895 47.180 ;
        RECT 44.435 47.170 44.665 47.320 ;
        RECT 44.425 46.430 44.795 47.170 ;
        RECT 47.725 46.990 48.155 51.960 ;
        RECT 48.665 51.950 48.895 52.015 ;
        RECT 49.805 51.950 50.035 52.015 ;
        RECT 48.605 46.950 49.005 51.950 ;
        RECT 49.685 46.950 50.085 51.950 ;
        RECT 50.595 51.920 50.825 52.015 ;
        RECT 55.045 51.970 55.275 52.075 ;
        RECT 50.535 46.950 50.965 51.920 ;
        RECT 54.915 50.250 55.285 51.970 ;
        RECT 55.835 51.850 56.065 52.075 ;
        RECT 59.125 51.940 59.355 51.995 ;
        RECT 55.045 50.075 55.275 50.250 ;
        RECT 55.825 50.170 56.195 51.850 ;
        RECT 55.835 50.075 56.065 50.170 ;
        RECT 55.195 49.630 55.915 49.890 ;
        RECT 48.155 46.580 48.615 46.810 ;
        RECT 50.085 46.690 50.545 46.810 ;
        RECT 49.935 46.580 50.545 46.690 ;
        RECT 52.965 46.610 53.735 47.680 ;
        RECT 55.055 47.450 55.775 47.710 ;
        RECT 54.895 47.160 55.125 47.300 ;
        RECT 43.645 46.320 43.875 46.410 ;
        RECT 44.435 46.320 44.665 46.430 ;
        RECT 49.935 46.410 50.515 46.580 ;
        RECT 54.755 46.390 55.145 47.160 ;
        RECT 55.685 47.150 55.915 47.300 ;
        RECT 55.675 46.410 56.045 47.150 ;
        RECT 58.975 46.970 59.405 51.940 ;
        RECT 59.915 51.930 60.145 51.995 ;
        RECT 61.055 51.930 61.285 51.995 ;
        RECT 59.855 46.930 60.255 51.930 ;
        RECT 60.935 46.930 61.335 51.930 ;
        RECT 61.845 51.900 62.075 51.995 ;
        RECT 66.265 51.960 66.495 52.065 ;
        RECT 61.785 46.930 62.215 51.900 ;
        RECT 66.135 50.240 66.505 51.960 ;
        RECT 67.055 51.840 67.285 52.065 ;
        RECT 70.345 51.930 70.575 51.985 ;
        RECT 66.265 50.065 66.495 50.240 ;
        RECT 67.045 50.160 67.415 51.840 ;
        RECT 67.055 50.065 67.285 50.160 ;
        RECT 66.415 49.620 67.135 49.880 ;
        RECT 59.405 46.560 59.865 46.790 ;
        RECT 61.335 46.670 61.795 46.790 ;
        RECT 61.185 46.560 61.795 46.670 ;
        RECT 64.185 46.600 64.955 47.670 ;
        RECT 66.275 47.440 66.995 47.700 ;
        RECT 66.115 47.150 66.345 47.290 ;
        RECT 54.895 46.300 55.125 46.390 ;
        RECT 55.685 46.300 55.915 46.410 ;
        RECT 61.185 46.390 61.765 46.560 ;
        RECT 65.975 46.380 66.365 47.150 ;
        RECT 66.905 47.140 67.135 47.290 ;
        RECT 66.895 46.400 67.265 47.140 ;
        RECT 70.195 46.960 70.625 51.930 ;
        RECT 71.135 51.920 71.365 51.985 ;
        RECT 72.275 51.920 72.505 51.985 ;
        RECT 71.075 46.920 71.475 51.920 ;
        RECT 72.155 46.920 72.555 51.920 ;
        RECT 73.065 51.890 73.295 51.985 ;
        RECT 77.505 51.950 77.735 52.055 ;
        RECT 73.005 46.920 73.435 51.890 ;
        RECT 77.375 50.230 77.745 51.950 ;
        RECT 78.295 51.830 78.525 52.055 ;
        RECT 81.585 51.920 81.815 51.975 ;
        RECT 77.505 50.055 77.735 50.230 ;
        RECT 78.285 50.150 78.655 51.830 ;
        RECT 78.295 50.055 78.525 50.150 ;
        RECT 77.655 49.610 78.375 49.870 ;
        RECT 70.625 46.550 71.085 46.780 ;
        RECT 72.555 46.660 73.015 46.780 ;
        RECT 72.405 46.550 73.015 46.660 ;
        RECT 75.425 46.590 76.195 47.660 ;
        RECT 77.515 47.430 78.235 47.690 ;
        RECT 77.355 47.140 77.585 47.280 ;
        RECT 66.115 46.290 66.345 46.380 ;
        RECT 66.905 46.290 67.135 46.400 ;
        RECT 72.405 46.380 72.985 46.550 ;
        RECT 77.215 46.370 77.605 47.140 ;
        RECT 78.145 47.130 78.375 47.280 ;
        RECT 78.135 46.390 78.505 47.130 ;
        RECT 81.435 46.950 81.865 51.920 ;
        RECT 82.375 51.910 82.605 51.975 ;
        RECT 83.515 51.910 83.745 51.975 ;
        RECT 82.315 46.910 82.715 51.910 ;
        RECT 83.395 46.910 83.795 51.910 ;
        RECT 84.305 51.880 84.535 51.975 ;
        RECT 88.755 51.960 88.985 52.065 ;
        RECT 84.245 46.910 84.675 51.880 ;
        RECT 88.625 50.240 88.995 51.960 ;
        RECT 89.545 51.840 89.775 52.065 ;
        RECT 92.835 51.930 93.065 51.985 ;
        RECT 88.755 50.065 88.985 50.240 ;
        RECT 89.535 50.160 89.905 51.840 ;
        RECT 89.545 50.065 89.775 50.160 ;
        RECT 88.905 49.620 89.625 49.880 ;
        RECT 81.865 46.540 82.325 46.770 ;
        RECT 83.795 46.650 84.255 46.770 ;
        RECT 83.645 46.540 84.255 46.650 ;
        RECT 86.675 46.600 87.445 47.670 ;
        RECT 88.765 47.440 89.485 47.700 ;
        RECT 88.605 47.150 88.835 47.290 ;
        RECT 77.355 46.280 77.585 46.370 ;
        RECT 78.145 46.280 78.375 46.390 ;
        RECT 83.645 46.370 84.225 46.540 ;
        RECT 88.465 46.380 88.855 47.150 ;
        RECT 89.395 47.140 89.625 47.290 ;
        RECT 89.385 46.400 89.755 47.140 ;
        RECT 92.685 46.960 93.115 51.930 ;
        RECT 93.625 51.920 93.855 51.985 ;
        RECT 94.765 51.920 94.995 51.985 ;
        RECT 93.565 46.920 93.965 51.920 ;
        RECT 94.645 46.920 95.045 51.920 ;
        RECT 95.555 51.890 95.785 51.985 ;
        RECT 100.035 51.950 100.265 52.055 ;
        RECT 95.495 46.920 95.925 51.890 ;
        RECT 99.905 50.230 100.275 51.950 ;
        RECT 100.825 51.830 101.055 52.055 ;
        RECT 104.115 51.920 104.345 51.975 ;
        RECT 100.035 50.055 100.265 50.230 ;
        RECT 100.815 50.150 101.185 51.830 ;
        RECT 100.825 50.055 101.055 50.150 ;
        RECT 100.185 49.610 100.905 49.870 ;
        RECT 93.115 46.550 93.575 46.780 ;
        RECT 95.045 46.660 95.505 46.780 ;
        RECT 94.895 46.550 95.505 46.660 ;
        RECT 97.955 46.590 98.725 47.660 ;
        RECT 100.045 47.430 100.765 47.690 ;
        RECT 99.885 47.140 100.115 47.280 ;
        RECT 88.605 46.290 88.835 46.380 ;
        RECT 89.395 46.290 89.625 46.400 ;
        RECT 94.895 46.380 95.475 46.550 ;
        RECT 99.745 46.370 100.135 47.140 ;
        RECT 100.675 47.130 100.905 47.280 ;
        RECT 100.665 46.390 101.035 47.130 ;
        RECT 103.965 46.950 104.395 51.920 ;
        RECT 104.905 51.910 105.135 51.975 ;
        RECT 106.045 51.910 106.275 51.975 ;
        RECT 104.845 46.910 105.245 51.910 ;
        RECT 105.925 46.910 106.325 51.910 ;
        RECT 106.835 51.880 107.065 51.975 ;
        RECT 111.305 51.950 111.535 52.055 ;
        RECT 106.775 46.910 107.205 51.880 ;
        RECT 111.175 50.230 111.545 51.950 ;
        RECT 112.095 51.830 112.325 52.055 ;
        RECT 115.385 51.920 115.615 51.975 ;
        RECT 111.305 50.055 111.535 50.230 ;
        RECT 112.085 50.150 112.455 51.830 ;
        RECT 112.095 50.055 112.325 50.150 ;
        RECT 111.455 49.610 112.175 49.870 ;
        RECT 104.395 46.540 104.855 46.770 ;
        RECT 106.325 46.650 106.785 46.770 ;
        RECT 106.175 46.540 106.785 46.650 ;
        RECT 109.225 46.590 109.995 47.660 ;
        RECT 111.315 47.430 112.035 47.690 ;
        RECT 111.155 47.140 111.385 47.280 ;
        RECT 99.885 46.280 100.115 46.370 ;
        RECT 100.675 46.280 100.905 46.390 ;
        RECT 106.175 46.370 106.755 46.540 ;
        RECT 111.015 46.370 111.405 47.140 ;
        RECT 111.945 47.130 112.175 47.280 ;
        RECT 111.935 46.390 112.305 47.130 ;
        RECT 115.235 46.950 115.665 51.920 ;
        RECT 116.175 51.910 116.405 51.975 ;
        RECT 117.315 51.910 117.545 51.975 ;
        RECT 116.115 46.910 116.515 51.910 ;
        RECT 117.195 46.910 117.595 51.910 ;
        RECT 118.105 51.880 118.335 51.975 ;
        RECT 122.555 51.950 122.785 52.055 ;
        RECT 118.045 46.910 118.475 51.880 ;
        RECT 122.425 50.230 122.795 51.950 ;
        RECT 123.345 51.830 123.575 52.055 ;
        RECT 126.635 51.920 126.865 51.975 ;
        RECT 122.555 50.055 122.785 50.230 ;
        RECT 123.335 50.150 123.705 51.830 ;
        RECT 123.345 50.055 123.575 50.150 ;
        RECT 122.705 49.610 123.425 49.870 ;
        RECT 115.665 46.540 116.125 46.770 ;
        RECT 117.595 46.650 118.055 46.770 ;
        RECT 117.445 46.540 118.055 46.650 ;
        RECT 120.475 46.590 121.245 47.660 ;
        RECT 122.565 47.430 123.285 47.690 ;
        RECT 122.405 47.140 122.635 47.280 ;
        RECT 111.155 46.280 111.385 46.370 ;
        RECT 111.945 46.280 112.175 46.390 ;
        RECT 117.445 46.370 118.025 46.540 ;
        RECT 122.265 46.370 122.655 47.140 ;
        RECT 123.195 47.130 123.425 47.280 ;
        RECT 123.185 46.390 123.555 47.130 ;
        RECT 126.485 46.950 126.915 51.920 ;
        RECT 127.425 51.910 127.655 51.975 ;
        RECT 128.565 51.910 128.795 51.975 ;
        RECT 127.365 46.910 127.765 51.910 ;
        RECT 128.445 46.910 128.845 51.910 ;
        RECT 129.355 51.880 129.585 51.975 ;
        RECT 129.295 46.910 129.725 51.880 ;
        RECT 126.915 46.540 127.375 46.770 ;
        RECT 128.845 46.650 129.305 46.770 ;
        RECT 128.695 46.540 129.305 46.650 ;
        RECT 122.405 46.280 122.635 46.370 ;
        RECT 123.195 46.280 123.425 46.390 ;
        RECT 128.695 46.370 129.275 46.540 ;
        RECT 21.505 45.950 21.965 46.180 ;
        RECT 32.705 45.960 33.165 46.190 ;
        RECT 43.925 45.930 44.385 46.160 ;
        RECT 55.175 45.910 55.635 46.140 ;
        RECT 66.395 45.900 66.855 46.130 ;
        RECT 77.635 45.890 78.095 46.120 ;
        RECT 88.885 45.900 89.345 46.130 ;
        RECT 100.165 45.890 100.625 46.120 ;
        RECT 111.435 45.890 111.895 46.120 ;
        RECT 122.685 45.890 123.145 46.120 ;
        RECT 29.055 45.020 41.225 45.030 ;
        RECT 17.855 45.005 41.225 45.020 ;
        RECT 15.900 45.000 41.225 45.005 ;
        RECT 15.900 44.980 52.445 45.000 ;
        RECT 15.900 44.970 63.695 44.980 ;
        RECT 15.900 44.960 74.915 44.970 ;
        RECT 85.235 44.960 97.405 44.970 ;
        RECT 15.900 43.880 131.205 44.960 ;
        RECT 15.900 43.870 30.025 43.880 ;
        RECT 15.900 43.855 18.690 43.870 ;
        RECT 15.900 41.620 17.050 43.855 ;
        RECT 40.275 43.850 131.205 43.880 ;
        RECT 51.525 43.830 131.205 43.850 ;
        RECT 62.745 43.820 131.205 43.830 ;
        RECT 73.985 43.810 86.155 43.820 ;
        RECT 96.515 43.810 131.205 43.820 ;
        RECT 29.015 43.330 41.185 43.340 ;
        RECT 17.815 43.310 41.185 43.330 ;
        RECT 142.830 43.320 144.150 43.340 ;
        RECT 17.815 43.290 52.405 43.310 ;
        RECT 140.750 43.300 144.150 43.320 ;
        RECT 17.815 43.280 63.655 43.290 ;
        RECT 119.895 43.280 144.150 43.300 ;
        RECT 17.815 43.270 74.875 43.280 ;
        RECT 85.195 43.270 97.365 43.280 ;
        RECT 108.685 43.270 144.150 43.280 ;
        RECT 17.815 42.180 144.150 43.270 ;
        RECT 18.755 42.150 144.150 42.180 ;
        RECT 18.755 42.120 131.165 42.150 ;
        RECT 18.755 42.090 109.655 42.120 ;
        RECT 18.755 42.080 98.445 42.090 ;
        RECT 41.325 42.070 98.445 42.080 ;
        RECT 142.830 42.070 144.150 42.150 ;
        RECT 41.325 42.060 87.205 42.070 ;
        RECT 75.035 42.050 87.205 42.060 ;
        RECT 15.900 41.540 19.685 41.620 ;
        RECT 142.070 41.610 146.210 41.640 ;
        RECT 119.855 41.590 146.210 41.610 ;
        RECT 108.645 41.550 146.210 41.590 ;
        RECT 15.900 41.520 42.165 41.540 ;
        RECT 97.445 41.530 146.210 41.550 ;
        RECT 15.900 41.510 75.875 41.520 ;
        RECT 86.235 41.510 146.210 41.530 ;
        RECT 15.900 40.500 146.210 41.510 ;
        RECT 15.900 40.480 142.320 40.500 ;
        RECT 15.900 40.470 140.920 40.480 ;
        RECT 18.715 40.460 140.920 40.470 ;
        RECT 142.070 40.460 142.250 40.480 ;
        RECT 18.715 40.440 120.815 40.460 ;
        RECT 18.715 40.400 109.615 40.440 ;
        RECT 18.715 40.390 98.405 40.400 ;
        RECT 41.285 40.380 98.405 40.390 ;
        RECT 41.285 40.370 87.165 40.380 ;
        RECT 74.995 40.360 87.165 40.370 ;
        RECT 26.775 39.230 27.235 39.460 ;
        RECT 38.055 39.230 38.515 39.460 ;
        RECT 49.345 39.210 49.805 39.440 ;
        RECT 60.565 39.210 61.025 39.440 ;
        RECT 71.765 39.210 72.225 39.440 ;
        RECT 83.055 39.200 83.515 39.430 ;
        RECT 94.295 39.220 94.755 39.450 ;
        RECT 105.505 39.240 105.965 39.470 ;
        RECT 116.705 39.280 117.165 39.510 ;
        RECT 127.915 39.300 128.375 39.530 ;
        RECT 20.645 38.810 21.225 38.980 ;
        RECT 26.495 38.960 26.725 39.070 ;
        RECT 27.285 38.980 27.515 39.070 ;
        RECT 20.615 38.700 21.225 38.810 ;
        RECT 20.615 38.580 21.075 38.700 ;
        RECT 22.545 38.580 23.005 38.810 ;
        RECT 20.195 33.470 20.625 38.440 ;
        RECT 20.335 33.375 20.565 33.470 ;
        RECT 21.075 33.440 21.475 38.440 ;
        RECT 22.155 33.440 22.555 38.440 ;
        RECT 21.125 33.375 21.355 33.440 ;
        RECT 22.265 33.375 22.495 33.440 ;
        RECT 23.005 33.430 23.435 38.400 ;
        RECT 26.365 38.220 26.735 38.960 ;
        RECT 26.495 38.070 26.725 38.220 ;
        RECT 27.265 38.210 27.655 38.980 ;
        RECT 31.925 38.810 32.505 38.980 ;
        RECT 37.775 38.960 38.005 39.070 ;
        RECT 38.565 38.980 38.795 39.070 ;
        RECT 27.285 38.070 27.515 38.210 ;
        RECT 26.635 37.660 27.355 37.920 ;
        RECT 28.675 37.690 29.445 38.760 ;
        RECT 31.895 38.700 32.505 38.810 ;
        RECT 31.895 38.580 32.355 38.700 ;
        RECT 33.825 38.580 34.285 38.810 ;
        RECT 26.495 35.480 27.215 35.740 ;
        RECT 26.345 35.200 26.575 35.295 ;
        RECT 26.215 33.520 26.585 35.200 ;
        RECT 27.135 35.120 27.365 35.295 ;
        RECT 23.055 33.375 23.285 33.430 ;
        RECT 26.345 33.295 26.575 33.520 ;
        RECT 27.125 33.400 27.495 35.120 ;
        RECT 31.475 33.470 31.905 38.440 ;
        RECT 27.135 33.295 27.365 33.400 ;
        RECT 31.615 33.375 31.845 33.470 ;
        RECT 32.355 33.440 32.755 38.440 ;
        RECT 33.435 33.440 33.835 38.440 ;
        RECT 32.405 33.375 32.635 33.440 ;
        RECT 33.545 33.375 33.775 33.440 ;
        RECT 34.285 33.430 34.715 38.400 ;
        RECT 37.645 38.220 38.015 38.960 ;
        RECT 37.775 38.070 38.005 38.220 ;
        RECT 38.545 38.210 38.935 38.980 ;
        RECT 43.215 38.790 43.795 38.960 ;
        RECT 49.065 38.940 49.295 39.050 ;
        RECT 49.855 38.960 50.085 39.050 ;
        RECT 38.565 38.070 38.795 38.210 ;
        RECT 37.915 37.660 38.635 37.920 ;
        RECT 39.955 37.690 40.725 38.760 ;
        RECT 43.185 38.680 43.795 38.790 ;
        RECT 43.185 38.560 43.645 38.680 ;
        RECT 45.115 38.560 45.575 38.790 ;
        RECT 37.775 35.480 38.495 35.740 ;
        RECT 37.625 35.200 37.855 35.295 ;
        RECT 37.495 33.520 37.865 35.200 ;
        RECT 38.415 35.120 38.645 35.295 ;
        RECT 34.335 33.375 34.565 33.430 ;
        RECT 37.625 33.295 37.855 33.520 ;
        RECT 38.405 33.400 38.775 35.120 ;
        RECT 42.765 33.450 43.195 38.420 ;
        RECT 38.415 33.295 38.645 33.400 ;
        RECT 42.905 33.355 43.135 33.450 ;
        RECT 43.645 33.420 44.045 38.420 ;
        RECT 44.725 33.420 45.125 38.420 ;
        RECT 43.695 33.355 43.925 33.420 ;
        RECT 44.835 33.355 45.065 33.420 ;
        RECT 45.575 33.410 46.005 38.380 ;
        RECT 48.935 38.200 49.305 38.940 ;
        RECT 49.065 38.050 49.295 38.200 ;
        RECT 49.835 38.190 50.225 38.960 ;
        RECT 54.435 38.790 55.015 38.960 ;
        RECT 60.285 38.940 60.515 39.050 ;
        RECT 61.075 38.960 61.305 39.050 ;
        RECT 49.855 38.050 50.085 38.190 ;
        RECT 49.205 37.640 49.925 37.900 ;
        RECT 51.245 37.670 52.015 38.740 ;
        RECT 54.405 38.680 55.015 38.790 ;
        RECT 54.405 38.560 54.865 38.680 ;
        RECT 56.335 38.560 56.795 38.790 ;
        RECT 49.065 35.460 49.785 35.720 ;
        RECT 48.915 35.180 49.145 35.275 ;
        RECT 48.785 33.500 49.155 35.180 ;
        RECT 49.705 35.100 49.935 35.275 ;
        RECT 45.625 33.355 45.855 33.410 ;
        RECT 48.915 33.275 49.145 33.500 ;
        RECT 49.695 33.380 50.065 35.100 ;
        RECT 53.985 33.450 54.415 38.420 ;
        RECT 49.705 33.275 49.935 33.380 ;
        RECT 54.125 33.355 54.355 33.450 ;
        RECT 54.865 33.420 55.265 38.420 ;
        RECT 55.945 33.420 56.345 38.420 ;
        RECT 54.915 33.355 55.145 33.420 ;
        RECT 56.055 33.355 56.285 33.420 ;
        RECT 56.795 33.410 57.225 38.380 ;
        RECT 60.155 38.200 60.525 38.940 ;
        RECT 60.285 38.050 60.515 38.200 ;
        RECT 61.055 38.190 61.445 38.960 ;
        RECT 65.635 38.790 66.215 38.960 ;
        RECT 71.485 38.940 71.715 39.050 ;
        RECT 72.275 38.960 72.505 39.050 ;
        RECT 61.075 38.050 61.305 38.190 ;
        RECT 60.425 37.640 61.145 37.900 ;
        RECT 62.465 37.670 63.235 38.740 ;
        RECT 65.605 38.680 66.215 38.790 ;
        RECT 65.605 38.560 66.065 38.680 ;
        RECT 67.535 38.560 67.995 38.790 ;
        RECT 60.285 35.460 61.005 35.720 ;
        RECT 60.135 35.180 60.365 35.275 ;
        RECT 60.005 33.500 60.375 35.180 ;
        RECT 60.925 35.100 61.155 35.275 ;
        RECT 56.845 33.355 57.075 33.410 ;
        RECT 60.135 33.275 60.365 33.500 ;
        RECT 60.915 33.380 61.285 35.100 ;
        RECT 65.185 33.450 65.615 38.420 ;
        RECT 60.925 33.275 61.155 33.380 ;
        RECT 65.325 33.355 65.555 33.450 ;
        RECT 66.065 33.420 66.465 38.420 ;
        RECT 67.145 33.420 67.545 38.420 ;
        RECT 66.115 33.355 66.345 33.420 ;
        RECT 67.255 33.355 67.485 33.420 ;
        RECT 67.995 33.410 68.425 38.380 ;
        RECT 71.355 38.200 71.725 38.940 ;
        RECT 71.485 38.050 71.715 38.200 ;
        RECT 72.255 38.190 72.645 38.960 ;
        RECT 76.925 38.780 77.505 38.950 ;
        RECT 82.775 38.930 83.005 39.040 ;
        RECT 83.565 38.950 83.795 39.040 ;
        RECT 72.275 38.050 72.505 38.190 ;
        RECT 71.625 37.640 72.345 37.900 ;
        RECT 73.665 37.670 74.435 38.740 ;
        RECT 76.895 38.670 77.505 38.780 ;
        RECT 76.895 38.550 77.355 38.670 ;
        RECT 78.825 38.550 79.285 38.780 ;
        RECT 71.485 35.460 72.205 35.720 ;
        RECT 71.335 35.180 71.565 35.275 ;
        RECT 71.205 33.500 71.575 35.180 ;
        RECT 72.125 35.100 72.355 35.275 ;
        RECT 68.045 33.355 68.275 33.410 ;
        RECT 71.335 33.275 71.565 33.500 ;
        RECT 72.115 33.380 72.485 35.100 ;
        RECT 76.475 33.440 76.905 38.410 ;
        RECT 72.125 33.275 72.355 33.380 ;
        RECT 76.615 33.345 76.845 33.440 ;
        RECT 77.355 33.410 77.755 38.410 ;
        RECT 78.435 33.410 78.835 38.410 ;
        RECT 77.405 33.345 77.635 33.410 ;
        RECT 78.545 33.345 78.775 33.410 ;
        RECT 79.285 33.400 79.715 38.370 ;
        RECT 82.645 38.190 83.015 38.930 ;
        RECT 82.775 38.040 83.005 38.190 ;
        RECT 83.545 38.180 83.935 38.950 ;
        RECT 88.165 38.800 88.745 38.970 ;
        RECT 94.015 38.950 94.245 39.060 ;
        RECT 94.805 38.970 95.035 39.060 ;
        RECT 83.565 38.040 83.795 38.180 ;
        RECT 82.915 37.630 83.635 37.890 ;
        RECT 84.955 37.660 85.725 38.730 ;
        RECT 88.135 38.690 88.745 38.800 ;
        RECT 88.135 38.570 88.595 38.690 ;
        RECT 90.065 38.570 90.525 38.800 ;
        RECT 82.775 35.450 83.495 35.710 ;
        RECT 82.625 35.170 82.855 35.265 ;
        RECT 82.495 33.490 82.865 35.170 ;
        RECT 83.415 35.090 83.645 35.265 ;
        RECT 79.335 33.345 79.565 33.400 ;
        RECT 82.625 33.265 82.855 33.490 ;
        RECT 83.405 33.370 83.775 35.090 ;
        RECT 87.715 33.460 88.145 38.430 ;
        RECT 83.415 33.265 83.645 33.370 ;
        RECT 87.855 33.365 88.085 33.460 ;
        RECT 88.595 33.430 88.995 38.430 ;
        RECT 89.675 33.430 90.075 38.430 ;
        RECT 88.645 33.365 88.875 33.430 ;
        RECT 89.785 33.365 90.015 33.430 ;
        RECT 90.525 33.420 90.955 38.390 ;
        RECT 93.885 38.210 94.255 38.950 ;
        RECT 94.015 38.060 94.245 38.210 ;
        RECT 94.785 38.200 95.175 38.970 ;
        RECT 99.375 38.820 99.955 38.990 ;
        RECT 105.225 38.970 105.455 39.080 ;
        RECT 106.015 38.990 106.245 39.080 ;
        RECT 94.805 38.060 95.035 38.200 ;
        RECT 94.155 37.650 94.875 37.910 ;
        RECT 96.195 37.680 96.965 38.750 ;
        RECT 99.345 38.710 99.955 38.820 ;
        RECT 99.345 38.590 99.805 38.710 ;
        RECT 101.275 38.590 101.735 38.820 ;
        RECT 94.015 35.470 94.735 35.730 ;
        RECT 93.865 35.190 94.095 35.285 ;
        RECT 93.735 33.510 94.105 35.190 ;
        RECT 94.655 35.110 94.885 35.285 ;
        RECT 90.575 33.365 90.805 33.420 ;
        RECT 93.865 33.285 94.095 33.510 ;
        RECT 94.645 33.390 95.015 35.110 ;
        RECT 98.925 33.480 99.355 38.450 ;
        RECT 94.655 33.285 94.885 33.390 ;
        RECT 99.065 33.385 99.295 33.480 ;
        RECT 99.805 33.450 100.205 38.450 ;
        RECT 100.885 33.450 101.285 38.450 ;
        RECT 99.855 33.385 100.085 33.450 ;
        RECT 100.995 33.385 101.225 33.450 ;
        RECT 101.735 33.440 102.165 38.410 ;
        RECT 105.095 38.230 105.465 38.970 ;
        RECT 105.225 38.080 105.455 38.230 ;
        RECT 105.995 38.220 106.385 38.990 ;
        RECT 110.575 38.860 111.155 39.030 ;
        RECT 116.425 39.010 116.655 39.120 ;
        RECT 117.215 39.030 117.445 39.120 ;
        RECT 106.015 38.080 106.245 38.220 ;
        RECT 105.365 37.670 106.085 37.930 ;
        RECT 107.405 37.700 108.175 38.770 ;
        RECT 110.545 38.750 111.155 38.860 ;
        RECT 110.545 38.630 111.005 38.750 ;
        RECT 112.475 38.630 112.935 38.860 ;
        RECT 105.225 35.490 105.945 35.750 ;
        RECT 105.075 35.210 105.305 35.305 ;
        RECT 104.945 33.530 105.315 35.210 ;
        RECT 105.865 35.130 106.095 35.305 ;
        RECT 101.785 33.385 102.015 33.440 ;
        RECT 105.075 33.305 105.305 33.530 ;
        RECT 105.855 33.410 106.225 35.130 ;
        RECT 110.125 33.520 110.555 38.490 ;
        RECT 110.265 33.425 110.495 33.520 ;
        RECT 111.005 33.490 111.405 38.490 ;
        RECT 112.085 33.490 112.485 38.490 ;
        RECT 111.055 33.425 111.285 33.490 ;
        RECT 112.195 33.425 112.425 33.490 ;
        RECT 112.935 33.480 113.365 38.450 ;
        RECT 116.295 38.270 116.665 39.010 ;
        RECT 116.425 38.120 116.655 38.270 ;
        RECT 117.195 38.260 117.585 39.030 ;
        RECT 121.785 38.880 122.365 39.050 ;
        RECT 127.635 39.030 127.865 39.140 ;
        RECT 128.425 39.050 128.655 39.140 ;
        RECT 117.215 38.120 117.445 38.260 ;
        RECT 116.565 37.710 117.285 37.970 ;
        RECT 118.605 37.740 119.375 38.810 ;
        RECT 121.755 38.770 122.365 38.880 ;
        RECT 121.755 38.650 122.215 38.770 ;
        RECT 123.685 38.650 124.145 38.880 ;
        RECT 116.425 35.530 117.145 35.790 ;
        RECT 116.275 35.250 116.505 35.345 ;
        RECT 116.145 33.570 116.515 35.250 ;
        RECT 117.065 35.170 117.295 35.345 ;
        RECT 112.985 33.425 113.215 33.480 ;
        RECT 105.865 33.305 106.095 33.410 ;
        RECT 116.275 33.345 116.505 33.570 ;
        RECT 117.055 33.450 117.425 35.170 ;
        RECT 121.335 33.540 121.765 38.510 ;
        RECT 117.065 33.345 117.295 33.450 ;
        RECT 121.475 33.445 121.705 33.540 ;
        RECT 122.215 33.510 122.615 38.510 ;
        RECT 123.295 33.510 123.695 38.510 ;
        RECT 122.265 33.445 122.495 33.510 ;
        RECT 123.405 33.445 123.635 33.510 ;
        RECT 124.145 33.500 124.575 38.470 ;
        RECT 127.505 38.290 127.875 39.030 ;
        RECT 127.635 38.140 127.865 38.290 ;
        RECT 128.405 38.280 128.795 39.050 ;
        RECT 128.425 38.140 128.655 38.280 ;
        RECT 127.775 37.730 128.495 37.990 ;
        RECT 129.815 37.760 130.585 38.830 ;
        RECT 142.850 37.630 144.170 38.900 ;
        RECT 127.635 35.550 128.355 35.810 ;
        RECT 127.485 35.270 127.715 35.365 ;
        RECT 127.355 33.590 127.725 35.270 ;
        RECT 128.275 35.190 128.505 35.365 ;
        RECT 124.195 33.445 124.425 33.500 ;
        RECT 127.485 33.365 127.715 33.590 ;
        RECT 128.265 33.470 128.635 35.190 ;
        RECT 128.275 33.365 128.505 33.470 ;
        RECT 20.615 32.940 21.075 33.170 ;
        RECT 22.545 33.130 23.005 33.170 ;
        RECT 22.485 32.850 23.115 33.130 ;
        RECT 26.625 32.860 27.085 33.090 ;
        RECT 31.895 32.940 32.355 33.170 ;
        RECT 33.825 33.130 34.285 33.170 ;
        RECT 33.765 32.850 34.395 33.130 ;
        RECT 37.905 32.860 38.365 33.090 ;
        RECT 43.185 32.920 43.645 33.150 ;
        RECT 45.115 33.110 45.575 33.150 ;
        RECT 45.055 32.830 45.685 33.110 ;
        RECT 49.195 32.840 49.655 33.070 ;
        RECT 54.405 32.920 54.865 33.150 ;
        RECT 56.335 33.110 56.795 33.150 ;
        RECT 56.275 32.830 56.905 33.110 ;
        RECT 60.415 32.840 60.875 33.070 ;
        RECT 65.605 32.920 66.065 33.150 ;
        RECT 67.535 33.110 67.995 33.150 ;
        RECT 67.475 32.830 68.105 33.110 ;
        RECT 71.615 32.840 72.075 33.070 ;
        RECT 76.895 32.910 77.355 33.140 ;
        RECT 78.825 33.100 79.285 33.140 ;
        RECT 78.765 32.820 79.395 33.100 ;
        RECT 82.905 32.830 83.365 33.060 ;
        RECT 88.135 32.930 88.595 33.160 ;
        RECT 90.065 33.120 90.525 33.160 ;
        RECT 90.005 32.840 90.635 33.120 ;
        RECT 94.145 32.850 94.605 33.080 ;
        RECT 99.345 32.950 99.805 33.180 ;
        RECT 101.275 33.140 101.735 33.180 ;
        RECT 101.215 32.860 101.845 33.140 ;
        RECT 105.355 32.870 105.815 33.100 ;
        RECT 110.545 32.990 111.005 33.220 ;
        RECT 112.475 33.180 112.935 33.220 ;
        RECT 112.415 32.900 113.045 33.180 ;
        RECT 116.555 32.910 117.015 33.140 ;
        RECT 121.755 33.010 122.215 33.240 ;
        RECT 123.685 33.200 124.145 33.240 ;
        RECT 123.625 32.920 124.255 33.200 ;
        RECT 127.765 32.930 128.225 33.160 ;
        RECT 23.185 30.880 27.925 31.180 ;
        RECT 34.465 30.880 39.205 31.180 ;
        RECT 45.755 30.860 50.495 31.160 ;
        RECT 56.975 30.860 61.715 31.160 ;
        RECT 68.175 30.860 72.915 31.160 ;
        RECT 79.465 30.850 84.205 31.150 ;
        RECT 90.705 30.870 95.445 31.170 ;
        RECT 101.915 30.890 106.655 31.190 ;
        RECT 113.115 30.930 117.855 31.230 ;
        RECT 124.325 30.950 129.065 31.250 ;
        RECT 19.485 20.270 19.905 30.160 ;
        RECT 19.585 20.090 19.815 20.270 ;
        RECT 20.805 20.260 21.175 30.210 ;
        RECT 20.875 20.090 21.105 20.260 ;
        RECT 21.935 20.220 22.305 30.170 ;
        RECT 27.255 20.270 27.615 30.190 ;
        RECT 30.765 20.270 31.185 30.160 ;
        RECT 22.015 20.090 22.245 20.220 ;
        RECT 27.305 20.090 27.535 20.270 ;
        RECT 30.865 20.090 31.095 20.270 ;
        RECT 32.085 20.260 32.455 30.210 ;
        RECT 32.155 20.090 32.385 20.260 ;
        RECT 33.215 20.220 33.585 30.170 ;
        RECT 38.535 20.270 38.895 30.190 ;
        RECT 33.295 20.090 33.525 20.220 ;
        RECT 38.585 20.090 38.815 20.270 ;
        RECT 42.055 20.250 42.475 30.140 ;
        RECT 42.155 20.070 42.385 20.250 ;
        RECT 43.375 20.240 43.745 30.190 ;
        RECT 43.445 20.070 43.675 20.240 ;
        RECT 44.505 20.200 44.875 30.150 ;
        RECT 49.825 20.250 50.185 30.170 ;
        RECT 53.275 20.250 53.695 30.140 ;
        RECT 44.585 20.070 44.815 20.200 ;
        RECT 49.875 20.070 50.105 20.250 ;
        RECT 53.375 20.070 53.605 20.250 ;
        RECT 54.595 20.240 54.965 30.190 ;
        RECT 54.665 20.070 54.895 20.240 ;
        RECT 55.725 20.200 56.095 30.150 ;
        RECT 61.045 20.250 61.405 30.170 ;
        RECT 64.475 20.250 64.895 30.140 ;
        RECT 55.805 20.070 56.035 20.200 ;
        RECT 61.095 20.070 61.325 20.250 ;
        RECT 64.575 20.070 64.805 20.250 ;
        RECT 65.795 20.240 66.165 30.190 ;
        RECT 65.865 20.070 66.095 20.240 ;
        RECT 66.925 20.200 67.295 30.150 ;
        RECT 72.245 20.250 72.605 30.170 ;
        RECT 67.005 20.070 67.235 20.200 ;
        RECT 72.295 20.070 72.525 20.250 ;
        RECT 75.765 20.240 76.185 30.130 ;
        RECT 75.865 20.060 76.095 20.240 ;
        RECT 77.085 20.230 77.455 30.180 ;
        RECT 77.155 20.060 77.385 20.230 ;
        RECT 78.215 20.190 78.585 30.140 ;
        RECT 83.535 20.240 83.895 30.160 ;
        RECT 87.005 20.260 87.425 30.150 ;
        RECT 78.295 20.060 78.525 20.190 ;
        RECT 83.585 20.060 83.815 20.240 ;
        RECT 87.105 20.080 87.335 20.260 ;
        RECT 88.325 20.250 88.695 30.200 ;
        RECT 88.395 20.080 88.625 20.250 ;
        RECT 89.455 20.210 89.825 30.160 ;
        RECT 94.775 20.260 95.135 30.180 ;
        RECT 98.215 20.280 98.635 30.170 ;
        RECT 89.535 20.080 89.765 20.210 ;
        RECT 94.825 20.080 95.055 20.260 ;
        RECT 98.315 20.100 98.545 20.280 ;
        RECT 99.535 20.270 99.905 30.220 ;
        RECT 99.605 20.100 99.835 20.270 ;
        RECT 100.665 20.230 101.035 30.180 ;
        RECT 105.985 20.280 106.345 30.200 ;
        RECT 109.415 20.320 109.835 30.210 ;
        RECT 100.745 20.100 100.975 20.230 ;
        RECT 106.035 20.100 106.265 20.280 ;
        RECT 109.515 20.140 109.745 20.320 ;
        RECT 110.735 20.310 111.105 30.260 ;
        RECT 110.805 20.140 111.035 20.310 ;
        RECT 111.865 20.270 112.235 30.220 ;
        RECT 117.185 20.320 117.545 30.240 ;
        RECT 120.625 20.340 121.045 30.230 ;
        RECT 111.945 20.140 112.175 20.270 ;
        RECT 117.235 20.140 117.465 20.320 ;
        RECT 120.725 20.160 120.955 20.340 ;
        RECT 121.945 20.330 122.315 30.280 ;
        RECT 122.015 20.160 122.245 20.330 ;
        RECT 123.075 20.290 123.445 30.240 ;
        RECT 128.395 20.340 128.755 30.260 ;
        RECT 123.155 20.160 123.385 20.290 ;
        RECT 128.445 20.160 128.675 20.340 ;
        RECT 132.345 20.170 132.755 30.180 ;
        RECT 137.735 30.120 137.965 30.130 ;
        RECT 132.445 20.130 132.675 20.170 ;
        RECT 137.665 20.080 138.055 30.120 ;
        RECT 19.775 19.610 20.925 19.920 ;
        RECT 22.185 19.620 27.335 19.900 ;
        RECT 31.055 19.610 32.205 19.920 ;
        RECT 33.465 19.620 38.615 19.900 ;
        RECT 42.345 19.590 43.495 19.900 ;
        RECT 44.755 19.600 49.905 19.880 ;
        RECT 53.565 19.590 54.715 19.900 ;
        RECT 55.975 19.600 61.125 19.880 ;
        RECT 64.765 19.590 65.915 19.900 ;
        RECT 67.175 19.600 72.325 19.880 ;
        RECT 76.055 19.580 77.205 19.890 ;
        RECT 78.465 19.590 83.615 19.870 ;
        RECT 87.295 19.600 88.445 19.910 ;
        RECT 89.705 19.610 94.855 19.890 ;
        RECT 98.505 19.620 99.655 19.930 ;
        RECT 100.915 19.630 106.065 19.910 ;
        RECT 109.705 19.660 110.855 19.970 ;
        RECT 112.115 19.670 117.265 19.950 ;
        RECT 120.915 19.680 122.065 19.990 ;
        RECT 123.325 19.690 128.475 19.970 ;
        RECT 132.635 19.640 138.025 19.930 ;
        RECT 142.940 19.110 144.080 37.630 ;
        RECT 13.940 18.460 17.635 18.530 ;
        RECT 117.755 18.510 131.425 18.530 ;
        RECT 106.545 18.470 131.425 18.510 ;
        RECT 13.940 18.440 41.565 18.460 ;
        RECT 95.345 18.450 131.425 18.470 ;
        RECT 13.940 18.430 75.275 18.440 ;
        RECT 84.135 18.430 131.425 18.450 ;
        RECT 13.940 17.380 131.425 18.430 ;
        RECT 142.890 17.990 144.140 19.110 ;
        RECT 145.070 18.880 146.210 40.500 ;
        RECT 145.030 17.960 146.250 18.880 ;
        RECT 13.950 17.370 15.100 17.380 ;
        RECT 16.615 17.360 120.215 17.380 ;
        RECT 16.615 17.320 109.015 17.360 ;
        RECT 16.615 17.310 97.805 17.320 ;
        RECT 39.185 17.300 97.805 17.310 ;
        RECT 39.185 17.290 86.565 17.300 ;
        RECT 72.895 17.280 86.565 17.290 ;
        RECT 117.765 16.950 140.620 16.960 ;
        RECT 142.040 16.950 148.010 16.980 ;
        RECT 117.765 16.940 148.010 16.950 ;
        RECT 106.555 16.900 148.010 16.940 ;
        RECT 16.625 16.870 41.575 16.890 ;
        RECT 95.355 16.880 148.010 16.900 ;
        RECT 16.625 16.860 75.285 16.870 ;
        RECT 84.145 16.860 148.010 16.880 ;
        RECT 16.625 15.840 148.010 16.860 ;
        RECT 16.625 15.820 142.660 15.840 ;
        RECT 16.625 15.810 140.620 15.820 ;
        RECT 142.040 15.810 142.660 15.820 ;
        RECT 16.625 15.790 120.225 15.810 ;
        RECT 16.625 15.750 109.025 15.790 ;
        RECT 16.625 15.740 97.815 15.750 ;
        RECT 39.195 15.730 97.815 15.740 ;
        RECT 39.195 15.720 86.575 15.730 ;
        RECT 72.905 15.710 86.575 15.720 ;
        RECT 131.215 15.460 132.585 15.470 ;
        RECT 12.290 15.390 17.625 15.450 ;
        RECT 117.795 15.440 132.785 15.460 ;
        RECT 106.585 15.400 132.785 15.440 ;
        RECT 12.290 15.370 41.585 15.390 ;
        RECT 95.385 15.380 132.785 15.400 ;
        RECT 12.290 15.360 75.295 15.370 ;
        RECT 84.175 15.360 132.785 15.380 ;
        RECT 12.290 14.320 132.785 15.360 ;
        RECT 142.905 15.040 144.045 15.050 ;
        RECT 12.290 14.310 131.445 14.320 ;
        RECT 12.290 14.300 120.235 14.310 ;
        RECT 12.320 14.280 13.470 14.300 ;
        RECT 16.655 14.290 120.235 14.300 ;
        RECT 16.655 14.250 109.035 14.290 ;
        RECT 16.655 14.240 97.825 14.250 ;
        RECT 39.225 14.230 97.825 14.240 ;
        RECT 39.225 14.220 86.585 14.230 ;
        RECT 72.935 14.210 86.585 14.220 ;
        RECT 142.850 13.920 144.100 15.040 ;
        RECT 145.020 14.870 146.160 14.980 ;
        RECT 144.980 13.950 146.200 14.870 ;
        RECT 16.965 13.800 17.435 13.810 ;
        RECT 10.800 13.780 17.435 13.800 ;
        RECT 10.800 13.720 17.555 13.780 ;
        RECT 117.845 13.770 131.445 13.790 ;
        RECT 106.635 13.730 131.445 13.770 ;
        RECT 10.800 13.700 41.585 13.720 ;
        RECT 95.435 13.710 131.445 13.730 ;
        RECT 10.800 13.690 75.295 13.700 ;
        RECT 84.225 13.690 131.445 13.710 ;
        RECT 10.800 12.650 131.445 13.690 ;
        RECT 16.705 12.640 131.445 12.650 ;
        RECT 16.705 12.620 120.235 12.640 ;
        RECT 16.705 12.580 109.035 12.620 ;
        RECT 16.705 12.570 97.825 12.580 ;
        RECT 39.275 12.560 97.825 12.570 ;
        RECT 39.275 12.550 86.585 12.560 ;
        RECT 72.985 12.540 86.585 12.550 ;
        RECT 128.755 12.240 130.465 12.250 ;
        RECT 117.545 12.220 119.255 12.230 ;
        RECT 106.345 12.180 108.055 12.190 ;
        RECT 27.615 12.170 29.325 12.180 ;
        RECT 38.895 12.170 40.605 12.180 ;
        RECT 25.675 11.030 29.325 12.170 ;
        RECT 36.955 11.030 40.605 12.170 ;
        RECT 95.135 12.160 96.845 12.170 ;
        RECT 50.185 12.150 51.895 12.160 ;
        RECT 61.405 12.150 63.115 12.160 ;
        RECT 72.605 12.150 74.315 12.160 ;
        RECT 25.675 11.020 27.625 11.030 ;
        RECT 36.955 11.020 38.905 11.030 ;
        RECT 48.245 11.010 51.895 12.150 ;
        RECT 59.465 11.010 63.115 12.150 ;
        RECT 70.665 11.010 74.315 12.150 ;
        RECT 83.895 12.140 85.605 12.150 ;
        RECT 48.245 11.000 50.195 11.010 ;
        RECT 59.465 11.000 61.415 11.010 ;
        RECT 70.665 11.000 72.615 11.010 ;
        RECT 81.955 11.000 85.605 12.140 ;
        RECT 93.195 11.020 96.845 12.160 ;
        RECT 104.405 11.040 108.055 12.180 ;
        RECT 115.605 11.080 119.255 12.220 ;
        RECT 126.815 11.100 130.465 12.240 ;
        RECT 126.815 11.090 128.765 11.100 ;
        RECT 115.605 11.070 117.555 11.080 ;
        RECT 104.405 11.030 106.355 11.040 ;
        RECT 93.195 11.010 95.145 11.020 ;
        RECT 81.955 10.990 83.905 11.000 ;
        RECT 142.905 8.580 144.045 13.920 ;
        RECT 74.420 7.440 144.045 8.580 ;
        RECT 74.420 1.410 75.560 7.440 ;
        RECT 145.020 6.630 146.160 13.950 ;
        RECT 93.650 5.490 146.160 6.630 ;
        RECT 93.650 1.480 94.790 5.490 ;
        RECT 146.870 4.560 148.010 15.840 ;
        RECT 113.130 3.420 148.010 4.560 ;
        RECT 113.130 1.610 114.270 3.420 ;
        RECT 149.460 2.770 150.600 64.660 ;
        RECT 131.940 1.880 150.600 2.770 ;
        RECT 131.800 1.630 150.600 1.880 ;
        RECT 74.290 0.160 75.680 1.410 ;
        RECT 93.500 0.230 94.890 1.480 ;
        RECT 112.900 0.360 114.290 1.610 ;
        RECT 131.800 1.380 133.490 1.630 ;
        RECT 151.730 1.420 152.870 66.900 ;
        RECT 131.800 0.430 133.540 1.380 ;
        RECT 113.130 0.330 114.270 0.360 ;
        RECT 151.600 0.300 152.970 1.420 ;
        RECT 93.650 0.150 94.790 0.230 ;
      LAYER met2 ;
        RECT 135.390 223.830 136.740 225.230 ;
        RECT 138.180 223.760 139.530 225.160 ;
        RECT 143.230 223.790 144.580 225.190 ;
        RECT 59.730 204.720 59.990 205.040 ;
        RECT 75.830 204.720 76.090 205.040 ;
        RECT 32.510 203.845 34.390 204.215 ;
        RECT 59.790 203.000 59.930 204.720 ;
        RECT 62.510 203.845 64.390 204.215 ;
        RECT 65.710 203.360 65.970 203.680 ;
        RECT 68.470 203.360 68.730 203.680 ;
        RECT 72.150 203.360 72.410 203.680 ;
        RECT 65.770 203.000 65.910 203.360 ;
        RECT 59.730 202.680 59.990 203.000 ;
        RECT 65.710 202.680 65.970 203.000 ;
        RECT 66.160 202.825 66.440 203.195 ;
        RECT 68.010 203.020 68.270 203.340 ;
        RECT 66.170 202.680 66.430 202.825 ;
        RECT 58.810 202.000 59.070 202.320 ;
        RECT 56.050 201.660 56.310 201.980 ;
        RECT 47.510 201.125 49.390 201.495 ;
        RECT 52.370 199.620 52.630 199.940 ;
        RECT 32.510 198.405 34.390 198.775 ;
        RECT 52.430 197.560 52.570 199.620 ;
        RECT 56.110 197.900 56.250 201.660 ;
        RECT 58.870 197.900 59.010 202.000 ;
        RECT 59.270 199.620 59.530 199.940 ;
        RECT 56.050 197.580 56.310 197.900 ;
        RECT 58.810 197.580 59.070 197.900 ;
        RECT 46.390 197.240 46.650 197.560 ;
        RECT 52.370 197.240 52.630 197.560 ;
        RECT 46.450 195.520 46.590 197.240 ;
        RECT 46.850 196.220 47.110 196.540 ;
        RECT 46.390 195.200 46.650 195.520 ;
        RECT 35.350 195.035 35.610 195.180 ;
        RECT 35.340 194.665 35.620 195.035 ;
        RECT 36.270 194.520 36.530 194.840 ;
        RECT 30.290 194.180 30.550 194.500 ;
        RECT 32.130 194.180 32.390 194.500 ;
        RECT 33.510 194.355 33.770 194.500 ;
        RECT 30.350 192.120 30.490 194.180 ;
        RECT 27.530 191.800 27.790 192.120 ;
        RECT 30.290 191.800 30.550 192.120 ;
        RECT 30.750 191.800 31.010 192.120 ;
        RECT 26.610 188.740 26.870 189.060 ;
        RECT 26.670 187.360 26.810 188.740 ;
        RECT 26.610 187.040 26.870 187.360 ;
        RECT 26.610 183.640 26.870 183.960 ;
        RECT 26.150 182.620 26.410 182.940 ;
        RECT 26.210 181.920 26.350 182.620 ;
        RECT 26.150 181.600 26.410 181.920 ;
        RECT 26.670 178.520 26.810 183.640 ;
        RECT 27.590 183.620 27.730 191.800 ;
        RECT 30.290 190.780 30.550 191.100 ;
        RECT 28.450 188.060 28.710 188.380 ;
        RECT 29.830 188.060 30.090 188.380 ;
        RECT 27.530 183.300 27.790 183.620 ;
        RECT 26.610 178.200 26.870 178.520 ;
        RECT 26.610 177.180 26.870 177.500 ;
        RECT 26.670 175.800 26.810 177.180 ;
        RECT 26.610 175.480 26.870 175.800 ;
        RECT 27.590 175.710 27.730 183.300 ;
        RECT 28.510 181.920 28.650 188.060 ;
        RECT 28.450 181.600 28.710 181.920 ;
        RECT 28.910 181.600 29.170 181.920 ;
        RECT 28.450 180.580 28.710 180.900 ;
        RECT 27.990 177.860 28.250 178.180 ;
        RECT 28.050 176.560 28.190 177.860 ;
        RECT 28.510 177.840 28.650 180.580 ;
        RECT 28.450 177.520 28.710 177.840 ;
        RECT 28.050 176.420 28.650 176.560 ;
        RECT 28.970 176.480 29.110 181.600 ;
        RECT 29.370 179.900 29.630 180.220 ;
        RECT 29.430 178.180 29.570 179.900 ;
        RECT 29.370 177.860 29.630 178.180 ;
        RECT 27.990 175.710 28.250 175.800 ;
        RECT 27.590 175.570 28.250 175.710 ;
        RECT 27.990 175.480 28.250 175.570 ;
        RECT 28.050 173.760 28.190 175.480 ;
        RECT 27.990 173.440 28.250 173.760 ;
        RECT 25.690 172.420 25.950 172.740 ;
        RECT 25.230 171.740 25.490 172.060 ;
        RECT 25.290 165.260 25.430 171.740 ;
        RECT 25.750 168.320 25.890 172.420 ;
        RECT 28.050 172.400 28.190 173.440 ;
        RECT 28.510 173.275 28.650 176.420 ;
        RECT 28.910 176.160 29.170 176.480 ;
        RECT 29.890 175.800 30.030 188.060 ;
        RECT 30.350 187.020 30.490 190.780 ;
        RECT 30.810 190.080 30.950 191.800 ;
        RECT 32.190 191.440 32.330 194.180 ;
        RECT 33.500 193.985 33.780 194.355 ;
        RECT 35.350 194.180 35.610 194.500 ;
        RECT 35.410 193.820 35.550 194.180 ;
        RECT 35.810 193.840 36.070 194.160 ;
        RECT 35.350 193.500 35.610 193.820 ;
        RECT 32.510 192.965 34.390 193.335 ;
        RECT 35.410 192.120 35.550 193.500 ;
        RECT 35.350 191.800 35.610 192.120 ;
        RECT 35.410 191.520 35.550 191.800 ;
        RECT 35.870 191.780 36.010 193.840 ;
        RECT 32.130 191.120 32.390 191.440 ;
        RECT 34.430 191.120 34.690 191.440 ;
        RECT 34.950 191.380 35.550 191.520 ;
        RECT 35.810 191.460 36.070 191.780 ;
        RECT 31.670 190.780 31.930 191.100 ;
        RECT 30.750 189.760 31.010 190.080 ;
        RECT 30.290 186.700 30.550 187.020 ;
        RECT 31.730 186.340 31.870 190.780 ;
        RECT 34.490 190.080 34.630 191.120 ;
        RECT 34.430 189.760 34.690 190.080 ;
        RECT 32.130 189.080 32.390 189.400 ;
        RECT 33.960 189.225 34.240 189.595 ;
        RECT 32.190 188.915 32.330 189.080 ;
        RECT 34.030 189.060 34.170 189.225 ;
        RECT 32.120 188.545 32.400 188.915 ;
        RECT 33.510 188.740 33.770 189.060 ;
        RECT 33.970 188.740 34.230 189.060 ;
        RECT 33.570 188.380 33.710 188.740 ;
        RECT 34.950 188.380 35.090 191.380 ;
        RECT 35.350 190.955 35.610 191.100 ;
        RECT 35.340 190.585 35.620 190.955 ;
        RECT 35.350 189.760 35.610 190.080 ;
        RECT 33.510 188.060 33.770 188.380 ;
        RECT 34.890 188.060 35.150 188.380 ;
        RECT 32.510 187.525 34.390 187.895 ;
        RECT 35.410 186.760 35.550 189.760 ;
        RECT 35.870 187.360 36.010 191.460 ;
        RECT 35.810 187.040 36.070 187.360 ;
        RECT 36.330 187.020 36.470 194.520 ;
        RECT 37.180 193.985 37.460 194.355 ;
        RECT 39.490 194.180 39.750 194.500 ;
        RECT 43.630 194.180 43.890 194.500 ;
        RECT 45.930 194.180 46.190 194.500 ;
        RECT 37.250 192.030 37.390 193.985 ;
        RECT 39.030 192.480 39.290 192.800 ;
        RECT 37.650 192.030 37.910 192.120 ;
        RECT 37.250 191.890 37.910 192.030 ;
        RECT 37.250 189.595 37.390 191.890 ;
        RECT 37.650 191.800 37.910 191.890 ;
        RECT 38.570 191.800 38.830 192.120 ;
        RECT 37.180 189.225 37.460 189.595 ;
        RECT 37.650 189.420 37.910 189.740 ;
        RECT 36.730 188.740 36.990 189.060 ;
        RECT 35.410 186.620 36.010 186.760 ;
        RECT 36.270 186.700 36.530 187.020 ;
        RECT 31.670 186.020 31.930 186.340 ;
        RECT 35.350 186.020 35.610 186.340 ;
        RECT 35.410 183.960 35.550 186.020 ;
        RECT 35.350 183.640 35.610 183.960 ;
        RECT 34.890 182.620 35.150 182.940 ;
        RECT 32.510 182.085 34.390 182.455 ;
        RECT 32.130 180.920 32.390 181.240 ;
        RECT 30.290 180.580 30.550 180.900 ;
        RECT 30.350 178.520 30.490 180.580 ;
        RECT 31.210 178.880 31.470 179.200 ;
        RECT 30.290 178.200 30.550 178.520 ;
        RECT 29.830 175.480 30.090 175.800 ;
        RECT 30.750 174.460 31.010 174.780 ;
        RECT 28.440 172.905 28.720 173.275 ;
        RECT 29.830 172.420 30.090 172.740 ;
        RECT 27.990 172.080 28.250 172.400 ;
        RECT 28.910 172.080 29.170 172.400 ;
        RECT 25.690 168.000 25.950 168.320 ;
        RECT 28.970 167.300 29.110 172.080 ;
        RECT 29.890 170.020 30.030 172.420 ;
        RECT 29.830 169.700 30.090 170.020 ;
        RECT 29.370 167.550 29.630 167.640 ;
        RECT 29.370 167.410 30.030 167.550 ;
        RECT 29.370 167.320 29.630 167.410 ;
        RECT 26.150 166.980 26.410 167.300 ;
        RECT 28.910 166.980 29.170 167.300 ;
        RECT 25.230 164.940 25.490 165.260 ;
        RECT 26.210 164.580 26.350 166.980 ;
        RECT 27.530 166.300 27.790 166.620 ;
        RECT 26.150 164.260 26.410 164.580 ;
        RECT 27.590 161.180 27.730 166.300 ;
        RECT 28.910 161.200 29.170 161.520 ;
        RECT 27.530 160.860 27.790 161.180 ;
        RECT 27.590 159.820 27.730 160.860 ;
        RECT 27.530 159.500 27.790 159.820 ;
        RECT 27.590 154.380 27.730 159.500 ;
        RECT 28.970 157.440 29.110 161.200 ;
        RECT 29.890 158.460 30.030 167.410 ;
        RECT 30.290 161.880 30.550 162.200 ;
        RECT 29.370 158.140 29.630 158.460 ;
        RECT 29.830 158.140 30.090 158.460 ;
        RECT 28.910 157.120 29.170 157.440 ;
        RECT 29.430 156.420 29.570 158.140 ;
        RECT 30.350 157.440 30.490 161.880 ;
        RECT 30.290 157.120 30.550 157.440 ;
        RECT 29.370 156.100 29.630 156.420 ;
        RECT 27.530 154.060 27.790 154.380 ;
        RECT 26.150 153.720 26.410 154.040 ;
        RECT 29.830 153.720 30.090 154.040 ;
        RECT 24.300 148.425 24.580 148.795 ;
        RECT 25.230 148.620 25.490 148.940 ;
        RECT 20.170 123.120 20.430 123.440 ;
        RECT 20.230 104.355 20.370 123.120 ;
        RECT 24.370 121.400 24.510 148.425 ;
        RECT 25.290 146.560 25.430 148.620 ;
        RECT 25.230 146.240 25.490 146.560 ;
        RECT 25.690 145.450 25.950 145.540 ;
        RECT 26.210 145.450 26.350 153.720 ;
        RECT 29.370 153.380 29.630 153.700 ;
        RECT 27.070 152.700 27.330 153.020 ;
        RECT 27.130 150.640 27.270 152.700 ;
        RECT 29.430 151.320 29.570 153.380 ;
        RECT 29.370 151.000 29.630 151.320 ;
        RECT 27.070 150.320 27.330 150.640 ;
        RECT 29.430 149.280 29.570 151.000 ;
        RECT 29.370 148.960 29.630 149.280 ;
        RECT 29.890 147.580 30.030 153.720 ;
        RECT 30.810 152.880 30.950 174.460 ;
        RECT 31.270 156.760 31.410 178.880 ;
        RECT 31.670 177.860 31.930 178.180 ;
        RECT 31.730 175.800 31.870 177.860 ;
        RECT 31.670 175.480 31.930 175.800 ;
        RECT 32.190 175.120 32.330 180.920 ;
        RECT 34.950 180.220 35.090 182.620 ;
        RECT 35.410 180.900 35.550 183.640 ;
        RECT 35.350 180.580 35.610 180.900 ;
        RECT 34.890 179.900 35.150 180.220 ;
        RECT 32.510 176.645 34.390 177.015 ;
        RECT 33.510 175.820 33.770 176.140 ;
        RECT 32.590 175.480 32.850 175.800 ;
        RECT 32.130 174.800 32.390 175.120 ;
        RECT 32.650 172.740 32.790 175.480 ;
        RECT 33.570 173.420 33.710 175.820 ;
        RECT 35.410 175.460 35.550 180.580 ;
        RECT 35.870 176.480 36.010 186.620 ;
        RECT 36.790 183.620 36.930 188.740 ;
        RECT 36.730 183.300 36.990 183.620 ;
        RECT 36.790 181.240 36.930 183.300 ;
        RECT 36.730 180.920 36.990 181.240 ;
        RECT 35.810 176.160 36.070 176.480 ;
        RECT 35.350 175.140 35.610 175.460 ;
        RECT 34.890 174.460 35.150 174.780 ;
        RECT 33.510 173.100 33.770 173.420 ;
        RECT 33.970 173.275 34.230 173.420 ;
        RECT 33.960 172.905 34.240 173.275 ;
        RECT 34.950 173.080 35.090 174.460 ;
        RECT 35.410 173.080 35.550 175.140 ;
        RECT 37.250 174.780 37.390 189.225 ;
        RECT 37.710 183.620 37.850 189.420 ;
        RECT 38.110 189.080 38.370 189.400 ;
        RECT 37.650 183.300 37.910 183.620 ;
        RECT 38.170 178.180 38.310 189.080 ;
        RECT 38.630 188.720 38.770 191.800 ;
        RECT 38.570 188.400 38.830 188.720 ;
        RECT 39.090 188.380 39.230 192.480 ;
        RECT 39.550 191.100 39.690 194.180 ;
        RECT 42.250 193.840 42.510 194.160 ;
        RECT 41.790 192.140 42.050 192.460 ;
        RECT 39.490 190.780 39.750 191.100 ;
        RECT 39.550 190.080 39.690 190.780 ;
        RECT 41.850 190.080 41.990 192.140 ;
        RECT 39.490 189.760 39.750 190.080 ;
        RECT 41.790 189.760 42.050 190.080 ;
        RECT 39.030 188.060 39.290 188.380 ;
        RECT 39.090 185.515 39.230 188.060 ;
        RECT 39.020 185.145 39.300 185.515 ;
        RECT 38.570 183.300 38.830 183.620 ;
        RECT 38.630 181.580 38.770 183.300 ;
        RECT 39.550 183.280 39.690 189.760 ;
        RECT 40.410 188.740 40.670 189.060 ;
        RECT 40.470 184.640 40.610 188.740 ;
        RECT 41.790 188.060 42.050 188.380 ;
        RECT 41.330 187.040 41.590 187.360 ;
        RECT 40.410 184.320 40.670 184.640 ;
        RECT 39.490 182.960 39.750 183.280 ;
        RECT 39.950 182.620 40.210 182.940 ;
        RECT 38.570 181.260 38.830 181.580 ;
        RECT 38.630 179.200 38.770 181.260 ;
        RECT 39.490 179.900 39.750 180.220 ;
        RECT 38.570 178.880 38.830 179.200 ;
        RECT 38.110 177.860 38.370 178.180 ;
        RECT 39.550 177.840 39.690 179.900 ;
        RECT 40.010 179.200 40.150 182.620 ;
        RECT 41.390 181.240 41.530 187.040 ;
        RECT 41.850 187.020 41.990 188.060 ;
        RECT 41.790 186.700 42.050 187.020 ;
        RECT 42.310 184.300 42.450 193.840 ;
        RECT 43.170 191.460 43.430 191.780 ;
        RECT 43.230 189.400 43.370 191.460 ;
        RECT 43.170 189.080 43.430 189.400 ;
        RECT 43.230 186.340 43.370 189.080 ;
        RECT 43.170 186.020 43.430 186.340 ;
        RECT 42.710 185.340 42.970 185.660 ;
        RECT 42.250 183.980 42.510 184.300 ;
        RECT 42.770 181.920 42.910 185.340 ;
        RECT 43.160 185.145 43.440 185.515 ;
        RECT 43.230 183.960 43.370 185.145 ;
        RECT 43.690 184.640 43.830 194.180 ;
        RECT 44.550 190.780 44.810 191.100 ;
        RECT 44.610 189.400 44.750 190.780 ;
        RECT 44.550 189.080 44.810 189.400 ;
        RECT 44.550 188.400 44.810 188.720 ;
        RECT 43.630 184.320 43.890 184.640 ;
        RECT 43.170 183.640 43.430 183.960 ;
        RECT 43.630 183.640 43.890 183.960 ;
        RECT 42.710 181.600 42.970 181.920 ;
        RECT 41.330 180.920 41.590 181.240 ;
        RECT 41.790 180.920 42.050 181.240 ;
        RECT 39.950 178.880 40.210 179.200 ;
        RECT 41.850 178.860 41.990 180.920 ;
        RECT 43.170 178.880 43.430 179.200 ;
        RECT 41.790 178.540 42.050 178.860 ;
        RECT 39.490 177.520 39.750 177.840 ;
        RECT 41.850 177.500 41.990 178.540 ;
        RECT 41.790 177.180 42.050 177.500 ;
        RECT 41.850 176.480 42.910 176.560 ;
        RECT 41.790 176.420 42.970 176.480 ;
        RECT 41.790 176.160 42.050 176.420 ;
        RECT 42.710 176.160 42.970 176.420 ;
        RECT 42.710 175.480 42.970 175.800 ;
        RECT 37.190 174.460 37.450 174.780 ;
        RECT 34.890 172.760 35.150 173.080 ;
        RECT 35.350 172.760 35.610 173.080 ;
        RECT 39.480 172.905 39.760 173.275 ;
        RECT 31.670 172.420 31.930 172.740 ;
        RECT 32.590 172.420 32.850 172.740 ;
        RECT 34.950 172.595 35.090 172.760 ;
        RECT 31.730 168.320 31.870 172.420 ;
        RECT 34.880 172.225 35.160 172.595 ;
        RECT 32.130 171.740 32.390 172.060 ;
        RECT 32.190 170.360 32.330 171.740 ;
        RECT 32.510 171.205 34.390 171.575 ;
        RECT 32.130 170.040 32.390 170.360 ;
        RECT 35.410 170.020 35.550 172.760 ;
        RECT 36.720 172.225 37.000 172.595 ;
        RECT 37.650 172.420 37.910 172.740 ;
        RECT 35.810 170.720 36.070 171.040 ;
        RECT 36.270 170.720 36.530 171.040 ;
        RECT 33.050 169.700 33.310 170.020 ;
        RECT 35.350 169.700 35.610 170.020 ;
        RECT 33.110 169.340 33.250 169.700 ;
        RECT 32.590 169.020 32.850 169.340 ;
        RECT 33.050 169.020 33.310 169.340 ;
        RECT 31.670 168.000 31.930 168.320 ;
        RECT 32.650 167.040 32.790 169.020 ;
        RECT 35.410 167.300 35.550 169.700 ;
        RECT 32.190 166.960 32.790 167.040 ;
        RECT 35.350 166.980 35.610 167.300 ;
        RECT 32.190 166.900 32.850 166.960 ;
        RECT 31.670 164.260 31.930 164.580 ;
        RECT 31.730 162.880 31.870 164.260 ;
        RECT 31.670 162.560 31.930 162.880 ;
        RECT 31.670 159.500 31.930 159.820 ;
        RECT 31.730 157.440 31.870 159.500 ;
        RECT 31.670 157.120 31.930 157.440 ;
        RECT 31.210 156.440 31.470 156.760 ;
        RECT 32.190 156.330 32.330 166.900 ;
        RECT 32.590 166.640 32.850 166.900 ;
        RECT 34.890 166.300 35.150 166.620 ;
        RECT 32.510 165.765 34.390 166.135 ;
        RECT 34.950 161.860 35.090 166.300 ;
        RECT 35.410 164.580 35.550 166.980 ;
        RECT 35.350 164.260 35.610 164.580 ;
        RECT 35.410 162.200 35.550 164.260 ;
        RECT 35.870 162.880 36.010 170.720 ;
        RECT 36.330 170.360 36.470 170.720 ;
        RECT 36.790 170.360 36.930 172.225 ;
        RECT 37.190 172.080 37.450 172.400 ;
        RECT 37.250 170.360 37.390 172.080 ;
        RECT 37.710 170.360 37.850 172.420 ;
        RECT 36.270 170.040 36.530 170.360 ;
        RECT 36.730 170.040 36.990 170.360 ;
        RECT 37.190 170.040 37.450 170.360 ;
        RECT 37.650 170.040 37.910 170.360 ;
        RECT 39.030 169.020 39.290 169.340 ;
        RECT 37.650 168.000 37.910 168.320 ;
        RECT 38.570 168.000 38.830 168.320 ;
        RECT 37.710 166.620 37.850 168.000 ;
        RECT 38.630 167.300 38.770 168.000 ;
        RECT 39.090 167.835 39.230 169.020 ;
        RECT 39.020 167.465 39.300 167.835 ;
        RECT 38.570 166.980 38.830 167.300 ;
        RECT 37.650 166.300 37.910 166.620 ;
        RECT 35.810 162.560 36.070 162.880 ;
        RECT 35.350 161.880 35.610 162.200 ;
        RECT 38.110 161.880 38.370 162.200 ;
        RECT 34.890 161.540 35.150 161.860 ;
        RECT 35.350 161.200 35.610 161.520 ;
        RECT 32.510 160.325 34.390 160.695 ;
        RECT 33.510 157.120 33.770 157.440 ;
        RECT 33.570 156.420 33.710 157.120 ;
        RECT 35.410 157.100 35.550 161.200 ;
        RECT 36.730 160.860 36.990 161.180 ;
        RECT 36.790 159.480 36.930 160.860 ;
        RECT 38.170 159.480 38.310 161.880 ;
        RECT 38.570 161.540 38.830 161.860 ;
        RECT 38.630 160.160 38.770 161.540 ;
        RECT 38.570 159.840 38.830 160.160 ;
        RECT 36.730 159.160 36.990 159.480 ;
        RECT 38.110 159.160 38.370 159.480 ;
        RECT 36.720 158.625 37.000 158.995 ;
        RECT 35.350 156.780 35.610 157.100 ;
        RECT 32.590 156.330 32.850 156.420 ;
        RECT 32.190 156.190 32.850 156.330 ;
        RECT 32.590 156.100 32.850 156.190 ;
        RECT 33.510 156.100 33.770 156.420 ;
        RECT 35.810 155.420 36.070 155.740 ;
        RECT 32.510 154.885 34.390 155.255 ;
        RECT 35.350 154.400 35.610 154.720 ;
        RECT 35.410 154.235 35.550 154.400 ;
        RECT 35.340 153.865 35.620 154.235 ;
        RECT 30.350 152.740 30.950 152.880 ;
        RECT 30.350 152.000 30.490 152.740 ;
        RECT 32.590 152.700 32.850 153.020 ;
        RECT 30.290 151.680 30.550 152.000 ;
        RECT 32.650 151.320 32.790 152.700 ;
        RECT 32.590 151.000 32.850 151.320 ;
        RECT 35.870 150.980 36.010 155.420 ;
        RECT 36.790 153.700 36.930 158.625 ;
        RECT 38.570 156.440 38.830 156.760 ;
        RECT 39.030 156.440 39.290 156.760 ;
        RECT 38.630 154.380 38.770 156.440 ;
        RECT 38.570 154.060 38.830 154.380 ;
        RECT 39.090 153.700 39.230 156.440 ;
        RECT 39.550 156.420 39.690 172.905 ;
        RECT 42.250 171.740 42.510 172.060 ;
        RECT 40.410 170.040 40.670 170.360 ;
        RECT 39.950 169.360 40.210 169.680 ;
        RECT 40.010 167.300 40.150 169.360 ;
        RECT 39.950 166.980 40.210 167.300 ;
        RECT 40.010 161.520 40.150 166.980 ;
        RECT 39.950 161.200 40.210 161.520 ;
        RECT 40.470 159.480 40.610 170.040 ;
        RECT 41.330 169.020 41.590 169.340 ;
        RECT 41.390 167.640 41.530 169.020 ;
        RECT 41.330 167.320 41.590 167.640 ;
        RECT 41.330 166.640 41.590 166.960 ;
        RECT 40.870 162.560 41.130 162.880 ;
        RECT 40.930 160.160 41.070 162.560 ;
        RECT 41.390 161.520 41.530 166.640 ;
        RECT 41.330 161.200 41.590 161.520 ;
        RECT 40.870 159.840 41.130 160.160 ;
        RECT 40.410 159.160 40.670 159.480 ;
        RECT 41.330 158.820 41.590 159.140 ;
        RECT 41.390 156.420 41.530 158.820 ;
        RECT 39.490 156.100 39.750 156.420 ;
        RECT 41.330 156.100 41.590 156.420 ;
        RECT 41.790 156.275 42.050 156.420 ;
        RECT 39.550 154.040 39.690 156.100 ;
        RECT 41.780 155.905 42.060 156.275 ;
        RECT 39.950 155.420 40.210 155.740 ;
        RECT 39.490 153.720 39.750 154.040 ;
        RECT 36.730 153.380 36.990 153.700 ;
        RECT 39.030 153.380 39.290 153.700 ;
        RECT 36.730 152.700 36.990 153.020 ;
        RECT 37.650 152.700 37.910 153.020 ;
        RECT 32.130 150.660 32.390 150.980 ;
        RECT 34.890 150.660 35.150 150.980 ;
        RECT 35.810 150.660 36.070 150.980 ;
        RECT 31.670 149.980 31.930 150.300 ;
        RECT 31.730 148.600 31.870 149.980 ;
        RECT 31.670 148.280 31.930 148.600 ;
        RECT 29.830 147.260 30.090 147.580 ;
        RECT 30.290 147.260 30.550 147.580 ;
        RECT 29.890 145.880 30.030 147.260 ;
        RECT 29.370 145.560 29.630 145.880 ;
        RECT 29.830 145.560 30.090 145.880 ;
        RECT 25.690 145.310 26.350 145.450 ;
        RECT 25.690 145.220 25.950 145.310 ;
        RECT 26.210 143.160 26.350 145.310 ;
        RECT 29.430 143.840 29.570 145.560 ;
        RECT 29.830 144.880 30.090 145.200 ;
        RECT 29.370 143.520 29.630 143.840 ;
        RECT 29.890 143.500 30.030 144.880 ;
        RECT 29.830 143.180 30.090 143.500 ;
        RECT 26.150 142.840 26.410 143.160 ;
        RECT 27.530 143.070 27.790 143.160 ;
        RECT 28.450 143.070 28.710 143.160 ;
        RECT 27.530 142.930 28.710 143.070 ;
        RECT 27.530 142.840 27.790 142.930 ;
        RECT 28.450 142.840 28.710 142.930 ;
        RECT 26.210 140.100 26.350 142.840 ;
        RECT 29.370 142.560 29.630 142.820 ;
        RECT 30.350 142.560 30.490 147.260 ;
        RECT 30.750 146.240 31.010 146.560 ;
        RECT 29.370 142.500 30.490 142.560 ;
        RECT 29.430 142.420 30.490 142.500 ;
        RECT 30.810 142.140 30.950 146.240 ;
        RECT 32.190 142.480 32.330 150.660 ;
        RECT 32.510 149.445 34.390 149.815 ;
        RECT 34.950 148.260 35.090 150.660 ;
        RECT 36.270 149.980 36.530 150.300 ;
        RECT 36.330 148.795 36.470 149.980 ;
        RECT 35.350 148.280 35.610 148.600 ;
        RECT 36.260 148.425 36.540 148.795 ;
        RECT 34.890 147.940 35.150 148.260 ;
        RECT 34.430 147.600 34.690 147.920 ;
        RECT 34.490 146.560 34.630 147.600 ;
        RECT 34.430 146.240 34.690 146.560 ;
        RECT 34.950 144.860 35.090 147.940 ;
        RECT 35.410 146.560 35.550 148.280 ;
        RECT 36.790 148.260 36.930 152.700 ;
        RECT 36.730 148.170 36.990 148.260 ;
        RECT 35.870 148.030 36.990 148.170 ;
        RECT 35.350 146.240 35.610 146.560 ;
        RECT 34.890 144.540 35.150 144.860 ;
        RECT 32.510 144.005 34.390 144.375 ;
        RECT 34.950 143.160 35.090 144.540 ;
        RECT 35.410 143.840 35.550 146.240 ;
        RECT 35.870 146.220 36.010 148.030 ;
        RECT 36.730 147.940 36.990 148.030 ;
        RECT 37.710 147.580 37.850 152.700 ;
        RECT 38.570 151.680 38.830 152.000 ;
        RECT 37.650 147.260 37.910 147.580 ;
        RECT 38.630 146.560 38.770 151.680 ;
        RECT 40.010 150.980 40.150 155.420 ;
        RECT 40.870 154.400 41.130 154.720 ;
        RECT 40.400 151.825 40.680 152.195 ;
        RECT 40.930 152.000 41.070 154.400 ;
        RECT 41.330 153.950 41.590 154.040 ;
        RECT 41.850 153.950 41.990 155.905 ;
        RECT 41.330 153.810 41.990 153.950 ;
        RECT 41.330 153.720 41.590 153.810 ;
        RECT 42.310 153.700 42.450 171.740 ;
        RECT 42.770 167.980 42.910 175.480 ;
        RECT 42.710 167.660 42.970 167.980 ;
        RECT 42.710 166.980 42.970 167.300 ;
        RECT 42.770 159.675 42.910 166.980 ;
        RECT 42.700 159.305 42.980 159.675 ;
        RECT 43.230 158.880 43.370 178.880 ;
        RECT 43.690 178.520 43.830 183.640 ;
        RECT 43.630 178.200 43.890 178.520 ;
        RECT 43.630 177.520 43.890 177.840 ;
        RECT 43.690 172.740 43.830 177.520 ;
        RECT 44.610 175.800 44.750 188.400 ;
        RECT 45.990 188.380 46.130 194.180 ;
        RECT 46.910 192.460 47.050 196.220 ;
        RECT 47.510 195.685 49.390 196.055 ;
        RECT 59.330 195.520 59.470 199.620 ;
        RECT 59.270 195.200 59.530 195.520 ;
        RECT 53.290 194.520 53.550 194.840 ;
        RECT 50.990 194.180 51.250 194.500 ;
        RECT 46.850 192.140 47.110 192.460 ;
        RECT 47.510 190.245 49.390 190.615 ;
        RECT 50.530 189.080 50.790 189.400 ;
        RECT 45.930 188.060 46.190 188.380 ;
        RECT 45.990 186.680 46.130 188.060 ;
        RECT 50.590 187.360 50.730 189.080 ;
        RECT 51.050 188.720 51.190 194.180 ;
        RECT 52.370 193.500 52.630 193.820 ;
        RECT 51.450 191.800 51.710 192.120 ;
        RECT 50.990 188.400 51.250 188.720 ;
        RECT 51.510 187.360 51.650 191.800 ;
        RECT 51.910 191.460 52.170 191.780 ;
        RECT 51.970 190.080 52.110 191.460 ;
        RECT 51.910 189.760 52.170 190.080 ;
        RECT 52.430 187.360 52.570 193.500 ;
        RECT 50.530 187.040 50.790 187.360 ;
        RECT 51.450 187.040 51.710 187.360 ;
        RECT 52.370 187.040 52.630 187.360 ;
        RECT 51.910 186.700 52.170 187.020 ;
        RECT 45.930 186.360 46.190 186.680 ;
        RECT 46.390 186.360 46.650 186.680 ;
        RECT 46.450 184.300 46.590 186.360 ;
        RECT 47.510 184.805 49.390 185.175 ;
        RECT 46.390 183.980 46.650 184.300 ;
        RECT 49.670 181.690 51.650 181.830 ;
        RECT 49.670 181.240 49.810 181.690 ;
        RECT 49.610 180.920 49.870 181.240 ;
        RECT 50.070 180.920 50.330 181.240 ;
        RECT 47.510 179.365 49.390 179.735 ;
        RECT 50.130 179.200 50.270 180.920 ;
        RECT 50.070 178.880 50.330 179.200 ;
        RECT 44.550 175.480 44.810 175.800 ;
        RECT 45.010 175.480 45.270 175.800 ;
        RECT 45.930 175.480 46.190 175.800 ;
        RECT 46.390 175.480 46.650 175.800 ;
        RECT 46.850 175.480 47.110 175.800 ;
        RECT 49.610 175.480 49.870 175.800 ;
        RECT 50.530 175.480 50.790 175.800 ;
        RECT 44.090 174.460 44.350 174.780 ;
        RECT 43.630 172.420 43.890 172.740 ;
        RECT 43.630 171.740 43.890 172.060 ;
        RECT 43.690 169.340 43.830 171.740 ;
        RECT 44.150 170.700 44.290 174.460 ;
        RECT 44.610 173.760 44.750 175.480 ;
        RECT 44.550 173.440 44.810 173.760 ;
        RECT 44.550 172.080 44.810 172.400 ;
        RECT 44.090 170.380 44.350 170.700 ;
        RECT 43.630 169.020 43.890 169.340 ;
        RECT 44.090 169.020 44.350 169.340 ;
        RECT 43.630 166.300 43.890 166.620 ;
        RECT 43.690 164.920 43.830 166.300 ;
        RECT 43.630 164.600 43.890 164.920 ;
        RECT 44.150 164.580 44.290 169.020 ;
        RECT 44.090 164.260 44.350 164.580 ;
        RECT 43.630 160.860 43.890 161.180 ;
        RECT 43.690 159.480 43.830 160.860 ;
        RECT 44.150 159.820 44.290 164.260 ;
        RECT 44.090 159.500 44.350 159.820 ;
        RECT 43.630 159.160 43.890 159.480 ;
        RECT 43.230 158.740 43.830 158.880 ;
        RECT 42.710 155.420 42.970 155.740 ;
        RECT 42.770 154.380 42.910 155.420 ;
        RECT 42.710 154.060 42.970 154.380 ;
        RECT 42.250 153.380 42.510 153.700 ;
        RECT 42.710 152.700 42.970 153.020 ;
        RECT 43.170 152.700 43.430 153.020 ;
        RECT 43.690 152.880 43.830 158.740 ;
        RECT 44.610 158.460 44.750 172.080 ;
        RECT 45.070 171.040 45.210 175.480 ;
        RECT 45.470 174.800 45.730 175.120 ;
        RECT 45.010 170.720 45.270 171.040 ;
        RECT 45.070 160.355 45.210 170.720 ;
        RECT 45.000 159.985 45.280 160.355 ;
        RECT 45.070 159.480 45.210 159.985 ;
        RECT 45.010 159.160 45.270 159.480 ;
        RECT 45.010 158.480 45.270 158.800 ;
        RECT 44.550 158.140 44.810 158.460 ;
        RECT 44.550 156.100 44.810 156.420 ;
        RECT 44.080 153.185 44.360 153.555 ;
        RECT 44.090 153.040 44.350 153.185 ;
        RECT 43.690 152.740 44.290 152.880 ;
        RECT 40.470 151.320 40.610 151.825 ;
        RECT 40.870 151.680 41.130 152.000 ;
        RECT 41.330 151.680 41.590 152.000 ;
        RECT 40.410 151.000 40.670 151.320 ;
        RECT 39.950 150.660 40.210 150.980 ;
        RECT 39.030 149.980 39.290 150.300 ;
        RECT 38.570 146.240 38.830 146.560 ;
        RECT 35.810 145.900 36.070 146.220 ;
        RECT 35.350 143.520 35.610 143.840 ;
        RECT 35.870 143.240 36.010 145.900 ;
        RECT 36.270 144.540 36.530 144.860 ;
        RECT 34.890 142.840 35.150 143.160 ;
        RECT 35.410 143.100 36.010 143.240 ;
        RECT 34.430 142.500 34.690 142.820 ;
        RECT 32.130 142.160 32.390 142.480 ;
        RECT 34.490 142.140 34.630 142.500 ;
        RECT 30.750 141.820 31.010 142.140 ;
        RECT 34.430 141.820 34.690 142.140 ;
        RECT 28.450 140.460 28.710 140.780 ;
        RECT 26.150 139.780 26.410 140.100 ;
        RECT 25.230 137.400 25.490 137.720 ;
        RECT 25.290 131.940 25.430 137.400 ;
        RECT 26.210 134.660 26.350 139.780 ;
        RECT 26.610 139.100 26.870 139.420 ;
        RECT 26.670 137.720 26.810 139.100 ;
        RECT 28.510 138.060 28.650 140.460 ;
        RECT 30.810 139.760 30.950 141.820 ;
        RECT 31.670 140.120 31.930 140.440 ;
        RECT 30.750 139.440 31.010 139.760 ;
        RECT 30.290 139.100 30.550 139.420 ;
        RECT 28.450 137.740 28.710 138.060 ;
        RECT 26.610 137.400 26.870 137.720 ;
        RECT 27.990 135.020 28.250 135.340 ;
        RECT 26.150 134.340 26.410 134.660 ;
        RECT 25.690 133.660 25.950 133.980 ;
        RECT 25.750 132.620 25.890 133.660 ;
        RECT 25.690 132.300 25.950 132.620 ;
        RECT 25.230 131.620 25.490 131.940 ;
        RECT 25.290 129.220 25.430 131.620 ;
        RECT 25.230 128.900 25.490 129.220 ;
        RECT 24.770 128.220 25.030 128.540 ;
        RECT 24.830 127.520 24.970 128.220 ;
        RECT 24.770 127.200 25.030 127.520 ;
        RECT 24.310 121.080 24.570 121.400 ;
        RECT 25.290 118.340 25.430 128.900 ;
        RECT 25.680 126.920 25.960 127.035 ;
        RECT 26.210 126.920 26.350 134.340 ;
        RECT 27.070 133.660 27.330 133.980 ;
        RECT 27.130 129.560 27.270 133.660 ;
        RECT 27.070 129.240 27.330 129.560 ;
        RECT 25.680 126.780 26.350 126.920 ;
        RECT 28.050 126.840 28.190 135.020 ;
        RECT 30.350 134.320 30.490 139.100 ;
        RECT 30.810 138.400 30.950 139.440 ;
        RECT 30.750 138.080 31.010 138.400 ;
        RECT 31.730 135.000 31.870 140.120 ;
        RECT 34.950 139.840 35.090 142.840 ;
        RECT 35.410 142.820 35.550 143.100 ;
        RECT 35.350 142.500 35.610 142.820 ;
        RECT 35.810 142.500 36.070 142.820 ;
        RECT 35.410 141.120 35.550 142.500 ;
        RECT 35.350 140.800 35.610 141.120 ;
        RECT 35.350 139.840 35.610 140.100 ;
        RECT 34.950 139.780 35.610 139.840 ;
        RECT 34.950 139.700 35.550 139.780 ;
        RECT 32.510 138.565 34.390 138.935 ;
        RECT 34.950 137.380 35.090 139.700 ;
        RECT 35.870 138.400 36.010 142.500 ;
        RECT 35.810 138.080 36.070 138.400 ;
        RECT 36.330 137.800 36.470 144.540 ;
        RECT 35.870 137.720 36.470 137.800 ;
        RECT 35.810 137.660 36.470 137.720 ;
        RECT 35.810 137.400 36.070 137.660 ;
        RECT 34.890 137.060 35.150 137.380 ;
        RECT 31.670 134.910 31.930 135.000 ;
        RECT 31.670 134.770 32.330 134.910 ;
        RECT 31.670 134.680 31.930 134.770 ;
        RECT 30.750 134.340 31.010 134.660 ;
        RECT 28.450 134.000 28.710 134.320 ;
        RECT 30.290 134.000 30.550 134.320 ;
        RECT 28.510 127.520 28.650 134.000 ;
        RECT 30.350 131.260 30.490 134.000 ;
        RECT 30.290 130.940 30.550 131.260 ;
        RECT 28.450 127.200 28.710 127.520 ;
        RECT 30.810 126.840 30.950 134.340 ;
        RECT 32.190 132.280 32.330 134.770 ;
        RECT 34.950 134.660 35.090 137.060 ;
        RECT 34.890 134.340 35.150 134.660 ;
        RECT 37.650 134.340 37.910 134.660 ;
        RECT 32.510 133.125 34.390 133.495 ;
        RECT 31.670 131.960 31.930 132.280 ;
        RECT 32.130 131.960 32.390 132.280 ;
        RECT 31.210 128.220 31.470 128.540 ;
        RECT 25.680 126.665 25.960 126.780 ;
        RECT 25.690 126.520 25.950 126.665 ;
        RECT 27.990 126.520 28.250 126.840 ;
        RECT 30.750 126.520 31.010 126.840 ;
        RECT 31.270 126.500 31.410 128.220 ;
        RECT 31.730 127.180 31.870 131.960 ;
        RECT 31.670 126.860 31.930 127.180 ;
        RECT 32.190 126.500 32.330 131.960 ;
        RECT 34.950 131.940 35.090 134.340 ;
        RECT 35.350 134.000 35.610 134.320 ;
        RECT 34.890 131.620 35.150 131.940 ;
        RECT 34.950 129.560 35.090 131.620 ;
        RECT 35.410 129.900 35.550 134.000 ;
        RECT 37.190 132.640 37.450 132.960 ;
        RECT 36.270 131.960 36.530 132.280 ;
        RECT 35.350 129.580 35.610 129.900 ;
        RECT 34.890 129.240 35.150 129.560 ;
        RECT 32.510 127.685 34.390 128.055 ;
        RECT 31.210 126.180 31.470 126.500 ;
        RECT 32.130 126.180 32.390 126.500 ;
        RECT 34.950 124.120 35.090 129.240 ;
        RECT 35.350 128.560 35.610 128.880 ;
        RECT 35.410 126.840 35.550 128.560 ;
        RECT 36.330 127.520 36.470 131.960 ;
        RECT 36.270 127.200 36.530 127.520 ;
        RECT 35.350 126.520 35.610 126.840 ;
        RECT 35.410 125.820 35.550 126.520 ;
        RECT 35.350 125.500 35.610 125.820 ;
        RECT 34.890 123.800 35.150 124.120 ;
        RECT 37.250 123.780 37.390 132.640 ;
        RECT 37.710 130.240 37.850 134.340 ;
        RECT 38.570 132.300 38.830 132.620 ;
        RECT 38.110 130.940 38.370 131.260 ;
        RECT 37.650 129.920 37.910 130.240 ;
        RECT 38.170 129.220 38.310 130.940 ;
        RECT 38.110 128.900 38.370 129.220 ;
        RECT 37.650 126.180 37.910 126.500 ;
        RECT 37.710 124.120 37.850 126.180 ;
        RECT 37.650 123.800 37.910 124.120 ;
        RECT 37.190 123.460 37.450 123.780 ;
        RECT 26.150 123.120 26.410 123.440 ;
        RECT 25.690 122.780 25.950 123.100 ;
        RECT 25.750 122.080 25.890 122.780 ;
        RECT 26.210 122.080 26.350 123.120 ;
        RECT 32.510 122.245 34.390 122.615 ;
        RECT 25.690 121.760 25.950 122.080 ;
        RECT 26.150 121.760 26.410 122.080 ;
        RECT 35.810 121.420 36.070 121.740 ;
        RECT 26.610 121.080 26.870 121.400 ;
        RECT 26.670 118.680 26.810 121.080 ;
        RECT 30.290 120.740 30.550 121.060 ;
        RECT 26.610 118.360 26.870 118.680 ;
        RECT 25.230 118.020 25.490 118.340 ;
        RECT 25.230 115.300 25.490 115.620 ;
        RECT 25.290 104.355 25.430 115.300 ;
        RECT 30.350 104.355 30.490 120.740 ;
        RECT 34.890 117.680 35.150 118.000 ;
        RECT 35.350 117.680 35.610 118.000 ;
        RECT 32.510 116.805 34.390 117.175 ;
        RECT 34.950 116.640 35.090 117.680 ;
        RECT 34.890 116.320 35.150 116.640 ;
        RECT 35.410 104.355 35.550 117.680 ;
        RECT 35.870 114.940 36.010 121.420 ;
        RECT 37.710 121.400 37.850 123.800 ;
        RECT 38.630 123.780 38.770 132.300 ;
        RECT 38.570 123.460 38.830 123.780 ;
        RECT 37.650 121.080 37.910 121.400 ;
        RECT 37.710 118.680 37.850 121.080 ;
        RECT 38.110 120.740 38.370 121.060 ;
        RECT 38.170 119.360 38.310 120.740 ;
        RECT 38.110 119.040 38.370 119.360 ;
        RECT 37.650 118.360 37.910 118.680 ;
        RECT 37.190 118.020 37.450 118.340 ;
        RECT 37.250 115.960 37.390 118.020 ;
        RECT 37.190 115.640 37.450 115.960 ;
        RECT 37.710 115.620 37.850 118.360 ;
        RECT 39.090 118.340 39.230 149.980 ;
        RECT 41.390 149.280 41.530 151.680 ;
        RECT 42.770 149.280 42.910 152.700 ;
        RECT 43.230 150.300 43.370 152.700 ;
        RECT 43.630 151.340 43.890 151.660 ;
        RECT 44.150 151.400 44.290 152.740 ;
        RECT 44.610 152.000 44.750 156.100 ;
        RECT 44.550 151.680 44.810 152.000 ;
        RECT 43.690 150.980 43.830 151.340 ;
        RECT 44.150 151.260 44.750 151.400 ;
        RECT 43.630 150.660 43.890 150.980 ;
        RECT 44.090 150.660 44.350 150.980 ;
        RECT 43.170 149.980 43.430 150.300 ;
        RECT 44.150 149.280 44.290 150.660 ;
        RECT 39.950 148.960 40.210 149.280 ;
        RECT 41.330 148.960 41.590 149.280 ;
        RECT 42.710 148.960 42.970 149.280 ;
        RECT 44.090 148.960 44.350 149.280 ;
        RECT 40.010 148.600 40.150 148.960 ;
        RECT 44.610 148.680 44.750 151.260 ;
        RECT 39.490 148.280 39.750 148.600 ;
        RECT 39.950 148.280 40.210 148.600 ;
        RECT 43.690 148.540 44.750 148.680 ;
        RECT 39.550 145.540 39.690 148.280 ;
        RECT 39.490 145.220 39.750 145.540 ;
        RECT 40.870 144.540 41.130 144.860 ;
        RECT 40.930 143.840 41.070 144.540 ;
        RECT 40.870 143.520 41.130 143.840 ;
        RECT 39.950 131.960 40.210 132.280 ;
        RECT 40.010 129.560 40.150 131.960 ;
        RECT 40.930 131.940 41.070 143.520 ;
        RECT 42.710 142.160 42.970 142.480 ;
        RECT 42.240 140.265 42.520 140.635 ;
        RECT 40.870 131.620 41.130 131.940 ;
        RECT 40.410 131.280 40.670 131.600 ;
        RECT 40.470 131.000 40.610 131.280 ;
        RECT 40.470 130.860 41.990 131.000 ;
        RECT 39.950 129.240 40.210 129.560 ;
        RECT 39.490 128.900 39.750 129.220 ;
        RECT 39.550 124.800 39.690 128.900 ;
        RECT 39.950 126.520 40.210 126.840 ;
        RECT 39.490 124.480 39.750 124.800 ;
        RECT 40.010 124.460 40.150 126.520 ;
        RECT 39.950 124.140 40.210 124.460 ;
        RECT 40.470 124.120 40.610 130.860 ;
        RECT 41.850 130.240 41.990 130.860 ;
        RECT 40.870 129.920 41.130 130.240 ;
        RECT 41.790 129.920 42.050 130.240 ;
        RECT 40.930 129.640 41.070 129.920 ;
        RECT 40.930 129.500 41.530 129.640 ;
        RECT 41.390 126.840 41.530 129.500 ;
        RECT 41.330 126.520 41.590 126.840 ;
        RECT 40.410 123.800 40.670 124.120 ;
        RECT 41.390 123.780 41.530 126.520 ;
        RECT 42.310 124.800 42.450 140.265 ;
        RECT 42.770 135.680 42.910 142.160 ;
        RECT 42.710 135.360 42.970 135.680 ;
        RECT 43.690 135.000 43.830 148.540 ;
        RECT 44.090 145.220 44.350 145.540 ;
        RECT 44.150 135.680 44.290 145.220 ;
        RECT 44.540 138.225 44.820 138.595 ;
        RECT 44.610 138.060 44.750 138.225 ;
        RECT 44.550 137.740 44.810 138.060 ;
        RECT 44.090 135.360 44.350 135.680 ;
        RECT 43.630 134.680 43.890 135.000 ;
        RECT 44.150 132.620 44.290 135.360 ;
        RECT 45.070 134.660 45.210 158.480 ;
        RECT 45.530 143.160 45.670 174.800 ;
        RECT 45.990 165.115 46.130 175.480 ;
        RECT 46.450 167.980 46.590 175.480 ;
        RECT 46.910 175.315 47.050 175.480 ;
        RECT 46.840 174.945 47.120 175.315 ;
        RECT 46.850 174.460 47.110 174.780 ;
        RECT 46.910 173.160 47.050 174.460 ;
        RECT 47.510 173.925 49.390 174.295 ;
        RECT 46.910 173.020 47.510 173.160 ;
        RECT 46.850 172.080 47.110 172.400 ;
        RECT 46.910 171.915 47.050 172.080 ;
        RECT 46.840 171.545 47.120 171.915 ;
        RECT 47.370 170.700 47.510 173.020 ;
        RECT 47.310 170.380 47.570 170.700 ;
        RECT 47.510 168.485 49.390 168.855 ;
        RECT 49.670 168.320 49.810 175.480 ;
        RECT 50.590 173.760 50.730 175.480 ;
        RECT 50.990 174.460 51.250 174.780 ;
        RECT 50.530 173.440 50.790 173.760 ;
        RECT 50.590 172.740 50.730 173.440 ;
        RECT 50.530 172.420 50.790 172.740 ;
        RECT 51.050 170.360 51.190 174.460 ;
        RECT 50.990 170.040 51.250 170.360 ;
        RECT 50.530 169.700 50.790 170.020 ;
        RECT 50.590 168.320 50.730 169.700 ;
        RECT 49.610 168.000 49.870 168.320 ;
        RECT 50.530 168.000 50.790 168.320 ;
        RECT 46.390 167.660 46.650 167.980 ;
        RECT 45.920 164.745 46.200 165.115 ;
        RECT 46.450 164.490 46.590 167.660 ;
        RECT 50.070 167.320 50.330 167.640 ;
        RECT 47.770 166.980 48.030 167.300 ;
        RECT 46.850 166.640 47.110 166.960 ;
        RECT 46.910 164.920 47.050 166.640 ;
        RECT 47.830 165.600 47.970 166.980 ;
        RECT 47.770 165.280 48.030 165.600 ;
        RECT 46.850 164.600 47.110 164.920 ;
        RECT 45.990 164.350 46.590 164.490 ;
        RECT 45.990 157.100 46.130 164.350 ;
        RECT 46.840 164.065 47.120 164.435 ;
        RECT 46.910 162.880 47.050 164.065 ;
        RECT 47.510 163.045 49.390 163.415 ;
        RECT 46.850 162.560 47.110 162.880 ;
        RECT 50.130 162.540 50.270 167.320 ;
        RECT 51.510 165.000 51.650 181.690 ;
        RECT 51.970 181.240 52.110 186.700 ;
        RECT 53.350 186.340 53.490 194.520 ;
        RECT 59.790 194.500 59.930 202.680 ;
        RECT 67.090 202.340 67.350 202.660 ;
        RECT 66.170 202.000 66.430 202.320 ;
        RECT 66.230 200.280 66.370 202.000 ;
        RECT 66.170 199.960 66.430 200.280 ;
        RECT 67.150 199.940 67.290 202.340 ;
        RECT 68.070 201.980 68.210 203.020 ;
        RECT 68.530 201.980 68.670 203.360 ;
        RECT 70.310 203.020 70.570 203.340 ;
        RECT 72.210 203.195 72.350 203.360 ;
        RECT 68.930 202.680 69.190 203.000 ;
        RECT 68.010 201.660 68.270 201.980 ;
        RECT 68.470 201.660 68.730 201.980 ;
        RECT 67.550 200.640 67.810 200.960 ;
        RECT 65.710 199.620 65.970 199.940 ;
        RECT 67.090 199.620 67.350 199.940 ;
        RECT 65.250 198.940 65.510 199.260 ;
        RECT 62.510 198.405 64.390 198.775 ;
        RECT 65.310 197.560 65.450 198.940 ;
        RECT 65.770 198.240 65.910 199.620 ;
        RECT 65.710 197.920 65.970 198.240 ;
        RECT 65.250 197.240 65.510 197.560 ;
        RECT 61.110 196.900 61.370 197.220 ;
        RECT 56.970 194.180 57.230 194.500 ;
        RECT 59.730 194.180 59.990 194.500 ;
        RECT 57.030 192.120 57.170 194.180 ;
        RECT 56.970 191.800 57.230 192.120 ;
        RECT 60.650 191.800 60.910 192.120 ;
        RECT 54.670 190.780 54.930 191.100 ;
        RECT 56.050 190.780 56.310 191.100 ;
        RECT 54.730 187.020 54.870 190.780 ;
        RECT 56.110 188.720 56.250 190.780 ;
        RECT 56.050 188.400 56.310 188.720 ;
        RECT 54.670 186.700 54.930 187.020 ;
        RECT 60.710 186.680 60.850 191.800 ;
        RECT 61.170 189.400 61.310 196.900 ;
        RECT 65.310 195.520 65.450 197.240 ;
        RECT 67.150 197.220 67.290 199.620 ;
        RECT 67.090 196.900 67.350 197.220 ;
        RECT 65.250 195.200 65.510 195.520 ;
        RECT 62.510 192.965 64.390 193.335 ;
        RECT 61.110 189.080 61.370 189.400 ;
        RECT 56.510 186.360 56.770 186.680 ;
        RECT 60.650 186.360 60.910 186.680 ;
        RECT 53.290 186.020 53.550 186.340 ;
        RECT 54.670 186.020 54.930 186.340 ;
        RECT 52.830 183.980 53.090 184.300 ;
        RECT 52.890 182.940 53.030 183.980 ;
        RECT 53.350 183.620 53.490 186.020 ;
        RECT 54.730 183.960 54.870 186.020 ;
        RECT 55.130 185.340 55.390 185.660 ;
        RECT 54.670 183.640 54.930 183.960 ;
        RECT 53.290 183.300 53.550 183.620 ;
        RECT 52.370 182.620 52.630 182.940 ;
        RECT 52.830 182.620 53.090 182.940 ;
        RECT 52.430 181.240 52.570 182.620 ;
        RECT 52.890 181.240 53.030 182.620 ;
        RECT 51.910 180.920 52.170 181.240 ;
        RECT 52.370 180.920 52.630 181.240 ;
        RECT 52.830 180.920 53.090 181.240 ;
        RECT 51.970 180.640 52.110 180.920 ;
        RECT 51.970 180.500 52.570 180.640 ;
        RECT 54.670 180.580 54.930 180.900 ;
        RECT 51.910 179.900 52.170 180.220 ;
        RECT 51.970 178.520 52.110 179.900 ;
        RECT 51.910 178.200 52.170 178.520 ;
        RECT 52.430 176.140 52.570 180.500 ;
        RECT 52.370 175.820 52.630 176.140 ;
        RECT 51.910 172.420 52.170 172.740 ;
        RECT 51.970 167.300 52.110 172.420 ;
        RECT 52.370 170.720 52.630 171.040 ;
        RECT 51.910 166.980 52.170 167.300 ;
        RECT 52.430 165.600 52.570 170.720 ;
        RECT 53.750 169.020 54.010 169.340 ;
        RECT 53.280 167.465 53.560 167.835 ;
        RECT 52.830 166.300 53.090 166.620 ;
        RECT 52.370 165.280 52.630 165.600 ;
        RECT 51.510 164.860 52.570 165.000 ;
        RECT 50.990 164.260 51.250 164.580 ;
        RECT 50.530 163.580 50.790 163.900 ;
        RECT 50.070 162.220 50.330 162.540 ;
        RECT 46.390 161.880 46.650 162.200 ;
        RECT 46.450 160.160 46.590 161.880 ;
        RECT 50.590 161.860 50.730 163.580 ;
        RECT 51.050 162.880 51.190 164.260 ;
        RECT 50.990 162.560 51.250 162.880 ;
        RECT 50.530 161.540 50.790 161.860 ;
        RECT 46.390 159.840 46.650 160.160 ;
        RECT 46.850 159.840 47.110 160.160 ;
        RECT 46.910 159.560 47.050 159.840 ;
        RECT 46.450 159.480 47.050 159.560 ;
        RECT 46.390 159.420 47.050 159.480 ;
        RECT 46.390 159.160 46.650 159.420 ;
        RECT 50.070 159.160 50.330 159.480 ;
        RECT 46.450 158.460 46.590 159.160 ;
        RECT 46.390 158.140 46.650 158.460 ;
        RECT 49.610 158.140 49.870 158.460 ;
        RECT 47.510 157.605 49.390 157.975 ;
        RECT 45.930 156.780 46.190 157.100 ;
        RECT 46.850 156.440 47.110 156.760 ;
        RECT 45.930 156.275 46.190 156.420 ;
        RECT 45.920 155.905 46.200 156.275 ;
        RECT 45.930 155.420 46.190 155.740 ;
        RECT 45.990 154.720 46.130 155.420 ;
        RECT 45.930 154.400 46.190 154.720 ;
        RECT 46.910 154.040 47.050 156.440 ;
        RECT 48.230 154.060 48.490 154.380 ;
        RECT 46.390 153.720 46.650 154.040 ;
        RECT 46.850 153.720 47.110 154.040 ;
        RECT 46.450 149.280 46.590 153.720 ;
        RECT 46.910 150.980 47.050 153.720 ;
        RECT 48.290 153.360 48.430 154.060 ;
        RECT 49.670 153.440 49.810 158.140 ;
        RECT 50.130 154.380 50.270 159.160 ;
        RECT 51.450 158.140 51.710 158.460 ;
        RECT 50.980 157.265 51.260 157.635 ;
        RECT 51.050 156.760 51.190 157.265 ;
        RECT 51.510 156.760 51.650 158.140 ;
        RECT 50.990 156.440 51.250 156.760 ;
        RECT 51.450 156.440 51.710 156.760 ;
        RECT 51.900 155.905 52.180 156.275 ;
        RECT 50.070 154.060 50.330 154.380 ;
        RECT 50.980 153.865 51.260 154.235 ;
        RECT 50.990 153.720 51.250 153.865 ;
        RECT 48.230 153.040 48.490 153.360 ;
        RECT 49.670 153.300 50.270 153.440 ;
        RECT 47.510 152.165 49.390 152.535 ;
        RECT 48.230 151.340 48.490 151.660 ;
        RECT 46.850 150.660 47.110 150.980 ;
        RECT 46.390 148.960 46.650 149.280 ;
        RECT 48.290 148.600 48.430 151.340 ;
        RECT 48.690 150.660 48.950 150.980 ;
        RECT 48.750 150.300 48.890 150.660 ;
        RECT 48.690 149.980 48.950 150.300 ;
        RECT 49.610 149.980 49.870 150.300 ;
        RECT 49.670 149.280 49.810 149.980 ;
        RECT 49.610 148.960 49.870 149.280 ;
        RECT 48.230 148.280 48.490 148.600 ;
        RECT 49.610 148.280 49.870 148.600 ;
        RECT 47.510 146.725 49.390 147.095 ;
        RECT 49.670 143.840 49.810 148.280 ;
        RECT 45.930 143.520 46.190 143.840 ;
        RECT 49.610 143.520 49.870 143.840 ;
        RECT 45.470 142.840 45.730 143.160 ;
        RECT 45.470 141.820 45.730 142.140 ;
        RECT 45.010 134.340 45.270 134.660 ;
        RECT 44.550 132.640 44.810 132.960 ;
        RECT 44.090 132.300 44.350 132.620 ;
        RECT 43.630 131.620 43.890 131.940 ;
        RECT 43.690 127.520 43.830 131.620 ;
        RECT 44.080 131.425 44.360 131.795 ;
        RECT 43.630 127.200 43.890 127.520 ;
        RECT 44.150 127.180 44.290 131.425 ;
        RECT 44.610 130.240 44.750 132.640 ;
        RECT 44.550 129.920 44.810 130.240 ;
        RECT 45.010 128.900 45.270 129.220 ;
        RECT 44.090 127.035 44.350 127.180 ;
        RECT 44.080 126.665 44.360 127.035 ;
        RECT 45.070 126.840 45.210 128.900 ;
        RECT 45.010 126.520 45.270 126.840 ;
        RECT 42.250 124.480 42.510 124.800 ;
        RECT 41.330 123.460 41.590 123.780 ;
        RECT 44.090 123.120 44.350 123.440 ;
        RECT 45.010 123.120 45.270 123.440 ;
        RECT 39.950 121.420 40.210 121.740 ;
        RECT 40.010 119.020 40.150 121.420 ;
        RECT 40.410 121.080 40.670 121.400 ;
        RECT 39.950 118.700 40.210 119.020 ;
        RECT 38.570 118.195 38.830 118.340 ;
        RECT 38.560 117.825 38.840 118.195 ;
        RECT 39.030 118.020 39.290 118.340 ;
        RECT 38.560 117.145 38.840 117.515 ;
        RECT 38.630 115.960 38.770 117.145 ;
        RECT 38.570 115.640 38.830 115.960 ;
        RECT 37.650 115.300 37.910 115.620 ;
        RECT 35.810 114.620 36.070 114.940 ;
        RECT 40.470 104.355 40.610 121.080 ;
        RECT 20.160 102.355 20.440 104.355 ;
        RECT 25.220 102.355 25.500 104.355 ;
        RECT 30.280 102.355 30.560 104.355 ;
        RECT 35.340 102.355 35.620 104.355 ;
        RECT 40.400 102.355 40.680 104.355 ;
        RECT 44.150 103.800 44.290 123.120 ;
        RECT 45.070 116.640 45.210 123.120 ;
        RECT 45.010 116.320 45.270 116.640 ;
        RECT 45.530 115.960 45.670 141.820 ;
        RECT 45.990 126.840 46.130 143.520 ;
        RECT 46.390 143.180 46.650 143.500 ;
        RECT 46.450 138.400 46.590 143.180 ;
        RECT 47.300 142.985 47.580 143.355 ;
        RECT 49.670 143.160 49.810 143.520 ;
        RECT 47.310 142.840 47.570 142.985 ;
        RECT 49.610 142.840 49.870 143.160 ;
        RECT 49.610 141.820 49.870 142.140 ;
        RECT 47.510 141.285 49.390 141.655 ;
        RECT 49.670 139.760 49.810 141.820 ;
        RECT 49.610 139.440 49.870 139.760 ;
        RECT 46.390 138.080 46.650 138.400 ;
        RECT 47.310 137.400 47.570 137.720 ;
        RECT 49.610 137.400 49.870 137.720 ;
        RECT 47.370 136.700 47.510 137.400 ;
        RECT 47.310 136.380 47.570 136.700 ;
        RECT 47.510 135.845 49.390 136.215 ;
        RECT 46.850 135.360 47.110 135.680 ;
        RECT 46.390 133.660 46.650 133.980 ;
        RECT 45.930 126.520 46.190 126.840 ;
        RECT 46.450 121.740 46.590 133.660 ;
        RECT 46.910 129.900 47.050 135.360 ;
        RECT 49.670 135.340 49.810 137.400 ;
        RECT 49.610 135.020 49.870 135.340 ;
        RECT 49.610 132.640 49.870 132.960 ;
        RECT 47.310 131.795 47.570 131.940 ;
        RECT 47.300 131.425 47.580 131.795 ;
        RECT 47.510 130.405 49.390 130.775 ;
        RECT 46.850 129.580 47.110 129.900 ;
        RECT 46.850 126.520 47.110 126.840 ;
        RECT 46.910 123.100 47.050 126.520 ;
        RECT 47.510 124.965 49.390 125.335 ;
        RECT 48.230 123.800 48.490 124.120 ;
        RECT 46.850 122.780 47.110 123.100 ;
        RECT 46.390 121.420 46.650 121.740 ;
        RECT 48.290 121.400 48.430 123.800 ;
        RECT 49.670 121.400 49.810 132.640 ;
        RECT 50.130 132.280 50.270 153.300 ;
        RECT 50.530 153.040 50.790 153.360 ;
        RECT 50.590 151.320 50.730 153.040 ;
        RECT 51.050 152.000 51.190 153.720 ;
        RECT 50.990 151.680 51.250 152.000 ;
        RECT 50.530 151.000 50.790 151.320 ;
        RECT 50.590 143.160 50.730 151.000 ;
        RECT 51.970 150.980 52.110 155.905 ;
        RECT 52.430 152.880 52.570 164.860 ;
        RECT 52.890 161.180 53.030 166.300 ;
        RECT 53.350 165.000 53.490 167.465 ;
        RECT 53.810 165.600 53.950 169.020 ;
        RECT 53.750 165.280 54.010 165.600 ;
        RECT 53.350 164.860 53.950 165.000 ;
        RECT 53.290 164.260 53.550 164.580 ;
        RECT 53.350 162.540 53.490 164.260 ;
        RECT 53.290 162.220 53.550 162.540 ;
        RECT 52.830 160.860 53.090 161.180 ;
        RECT 52.890 160.160 53.030 160.860 ;
        RECT 52.830 159.840 53.090 160.160 ;
        RECT 52.820 155.905 53.100 156.275 ;
        RECT 52.890 154.040 53.030 155.905 ;
        RECT 52.830 153.720 53.090 154.040 ;
        RECT 53.290 153.720 53.550 154.040 ;
        RECT 52.430 152.740 53.030 152.880 ;
        RECT 51.910 150.660 52.170 150.980 ;
        RECT 52.370 150.320 52.630 150.640 ;
        RECT 51.910 149.980 52.170 150.300 ;
        RECT 51.970 145.540 52.110 149.980 ;
        RECT 51.910 145.220 52.170 145.540 ;
        RECT 52.430 145.280 52.570 150.320 ;
        RECT 52.890 145.880 53.030 152.740 ;
        RECT 53.350 152.000 53.490 153.720 ;
        RECT 53.290 151.680 53.550 152.000 ;
        RECT 52.830 145.560 53.090 145.880 ;
        RECT 53.810 145.540 53.950 164.860 ;
        RECT 54.210 156.440 54.470 156.760 ;
        RECT 54.270 151.660 54.410 156.440 ;
        RECT 54.210 151.340 54.470 151.660 ;
        RECT 52.430 145.140 53.030 145.280 ;
        RECT 53.750 145.220 54.010 145.540 ;
        RECT 52.370 144.540 52.630 144.860 ;
        RECT 50.530 142.840 50.790 143.160 ;
        RECT 51.910 141.820 52.170 142.140 ;
        RECT 50.530 137.060 50.790 137.380 ;
        RECT 50.590 135.340 50.730 137.060 ;
        RECT 50.990 136.720 51.250 137.040 ;
        RECT 50.530 135.020 50.790 135.340 ;
        RECT 51.050 134.660 51.190 136.720 ;
        RECT 50.990 134.340 51.250 134.660 ;
        RECT 50.990 133.660 51.250 133.980 ;
        RECT 51.450 133.660 51.710 133.980 ;
        RECT 51.050 132.960 51.190 133.660 ;
        RECT 50.990 132.640 51.250 132.960 ;
        RECT 50.070 131.960 50.330 132.280 ;
        RECT 50.070 130.940 50.330 131.260 ;
        RECT 50.130 126.500 50.270 130.940 ;
        RECT 51.050 130.240 51.190 132.640 ;
        RECT 51.510 132.620 51.650 133.660 ;
        RECT 51.450 132.300 51.710 132.620 ;
        RECT 51.970 132.280 52.110 141.820 ;
        RECT 51.910 131.960 52.170 132.280 ;
        RECT 50.990 129.920 51.250 130.240 ;
        RECT 52.430 129.220 52.570 144.540 ;
        RECT 52.890 142.820 53.030 145.140 ;
        RECT 53.750 143.520 54.010 143.840 ;
        RECT 52.830 142.500 53.090 142.820 ;
        RECT 52.890 141.120 53.030 142.500 ;
        RECT 52.830 140.800 53.090 141.120 ;
        RECT 53.810 136.700 53.950 143.520 ;
        RECT 54.730 141.120 54.870 180.580 ;
        RECT 55.190 152.880 55.330 185.340 ;
        RECT 56.050 184.320 56.310 184.640 ;
        RECT 56.110 183.960 56.250 184.320 ;
        RECT 56.050 183.640 56.310 183.960 ;
        RECT 56.110 180.900 56.250 183.640 ;
        RECT 56.570 181.920 56.710 186.360 ;
        RECT 60.190 185.680 60.450 186.000 ;
        RECT 58.810 185.340 59.070 185.660 ;
        RECT 59.730 185.340 59.990 185.660 ;
        RECT 58.870 181.920 59.010 185.340 ;
        RECT 59.790 183.960 59.930 185.340 ;
        RECT 59.730 183.640 59.990 183.960 ;
        RECT 60.250 183.280 60.390 185.680 ;
        RECT 60.190 182.960 60.450 183.280 ;
        RECT 59.730 182.620 59.990 182.940 ;
        RECT 56.510 181.600 56.770 181.920 ;
        RECT 58.810 181.600 59.070 181.920 ;
        RECT 57.430 181.260 57.690 181.580 ;
        RECT 56.970 180.920 57.230 181.240 ;
        RECT 56.050 180.580 56.310 180.900 ;
        RECT 57.030 178.860 57.170 180.920 ;
        RECT 56.970 178.540 57.230 178.860 ;
        RECT 56.970 177.860 57.230 178.180 ;
        RECT 57.030 175.800 57.170 177.860 ;
        RECT 57.490 175.800 57.630 181.260 ;
        RECT 58.350 180.580 58.610 180.900 ;
        RECT 57.890 179.900 58.150 180.220 ;
        RECT 57.950 178.520 58.090 179.900 ;
        RECT 58.410 178.520 58.550 180.580 ;
        RECT 57.890 178.200 58.150 178.520 ;
        RECT 58.350 178.200 58.610 178.520 ;
        RECT 59.790 175.800 59.930 182.620 ;
        RECT 60.190 179.900 60.450 180.220 ;
        RECT 60.250 175.800 60.390 179.900 ;
        RECT 60.710 178.180 60.850 186.360 ;
        RECT 61.170 183.960 61.310 189.080 ;
        RECT 62.510 187.525 64.390 187.895 ;
        RECT 64.320 186.505 64.600 186.875 ;
        RECT 64.790 186.590 65.050 186.680 ;
        RECT 65.310 186.590 65.450 195.200 ;
        RECT 66.170 193.840 66.430 194.160 ;
        RECT 65.710 191.800 65.970 192.120 ;
        RECT 63.870 185.515 64.130 185.660 ;
        RECT 63.860 185.145 64.140 185.515 ;
        RECT 61.110 183.640 61.370 183.960 ;
        RECT 61.170 180.810 61.310 183.640 ;
        RECT 64.390 183.620 64.530 186.505 ;
        RECT 64.790 186.450 65.450 186.590 ;
        RECT 64.790 186.360 65.050 186.450 ;
        RECT 64.850 183.620 64.990 186.360 ;
        RECT 65.250 185.340 65.510 185.660 ;
        RECT 65.310 184.640 65.450 185.340 ;
        RECT 65.250 184.320 65.510 184.640 ;
        RECT 64.330 183.300 64.590 183.620 ;
        RECT 64.790 183.300 65.050 183.620 ;
        RECT 62.510 182.085 64.390 182.455 ;
        RECT 62.950 181.260 63.210 181.580 ;
        RECT 61.570 180.810 61.830 180.900 ;
        RECT 61.170 180.670 61.830 180.810 ;
        RECT 60.650 177.860 60.910 178.180 ;
        RECT 56.970 175.480 57.230 175.800 ;
        RECT 57.430 175.480 57.690 175.800 ;
        RECT 59.730 175.480 59.990 175.800 ;
        RECT 60.190 175.480 60.450 175.800 ;
        RECT 56.510 173.100 56.770 173.420 ;
        RECT 55.580 159.985 55.860 160.355 ;
        RECT 56.570 160.240 56.710 173.100 ;
        RECT 57.030 172.400 57.170 175.480 ;
        RECT 58.350 174.460 58.610 174.780 ;
        RECT 56.970 172.080 57.230 172.400 ;
        RECT 57.030 170.700 57.170 172.080 ;
        RECT 56.970 170.380 57.230 170.700 ;
        RECT 56.970 164.260 57.230 164.580 ;
        RECT 57.030 161.860 57.170 164.260 ;
        RECT 56.970 161.540 57.230 161.860 ;
        RECT 57.430 161.200 57.690 161.520 ;
        RECT 56.110 160.100 56.710 160.240 ;
        RECT 55.650 159.480 55.790 159.985 ;
        RECT 55.590 159.160 55.850 159.480 ;
        RECT 55.590 156.100 55.850 156.420 ;
        RECT 56.110 156.275 56.250 160.100 ;
        RECT 56.500 159.305 56.780 159.675 ;
        RECT 57.490 159.480 57.630 161.200 ;
        RECT 56.510 159.160 56.770 159.305 ;
        RECT 57.430 159.160 57.690 159.480 ;
        RECT 57.490 158.800 57.630 159.160 ;
        RECT 57.430 158.480 57.690 158.800 ;
        RECT 57.490 157.440 57.630 158.480 ;
        RECT 57.430 157.120 57.690 157.440 ;
        RECT 56.510 156.780 56.770 157.100 ;
        RECT 55.650 153.700 55.790 156.100 ;
        RECT 56.040 155.905 56.320 156.275 ;
        RECT 56.050 154.290 56.310 154.380 ;
        RECT 56.570 154.290 56.710 156.780 ;
        RECT 57.430 156.100 57.690 156.420 ;
        RECT 56.970 155.420 57.230 155.740 ;
        RECT 57.030 154.380 57.170 155.420 ;
        RECT 56.050 154.150 56.710 154.290 ;
        RECT 56.050 154.060 56.310 154.150 ;
        RECT 56.970 154.060 57.230 154.380 ;
        RECT 55.590 153.380 55.850 153.700 ;
        RECT 57.490 153.360 57.630 156.100 ;
        RECT 57.430 153.040 57.690 153.360 ;
        RECT 55.190 152.740 55.790 152.880 ;
        RECT 55.130 144.540 55.390 144.860 ;
        RECT 54.670 140.800 54.930 141.120 ;
        RECT 54.670 140.120 54.930 140.440 ;
        RECT 53.750 136.380 54.010 136.700 ;
        RECT 53.810 132.280 53.950 136.380 ;
        RECT 54.210 132.870 54.470 132.960 ;
        RECT 54.730 132.870 54.870 140.120 ;
        RECT 54.210 132.730 54.870 132.870 ;
        RECT 54.210 132.640 54.470 132.730 ;
        RECT 53.750 131.960 54.010 132.280 ;
        RECT 52.370 128.900 52.630 129.220 ;
        RECT 53.810 127.520 53.950 131.960 ;
        RECT 53.750 127.200 54.010 127.520 ;
        RECT 50.070 126.180 50.330 126.500 ;
        RECT 51.450 123.120 51.710 123.440 ;
        RECT 51.510 122.080 51.650 123.120 ;
        RECT 55.190 122.080 55.330 144.540 ;
        RECT 55.650 131.600 55.790 152.740 ;
        RECT 56.050 152.700 56.310 153.020 ;
        RECT 57.490 152.880 57.630 153.040 ;
        RECT 57.490 152.740 58.090 152.880 ;
        RECT 56.110 148.600 56.250 152.700 ;
        RECT 57.430 149.980 57.690 150.300 ;
        RECT 56.050 148.280 56.310 148.600 ;
        RECT 56.970 148.280 57.230 148.600 ;
        RECT 56.050 145.900 56.310 146.220 ;
        RECT 56.110 143.160 56.250 145.900 ;
        RECT 56.050 142.840 56.310 143.160 ;
        RECT 57.030 140.440 57.170 148.280 ;
        RECT 57.490 148.170 57.630 149.980 ;
        RECT 57.950 148.940 58.090 152.740 ;
        RECT 57.890 148.620 58.150 148.940 ;
        RECT 57.490 148.030 58.090 148.170 ;
        RECT 57.950 145.200 58.090 148.030 ;
        RECT 58.410 145.880 58.550 174.460 ;
        RECT 60.710 173.080 60.850 177.860 ;
        RECT 61.170 177.840 61.310 180.670 ;
        RECT 61.570 180.580 61.830 180.670 ;
        RECT 63.010 179.200 63.150 181.260 ;
        RECT 64.790 179.900 65.050 180.220 ;
        RECT 64.850 179.200 64.990 179.900 ;
        RECT 62.950 178.880 63.210 179.200 ;
        RECT 64.790 178.880 65.050 179.200 ;
        RECT 61.570 178.540 61.830 178.860 ;
        RECT 62.030 178.540 62.290 178.860 ;
        RECT 61.110 177.520 61.370 177.840 ;
        RECT 61.630 175.800 61.770 178.540 ;
        RECT 62.090 176.140 62.230 178.540 ;
        RECT 65.310 178.520 65.450 184.320 ;
        RECT 65.250 178.200 65.510 178.520 ;
        RECT 64.790 177.860 65.050 178.180 ;
        RECT 62.510 176.645 64.390 177.015 ;
        RECT 64.850 176.480 64.990 177.860 ;
        RECT 64.790 176.160 65.050 176.480 ;
        RECT 62.030 175.820 62.290 176.140 ;
        RECT 61.570 175.480 61.830 175.800 ;
        RECT 64.790 173.100 65.050 173.420 ;
        RECT 60.650 172.760 60.910 173.080 ;
        RECT 60.190 172.420 60.450 172.740 ;
        RECT 59.270 171.740 59.530 172.060 ;
        RECT 59.330 166.870 59.470 171.740 ;
        RECT 60.250 170.360 60.390 172.420 ;
        RECT 60.650 171.740 60.910 172.060 ;
        RECT 60.190 170.040 60.450 170.360 ;
        RECT 59.730 169.760 59.990 170.020 ;
        RECT 59.730 169.700 60.390 169.760 ;
        RECT 59.790 169.620 60.390 169.700 ;
        RECT 59.730 169.020 59.990 169.340 ;
        RECT 59.790 167.640 59.930 169.020 ;
        RECT 59.730 167.320 59.990 167.640 ;
        RECT 59.730 166.870 59.990 166.960 ;
        RECT 59.330 166.730 59.990 166.870 ;
        RECT 59.730 166.640 59.990 166.730 ;
        RECT 58.810 158.140 59.070 158.460 ;
        RECT 58.350 145.560 58.610 145.880 ;
        RECT 58.870 145.540 59.010 158.140 ;
        RECT 59.270 153.380 59.530 153.700 ;
        RECT 59.330 148.600 59.470 153.380 ;
        RECT 59.790 148.600 59.930 166.640 ;
        RECT 60.250 156.420 60.390 169.620 ;
        RECT 60.710 165.260 60.850 171.740 ;
        RECT 62.510 171.205 64.390 171.575 ;
        RECT 64.850 170.020 64.990 173.100 ;
        RECT 65.310 172.740 65.450 178.200 ;
        RECT 65.770 173.420 65.910 191.800 ;
        RECT 66.230 191.100 66.370 193.840 ;
        RECT 66.170 190.780 66.430 191.100 ;
        RECT 66.230 188.120 66.370 190.780 ;
        RECT 66.230 187.980 66.830 188.120 ;
        RECT 66.170 187.040 66.430 187.360 ;
        RECT 66.230 184.640 66.370 187.040 ;
        RECT 66.690 186.000 66.830 187.980 ;
        RECT 66.630 185.680 66.890 186.000 ;
        RECT 66.170 184.320 66.430 184.640 ;
        RECT 67.090 178.880 67.350 179.200 ;
        RECT 67.150 175.460 67.290 178.880 ;
        RECT 67.090 175.140 67.350 175.460 ;
        RECT 67.610 175.120 67.750 200.640 ;
        RECT 68.070 197.900 68.210 201.660 ;
        RECT 68.470 199.620 68.730 199.940 ;
        RECT 68.010 197.580 68.270 197.900 ;
        RECT 68.530 197.220 68.670 199.620 ;
        RECT 68.010 196.900 68.270 197.220 ;
        RECT 68.470 196.900 68.730 197.220 ;
        RECT 68.070 194.160 68.210 196.900 ;
        RECT 68.530 194.840 68.670 196.900 ;
        RECT 68.990 195.520 69.130 202.680 ;
        RECT 69.850 201.660 70.110 201.980 ;
        RECT 69.390 199.620 69.650 199.940 ;
        RECT 68.930 195.200 69.190 195.520 ;
        RECT 68.470 194.520 68.730 194.840 ;
        RECT 68.010 193.840 68.270 194.160 ;
        RECT 68.470 193.840 68.730 194.160 ;
        RECT 68.070 189.400 68.210 193.840 ;
        RECT 68.530 189.480 68.670 193.840 ;
        RECT 69.450 193.820 69.590 199.620 ;
        RECT 69.910 198.240 70.050 201.660 ;
        RECT 69.850 197.920 70.110 198.240 ;
        RECT 69.910 195.180 70.050 197.920 ;
        RECT 69.850 194.860 70.110 195.180 ;
        RECT 69.390 193.500 69.650 193.820 ;
        RECT 69.450 192.460 69.590 193.500 ;
        RECT 69.390 192.140 69.650 192.460 ;
        RECT 69.910 189.740 70.050 194.860 ;
        RECT 70.370 194.500 70.510 203.020 ;
        RECT 72.140 202.825 72.420 203.195 ;
        RECT 75.890 203.000 76.030 204.720 ;
        RECT 92.510 203.845 94.390 204.215 ;
        RECT 80.890 203.360 81.150 203.680 ;
        RECT 75.830 202.680 76.090 203.000 ;
        RECT 75.370 202.340 75.630 202.660 ;
        RECT 74.910 201.660 75.170 201.980 ;
        RECT 70.770 198.940 71.030 199.260 ;
        RECT 70.830 197.560 70.970 198.940 ;
        RECT 70.770 197.240 71.030 197.560 ;
        RECT 70.830 195.520 70.970 197.240 ;
        RECT 73.070 196.220 73.330 196.540 ;
        RECT 70.770 195.200 71.030 195.520 ;
        RECT 70.310 194.180 70.570 194.500 ;
        RECT 70.370 192.800 70.510 194.180 ;
        RECT 70.310 192.710 70.570 192.800 ;
        RECT 70.310 192.570 70.970 192.710 ;
        RECT 70.310 192.480 70.570 192.570 ;
        RECT 70.830 191.780 70.970 192.570 ;
        RECT 73.130 192.460 73.270 196.220 ;
        RECT 74.970 194.160 75.110 201.660 ;
        RECT 75.430 198.240 75.570 202.340 ;
        RECT 75.890 200.960 76.030 202.680 ;
        RECT 79.970 202.000 80.230 202.320 ;
        RECT 76.750 201.660 77.010 201.980 ;
        RECT 79.510 201.660 79.770 201.980 ;
        RECT 75.830 200.640 76.090 200.960 ;
        RECT 75.370 197.920 75.630 198.240 ;
        RECT 75.890 197.640 76.030 200.640 ;
        RECT 76.810 199.600 76.950 201.660 ;
        RECT 77.510 201.125 79.390 201.495 ;
        RECT 79.570 200.620 79.710 201.660 ;
        RECT 79.510 200.300 79.770 200.620 ;
        RECT 80.030 199.940 80.170 202.000 ;
        RECT 80.950 200.620 81.090 203.360 ;
        RECT 96.990 202.680 97.250 203.000 ;
        RECT 101.590 202.680 101.850 203.000 ;
        RECT 95.610 201.660 95.870 201.980 ;
        RECT 80.890 200.300 81.150 200.620 ;
        RECT 80.430 199.960 80.690 200.280 ;
        RECT 79.970 199.620 80.230 199.940 ;
        RECT 76.750 199.280 77.010 199.600 ;
        RECT 79.970 198.940 80.230 199.260 ;
        RECT 75.890 197.500 76.490 197.640 ;
        RECT 74.910 193.840 75.170 194.160 ;
        RECT 76.350 193.820 76.490 197.500 ;
        RECT 76.750 196.220 77.010 196.540 ;
        RECT 76.290 193.500 76.550 193.820 ;
        RECT 76.350 192.460 76.490 193.500 ;
        RECT 76.810 192.800 76.950 196.220 ;
        RECT 77.510 195.685 79.390 196.055 ;
        RECT 80.030 195.180 80.170 198.940 ;
        RECT 80.490 198.240 80.630 199.960 ;
        RECT 80.430 197.920 80.690 198.240 ;
        RECT 80.490 195.520 80.630 197.920 ;
        RECT 80.430 195.200 80.690 195.520 ;
        RECT 79.970 194.860 80.230 195.180 ;
        RECT 80.950 194.500 81.090 200.300 ;
        RECT 91.010 199.620 91.270 199.940 ;
        RECT 87.330 199.280 87.590 199.600 ;
        RECT 86.410 198.940 86.670 199.260 ;
        RECT 86.470 197.900 86.610 198.940 ;
        RECT 81.810 197.580 82.070 197.900 ;
        RECT 86.410 197.580 86.670 197.900 ;
        RECT 81.870 195.520 82.010 197.580 ;
        RECT 87.390 197.220 87.530 199.280 ;
        RECT 89.630 198.940 89.890 199.260 ;
        RECT 87.330 196.900 87.590 197.220 ;
        RECT 89.170 196.900 89.430 197.220 ;
        RECT 81.810 195.200 82.070 195.520 ;
        RECT 87.390 194.500 87.530 196.900 ;
        RECT 89.230 194.840 89.370 196.900 ;
        RECT 89.170 194.520 89.430 194.840 ;
        RECT 79.970 194.180 80.230 194.500 ;
        RECT 80.890 194.180 81.150 194.500 ;
        RECT 87.330 194.180 87.590 194.500 ;
        RECT 79.510 193.500 79.770 193.820 ;
        RECT 76.750 192.480 77.010 192.800 ;
        RECT 79.570 192.460 79.710 193.500 ;
        RECT 80.030 192.800 80.170 194.180 ;
        RECT 80.950 193.820 81.090 194.180 ;
        RECT 80.890 193.500 81.150 193.820 ;
        RECT 86.010 193.420 87.070 193.560 ;
        RECT 79.970 192.480 80.230 192.800 ;
        RECT 86.010 192.460 86.150 193.420 ;
        RECT 86.930 192.800 87.070 193.420 ;
        RECT 86.410 192.480 86.670 192.800 ;
        RECT 86.870 192.480 87.130 192.800 ;
        RECT 73.070 192.140 73.330 192.460 ;
        RECT 76.290 192.140 76.550 192.460 ;
        RECT 79.510 192.140 79.770 192.460 ;
        RECT 80.430 192.140 80.690 192.460 ;
        RECT 85.950 192.140 86.210 192.460 ;
        RECT 73.990 191.800 74.250 192.120 ;
        RECT 70.770 191.460 71.030 191.780 ;
        RECT 68.010 189.080 68.270 189.400 ;
        RECT 68.530 189.340 69.590 189.480 ;
        RECT 69.850 189.420 70.110 189.740 ;
        RECT 68.070 188.380 68.210 189.080 ;
        RECT 68.470 188.400 68.730 188.720 ;
        RECT 68.010 188.060 68.270 188.380 ;
        RECT 68.070 187.020 68.210 188.060 ;
        RECT 68.010 186.700 68.270 187.020 ;
        RECT 68.010 183.300 68.270 183.620 ;
        RECT 68.070 178.180 68.210 183.300 ;
        RECT 68.010 177.860 68.270 178.180 ;
        RECT 68.530 175.460 68.670 188.400 ;
        RECT 68.930 183.640 69.190 183.960 ;
        RECT 68.990 181.240 69.130 183.640 ;
        RECT 68.930 180.920 69.190 181.240 ;
        RECT 68.930 177.180 69.190 177.500 ;
        RECT 68.470 175.140 68.730 175.460 ;
        RECT 67.550 174.800 67.810 175.120 ;
        RECT 65.710 173.100 65.970 173.420 ;
        RECT 66.630 172.760 66.890 173.080 ;
        RECT 68.000 172.905 68.280 173.275 ;
        RECT 65.250 172.420 65.510 172.740 ;
        RECT 64.790 169.700 65.050 170.020 ;
        RECT 61.110 169.360 61.370 169.680 ;
        RECT 63.410 169.360 63.670 169.680 ;
        RECT 61.170 167.640 61.310 169.360 ;
        RECT 62.030 169.020 62.290 169.340 ;
        RECT 61.110 167.320 61.370 167.640 ;
        RECT 60.650 164.940 60.910 165.260 ;
        RECT 61.170 164.580 61.310 167.320 ;
        RECT 62.090 165.600 62.230 169.020 ;
        RECT 63.470 168.320 63.610 169.360 ;
        RECT 63.410 168.000 63.670 168.320 ;
        RECT 62.510 165.765 64.390 166.135 ;
        RECT 62.030 165.280 62.290 165.600 ;
        RECT 60.650 164.260 60.910 164.580 ;
        RECT 61.110 164.260 61.370 164.580 ;
        RECT 60.710 162.200 60.850 164.260 ;
        RECT 61.110 163.580 61.370 163.900 ;
        RECT 64.330 163.580 64.590 163.900 ;
        RECT 61.170 162.200 61.310 163.580 ;
        RECT 64.390 162.540 64.530 163.580 ;
        RECT 64.330 162.220 64.590 162.540 ;
        RECT 64.790 162.220 65.050 162.540 ;
        RECT 65.310 162.280 65.450 172.420 ;
        RECT 65.710 172.080 65.970 172.400 ;
        RECT 65.770 170.360 65.910 172.080 ;
        RECT 65.710 170.040 65.970 170.360 ;
        RECT 65.770 167.300 65.910 170.040 ;
        RECT 66.690 170.020 66.830 172.760 ;
        RECT 66.630 169.700 66.890 170.020 ;
        RECT 65.710 166.980 65.970 167.300 ;
        RECT 60.650 161.880 60.910 162.200 ;
        RECT 61.110 161.880 61.370 162.200 ;
        RECT 64.390 161.860 64.530 162.220 ;
        RECT 64.330 161.540 64.590 161.860 ;
        RECT 64.850 161.520 64.990 162.220 ;
        RECT 65.310 162.140 65.910 162.280 ;
        RECT 65.250 161.540 65.510 161.860 ;
        RECT 64.790 161.200 65.050 161.520 ;
        RECT 62.030 160.860 62.290 161.180 ;
        RECT 61.560 158.625 61.840 158.995 ;
        RECT 61.570 158.480 61.830 158.625 ;
        RECT 60.190 156.100 60.450 156.420 ;
        RECT 61.570 151.680 61.830 152.000 ;
        RECT 61.630 150.980 61.770 151.680 ;
        RECT 61.570 150.660 61.830 150.980 ;
        RECT 60.650 150.320 60.910 150.640 ;
        RECT 61.110 150.320 61.370 150.640 ;
        RECT 59.270 148.280 59.530 148.600 ;
        RECT 59.730 148.280 59.990 148.600 ;
        RECT 58.810 145.220 59.070 145.540 ;
        RECT 57.430 144.880 57.690 145.200 ;
        RECT 57.890 144.880 58.150 145.200 ;
        RECT 57.490 143.840 57.630 144.880 ;
        RECT 57.430 143.520 57.690 143.840 ;
        RECT 57.950 143.160 58.090 144.880 ;
        RECT 58.350 143.520 58.610 143.840 ;
        RECT 57.890 142.840 58.150 143.160 ;
        RECT 56.970 140.120 57.230 140.440 ;
        RECT 57.030 138.400 57.170 140.120 ;
        RECT 56.970 138.080 57.230 138.400 ;
        RECT 57.030 134.660 57.170 138.080 ;
        RECT 57.950 137.380 58.090 142.840 ;
        RECT 58.410 140.100 58.550 143.520 ;
        RECT 58.810 142.840 59.070 143.160 ;
        RECT 58.870 142.480 59.010 142.840 ;
        RECT 58.810 142.160 59.070 142.480 ;
        RECT 58.810 140.800 59.070 141.120 ;
        RECT 59.270 140.800 59.530 141.120 ;
        RECT 58.870 140.635 59.010 140.800 ;
        RECT 58.800 140.265 59.080 140.635 ;
        RECT 58.350 139.780 58.610 140.100 ;
        RECT 58.810 139.440 59.070 139.760 ;
        RECT 58.870 138.400 59.010 139.440 ;
        RECT 58.810 138.080 59.070 138.400 ;
        RECT 58.810 137.400 59.070 137.720 ;
        RECT 57.890 137.060 58.150 137.380 ;
        RECT 57.950 134.660 58.090 137.060 ;
        RECT 58.870 135.340 59.010 137.400 ;
        RECT 58.810 135.020 59.070 135.340 ;
        RECT 56.970 134.570 57.230 134.660 ;
        RECT 56.970 134.430 57.630 134.570 ;
        RECT 56.970 134.340 57.230 134.430 ;
        RECT 56.970 132.640 57.230 132.960 ;
        RECT 55.590 131.280 55.850 131.600 ;
        RECT 56.510 126.180 56.770 126.500 ;
        RECT 56.570 124.800 56.710 126.180 ;
        RECT 56.510 124.480 56.770 124.800 ;
        RECT 57.030 123.780 57.170 132.640 ;
        RECT 57.490 129.560 57.630 134.430 ;
        RECT 57.890 134.340 58.150 134.660 ;
        RECT 59.330 132.360 59.470 140.800 ;
        RECT 59.790 140.100 59.930 148.280 ;
        RECT 60.190 146.240 60.450 146.560 ;
        RECT 59.730 139.780 59.990 140.100 ;
        RECT 59.790 135.340 59.930 139.780 ;
        RECT 59.730 135.020 59.990 135.340 ;
        RECT 59.730 133.660 59.990 133.980 ;
        RECT 58.870 132.220 59.470 132.360 ;
        RECT 59.790 132.280 59.930 133.660 ;
        RECT 57.430 129.240 57.690 129.560 ;
        RECT 57.490 126.500 57.630 129.240 ;
        RECT 57.430 126.180 57.690 126.500 ;
        RECT 57.490 124.120 57.630 126.180 ;
        RECT 57.430 123.800 57.690 124.120 ;
        RECT 58.870 123.780 59.010 132.220 ;
        RECT 59.730 131.960 59.990 132.280 ;
        RECT 59.730 129.240 59.990 129.560 ;
        RECT 59.270 128.220 59.530 128.540 ;
        RECT 59.330 127.520 59.470 128.220 ;
        RECT 59.790 127.520 59.930 129.240 ;
        RECT 59.270 127.200 59.530 127.520 ;
        RECT 59.730 127.200 59.990 127.520 ;
        RECT 60.250 123.780 60.390 146.240 ;
        RECT 60.710 142.820 60.850 150.320 ;
        RECT 61.170 149.280 61.310 150.320 ;
        RECT 61.110 148.960 61.370 149.280 ;
        RECT 61.110 143.180 61.370 143.500 ;
        RECT 60.650 142.500 60.910 142.820 ;
        RECT 60.710 137.720 60.850 142.500 ;
        RECT 61.170 142.140 61.310 143.180 ;
        RECT 61.630 143.160 61.770 150.660 ;
        RECT 62.090 143.840 62.230 160.860 ;
        RECT 62.510 160.325 64.390 160.695 ;
        RECT 64.850 159.140 64.990 161.200 ;
        RECT 65.310 159.820 65.450 161.540 ;
        RECT 65.250 159.500 65.510 159.820 ;
        RECT 65.770 159.480 65.910 162.140 ;
        RECT 65.710 159.160 65.970 159.480 ;
        RECT 64.790 158.820 65.050 159.140 ;
        RECT 62.490 158.480 62.750 158.800 ;
        RECT 62.550 157.635 62.690 158.480 ;
        RECT 62.480 157.265 62.760 157.635 ;
        RECT 65.770 156.420 65.910 159.160 ;
        RECT 65.710 156.100 65.970 156.420 ;
        RECT 64.790 155.420 65.050 155.740 ;
        RECT 65.710 155.420 65.970 155.740 ;
        RECT 62.510 154.885 64.390 155.255 ;
        RECT 64.850 153.700 64.990 155.420 ;
        RECT 64.790 153.380 65.050 153.700 ;
        RECT 65.770 152.000 65.910 155.420 ;
        RECT 66.170 153.720 66.430 154.040 ;
        RECT 65.710 151.680 65.970 152.000 ;
        RECT 64.330 151.340 64.590 151.660 ;
        RECT 64.390 150.720 64.530 151.340 ;
        RECT 64.390 150.580 64.990 150.720 ;
        RECT 62.510 149.445 64.390 149.815 ;
        RECT 64.850 148.680 64.990 150.580 ;
        RECT 63.930 148.540 64.990 148.680 ;
        RECT 63.930 148.260 64.070 148.540 ;
        RECT 63.870 147.940 64.130 148.260 ;
        RECT 63.930 145.540 64.070 147.940 ;
        RECT 66.230 147.920 66.370 153.720 ;
        RECT 64.330 147.600 64.590 147.920 ;
        RECT 66.170 147.600 66.430 147.920 ;
        RECT 64.390 146.220 64.530 147.600 ;
        RECT 66.690 146.640 66.830 169.700 ;
        RECT 68.070 168.320 68.210 172.905 ;
        RECT 68.010 168.000 68.270 168.320 ;
        RECT 67.550 165.280 67.810 165.600 ;
        RECT 67.090 164.940 67.350 165.260 ;
        RECT 67.150 162.880 67.290 164.940 ;
        RECT 67.090 162.560 67.350 162.880 ;
        RECT 67.610 154.235 67.750 165.280 ;
        RECT 68.070 163.900 68.210 168.000 ;
        RECT 68.530 167.300 68.670 175.140 ;
        RECT 68.470 166.980 68.730 167.300 ;
        RECT 68.010 163.580 68.270 163.900 ;
        RECT 68.010 159.500 68.270 159.820 ;
        RECT 68.070 156.275 68.210 159.500 ;
        RECT 68.530 156.760 68.670 166.980 ;
        RECT 68.470 156.440 68.730 156.760 ;
        RECT 68.000 155.905 68.280 156.275 ;
        RECT 68.010 155.420 68.270 155.740 ;
        RECT 67.540 153.865 67.820 154.235 ;
        RECT 67.610 153.360 67.750 153.865 ;
        RECT 67.550 153.040 67.810 153.360 ;
        RECT 68.070 150.300 68.210 155.420 ;
        RECT 68.470 153.720 68.730 154.040 ;
        RECT 68.010 149.980 68.270 150.300 ;
        RECT 68.070 148.260 68.210 149.980 ;
        RECT 67.550 147.940 67.810 148.260 ;
        RECT 68.010 147.940 68.270 148.260 ;
        RECT 67.090 147.260 67.350 147.580 ;
        RECT 65.770 146.500 66.830 146.640 ;
        RECT 64.330 145.900 64.590 146.220 ;
        RECT 63.870 145.220 64.130 145.540 ;
        RECT 64.790 144.880 65.050 145.200 ;
        RECT 62.510 144.005 64.390 144.375 ;
        RECT 62.030 143.520 62.290 143.840 ;
        RECT 63.410 143.180 63.670 143.500 ;
        RECT 61.570 142.840 61.830 143.160 ;
        RECT 61.110 141.820 61.370 142.140 ;
        RECT 61.630 137.720 61.770 142.840 ;
        RECT 63.470 141.120 63.610 143.180 ;
        RECT 64.850 141.120 64.990 144.880 ;
        RECT 65.250 144.540 65.510 144.860 ;
        RECT 65.310 142.140 65.450 144.540 ;
        RECT 65.250 141.820 65.510 142.140 ;
        RECT 63.410 140.800 63.670 141.120 ;
        RECT 64.790 140.800 65.050 141.120 ;
        RECT 62.510 138.565 64.390 138.935 ;
        RECT 64.850 138.060 64.990 140.800 ;
        RECT 65.310 138.400 65.450 141.820 ;
        RECT 65.250 138.080 65.510 138.400 ;
        RECT 64.790 137.740 65.050 138.060 ;
        RECT 60.650 137.400 60.910 137.720 ;
        RECT 61.570 137.400 61.830 137.720 ;
        RECT 65.250 137.400 65.510 137.720 ;
        RECT 60.710 135.680 60.850 137.400 ;
        RECT 64.790 137.060 65.050 137.380 ;
        RECT 64.850 135.680 64.990 137.060 ;
        RECT 60.650 135.360 60.910 135.680 ;
        RECT 64.790 135.360 65.050 135.680 ;
        RECT 60.650 134.680 60.910 135.000 ;
        RECT 60.710 126.840 60.850 134.680 ;
        RECT 62.510 133.125 64.390 133.495 ;
        RECT 64.850 132.960 64.990 135.360 ;
        RECT 64.790 132.640 65.050 132.960 ;
        RECT 63.410 131.620 63.670 131.940 ;
        RECT 61.570 130.940 61.830 131.260 ;
        RECT 61.630 126.840 61.770 130.940 ;
        RECT 63.470 130.240 63.610 131.620 ;
        RECT 65.310 131.600 65.450 137.400 ;
        RECT 65.250 131.280 65.510 131.600 ;
        RECT 65.770 130.240 65.910 146.500 ;
        RECT 66.170 145.900 66.430 146.220 ;
        RECT 66.230 137.720 66.370 145.900 ;
        RECT 66.620 145.705 66.900 146.075 ;
        RECT 66.690 145.540 66.830 145.705 ;
        RECT 66.630 145.220 66.890 145.540 ;
        RECT 66.690 140.100 66.830 145.220 ;
        RECT 66.630 139.780 66.890 140.100 ;
        RECT 67.150 138.400 67.290 147.260 ;
        RECT 67.610 144.860 67.750 147.940 ;
        RECT 67.550 144.540 67.810 144.860 ;
        RECT 68.010 144.540 68.270 144.860 ;
        RECT 67.610 140.780 67.750 144.540 ;
        RECT 68.070 143.160 68.210 144.540 ;
        RECT 68.010 142.840 68.270 143.160 ;
        RECT 67.550 140.460 67.810 140.780 ;
        RECT 68.530 140.440 68.670 153.720 ;
        RECT 68.990 148.600 69.130 177.180 ;
        RECT 69.450 156.420 69.590 189.340 ;
        RECT 69.910 187.360 70.050 189.420 ;
        RECT 70.830 189.400 70.970 191.460 ;
        RECT 72.150 190.780 72.410 191.100 ;
        RECT 70.770 189.080 71.030 189.400 ;
        RECT 70.310 188.060 70.570 188.380 ;
        RECT 69.850 187.040 70.110 187.360 ;
        RECT 69.910 186.680 70.050 187.040 ;
        RECT 69.850 186.360 70.110 186.680 ;
        RECT 69.910 184.300 70.050 186.360 ;
        RECT 69.850 183.980 70.110 184.300 ;
        RECT 69.850 183.475 70.110 183.620 ;
        RECT 70.370 183.530 70.510 188.060 ;
        RECT 70.830 187.360 70.970 189.080 ;
        RECT 72.210 189.060 72.350 190.780 ;
        RECT 74.050 189.060 74.190 191.800 ;
        RECT 79.510 191.460 79.770 191.780 ;
        RECT 77.510 190.245 79.390 190.615 ;
        RECT 71.230 188.740 71.490 189.060 ;
        RECT 72.150 188.740 72.410 189.060 ;
        RECT 73.990 188.740 74.250 189.060 ;
        RECT 71.290 188.380 71.430 188.740 ;
        RECT 71.230 188.060 71.490 188.380 ;
        RECT 70.770 187.040 71.030 187.360 ;
        RECT 70.830 186.340 70.970 187.040 ;
        RECT 71.680 186.505 71.960 186.875 ;
        RECT 71.690 186.360 71.950 186.505 ;
        RECT 70.770 186.020 71.030 186.340 ;
        RECT 70.830 184.640 70.970 186.020 ;
        RECT 71.230 185.340 71.490 185.660 ;
        RECT 70.770 184.320 71.030 184.640 ;
        RECT 70.770 183.530 71.030 183.620 ;
        RECT 69.840 183.105 70.120 183.475 ;
        RECT 70.370 183.390 71.030 183.530 ;
        RECT 70.770 183.300 71.030 183.390 ;
        RECT 70.770 182.620 71.030 182.940 ;
        RECT 70.830 181.920 70.970 182.620 ;
        RECT 70.770 181.600 71.030 181.920 ;
        RECT 70.770 180.920 71.030 181.240 ;
        RECT 70.310 180.580 70.570 180.900 ;
        RECT 69.850 179.900 70.110 180.220 ;
        RECT 69.910 179.200 70.050 179.900 ;
        RECT 69.850 178.880 70.110 179.200 ;
        RECT 69.850 177.860 70.110 178.180 ;
        RECT 69.910 175.880 70.050 177.860 ;
        RECT 70.370 176.480 70.510 180.580 ;
        RECT 70.830 178.860 70.970 180.920 ;
        RECT 70.770 178.540 71.030 178.860 ;
        RECT 70.830 177.840 70.970 178.540 ;
        RECT 70.770 177.520 71.030 177.840 ;
        RECT 70.310 176.160 70.570 176.480 ;
        RECT 69.910 175.800 70.510 175.880 ;
        RECT 69.910 175.740 70.570 175.800 ;
        RECT 70.310 175.480 70.570 175.740 ;
        RECT 70.310 174.800 70.570 175.120 ;
        RECT 69.850 174.460 70.110 174.780 ;
        RECT 69.910 171.040 70.050 174.460 ;
        RECT 69.850 170.720 70.110 171.040 ;
        RECT 69.910 167.300 70.050 170.720 ;
        RECT 70.370 167.980 70.510 174.800 ;
        RECT 70.770 169.700 71.030 170.020 ;
        RECT 70.830 168.320 70.970 169.700 ;
        RECT 70.770 168.000 71.030 168.320 ;
        RECT 70.310 167.660 70.570 167.980 ;
        RECT 70.370 167.300 70.510 167.660 ;
        RECT 69.850 166.980 70.110 167.300 ;
        RECT 70.310 166.980 70.570 167.300 ;
        RECT 71.290 165.260 71.430 185.340 ;
        RECT 72.210 183.960 72.350 188.740 ;
        RECT 73.070 188.400 73.330 188.720 ;
        RECT 75.830 188.400 76.090 188.720 ;
        RECT 72.150 183.640 72.410 183.960 ;
        RECT 72.610 183.640 72.870 183.960 ;
        RECT 71.690 182.620 71.950 182.940 ;
        RECT 71.750 181.240 71.890 182.620 ;
        RECT 72.150 181.600 72.410 181.920 ;
        RECT 72.210 181.240 72.350 181.600 ;
        RECT 71.690 180.920 71.950 181.240 ;
        RECT 72.150 180.920 72.410 181.240 ;
        RECT 71.690 180.240 71.950 180.560 ;
        RECT 71.750 178.180 71.890 180.240 ;
        RECT 72.210 179.200 72.350 180.920 ;
        RECT 72.150 178.880 72.410 179.200 ;
        RECT 72.210 178.180 72.350 178.880 ;
        RECT 71.690 177.860 71.950 178.180 ;
        RECT 72.150 177.860 72.410 178.180 ;
        RECT 72.670 175.460 72.810 183.640 ;
        RECT 73.130 183.280 73.270 188.400 ;
        RECT 75.890 186.680 76.030 188.400 ;
        RECT 74.450 186.360 74.710 186.680 ;
        RECT 75.830 186.360 76.090 186.680 ;
        RECT 74.510 184.640 74.650 186.360 ;
        RECT 75.370 185.680 75.630 186.000 ;
        RECT 74.450 184.320 74.710 184.640 ;
        RECT 75.430 183.960 75.570 185.680 ;
        RECT 79.570 185.660 79.710 191.460 ;
        RECT 80.490 188.380 80.630 192.140 ;
        RECT 86.470 192.120 86.610 192.480 ;
        RECT 86.410 191.800 86.670 192.120 ;
        RECT 86.870 191.800 87.130 192.120 ;
        RECT 81.350 191.460 81.610 191.780 ;
        RECT 80.430 188.060 80.690 188.380 ;
        RECT 76.750 185.340 77.010 185.660 ;
        RECT 79.510 185.340 79.770 185.660 ;
        RECT 76.810 183.960 76.950 185.340 ;
        RECT 77.510 184.805 79.390 185.175 ;
        RECT 75.370 183.640 75.630 183.960 ;
        RECT 76.750 183.640 77.010 183.960 ;
        RECT 73.530 183.475 73.790 183.620 ;
        RECT 73.070 182.960 73.330 183.280 ;
        RECT 73.520 183.105 73.800 183.475 ;
        RECT 79.570 183.280 79.710 185.340 ;
        RECT 79.510 182.960 79.770 183.280 ;
        RECT 78.130 182.620 78.390 182.940 ;
        RECT 78.190 181.920 78.330 182.620 ;
        RECT 78.130 181.600 78.390 181.920 ;
        RECT 75.370 181.260 75.630 181.580 ;
        RECT 74.450 180.920 74.710 181.240 ;
        RECT 74.510 178.180 74.650 180.920 ;
        RECT 74.450 177.860 74.710 178.180 ;
        RECT 73.990 177.355 74.250 177.500 ;
        RECT 73.980 176.985 74.260 177.355 ;
        RECT 74.910 177.180 75.170 177.500 ;
        RECT 74.450 175.480 74.710 175.800 ;
        RECT 72.610 175.140 72.870 175.460 ;
        RECT 72.150 174.800 72.410 175.120 ;
        RECT 72.210 172.400 72.350 174.800 ;
        RECT 72.150 172.080 72.410 172.400 ;
        RECT 71.690 171.740 71.950 172.060 ;
        RECT 71.750 170.020 71.890 171.740 ;
        RECT 72.670 171.120 72.810 175.140 ;
        RECT 73.990 174.460 74.250 174.780 ;
        RECT 74.050 173.080 74.190 174.460 ;
        RECT 73.990 172.760 74.250 173.080 ;
        RECT 72.670 170.980 74.190 171.120 ;
        RECT 74.510 171.040 74.650 175.480 ;
        RECT 73.530 170.040 73.790 170.360 ;
        RECT 71.690 169.700 71.950 170.020 ;
        RECT 71.750 166.960 71.890 169.700 ;
        RECT 73.590 169.340 73.730 170.040 ;
        RECT 73.530 169.020 73.790 169.340 ;
        RECT 73.590 167.300 73.730 169.020 ;
        RECT 73.530 166.980 73.790 167.300 ;
        RECT 71.690 166.640 71.950 166.960 ;
        RECT 71.230 164.940 71.490 165.260 ;
        RECT 70.770 164.600 71.030 164.920 ;
        RECT 70.830 161.860 70.970 164.600 ;
        RECT 70.770 161.540 71.030 161.860 ;
        RECT 70.310 160.860 70.570 161.180 ;
        RECT 69.390 156.100 69.650 156.420 ;
        RECT 69.850 155.420 70.110 155.740 ;
        RECT 69.390 150.320 69.650 150.640 ;
        RECT 69.450 149.280 69.590 150.320 ;
        RECT 69.910 149.280 70.050 155.420 ;
        RECT 69.390 148.960 69.650 149.280 ;
        RECT 69.850 148.960 70.110 149.280 ;
        RECT 68.930 148.280 69.190 148.600 ;
        RECT 69.390 147.600 69.650 147.920 ;
        RECT 69.450 145.880 69.590 147.600 ;
        RECT 69.850 147.260 70.110 147.580 ;
        RECT 69.390 145.560 69.650 145.880 ;
        RECT 69.450 143.500 69.590 145.560 ;
        RECT 69.390 143.180 69.650 143.500 ;
        RECT 69.910 142.560 70.050 147.260 ;
        RECT 70.370 143.840 70.510 160.860 ;
        RECT 70.830 160.160 70.970 161.540 ;
        RECT 70.770 159.840 71.030 160.160 ;
        RECT 70.770 159.160 71.030 159.480 ;
        RECT 70.830 156.160 70.970 159.160 ;
        RECT 71.290 157.440 71.430 164.940 ;
        RECT 71.750 164.920 71.890 166.640 ;
        RECT 72.150 166.300 72.410 166.620 ;
        RECT 72.210 164.920 72.350 166.300 ;
        RECT 71.690 164.600 71.950 164.920 ;
        RECT 72.150 164.600 72.410 164.920 ;
        RECT 72.610 164.600 72.870 164.920 ;
        RECT 72.670 164.320 72.810 164.600 ;
        RECT 71.690 163.920 71.950 164.240 ;
        RECT 72.210 164.180 72.810 164.320 ;
        RECT 71.750 162.540 71.890 163.920 ;
        RECT 71.690 162.220 71.950 162.540 ;
        RECT 71.750 159.140 71.890 162.220 ;
        RECT 72.210 161.860 72.350 164.180 ;
        RECT 72.610 163.580 72.870 163.900 ;
        RECT 72.150 161.540 72.410 161.860 ;
        RECT 72.210 159.480 72.350 161.540 ;
        RECT 72.150 159.160 72.410 159.480 ;
        RECT 71.690 158.820 71.950 159.140 ;
        RECT 71.690 158.140 71.950 158.460 ;
        RECT 71.230 157.120 71.490 157.440 ;
        RECT 71.290 156.760 71.430 157.120 ;
        RECT 71.230 156.440 71.490 156.760 ;
        RECT 70.830 156.080 71.430 156.160 ;
        RECT 70.830 156.020 71.490 156.080 ;
        RECT 71.230 155.760 71.490 156.020 ;
        RECT 70.770 150.660 71.030 150.980 ;
        RECT 70.310 143.520 70.570 143.840 ;
        RECT 70.310 143.070 70.570 143.160 ;
        RECT 70.830 143.070 70.970 150.660 ;
        RECT 71.230 149.980 71.490 150.300 ;
        RECT 70.310 142.930 70.970 143.070 ;
        RECT 70.310 142.840 70.570 142.930 ;
        RECT 69.910 142.420 70.510 142.560 ;
        RECT 68.470 140.120 68.730 140.440 ;
        RECT 67.090 138.080 67.350 138.400 ;
        RECT 66.170 137.400 66.430 137.720 ;
        RECT 67.550 137.060 67.810 137.380 ;
        RECT 66.170 136.380 66.430 136.700 ;
        RECT 66.230 132.280 66.370 136.380 ;
        RECT 67.610 132.280 67.750 137.060 ;
        RECT 66.170 131.960 66.430 132.280 ;
        RECT 67.550 131.960 67.810 132.280 ;
        RECT 66.170 130.940 66.430 131.260 ;
        RECT 63.410 129.920 63.670 130.240 ;
        RECT 65.710 129.920 65.970 130.240 ;
        RECT 64.790 128.560 65.050 128.880 ;
        RECT 62.510 127.685 64.390 128.055 ;
        RECT 64.850 127.520 64.990 128.560 ;
        RECT 64.790 127.200 65.050 127.520 ;
        RECT 65.770 127.180 65.910 129.920 ;
        RECT 65.710 126.860 65.970 127.180 ;
        RECT 66.230 126.840 66.370 130.940 ;
        RECT 60.650 126.520 60.910 126.840 ;
        RECT 61.570 126.520 61.830 126.840 ;
        RECT 66.170 126.520 66.430 126.840 ;
        RECT 61.110 123.800 61.370 124.120 ;
        RECT 56.970 123.460 57.230 123.780 ;
        RECT 58.810 123.460 59.070 123.780 ;
        RECT 60.190 123.460 60.450 123.780 ;
        RECT 55.590 122.780 55.850 123.100 ;
        RECT 59.730 122.780 59.990 123.100 ;
        RECT 51.450 121.760 51.710 122.080 ;
        RECT 55.130 121.760 55.390 122.080 ;
        RECT 55.650 121.400 55.790 122.780 ;
        RECT 48.230 121.080 48.490 121.400 ;
        RECT 49.610 121.080 49.870 121.400 ;
        RECT 55.590 121.080 55.850 121.400 ;
        RECT 46.850 120.740 47.110 121.060 ;
        RECT 56.970 120.740 57.230 121.060 ;
        RECT 46.910 116.640 47.050 120.740 ;
        RECT 49.610 120.060 49.870 120.380 ;
        RECT 54.210 120.060 54.470 120.380 ;
        RECT 47.510 119.525 49.390 119.895 ;
        RECT 49.670 118.000 49.810 120.060 ;
        RECT 54.270 119.020 54.410 120.060 ;
        RECT 54.210 118.700 54.470 119.020 ;
        RECT 50.530 118.360 50.790 118.680 ;
        RECT 49.610 117.680 49.870 118.000 ;
        RECT 46.850 116.320 47.110 116.640 ;
        RECT 45.470 115.640 45.730 115.960 ;
        RECT 47.510 114.085 49.390 114.455 ;
        RECT 50.590 104.355 50.730 118.360 ;
        RECT 55.590 117.340 55.850 117.660 ;
        RECT 55.650 104.355 55.790 117.340 ;
        RECT 57.030 116.300 57.170 120.740 ;
        RECT 59.790 118.680 59.930 122.780 ;
        RECT 61.170 121.060 61.310 123.800 ;
        RECT 67.090 122.780 67.350 123.100 ;
        RECT 62.510 122.245 64.390 122.615 ;
        RECT 67.150 121.740 67.290 122.780 ;
        RECT 68.530 121.990 68.670 140.120 ;
        RECT 69.850 139.780 70.110 140.100 ;
        RECT 69.910 137.720 70.050 139.780 ;
        RECT 69.850 137.400 70.110 137.720 ;
        RECT 68.930 136.720 69.190 137.040 ;
        RECT 68.990 131.260 69.130 136.720 ;
        RECT 69.850 136.380 70.110 136.700 ;
        RECT 69.390 134.340 69.650 134.660 ;
        RECT 69.450 132.960 69.590 134.340 ;
        RECT 69.910 132.960 70.050 136.380 ;
        RECT 69.390 132.640 69.650 132.960 ;
        RECT 69.850 132.640 70.110 132.960 ;
        RECT 68.930 130.940 69.190 131.260 ;
        RECT 69.390 128.900 69.650 129.220 ;
        RECT 69.450 127.520 69.590 128.900 ;
        RECT 69.390 127.200 69.650 127.520 ;
        RECT 70.370 123.780 70.510 142.420 ;
        RECT 70.830 140.440 70.970 142.930 ;
        RECT 70.770 140.120 71.030 140.440 ;
        RECT 70.830 134.660 70.970 140.120 ;
        RECT 70.770 134.340 71.030 134.660 ;
        RECT 70.830 129.220 70.970 134.340 ;
        RECT 70.770 128.900 71.030 129.220 ;
        RECT 70.770 128.220 71.030 128.540 ;
        RECT 70.830 127.520 70.970 128.220 ;
        RECT 70.770 127.200 71.030 127.520 ;
        RECT 70.310 123.460 70.570 123.780 ;
        RECT 69.390 121.990 69.650 122.080 ;
        RECT 68.530 121.850 69.650 121.990 ;
        RECT 69.390 121.760 69.650 121.850 ;
        RECT 62.030 121.420 62.290 121.740 ;
        RECT 67.090 121.420 67.350 121.740 ;
        RECT 60.650 120.740 60.910 121.060 ;
        RECT 61.110 120.740 61.370 121.060 ;
        RECT 59.730 118.360 59.990 118.680 ;
        RECT 57.430 117.680 57.690 118.000 ;
        RECT 57.490 116.640 57.630 117.680 ;
        RECT 57.430 116.320 57.690 116.640 ;
        RECT 56.970 115.980 57.230 116.300 ;
        RECT 60.710 104.355 60.850 120.740 ;
        RECT 61.170 118.340 61.310 120.740 ;
        RECT 61.110 118.020 61.370 118.340 ;
        RECT 62.090 116.640 62.230 121.420 ;
        RECT 71.290 121.400 71.430 149.980 ;
        RECT 71.750 148.600 71.890 158.140 ;
        RECT 72.150 155.420 72.410 155.740 ;
        RECT 72.210 154.380 72.350 155.420 ;
        RECT 72.150 154.060 72.410 154.380 ;
        RECT 72.670 150.980 72.810 163.580 ;
        RECT 73.070 160.860 73.330 161.180 ;
        RECT 72.610 150.660 72.870 150.980 ;
        RECT 71.690 148.280 71.950 148.600 ;
        RECT 71.690 145.900 71.950 146.220 ;
        RECT 71.750 143.160 71.890 145.900 ;
        RECT 73.130 145.280 73.270 160.860 ;
        RECT 73.590 159.480 73.730 166.980 ;
        RECT 73.530 159.160 73.790 159.480 ;
        RECT 74.050 157.100 74.190 170.980 ;
        RECT 74.450 170.720 74.710 171.040 ;
        RECT 74.970 170.440 75.110 177.180 ;
        RECT 74.510 170.300 75.110 170.440 ;
        RECT 73.990 156.780 74.250 157.100 ;
        RECT 74.050 154.040 74.190 156.780 ;
        RECT 73.990 153.720 74.250 154.040 ;
        RECT 73.530 151.680 73.790 152.000 ;
        RECT 72.670 145.140 73.270 145.280 ;
        RECT 71.690 142.840 71.950 143.160 ;
        RECT 72.150 142.840 72.410 143.160 ;
        RECT 71.680 142.305 71.960 142.675 ;
        RECT 71.690 142.160 71.950 142.305 ;
        RECT 72.210 142.140 72.350 142.840 ;
        RECT 72.150 141.820 72.410 142.140 ;
        RECT 71.690 138.080 71.950 138.400 ;
        RECT 71.750 132.960 71.890 138.080 ;
        RECT 72.670 137.720 72.810 145.140 ;
        RECT 73.590 141.120 73.730 151.680 ;
        RECT 73.990 151.340 74.250 151.660 ;
        RECT 74.050 148.510 74.190 151.340 ;
        RECT 74.510 151.320 74.650 170.300 ;
        RECT 74.910 166.300 75.170 166.620 ;
        RECT 74.970 164.920 75.110 166.300 ;
        RECT 74.910 164.600 75.170 164.920 ;
        RECT 74.910 159.160 75.170 159.480 ;
        RECT 74.970 156.760 75.110 159.160 ;
        RECT 74.910 156.440 75.170 156.760 ;
        RECT 74.450 151.000 74.710 151.320 ;
        RECT 74.450 148.510 74.710 148.600 ;
        RECT 74.050 148.370 74.710 148.510 ;
        RECT 74.450 148.280 74.710 148.370 ;
        RECT 74.510 145.540 74.650 148.280 ;
        RECT 74.450 145.220 74.710 145.540 ;
        RECT 74.510 142.675 74.650 145.220 ;
        RECT 74.910 144.540 75.170 144.860 ;
        RECT 74.970 143.500 75.110 144.540 ;
        RECT 74.910 143.180 75.170 143.500 ;
        RECT 75.430 142.820 75.570 181.260 ;
        RECT 76.290 180.580 76.550 180.900 ;
        RECT 75.830 178.880 76.090 179.200 ;
        RECT 75.890 178.180 76.030 178.880 ;
        RECT 76.350 178.180 76.490 180.580 ;
        RECT 77.510 179.365 79.390 179.735 ;
        RECT 79.570 178.860 79.710 182.960 ;
        RECT 79.510 178.540 79.770 178.860 ;
        RECT 80.490 178.180 80.630 188.060 ;
        RECT 81.410 183.960 81.550 191.460 ;
        RECT 83.190 190.780 83.450 191.100 ;
        RECT 85.490 190.780 85.750 191.100 ;
        RECT 83.250 188.720 83.390 190.780 ;
        RECT 85.550 189.400 85.690 190.780 ;
        RECT 85.490 189.080 85.750 189.400 ;
        RECT 83.190 188.400 83.450 188.720 ;
        RECT 86.930 186.680 87.070 191.800 ;
        RECT 87.390 189.060 87.530 194.180 ;
        RECT 88.710 191.460 88.970 191.780 ;
        RECT 88.770 189.400 88.910 191.460 ;
        RECT 88.710 189.080 88.970 189.400 ;
        RECT 87.330 188.740 87.590 189.060 ;
        RECT 87.790 188.740 88.050 189.060 ;
        RECT 86.870 186.360 87.130 186.680 ;
        RECT 84.570 186.020 84.830 186.340 ;
        RECT 84.630 184.640 84.770 186.020 ;
        RECT 86.410 185.340 86.670 185.660 ;
        RECT 84.570 184.320 84.830 184.640 ;
        RECT 86.470 183.960 86.610 185.340 ;
        RECT 81.350 183.640 81.610 183.960 ;
        RECT 86.410 183.640 86.670 183.960 ;
        RECT 84.570 183.300 84.830 183.620 ;
        RECT 84.110 182.620 84.370 182.940 ;
        RECT 83.650 181.260 83.910 181.580 ;
        RECT 83.710 178.860 83.850 181.260 ;
        RECT 83.650 178.540 83.910 178.860 ;
        RECT 84.170 178.520 84.310 182.620 ;
        RECT 84.630 179.200 84.770 183.300 ;
        RECT 86.930 183.190 87.070 186.360 ;
        RECT 87.390 186.340 87.530 188.740 ;
        RECT 87.330 186.020 87.590 186.340 ;
        RECT 86.470 183.050 87.070 183.190 ;
        RECT 85.950 182.620 86.210 182.940 ;
        RECT 86.010 181.580 86.150 182.620 ;
        RECT 85.950 181.260 86.210 181.580 ;
        RECT 84.570 178.880 84.830 179.200 ;
        RECT 84.110 178.200 84.370 178.520 ;
        RECT 86.470 178.180 86.610 183.050 ;
        RECT 87.390 180.900 87.530 186.020 ;
        RECT 87.850 185.660 87.990 188.740 ;
        RECT 88.710 187.040 88.970 187.360 ;
        RECT 87.790 185.340 88.050 185.660 ;
        RECT 88.770 183.620 88.910 187.040 ;
        RECT 88.710 183.300 88.970 183.620 ;
        RECT 88.710 182.620 88.970 182.940 ;
        RECT 87.780 181.065 88.060 181.435 ;
        RECT 87.330 180.810 87.590 180.900 ;
        RECT 86.930 180.670 87.590 180.810 ;
        RECT 75.830 177.860 76.090 178.180 ;
        RECT 76.290 177.860 76.550 178.180 ;
        RECT 80.430 177.860 80.690 178.180 ;
        RECT 86.410 177.860 86.670 178.180 ;
        RECT 85.030 177.520 85.290 177.840 ;
        RECT 80.430 175.480 80.690 175.800 ;
        RECT 79.510 174.460 79.770 174.780 ;
        RECT 77.510 173.925 79.390 174.295 ;
        RECT 79.570 170.700 79.710 174.460 ;
        RECT 80.490 173.955 80.630 175.480 ;
        RECT 80.420 173.585 80.700 173.955 ;
        RECT 83.650 172.420 83.910 172.740 ;
        RECT 79.510 170.380 79.770 170.700 ;
        RECT 75.830 169.700 76.090 170.020 ;
        RECT 75.890 165.600 76.030 169.700 ;
        RECT 83.190 169.020 83.450 169.340 ;
        RECT 77.510 168.485 79.390 168.855 ;
        RECT 78.590 167.320 78.850 167.640 ;
        RECT 76.750 166.300 77.010 166.620 ;
        RECT 75.830 165.280 76.090 165.600 ;
        RECT 76.810 164.920 76.950 166.300 ;
        RECT 76.750 164.600 77.010 164.920 ;
        RECT 76.810 162.200 76.950 164.600 ;
        RECT 78.650 164.580 78.790 167.320 ;
        RECT 79.510 166.640 79.770 166.960 ;
        RECT 79.570 164.920 79.710 166.640 ;
        RECT 79.510 164.600 79.770 164.920 ;
        RECT 78.590 164.260 78.850 164.580 ;
        RECT 77.510 163.045 79.390 163.415 ;
        RECT 79.570 162.880 79.710 164.600 ;
        RECT 82.730 163.920 82.990 164.240 ;
        RECT 79.970 163.580 80.230 163.900 ;
        RECT 79.510 162.560 79.770 162.880 ;
        RECT 76.750 161.880 77.010 162.200 ;
        RECT 79.050 161.200 79.310 161.520 ;
        RECT 78.590 160.860 78.850 161.180 ;
        RECT 78.650 158.800 78.790 160.860 ;
        RECT 79.110 159.820 79.250 161.200 ;
        RECT 79.050 159.500 79.310 159.820 ;
        RECT 80.030 159.480 80.170 163.580 ;
        RECT 82.790 162.880 82.930 163.920 ;
        RECT 83.250 163.900 83.390 169.020 ;
        RECT 83.190 163.580 83.450 163.900 ;
        RECT 82.730 162.560 82.990 162.880 ;
        RECT 83.710 162.200 83.850 172.420 ;
        RECT 84.110 169.020 84.370 169.340 ;
        RECT 84.170 167.640 84.310 169.020 ;
        RECT 85.090 167.720 85.230 177.520 ;
        RECT 86.930 174.780 87.070 180.670 ;
        RECT 87.330 180.580 87.590 180.670 ;
        RECT 87.850 179.960 87.990 181.065 ;
        RECT 87.390 179.820 87.990 179.960 ;
        RECT 86.870 174.460 87.130 174.780 ;
        RECT 86.930 172.740 87.070 174.460 ;
        RECT 86.870 172.420 87.130 172.740 ;
        RECT 85.490 169.700 85.750 170.020 ;
        RECT 85.550 169.340 85.690 169.700 ;
        RECT 85.490 169.020 85.750 169.340 ;
        RECT 84.630 167.640 85.230 167.720 ;
        RECT 84.110 167.320 84.370 167.640 ;
        RECT 84.570 167.580 85.230 167.640 ;
        RECT 84.570 167.320 84.830 167.580 ;
        RECT 85.950 166.300 86.210 166.620 ;
        RECT 85.030 164.940 85.290 165.260 ;
        RECT 85.090 162.880 85.230 164.940 ;
        RECT 85.030 162.560 85.290 162.880 ;
        RECT 83.650 161.880 83.910 162.200 ;
        RECT 86.010 161.860 86.150 166.300 ;
        RECT 81.810 161.540 82.070 161.860 ;
        RECT 85.950 161.540 86.210 161.860 ;
        RECT 81.870 160.160 82.010 161.540 ;
        RECT 83.190 161.200 83.450 161.520 ;
        RECT 81.810 159.840 82.070 160.160 ;
        RECT 82.730 159.840 82.990 160.160 ;
        RECT 79.970 159.160 80.230 159.480 ;
        RECT 82.270 159.160 82.530 159.480 ;
        RECT 78.590 158.480 78.850 158.800 ;
        RECT 77.510 157.605 79.390 157.975 ;
        RECT 79.970 156.100 80.230 156.420 ;
        RECT 78.130 155.420 78.390 155.740 ;
        RECT 78.190 154.380 78.330 155.420 ;
        RECT 78.130 154.060 78.390 154.380 ;
        RECT 79.510 152.700 79.770 153.020 ;
        RECT 77.510 152.165 79.390 152.535 ;
        RECT 75.830 150.660 76.090 150.980 ;
        RECT 78.590 150.660 78.850 150.980 ;
        RECT 75.890 148.940 76.030 150.660 ;
        RECT 75.830 148.620 76.090 148.940 ;
        RECT 75.890 145.540 76.030 148.620 ;
        RECT 78.650 148.260 78.790 150.660 ;
        RECT 79.570 150.640 79.710 152.700 ;
        RECT 79.510 150.320 79.770 150.640 ;
        RECT 80.030 148.600 80.170 156.100 ;
        RECT 82.330 152.000 82.470 159.160 ;
        RECT 82.790 156.760 82.930 159.840 ;
        RECT 83.250 159.820 83.390 161.200 ;
        RECT 83.190 159.500 83.450 159.820 ;
        RECT 84.570 158.140 84.830 158.460 ;
        RECT 82.730 156.440 82.990 156.760 ;
        RECT 83.650 155.420 83.910 155.740 ;
        RECT 82.270 151.680 82.530 152.000 ;
        RECT 83.710 150.640 83.850 155.420 ;
        RECT 84.630 154.040 84.770 158.140 ;
        RECT 87.390 156.760 87.530 179.820 ;
        RECT 87.790 177.860 88.050 178.180 ;
        RECT 87.850 172.740 87.990 177.860 ;
        RECT 88.250 177.180 88.510 177.500 ;
        RECT 88.310 176.140 88.450 177.180 ;
        RECT 88.250 175.820 88.510 176.140 ;
        RECT 88.250 175.140 88.510 175.460 ;
        RECT 87.790 172.420 88.050 172.740 ;
        RECT 88.310 172.400 88.450 175.140 ;
        RECT 88.250 172.080 88.510 172.400 ;
        RECT 88.310 171.040 88.450 172.080 ;
        RECT 88.250 170.720 88.510 171.040 ;
        RECT 87.790 164.260 88.050 164.580 ;
        RECT 87.850 162.880 87.990 164.260 ;
        RECT 87.790 162.560 88.050 162.880 ;
        RECT 88.310 161.520 88.450 170.720 ;
        RECT 88.250 161.200 88.510 161.520 ;
        RECT 88.250 157.120 88.510 157.440 ;
        RECT 85.030 156.440 85.290 156.760 ;
        RECT 87.330 156.440 87.590 156.760 ;
        RECT 85.090 154.720 85.230 156.440 ;
        RECT 87.790 155.420 88.050 155.740 ;
        RECT 85.030 154.400 85.290 154.720 ;
        RECT 84.570 153.720 84.830 154.040 ;
        RECT 85.090 152.880 85.230 154.400 ;
        RECT 87.850 154.040 87.990 155.420 ;
        RECT 87.790 153.720 88.050 154.040 ;
        RECT 86.410 153.380 86.670 153.700 ;
        RECT 85.090 152.740 85.690 152.880 ;
        RECT 85.550 151.320 85.690 152.740 ;
        RECT 85.490 151.000 85.750 151.320 ;
        RECT 83.650 150.320 83.910 150.640 ;
        RECT 80.890 149.980 81.150 150.300 ;
        RECT 79.970 148.280 80.230 148.600 ;
        RECT 78.590 147.940 78.850 148.260 ;
        RECT 77.510 146.725 79.390 147.095 ;
        RECT 78.130 145.900 78.390 146.220 ;
        RECT 75.830 145.220 76.090 145.540 ;
        RECT 74.440 142.305 74.720 142.675 ;
        RECT 75.370 142.500 75.630 142.820 ;
        RECT 75.890 142.480 76.030 145.220 ;
        RECT 78.190 143.840 78.330 145.900 ;
        RECT 80.950 145.540 81.090 149.980 ;
        RECT 83.650 147.940 83.910 148.260 ;
        RECT 80.890 145.220 81.150 145.540 ;
        RECT 81.350 144.880 81.610 145.200 ;
        RECT 81.410 143.840 81.550 144.880 ;
        RECT 78.130 143.520 78.390 143.840 ;
        RECT 81.350 143.520 81.610 143.840 ;
        RECT 83.190 143.180 83.450 143.500 ;
        RECT 75.830 142.160 76.090 142.480 ;
        RECT 73.990 141.820 74.250 142.140 ;
        RECT 74.910 141.820 75.170 142.140 ;
        RECT 76.750 141.820 77.010 142.140 ;
        RECT 73.530 140.800 73.790 141.120 ;
        RECT 73.530 139.440 73.790 139.760 ;
        RECT 73.060 138.225 73.340 138.595 ;
        RECT 73.130 137.720 73.270 138.225 ;
        RECT 72.610 137.400 72.870 137.720 ;
        RECT 73.070 137.400 73.330 137.720 ;
        RECT 73.590 137.040 73.730 139.440 ;
        RECT 74.050 138.060 74.190 141.820 ;
        RECT 73.990 137.740 74.250 138.060 ;
        RECT 74.970 137.380 75.110 141.820 ;
        RECT 76.290 137.400 76.550 137.720 ;
        RECT 74.910 137.060 75.170 137.380 ;
        RECT 72.150 136.720 72.410 137.040 ;
        RECT 73.530 136.720 73.790 137.040 ;
        RECT 71.690 132.640 71.950 132.960 ;
        RECT 71.750 129.900 71.890 132.640 ;
        RECT 71.690 129.580 71.950 129.900 ;
        RECT 72.210 121.740 72.350 136.720 ;
        RECT 73.590 132.280 73.730 136.720 ;
        RECT 76.350 135.680 76.490 137.400 ;
        RECT 76.290 135.360 76.550 135.680 ;
        RECT 74.450 134.000 74.710 134.320 ;
        RECT 73.530 131.960 73.790 132.280 ;
        RECT 73.590 131.600 73.730 131.960 ;
        RECT 73.530 131.280 73.790 131.600 ;
        RECT 74.510 127.520 74.650 134.000 ;
        RECT 76.290 132.300 76.550 132.620 ;
        RECT 75.830 131.680 76.090 131.940 ;
        RECT 76.350 131.680 76.490 132.300 ;
        RECT 75.830 131.620 76.490 131.680 ;
        RECT 75.890 131.540 76.490 131.620 ;
        RECT 76.350 127.520 76.490 131.540 ;
        RECT 74.450 127.200 74.710 127.520 ;
        RECT 76.290 127.200 76.550 127.520 ;
        RECT 73.990 125.500 74.250 125.820 ;
        RECT 72.150 121.420 72.410 121.740 ;
        RECT 74.050 121.400 74.190 125.500 ;
        RECT 76.810 122.080 76.950 141.820 ;
        RECT 77.510 141.285 79.390 141.655 ;
        RECT 83.250 141.120 83.390 143.180 ;
        RECT 83.710 142.560 83.850 147.940 ;
        RECT 85.550 146.220 85.690 151.000 ;
        RECT 86.470 148.600 86.610 153.380 ;
        RECT 87.790 149.980 88.050 150.300 ;
        RECT 87.850 148.600 87.990 149.980 ;
        RECT 86.410 148.280 86.670 148.600 ;
        RECT 87.790 148.280 88.050 148.600 ;
        RECT 85.490 145.900 85.750 146.220 ;
        RECT 87.790 145.220 88.050 145.540 ;
        RECT 84.570 144.540 84.830 144.860 ;
        RECT 84.630 143.160 84.770 144.540 ;
        RECT 84.570 142.840 84.830 143.160 ;
        RECT 85.490 142.730 85.750 142.820 ;
        RECT 85.090 142.590 85.750 142.730 ;
        RECT 83.710 142.420 84.770 142.560 ;
        RECT 83.190 140.800 83.450 141.120 ;
        RECT 80.880 140.265 81.160 140.635 ;
        RECT 80.950 140.100 81.090 140.265 ;
        RECT 84.630 140.100 84.770 142.420 ;
        RECT 80.890 139.780 81.150 140.100 ;
        RECT 82.730 139.780 82.990 140.100 ;
        RECT 84.570 139.780 84.830 140.100 ;
        RECT 82.790 137.720 82.930 139.780 ;
        RECT 84.630 138.060 84.770 139.780 ;
        RECT 84.570 137.740 84.830 138.060 ;
        RECT 82.730 137.400 82.990 137.720 ;
        RECT 85.090 137.380 85.230 142.590 ;
        RECT 85.490 142.500 85.750 142.590 ;
        RECT 87.320 140.265 87.600 140.635 ;
        RECT 87.390 139.760 87.530 140.265 ;
        RECT 87.330 139.440 87.590 139.760 ;
        RECT 85.490 137.740 85.750 138.060 ;
        RECT 84.570 137.060 84.830 137.380 ;
        RECT 85.030 137.060 85.290 137.380 ;
        RECT 79.970 136.380 80.230 136.700 ;
        RECT 77.510 135.845 79.390 136.215 ;
        RECT 79.050 132.870 79.310 132.960 ;
        RECT 79.050 132.730 79.710 132.870 ;
        RECT 79.050 132.640 79.310 132.730 ;
        RECT 77.510 130.405 79.390 130.775 ;
        RECT 77.510 124.965 79.390 125.335 ;
        RECT 79.570 123.780 79.710 132.730 ;
        RECT 80.030 132.620 80.170 136.380 ;
        RECT 82.730 134.680 82.990 135.000 ;
        RECT 82.790 132.960 82.930 134.680 ;
        RECT 82.730 132.640 82.990 132.960 ;
        RECT 79.970 132.300 80.230 132.620 ;
        RECT 84.630 132.180 84.770 137.060 ;
        RECT 85.090 134.660 85.230 137.060 ;
        RECT 85.550 134.660 85.690 137.740 ;
        RECT 85.030 134.340 85.290 134.660 ;
        RECT 85.490 134.340 85.750 134.660 ;
        RECT 84.630 132.040 85.230 132.180 ;
        RECT 81.350 131.620 81.610 131.940 ;
        RECT 79.970 130.940 80.230 131.260 ;
        RECT 80.030 129.560 80.170 130.940 ;
        RECT 81.410 130.240 81.550 131.620 ;
        RECT 83.650 131.280 83.910 131.600 ;
        RECT 84.570 131.280 84.830 131.600 ;
        RECT 81.350 129.920 81.610 130.240 ;
        RECT 79.970 129.240 80.230 129.560 ;
        RECT 83.710 128.540 83.850 131.280 ;
        RECT 84.630 129.560 84.770 131.280 ;
        RECT 85.090 129.900 85.230 132.040 ;
        RECT 85.490 131.960 85.750 132.280 ;
        RECT 85.030 129.580 85.290 129.900 ;
        RECT 84.570 129.240 84.830 129.560 ;
        RECT 84.110 128.560 84.370 128.880 ;
        RECT 80.430 128.220 80.690 128.540 ;
        RECT 83.650 128.220 83.910 128.540 ;
        RECT 80.490 127.180 80.630 128.220 ;
        RECT 83.710 127.520 83.850 128.220 ;
        RECT 83.650 127.200 83.910 127.520 ;
        RECT 80.430 126.860 80.690 127.180 ;
        RECT 84.170 126.840 84.310 128.560 ;
        RECT 85.550 127.180 85.690 131.960 ;
        RECT 87.850 131.600 87.990 145.220 ;
        RECT 88.310 141.120 88.450 157.120 ;
        RECT 88.770 148.600 88.910 182.620 ;
        RECT 89.230 181.240 89.370 194.520 ;
        RECT 89.690 194.500 89.830 198.940 ;
        RECT 91.070 196.540 91.210 199.620 ;
        RECT 92.510 198.405 94.390 198.775 ;
        RECT 95.670 197.900 95.810 201.660 ;
        RECT 97.050 200.960 97.190 202.680 ;
        RECT 98.370 201.660 98.630 201.980 ;
        RECT 99.290 201.660 99.550 201.980 ;
        RECT 101.130 201.660 101.390 201.980 ;
        RECT 96.990 200.640 97.250 200.960 ;
        RECT 97.450 199.620 97.710 199.940 ;
        RECT 95.610 197.580 95.870 197.900 ;
        RECT 90.550 196.220 90.810 196.540 ;
        RECT 91.010 196.220 91.270 196.540 ;
        RECT 89.630 194.180 89.890 194.500 ;
        RECT 90.610 191.780 90.750 196.220 ;
        RECT 90.550 191.460 90.810 191.780 ;
        RECT 91.070 191.440 91.210 196.220 ;
        RECT 96.990 194.520 97.250 194.840 ;
        RECT 94.690 193.840 94.950 194.160 ;
        RECT 92.510 192.965 94.390 193.335 ;
        RECT 94.750 192.800 94.890 193.840 ;
        RECT 94.690 192.480 94.950 192.800 ;
        RECT 94.230 191.460 94.490 191.780 ;
        RECT 96.530 191.460 96.790 191.780 ;
        RECT 91.010 191.120 91.270 191.440 ;
        RECT 94.290 189.400 94.430 191.460 ;
        RECT 94.230 189.080 94.490 189.400 ;
        RECT 96.070 188.060 96.330 188.380 ;
        RECT 92.510 187.525 94.390 187.895 ;
        RECT 95.150 187.040 95.410 187.360 ;
        RECT 92.850 184.320 93.110 184.640 ;
        RECT 90.090 183.980 90.350 184.300 ;
        RECT 89.630 183.300 89.890 183.620 ;
        RECT 89.690 181.240 89.830 183.300 ;
        RECT 89.170 180.920 89.430 181.240 ;
        RECT 89.630 180.920 89.890 181.240 ;
        RECT 90.150 173.760 90.290 183.980 ;
        RECT 92.910 183.620 93.050 184.320 ;
        RECT 95.210 183.960 95.350 187.040 ;
        RECT 95.150 183.640 95.410 183.960 ;
        RECT 96.130 183.620 96.270 188.060 ;
        RECT 96.590 183.960 96.730 191.460 ;
        RECT 97.050 187.360 97.190 194.520 ;
        RECT 97.510 192.800 97.650 199.620 ;
        RECT 98.430 197.900 98.570 201.660 ;
        RECT 98.830 200.640 99.090 200.960 ;
        RECT 98.370 197.580 98.630 197.900 ;
        RECT 98.890 195.520 99.030 200.640 ;
        RECT 98.830 195.200 99.090 195.520 ;
        RECT 98.370 194.180 98.630 194.500 ;
        RECT 97.450 192.480 97.710 192.800 ;
        RECT 96.990 187.040 97.250 187.360 ;
        RECT 97.910 185.680 98.170 186.000 ;
        RECT 96.530 183.640 96.790 183.960 ;
        RECT 91.470 183.475 91.730 183.620 ;
        RECT 90.550 182.960 90.810 183.280 ;
        RECT 91.460 183.105 91.740 183.475 ;
        RECT 92.850 183.300 93.110 183.620 ;
        RECT 93.310 183.300 93.570 183.620 ;
        RECT 96.070 183.300 96.330 183.620 ;
        RECT 90.610 181.240 90.750 182.960 ;
        RECT 91.010 181.600 91.270 181.920 ;
        RECT 90.550 180.920 90.810 181.240 ;
        RECT 90.550 177.860 90.810 178.180 ;
        RECT 90.090 173.440 90.350 173.760 ;
        RECT 90.610 173.420 90.750 177.860 ;
        RECT 89.170 173.100 89.430 173.420 ;
        RECT 90.550 173.100 90.810 173.420 ;
        RECT 89.230 164.920 89.370 173.100 ;
        RECT 90.090 172.080 90.350 172.400 ;
        RECT 89.630 169.020 89.890 169.340 ;
        RECT 89.690 167.640 89.830 169.020 ;
        RECT 89.630 167.320 89.890 167.640 ;
        RECT 89.690 164.920 89.830 167.320 ;
        RECT 90.150 166.960 90.290 172.080 ;
        RECT 90.090 166.640 90.350 166.960 ;
        RECT 90.610 165.260 90.750 173.100 ;
        RECT 91.070 167.300 91.210 181.600 ;
        RECT 91.530 181.580 91.670 183.105 ;
        RECT 93.370 182.940 93.510 183.300 ;
        RECT 93.310 182.620 93.570 182.940 ;
        RECT 92.510 182.085 94.390 182.455 ;
        RECT 96.060 182.425 96.340 182.795 ;
        RECT 96.530 182.620 96.790 182.940 ;
        RECT 91.470 181.260 91.730 181.580 ;
        RECT 95.150 180.920 95.410 181.240 ;
        RECT 91.930 180.580 92.190 180.900 ;
        RECT 91.460 172.905 91.740 173.275 ;
        RECT 91.530 170.700 91.670 172.905 ;
        RECT 91.470 170.380 91.730 170.700 ;
        RECT 91.990 169.930 92.130 180.580 ;
        RECT 94.690 180.240 94.950 180.560 ;
        RECT 94.750 178.180 94.890 180.240 ;
        RECT 94.690 177.860 94.950 178.180 ;
        RECT 92.510 176.645 94.390 177.015 ;
        RECT 92.510 171.205 94.390 171.575 ;
        RECT 94.750 170.020 94.890 177.860 ;
        RECT 95.210 176.480 95.350 180.920 ;
        RECT 95.610 180.580 95.870 180.900 ;
        RECT 95.670 179.200 95.810 180.580 ;
        RECT 95.610 178.880 95.870 179.200 ;
        RECT 96.130 178.600 96.270 182.425 ;
        RECT 95.670 178.460 96.270 178.600 ;
        RECT 95.150 176.160 95.410 176.480 ;
        RECT 91.530 169.790 92.130 169.930 ;
        RECT 91.010 166.980 91.270 167.300 ;
        RECT 90.550 164.940 90.810 165.260 ;
        RECT 89.170 164.600 89.430 164.920 ;
        RECT 89.630 164.600 89.890 164.920 ;
        RECT 89.690 159.140 89.830 164.600 ;
        RECT 91.010 163.580 91.270 163.900 ;
        RECT 90.550 162.220 90.810 162.540 ;
        RECT 90.090 159.500 90.350 159.820 ;
        RECT 89.630 158.820 89.890 159.140 ;
        RECT 89.160 157.945 89.440 158.315 ;
        RECT 89.230 156.420 89.370 157.945 ;
        RECT 89.170 156.100 89.430 156.420 ;
        RECT 90.150 154.720 90.290 159.500 ;
        RECT 90.610 156.760 90.750 162.220 ;
        RECT 91.070 161.860 91.210 163.580 ;
        RECT 91.010 161.540 91.270 161.860 ;
        RECT 91.010 160.860 91.270 161.180 ;
        RECT 90.550 156.440 90.810 156.760 ;
        RECT 90.550 155.420 90.810 155.740 ;
        RECT 90.090 154.400 90.350 154.720 ;
        RECT 89.630 152.700 89.890 153.020 ;
        RECT 88.710 148.280 88.970 148.600 ;
        RECT 89.690 148.260 89.830 152.700 ;
        RECT 89.630 147.940 89.890 148.260 ;
        RECT 90.090 147.600 90.350 147.920 ;
        RECT 89.630 147.260 89.890 147.580 ;
        RECT 89.690 146.560 89.830 147.260 ;
        RECT 89.630 146.240 89.890 146.560 ;
        RECT 88.710 145.220 88.970 145.540 ;
        RECT 88.250 140.800 88.510 141.120 ;
        RECT 88.770 140.780 88.910 145.220 ;
        RECT 89.630 143.180 89.890 143.500 ;
        RECT 88.710 140.460 88.970 140.780 ;
        RECT 89.690 139.840 89.830 143.180 ;
        RECT 90.150 141.120 90.290 147.600 ;
        RECT 90.090 140.800 90.350 141.120 ;
        RECT 89.230 139.700 89.830 139.840 ;
        RECT 88.710 137.740 88.970 138.060 ;
        RECT 88.770 135.680 88.910 137.740 ;
        RECT 89.230 135.680 89.370 139.700 ;
        RECT 89.630 137.060 89.890 137.380 ;
        RECT 89.690 135.680 89.830 137.060 ;
        RECT 88.710 135.360 88.970 135.680 ;
        RECT 89.170 135.360 89.430 135.680 ;
        RECT 89.630 135.360 89.890 135.680 ;
        RECT 88.710 134.340 88.970 134.660 ;
        RECT 88.770 132.960 88.910 134.340 ;
        RECT 88.710 132.640 88.970 132.960 ;
        RECT 88.250 132.300 88.510 132.620 ;
        RECT 87.790 131.280 88.050 131.600 ;
        RECT 87.850 128.960 87.990 131.280 ;
        RECT 88.310 130.240 88.450 132.300 ;
        RECT 88.250 129.920 88.510 130.240 ;
        RECT 87.850 128.880 88.450 128.960 ;
        RECT 87.850 128.820 88.510 128.880 ;
        RECT 88.250 128.560 88.510 128.820 ;
        RECT 85.490 126.860 85.750 127.180 ;
        RECT 84.110 126.520 84.370 126.840 ;
        RECT 79.970 126.180 80.230 126.500 ;
        RECT 80.030 124.800 80.170 126.180 ;
        RECT 79.970 124.480 80.230 124.800 ;
        RECT 79.510 123.460 79.770 123.780 ;
        RECT 79.970 123.120 80.230 123.440 ;
        RECT 76.750 121.760 77.010 122.080 ;
        RECT 75.830 121.420 76.090 121.740 ;
        RECT 71.230 121.080 71.490 121.400 ;
        RECT 73.990 121.080 74.250 121.400 ;
        RECT 75.370 120.740 75.630 121.060 ;
        RECT 70.770 120.060 71.030 120.380 ;
        RECT 71.230 120.060 71.490 120.380 ;
        RECT 72.610 120.060 72.870 120.380 ;
        RECT 70.830 118.680 70.970 120.060 ;
        RECT 70.770 118.360 71.030 118.680 ;
        RECT 65.250 118.020 65.510 118.340 ;
        RECT 62.510 116.805 64.390 117.175 ;
        RECT 65.310 116.640 65.450 118.020 ;
        RECT 65.710 117.340 65.970 117.660 ;
        RECT 62.030 116.320 62.290 116.640 ;
        RECT 65.250 116.320 65.510 116.640 ;
        RECT 65.770 104.355 65.910 117.340 ;
        RECT 71.290 116.300 71.430 120.060 ;
        RECT 72.670 118.680 72.810 120.060 ;
        RECT 72.610 118.360 72.870 118.680 ;
        RECT 72.610 117.680 72.870 118.000 ;
        RECT 73.530 117.680 73.790 118.000 ;
        RECT 71.230 115.980 71.490 116.300 ;
        RECT 70.830 104.355 71.430 104.480 ;
        RECT 45.460 103.800 45.740 104.355 ;
        RECT 44.150 103.660 45.740 103.800 ;
        RECT 45.460 102.355 45.740 103.660 ;
        RECT 50.520 102.355 50.800 104.355 ;
        RECT 55.580 102.355 55.860 104.355 ;
        RECT 60.640 102.355 60.920 104.355 ;
        RECT 65.700 102.355 65.980 104.355 ;
        RECT 70.760 104.340 71.430 104.355 ;
        RECT 70.760 102.355 71.040 104.340 ;
        RECT 71.290 103.800 71.430 104.340 ;
        RECT 72.670 103.800 72.810 117.680 ;
        RECT 73.590 116.640 73.730 117.680 ;
        RECT 73.530 116.320 73.790 116.640 ;
        RECT 75.430 116.040 75.570 120.740 ;
        RECT 75.890 116.640 76.030 121.420 ;
        RECT 77.510 119.525 79.390 119.895 ;
        RECT 76.750 117.340 77.010 117.660 ;
        RECT 75.830 116.320 76.090 116.640 ;
        RECT 75.430 115.900 76.030 116.040 ;
        RECT 76.810 115.960 76.950 117.340 ;
        RECT 75.890 104.355 76.030 115.900 ;
        RECT 76.750 115.640 77.010 115.960 ;
        RECT 80.030 114.940 80.170 123.120 ;
        RECT 83.650 122.780 83.910 123.100 ;
        RECT 83.710 121.740 83.850 122.780 ;
        RECT 84.170 121.740 84.310 126.520 ;
        RECT 90.610 124.120 90.750 155.420 ;
        RECT 91.070 148.600 91.210 160.860 ;
        RECT 91.530 156.760 91.670 169.790 ;
        RECT 94.690 169.700 94.950 170.020 ;
        RECT 95.210 168.400 95.350 176.160 ;
        RECT 95.670 170.440 95.810 178.460 ;
        RECT 96.070 177.520 96.330 177.840 ;
        RECT 96.130 171.040 96.270 177.520 ;
        RECT 96.070 170.720 96.330 171.040 ;
        RECT 95.670 170.300 96.270 170.440 ;
        RECT 95.610 169.700 95.870 170.020 ;
        RECT 92.390 168.000 92.650 168.320 ;
        RECT 94.750 168.260 95.350 168.400 ;
        RECT 95.670 168.320 95.810 169.700 ;
        RECT 92.450 166.870 92.590 168.000 ;
        RECT 91.990 166.730 92.590 166.870 ;
        RECT 91.990 161.860 92.130 166.730 ;
        RECT 92.510 165.765 94.390 166.135 ;
        RECT 93.770 165.280 94.030 165.600 ;
        RECT 93.830 164.920 93.970 165.280 ;
        RECT 94.750 165.000 94.890 168.260 ;
        RECT 95.610 168.000 95.870 168.320 ;
        RECT 96.130 167.720 96.270 170.300 ;
        RECT 95.150 167.320 95.410 167.640 ;
        RECT 95.670 167.580 96.270 167.720 ;
        RECT 95.210 165.600 95.350 167.320 ;
        RECT 95.150 165.280 95.410 165.600 ;
        RECT 92.390 164.600 92.650 164.920 ;
        RECT 93.770 164.600 94.030 164.920 ;
        RECT 94.750 164.860 95.350 165.000 ;
        RECT 92.450 162.880 92.590 164.600 ;
        RECT 92.390 162.560 92.650 162.880 ;
        RECT 93.830 161.860 93.970 164.600 ;
        RECT 94.230 163.920 94.490 164.240 ;
        RECT 94.290 162.880 94.430 163.920 ;
        RECT 94.230 162.560 94.490 162.880 ;
        RECT 94.290 161.860 94.430 162.560 ;
        RECT 95.210 161.860 95.350 164.860 ;
        RECT 91.930 161.540 92.190 161.860 ;
        RECT 93.770 161.540 94.030 161.860 ;
        RECT 94.230 161.540 94.490 161.860 ;
        RECT 94.690 161.540 94.950 161.860 ;
        RECT 95.150 161.540 95.410 161.860 ;
        RECT 91.930 160.860 92.190 161.180 ;
        RECT 91.470 156.440 91.730 156.760 ;
        RECT 91.990 156.330 92.130 160.860 ;
        RECT 92.510 160.325 94.390 160.695 ;
        RECT 93.770 159.840 94.030 160.160 ;
        RECT 92.390 157.120 92.650 157.440 ;
        RECT 92.450 156.840 92.590 157.120 ;
        RECT 93.310 156.840 93.570 157.100 ;
        RECT 92.450 156.780 93.570 156.840 ;
        RECT 92.450 156.700 93.510 156.780 ;
        RECT 93.830 156.760 93.970 159.840 ;
        RECT 94.750 159.480 94.890 161.540 ;
        RECT 94.690 159.160 94.950 159.480 ;
        RECT 95.670 158.800 95.810 167.580 ;
        RECT 96.590 164.320 96.730 182.620 ;
        RECT 97.450 179.900 97.710 180.220 ;
        RECT 96.990 177.180 97.250 177.500 ;
        RECT 97.050 176.140 97.190 177.180 ;
        RECT 97.510 176.140 97.650 179.900 ;
        RECT 97.970 177.840 98.110 185.680 ;
        RECT 97.910 177.520 98.170 177.840 ;
        RECT 96.990 175.820 97.250 176.140 ;
        RECT 97.450 175.820 97.710 176.140 ;
        RECT 98.430 175.800 98.570 194.180 ;
        RECT 99.350 188.720 99.490 201.660 ;
        RECT 101.190 199.600 101.330 201.660 ;
        RECT 101.650 200.280 101.790 202.680 ;
        RECT 104.350 202.340 104.610 202.660 ;
        RECT 102.970 200.640 103.230 200.960 ;
        RECT 101.590 199.960 101.850 200.280 ;
        RECT 101.130 199.280 101.390 199.600 ;
        RECT 99.750 198.940 100.010 199.260 ;
        RECT 99.810 197.900 99.950 198.940 ;
        RECT 99.750 197.580 100.010 197.900 ;
        RECT 100.670 197.240 100.930 197.560 ;
        RECT 99.750 196.900 100.010 197.220 ;
        RECT 99.810 194.500 99.950 196.900 ;
        RECT 99.750 194.180 100.010 194.500 ;
        RECT 100.210 194.180 100.470 194.500 ;
        RECT 100.270 189.400 100.410 194.180 ;
        RECT 100.730 190.080 100.870 197.240 ;
        RECT 101.130 196.900 101.390 197.220 ;
        RECT 101.190 191.780 101.330 196.900 ;
        RECT 101.650 196.540 101.790 199.960 ;
        RECT 103.030 197.220 103.170 200.640 ;
        RECT 104.410 198.240 104.550 202.340 ;
        RECT 106.650 201.660 106.910 201.980 ;
        RECT 106.710 199.940 106.850 201.660 ;
        RECT 107.510 201.125 109.390 201.495 ;
        RECT 106.650 199.620 106.910 199.940 ;
        RECT 105.270 199.280 105.530 199.600 ;
        RECT 104.350 197.920 104.610 198.240 ;
        RECT 102.970 196.900 103.230 197.220 ;
        RECT 104.350 196.900 104.610 197.220 ;
        RECT 101.590 196.220 101.850 196.540 ;
        RECT 102.510 193.500 102.770 193.820 ;
        RECT 102.570 192.800 102.710 193.500 ;
        RECT 102.510 192.480 102.770 192.800 ;
        RECT 101.130 191.460 101.390 191.780 ;
        RECT 102.050 191.460 102.310 191.780 ;
        RECT 100.670 189.760 100.930 190.080 ;
        RECT 101.190 189.740 101.330 191.460 ;
        RECT 101.130 189.480 101.390 189.740 ;
        RECT 101.130 189.420 101.790 189.480 ;
        RECT 100.210 189.080 100.470 189.400 ;
        RECT 101.190 189.340 101.790 189.420 ;
        RECT 99.290 188.400 99.550 188.720 ;
        RECT 99.750 186.360 100.010 186.680 ;
        RECT 99.810 185.660 99.950 186.360 ;
        RECT 99.290 185.340 99.550 185.660 ;
        RECT 99.750 185.340 100.010 185.660 ;
        RECT 99.350 184.640 99.490 185.340 ;
        RECT 99.290 184.320 99.550 184.640 ;
        RECT 100.270 184.300 100.410 189.080 ;
        RECT 101.130 188.060 101.390 188.380 ;
        RECT 100.210 183.980 100.470 184.300 ;
        RECT 101.190 183.280 101.330 188.060 ;
        RECT 101.650 183.960 101.790 189.340 ;
        RECT 102.110 189.060 102.250 191.460 ;
        RECT 102.510 190.780 102.770 191.100 ;
        RECT 102.050 188.740 102.310 189.060 ;
        RECT 102.570 187.360 102.710 190.780 ;
        RECT 102.510 187.040 102.770 187.360 ;
        RECT 102.050 185.340 102.310 185.660 ;
        RECT 101.590 183.640 101.850 183.960 ;
        RECT 101.130 182.960 101.390 183.280 ;
        RECT 99.750 182.620 100.010 182.940 ;
        RECT 100.670 182.620 100.930 182.940 ;
        RECT 99.810 177.500 99.950 182.620 ;
        RECT 100.210 177.860 100.470 178.180 ;
        RECT 99.750 177.180 100.010 177.500 ;
        RECT 98.370 175.480 98.630 175.800 ;
        RECT 97.900 171.545 98.180 171.915 ;
        RECT 97.970 170.360 98.110 171.545 ;
        RECT 97.910 170.040 98.170 170.360 ;
        RECT 97.450 169.020 97.710 169.340 ;
        RECT 97.510 164.920 97.650 169.020 ;
        RECT 98.430 167.720 98.570 175.480 ;
        RECT 98.830 174.460 99.090 174.780 ;
        RECT 98.890 172.400 99.030 174.460 ;
        RECT 98.830 172.080 99.090 172.400 ;
        RECT 99.810 171.040 99.950 177.180 ;
        RECT 99.750 170.720 100.010 171.040 ;
        RECT 98.830 169.020 99.090 169.340 ;
        RECT 97.970 167.640 98.570 167.720 ;
        RECT 97.910 167.580 98.570 167.640 ;
        RECT 97.910 167.320 98.170 167.580 ;
        RECT 97.450 164.600 97.710 164.920 ;
        RECT 96.590 164.180 97.650 164.320 ;
        RECT 96.070 163.580 96.330 163.900 ;
        RECT 96.990 163.580 97.250 163.900 ;
        RECT 95.610 158.480 95.870 158.800 ;
        RECT 94.690 158.140 94.950 158.460 ;
        RECT 93.770 156.440 94.030 156.760 ;
        RECT 92.390 156.330 92.650 156.420 ;
        RECT 91.990 156.190 92.650 156.330 ;
        RECT 92.390 156.100 92.650 156.190 ;
        RECT 91.930 155.420 92.190 155.740 ;
        RECT 91.990 154.720 92.130 155.420 ;
        RECT 92.510 154.885 94.390 155.255 ;
        RECT 91.930 154.400 92.190 154.720 ;
        RECT 94.750 154.380 94.890 158.140 ;
        RECT 95.610 156.780 95.870 157.100 ;
        RECT 95.150 155.420 95.410 155.740 ;
        RECT 95.210 154.380 95.350 155.420 ;
        RECT 94.690 154.060 94.950 154.380 ;
        RECT 95.150 154.060 95.410 154.380 ;
        RECT 95.670 153.610 95.810 156.780 ;
        RECT 96.130 154.040 96.270 163.580 ;
        RECT 96.530 161.200 96.790 161.520 ;
        RECT 96.590 159.480 96.730 161.200 ;
        RECT 96.530 159.160 96.790 159.480 ;
        RECT 96.530 158.315 96.790 158.460 ;
        RECT 96.520 157.945 96.800 158.315 ;
        RECT 96.530 156.780 96.790 157.100 ;
        RECT 96.590 156.420 96.730 156.780 ;
        RECT 96.530 156.100 96.790 156.420 ;
        RECT 96.070 153.720 96.330 154.040 ;
        RECT 94.750 153.470 95.810 153.610 ;
        RECT 94.230 153.040 94.490 153.360 ;
        RECT 91.470 152.700 91.730 153.020 ;
        RECT 91.010 148.280 91.270 148.600 ;
        RECT 91.530 148.000 91.670 152.700 ;
        RECT 94.290 151.320 94.430 153.040 ;
        RECT 94.230 151.000 94.490 151.320 ;
        RECT 91.930 150.660 92.190 150.980 ;
        RECT 91.990 148.850 92.130 150.660 ;
        RECT 92.510 149.445 94.390 149.815 ;
        RECT 93.310 148.960 93.570 149.280 ;
        RECT 92.390 148.850 92.650 148.940 ;
        RECT 91.990 148.710 92.650 148.850 ;
        RECT 92.390 148.620 92.650 148.710 ;
        RECT 93.370 148.600 93.510 148.960 ;
        RECT 93.310 148.280 93.570 148.600 ;
        RECT 94.230 148.280 94.490 148.600 ;
        RECT 91.530 147.860 92.130 148.000 ;
        RECT 91.470 147.260 91.730 147.580 ;
        RECT 91.010 144.540 91.270 144.860 ;
        RECT 91.070 143.840 91.210 144.540 ;
        RECT 91.010 143.520 91.270 143.840 ;
        RECT 91.010 136.380 91.270 136.700 ;
        RECT 91.070 134.660 91.210 136.380 ;
        RECT 91.010 134.340 91.270 134.660 ;
        RECT 91.010 130.940 91.270 131.260 ;
        RECT 91.070 129.900 91.210 130.940 ;
        RECT 91.010 129.580 91.270 129.900 ;
        RECT 90.550 123.800 90.810 124.120 ;
        RECT 91.530 123.780 91.670 147.260 ;
        RECT 91.990 137.120 92.130 147.860 ;
        RECT 94.290 145.200 94.430 148.280 ;
        RECT 94.750 145.880 94.890 153.470 ;
        RECT 95.150 152.700 95.410 153.020 ;
        RECT 95.610 152.700 95.870 153.020 ;
        RECT 94.690 145.560 94.950 145.880 ;
        RECT 94.230 144.880 94.490 145.200 ;
        RECT 94.690 144.540 94.950 144.860 ;
        RECT 92.510 144.005 94.390 144.375 ;
        RECT 93.770 141.820 94.030 142.140 ;
        RECT 93.830 141.120 93.970 141.820 ;
        RECT 93.770 140.800 94.030 141.120 ;
        RECT 92.510 138.565 94.390 138.935 ;
        RECT 94.750 137.720 94.890 144.540 ;
        RECT 95.210 141.120 95.350 152.700 ;
        RECT 95.670 148.000 95.810 152.700 ;
        RECT 96.070 150.320 96.330 150.640 ;
        RECT 96.130 149.280 96.270 150.320 ;
        RECT 96.070 148.960 96.330 149.280 ;
        RECT 96.070 148.510 96.330 148.600 ;
        RECT 97.050 148.510 97.190 163.580 ;
        RECT 96.070 148.370 97.190 148.510 ;
        RECT 96.070 148.280 96.330 148.370 ;
        RECT 97.510 148.260 97.650 164.180 ;
        RECT 97.910 163.920 98.170 164.240 ;
        RECT 97.970 161.860 98.110 163.920 ;
        RECT 98.430 162.540 98.570 167.580 ;
        RECT 98.890 164.920 99.030 169.020 ;
        RECT 100.270 168.320 100.410 177.860 ;
        RECT 100.210 168.000 100.470 168.320 ;
        RECT 99.290 166.980 99.550 167.300 ;
        RECT 98.830 164.600 99.090 164.920 ;
        RECT 99.350 164.320 99.490 166.980 ;
        RECT 99.750 166.300 100.010 166.620 ;
        RECT 98.890 164.240 99.490 164.320 ;
        RECT 98.830 164.180 99.490 164.240 ;
        RECT 98.830 163.920 99.090 164.180 ;
        RECT 98.370 162.220 98.630 162.540 ;
        RECT 97.910 161.540 98.170 161.860 ;
        RECT 97.970 160.160 98.110 161.540 ;
        RECT 97.910 159.840 98.170 160.160 ;
        RECT 98.890 159.480 99.030 163.920 ;
        RECT 99.810 163.810 99.950 166.300 ;
        RECT 99.350 163.670 99.950 163.810 ;
        RECT 99.350 161.860 99.490 163.670 ;
        RECT 99.290 161.540 99.550 161.860 ;
        RECT 97.910 159.390 98.170 159.480 ;
        RECT 97.910 159.250 98.570 159.390 ;
        RECT 97.910 159.160 98.170 159.250 ;
        RECT 97.910 158.480 98.170 158.800 ;
        RECT 97.970 154.630 98.110 158.480 ;
        RECT 98.430 157.440 98.570 159.250 ;
        RECT 98.830 159.160 99.090 159.480 ;
        RECT 99.750 159.160 100.010 159.480 ;
        RECT 98.370 157.120 98.630 157.440 ;
        RECT 99.290 157.120 99.550 157.440 ;
        RECT 99.350 156.420 99.490 157.120 ;
        RECT 99.810 156.955 99.950 159.160 ;
        RECT 100.210 158.820 100.470 159.140 ;
        RECT 99.740 156.585 100.020 156.955 ;
        RECT 99.290 156.100 99.550 156.420 ;
        RECT 99.750 156.330 100.010 156.420 ;
        RECT 100.270 156.330 100.410 158.820 ;
        RECT 99.750 156.190 100.410 156.330 ;
        RECT 99.750 156.100 100.010 156.190 ;
        RECT 97.970 154.490 98.570 154.630 ;
        RECT 97.910 153.720 98.170 154.040 ;
        RECT 97.970 152.000 98.110 153.720 ;
        RECT 98.430 153.700 98.570 154.490 ;
        RECT 98.370 153.380 98.630 153.700 ;
        RECT 98.370 152.700 98.630 153.020 ;
        RECT 97.910 151.680 98.170 152.000 ;
        RECT 97.910 151.000 98.170 151.320 ;
        RECT 97.970 148.940 98.110 151.000 ;
        RECT 97.910 148.620 98.170 148.940 ;
        RECT 95.670 147.860 96.270 148.000 ;
        RECT 97.450 147.940 97.710 148.260 ;
        RECT 95.610 142.500 95.870 142.820 ;
        RECT 95.150 140.800 95.410 141.120 ;
        RECT 95.670 138.400 95.810 142.500 ;
        RECT 95.610 138.080 95.870 138.400 ;
        RECT 94.690 137.400 94.950 137.720 ;
        RECT 91.990 136.980 95.810 137.120 ;
        RECT 91.930 134.680 92.190 135.000 ;
        RECT 91.990 129.470 92.130 134.680 ;
        RECT 95.150 134.000 95.410 134.320 ;
        RECT 92.510 133.125 94.390 133.495 ;
        RECT 95.210 132.960 95.350 134.000 ;
        RECT 95.150 132.640 95.410 132.960 ;
        RECT 92.390 131.620 92.650 131.940 ;
        RECT 94.230 131.620 94.490 131.940 ;
        RECT 92.450 130.240 92.590 131.620 ;
        RECT 92.390 129.920 92.650 130.240 ;
        RECT 92.390 129.470 92.650 129.560 ;
        RECT 91.990 129.330 92.650 129.470 ;
        RECT 92.390 129.240 92.650 129.330 ;
        RECT 94.290 128.960 94.430 131.620 ;
        RECT 94.290 128.880 94.890 128.960 ;
        RECT 94.230 128.820 94.890 128.880 ;
        RECT 94.230 128.560 94.490 128.820 ;
        RECT 91.930 128.220 92.190 128.540 ;
        RECT 91.990 126.840 92.130 128.220 ;
        RECT 92.510 127.685 94.390 128.055 ;
        RECT 94.750 126.840 94.890 128.820 ;
        RECT 91.930 126.520 92.190 126.840 ;
        RECT 94.690 126.520 94.950 126.840 ;
        RECT 91.470 123.460 91.730 123.780 ;
        RECT 95.670 123.440 95.810 136.980 ;
        RECT 96.130 123.780 96.270 147.860 ;
        RECT 96.990 147.260 97.250 147.580 ;
        RECT 97.910 147.260 98.170 147.580 ;
        RECT 96.530 145.220 96.790 145.540 ;
        RECT 96.590 138.060 96.730 145.220 ;
        RECT 97.050 143.840 97.190 147.260 ;
        RECT 97.450 145.220 97.710 145.540 ;
        RECT 96.990 143.520 97.250 143.840 ;
        RECT 97.510 143.160 97.650 145.220 ;
        RECT 97.450 143.070 97.710 143.160 ;
        RECT 97.050 142.930 97.710 143.070 ;
        RECT 97.050 140.100 97.190 142.930 ;
        RECT 97.450 142.840 97.710 142.930 ;
        RECT 97.450 142.160 97.710 142.480 ;
        RECT 96.990 139.780 97.250 140.100 ;
        RECT 96.530 137.740 96.790 138.060 ;
        RECT 96.530 137.060 96.790 137.380 ;
        RECT 96.590 131.940 96.730 137.060 ;
        RECT 97.510 135.000 97.650 142.160 ;
        RECT 97.450 134.680 97.710 135.000 ;
        RECT 97.510 132.960 97.650 134.680 ;
        RECT 97.450 132.640 97.710 132.960 ;
        RECT 96.530 131.620 96.790 131.940 ;
        RECT 96.590 129.560 96.730 131.620 ;
        RECT 96.530 129.240 96.790 129.560 ;
        RECT 96.070 123.460 96.330 123.780 ;
        RECT 95.610 123.120 95.870 123.440 ;
        RECT 96.530 122.780 96.790 123.100 ;
        RECT 97.450 122.780 97.710 123.100 ;
        RECT 92.510 122.245 94.390 122.615 ;
        RECT 96.590 121.740 96.730 122.780 ;
        RECT 83.650 121.420 83.910 121.740 ;
        RECT 84.110 121.420 84.370 121.740 ;
        RECT 88.710 121.420 88.970 121.740 ;
        RECT 96.530 121.420 96.790 121.740 ;
        RECT 84.170 119.020 84.310 121.420 ;
        RECT 87.330 120.060 87.590 120.380 ;
        RECT 84.110 118.700 84.370 119.020 ;
        RECT 87.390 118.680 87.530 120.060 ;
        RECT 87.330 118.360 87.590 118.680 ;
        RECT 84.110 118.020 84.370 118.340 ;
        RECT 86.870 118.250 87.130 118.340 ;
        RECT 86.010 118.110 87.130 118.250 ;
        RECT 83.650 117.340 83.910 117.660 ;
        RECT 83.710 115.960 83.850 117.340 ;
        RECT 84.170 116.040 84.310 118.020 ;
        RECT 85.030 117.340 85.290 117.660 ;
        RECT 85.090 116.300 85.230 117.340 ;
        RECT 84.170 115.960 84.770 116.040 ;
        RECT 85.030 115.980 85.290 116.300 ;
        RECT 83.650 115.640 83.910 115.960 ;
        RECT 84.170 115.900 84.830 115.960 ;
        RECT 80.890 115.300 81.150 115.620 ;
        RECT 79.970 114.620 80.230 114.940 ;
        RECT 77.510 114.085 79.390 114.455 ;
        RECT 80.950 104.355 81.090 115.300 ;
        RECT 84.170 114.940 84.310 115.900 ;
        RECT 84.570 115.640 84.830 115.900 ;
        RECT 84.110 114.620 84.370 114.940 ;
        RECT 86.010 104.355 86.150 118.110 ;
        RECT 86.870 118.020 87.130 118.110 ;
        RECT 88.770 116.640 88.910 121.420 ;
        RECT 91.010 120.400 91.270 120.720 ;
        RECT 88.710 116.320 88.970 116.640 ;
        RECT 91.070 104.355 91.210 120.400 ;
        RECT 92.510 116.805 94.390 117.175 ;
        RECT 97.510 116.640 97.650 122.780 ;
        RECT 97.970 121.740 98.110 147.260 ;
        RECT 98.430 146.560 98.570 152.700 ;
        RECT 98.830 150.890 99.090 150.980 ;
        RECT 99.350 150.890 99.490 156.100 ;
        RECT 100.270 151.320 100.410 156.190 ;
        RECT 100.730 154.380 100.870 182.620 ;
        RECT 102.110 178.180 102.250 185.340 ;
        RECT 103.030 184.300 103.170 196.900 ;
        RECT 104.410 192.800 104.550 196.900 ;
        RECT 105.330 195.520 105.470 199.280 ;
        RECT 105.730 196.220 105.990 196.540 ;
        RECT 107.110 196.220 107.370 196.540 ;
        RECT 109.870 196.220 110.130 196.540 ;
        RECT 105.790 195.520 105.930 196.220 ;
        RECT 105.270 195.200 105.530 195.520 ;
        RECT 105.730 195.200 105.990 195.520 ;
        RECT 104.350 192.480 104.610 192.800 ;
        RECT 104.350 191.460 104.610 191.780 ;
        RECT 104.410 184.640 104.550 191.460 ;
        RECT 105.330 186.340 105.470 195.200 ;
        RECT 107.170 188.720 107.310 196.220 ;
        RECT 107.510 195.685 109.390 196.055 ;
        RECT 109.930 195.180 110.070 196.220 ;
        RECT 109.870 194.860 110.130 195.180 ;
        RECT 111.710 193.500 111.970 193.820 ;
        RECT 111.770 191.780 111.910 193.500 ;
        RECT 111.710 191.460 111.970 191.780 ;
        RECT 107.510 190.245 109.390 190.615 ;
        RECT 110.330 188.740 110.590 189.060 ;
        RECT 111.250 188.740 111.510 189.060 ;
        RECT 107.110 188.400 107.370 188.720 ;
        RECT 109.870 187.040 110.130 187.360 ;
        RECT 105.270 186.020 105.530 186.340 ;
        RECT 107.510 184.805 109.390 185.175 ;
        RECT 104.350 184.320 104.610 184.640 ;
        RECT 102.970 183.980 103.230 184.300 ;
        RECT 107.110 183.980 107.370 184.300 ;
        RECT 107.170 183.620 107.310 183.980 ;
        RECT 106.190 183.300 106.450 183.620 ;
        RECT 106.650 183.300 106.910 183.620 ;
        RECT 107.110 183.300 107.370 183.620 ;
        RECT 108.950 183.475 109.210 183.620 ;
        RECT 106.250 181.920 106.390 183.300 ;
        RECT 106.710 181.920 106.850 183.300 ;
        RECT 108.940 183.105 109.220 183.475 ;
        RECT 109.010 182.940 109.150 183.105 ;
        RECT 107.110 182.620 107.370 182.940 ;
        RECT 108.490 182.795 108.750 182.940 ;
        RECT 106.190 181.600 106.450 181.920 ;
        RECT 106.650 181.600 106.910 181.920 ;
        RECT 104.350 181.435 104.610 181.580 ;
        RECT 104.340 181.065 104.620 181.435 ;
        RECT 107.170 181.240 107.310 182.620 ;
        RECT 108.480 182.425 108.760 182.795 ;
        RECT 108.950 182.620 109.210 182.940 ;
        RECT 109.010 181.240 109.150 182.620 ;
        RECT 107.110 180.920 107.370 181.240 ;
        RECT 108.950 180.920 109.210 181.240 ;
        RECT 103.430 179.900 103.690 180.220 ;
        RECT 102.050 177.860 102.310 178.180 ;
        RECT 103.490 177.500 103.630 179.900 ;
        RECT 107.510 179.365 109.390 179.735 ;
        RECT 101.130 177.180 101.390 177.500 ;
        RECT 102.050 177.180 102.310 177.500 ;
        RECT 103.430 177.180 103.690 177.500 ;
        RECT 101.190 176.140 101.330 177.180 ;
        RECT 101.130 175.820 101.390 176.140 ;
        RECT 101.590 175.480 101.850 175.800 ;
        RECT 101.130 170.040 101.390 170.360 ;
        RECT 101.190 169.340 101.330 170.040 ;
        RECT 101.130 169.020 101.390 169.340 ;
        RECT 101.190 164.920 101.330 169.020 ;
        RECT 101.130 164.600 101.390 164.920 ;
        RECT 101.190 161.860 101.330 164.600 ;
        RECT 101.130 161.540 101.390 161.860 ;
        RECT 100.670 154.060 100.930 154.380 ;
        RECT 101.190 154.040 101.330 161.540 ;
        RECT 101.650 158.800 101.790 175.480 ;
        RECT 102.110 172.740 102.250 177.180 ;
        RECT 102.970 175.140 103.230 175.460 ;
        RECT 102.510 172.760 102.770 173.080 ;
        RECT 102.050 172.420 102.310 172.740 ;
        RECT 102.050 169.700 102.310 170.020 ;
        RECT 102.110 167.640 102.250 169.700 ;
        RECT 102.050 167.320 102.310 167.640 ;
        RECT 102.570 165.600 102.710 172.760 ;
        RECT 103.030 172.060 103.170 175.140 ;
        RECT 102.970 171.740 103.230 172.060 ;
        RECT 102.970 170.040 103.230 170.360 ;
        RECT 103.030 167.640 103.170 170.040 ;
        RECT 102.970 167.320 103.230 167.640 ;
        RECT 102.970 166.640 103.230 166.960 ;
        RECT 102.510 165.280 102.770 165.600 ;
        RECT 103.030 159.480 103.170 166.640 ;
        RECT 103.490 166.620 103.630 177.180 ;
        RECT 109.930 175.800 110.070 187.040 ;
        RECT 110.390 186.340 110.530 188.740 ;
        RECT 110.790 188.060 111.050 188.380 ;
        RECT 110.330 186.020 110.590 186.340 ;
        RECT 110.390 179.200 110.530 186.020 ;
        RECT 110.330 178.880 110.590 179.200 ;
        RECT 110.850 177.840 110.990 188.060 ;
        RECT 111.310 181.920 111.450 188.740 ;
        RECT 111.770 184.300 111.910 191.460 ;
        RECT 111.710 183.980 111.970 184.300 ;
        RECT 111.250 181.600 111.510 181.920 ;
        RECT 110.790 177.520 111.050 177.840 ;
        RECT 109.870 175.480 110.130 175.800 ;
        RECT 104.350 174.460 104.610 174.780 ;
        RECT 110.790 174.460 111.050 174.780 ;
        RECT 103.430 166.300 103.690 166.620 ;
        RECT 103.430 164.940 103.690 165.260 ;
        RECT 103.490 162.880 103.630 164.940 ;
        RECT 103.430 162.560 103.690 162.880 ;
        RECT 104.410 162.200 104.550 174.460 ;
        RECT 107.510 173.925 109.390 174.295 ;
        RECT 110.330 172.080 110.590 172.400 ;
        RECT 105.270 169.700 105.530 170.020 ;
        RECT 104.350 161.880 104.610 162.200 ;
        RECT 105.330 160.160 105.470 169.700 ;
        RECT 110.390 169.340 110.530 172.080 ;
        RECT 110.850 170.020 110.990 174.460 ;
        RECT 135.630 173.380 136.780 174.600 ;
        RECT 111.250 172.420 111.510 172.740 ;
        RECT 111.710 172.420 111.970 172.740 ;
        RECT 111.310 170.360 111.450 172.420 ;
        RECT 111.770 171.915 111.910 172.420 ;
        RECT 112.160 172.225 112.440 172.595 ;
        RECT 111.700 171.545 111.980 171.915 ;
        RECT 111.250 170.040 111.510 170.360 ;
        RECT 110.790 169.700 111.050 170.020 ;
        RECT 110.330 169.020 110.590 169.340 ;
        RECT 107.510 168.485 109.390 168.855 ;
        RECT 106.650 166.640 106.910 166.960 ;
        RECT 106.190 163.580 106.450 163.900 ;
        RECT 106.250 161.520 106.390 163.580 ;
        RECT 106.190 161.200 106.450 161.520 ;
        RECT 103.430 159.840 103.690 160.160 ;
        RECT 105.270 159.840 105.530 160.160 ;
        RECT 105.730 159.840 105.990 160.160 ;
        RECT 102.970 159.160 103.230 159.480 ;
        RECT 101.590 158.480 101.850 158.800 ;
        RECT 103.490 157.100 103.630 159.840 ;
        RECT 103.890 158.820 104.150 159.140 ;
        RECT 101.580 156.585 101.860 156.955 ;
        RECT 103.430 156.780 103.690 157.100 ;
        RECT 103.950 156.760 104.090 158.820 ;
        RECT 105.270 158.140 105.530 158.460 ;
        RECT 105.330 156.760 105.470 158.140 ;
        RECT 101.650 156.420 101.790 156.585 ;
        RECT 103.890 156.440 104.150 156.760 ;
        RECT 105.270 156.440 105.530 156.760 ;
        RECT 101.590 156.100 101.850 156.420 ;
        RECT 101.130 153.720 101.390 154.040 ;
        RECT 100.210 151.000 100.470 151.320 ;
        RECT 101.190 150.980 101.330 153.720 ;
        RECT 101.650 151.660 101.790 156.100 ;
        RECT 101.590 151.340 101.850 151.660 ;
        RECT 103.950 151.320 104.090 156.440 ;
        RECT 105.790 156.420 105.930 159.840 ;
        RECT 105.730 156.100 105.990 156.420 ;
        RECT 104.350 155.420 104.610 155.740 ;
        RECT 104.410 153.020 104.550 155.420 ;
        RECT 106.190 154.400 106.450 154.720 ;
        RECT 104.350 152.700 104.610 153.020 ;
        RECT 103.890 151.000 104.150 151.320 ;
        RECT 98.830 150.750 99.490 150.890 ;
        RECT 98.830 150.660 99.090 150.750 ;
        RECT 101.130 150.660 101.390 150.980 ;
        RECT 102.050 150.720 102.310 150.980 ;
        RECT 103.950 150.720 104.090 151.000 ;
        RECT 104.410 150.980 104.550 152.700 ;
        RECT 101.650 150.660 102.310 150.720 ;
        RECT 101.650 150.580 102.250 150.660 ;
        RECT 103.490 150.580 104.090 150.720 ;
        RECT 104.350 150.660 104.610 150.980 ;
        RECT 101.650 150.300 101.790 150.580 ;
        RECT 101.590 149.980 101.850 150.300 ;
        RECT 102.050 149.980 102.310 150.300 ;
        RECT 102.110 148.940 102.250 149.980 ;
        RECT 102.050 148.620 102.310 148.940 ;
        RECT 98.370 146.240 98.630 146.560 ;
        RECT 103.490 146.220 103.630 150.580 ;
        RECT 103.890 149.980 104.150 150.300 ;
        RECT 103.950 147.580 104.090 149.980 ;
        RECT 103.890 147.260 104.150 147.580 ;
        RECT 103.430 145.900 103.690 146.220 ;
        RECT 103.950 145.540 104.090 147.260 ;
        RECT 98.830 145.220 99.090 145.540 ;
        RECT 103.890 145.220 104.150 145.540 ;
        RECT 98.370 139.100 98.630 139.420 ;
        RECT 98.430 138.400 98.570 139.100 ;
        RECT 98.370 138.080 98.630 138.400 ;
        RECT 98.890 131.940 99.030 145.220 ;
        RECT 103.430 144.540 103.690 144.860 ;
        RECT 103.490 143.840 103.630 144.540 ;
        RECT 103.430 143.520 103.690 143.840 ;
        RECT 105.730 142.500 105.990 142.820 ;
        RECT 101.130 141.820 101.390 142.140 ;
        RECT 101.190 140.440 101.330 141.820 ;
        RECT 101.130 140.120 101.390 140.440 ;
        RECT 101.190 135.000 101.330 140.120 ;
        RECT 102.050 139.780 102.310 140.100 ;
        RECT 102.110 137.630 102.250 139.780 ;
        RECT 104.350 139.440 104.610 139.760 ;
        RECT 104.410 137.720 104.550 139.440 ;
        RECT 105.790 137.720 105.930 142.500 ;
        RECT 102.510 137.630 102.770 137.720 ;
        RECT 102.110 137.490 102.770 137.630 ;
        RECT 102.510 137.400 102.770 137.490 ;
        RECT 104.350 137.400 104.610 137.720 ;
        RECT 105.730 137.630 105.990 137.720 ;
        RECT 105.330 137.490 105.990 137.630 ;
        RECT 102.570 135.680 102.710 137.400 ;
        RECT 102.510 135.360 102.770 135.680 ;
        RECT 101.130 134.680 101.390 135.000 ;
        RECT 99.290 134.340 99.550 134.660 ;
        RECT 98.830 131.620 99.090 131.940 ;
        RECT 98.370 130.940 98.630 131.260 ;
        RECT 98.430 129.220 98.570 130.940 ;
        RECT 98.890 129.220 99.030 131.620 ;
        RECT 99.350 130.240 99.490 134.340 ;
        RECT 101.190 132.620 101.330 134.680 ;
        RECT 101.130 132.300 101.390 132.620 ;
        RECT 99.290 129.920 99.550 130.240 ;
        RECT 98.370 128.900 98.630 129.220 ;
        RECT 98.830 128.900 99.090 129.220 ;
        RECT 101.190 128.880 101.330 132.300 ;
        RECT 102.570 129.560 102.710 135.360 ;
        RECT 104.350 132.300 104.610 132.620 ;
        RECT 104.410 130.240 104.550 132.300 ;
        RECT 105.330 131.260 105.470 137.490 ;
        RECT 105.730 137.400 105.990 137.490 ;
        RECT 105.730 134.000 105.990 134.320 ;
        RECT 105.270 130.940 105.530 131.260 ;
        RECT 104.350 129.920 104.610 130.240 ;
        RECT 102.510 129.240 102.770 129.560 ;
        RECT 105.330 129.220 105.470 130.940 ;
        RECT 105.790 130.240 105.930 134.000 ;
        RECT 106.250 132.180 106.390 154.400 ;
        RECT 106.710 142.820 106.850 166.640 ;
        RECT 111.310 164.920 111.450 170.040 ;
        RECT 111.770 167.300 111.910 171.545 ;
        RECT 112.230 170.700 112.370 172.225 ;
        RECT 112.170 170.380 112.430 170.700 ;
        RECT 133.750 170.070 134.880 172.730 ;
        RECT 111.710 166.980 111.970 167.300 ;
        RECT 135.630 166.640 136.740 173.380 ;
        RECT 135.630 165.420 136.780 166.640 ;
        RECT 111.250 164.600 111.510 164.920 ;
        RECT 109.870 164.260 110.130 164.580 ;
        RECT 107.510 163.045 109.390 163.415 ;
        RECT 108.030 160.860 108.290 161.180 ;
        RECT 108.090 160.160 108.230 160.860 ;
        RECT 109.930 160.160 110.070 164.260 ;
        RECT 108.030 159.840 108.290 160.160 ;
        RECT 109.870 159.840 110.130 160.160 ;
        RECT 110.330 159.160 110.590 159.480 ;
        RECT 107.510 157.605 109.390 157.975 ;
        RECT 110.390 157.440 110.530 159.160 ;
        RECT 110.330 157.120 110.590 157.440 ;
        RECT 109.870 155.420 110.130 155.740 ;
        RECT 109.930 154.040 110.070 155.420 ;
        RECT 109.870 153.720 110.130 154.040 ;
        RECT 111.250 153.720 111.510 154.040 ;
        RECT 107.510 152.165 109.390 152.535 ;
        RECT 109.870 149.980 110.130 150.300 ;
        RECT 109.930 148.600 110.070 149.980 ;
        RECT 111.310 148.600 111.450 153.720 ;
        RECT 109.870 148.280 110.130 148.600 ;
        RECT 111.250 148.280 111.510 148.600 ;
        RECT 107.510 146.725 109.390 147.095 ;
        RECT 109.410 144.540 109.670 144.860 ;
        RECT 109.470 143.160 109.610 144.540 ;
        RECT 109.410 142.840 109.670 143.160 ;
        RECT 111.310 142.820 111.450 148.280 ;
        RECT 106.650 142.500 106.910 142.820 ;
        RECT 111.250 142.500 111.510 142.820 ;
        RECT 107.510 141.285 109.390 141.655 ;
        RECT 108.030 140.120 108.290 140.440 ;
        RECT 108.090 138.400 108.230 140.120 ;
        RECT 111.310 140.100 111.450 142.500 ;
        RECT 135.630 141.200 136.780 141.270 ;
        RECT 135.630 140.180 136.800 141.200 ;
        RECT 111.250 139.780 111.510 140.100 ;
        RECT 108.030 138.080 108.290 138.400 ;
        RECT 109.870 136.380 110.130 136.700 ;
        RECT 107.510 135.845 109.390 136.215 ;
        RECT 109.930 135.000 110.070 136.380 ;
        RECT 111.310 135.000 111.450 139.780 ;
        RECT 132.560 138.140 135.160 140.060 ;
        RECT 109.870 134.680 110.130 135.000 ;
        RECT 111.250 134.680 111.510 135.000 ;
        RECT 135.640 133.320 136.800 140.180 ;
        RECT 107.570 132.180 107.830 132.280 ;
        RECT 106.250 132.040 106.850 132.180 ;
        RECT 105.730 129.920 105.990 130.240 ;
        RECT 105.270 128.900 105.530 129.220 ;
        RECT 101.130 128.560 101.390 128.880 ;
        RECT 99.750 124.140 100.010 124.460 ;
        RECT 98.830 122.780 99.090 123.100 ;
        RECT 98.890 121.740 99.030 122.780 ;
        RECT 97.910 121.420 98.170 121.740 ;
        RECT 98.830 121.420 99.090 121.740 ;
        RECT 97.910 120.740 98.170 121.060 ;
        RECT 97.970 118.680 98.110 120.740 ;
        RECT 98.370 120.060 98.630 120.380 ;
        RECT 97.910 118.360 98.170 118.680 ;
        RECT 97.450 116.320 97.710 116.640 ;
        RECT 97.970 115.620 98.110 118.360 ;
        RECT 98.430 116.300 98.570 120.060 ;
        RECT 99.810 118.680 99.950 124.140 ;
        RECT 101.190 124.120 101.330 128.560 ;
        RECT 106.710 126.840 106.850 132.040 ;
        RECT 107.170 132.040 107.830 132.180 ;
        RECT 107.170 130.240 107.310 132.040 ;
        RECT 107.570 131.960 107.830 132.040 ;
        RECT 107.510 130.405 109.390 130.775 ;
        RECT 107.110 129.920 107.370 130.240 ;
        RECT 106.190 126.520 106.450 126.840 ;
        RECT 106.650 126.520 106.910 126.840 ;
        RECT 111.710 126.520 111.970 126.840 ;
        RECT 102.970 125.840 103.230 126.160 ;
        RECT 103.030 124.120 103.170 125.840 ;
        RECT 106.250 124.800 106.390 126.520 ;
        RECT 106.650 125.500 106.910 125.820 ;
        RECT 106.190 124.480 106.450 124.800 ;
        RECT 101.130 123.800 101.390 124.120 ;
        RECT 102.970 123.800 103.230 124.120 ;
        RECT 101.190 121.400 101.330 123.800 ;
        RECT 102.050 122.780 102.310 123.100 ;
        RECT 101.130 121.080 101.390 121.400 ;
        RECT 99.750 118.360 100.010 118.680 ;
        RECT 102.110 118.000 102.250 122.780 ;
        RECT 106.250 121.480 106.390 124.480 ;
        RECT 106.710 123.440 106.850 125.500 ;
        RECT 107.510 124.965 109.390 125.335 ;
        RECT 106.650 123.120 106.910 123.440 ;
        RECT 106.250 121.340 106.850 121.480 ;
        RECT 109.870 121.420 110.130 121.740 ;
        RECT 106.190 120.740 106.450 121.060 ;
        RECT 102.050 117.680 102.310 118.000 ;
        RECT 101.130 117.340 101.390 117.660 ;
        RECT 98.370 115.980 98.630 116.300 ;
        RECT 96.070 115.300 96.330 115.620 ;
        RECT 97.910 115.300 98.170 115.620 ;
        RECT 96.130 104.355 96.270 115.300 ;
        RECT 101.190 104.355 101.330 117.340 ;
        RECT 106.250 104.355 106.390 120.740 ;
        RECT 106.710 119.360 106.850 121.340 ;
        RECT 107.510 119.525 109.390 119.895 ;
        RECT 109.930 119.360 110.070 121.420 ;
        RECT 106.650 119.040 106.910 119.360 ;
        RECT 109.870 119.040 110.130 119.360 ;
        RECT 106.710 118.340 106.850 119.040 ;
        RECT 106.650 118.020 106.910 118.340 ;
        RECT 111.770 118.195 111.910 126.520 ;
        RECT 116.310 123.120 116.570 123.440 ;
        RECT 111.700 117.825 111.980 118.195 ;
        RECT 110.790 117.340 111.050 117.660 ;
        RECT 110.850 116.300 110.990 117.340 ;
        RECT 110.790 115.980 111.050 116.300 ;
        RECT 111.710 115.300 111.970 115.620 ;
        RECT 107.510 114.085 109.390 114.455 ;
        RECT 71.290 103.660 72.810 103.800 ;
        RECT 75.820 102.355 76.100 104.355 ;
        RECT 80.880 102.355 81.160 104.355 ;
        RECT 85.940 102.355 86.220 104.355 ;
        RECT 91.000 102.355 91.280 104.355 ;
        RECT 96.060 102.355 96.340 104.355 ;
        RECT 101.120 102.355 101.400 104.355 ;
        RECT 106.180 102.355 106.460 104.355 ;
        RECT 111.240 103.800 111.520 104.355 ;
        RECT 111.770 103.800 111.910 115.300 ;
        RECT 116.370 104.355 116.510 123.120 ;
        RECT 129.750 105.580 133.160 106.650 ;
        RECT 111.240 103.660 111.910 103.800 ;
        RECT 111.240 102.355 111.520 103.660 ;
        RECT 116.300 102.355 116.580 104.355 ;
        RECT 13.920 85.550 15.140 89.420 ;
        RECT 19.910 85.980 21.130 89.850 ;
        RECT 67.730 89.640 68.670 89.840 ;
        RECT 25.730 85.120 26.950 88.990 ;
        RECT 31.780 85.510 33.000 89.380 ;
        RECT 37.750 88.780 38.970 89.290 ;
        RECT 37.680 88.620 38.970 88.780 ;
        RECT 43.810 88.630 45.030 89.530 ;
        RECT 49.740 88.640 50.960 89.040 ;
        RECT 37.680 86.810 39.070 88.620 ;
        RECT 37.750 85.420 38.970 86.810 ;
        RECT 43.810 86.720 45.140 88.630 ;
        RECT 49.740 86.920 51.010 88.640 ;
        RECT 43.810 85.660 45.030 86.720 ;
        RECT 49.740 85.170 50.960 86.920 ;
        RECT 55.530 85.320 56.750 89.190 ;
        RECT 61.720 88.640 62.940 88.870 ;
        RECT 61.720 86.600 63.130 88.640 ;
        RECT 61.720 85.000 62.940 86.600 ;
        RECT 67.580 85.770 68.800 89.640 ;
        RECT 73.850 84.290 75.070 88.160 ;
        RECT 79.730 84.310 80.950 88.180 ;
        RECT 74.090 80.440 74.370 84.290 ;
        RECT 20.140 80.160 74.370 80.440 ;
        RECT 20.140 75.650 20.420 80.160 ;
        RECT 80.070 79.800 80.350 84.310 ;
        RECT 85.470 84.100 86.690 87.970 ;
        RECT 91.460 84.500 92.680 88.320 ;
        RECT 97.600 84.630 98.820 88.240 ;
        RECT 103.650 84.740 104.870 88.610 ;
        RECT 109.620 85.420 110.840 89.290 ;
        RECT 115.740 85.700 116.960 89.570 ;
        RECT 121.520 85.700 122.740 89.570 ;
        RECT 31.380 79.520 80.350 79.800 ;
        RECT 31.380 75.850 31.660 79.520 ;
        RECT 86.050 79.170 86.330 84.100 ;
        RECT 42.510 78.890 86.330 79.170 ;
        RECT 3.960 71.320 6.050 73.240 ;
        RECT 19.330 73.120 21.890 75.650 ;
        RECT 28.185 73.180 30.255 74.460 ;
        RECT 30.670 73.320 33.230 75.850 ;
        RECT 42.510 75.750 42.790 78.890 ;
        RECT 92.030 78.570 92.310 84.500 ;
        RECT 53.830 78.290 92.310 78.570 ;
        RECT 53.830 75.820 54.110 78.290 ;
        RECT 98.010 77.990 98.290 84.630 ;
        RECT 64.900 77.710 98.290 77.990 ;
        RECT 19.005 71.800 19.865 72.640 ;
        RECT 15.560 68.610 16.990 71.210 ;
        RECT 19.305 68.570 19.845 71.800 ;
        RECT 20.145 70.600 20.555 73.120 ;
        RECT 30.205 71.810 31.065 72.650 ;
        RECT 19.325 47.770 19.825 68.570 ;
        RECT 20.165 49.090 20.555 70.600 ;
        RECT 20.955 70.010 21.845 70.740 ;
        RECT 21.055 65.190 21.315 70.010 ;
        RECT 22.695 68.620 25.405 69.470 ;
        RECT 22.895 65.840 24.825 68.620 ;
        RECT 30.505 68.580 31.045 71.810 ;
        RECT 31.345 70.610 31.755 73.320 ;
        RECT 39.475 73.150 41.545 74.430 ;
        RECT 41.910 73.220 44.470 75.750 ;
        RECT 41.425 71.780 42.285 72.620 ;
        RECT 27.795 67.130 28.915 67.810 ;
        RECT 28.075 65.850 28.745 67.130 ;
        RECT 21.455 65.460 26.505 65.840 ;
        RECT 27.865 65.440 28.915 65.850 ;
        RECT 21.055 63.640 21.435 65.190 ;
        RECT 21.175 55.800 21.435 63.640 ;
        RECT 26.485 63.200 26.755 65.240 ;
        RECT 27.615 63.200 27.885 65.200 ;
        RECT 26.485 56.510 27.885 63.200 ;
        RECT 21.085 55.290 21.445 55.800 ;
        RECT 21.065 54.860 21.445 55.290 ;
        RECT 26.485 55.190 26.755 56.510 ;
        RECT 27.615 55.150 27.885 56.510 ;
        RECT 28.885 55.260 29.205 65.190 ;
        RECT 28.885 55.200 29.215 55.260 ;
        RECT 21.065 54.580 21.315 54.860 ;
        RECT 20.865 54.180 25.505 54.580 ;
        RECT 26.405 54.290 27.535 54.300 ;
        RECT 28.895 54.290 29.215 55.200 ;
        RECT 21.065 52.060 21.315 54.180 ;
        RECT 25.765 53.490 26.125 54.110 ;
        RECT 25.845 52.610 26.105 53.490 ;
        RECT 26.385 53.240 29.215 54.290 ;
        RECT 25.675 52.230 26.205 52.610 ;
        RECT 21.065 51.970 21.565 52.060 ;
        RECT 21.055 51.240 21.565 51.970 ;
        RECT 21.295 50.240 21.565 51.240 ;
        RECT 22.205 50.990 22.475 51.940 ;
        RECT 22.205 50.840 22.675 50.990 ;
        RECT 22.205 50.160 22.765 50.840 ;
        RECT 22.285 50.150 22.765 50.160 ;
        RECT 21.575 49.620 22.195 49.980 ;
        RECT 21.615 49.090 22.045 49.620 ;
        RECT 20.165 48.670 22.045 49.090 ;
        RECT 22.535 48.960 22.765 50.150 ;
        RECT 21.615 47.800 22.045 48.670 ;
        RECT 22.455 48.360 22.835 48.960 ;
        RECT 19.325 47.060 20.015 47.770 ;
        RECT 21.435 47.440 22.055 47.800 ;
        RECT 21.135 47.060 21.425 47.250 ;
        RECT 19.325 46.620 21.425 47.060 ;
        RECT 19.325 46.600 20.015 46.620 ;
        RECT 21.135 46.380 21.425 46.620 ;
        RECT 22.055 46.990 22.325 47.240 ;
        RECT 22.535 46.990 22.765 48.360 ;
        RECT 25.355 47.010 25.685 52.030 ;
        RECT 26.405 52.020 27.535 53.240 ;
        RECT 28.895 53.220 29.215 53.240 ;
        RECT 22.055 46.880 22.765 46.990 ;
        RECT 25.345 46.960 25.685 47.010 ;
        RECT 26.235 47.780 27.615 52.020 ;
        RECT 22.055 46.570 22.715 46.880 ;
        RECT 22.055 46.400 22.325 46.570 ;
        RECT 25.345 45.000 25.625 46.960 ;
        RECT 26.235 46.920 26.535 47.780 ;
        RECT 27.315 46.920 27.615 47.780 ;
        RECT 28.165 46.920 28.495 51.990 ;
        RECT 27.565 46.380 28.045 46.760 ;
        RECT 27.665 45.760 27.915 46.380 ;
        RECT 27.565 45.160 27.945 45.760 ;
        RECT 24.825 44.230 25.925 45.000 ;
        RECT 28.215 44.930 28.495 46.920 ;
        RECT 30.525 47.780 31.025 68.580 ;
        RECT 31.365 49.100 31.755 70.610 ;
        RECT 32.155 70.020 33.045 70.750 ;
        RECT 32.255 65.200 32.515 70.020 ;
        RECT 33.895 68.630 36.605 69.480 ;
        RECT 34.095 65.850 36.025 68.630 ;
        RECT 41.725 68.550 42.265 71.780 ;
        RECT 42.565 70.580 42.975 73.220 ;
        RECT 50.055 73.090 52.125 74.370 ;
        RECT 53.150 73.290 55.710 75.820 ;
        RECT 64.900 75.810 65.180 77.710 ;
        RECT 103.990 77.230 104.270 84.740 ;
        RECT 76.140 76.950 104.270 77.230 ;
        RECT 52.675 71.760 53.535 72.600 ;
        RECT 38.995 67.140 40.115 67.820 ;
        RECT 39.275 65.860 39.945 67.140 ;
        RECT 32.655 65.470 37.705 65.850 ;
        RECT 39.065 65.450 40.115 65.860 ;
        RECT 32.255 63.650 32.635 65.200 ;
        RECT 32.375 55.810 32.635 63.650 ;
        RECT 37.685 63.210 37.955 65.250 ;
        RECT 38.815 63.210 39.085 65.210 ;
        RECT 37.685 56.520 39.085 63.210 ;
        RECT 32.285 55.300 32.645 55.810 ;
        RECT 32.265 54.870 32.645 55.300 ;
        RECT 37.685 55.200 37.955 56.520 ;
        RECT 38.815 55.160 39.085 56.520 ;
        RECT 40.085 55.270 40.405 65.200 ;
        RECT 40.085 55.210 40.415 55.270 ;
        RECT 32.265 54.590 32.515 54.870 ;
        RECT 32.065 54.190 36.705 54.590 ;
        RECT 37.605 54.300 38.735 54.310 ;
        RECT 40.095 54.300 40.415 55.210 ;
        RECT 32.265 52.070 32.515 54.190 ;
        RECT 36.965 53.500 37.325 54.120 ;
        RECT 37.045 52.620 37.305 53.500 ;
        RECT 37.585 53.250 40.415 54.300 ;
        RECT 36.875 52.240 37.405 52.620 ;
        RECT 32.265 51.980 32.765 52.070 ;
        RECT 32.255 51.250 32.765 51.980 ;
        RECT 32.495 50.250 32.765 51.250 ;
        RECT 33.405 51.000 33.675 51.950 ;
        RECT 33.405 50.850 33.875 51.000 ;
        RECT 33.405 50.170 33.965 50.850 ;
        RECT 33.485 50.160 33.965 50.170 ;
        RECT 32.775 49.630 33.395 49.990 ;
        RECT 32.815 49.100 33.245 49.630 ;
        RECT 31.365 48.680 33.245 49.100 ;
        RECT 33.735 48.970 33.965 50.160 ;
        RECT 32.815 47.810 33.245 48.680 ;
        RECT 33.655 48.370 34.035 48.970 ;
        RECT 30.525 47.070 31.215 47.780 ;
        RECT 32.635 47.450 33.255 47.810 ;
        RECT 32.335 47.070 32.625 47.260 ;
        RECT 30.525 46.630 32.625 47.070 ;
        RECT 30.525 46.610 31.215 46.630 ;
        RECT 32.335 46.390 32.625 46.630 ;
        RECT 33.255 47.000 33.525 47.250 ;
        RECT 33.735 47.000 33.965 48.370 ;
        RECT 36.555 47.020 36.885 52.040 ;
        RECT 37.605 52.030 38.735 53.250 ;
        RECT 40.095 53.230 40.415 53.250 ;
        RECT 33.255 46.890 33.965 47.000 ;
        RECT 36.545 46.970 36.885 47.020 ;
        RECT 37.435 47.790 38.815 52.030 ;
        RECT 33.255 46.580 33.915 46.890 ;
        RECT 33.255 46.410 33.525 46.580 ;
        RECT 36.545 45.010 36.825 46.970 ;
        RECT 37.435 46.930 37.735 47.790 ;
        RECT 38.515 46.930 38.815 47.790 ;
        RECT 39.365 46.930 39.695 52.000 ;
        RECT 38.765 46.390 39.245 46.770 ;
        RECT 38.865 45.770 39.115 46.390 ;
        RECT 38.765 45.170 39.145 45.770 ;
        RECT 28.215 43.200 28.515 44.930 ;
        RECT 36.025 44.240 37.125 45.010 ;
        RECT 39.415 44.940 39.695 46.930 ;
        RECT 41.745 47.750 42.245 68.550 ;
        RECT 42.585 49.070 42.975 70.580 ;
        RECT 43.375 69.990 44.265 70.720 ;
        RECT 43.475 65.170 43.735 69.990 ;
        RECT 45.115 68.600 47.825 69.450 ;
        RECT 45.315 65.820 47.245 68.600 ;
        RECT 52.975 68.530 53.515 71.760 ;
        RECT 53.815 70.560 54.225 73.290 ;
        RECT 61.475 73.120 63.545 74.400 ;
        RECT 64.400 73.280 66.960 75.810 ;
        RECT 76.140 75.740 76.420 76.950 ;
        RECT 109.970 76.610 110.250 85.420 ;
        RECT 87.580 76.330 110.250 76.610 ;
        RECT 87.580 75.760 87.860 76.330 ;
        RECT 115.950 76.030 116.230 85.700 ;
        RECT 98.850 75.840 116.230 76.030 ;
        RECT 63.895 71.750 64.755 72.590 ;
        RECT 50.215 67.110 51.335 67.790 ;
        RECT 50.495 65.830 51.165 67.110 ;
        RECT 43.875 65.440 48.925 65.820 ;
        RECT 50.285 65.420 51.335 65.830 ;
        RECT 43.475 63.620 43.855 65.170 ;
        RECT 43.595 55.780 43.855 63.620 ;
        RECT 48.905 63.180 49.175 65.220 ;
        RECT 50.035 63.180 50.305 65.180 ;
        RECT 48.905 56.490 50.305 63.180 ;
        RECT 43.505 55.270 43.865 55.780 ;
        RECT 43.485 54.840 43.865 55.270 ;
        RECT 48.905 55.170 49.175 56.490 ;
        RECT 50.035 55.130 50.305 56.490 ;
        RECT 51.305 55.240 51.625 65.170 ;
        RECT 51.305 55.180 51.635 55.240 ;
        RECT 43.485 54.560 43.735 54.840 ;
        RECT 43.285 54.160 47.925 54.560 ;
        RECT 48.825 54.270 49.955 54.280 ;
        RECT 51.315 54.270 51.635 55.180 ;
        RECT 43.485 52.040 43.735 54.160 ;
        RECT 48.185 53.470 48.545 54.090 ;
        RECT 48.265 52.590 48.525 53.470 ;
        RECT 48.805 53.220 51.635 54.270 ;
        RECT 48.095 52.210 48.625 52.590 ;
        RECT 43.485 51.950 43.985 52.040 ;
        RECT 43.475 51.220 43.985 51.950 ;
        RECT 43.715 50.220 43.985 51.220 ;
        RECT 44.625 50.970 44.895 51.920 ;
        RECT 44.625 50.820 45.095 50.970 ;
        RECT 44.625 50.140 45.185 50.820 ;
        RECT 44.705 50.130 45.185 50.140 ;
        RECT 43.995 49.600 44.615 49.960 ;
        RECT 44.035 49.070 44.465 49.600 ;
        RECT 42.585 48.650 44.465 49.070 ;
        RECT 44.955 48.940 45.185 50.130 ;
        RECT 44.035 47.780 44.465 48.650 ;
        RECT 44.875 48.340 45.255 48.940 ;
        RECT 41.745 47.040 42.435 47.750 ;
        RECT 43.855 47.420 44.475 47.780 ;
        RECT 43.555 47.040 43.845 47.230 ;
        RECT 41.745 46.600 43.845 47.040 ;
        RECT 41.745 46.580 42.435 46.600 ;
        RECT 43.555 46.360 43.845 46.600 ;
        RECT 44.475 46.970 44.745 47.220 ;
        RECT 44.955 46.970 45.185 48.340 ;
        RECT 47.775 46.990 48.105 52.010 ;
        RECT 48.825 52.000 49.955 53.220 ;
        RECT 51.315 53.200 51.635 53.220 ;
        RECT 44.475 46.860 45.185 46.970 ;
        RECT 47.765 46.940 48.105 46.990 ;
        RECT 48.655 47.760 50.035 52.000 ;
        RECT 44.475 46.550 45.135 46.860 ;
        RECT 44.475 46.380 44.745 46.550 ;
        RECT 47.765 44.980 48.045 46.940 ;
        RECT 48.655 46.900 48.955 47.760 ;
        RECT 49.735 46.900 50.035 47.760 ;
        RECT 50.585 46.900 50.915 51.970 ;
        RECT 49.985 46.360 50.465 46.740 ;
        RECT 50.085 45.740 50.335 46.360 ;
        RECT 49.985 45.140 50.365 45.740 ;
        RECT 39.415 43.210 39.715 44.940 ;
        RECT 47.245 44.210 48.345 44.980 ;
        RECT 50.635 44.910 50.915 46.900 ;
        RECT 52.995 47.730 53.495 68.530 ;
        RECT 53.835 49.050 54.225 70.560 ;
        RECT 54.625 69.970 55.515 70.700 ;
        RECT 54.725 65.150 54.985 69.970 ;
        RECT 56.365 68.580 59.075 69.430 ;
        RECT 56.565 65.800 58.495 68.580 ;
        RECT 64.195 68.520 64.735 71.750 ;
        RECT 65.035 70.550 65.445 73.280 ;
        RECT 72.585 73.130 74.655 74.410 ;
        RECT 75.550 73.210 78.110 75.740 ;
        RECT 75.135 71.740 75.995 72.580 ;
        RECT 61.465 67.090 62.585 67.770 ;
        RECT 61.745 65.810 62.415 67.090 ;
        RECT 55.125 65.420 60.175 65.800 ;
        RECT 61.535 65.400 62.585 65.810 ;
        RECT 54.725 63.600 55.105 65.150 ;
        RECT 54.845 55.760 55.105 63.600 ;
        RECT 60.155 63.160 60.425 65.200 ;
        RECT 61.285 63.160 61.555 65.160 ;
        RECT 60.155 56.470 61.555 63.160 ;
        RECT 54.755 55.250 55.115 55.760 ;
        RECT 54.735 54.820 55.115 55.250 ;
        RECT 60.155 55.150 60.425 56.470 ;
        RECT 61.285 55.110 61.555 56.470 ;
        RECT 62.555 55.220 62.875 65.150 ;
        RECT 62.555 55.160 62.885 55.220 ;
        RECT 54.735 54.540 54.985 54.820 ;
        RECT 54.535 54.140 59.175 54.540 ;
        RECT 60.075 54.250 61.205 54.260 ;
        RECT 62.565 54.250 62.885 55.160 ;
        RECT 54.735 52.020 54.985 54.140 ;
        RECT 59.435 53.450 59.795 54.070 ;
        RECT 59.515 52.570 59.775 53.450 ;
        RECT 60.055 53.200 62.885 54.250 ;
        RECT 59.345 52.190 59.875 52.570 ;
        RECT 54.735 51.930 55.235 52.020 ;
        RECT 54.725 51.200 55.235 51.930 ;
        RECT 54.965 50.200 55.235 51.200 ;
        RECT 55.875 50.950 56.145 51.900 ;
        RECT 55.875 50.800 56.345 50.950 ;
        RECT 55.875 50.120 56.435 50.800 ;
        RECT 55.955 50.110 56.435 50.120 ;
        RECT 55.245 49.580 55.865 49.940 ;
        RECT 55.285 49.050 55.715 49.580 ;
        RECT 53.835 48.630 55.715 49.050 ;
        RECT 56.205 48.920 56.435 50.110 ;
        RECT 55.285 47.760 55.715 48.630 ;
        RECT 56.125 48.320 56.505 48.920 ;
        RECT 52.995 47.020 53.685 47.730 ;
        RECT 55.105 47.400 55.725 47.760 ;
        RECT 54.805 47.020 55.095 47.210 ;
        RECT 52.995 46.580 55.095 47.020 ;
        RECT 52.995 46.560 53.685 46.580 ;
        RECT 54.805 46.340 55.095 46.580 ;
        RECT 55.725 46.950 55.995 47.200 ;
        RECT 56.205 46.950 56.435 48.320 ;
        RECT 59.025 46.970 59.355 51.990 ;
        RECT 60.075 51.980 61.205 53.200 ;
        RECT 62.565 53.180 62.885 53.200 ;
        RECT 55.725 46.840 56.435 46.950 ;
        RECT 59.015 46.920 59.355 46.970 ;
        RECT 59.905 47.740 61.285 51.980 ;
        RECT 55.725 46.530 56.385 46.840 ;
        RECT 55.725 46.360 55.995 46.530 ;
        RECT 59.015 44.960 59.295 46.920 ;
        RECT 59.905 46.880 60.205 47.740 ;
        RECT 60.985 46.880 61.285 47.740 ;
        RECT 61.835 46.880 62.165 51.950 ;
        RECT 61.235 46.340 61.715 46.720 ;
        RECT 61.335 45.720 61.585 46.340 ;
        RECT 61.235 45.120 61.615 45.720 ;
        RECT 19.865 42.210 21.245 42.780 ;
        RECT 27.495 42.630 28.875 43.200 ;
        RECT 31.145 42.210 32.525 42.780 ;
        RECT 38.695 42.640 40.075 43.210 ;
        RECT 50.635 43.180 50.935 44.910 ;
        RECT 58.495 44.190 59.595 44.960 ;
        RECT 61.885 44.890 62.165 46.880 ;
        RECT 64.215 47.720 64.715 68.520 ;
        RECT 65.055 49.040 65.445 70.550 ;
        RECT 65.845 69.960 66.735 70.690 ;
        RECT 65.945 65.140 66.205 69.960 ;
        RECT 67.585 68.570 70.295 69.420 ;
        RECT 67.785 65.790 69.715 68.570 ;
        RECT 75.435 68.510 75.975 71.740 ;
        RECT 76.275 70.540 76.685 73.210 ;
        RECT 83.855 73.120 85.925 74.400 ;
        RECT 86.850 73.230 89.410 75.760 ;
        RECT 98.150 75.750 116.230 75.840 ;
        RECT 86.385 71.750 87.245 72.590 ;
        RECT 72.685 67.080 73.805 67.760 ;
        RECT 72.965 65.800 73.635 67.080 ;
        RECT 66.345 65.410 71.395 65.790 ;
        RECT 72.755 65.390 73.805 65.800 ;
        RECT 65.945 63.590 66.325 65.140 ;
        RECT 66.065 55.750 66.325 63.590 ;
        RECT 71.375 63.150 71.645 65.190 ;
        RECT 72.505 63.150 72.775 65.150 ;
        RECT 71.375 56.460 72.775 63.150 ;
        RECT 65.975 55.240 66.335 55.750 ;
        RECT 65.955 54.810 66.335 55.240 ;
        RECT 71.375 55.140 71.645 56.460 ;
        RECT 72.505 55.100 72.775 56.460 ;
        RECT 73.775 55.210 74.095 65.140 ;
        RECT 73.775 55.150 74.105 55.210 ;
        RECT 65.955 54.530 66.205 54.810 ;
        RECT 65.755 54.130 70.395 54.530 ;
        RECT 71.295 54.240 72.425 54.250 ;
        RECT 73.785 54.240 74.105 55.150 ;
        RECT 65.955 52.010 66.205 54.130 ;
        RECT 70.655 53.440 71.015 54.060 ;
        RECT 70.735 52.560 70.995 53.440 ;
        RECT 71.275 53.190 74.105 54.240 ;
        RECT 70.565 52.180 71.095 52.560 ;
        RECT 65.955 51.920 66.455 52.010 ;
        RECT 65.945 51.190 66.455 51.920 ;
        RECT 66.185 50.190 66.455 51.190 ;
        RECT 67.095 50.940 67.365 51.890 ;
        RECT 67.095 50.790 67.565 50.940 ;
        RECT 67.095 50.110 67.655 50.790 ;
        RECT 67.175 50.100 67.655 50.110 ;
        RECT 66.465 49.570 67.085 49.930 ;
        RECT 66.505 49.040 66.935 49.570 ;
        RECT 65.055 48.620 66.935 49.040 ;
        RECT 67.425 48.910 67.655 50.100 ;
        RECT 66.505 47.750 66.935 48.620 ;
        RECT 67.345 48.310 67.725 48.910 ;
        RECT 64.215 47.010 64.905 47.720 ;
        RECT 66.325 47.390 66.945 47.750 ;
        RECT 66.025 47.010 66.315 47.200 ;
        RECT 64.215 46.570 66.315 47.010 ;
        RECT 64.215 46.550 64.905 46.570 ;
        RECT 66.025 46.330 66.315 46.570 ;
        RECT 66.945 46.940 67.215 47.190 ;
        RECT 67.425 46.940 67.655 48.310 ;
        RECT 70.245 46.960 70.575 51.980 ;
        RECT 71.295 51.970 72.425 53.190 ;
        RECT 73.785 53.170 74.105 53.190 ;
        RECT 66.945 46.830 67.655 46.940 ;
        RECT 70.235 46.910 70.575 46.960 ;
        RECT 71.125 47.730 72.505 51.970 ;
        RECT 66.945 46.520 67.605 46.830 ;
        RECT 66.945 46.350 67.215 46.520 ;
        RECT 70.235 44.950 70.515 46.910 ;
        RECT 71.125 46.870 71.425 47.730 ;
        RECT 72.205 46.870 72.505 47.730 ;
        RECT 73.055 46.870 73.385 51.940 ;
        RECT 72.455 46.330 72.935 46.710 ;
        RECT 72.555 45.710 72.805 46.330 ;
        RECT 72.455 45.110 72.835 45.710 ;
        RECT 20.225 40.480 20.525 42.210 ;
        RECT 20.245 38.490 20.525 40.480 ;
        RECT 22.815 40.410 23.915 41.180 ;
        RECT 31.505 40.480 31.805 42.210 ;
        RECT 42.435 42.190 43.815 42.760 ;
        RECT 49.915 42.610 51.295 43.180 ;
        RECT 61.885 43.160 62.185 44.890 ;
        RECT 69.715 44.180 70.815 44.950 ;
        RECT 73.105 44.880 73.385 46.870 ;
        RECT 75.455 47.710 75.955 68.510 ;
        RECT 76.295 49.030 76.685 70.540 ;
        RECT 77.085 69.950 77.975 70.680 ;
        RECT 77.185 65.130 77.445 69.950 ;
        RECT 78.825 68.560 81.535 69.410 ;
        RECT 79.025 65.780 80.955 68.560 ;
        RECT 86.685 68.520 87.225 71.750 ;
        RECT 87.525 70.550 87.935 73.230 ;
        RECT 95.045 73.060 97.115 74.340 ;
        RECT 98.150 73.310 100.710 75.750 ;
        RECT 109.390 75.480 111.950 75.560 ;
        RECT 121.930 75.480 122.210 85.700 ;
        RECT 127.550 85.510 128.770 89.380 ;
        RECT 127.910 76.040 128.190 85.510 ;
        RECT 133.380 76.580 136.010 77.880 ;
        RECT 137.240 76.560 139.870 77.860 ;
        RECT 109.390 75.200 122.210 75.480 ;
        RECT 97.665 71.740 98.525 72.580 ;
        RECT 83.925 67.070 85.045 67.750 ;
        RECT 84.205 65.790 84.875 67.070 ;
        RECT 77.585 65.400 82.635 65.780 ;
        RECT 83.995 65.380 85.045 65.790 ;
        RECT 77.185 63.580 77.565 65.130 ;
        RECT 77.305 55.740 77.565 63.580 ;
        RECT 82.615 63.140 82.885 65.180 ;
        RECT 83.745 63.140 84.015 65.140 ;
        RECT 82.615 56.450 84.015 63.140 ;
        RECT 77.215 55.230 77.575 55.740 ;
        RECT 77.195 54.800 77.575 55.230 ;
        RECT 82.615 55.130 82.885 56.450 ;
        RECT 83.745 55.090 84.015 56.450 ;
        RECT 85.015 55.200 85.335 65.130 ;
        RECT 85.015 55.140 85.345 55.200 ;
        RECT 77.195 54.520 77.445 54.800 ;
        RECT 76.995 54.120 81.635 54.520 ;
        RECT 82.535 54.230 83.665 54.240 ;
        RECT 85.025 54.230 85.345 55.140 ;
        RECT 77.195 52.000 77.445 54.120 ;
        RECT 81.895 53.430 82.255 54.050 ;
        RECT 81.975 52.550 82.235 53.430 ;
        RECT 82.515 53.180 85.345 54.230 ;
        RECT 81.805 52.170 82.335 52.550 ;
        RECT 77.195 51.910 77.695 52.000 ;
        RECT 77.185 51.180 77.695 51.910 ;
        RECT 77.425 50.180 77.695 51.180 ;
        RECT 78.335 50.930 78.605 51.880 ;
        RECT 78.335 50.780 78.805 50.930 ;
        RECT 78.335 50.100 78.895 50.780 ;
        RECT 78.415 50.090 78.895 50.100 ;
        RECT 77.705 49.560 78.325 49.920 ;
        RECT 77.745 49.030 78.175 49.560 ;
        RECT 76.295 48.610 78.175 49.030 ;
        RECT 78.665 48.900 78.895 50.090 ;
        RECT 77.745 47.740 78.175 48.610 ;
        RECT 78.585 48.300 78.965 48.900 ;
        RECT 75.455 47.000 76.145 47.710 ;
        RECT 77.565 47.380 78.185 47.740 ;
        RECT 77.265 47.000 77.555 47.190 ;
        RECT 75.455 46.560 77.555 47.000 ;
        RECT 75.455 46.540 76.145 46.560 ;
        RECT 77.265 46.320 77.555 46.560 ;
        RECT 78.185 46.930 78.455 47.180 ;
        RECT 78.665 46.930 78.895 48.300 ;
        RECT 81.485 46.950 81.815 51.970 ;
        RECT 82.535 51.960 83.665 53.180 ;
        RECT 85.025 53.160 85.345 53.180 ;
        RECT 78.185 46.820 78.895 46.930 ;
        RECT 81.475 46.900 81.815 46.950 ;
        RECT 82.365 47.720 83.745 51.960 ;
        RECT 78.185 46.510 78.845 46.820 ;
        RECT 78.185 46.340 78.455 46.510 ;
        RECT 81.475 44.940 81.755 46.900 ;
        RECT 82.365 46.860 82.665 47.720 ;
        RECT 83.445 46.860 83.745 47.720 ;
        RECT 84.295 46.860 84.625 51.930 ;
        RECT 83.695 46.320 84.175 46.700 ;
        RECT 83.795 45.700 84.045 46.320 ;
        RECT 83.695 45.100 84.075 45.700 ;
        RECT 53.655 42.190 55.035 42.760 ;
        RECT 61.165 42.590 62.545 43.160 ;
        RECT 73.105 43.150 73.405 44.880 ;
        RECT 80.955 44.170 82.055 44.940 ;
        RECT 84.345 44.870 84.625 46.860 ;
        RECT 86.705 47.720 87.205 68.520 ;
        RECT 87.545 49.040 87.935 70.550 ;
        RECT 88.335 69.960 89.225 70.690 ;
        RECT 88.435 65.140 88.695 69.960 ;
        RECT 90.075 68.570 92.785 69.420 ;
        RECT 90.275 65.790 92.205 68.570 ;
        RECT 97.965 68.510 98.505 71.740 ;
        RECT 98.805 70.540 99.215 73.310 ;
        RECT 106.455 73.110 108.525 74.390 ;
        RECT 109.390 73.030 111.950 75.200 ;
        RECT 125.760 74.810 128.190 76.040 ;
        RECT 121.290 74.790 128.190 74.810 ;
        RECT 120.600 74.530 128.190 74.790 ;
        RECT 117.655 73.110 119.725 74.390 ;
        RECT 120.600 73.180 128.160 74.530 ;
        RECT 129.505 73.190 131.575 74.470 ;
        RECT 120.600 73.110 126.160 73.180 ;
        RECT 108.935 71.740 109.795 72.580 ;
        RECT 95.175 67.080 96.295 67.760 ;
        RECT 95.455 65.800 96.125 67.080 ;
        RECT 88.835 65.410 93.885 65.790 ;
        RECT 95.245 65.390 96.295 65.800 ;
        RECT 88.435 63.590 88.815 65.140 ;
        RECT 88.555 55.750 88.815 63.590 ;
        RECT 93.865 63.150 94.135 65.190 ;
        RECT 94.995 63.150 95.265 65.150 ;
        RECT 93.865 56.460 95.265 63.150 ;
        RECT 88.465 55.240 88.825 55.750 ;
        RECT 88.445 54.810 88.825 55.240 ;
        RECT 93.865 55.140 94.135 56.460 ;
        RECT 94.995 55.100 95.265 56.460 ;
        RECT 96.265 55.210 96.585 65.140 ;
        RECT 96.265 55.150 96.595 55.210 ;
        RECT 88.445 54.530 88.695 54.810 ;
        RECT 88.245 54.130 92.885 54.530 ;
        RECT 93.785 54.240 94.915 54.250 ;
        RECT 96.275 54.240 96.595 55.150 ;
        RECT 88.445 52.010 88.695 54.130 ;
        RECT 93.145 53.440 93.505 54.060 ;
        RECT 93.225 52.560 93.485 53.440 ;
        RECT 93.765 53.190 96.595 54.240 ;
        RECT 93.055 52.180 93.585 52.560 ;
        RECT 88.445 51.920 88.945 52.010 ;
        RECT 88.435 51.190 88.945 51.920 ;
        RECT 88.675 50.190 88.945 51.190 ;
        RECT 89.585 50.940 89.855 51.890 ;
        RECT 89.585 50.790 90.055 50.940 ;
        RECT 89.585 50.110 90.145 50.790 ;
        RECT 89.665 50.100 90.145 50.110 ;
        RECT 88.955 49.570 89.575 49.930 ;
        RECT 88.995 49.040 89.425 49.570 ;
        RECT 87.545 48.620 89.425 49.040 ;
        RECT 89.915 48.910 90.145 50.100 ;
        RECT 88.995 47.750 89.425 48.620 ;
        RECT 89.835 48.310 90.215 48.910 ;
        RECT 86.705 47.010 87.395 47.720 ;
        RECT 88.815 47.390 89.435 47.750 ;
        RECT 88.515 47.010 88.805 47.200 ;
        RECT 86.705 46.570 88.805 47.010 ;
        RECT 86.705 46.550 87.395 46.570 ;
        RECT 88.515 46.330 88.805 46.570 ;
        RECT 89.435 46.940 89.705 47.190 ;
        RECT 89.915 46.940 90.145 48.310 ;
        RECT 92.735 46.960 93.065 51.980 ;
        RECT 93.785 51.970 94.915 53.190 ;
        RECT 96.275 53.170 96.595 53.190 ;
        RECT 89.435 46.830 90.145 46.940 ;
        RECT 92.725 46.910 93.065 46.960 ;
        RECT 93.615 47.730 94.995 51.970 ;
        RECT 89.435 46.520 90.095 46.830 ;
        RECT 89.435 46.350 89.705 46.520 ;
        RECT 92.725 44.950 93.005 46.910 ;
        RECT 93.615 46.870 93.915 47.730 ;
        RECT 94.695 46.870 94.995 47.730 ;
        RECT 95.545 46.870 95.875 51.940 ;
        RECT 94.945 46.330 95.425 46.710 ;
        RECT 95.045 45.710 95.295 46.330 ;
        RECT 94.945 45.110 95.325 45.710 ;
        RECT 64.855 42.190 66.235 42.760 ;
        RECT 72.385 42.580 73.765 43.150 ;
        RECT 84.345 43.140 84.645 44.870 ;
        RECT 92.205 44.180 93.305 44.950 ;
        RECT 95.595 44.880 95.875 46.870 ;
        RECT 97.985 47.710 98.485 68.510 ;
        RECT 98.825 49.030 99.215 70.540 ;
        RECT 99.615 69.950 100.505 70.680 ;
        RECT 99.715 65.130 99.975 69.950 ;
        RECT 101.355 68.560 104.065 69.410 ;
        RECT 101.555 65.780 103.485 68.560 ;
        RECT 109.235 68.510 109.775 71.740 ;
        RECT 110.075 70.540 110.485 73.030 ;
        RECT 120.185 71.740 121.045 72.580 ;
        RECT 106.455 67.070 107.575 67.750 ;
        RECT 106.735 65.790 107.405 67.070 ;
        RECT 100.115 65.400 105.165 65.780 ;
        RECT 106.525 65.380 107.575 65.790 ;
        RECT 99.715 63.580 100.095 65.130 ;
        RECT 99.835 55.740 100.095 63.580 ;
        RECT 105.145 63.140 105.415 65.180 ;
        RECT 106.275 63.140 106.545 65.140 ;
        RECT 105.145 56.450 106.545 63.140 ;
        RECT 99.745 55.230 100.105 55.740 ;
        RECT 99.725 54.800 100.105 55.230 ;
        RECT 105.145 55.130 105.415 56.450 ;
        RECT 106.275 55.090 106.545 56.450 ;
        RECT 107.545 55.200 107.865 65.130 ;
        RECT 107.545 55.140 107.875 55.200 ;
        RECT 99.725 54.520 99.975 54.800 ;
        RECT 99.525 54.120 104.165 54.520 ;
        RECT 105.065 54.230 106.195 54.240 ;
        RECT 107.555 54.230 107.875 55.140 ;
        RECT 99.725 52.000 99.975 54.120 ;
        RECT 104.425 53.430 104.785 54.050 ;
        RECT 104.505 52.550 104.765 53.430 ;
        RECT 105.045 53.180 107.875 54.230 ;
        RECT 104.335 52.170 104.865 52.550 ;
        RECT 99.725 51.910 100.225 52.000 ;
        RECT 99.715 51.180 100.225 51.910 ;
        RECT 99.955 50.180 100.225 51.180 ;
        RECT 100.865 50.930 101.135 51.880 ;
        RECT 100.865 50.780 101.335 50.930 ;
        RECT 100.865 50.100 101.425 50.780 ;
        RECT 100.945 50.090 101.425 50.100 ;
        RECT 100.235 49.560 100.855 49.920 ;
        RECT 100.275 49.030 100.705 49.560 ;
        RECT 98.825 48.610 100.705 49.030 ;
        RECT 101.195 48.900 101.425 50.090 ;
        RECT 100.275 47.740 100.705 48.610 ;
        RECT 101.115 48.300 101.495 48.900 ;
        RECT 97.985 47.000 98.675 47.710 ;
        RECT 100.095 47.380 100.715 47.740 ;
        RECT 99.795 47.000 100.085 47.190 ;
        RECT 97.985 46.560 100.085 47.000 ;
        RECT 97.985 46.540 98.675 46.560 ;
        RECT 99.795 46.320 100.085 46.560 ;
        RECT 100.715 46.930 100.985 47.180 ;
        RECT 101.195 46.930 101.425 48.300 ;
        RECT 104.015 46.950 104.345 51.970 ;
        RECT 105.065 51.960 106.195 53.180 ;
        RECT 107.555 53.160 107.875 53.180 ;
        RECT 100.715 46.820 101.425 46.930 ;
        RECT 104.005 46.900 104.345 46.950 ;
        RECT 104.895 47.720 106.275 51.960 ;
        RECT 100.715 46.510 101.375 46.820 ;
        RECT 100.715 46.340 100.985 46.510 ;
        RECT 104.005 44.940 104.285 46.900 ;
        RECT 104.895 46.860 105.195 47.720 ;
        RECT 105.975 46.860 106.275 47.720 ;
        RECT 106.825 46.860 107.155 51.930 ;
        RECT 106.225 46.320 106.705 46.700 ;
        RECT 106.325 45.700 106.575 46.320 ;
        RECT 106.225 45.100 106.605 45.700 ;
        RECT 95.595 43.150 95.895 44.880 ;
        RECT 103.485 44.170 104.585 44.940 ;
        RECT 106.875 44.870 107.155 46.860 ;
        RECT 109.255 47.710 109.755 68.510 ;
        RECT 110.095 49.030 110.485 70.540 ;
        RECT 110.885 69.950 111.775 70.680 ;
        RECT 110.985 65.130 111.245 69.950 ;
        RECT 112.625 68.560 115.335 69.410 ;
        RECT 112.825 65.780 114.755 68.560 ;
        RECT 120.485 68.510 121.025 71.740 ;
        RECT 121.325 70.540 121.735 73.110 ;
        RECT 132.925 70.810 133.225 70.900 ;
        RECT 117.725 67.070 118.845 67.750 ;
        RECT 118.005 65.790 118.675 67.070 ;
        RECT 111.385 65.400 116.435 65.780 ;
        RECT 117.795 65.380 118.845 65.790 ;
        RECT 110.985 63.580 111.365 65.130 ;
        RECT 111.105 55.740 111.365 63.580 ;
        RECT 116.415 63.140 116.685 65.180 ;
        RECT 117.545 63.140 117.815 65.140 ;
        RECT 116.415 56.450 117.815 63.140 ;
        RECT 111.015 55.230 111.375 55.740 ;
        RECT 110.995 54.800 111.375 55.230 ;
        RECT 116.415 55.130 116.685 56.450 ;
        RECT 117.545 55.090 117.815 56.450 ;
        RECT 118.815 55.200 119.135 65.130 ;
        RECT 118.815 55.140 119.145 55.200 ;
        RECT 110.995 54.520 111.245 54.800 ;
        RECT 110.795 54.120 115.435 54.520 ;
        RECT 116.335 54.230 117.465 54.240 ;
        RECT 118.825 54.230 119.145 55.140 ;
        RECT 110.995 52.000 111.245 54.120 ;
        RECT 115.695 53.430 116.055 54.050 ;
        RECT 115.775 52.550 116.035 53.430 ;
        RECT 116.315 53.180 119.145 54.230 ;
        RECT 115.605 52.170 116.135 52.550 ;
        RECT 110.995 51.910 111.495 52.000 ;
        RECT 110.985 51.180 111.495 51.910 ;
        RECT 111.225 50.180 111.495 51.180 ;
        RECT 112.135 50.930 112.405 51.880 ;
        RECT 112.135 50.780 112.605 50.930 ;
        RECT 112.135 50.100 112.695 50.780 ;
        RECT 112.215 50.090 112.695 50.100 ;
        RECT 111.505 49.560 112.125 49.920 ;
        RECT 111.545 49.030 111.975 49.560 ;
        RECT 110.095 48.610 111.975 49.030 ;
        RECT 112.465 48.900 112.695 50.090 ;
        RECT 111.545 47.740 111.975 48.610 ;
        RECT 112.385 48.300 112.765 48.900 ;
        RECT 109.255 47.000 109.945 47.710 ;
        RECT 111.365 47.380 111.985 47.740 ;
        RECT 111.065 47.000 111.355 47.190 ;
        RECT 109.255 46.560 111.355 47.000 ;
        RECT 109.255 46.540 109.945 46.560 ;
        RECT 111.065 46.320 111.355 46.560 ;
        RECT 111.985 46.930 112.255 47.180 ;
        RECT 112.465 46.930 112.695 48.300 ;
        RECT 115.285 46.950 115.615 51.970 ;
        RECT 116.335 51.960 117.465 53.180 ;
        RECT 118.825 53.160 119.145 53.180 ;
        RECT 111.985 46.820 112.695 46.930 ;
        RECT 115.275 46.900 115.615 46.950 ;
        RECT 116.165 47.720 117.545 51.960 ;
        RECT 111.985 46.510 112.645 46.820 ;
        RECT 111.985 46.340 112.255 46.510 ;
        RECT 115.275 44.940 115.555 46.900 ;
        RECT 116.165 46.860 116.465 47.720 ;
        RECT 117.245 46.860 117.545 47.720 ;
        RECT 118.095 46.860 118.425 51.930 ;
        RECT 117.495 46.320 117.975 46.700 ;
        RECT 117.595 45.700 117.845 46.320 ;
        RECT 117.495 45.100 117.875 45.700 ;
        RECT 20.795 39.650 21.175 40.250 ;
        RECT 20.825 39.030 21.075 39.650 ;
        RECT 20.695 38.650 21.175 39.030 ;
        RECT 20.245 33.420 20.575 38.490 ;
        RECT 21.125 37.630 21.425 38.490 ;
        RECT 22.205 37.630 22.505 38.490 ;
        RECT 23.115 38.450 23.395 40.410 ;
        RECT 26.415 38.840 26.685 39.010 ;
        RECT 26.025 38.530 26.685 38.840 ;
        RECT 21.125 33.390 22.505 37.630 ;
        RECT 23.055 38.400 23.395 38.450 ;
        RECT 25.975 38.420 26.685 38.530 ;
        RECT 19.525 32.170 19.845 32.190 ;
        RECT 21.205 32.170 22.335 33.390 ;
        RECT 23.055 33.380 23.385 38.400 ;
        RECT 25.975 37.050 26.205 38.420 ;
        RECT 26.415 38.170 26.685 38.420 ;
        RECT 27.315 38.790 27.605 39.030 ;
        RECT 28.725 38.790 29.415 38.810 ;
        RECT 27.315 38.350 29.415 38.790 ;
        RECT 27.315 38.160 27.605 38.350 ;
        RECT 26.685 37.610 27.305 37.970 ;
        RECT 28.725 37.640 29.415 38.350 ;
        RECT 25.905 36.450 26.285 37.050 ;
        RECT 26.695 36.740 27.125 37.610 ;
        RECT 25.975 35.260 26.205 36.450 ;
        RECT 26.695 36.320 28.575 36.740 ;
        RECT 26.695 35.790 27.125 36.320 ;
        RECT 26.545 35.430 27.165 35.790 ;
        RECT 25.975 35.250 26.455 35.260 ;
        RECT 25.975 34.570 26.535 35.250 ;
        RECT 26.065 34.420 26.535 34.570 ;
        RECT 26.265 33.470 26.535 34.420 ;
        RECT 27.175 34.170 27.445 35.170 ;
        RECT 27.175 33.440 27.685 34.170 ;
        RECT 27.175 33.350 27.675 33.440 ;
        RECT 22.535 32.800 23.065 33.180 ;
        RECT 19.525 31.120 22.355 32.170 ;
        RECT 22.635 31.920 22.895 32.800 ;
        RECT 22.615 31.300 22.975 31.920 ;
        RECT 27.425 31.230 27.675 33.350 ;
        RECT 19.525 30.210 19.845 31.120 ;
        RECT 21.205 31.110 22.335 31.120 ;
        RECT 23.235 30.830 27.875 31.230 ;
        RECT 27.425 30.550 27.675 30.830 ;
        RECT 19.525 30.150 19.855 30.210 ;
        RECT 19.535 20.220 19.855 30.150 ;
        RECT 20.855 28.900 21.125 30.260 ;
        RECT 21.985 28.900 22.255 30.220 ;
        RECT 27.295 30.120 27.675 30.550 ;
        RECT 27.295 29.610 27.655 30.120 ;
        RECT 20.855 22.210 22.255 28.900 ;
        RECT 20.855 20.210 21.125 22.210 ;
        RECT 21.985 20.170 22.255 22.210 ;
        RECT 27.305 21.770 27.565 29.610 ;
        RECT 27.305 20.220 27.685 21.770 ;
        RECT 19.825 19.560 20.875 19.970 ;
        RECT 22.235 19.570 27.285 19.950 ;
        RECT 19.995 18.280 20.665 19.560 ;
        RECT 19.825 17.600 20.945 18.280 ;
        RECT 23.915 16.790 25.845 19.570 ;
        RECT 23.335 15.940 26.045 16.790 ;
        RECT 27.425 15.400 27.685 20.220 ;
        RECT 26.895 14.670 27.785 15.400 ;
        RECT 28.185 14.810 28.575 36.320 ;
        RECT 28.915 16.840 29.415 37.640 ;
        RECT 31.525 38.490 31.805 40.480 ;
        RECT 34.095 40.410 35.195 41.180 ;
        RECT 42.795 40.460 43.095 42.190 ;
        RECT 32.075 39.650 32.455 40.250 ;
        RECT 32.105 39.030 32.355 39.650 ;
        RECT 31.975 38.650 32.455 39.030 ;
        RECT 31.525 33.420 31.855 38.490 ;
        RECT 32.405 37.630 32.705 38.490 ;
        RECT 33.485 37.630 33.785 38.490 ;
        RECT 34.395 38.450 34.675 40.410 ;
        RECT 37.695 38.840 37.965 39.010 ;
        RECT 37.305 38.530 37.965 38.840 ;
        RECT 32.405 33.390 33.785 37.630 ;
        RECT 34.335 38.400 34.675 38.450 ;
        RECT 37.255 38.420 37.965 38.530 ;
        RECT 30.805 32.170 31.125 32.190 ;
        RECT 32.485 32.170 33.615 33.390 ;
        RECT 34.335 33.380 34.665 38.400 ;
        RECT 37.255 37.050 37.485 38.420 ;
        RECT 37.695 38.170 37.965 38.420 ;
        RECT 38.595 38.790 38.885 39.030 ;
        RECT 40.005 38.790 40.695 38.810 ;
        RECT 38.595 38.350 40.695 38.790 ;
        RECT 38.595 38.160 38.885 38.350 ;
        RECT 37.965 37.610 38.585 37.970 ;
        RECT 40.005 37.640 40.695 38.350 ;
        RECT 37.185 36.450 37.565 37.050 ;
        RECT 37.975 36.740 38.405 37.610 ;
        RECT 37.255 35.260 37.485 36.450 ;
        RECT 37.975 36.320 39.855 36.740 ;
        RECT 37.975 35.790 38.405 36.320 ;
        RECT 37.825 35.430 38.445 35.790 ;
        RECT 37.255 35.250 37.735 35.260 ;
        RECT 37.255 34.570 37.815 35.250 ;
        RECT 37.345 34.420 37.815 34.570 ;
        RECT 37.545 33.470 37.815 34.420 ;
        RECT 38.455 34.170 38.725 35.170 ;
        RECT 38.455 33.440 38.965 34.170 ;
        RECT 38.455 33.350 38.955 33.440 ;
        RECT 33.815 32.800 34.345 33.180 ;
        RECT 30.805 31.120 33.635 32.170 ;
        RECT 33.915 31.920 34.175 32.800 ;
        RECT 33.895 31.300 34.255 31.920 ;
        RECT 38.705 31.230 38.955 33.350 ;
        RECT 30.805 30.210 31.125 31.120 ;
        RECT 32.485 31.110 33.615 31.120 ;
        RECT 34.515 30.830 39.155 31.230 ;
        RECT 38.705 30.550 38.955 30.830 ;
        RECT 30.805 30.150 31.135 30.210 ;
        RECT 30.815 20.220 31.135 30.150 ;
        RECT 32.135 28.900 32.405 30.260 ;
        RECT 33.265 28.900 33.535 30.220 ;
        RECT 38.575 30.120 38.955 30.550 ;
        RECT 38.575 29.610 38.935 30.120 ;
        RECT 32.135 22.210 33.535 28.900 ;
        RECT 32.135 20.210 32.405 22.210 ;
        RECT 33.265 20.170 33.535 22.210 ;
        RECT 38.585 21.770 38.845 29.610 ;
        RECT 38.585 20.220 38.965 21.770 ;
        RECT 31.105 19.560 32.155 19.970 ;
        RECT 33.515 19.570 38.565 19.950 ;
        RECT 31.275 18.280 31.945 19.560 ;
        RECT 31.105 17.600 32.225 18.280 ;
        RECT 28.185 12.290 28.595 14.810 ;
        RECT 28.895 13.610 29.435 16.840 ;
        RECT 35.195 16.790 37.125 19.570 ;
        RECT 34.615 15.940 37.325 16.790 ;
        RECT 38.705 15.400 38.965 20.220 ;
        RECT 38.175 14.670 39.065 15.400 ;
        RECT 39.465 14.810 39.855 36.320 ;
        RECT 40.195 16.840 40.695 37.640 ;
        RECT 42.815 38.470 43.095 40.460 ;
        RECT 45.385 40.390 46.485 41.160 ;
        RECT 54.015 40.460 54.315 42.190 ;
        RECT 43.365 39.630 43.745 40.230 ;
        RECT 43.395 39.010 43.645 39.630 ;
        RECT 43.265 38.630 43.745 39.010 ;
        RECT 42.815 33.400 43.145 38.470 ;
        RECT 43.695 37.610 43.995 38.470 ;
        RECT 44.775 37.610 45.075 38.470 ;
        RECT 45.685 38.430 45.965 40.390 ;
        RECT 48.985 38.820 49.255 38.990 ;
        RECT 48.595 38.510 49.255 38.820 ;
        RECT 43.695 33.370 45.075 37.610 ;
        RECT 45.625 38.380 45.965 38.430 ;
        RECT 48.545 38.400 49.255 38.510 ;
        RECT 42.095 32.150 42.415 32.170 ;
        RECT 43.775 32.150 44.905 33.370 ;
        RECT 45.625 33.360 45.955 38.380 ;
        RECT 48.545 37.030 48.775 38.400 ;
        RECT 48.985 38.150 49.255 38.400 ;
        RECT 49.885 38.770 50.175 39.010 ;
        RECT 51.295 38.770 51.985 38.790 ;
        RECT 49.885 38.330 51.985 38.770 ;
        RECT 49.885 38.140 50.175 38.330 ;
        RECT 49.255 37.590 49.875 37.950 ;
        RECT 51.295 37.620 51.985 38.330 ;
        RECT 48.475 36.430 48.855 37.030 ;
        RECT 49.265 36.720 49.695 37.590 ;
        RECT 48.545 35.240 48.775 36.430 ;
        RECT 49.265 36.300 51.145 36.720 ;
        RECT 49.265 35.770 49.695 36.300 ;
        RECT 49.115 35.410 49.735 35.770 ;
        RECT 48.545 35.230 49.025 35.240 ;
        RECT 48.545 34.550 49.105 35.230 ;
        RECT 48.635 34.400 49.105 34.550 ;
        RECT 48.835 33.450 49.105 34.400 ;
        RECT 49.745 34.150 50.015 35.150 ;
        RECT 49.745 33.420 50.255 34.150 ;
        RECT 49.745 33.330 50.245 33.420 ;
        RECT 45.105 32.780 45.635 33.160 ;
        RECT 42.095 31.100 44.925 32.150 ;
        RECT 45.205 31.900 45.465 32.780 ;
        RECT 45.185 31.280 45.545 31.900 ;
        RECT 49.995 31.210 50.245 33.330 ;
        RECT 42.095 30.190 42.415 31.100 ;
        RECT 43.775 31.090 44.905 31.100 ;
        RECT 45.805 30.810 50.445 31.210 ;
        RECT 49.995 30.530 50.245 30.810 ;
        RECT 42.095 30.130 42.425 30.190 ;
        RECT 42.105 20.200 42.425 30.130 ;
        RECT 43.425 28.880 43.695 30.240 ;
        RECT 44.555 28.880 44.825 30.200 ;
        RECT 49.865 30.100 50.245 30.530 ;
        RECT 49.865 29.590 50.225 30.100 ;
        RECT 43.425 22.190 44.825 28.880 ;
        RECT 43.425 20.190 43.695 22.190 ;
        RECT 44.555 20.150 44.825 22.190 ;
        RECT 49.875 21.750 50.135 29.590 ;
        RECT 49.875 20.200 50.255 21.750 ;
        RECT 42.395 19.540 43.445 19.950 ;
        RECT 44.805 19.550 49.855 19.930 ;
        RECT 42.565 18.260 43.235 19.540 ;
        RECT 42.395 17.580 43.515 18.260 ;
        RECT 28.875 12.770 29.735 13.610 ;
        RECT 28.185 11.950 30.415 12.290 ;
        RECT 39.465 11.990 39.875 14.810 ;
        RECT 40.175 13.610 40.715 16.840 ;
        RECT 46.485 16.770 48.415 19.550 ;
        RECT 45.905 15.920 48.615 16.770 ;
        RECT 49.995 15.380 50.255 20.200 ;
        RECT 49.465 14.650 50.355 15.380 ;
        RECT 50.755 14.790 51.145 36.300 ;
        RECT 51.485 16.820 51.985 37.620 ;
        RECT 54.035 38.470 54.315 40.460 ;
        RECT 56.605 40.390 57.705 41.160 ;
        RECT 65.215 40.460 65.515 42.190 ;
        RECT 76.145 42.180 77.525 42.750 ;
        RECT 83.625 42.570 85.005 43.140 ;
        RECT 87.385 42.200 88.765 42.770 ;
        RECT 94.875 42.580 96.255 43.150 ;
        RECT 106.875 43.140 107.175 44.870 ;
        RECT 114.755 44.170 115.855 44.940 ;
        RECT 118.145 44.870 118.425 46.860 ;
        RECT 120.505 47.710 121.005 68.510 ;
        RECT 121.345 49.030 121.735 70.540 ;
        RECT 122.135 69.950 123.025 70.680 ;
        RECT 132.615 70.040 134.265 70.810 ;
        RECT 122.235 65.130 122.495 69.950 ;
        RECT 123.875 68.560 126.585 69.410 ;
        RECT 124.075 65.780 126.005 68.560 ;
        RECT 128.975 67.070 130.095 67.750 ;
        RECT 129.255 65.790 129.925 67.070 ;
        RECT 122.635 65.400 127.685 65.780 ;
        RECT 129.045 65.380 130.095 65.790 ;
        RECT 132.925 65.180 133.225 70.040 ;
        RECT 137.675 68.690 139.075 69.460 ;
        RECT 138.385 65.740 138.645 68.690 ;
        RECT 149.410 68.420 150.690 69.620 ;
        RECT 149.480 65.810 150.640 68.420 ;
        RECT 133.365 65.380 138.645 65.740 ;
        RECT 122.235 63.580 122.615 65.130 ;
        RECT 122.355 55.740 122.615 63.580 ;
        RECT 127.665 63.140 127.935 65.180 ;
        RECT 128.795 63.140 129.065 65.140 ;
        RECT 127.665 56.450 129.065 63.140 ;
        RECT 122.265 55.230 122.625 55.740 ;
        RECT 122.245 54.800 122.625 55.230 ;
        RECT 127.665 55.130 127.935 56.450 ;
        RECT 128.795 55.090 129.065 56.450 ;
        RECT 130.065 55.200 130.385 65.130 ;
        RECT 132.925 61.010 133.355 65.180 ;
        RECT 138.385 65.150 138.645 65.380 ;
        RECT 138.385 64.770 138.675 65.150 ;
        RECT 130.065 55.140 130.395 55.200 ;
        RECT 133.055 55.190 133.355 61.010 ;
        RECT 122.245 54.520 122.495 54.800 ;
        RECT 122.045 54.120 126.685 54.520 ;
        RECT 127.585 54.230 128.715 54.240 ;
        RECT 130.075 54.230 130.395 55.140 ;
        RECT 138.395 55.080 138.675 64.770 ;
        RECT 149.390 64.610 150.670 65.810 ;
        RECT 122.245 52.000 122.495 54.120 ;
        RECT 126.945 53.430 127.305 54.050 ;
        RECT 127.025 52.550 127.285 53.430 ;
        RECT 127.565 53.180 130.395 54.230 ;
        RECT 126.855 52.170 127.385 52.550 ;
        RECT 122.245 51.910 122.745 52.000 ;
        RECT 122.235 51.180 122.745 51.910 ;
        RECT 122.475 50.180 122.745 51.180 ;
        RECT 123.385 50.930 123.655 51.880 ;
        RECT 123.385 50.780 123.855 50.930 ;
        RECT 123.385 50.100 123.945 50.780 ;
        RECT 123.465 50.090 123.945 50.100 ;
        RECT 122.755 49.560 123.375 49.920 ;
        RECT 122.795 49.030 123.225 49.560 ;
        RECT 121.345 48.610 123.225 49.030 ;
        RECT 123.715 48.900 123.945 50.090 ;
        RECT 122.795 47.740 123.225 48.610 ;
        RECT 123.635 48.300 124.015 48.900 ;
        RECT 120.505 47.000 121.195 47.710 ;
        RECT 122.615 47.380 123.235 47.740 ;
        RECT 122.315 47.000 122.605 47.190 ;
        RECT 120.505 46.560 122.605 47.000 ;
        RECT 120.505 46.540 121.195 46.560 ;
        RECT 122.315 46.320 122.605 46.560 ;
        RECT 123.235 46.930 123.505 47.180 ;
        RECT 123.715 46.930 123.945 48.300 ;
        RECT 126.535 46.950 126.865 51.970 ;
        RECT 127.585 51.960 128.715 53.180 ;
        RECT 130.075 53.160 130.395 53.180 ;
        RECT 123.235 46.820 123.945 46.930 ;
        RECT 126.525 46.900 126.865 46.950 ;
        RECT 127.415 47.720 128.795 51.960 ;
        RECT 123.235 46.510 123.895 46.820 ;
        RECT 123.235 46.340 123.505 46.510 ;
        RECT 126.525 44.940 126.805 46.900 ;
        RECT 127.415 46.860 127.715 47.720 ;
        RECT 128.495 46.860 128.795 47.720 ;
        RECT 129.345 46.860 129.675 51.930 ;
        RECT 128.745 46.320 129.225 46.700 ;
        RECT 128.845 45.700 129.095 46.320 ;
        RECT 128.745 45.100 129.125 45.700 ;
        RECT 118.145 43.140 118.445 44.870 ;
        RECT 126.005 44.170 127.105 44.940 ;
        RECT 129.395 44.870 129.675 46.860 ;
        RECT 129.395 43.140 129.695 44.870 ;
        RECT 98.595 42.220 99.975 42.790 ;
        RECT 106.155 42.570 107.535 43.140 ;
        RECT 109.795 42.260 111.175 42.830 ;
        RECT 117.425 42.570 118.805 43.140 ;
        RECT 121.005 42.280 122.385 42.850 ;
        RECT 128.675 42.570 130.055 43.140 ;
        RECT 54.585 39.630 54.965 40.230 ;
        RECT 54.615 39.010 54.865 39.630 ;
        RECT 54.485 38.630 54.965 39.010 ;
        RECT 54.035 33.400 54.365 38.470 ;
        RECT 54.915 37.610 55.215 38.470 ;
        RECT 55.995 37.610 56.295 38.470 ;
        RECT 56.905 38.430 57.185 40.390 ;
        RECT 60.205 38.820 60.475 38.990 ;
        RECT 59.815 38.510 60.475 38.820 ;
        RECT 54.915 33.370 56.295 37.610 ;
        RECT 56.845 38.380 57.185 38.430 ;
        RECT 59.765 38.400 60.475 38.510 ;
        RECT 53.315 32.150 53.635 32.170 ;
        RECT 54.995 32.150 56.125 33.370 ;
        RECT 56.845 33.360 57.175 38.380 ;
        RECT 59.765 37.030 59.995 38.400 ;
        RECT 60.205 38.150 60.475 38.400 ;
        RECT 61.105 38.770 61.395 39.010 ;
        RECT 62.515 38.770 63.205 38.790 ;
        RECT 61.105 38.330 63.205 38.770 ;
        RECT 61.105 38.140 61.395 38.330 ;
        RECT 60.475 37.590 61.095 37.950 ;
        RECT 62.515 37.620 63.205 38.330 ;
        RECT 59.695 36.430 60.075 37.030 ;
        RECT 60.485 36.720 60.915 37.590 ;
        RECT 59.765 35.240 59.995 36.430 ;
        RECT 60.485 36.300 62.365 36.720 ;
        RECT 60.485 35.770 60.915 36.300 ;
        RECT 60.335 35.410 60.955 35.770 ;
        RECT 59.765 35.230 60.245 35.240 ;
        RECT 59.765 34.550 60.325 35.230 ;
        RECT 59.855 34.400 60.325 34.550 ;
        RECT 60.055 33.450 60.325 34.400 ;
        RECT 60.965 34.150 61.235 35.150 ;
        RECT 60.965 33.420 61.475 34.150 ;
        RECT 60.965 33.330 61.465 33.420 ;
        RECT 56.325 32.780 56.855 33.160 ;
        RECT 53.315 31.100 56.145 32.150 ;
        RECT 56.425 31.900 56.685 32.780 ;
        RECT 56.405 31.280 56.765 31.900 ;
        RECT 61.215 31.210 61.465 33.330 ;
        RECT 53.315 30.190 53.635 31.100 ;
        RECT 54.995 31.090 56.125 31.100 ;
        RECT 57.025 30.810 61.665 31.210 ;
        RECT 61.215 30.530 61.465 30.810 ;
        RECT 53.315 30.130 53.645 30.190 ;
        RECT 53.325 20.200 53.645 30.130 ;
        RECT 54.645 28.880 54.915 30.240 ;
        RECT 55.775 28.880 56.045 30.200 ;
        RECT 61.085 30.100 61.465 30.530 ;
        RECT 61.085 29.590 61.445 30.100 ;
        RECT 54.645 22.190 56.045 28.880 ;
        RECT 54.645 20.190 54.915 22.190 ;
        RECT 55.775 20.150 56.045 22.190 ;
        RECT 61.095 21.750 61.355 29.590 ;
        RECT 61.095 20.200 61.475 21.750 ;
        RECT 53.615 19.540 54.665 19.950 ;
        RECT 56.025 19.550 61.075 19.930 ;
        RECT 53.785 18.260 54.455 19.540 ;
        RECT 53.615 17.580 54.735 18.260 ;
        RECT 40.155 12.770 41.015 13.610 ;
        RECT 50.755 12.170 51.165 14.790 ;
        RECT 51.465 13.590 52.005 16.820 ;
        RECT 57.705 16.770 59.635 19.550 ;
        RECT 57.125 15.920 59.835 16.770 ;
        RECT 61.215 15.380 61.475 20.200 ;
        RECT 60.685 14.650 61.575 15.380 ;
        RECT 61.975 14.790 62.365 36.300 ;
        RECT 62.705 16.820 63.205 37.620 ;
        RECT 65.235 38.470 65.515 40.460 ;
        RECT 67.805 40.390 68.905 41.160 ;
        RECT 76.505 40.450 76.805 42.180 ;
        RECT 65.785 39.630 66.165 40.230 ;
        RECT 65.815 39.010 66.065 39.630 ;
        RECT 65.685 38.630 66.165 39.010 ;
        RECT 65.235 33.400 65.565 38.470 ;
        RECT 66.115 37.610 66.415 38.470 ;
        RECT 67.195 37.610 67.495 38.470 ;
        RECT 68.105 38.430 68.385 40.390 ;
        RECT 71.405 38.820 71.675 38.990 ;
        RECT 71.015 38.510 71.675 38.820 ;
        RECT 66.115 33.370 67.495 37.610 ;
        RECT 68.045 38.380 68.385 38.430 ;
        RECT 70.965 38.400 71.675 38.510 ;
        RECT 64.515 32.150 64.835 32.170 ;
        RECT 66.195 32.150 67.325 33.370 ;
        RECT 68.045 33.360 68.375 38.380 ;
        RECT 70.965 37.030 71.195 38.400 ;
        RECT 71.405 38.150 71.675 38.400 ;
        RECT 72.305 38.770 72.595 39.010 ;
        RECT 73.715 38.770 74.405 38.790 ;
        RECT 72.305 38.330 74.405 38.770 ;
        RECT 72.305 38.140 72.595 38.330 ;
        RECT 71.675 37.590 72.295 37.950 ;
        RECT 73.715 37.620 74.405 38.330 ;
        RECT 70.895 36.430 71.275 37.030 ;
        RECT 71.685 36.720 72.115 37.590 ;
        RECT 70.965 35.240 71.195 36.430 ;
        RECT 71.685 36.300 73.565 36.720 ;
        RECT 71.685 35.770 72.115 36.300 ;
        RECT 71.535 35.410 72.155 35.770 ;
        RECT 70.965 35.230 71.445 35.240 ;
        RECT 70.965 34.550 71.525 35.230 ;
        RECT 71.055 34.400 71.525 34.550 ;
        RECT 71.255 33.450 71.525 34.400 ;
        RECT 72.165 34.150 72.435 35.150 ;
        RECT 72.165 33.420 72.675 34.150 ;
        RECT 72.165 33.330 72.665 33.420 ;
        RECT 67.525 32.780 68.055 33.160 ;
        RECT 64.515 31.100 67.345 32.150 ;
        RECT 67.625 31.900 67.885 32.780 ;
        RECT 67.605 31.280 67.965 31.900 ;
        RECT 72.415 31.210 72.665 33.330 ;
        RECT 64.515 30.190 64.835 31.100 ;
        RECT 66.195 31.090 67.325 31.100 ;
        RECT 68.225 30.810 72.865 31.210 ;
        RECT 72.415 30.530 72.665 30.810 ;
        RECT 64.515 30.130 64.845 30.190 ;
        RECT 64.525 20.200 64.845 30.130 ;
        RECT 65.845 28.880 66.115 30.240 ;
        RECT 66.975 28.880 67.245 30.200 ;
        RECT 72.285 30.100 72.665 30.530 ;
        RECT 72.285 29.590 72.645 30.100 ;
        RECT 65.845 22.190 67.245 28.880 ;
        RECT 65.845 20.190 66.115 22.190 ;
        RECT 66.975 20.150 67.245 22.190 ;
        RECT 72.295 21.750 72.555 29.590 ;
        RECT 72.295 20.200 72.675 21.750 ;
        RECT 64.815 19.540 65.865 19.950 ;
        RECT 67.225 19.550 72.275 19.930 ;
        RECT 64.985 18.260 65.655 19.540 ;
        RECT 64.815 17.580 65.935 18.260 ;
        RECT 51.445 12.750 52.305 13.590 ;
        RECT 27.865 11.130 30.415 11.950 ;
        RECT 28.395 11.090 30.415 11.130 ;
        RECT 39.115 10.980 41.565 11.990 ;
        RECT 50.335 10.970 52.355 12.170 ;
        RECT 61.975 12.160 62.385 14.790 ;
        RECT 62.685 13.590 63.225 16.820 ;
        RECT 68.905 16.770 70.835 19.550 ;
        RECT 68.325 15.920 71.035 16.770 ;
        RECT 72.415 15.380 72.675 20.200 ;
        RECT 71.885 14.650 72.775 15.380 ;
        RECT 73.175 14.790 73.565 36.300 ;
        RECT 73.905 16.820 74.405 37.620 ;
        RECT 76.525 38.460 76.805 40.450 ;
        RECT 79.095 40.380 80.195 41.150 ;
        RECT 87.745 40.470 88.045 42.200 ;
        RECT 77.075 39.620 77.455 40.220 ;
        RECT 77.105 39.000 77.355 39.620 ;
        RECT 76.975 38.620 77.455 39.000 ;
        RECT 76.525 33.390 76.855 38.460 ;
        RECT 77.405 37.600 77.705 38.460 ;
        RECT 78.485 37.600 78.785 38.460 ;
        RECT 79.395 38.420 79.675 40.380 ;
        RECT 82.695 38.810 82.965 38.980 ;
        RECT 82.305 38.500 82.965 38.810 ;
        RECT 77.405 33.360 78.785 37.600 ;
        RECT 79.335 38.370 79.675 38.420 ;
        RECT 82.255 38.390 82.965 38.500 ;
        RECT 75.805 32.140 76.125 32.160 ;
        RECT 77.485 32.140 78.615 33.360 ;
        RECT 79.335 33.350 79.665 38.370 ;
        RECT 82.255 37.020 82.485 38.390 ;
        RECT 82.695 38.140 82.965 38.390 ;
        RECT 83.595 38.760 83.885 39.000 ;
        RECT 85.005 38.760 85.695 38.780 ;
        RECT 83.595 38.320 85.695 38.760 ;
        RECT 83.595 38.130 83.885 38.320 ;
        RECT 82.965 37.580 83.585 37.940 ;
        RECT 85.005 37.610 85.695 38.320 ;
        RECT 82.185 36.420 82.565 37.020 ;
        RECT 82.975 36.710 83.405 37.580 ;
        RECT 82.255 35.230 82.485 36.420 ;
        RECT 82.975 36.290 84.855 36.710 ;
        RECT 82.975 35.760 83.405 36.290 ;
        RECT 82.825 35.400 83.445 35.760 ;
        RECT 82.255 35.220 82.735 35.230 ;
        RECT 82.255 34.540 82.815 35.220 ;
        RECT 82.345 34.390 82.815 34.540 ;
        RECT 82.545 33.440 82.815 34.390 ;
        RECT 83.455 34.140 83.725 35.140 ;
        RECT 83.455 33.410 83.965 34.140 ;
        RECT 83.455 33.320 83.955 33.410 ;
        RECT 78.815 32.770 79.345 33.150 ;
        RECT 75.805 31.090 78.635 32.140 ;
        RECT 78.915 31.890 79.175 32.770 ;
        RECT 78.895 31.270 79.255 31.890 ;
        RECT 83.705 31.200 83.955 33.320 ;
        RECT 75.805 30.180 76.125 31.090 ;
        RECT 77.485 31.080 78.615 31.090 ;
        RECT 79.515 30.800 84.155 31.200 ;
        RECT 83.705 30.520 83.955 30.800 ;
        RECT 75.805 30.120 76.135 30.180 ;
        RECT 75.815 20.190 76.135 30.120 ;
        RECT 77.135 28.870 77.405 30.230 ;
        RECT 78.265 28.870 78.535 30.190 ;
        RECT 83.575 30.090 83.955 30.520 ;
        RECT 83.575 29.580 83.935 30.090 ;
        RECT 77.135 22.180 78.535 28.870 ;
        RECT 77.135 20.180 77.405 22.180 ;
        RECT 78.265 20.140 78.535 22.180 ;
        RECT 83.585 21.740 83.845 29.580 ;
        RECT 83.585 20.190 83.965 21.740 ;
        RECT 76.105 19.530 77.155 19.940 ;
        RECT 78.515 19.540 83.565 19.920 ;
        RECT 76.275 18.250 76.945 19.530 ;
        RECT 76.105 17.570 77.225 18.250 ;
        RECT 62.665 12.750 63.525 13.590 ;
        RECT 73.175 12.190 73.585 14.790 ;
        RECT 73.885 13.590 74.425 16.820 ;
        RECT 80.195 16.760 82.125 19.540 ;
        RECT 79.615 15.910 82.325 16.760 ;
        RECT 83.705 15.370 83.965 20.190 ;
        RECT 83.175 14.640 84.065 15.370 ;
        RECT 84.465 14.780 84.855 36.290 ;
        RECT 85.195 16.810 85.695 37.610 ;
        RECT 87.765 38.480 88.045 40.470 ;
        RECT 90.335 40.400 91.435 41.170 ;
        RECT 98.955 40.490 99.255 42.220 ;
        RECT 88.315 39.640 88.695 40.240 ;
        RECT 88.345 39.020 88.595 39.640 ;
        RECT 88.215 38.640 88.695 39.020 ;
        RECT 87.765 33.410 88.095 38.480 ;
        RECT 88.645 37.620 88.945 38.480 ;
        RECT 89.725 37.620 90.025 38.480 ;
        RECT 90.635 38.440 90.915 40.400 ;
        RECT 93.935 38.830 94.205 39.000 ;
        RECT 93.545 38.520 94.205 38.830 ;
        RECT 88.645 33.380 90.025 37.620 ;
        RECT 90.575 38.390 90.915 38.440 ;
        RECT 93.495 38.410 94.205 38.520 ;
        RECT 87.045 32.160 87.365 32.180 ;
        RECT 88.725 32.160 89.855 33.380 ;
        RECT 90.575 33.370 90.905 38.390 ;
        RECT 93.495 37.040 93.725 38.410 ;
        RECT 93.935 38.160 94.205 38.410 ;
        RECT 94.835 38.780 95.125 39.020 ;
        RECT 96.245 38.780 96.935 38.800 ;
        RECT 94.835 38.340 96.935 38.780 ;
        RECT 94.835 38.150 95.125 38.340 ;
        RECT 94.205 37.600 94.825 37.960 ;
        RECT 96.245 37.630 96.935 38.340 ;
        RECT 93.425 36.440 93.805 37.040 ;
        RECT 94.215 36.730 94.645 37.600 ;
        RECT 93.495 35.250 93.725 36.440 ;
        RECT 94.215 36.310 96.095 36.730 ;
        RECT 94.215 35.780 94.645 36.310 ;
        RECT 94.065 35.420 94.685 35.780 ;
        RECT 93.495 35.240 93.975 35.250 ;
        RECT 93.495 34.560 94.055 35.240 ;
        RECT 93.585 34.410 94.055 34.560 ;
        RECT 93.785 33.460 94.055 34.410 ;
        RECT 94.695 34.160 94.965 35.160 ;
        RECT 94.695 33.430 95.205 34.160 ;
        RECT 94.695 33.340 95.195 33.430 ;
        RECT 90.055 32.790 90.585 33.170 ;
        RECT 87.045 31.110 89.875 32.160 ;
        RECT 90.155 31.910 90.415 32.790 ;
        RECT 90.135 31.290 90.495 31.910 ;
        RECT 94.945 31.220 95.195 33.340 ;
        RECT 87.045 30.200 87.365 31.110 ;
        RECT 88.725 31.100 89.855 31.110 ;
        RECT 90.755 30.820 95.395 31.220 ;
        RECT 94.945 30.540 95.195 30.820 ;
        RECT 87.045 30.140 87.375 30.200 ;
        RECT 87.055 20.210 87.375 30.140 ;
        RECT 88.375 28.890 88.645 30.250 ;
        RECT 89.505 28.890 89.775 30.210 ;
        RECT 94.815 30.110 95.195 30.540 ;
        RECT 94.815 29.600 95.175 30.110 ;
        RECT 88.375 22.200 89.775 28.890 ;
        RECT 88.375 20.200 88.645 22.200 ;
        RECT 89.505 20.160 89.775 22.200 ;
        RECT 94.825 21.760 95.085 29.600 ;
        RECT 94.825 20.210 95.205 21.760 ;
        RECT 87.345 19.550 88.395 19.960 ;
        RECT 89.755 19.560 94.805 19.940 ;
        RECT 87.515 18.270 88.185 19.550 ;
        RECT 87.345 17.590 88.465 18.270 ;
        RECT 73.865 12.750 74.725 13.590 ;
        RECT 61.415 10.960 63.435 12.160 ;
        RECT 72.725 10.990 74.745 12.190 ;
        RECT 84.465 12.180 84.875 14.780 ;
        RECT 85.175 13.580 85.715 16.810 ;
        RECT 91.435 16.780 93.365 19.560 ;
        RECT 90.855 15.930 93.565 16.780 ;
        RECT 94.945 15.390 95.205 20.210 ;
        RECT 94.415 14.660 95.305 15.390 ;
        RECT 95.705 14.800 96.095 36.310 ;
        RECT 96.435 16.830 96.935 37.630 ;
        RECT 98.975 38.500 99.255 40.490 ;
        RECT 101.545 40.420 102.645 41.190 ;
        RECT 110.155 40.530 110.455 42.260 ;
        RECT 99.525 39.660 99.905 40.260 ;
        RECT 99.555 39.040 99.805 39.660 ;
        RECT 99.425 38.660 99.905 39.040 ;
        RECT 98.975 33.430 99.305 38.500 ;
        RECT 99.855 37.640 100.155 38.500 ;
        RECT 100.935 37.640 101.235 38.500 ;
        RECT 101.845 38.460 102.125 40.420 ;
        RECT 105.145 38.850 105.415 39.020 ;
        RECT 104.755 38.540 105.415 38.850 ;
        RECT 99.855 33.400 101.235 37.640 ;
        RECT 101.785 38.410 102.125 38.460 ;
        RECT 104.705 38.430 105.415 38.540 ;
        RECT 98.255 32.180 98.575 32.200 ;
        RECT 99.935 32.180 101.065 33.400 ;
        RECT 101.785 33.390 102.115 38.410 ;
        RECT 104.705 37.060 104.935 38.430 ;
        RECT 105.145 38.180 105.415 38.430 ;
        RECT 106.045 38.800 106.335 39.040 ;
        RECT 107.455 38.800 108.145 38.820 ;
        RECT 106.045 38.360 108.145 38.800 ;
        RECT 106.045 38.170 106.335 38.360 ;
        RECT 105.415 37.620 106.035 37.980 ;
        RECT 107.455 37.650 108.145 38.360 ;
        RECT 104.635 36.460 105.015 37.060 ;
        RECT 105.425 36.750 105.855 37.620 ;
        RECT 104.705 35.270 104.935 36.460 ;
        RECT 105.425 36.330 107.305 36.750 ;
        RECT 105.425 35.800 105.855 36.330 ;
        RECT 105.275 35.440 105.895 35.800 ;
        RECT 104.705 35.260 105.185 35.270 ;
        RECT 104.705 34.580 105.265 35.260 ;
        RECT 104.795 34.430 105.265 34.580 ;
        RECT 104.995 33.480 105.265 34.430 ;
        RECT 105.905 34.180 106.175 35.180 ;
        RECT 105.905 33.450 106.415 34.180 ;
        RECT 105.905 33.360 106.405 33.450 ;
        RECT 101.265 32.810 101.795 33.190 ;
        RECT 98.255 31.130 101.085 32.180 ;
        RECT 101.365 31.930 101.625 32.810 ;
        RECT 101.345 31.310 101.705 31.930 ;
        RECT 106.155 31.240 106.405 33.360 ;
        RECT 98.255 30.220 98.575 31.130 ;
        RECT 99.935 31.120 101.065 31.130 ;
        RECT 101.965 30.840 106.605 31.240 ;
        RECT 106.155 30.560 106.405 30.840 ;
        RECT 98.255 30.160 98.585 30.220 ;
        RECT 98.265 20.230 98.585 30.160 ;
        RECT 99.585 28.910 99.855 30.270 ;
        RECT 100.715 28.910 100.985 30.230 ;
        RECT 106.025 30.130 106.405 30.560 ;
        RECT 106.025 29.620 106.385 30.130 ;
        RECT 99.585 22.220 100.985 28.910 ;
        RECT 99.585 20.220 99.855 22.220 ;
        RECT 100.715 20.180 100.985 22.220 ;
        RECT 106.035 21.780 106.295 29.620 ;
        RECT 106.035 20.230 106.415 21.780 ;
        RECT 98.555 19.570 99.605 19.980 ;
        RECT 100.965 19.580 106.015 19.960 ;
        RECT 98.725 18.290 99.395 19.570 ;
        RECT 98.555 17.610 99.675 18.290 ;
        RECT 85.155 12.740 86.015 13.580 ;
        RECT 95.705 12.180 96.115 14.800 ;
        RECT 96.415 13.600 96.955 16.830 ;
        RECT 102.645 16.800 104.575 19.580 ;
        RECT 102.065 15.950 104.775 16.800 ;
        RECT 106.155 15.410 106.415 20.230 ;
        RECT 105.625 14.680 106.515 15.410 ;
        RECT 106.915 14.820 107.305 36.330 ;
        RECT 107.645 16.850 108.145 37.650 ;
        RECT 110.175 38.540 110.455 40.530 ;
        RECT 112.745 40.460 113.845 41.230 ;
        RECT 121.365 40.550 121.665 42.280 ;
        RECT 142.880 42.020 144.100 43.390 ;
        RECT 110.725 39.700 111.105 40.300 ;
        RECT 110.755 39.080 111.005 39.700 ;
        RECT 110.625 38.700 111.105 39.080 ;
        RECT 110.175 33.470 110.505 38.540 ;
        RECT 111.055 37.680 111.355 38.540 ;
        RECT 112.135 37.680 112.435 38.540 ;
        RECT 113.045 38.500 113.325 40.460 ;
        RECT 116.345 38.890 116.615 39.060 ;
        RECT 115.955 38.580 116.615 38.890 ;
        RECT 111.055 33.440 112.435 37.680 ;
        RECT 112.985 38.450 113.325 38.500 ;
        RECT 115.905 38.470 116.615 38.580 ;
        RECT 109.455 32.220 109.775 32.240 ;
        RECT 111.135 32.220 112.265 33.440 ;
        RECT 112.985 33.430 113.315 38.450 ;
        RECT 115.905 37.100 116.135 38.470 ;
        RECT 116.345 38.220 116.615 38.470 ;
        RECT 117.245 38.840 117.535 39.080 ;
        RECT 118.655 38.840 119.345 38.860 ;
        RECT 117.245 38.400 119.345 38.840 ;
        RECT 117.245 38.210 117.535 38.400 ;
        RECT 116.615 37.660 117.235 38.020 ;
        RECT 118.655 37.690 119.345 38.400 ;
        RECT 115.835 36.500 116.215 37.100 ;
        RECT 116.625 36.790 117.055 37.660 ;
        RECT 115.905 35.310 116.135 36.500 ;
        RECT 116.625 36.370 118.505 36.790 ;
        RECT 116.625 35.840 117.055 36.370 ;
        RECT 116.475 35.480 117.095 35.840 ;
        RECT 115.905 35.300 116.385 35.310 ;
        RECT 115.905 34.620 116.465 35.300 ;
        RECT 115.995 34.470 116.465 34.620 ;
        RECT 116.195 33.520 116.465 34.470 ;
        RECT 117.105 34.220 117.375 35.220 ;
        RECT 117.105 33.490 117.615 34.220 ;
        RECT 117.105 33.400 117.605 33.490 ;
        RECT 112.465 32.850 112.995 33.230 ;
        RECT 109.455 31.170 112.285 32.220 ;
        RECT 112.565 31.970 112.825 32.850 ;
        RECT 112.545 31.350 112.905 31.970 ;
        RECT 117.355 31.280 117.605 33.400 ;
        RECT 109.455 30.260 109.775 31.170 ;
        RECT 111.135 31.160 112.265 31.170 ;
        RECT 113.165 30.880 117.805 31.280 ;
        RECT 117.355 30.600 117.605 30.880 ;
        RECT 109.455 30.200 109.785 30.260 ;
        RECT 109.465 20.270 109.785 30.200 ;
        RECT 110.785 28.950 111.055 30.310 ;
        RECT 111.915 28.950 112.185 30.270 ;
        RECT 117.225 30.170 117.605 30.600 ;
        RECT 117.225 29.660 117.585 30.170 ;
        RECT 110.785 22.260 112.185 28.950 ;
        RECT 110.785 20.260 111.055 22.260 ;
        RECT 111.915 20.220 112.185 22.260 ;
        RECT 117.235 21.820 117.495 29.660 ;
        RECT 117.235 20.270 117.615 21.820 ;
        RECT 109.755 19.610 110.805 20.020 ;
        RECT 112.165 19.620 117.215 20.000 ;
        RECT 109.925 18.330 110.595 19.610 ;
        RECT 109.755 17.650 110.875 18.330 ;
        RECT 96.395 12.760 97.255 13.600 ;
        RECT 106.915 12.230 107.325 14.820 ;
        RECT 107.625 13.620 108.165 16.850 ;
        RECT 113.845 16.840 115.775 19.620 ;
        RECT 113.265 15.990 115.975 16.840 ;
        RECT 117.355 15.450 117.615 20.270 ;
        RECT 116.825 14.720 117.715 15.450 ;
        RECT 118.115 14.860 118.505 36.370 ;
        RECT 118.845 16.890 119.345 37.690 ;
        RECT 121.385 38.560 121.665 40.550 ;
        RECT 123.955 40.480 125.055 41.250 ;
        RECT 121.935 39.720 122.315 40.320 ;
        RECT 121.965 39.100 122.215 39.720 ;
        RECT 121.835 38.720 122.315 39.100 ;
        RECT 121.385 33.490 121.715 38.560 ;
        RECT 122.265 37.700 122.565 38.560 ;
        RECT 123.345 37.700 123.645 38.560 ;
        RECT 124.255 38.520 124.535 40.480 ;
        RECT 127.555 38.910 127.825 39.080 ;
        RECT 127.165 38.600 127.825 38.910 ;
        RECT 122.265 33.460 123.645 37.700 ;
        RECT 124.195 38.470 124.535 38.520 ;
        RECT 127.115 38.490 127.825 38.600 ;
        RECT 120.665 32.240 120.985 32.260 ;
        RECT 122.345 32.240 123.475 33.460 ;
        RECT 124.195 33.450 124.525 38.470 ;
        RECT 127.115 37.120 127.345 38.490 ;
        RECT 127.555 38.240 127.825 38.490 ;
        RECT 128.455 38.860 128.745 39.100 ;
        RECT 142.940 38.950 144.100 42.020 ;
        RECT 129.865 38.860 130.555 38.880 ;
        RECT 128.455 38.420 130.555 38.860 ;
        RECT 128.455 38.230 128.745 38.420 ;
        RECT 127.825 37.680 128.445 38.040 ;
        RECT 129.865 37.710 130.555 38.420 ;
        RECT 127.045 36.520 127.425 37.120 ;
        RECT 127.835 36.810 128.265 37.680 ;
        RECT 127.115 35.330 127.345 36.520 ;
        RECT 127.835 36.390 129.715 36.810 ;
        RECT 127.835 35.860 128.265 36.390 ;
        RECT 127.685 35.500 128.305 35.860 ;
        RECT 127.115 35.320 127.595 35.330 ;
        RECT 127.115 34.640 127.675 35.320 ;
        RECT 127.205 34.490 127.675 34.640 ;
        RECT 127.405 33.540 127.675 34.490 ;
        RECT 128.315 34.240 128.585 35.240 ;
        RECT 128.315 33.510 128.825 34.240 ;
        RECT 128.315 33.420 128.815 33.510 ;
        RECT 123.675 32.870 124.205 33.250 ;
        RECT 120.665 31.190 123.495 32.240 ;
        RECT 123.775 31.990 124.035 32.870 ;
        RECT 123.755 31.370 124.115 31.990 ;
        RECT 128.565 31.300 128.815 33.420 ;
        RECT 120.665 30.280 120.985 31.190 ;
        RECT 122.345 31.180 123.475 31.190 ;
        RECT 124.375 30.900 129.015 31.300 ;
        RECT 128.565 30.620 128.815 30.900 ;
        RECT 120.665 30.220 120.995 30.280 ;
        RECT 120.675 20.290 120.995 30.220 ;
        RECT 121.995 28.970 122.265 30.330 ;
        RECT 123.125 28.970 123.395 30.290 ;
        RECT 128.435 30.190 128.815 30.620 ;
        RECT 128.435 29.680 128.795 30.190 ;
        RECT 121.995 22.280 123.395 28.970 ;
        RECT 121.995 20.280 122.265 22.280 ;
        RECT 123.125 20.240 123.395 22.280 ;
        RECT 128.445 21.840 128.705 29.680 ;
        RECT 128.445 20.290 128.825 21.840 ;
        RECT 120.965 19.630 122.015 20.040 ;
        RECT 123.375 19.640 128.425 20.020 ;
        RECT 121.135 18.350 121.805 19.630 ;
        RECT 120.965 17.670 122.085 18.350 ;
        RECT 107.605 12.780 108.465 13.620 ;
        RECT 118.115 12.230 118.525 14.860 ;
        RECT 118.825 13.660 119.365 16.890 ;
        RECT 125.055 16.860 126.985 19.640 ;
        RECT 124.475 16.010 127.185 16.860 ;
        RECT 128.565 15.470 128.825 20.290 ;
        RECT 128.035 14.740 128.925 15.470 ;
        RECT 129.325 14.880 129.715 36.390 ;
        RECT 130.055 16.910 130.555 37.710 ;
        RECT 142.900 37.580 144.120 38.950 ;
        RECT 132.395 24.340 132.705 30.230 ;
        RECT 132.195 20.120 132.705 24.340 ;
        RECT 118.805 12.820 119.665 13.660 ;
        RECT 129.325 12.260 129.735 14.880 ;
        RECT 130.035 13.680 130.575 16.910 ;
        RECT 132.195 15.510 132.505 20.120 ;
        RECT 137.715 19.980 138.005 30.170 ;
        RECT 132.685 19.590 138.005 19.980 ;
        RECT 137.715 16.940 138.005 19.590 ;
        RECT 142.940 17.940 144.090 19.160 ;
        RECT 145.080 18.760 146.200 18.930 ;
        RECT 137.395 15.890 138.295 16.940 ;
        RECT 137.715 15.720 138.005 15.890 ;
        RECT 131.975 14.270 132.735 15.510 ;
        RECT 142.940 15.090 144.050 17.940 ;
        RECT 142.900 13.870 144.050 15.090 ;
        RECT 145.070 14.920 146.200 18.760 ;
        RECT 145.030 13.970 146.200 14.920 ;
        RECT 145.030 13.900 146.150 13.970 ;
        RECT 130.015 12.840 130.875 13.680 ;
        RECT 83.845 10.980 85.865 12.180 ;
        RECT 95.145 10.980 97.165 12.180 ;
        RECT 106.335 11.030 108.355 12.230 ;
        RECT 117.565 11.030 119.585 12.230 ;
        RECT 128.865 11.060 130.885 12.260 ;
        RECT 74.340 0.110 75.630 1.460 ;
        RECT 93.550 0.180 94.840 1.530 ;
        RECT 112.950 0.310 114.240 1.660 ;
        RECT 131.850 0.380 133.490 1.930 ;
        RECT 151.650 0.250 152.920 1.470 ;
      LAYER met3 ;
        RECT 135.340 223.855 136.790 225.205 ;
        RECT 138.130 223.785 139.580 225.135 ;
        RECT 143.180 223.815 144.630 225.165 ;
        RECT 32.460 203.865 34.440 204.195 ;
        RECT 62.460 203.865 64.440 204.195 ;
        RECT 92.460 203.865 94.440 204.195 ;
        RECT 66.135 203.160 66.465 203.175 ;
        RECT 72.115 203.160 72.445 203.175 ;
        RECT 66.135 202.860 72.445 203.160 ;
        RECT 66.135 202.845 66.465 202.860 ;
        RECT 72.115 202.845 72.445 202.860 ;
        RECT 47.460 201.145 49.440 201.475 ;
        RECT 77.460 201.145 79.440 201.475 ;
        RECT 107.460 201.145 109.440 201.475 ;
        RECT 32.460 198.425 34.440 198.755 ;
        RECT 62.460 198.425 64.440 198.755 ;
        RECT 92.460 198.425 94.440 198.755 ;
        RECT 47.460 195.705 49.440 196.035 ;
        RECT 77.460 195.705 79.440 196.035 ;
        RECT 107.460 195.705 109.440 196.035 ;
        RECT 35.315 195.000 35.645 195.015 ;
        RECT 40.120 195.000 40.500 195.010 ;
        RECT 35.315 194.700 40.500 195.000 ;
        RECT 35.315 194.685 35.645 194.700 ;
        RECT 40.120 194.690 40.500 194.700 ;
        RECT 33.475 194.320 33.805 194.335 ;
        RECT 37.155 194.320 37.485 194.335 ;
        RECT 33.475 194.020 37.485 194.320 ;
        RECT 33.475 194.005 33.805 194.020 ;
        RECT 37.155 194.005 37.485 194.020 ;
        RECT 32.460 192.985 34.440 193.315 ;
        RECT 62.460 192.985 64.440 193.315 ;
        RECT 92.460 192.985 94.440 193.315 ;
        RECT 35.315 190.920 35.645 190.935 ;
        RECT 36.440 190.920 36.820 190.930 ;
        RECT 35.315 190.620 36.820 190.920 ;
        RECT 35.315 190.605 35.645 190.620 ;
        RECT 36.440 190.610 36.820 190.620 ;
        RECT 47.460 190.265 49.440 190.595 ;
        RECT 77.460 190.265 79.440 190.595 ;
        RECT 107.460 190.265 109.440 190.595 ;
        RECT 33.935 189.560 34.265 189.575 ;
        RECT 37.155 189.560 37.485 189.575 ;
        RECT 33.935 189.260 37.485 189.560 ;
        RECT 33.935 189.245 34.265 189.260 ;
        RECT 37.155 189.245 37.485 189.260 ;
        RECT 32.095 188.880 32.425 188.895 ;
        RECT 45.640 188.880 46.020 188.890 ;
        RECT 32.095 188.580 46.020 188.880 ;
        RECT 32.095 188.565 32.425 188.580 ;
        RECT 45.640 188.570 46.020 188.580 ;
        RECT 32.460 187.545 34.440 187.875 ;
        RECT 62.460 187.545 64.440 187.875 ;
        RECT 92.460 187.545 94.440 187.875 ;
        RECT 64.295 186.840 64.625 186.855 ;
        RECT 71.655 186.840 71.985 186.855 ;
        RECT 64.295 186.540 71.985 186.840 ;
        RECT 64.295 186.525 64.625 186.540 ;
        RECT 71.655 186.525 71.985 186.540 ;
        RECT 38.995 185.480 39.325 185.495 ;
        RECT 43.135 185.480 43.465 185.495 ;
        RECT 38.995 185.180 43.465 185.480 ;
        RECT 38.995 185.165 39.325 185.180 ;
        RECT 43.135 185.165 43.465 185.180 ;
        RECT 63.835 185.480 64.165 185.495 ;
        RECT 65.880 185.480 66.260 185.490 ;
        RECT 63.835 185.180 66.260 185.480 ;
        RECT 63.835 185.165 64.165 185.180 ;
        RECT 65.880 185.170 66.260 185.180 ;
        RECT 47.460 184.825 49.440 185.155 ;
        RECT 77.460 184.825 79.440 185.155 ;
        RECT 107.460 184.825 109.440 185.155 ;
        RECT 69.815 183.440 70.145 183.455 ;
        RECT 73.495 183.440 73.825 183.455 ;
        RECT 69.815 183.140 73.825 183.440 ;
        RECT 69.815 183.125 70.145 183.140 ;
        RECT 73.495 183.125 73.825 183.140 ;
        RECT 91.435 183.440 91.765 183.455 ;
        RECT 108.915 183.440 109.245 183.455 ;
        RECT 91.435 183.140 109.245 183.440 ;
        RECT 91.435 183.125 91.765 183.140 ;
        RECT 108.915 183.125 109.245 183.140 ;
        RECT 96.035 182.760 96.365 182.775 ;
        RECT 108.455 182.760 108.785 182.775 ;
        RECT 96.035 182.460 108.785 182.760 ;
        RECT 96.035 182.445 96.365 182.460 ;
        RECT 108.455 182.445 108.785 182.460 ;
        RECT 32.460 182.105 34.440 182.435 ;
        RECT 62.460 182.105 64.440 182.435 ;
        RECT 92.460 182.105 94.440 182.435 ;
        RECT 87.755 181.400 88.085 181.415 ;
        RECT 104.315 181.400 104.645 181.415 ;
        RECT 87.755 181.100 104.645 181.400 ;
        RECT 87.755 181.085 88.085 181.100 ;
        RECT 104.315 181.085 104.645 181.100 ;
        RECT 47.460 179.385 49.440 179.715 ;
        RECT 77.460 179.385 79.440 179.715 ;
        RECT 107.460 179.385 109.440 179.715 ;
        RECT 73.240 177.320 73.620 177.330 ;
        RECT 73.955 177.320 74.285 177.335 ;
        RECT 73.240 177.020 74.285 177.320 ;
        RECT 73.240 177.010 73.620 177.020 ;
        RECT 73.955 177.005 74.285 177.020 ;
        RECT 32.460 176.665 34.440 176.995 ;
        RECT 62.460 176.665 64.440 176.995 ;
        RECT 92.460 176.665 94.440 176.995 ;
        RECT 46.815 175.280 47.145 175.295 ;
        RECT 46.600 174.965 47.145 175.280 ;
        RECT 28.415 173.240 28.745 173.255 ;
        RECT 33.935 173.240 34.265 173.255 ;
        RECT 28.415 172.940 34.265 173.240 ;
        RECT 28.415 172.925 28.745 172.940 ;
        RECT 33.935 172.925 34.265 172.940 ;
        RECT 39.455 173.240 39.785 173.255 ;
        RECT 46.600 173.240 46.900 174.965 ;
        RECT 47.460 173.945 49.440 174.275 ;
        RECT 77.460 173.945 79.440 174.275 ;
        RECT 107.460 173.945 109.440 174.275 ;
        RECT 80.395 173.920 80.725 173.935 ;
        RECT 80.395 173.605 80.940 173.920 ;
        RECT 67.975 173.240 68.305 173.255 ;
        RECT 80.640 173.250 80.940 173.605 ;
        RECT 39.455 172.940 68.305 173.240 ;
        RECT 39.455 172.925 39.785 172.940 ;
        RECT 67.975 172.925 68.305 172.940 ;
        RECT 80.600 173.240 80.980 173.250 ;
        RECT 91.435 173.240 91.765 173.255 ;
        RECT 80.600 172.940 91.765 173.240 ;
        RECT 80.600 172.930 80.980 172.940 ;
        RECT 91.435 172.925 91.765 172.940 ;
        RECT 34.855 172.560 35.185 172.575 ;
        RECT 36.695 172.560 37.025 172.575 ;
        RECT 34.855 172.260 37.025 172.560 ;
        RECT 34.855 172.245 35.185 172.260 ;
        RECT 36.695 172.245 37.025 172.260 ;
        RECT 112.135 172.560 112.465 172.575 ;
        RECT 116.970 172.560 118.970 172.710 ;
        RECT 112.135 172.260 118.970 172.560 ;
        RECT 133.700 172.500 134.930 172.705 ;
        RECT 112.135 172.245 112.465 172.260 ;
        RECT 116.970 172.110 118.970 172.260 ;
        RECT 46.815 171.890 47.145 171.895 ;
        RECT 46.560 171.880 47.145 171.890 ;
        RECT 97.875 171.880 98.205 171.895 ;
        RECT 111.675 171.880 112.005 171.895 ;
        RECT 46.560 171.580 47.370 171.880 ;
        RECT 97.875 171.580 112.005 171.880 ;
        RECT 46.560 171.570 47.145 171.580 ;
        RECT 46.815 171.565 47.145 171.570 ;
        RECT 97.875 171.565 98.205 171.580 ;
        RECT 111.675 171.565 112.005 171.580 ;
        RECT 32.460 171.225 34.440 171.555 ;
        RECT 62.460 171.225 64.440 171.555 ;
        RECT 92.460 171.225 94.440 171.555 ;
        RECT 129.030 170.130 134.930 172.500 ;
        RECT 133.700 170.095 134.930 170.130 ;
        RECT 47.460 168.505 49.440 168.835 ;
        RECT 77.460 168.505 79.440 168.835 ;
        RECT 107.460 168.505 109.440 168.835 ;
        RECT 38.995 167.800 39.325 167.815 ;
        RECT 53.255 167.800 53.585 167.815 ;
        RECT 38.995 167.500 53.585 167.800 ;
        RECT 38.995 167.485 39.325 167.500 ;
        RECT 53.255 167.485 53.585 167.500 ;
        RECT 32.460 165.785 34.440 166.115 ;
        RECT 62.460 165.785 64.440 166.115 ;
        RECT 92.460 165.785 94.440 166.115 ;
        RECT 45.895 165.080 46.225 165.095 ;
        RECT 45.895 164.780 46.900 165.080 ;
        RECT 45.895 164.765 46.225 164.780 ;
        RECT 46.600 164.415 46.900 164.780 ;
        RECT 46.600 164.100 47.145 164.415 ;
        RECT 46.815 164.085 47.145 164.100 ;
        RECT 47.460 163.065 49.440 163.395 ;
        RECT 77.460 163.065 79.440 163.395 ;
        RECT 107.460 163.065 109.440 163.395 ;
        RECT 32.460 160.345 34.440 160.675 ;
        RECT 62.460 160.345 64.440 160.675 ;
        RECT 92.460 160.345 94.440 160.675 ;
        RECT 44.975 160.320 45.305 160.335 ;
        RECT 55.555 160.320 55.885 160.335 ;
        RECT 44.975 160.020 55.885 160.320 ;
        RECT 44.975 160.005 45.305 160.020 ;
        RECT 55.555 160.005 55.885 160.020 ;
        RECT 42.675 159.640 43.005 159.655 ;
        RECT 56.475 159.640 56.805 159.655 ;
        RECT 42.675 159.340 56.805 159.640 ;
        RECT 42.675 159.325 43.005 159.340 ;
        RECT 56.475 159.325 56.805 159.340 ;
        RECT 36.695 158.970 37.025 158.975 ;
        RECT 36.440 158.960 37.025 158.970 ;
        RECT 36.240 158.660 37.025 158.960 ;
        RECT 36.440 158.650 37.025 158.660 ;
        RECT 46.560 158.960 46.940 158.970 ;
        RECT 61.535 158.960 61.865 158.975 ;
        RECT 80.600 158.960 80.980 158.970 ;
        RECT 46.560 158.660 80.980 158.960 ;
        RECT 46.560 158.650 46.940 158.660 ;
        RECT 36.695 158.645 37.025 158.650 ;
        RECT 61.535 158.645 61.865 158.660 ;
        RECT 80.600 158.650 80.980 158.660 ;
        RECT 89.135 158.280 89.465 158.295 ;
        RECT 96.495 158.280 96.825 158.295 ;
        RECT 89.135 157.980 96.825 158.280 ;
        RECT 89.135 157.965 89.465 157.980 ;
        RECT 96.495 157.965 96.825 157.980 ;
        RECT 47.460 157.625 49.440 157.955 ;
        RECT 77.460 157.625 79.440 157.955 ;
        RECT 107.460 157.625 109.440 157.955 ;
        RECT 50.955 157.600 51.285 157.615 ;
        RECT 62.455 157.600 62.785 157.615 ;
        RECT 50.955 157.300 62.785 157.600 ;
        RECT 50.955 157.285 51.285 157.300 ;
        RECT 62.455 157.285 62.785 157.300 ;
        RECT 99.715 156.920 100.045 156.935 ;
        RECT 101.555 156.920 101.885 156.935 ;
        RECT 56.720 156.620 101.885 156.920 ;
        RECT 41.755 156.240 42.085 156.255 ;
        RECT 45.895 156.240 46.225 156.255 ;
        RECT 41.755 155.940 46.225 156.240 ;
        RECT 41.755 155.925 42.085 155.940 ;
        RECT 45.895 155.925 46.225 155.940 ;
        RECT 51.875 156.240 52.205 156.255 ;
        RECT 52.795 156.240 53.125 156.255 ;
        RECT 56.015 156.240 56.345 156.255 ;
        RECT 56.720 156.240 57.020 156.620 ;
        RECT 99.715 156.605 100.045 156.620 ;
        RECT 101.555 156.605 101.885 156.620 ;
        RECT 51.875 155.940 57.020 156.240 ;
        RECT 67.975 156.240 68.305 156.255 ;
        RECT 101.760 156.240 102.140 156.250 ;
        RECT 67.975 155.940 102.140 156.240 ;
        RECT 51.875 155.925 52.205 155.940 ;
        RECT 52.795 155.925 53.125 155.940 ;
        RECT 56.015 155.925 56.345 155.940 ;
        RECT 67.975 155.925 68.305 155.940 ;
        RECT 101.760 155.930 102.140 155.940 ;
        RECT 32.460 154.905 34.440 155.235 ;
        RECT 62.460 154.905 64.440 155.235 ;
        RECT 92.460 154.905 94.440 155.235 ;
        RECT 35.315 154.200 35.645 154.215 ;
        RECT 38.280 154.200 38.660 154.210 ;
        RECT 35.315 153.900 38.660 154.200 ;
        RECT 35.315 153.885 35.645 153.900 ;
        RECT 38.280 153.890 38.660 153.900 ;
        RECT 50.955 154.200 51.285 154.215 ;
        RECT 67.515 154.200 67.845 154.215 ;
        RECT 50.955 153.900 67.845 154.200 ;
        RECT 50.955 153.885 51.285 153.900 ;
        RECT 67.515 153.885 67.845 153.900 ;
        RECT 39.200 153.520 39.580 153.530 ;
        RECT 44.055 153.520 44.385 153.535 ;
        RECT 39.200 153.220 44.385 153.520 ;
        RECT 39.200 153.210 39.580 153.220 ;
        RECT 44.055 153.205 44.385 153.220 ;
        RECT 47.460 152.185 49.440 152.515 ;
        RECT 77.460 152.185 79.440 152.515 ;
        RECT 107.460 152.185 109.440 152.515 ;
        RECT 40.375 152.170 40.705 152.175 ;
        RECT 40.120 152.160 40.705 152.170 ;
        RECT 39.920 151.860 40.705 152.160 ;
        RECT 40.120 151.850 40.705 151.860 ;
        RECT 40.375 151.845 40.705 151.850 ;
        RECT 32.460 149.465 34.440 149.795 ;
        RECT 62.460 149.465 64.440 149.795 ;
        RECT 92.460 149.465 94.440 149.795 ;
        RECT 24.275 148.760 24.605 148.775 ;
        RECT 36.235 148.760 36.565 148.775 ;
        RECT 24.275 148.460 36.565 148.760 ;
        RECT 24.275 148.445 24.605 148.460 ;
        RECT 36.235 148.445 36.565 148.460 ;
        RECT 47.460 146.745 49.440 147.075 ;
        RECT 77.460 146.745 79.440 147.075 ;
        RECT 107.460 146.745 109.440 147.075 ;
        RECT 65.880 146.040 66.260 146.050 ;
        RECT 66.595 146.040 66.925 146.055 ;
        RECT 65.880 145.740 66.925 146.040 ;
        RECT 65.880 145.730 66.260 145.740 ;
        RECT 66.595 145.725 66.925 145.740 ;
        RECT 101.760 145.360 102.140 145.370 ;
        RECT 116.970 145.360 118.970 145.510 ;
        RECT 101.760 145.060 118.970 145.360 ;
        RECT 101.760 145.050 102.140 145.060 ;
        RECT 116.970 144.910 118.970 145.060 ;
        RECT 32.460 144.025 34.440 144.355 ;
        RECT 62.460 144.025 64.440 144.355 ;
        RECT 92.460 144.025 94.440 144.355 ;
        RECT 45.640 143.320 46.020 143.330 ;
        RECT 47.275 143.320 47.605 143.335 ;
        RECT 45.640 143.020 47.605 143.320 ;
        RECT 45.640 143.010 46.020 143.020 ;
        RECT 47.275 143.005 47.605 143.020 ;
        RECT 71.655 142.640 71.985 142.655 ;
        RECT 74.415 142.640 74.745 142.655 ;
        RECT 71.655 142.340 74.745 142.640 ;
        RECT 71.655 142.325 71.985 142.340 ;
        RECT 74.415 142.325 74.745 142.340 ;
        RECT 47.460 141.305 49.440 141.635 ;
        RECT 77.460 141.305 79.440 141.635 ;
        RECT 107.460 141.305 109.440 141.635 ;
        RECT 42.215 140.600 42.545 140.615 ;
        RECT 58.775 140.600 59.105 140.615 ;
        RECT 80.855 140.610 81.185 140.615 ;
        RECT 42.215 140.300 59.105 140.600 ;
        RECT 42.215 140.285 42.545 140.300 ;
        RECT 58.775 140.285 59.105 140.300 ;
        RECT 80.600 140.600 81.185 140.610 ;
        RECT 87.295 140.600 87.625 140.615 ;
        RECT 80.600 140.300 87.625 140.600 ;
        RECT 80.600 140.290 81.185 140.300 ;
        RECT 80.855 140.285 81.185 140.290 ;
        RECT 87.295 140.285 87.625 140.300 ;
        RECT 32.460 138.585 34.440 138.915 ;
        RECT 62.460 138.585 64.440 138.915 ;
        RECT 92.460 138.585 94.440 138.915 ;
        RECT 44.515 138.560 44.845 138.575 ;
        RECT 73.035 138.570 73.365 138.575 ;
        RECT 46.560 138.560 46.940 138.570 ;
        RECT 44.515 138.260 46.940 138.560 ;
        RECT 44.515 138.245 44.845 138.260 ;
        RECT 46.560 138.250 46.940 138.260 ;
        RECT 73.035 138.560 73.620 138.570 ;
        RECT 73.035 138.260 73.820 138.560 ;
        RECT 73.035 138.250 73.620 138.260 ;
        RECT 73.035 138.245 73.365 138.250 ;
        RECT 132.510 138.165 135.210 140.035 ;
        RECT 47.460 135.865 49.440 136.195 ;
        RECT 77.460 135.865 79.440 136.195 ;
        RECT 107.460 135.865 109.440 136.195 ;
        RECT 32.460 133.145 34.440 133.475 ;
        RECT 62.460 133.145 64.440 133.475 ;
        RECT 92.460 133.145 94.440 133.475 ;
        RECT 44.055 131.760 44.385 131.775 ;
        RECT 47.275 131.760 47.605 131.775 ;
        RECT 44.055 131.460 47.605 131.760 ;
        RECT 44.055 131.445 44.385 131.460 ;
        RECT 47.275 131.445 47.605 131.460 ;
        RECT 47.460 130.425 49.440 130.755 ;
        RECT 77.460 130.425 79.440 130.755 ;
        RECT 107.460 130.425 109.440 130.755 ;
        RECT 32.460 127.705 34.440 128.035 ;
        RECT 62.460 127.705 64.440 128.035 ;
        RECT 92.460 127.705 94.440 128.035 ;
        RECT 25.655 127.000 25.985 127.015 ;
        RECT 44.055 127.000 44.385 127.015 ;
        RECT 25.655 126.700 44.385 127.000 ;
        RECT 25.655 126.685 25.985 126.700 ;
        RECT 44.055 126.685 44.385 126.700 ;
        RECT 47.460 124.985 49.440 125.315 ;
        RECT 77.460 124.985 79.440 125.315 ;
        RECT 107.460 124.985 109.440 125.315 ;
        RECT 32.460 122.265 34.440 122.595 ;
        RECT 62.460 122.265 64.440 122.595 ;
        RECT 92.460 122.265 94.440 122.595 ;
        RECT 47.460 119.545 49.440 119.875 ;
        RECT 77.460 119.545 79.440 119.875 ;
        RECT 107.460 119.545 109.440 119.875 ;
        RECT 38.535 118.170 38.865 118.175 ;
        RECT 38.280 118.160 38.865 118.170 ;
        RECT 38.080 117.860 38.865 118.160 ;
        RECT 38.280 117.850 38.865 117.860 ;
        RECT 38.535 117.845 38.865 117.850 ;
        RECT 111.675 118.160 112.005 118.175 ;
        RECT 116.970 118.160 118.970 118.310 ;
        RECT 111.675 117.860 118.970 118.160 ;
        RECT 111.675 117.845 112.005 117.860 ;
        RECT 116.970 117.710 118.970 117.860 ;
        RECT 38.535 117.480 38.865 117.495 ;
        RECT 39.200 117.480 39.580 117.490 ;
        RECT 38.535 117.180 39.580 117.480 ;
        RECT 38.535 117.165 38.865 117.180 ;
        RECT 39.200 117.170 39.580 117.180 ;
        RECT 32.460 116.825 34.440 117.155 ;
        RECT 62.460 116.825 64.440 117.155 ;
        RECT 92.460 116.825 94.440 117.155 ;
        RECT 47.460 114.105 49.440 114.435 ;
        RECT 77.460 114.105 79.440 114.435 ;
        RECT 107.460 114.105 109.440 114.435 ;
        RECT 129.700 105.605 133.210 106.625 ;
        RECT 37.630 88.620 38.970 88.755 ;
        RECT 13.950 87.980 14.980 88.515 ;
        RECT 13.950 87.500 14.990 87.980 ;
        RECT 13.950 87.175 14.980 87.500 ;
        RECT 14.070 86.570 14.810 87.175 ;
        RECT 20.050 87.105 20.920 88.515 ;
        RECT 14.070 75.715 14.700 86.570 ;
        RECT 20.170 77.115 20.800 87.105 ;
        RECT 25.910 87.055 26.860 88.515 ;
        RECT 26.070 78.385 26.700 87.055 ;
        RECT 31.730 86.965 32.910 88.585 ;
        RECT 32.005 79.615 32.635 86.965 ;
        RECT 37.630 86.835 39.120 88.620 ;
        RECT 38.060 81.125 38.690 86.835 ;
        RECT 43.790 86.745 45.190 88.605 ;
        RECT 49.710 86.945 51.060 88.615 ;
        RECT 44.175 82.625 44.805 86.745 ;
        RECT 50.070 83.875 50.700 86.945 ;
        RECT 55.530 86.785 56.750 88.545 ;
        RECT 55.825 85.115 56.455 86.785 ;
        RECT 61.670 86.625 63.180 88.615 ;
        RECT 67.680 88.305 68.720 89.815 ;
        RECT 67.885 87.225 68.515 88.305 ;
        RECT 62.110 86.175 62.740 86.625 ;
        RECT 67.885 86.595 130.605 87.225 ;
        RECT 62.110 85.545 118.855 86.175 ;
        RECT 55.825 84.485 107.605 85.115 ;
        RECT 50.070 83.245 96.285 83.875 ;
        RECT 44.175 81.995 85.055 82.625 ;
        RECT 38.060 80.495 73.765 81.125 ;
        RECT 32.005 78.985 62.635 79.615 ;
        RECT 26.070 77.755 51.245 78.385 ;
        RECT 20.170 76.485 40.645 77.115 ;
        RECT 14.070 75.660 29.295 75.715 ;
        RECT 40.015 75.710 40.645 76.485 ;
        RECT 14.070 75.085 30.410 75.660 ;
        RECT 27.850 74.670 30.410 75.085 ;
        RECT 3.910 71.345 6.100 73.215 ;
        RECT 27.850 73.120 30.450 74.670 ;
        RECT 39.060 74.510 41.620 75.710 ;
        RECT 50.615 75.580 51.245 77.755 ;
        RECT 62.005 75.690 62.635 78.985 ;
        RECT 49.930 74.650 52.490 75.580 ;
        RECT 0.970 70.330 3.070 70.430 ;
        RECT 15.510 70.330 17.040 71.185 ;
        RECT 0.960 68.750 17.040 70.330 ;
        RECT 0.970 68.710 3.070 68.750 ;
        RECT 15.510 68.635 17.040 68.750 ;
        RECT 20.145 54.060 20.605 54.135 ;
        RECT 25.715 54.060 26.175 54.085 ;
        RECT 20.145 53.620 26.175 54.060 ;
        RECT 20.145 53.565 20.605 53.620 ;
        RECT 25.715 53.515 26.175 53.620 ;
        RECT 22.405 48.870 22.885 48.935 ;
        RECT 22.405 48.550 24.205 48.870 ;
        RECT 22.405 48.385 22.885 48.550 ;
        RECT 23.635 45.710 24.195 48.550 ;
        RECT 27.515 45.710 27.995 45.735 ;
        RECT 23.635 45.290 27.995 45.710 ;
        RECT 23.635 45.280 24.195 45.290 ;
        RECT 27.515 45.185 27.995 45.290 ;
        RECT 20.745 40.120 21.225 40.225 ;
        RECT 24.545 40.120 25.105 40.130 ;
        RECT 20.745 39.700 25.105 40.120 ;
        RECT 20.745 39.675 21.225 39.700 ;
        RECT 24.545 36.860 25.105 39.700 ;
        RECT 25.855 36.860 26.335 37.025 ;
        RECT 24.535 36.540 26.335 36.860 ;
        RECT 25.855 36.475 26.335 36.540 ;
        RECT 22.565 31.790 23.025 31.895 ;
        RECT 28.135 31.790 28.595 31.845 ;
        RECT 22.565 31.350 28.595 31.790 ;
        RECT 22.565 31.325 23.025 31.350 ;
        RECT 28.135 31.275 28.595 31.350 ;
        RECT 29.765 12.265 30.255 73.120 ;
        RECT 38.960 73.080 41.730 74.510 ;
        RECT 31.345 54.070 31.805 54.145 ;
        RECT 36.915 54.070 37.375 54.095 ;
        RECT 31.345 53.630 37.375 54.070 ;
        RECT 31.345 53.575 31.805 53.630 ;
        RECT 36.915 53.525 37.375 53.630 ;
        RECT 33.605 48.880 34.085 48.945 ;
        RECT 33.605 48.560 35.405 48.880 ;
        RECT 33.605 48.395 34.085 48.560 ;
        RECT 34.835 45.720 35.395 48.560 ;
        RECT 38.715 45.720 39.195 45.745 ;
        RECT 34.835 45.300 39.195 45.720 ;
        RECT 34.835 45.290 35.395 45.300 ;
        RECT 38.715 45.195 39.195 45.300 ;
        RECT 32.025 40.120 32.505 40.225 ;
        RECT 35.825 40.120 36.385 40.130 ;
        RECT 32.025 39.700 36.385 40.120 ;
        RECT 32.025 39.675 32.505 39.700 ;
        RECT 35.825 36.860 36.385 39.700 ;
        RECT 37.135 36.860 37.615 37.025 ;
        RECT 35.815 36.540 37.615 36.860 ;
        RECT 37.135 36.475 37.615 36.540 ;
        RECT 33.845 31.790 34.305 31.895 ;
        RECT 39.415 31.790 39.875 31.845 ;
        RECT 33.845 31.350 39.875 31.790 ;
        RECT 33.845 31.325 34.305 31.350 ;
        RECT 39.415 31.275 39.875 31.350 ;
        RECT 41.055 12.360 41.545 73.080 ;
        RECT 49.930 73.030 52.530 74.650 ;
        RECT 61.330 74.530 63.890 75.690 ;
        RECT 73.135 75.580 73.765 80.495 ;
        RECT 84.425 75.690 85.055 81.995 ;
        RECT 72.340 74.980 74.900 75.580 ;
        RECT 42.565 54.040 43.025 54.115 ;
        RECT 48.135 54.040 48.595 54.065 ;
        RECT 42.565 53.600 48.595 54.040 ;
        RECT 42.565 53.545 43.025 53.600 ;
        RECT 48.135 53.495 48.595 53.600 ;
        RECT 44.825 48.850 45.305 48.915 ;
        RECT 44.825 48.530 46.625 48.850 ;
        RECT 44.825 48.365 45.305 48.530 ;
        RECT 46.055 45.690 46.615 48.530 ;
        RECT 49.935 45.690 50.415 45.715 ;
        RECT 46.055 45.270 50.415 45.690 ;
        RECT 46.055 45.260 46.615 45.270 ;
        RECT 49.935 45.165 50.415 45.270 ;
        RECT 43.315 40.100 43.795 40.205 ;
        RECT 47.115 40.100 47.675 40.110 ;
        RECT 43.315 39.680 47.675 40.100 ;
        RECT 43.315 39.655 43.795 39.680 ;
        RECT 47.115 36.840 47.675 39.680 ;
        RECT 48.425 36.840 48.905 37.005 ;
        RECT 47.105 36.520 48.905 36.840 ;
        RECT 48.425 36.455 48.905 36.520 ;
        RECT 45.135 31.770 45.595 31.875 ;
        RECT 50.705 31.770 51.165 31.825 ;
        RECT 45.135 31.330 51.165 31.770 ;
        RECT 45.135 31.305 45.595 31.330 ;
        RECT 50.705 31.255 51.165 31.330 ;
        RECT 41.055 12.350 41.555 12.360 ;
        RECT 28.345 11.115 30.465 12.265 ;
        RECT 41.065 11.965 41.555 12.350 ;
        RECT 51.635 12.145 52.125 73.030 ;
        RECT 61.260 73.010 64.060 74.530 ;
        RECT 72.340 73.050 75.020 74.980 ;
        RECT 83.730 74.540 86.290 75.690 ;
        RECT 95.655 75.580 96.285 83.245 ;
        RECT 106.975 75.640 107.605 84.485 ;
        RECT 118.225 75.650 118.855 85.545 ;
        RECT 129.975 75.650 130.605 86.595 ;
        RECT 133.330 76.605 136.060 77.855 ;
        RECT 137.190 76.585 139.920 77.835 ;
        RECT 53.815 54.020 54.275 54.095 ;
        RECT 59.385 54.020 59.845 54.045 ;
        RECT 53.815 53.580 59.845 54.020 ;
        RECT 53.815 53.525 54.275 53.580 ;
        RECT 59.385 53.475 59.845 53.580 ;
        RECT 56.075 48.830 56.555 48.895 ;
        RECT 56.075 48.510 57.875 48.830 ;
        RECT 56.075 48.345 56.555 48.510 ;
        RECT 57.305 45.670 57.865 48.510 ;
        RECT 61.185 45.670 61.665 45.695 ;
        RECT 57.305 45.250 61.665 45.670 ;
        RECT 57.305 45.240 57.865 45.250 ;
        RECT 61.185 45.145 61.665 45.250 ;
        RECT 54.535 40.100 55.015 40.205 ;
        RECT 58.335 40.100 58.895 40.110 ;
        RECT 54.535 39.680 58.895 40.100 ;
        RECT 54.535 39.655 55.015 39.680 ;
        RECT 58.335 36.840 58.895 39.680 ;
        RECT 59.645 36.840 60.125 37.005 ;
        RECT 58.325 36.520 60.125 36.840 ;
        RECT 59.645 36.455 60.125 36.520 ;
        RECT 56.355 31.770 56.815 31.875 ;
        RECT 61.925 31.770 62.385 31.825 ;
        RECT 56.355 31.330 62.385 31.770 ;
        RECT 56.355 31.305 56.815 31.330 ;
        RECT 61.925 31.255 62.385 31.330 ;
        RECT 29.765 11.100 30.255 11.115 ;
        RECT 39.065 11.005 41.615 11.965 ;
        RECT 50.285 10.995 52.405 12.145 ;
        RECT 62.915 12.135 63.405 73.010 ;
        RECT 65.035 54.010 65.495 54.085 ;
        RECT 70.605 54.010 71.065 54.035 ;
        RECT 65.035 53.570 71.065 54.010 ;
        RECT 65.035 53.515 65.495 53.570 ;
        RECT 70.605 53.465 71.065 53.570 ;
        RECT 67.295 48.820 67.775 48.885 ;
        RECT 67.295 48.500 69.095 48.820 ;
        RECT 67.295 48.335 67.775 48.500 ;
        RECT 68.525 45.660 69.085 48.500 ;
        RECT 72.405 45.660 72.885 45.685 ;
        RECT 68.525 45.240 72.885 45.660 ;
        RECT 68.525 45.230 69.085 45.240 ;
        RECT 72.405 45.135 72.885 45.240 ;
        RECT 65.735 40.100 66.215 40.205 ;
        RECT 69.535 40.100 70.095 40.110 ;
        RECT 65.735 39.680 70.095 40.100 ;
        RECT 65.735 39.655 66.215 39.680 ;
        RECT 69.535 36.840 70.095 39.680 ;
        RECT 70.845 36.840 71.325 37.005 ;
        RECT 69.525 36.520 71.325 36.840 ;
        RECT 70.845 36.455 71.325 36.520 ;
        RECT 67.555 31.770 68.015 31.875 ;
        RECT 73.125 31.770 73.585 31.825 ;
        RECT 67.555 31.330 73.585 31.770 ;
        RECT 67.555 31.305 68.015 31.330 ;
        RECT 73.125 31.255 73.585 31.330 ;
        RECT 74.055 12.165 74.545 73.050 ;
        RECT 83.690 73.000 86.290 74.540 ;
        RECT 94.960 74.710 97.520 75.580 ;
        RECT 94.960 73.020 97.570 74.710 ;
        RECT 106.340 74.460 108.900 75.640 ;
        RECT 117.470 74.720 120.030 75.650 ;
        RECT 76.275 54.000 76.735 54.075 ;
        RECT 81.845 54.000 82.305 54.025 ;
        RECT 76.275 53.560 82.305 54.000 ;
        RECT 76.275 53.505 76.735 53.560 ;
        RECT 81.845 53.455 82.305 53.560 ;
        RECT 78.535 48.810 79.015 48.875 ;
        RECT 78.535 48.490 80.335 48.810 ;
        RECT 78.535 48.325 79.015 48.490 ;
        RECT 79.765 45.650 80.325 48.490 ;
        RECT 83.645 45.650 84.125 45.675 ;
        RECT 79.765 45.230 84.125 45.650 ;
        RECT 79.765 45.220 80.325 45.230 ;
        RECT 83.645 45.125 84.125 45.230 ;
        RECT 77.025 40.090 77.505 40.195 ;
        RECT 80.825 40.090 81.385 40.100 ;
        RECT 77.025 39.670 81.385 40.090 ;
        RECT 77.025 39.645 77.505 39.670 ;
        RECT 80.825 36.830 81.385 39.670 ;
        RECT 82.135 36.830 82.615 36.995 ;
        RECT 80.815 36.510 82.615 36.830 ;
        RECT 82.135 36.445 82.615 36.510 ;
        RECT 78.845 31.760 79.305 31.865 ;
        RECT 84.415 31.760 84.875 31.815 ;
        RECT 78.845 31.320 84.875 31.760 ;
        RECT 78.845 31.295 79.305 31.320 ;
        RECT 84.415 31.245 84.875 31.320 ;
        RECT 61.365 10.985 63.485 12.135 ;
        RECT 72.675 11.015 74.795 12.165 ;
        RECT 85.375 12.155 85.865 73.000 ;
        RECT 87.525 54.010 87.985 54.085 ;
        RECT 93.095 54.010 93.555 54.035 ;
        RECT 87.525 53.570 93.555 54.010 ;
        RECT 87.525 53.515 87.985 53.570 ;
        RECT 93.095 53.465 93.555 53.570 ;
        RECT 89.785 48.820 90.265 48.885 ;
        RECT 89.785 48.500 91.585 48.820 ;
        RECT 89.785 48.335 90.265 48.500 ;
        RECT 91.015 45.660 91.575 48.500 ;
        RECT 94.895 45.660 95.375 45.685 ;
        RECT 91.015 45.240 95.375 45.660 ;
        RECT 91.015 45.230 91.575 45.240 ;
        RECT 94.895 45.135 95.375 45.240 ;
        RECT 88.265 40.110 88.745 40.215 ;
        RECT 92.065 40.110 92.625 40.120 ;
        RECT 88.265 39.690 92.625 40.110 ;
        RECT 88.265 39.665 88.745 39.690 ;
        RECT 92.065 36.850 92.625 39.690 ;
        RECT 93.375 36.850 93.855 37.015 ;
        RECT 92.055 36.530 93.855 36.850 ;
        RECT 93.375 36.465 93.855 36.530 ;
        RECT 90.085 31.780 90.545 31.885 ;
        RECT 95.655 31.780 96.115 31.835 ;
        RECT 90.085 31.340 96.115 31.780 ;
        RECT 90.085 31.315 90.545 31.340 ;
        RECT 95.655 31.265 96.115 31.340 ;
        RECT 96.605 12.155 97.095 73.020 ;
        RECT 106.150 73.000 109.060 74.460 ;
        RECT 117.470 73.070 120.000 74.720 ;
        RECT 129.290 74.650 131.850 75.650 ;
        RECT 129.300 73.140 131.820 74.650 ;
        RECT 98.805 54.000 99.265 54.075 ;
        RECT 104.375 54.000 104.835 54.025 ;
        RECT 98.805 53.560 104.835 54.000 ;
        RECT 98.805 53.505 99.265 53.560 ;
        RECT 104.375 53.455 104.835 53.560 ;
        RECT 101.065 48.810 101.545 48.875 ;
        RECT 101.065 48.490 102.865 48.810 ;
        RECT 101.065 48.325 101.545 48.490 ;
        RECT 102.295 45.650 102.855 48.490 ;
        RECT 106.175 45.650 106.655 45.675 ;
        RECT 102.295 45.230 106.655 45.650 ;
        RECT 102.295 45.220 102.855 45.230 ;
        RECT 106.175 45.125 106.655 45.230 ;
        RECT 99.475 40.130 99.955 40.235 ;
        RECT 103.275 40.130 103.835 40.140 ;
        RECT 99.475 39.710 103.835 40.130 ;
        RECT 99.475 39.685 99.955 39.710 ;
        RECT 103.275 36.870 103.835 39.710 ;
        RECT 104.585 36.870 105.065 37.035 ;
        RECT 103.265 36.550 105.065 36.870 ;
        RECT 104.585 36.485 105.065 36.550 ;
        RECT 101.295 31.800 101.755 31.905 ;
        RECT 106.865 31.800 107.325 31.855 ;
        RECT 101.295 31.360 107.325 31.800 ;
        RECT 101.295 31.335 101.755 31.360 ;
        RECT 106.865 31.285 107.325 31.360 ;
        RECT 107.865 12.205 108.355 73.000 ;
        RECT 110.075 54.000 110.535 54.075 ;
        RECT 115.645 54.000 116.105 54.025 ;
        RECT 110.075 53.560 116.105 54.000 ;
        RECT 110.075 53.505 110.535 53.560 ;
        RECT 115.645 53.455 116.105 53.560 ;
        RECT 112.335 48.810 112.815 48.875 ;
        RECT 112.335 48.490 114.135 48.810 ;
        RECT 112.335 48.325 112.815 48.490 ;
        RECT 113.565 45.650 114.125 48.490 ;
        RECT 117.445 45.650 117.925 45.675 ;
        RECT 113.565 45.230 117.925 45.650 ;
        RECT 113.565 45.220 114.125 45.230 ;
        RECT 117.445 45.125 117.925 45.230 ;
        RECT 110.675 40.170 111.155 40.275 ;
        RECT 114.475 40.170 115.035 40.180 ;
        RECT 110.675 39.750 115.035 40.170 ;
        RECT 110.675 39.725 111.155 39.750 ;
        RECT 114.475 36.910 115.035 39.750 ;
        RECT 115.785 36.910 116.265 37.075 ;
        RECT 114.465 36.590 116.265 36.910 ;
        RECT 115.785 36.525 116.265 36.590 ;
        RECT 112.495 31.840 112.955 31.945 ;
        RECT 118.065 31.840 118.525 31.895 ;
        RECT 112.495 31.400 118.525 31.840 ;
        RECT 112.495 31.375 112.955 31.400 ;
        RECT 118.065 31.325 118.525 31.400 ;
        RECT 119.085 12.205 119.575 73.070 ;
        RECT 121.325 54.000 121.785 54.075 ;
        RECT 126.895 54.000 127.355 54.025 ;
        RECT 121.325 53.560 127.355 54.000 ;
        RECT 121.325 53.505 121.785 53.560 ;
        RECT 126.895 53.455 127.355 53.560 ;
        RECT 123.585 48.810 124.065 48.875 ;
        RECT 123.585 48.490 125.385 48.810 ;
        RECT 123.585 48.325 124.065 48.490 ;
        RECT 124.815 45.650 125.375 48.490 ;
        RECT 128.695 45.650 129.175 45.675 ;
        RECT 124.815 45.230 129.175 45.650 ;
        RECT 124.815 45.220 125.375 45.230 ;
        RECT 128.695 45.125 129.175 45.230 ;
        RECT 121.885 40.190 122.365 40.295 ;
        RECT 125.685 40.190 126.245 40.200 ;
        RECT 121.885 39.770 126.245 40.190 ;
        RECT 121.885 39.745 122.365 39.770 ;
        RECT 125.685 36.930 126.245 39.770 ;
        RECT 126.995 36.930 127.475 37.095 ;
        RECT 125.675 36.610 127.475 36.930 ;
        RECT 126.995 36.545 127.475 36.610 ;
        RECT 123.705 31.860 124.165 31.965 ;
        RECT 129.275 31.860 129.735 31.915 ;
        RECT 123.705 31.420 129.735 31.860 ;
        RECT 123.705 31.395 124.165 31.420 ;
        RECT 129.275 31.345 129.735 31.420 ;
        RECT 130.335 12.235 130.825 73.140 ;
        RECT 74.055 11.010 74.545 11.015 ;
        RECT 83.795 11.005 85.915 12.155 ;
        RECT 95.095 11.005 97.215 12.155 ;
        RECT 106.285 11.055 108.405 12.205 ;
        RECT 117.515 11.055 119.635 12.205 ;
        RECT 128.815 11.085 130.935 12.235 ;
        RECT 107.865 11.010 108.355 11.055 ;
        RECT 119.085 11.050 119.575 11.055 ;
        RECT 85.375 11.000 85.865 11.005 ;
        RECT 96.605 10.980 97.095 11.005 ;
        RECT 74.290 0.135 75.680 1.435 ;
        RECT 93.500 0.205 94.890 1.505 ;
        RECT 112.900 0.335 114.290 1.635 ;
        RECT 131.800 0.405 133.540 1.905 ;
        RECT 151.600 0.275 152.970 1.445 ;
      LAYER met4 ;
        RECT 30.420 225.130 30.670 225.140 ;
        RECT 30.300 224.760 30.670 225.130 ;
        RECT 30.970 224.760 33.430 225.140 ;
        RECT 33.730 224.760 36.190 225.140 ;
        RECT 36.490 224.760 38.950 225.140 ;
        RECT 39.250 224.760 41.710 225.140 ;
        RECT 42.010 224.760 44.470 225.140 ;
        RECT 44.770 224.760 47.230 225.140 ;
        RECT 47.530 224.760 49.990 225.140 ;
        RECT 50.290 224.760 52.750 225.140 ;
        RECT 53.050 224.760 55.510 225.140 ;
        RECT 55.810 224.760 58.270 225.140 ;
        RECT 58.570 224.760 61.030 225.140 ;
        RECT 61.330 224.760 63.790 225.140 ;
        RECT 64.090 224.760 66.550 225.140 ;
        RECT 66.850 224.760 69.310 225.140 ;
        RECT 69.610 224.760 72.070 225.140 ;
        RECT 72.370 224.760 74.830 225.140 ;
        RECT 75.130 224.760 77.590 225.140 ;
        RECT 77.890 224.760 80.350 225.140 ;
        RECT 80.650 224.760 83.110 225.140 ;
        RECT 83.410 224.760 85.870 225.140 ;
        RECT 86.170 224.760 88.630 225.140 ;
        RECT 88.930 224.760 91.390 225.140 ;
        RECT 91.690 224.760 94.150 225.140 ;
        RECT 94.450 224.760 96.910 225.140 ;
        RECT 97.210 224.760 99.670 225.140 ;
        RECT 99.970 224.760 102.430 225.140 ;
        RECT 102.730 224.760 105.190 225.140 ;
        RECT 105.490 224.760 107.950 225.140 ;
        RECT 108.250 224.760 110.710 225.140 ;
        RECT 111.010 224.760 113.470 225.140 ;
        RECT 113.770 224.760 116.230 225.140 ;
        RECT 116.530 224.760 118.990 225.140 ;
        RECT 119.290 224.760 121.750 225.140 ;
        RECT 122.050 224.760 124.510 225.140 ;
        RECT 124.810 224.760 127.270 225.140 ;
        RECT 127.570 224.760 130.030 225.140 ;
        RECT 130.330 224.760 132.790 225.140 ;
        RECT 133.090 224.760 133.520 225.140 ;
        RECT 30.300 224.240 133.520 224.760 ;
        RECT 135.385 224.760 135.550 225.185 ;
        RECT 135.850 224.760 136.745 225.185 ;
        RECT 30.300 219.100 31.660 224.240 ;
        RECT 135.385 223.875 136.745 224.760 ;
        RECT 138.175 224.760 138.310 225.115 ;
        RECT 138.610 224.760 139.535 225.115 ;
        RECT 138.175 223.805 139.535 224.760 ;
        RECT 143.225 224.760 143.830 225.145 ;
        RECT 144.130 224.760 144.585 225.145 ;
        RECT 143.225 223.835 144.585 224.760 ;
        RECT 6.000 218.040 31.660 219.100 ;
        RECT 30.300 217.960 31.660 218.040 ;
        RECT 32.450 114.030 34.450 204.270 ;
        RECT 40.145 194.685 40.475 195.015 ;
        RECT 36.465 190.605 36.795 190.935 ;
        RECT 36.480 158.975 36.780 190.605 ;
        RECT 36.465 158.645 36.795 158.975 ;
        RECT 38.305 153.885 38.635 154.215 ;
        RECT 38.320 118.175 38.620 153.885 ;
        RECT 39.225 153.205 39.555 153.535 ;
        RECT 38.305 117.845 38.635 118.175 ;
        RECT 39.240 117.495 39.540 153.205 ;
        RECT 40.160 152.175 40.460 194.685 ;
        RECT 45.665 188.565 45.995 188.895 ;
        RECT 40.145 151.845 40.475 152.175 ;
        RECT 45.680 143.335 45.980 188.565 ;
        RECT 46.585 171.565 46.915 171.895 ;
        RECT 46.600 158.975 46.900 171.565 ;
        RECT 46.585 158.645 46.915 158.975 ;
        RECT 45.665 143.005 45.995 143.335 ;
        RECT 46.600 138.575 46.900 158.645 ;
        RECT 46.585 138.245 46.915 138.575 ;
        RECT 39.225 117.165 39.555 117.495 ;
        RECT 47.450 114.030 49.450 204.270 ;
        RECT 62.450 114.030 64.450 204.270 ;
        RECT 65.905 185.165 66.235 185.495 ;
        RECT 65.920 146.055 66.220 185.165 ;
        RECT 73.265 177.005 73.595 177.335 ;
        RECT 65.905 145.725 66.235 146.055 ;
        RECT 73.280 138.575 73.580 177.005 ;
        RECT 73.265 138.245 73.595 138.575 ;
        RECT 77.450 114.030 79.450 204.270 ;
        RECT 80.625 172.925 80.955 173.255 ;
        RECT 80.640 158.975 80.940 172.925 ;
        RECT 80.625 158.645 80.955 158.975 ;
        RECT 80.640 140.615 80.940 158.645 ;
        RECT 80.625 140.285 80.955 140.615 ;
        RECT 92.450 114.030 94.450 204.270 ;
        RECT 101.785 155.925 102.115 156.255 ;
        RECT 101.800 145.375 102.100 155.925 ;
        RECT 101.785 145.045 102.115 145.375 ;
        RECT 107.450 114.030 109.450 204.270 ;
        RECT 118.110 97.700 120.130 99.670 ;
        RECT 121.810 97.750 123.830 99.720 ;
        RECT 118.130 93.980 120.130 97.700 ;
        RECT 121.820 96.830 123.820 97.750 ;
        RECT 121.820 94.830 139.410 96.830 ;
        RECT 118.130 91.980 135.580 93.980 ;
        RECT 133.580 77.835 135.580 91.980 ;
        RECT 133.375 76.625 136.015 77.835 ;
        RECT 137.410 77.815 139.410 94.830 ;
        RECT 137.235 76.605 139.875 77.815 ;
        RECT 3.955 71.365 4.000 73.195 ;
        RECT 6.000 71.365 6.055 73.195 ;
        RECT 3.000 68.705 3.025 70.435 ;
        RECT 15.555 68.655 16.995 71.165 ;
        RECT 74.335 1.000 75.635 1.415 ;
        RECT 74.335 0.155 74.530 1.000 ;
        RECT 75.430 0.155 75.635 1.000 ;
        RECT 93.545 1.000 94.845 1.485 ;
        RECT 93.545 0.225 93.850 1.000 ;
        RECT 94.750 0.225 94.845 1.000 ;
        RECT 112.945 1.000 114.245 1.615 ;
        RECT 112.945 0.355 113.170 1.000 ;
        RECT 114.070 0.355 114.245 1.000 ;
        RECT 131.845 1.000 133.495 1.885 ;
        RECT 131.845 0.425 132.490 1.000 ;
        RECT 133.390 0.425 133.495 1.000 ;
        RECT 151.645 1.000 152.925 1.425 ;
        RECT 151.645 0.295 151.810 1.000 ;
        RECT 152.710 0.295 152.925 1.000 ;
  END
END tt_um_08_sws
END LIBRARY

